module basic_2500_25000_3000_50_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_1344,In_1745);
nand U1 (N_1,In_665,In_204);
nand U2 (N_2,In_596,In_2326);
nor U3 (N_3,In_1182,In_50);
xor U4 (N_4,In_598,In_1088);
or U5 (N_5,In_733,In_66);
or U6 (N_6,In_1106,In_1181);
nand U7 (N_7,In_1414,In_1719);
xor U8 (N_8,In_2113,In_502);
nor U9 (N_9,In_2086,In_1354);
nand U10 (N_10,In_1062,In_1657);
xnor U11 (N_11,In_977,In_837);
nand U12 (N_12,In_1534,In_2203);
xor U13 (N_13,In_376,In_1495);
xor U14 (N_14,In_1353,In_2374);
nor U15 (N_15,In_526,In_258);
nor U16 (N_16,In_2115,In_708);
nor U17 (N_17,In_1685,In_2061);
and U18 (N_18,In_992,In_1468);
nand U19 (N_19,In_692,In_390);
xor U20 (N_20,In_1663,In_2010);
nand U21 (N_21,In_1336,In_2148);
nor U22 (N_22,In_874,In_2153);
nand U23 (N_23,In_1377,In_1989);
or U24 (N_24,In_1319,In_2121);
or U25 (N_25,In_111,In_2058);
xor U26 (N_26,In_1008,In_2275);
nand U27 (N_27,In_736,In_1011);
and U28 (N_28,In_673,In_2371);
and U29 (N_29,In_2319,In_2361);
xnor U30 (N_30,In_532,In_75);
or U31 (N_31,In_215,In_1476);
or U32 (N_32,In_1981,In_1766);
or U33 (N_33,In_651,In_1574);
nand U34 (N_34,In_1725,In_1120);
nor U35 (N_35,In_712,In_264);
xor U36 (N_36,In_779,In_1603);
xor U37 (N_37,In_2088,In_2483);
xnor U38 (N_38,In_2256,In_122);
nand U39 (N_39,In_450,In_1091);
and U40 (N_40,In_261,In_1598);
or U41 (N_41,In_2313,In_1596);
xnor U42 (N_42,In_420,In_179);
xnor U43 (N_43,In_1112,In_1847);
xor U44 (N_44,In_897,In_1591);
and U45 (N_45,In_1801,In_1142);
nor U46 (N_46,In_1231,In_57);
nand U47 (N_47,In_43,In_2026);
or U48 (N_48,In_2266,In_769);
and U49 (N_49,In_302,In_395);
nand U50 (N_50,In_2224,In_2478);
nor U51 (N_51,In_1079,In_1892);
nand U52 (N_52,In_340,In_842);
nand U53 (N_53,In_2355,In_1520);
nand U54 (N_54,In_167,In_1310);
xor U55 (N_55,In_448,In_1679);
nor U56 (N_56,In_1540,In_2427);
nor U57 (N_57,In_377,In_875);
or U58 (N_58,In_1964,In_1479);
nor U59 (N_59,In_949,In_455);
and U60 (N_60,In_1589,In_2401);
xnor U61 (N_61,In_2166,In_2068);
or U62 (N_62,In_1423,In_1125);
nor U63 (N_63,In_2450,In_431);
and U64 (N_64,In_1727,In_937);
xnor U65 (N_65,In_705,In_2381);
or U66 (N_66,In_1483,In_808);
and U67 (N_67,In_1699,In_476);
nand U68 (N_68,In_1929,In_506);
nand U69 (N_69,In_2336,In_1060);
or U70 (N_70,In_373,In_2150);
and U71 (N_71,In_558,In_2073);
xor U72 (N_72,In_2156,In_946);
and U73 (N_73,In_24,In_2155);
nor U74 (N_74,In_953,In_1938);
nor U75 (N_75,In_1641,In_2340);
xnor U76 (N_76,In_109,In_2395);
nand U77 (N_77,In_499,In_934);
nand U78 (N_78,In_656,In_2096);
xor U79 (N_79,In_1921,In_324);
and U80 (N_80,In_312,In_905);
nand U81 (N_81,In_2105,In_1782);
xor U82 (N_82,In_2403,In_18);
or U83 (N_83,In_758,In_473);
nor U84 (N_84,In_2257,In_1979);
xnor U85 (N_85,In_1849,In_467);
nor U86 (N_86,In_1119,In_828);
nand U87 (N_87,In_17,In_387);
nor U88 (N_88,In_1568,In_393);
xnor U89 (N_89,In_216,In_784);
and U90 (N_90,In_1058,In_670);
or U91 (N_91,In_2376,In_1232);
and U92 (N_92,In_1105,In_2345);
nor U93 (N_93,In_238,In_1269);
and U94 (N_94,In_418,In_2463);
and U95 (N_95,In_1444,In_1493);
nor U96 (N_96,In_1016,In_576);
xnor U97 (N_97,In_68,In_161);
nor U98 (N_98,In_855,In_2335);
xnor U99 (N_99,In_273,In_1285);
nand U100 (N_100,In_2382,In_2302);
nand U101 (N_101,In_1917,In_2173);
xor U102 (N_102,In_1180,In_2200);
or U103 (N_103,In_1013,In_359);
xor U104 (N_104,In_422,In_945);
and U105 (N_105,In_990,In_1029);
xnor U106 (N_106,In_1653,In_1683);
nand U107 (N_107,In_1823,In_2069);
or U108 (N_108,In_2139,In_1099);
xor U109 (N_109,In_1150,In_1368);
and U110 (N_110,In_592,In_2269);
nand U111 (N_111,In_1398,In_1096);
nor U112 (N_112,In_1910,In_1742);
nor U113 (N_113,In_2220,In_1951);
xor U114 (N_114,In_2074,In_1983);
xnor U115 (N_115,In_1006,In_48);
and U116 (N_116,In_972,In_2038);
or U117 (N_117,In_589,In_1484);
and U118 (N_118,In_405,In_2186);
nand U119 (N_119,In_906,In_162);
and U120 (N_120,In_1010,In_727);
or U121 (N_121,In_921,In_1654);
or U122 (N_122,In_1889,In_768);
nor U123 (N_123,In_236,In_1404);
nor U124 (N_124,In_1138,In_1928);
nand U125 (N_125,In_2480,In_1051);
xnor U126 (N_126,In_1824,In_351);
xor U127 (N_127,In_739,In_2177);
or U128 (N_128,In_2067,In_345);
nor U129 (N_129,In_2090,In_1140);
or U130 (N_130,In_1937,In_299);
nor U131 (N_131,In_1372,In_757);
nand U132 (N_132,In_1092,In_1521);
or U133 (N_133,In_110,In_2431);
and U134 (N_134,In_1048,In_2218);
and U135 (N_135,In_1785,In_267);
nor U136 (N_136,In_1316,In_2352);
nor U137 (N_137,In_646,In_1570);
or U138 (N_138,In_1959,In_1973);
nor U139 (N_139,In_879,In_285);
and U140 (N_140,In_1244,In_1557);
nand U141 (N_141,In_1763,In_1332);
and U142 (N_142,In_1798,In_1815);
and U143 (N_143,In_1582,In_1385);
xor U144 (N_144,In_2097,In_979);
xnor U145 (N_145,In_1390,In_525);
nor U146 (N_146,In_1518,In_1754);
nor U147 (N_147,In_569,In_771);
and U148 (N_148,In_791,In_831);
or U149 (N_149,In_2454,In_271);
or U150 (N_150,In_1831,In_691);
xnor U151 (N_151,In_631,In_363);
and U152 (N_152,In_2064,In_1159);
nor U153 (N_153,In_2466,In_1696);
xnor U154 (N_154,In_427,In_1834);
nor U155 (N_155,In_696,In_1194);
xor U156 (N_156,In_1173,In_827);
nor U157 (N_157,In_1408,In_1121);
xor U158 (N_158,In_871,In_2042);
nand U159 (N_159,In_1756,In_263);
or U160 (N_160,In_1562,In_257);
and U161 (N_161,In_2461,In_2223);
xor U162 (N_162,In_2031,In_2495);
or U163 (N_163,In_1475,In_279);
xor U164 (N_164,In_918,In_195);
nor U165 (N_165,In_1774,In_2240);
nor U166 (N_166,In_1949,In_588);
xor U167 (N_167,In_1104,In_862);
xnor U168 (N_168,In_1729,In_25);
xnor U169 (N_169,In_78,In_517);
nand U170 (N_170,In_2037,In_688);
nand U171 (N_171,In_1758,In_1552);
or U172 (N_172,In_711,In_136);
nor U173 (N_173,In_1649,In_821);
nor U174 (N_174,In_986,In_382);
nand U175 (N_175,In_1465,In_2125);
nor U176 (N_176,In_1531,In_1623);
nor U177 (N_177,In_516,In_1790);
or U178 (N_178,In_1097,In_510);
and U179 (N_179,In_1076,In_2481);
and U180 (N_180,In_1075,In_907);
nand U181 (N_181,In_2285,In_1481);
nand U182 (N_182,In_1057,In_1571);
xor U183 (N_183,In_737,In_1644);
and U184 (N_184,In_1590,In_2228);
or U185 (N_185,In_323,In_2050);
nand U186 (N_186,In_1210,In_2255);
xnor U187 (N_187,In_1965,In_2410);
and U188 (N_188,In_1219,In_1373);
xor U189 (N_189,In_184,In_1100);
nor U190 (N_190,In_2063,In_106);
or U191 (N_191,In_1433,In_529);
or U192 (N_192,In_647,In_2017);
nand U193 (N_193,In_2124,In_1019);
and U194 (N_194,In_1186,In_775);
nor U195 (N_195,In_1869,In_1982);
and U196 (N_196,In_1975,In_45);
or U197 (N_197,In_507,In_1734);
nand U198 (N_198,In_2099,In_2062);
nor U199 (N_199,In_409,In_1205);
xor U200 (N_200,In_2225,In_960);
nor U201 (N_201,In_649,In_1496);
nor U202 (N_202,In_930,In_1530);
xnor U203 (N_203,In_2211,In_1887);
nor U204 (N_204,In_1751,In_2066);
nor U205 (N_205,In_441,In_1328);
or U206 (N_206,In_146,In_346);
or U207 (N_207,In_2023,In_668);
nand U208 (N_208,In_817,In_7);
and U209 (N_209,In_1208,In_1897);
or U210 (N_210,In_911,In_535);
or U211 (N_211,In_1512,In_1948);
xor U212 (N_212,In_1884,In_1477);
xnor U213 (N_213,In_604,In_1737);
and U214 (N_214,In_745,In_443);
or U215 (N_215,In_880,In_851);
nor U216 (N_216,In_79,In_732);
xnor U217 (N_217,In_339,In_483);
xor U218 (N_218,In_2411,In_1626);
xor U219 (N_219,In_1797,In_2264);
nor U220 (N_220,In_962,In_1893);
and U221 (N_221,In_710,In_504);
and U222 (N_222,In_2405,In_70);
xor U223 (N_223,In_428,In_1473);
nand U224 (N_224,In_1126,In_2191);
nor U225 (N_225,In_259,In_335);
or U226 (N_226,In_243,In_546);
nand U227 (N_227,In_298,In_1559);
xor U228 (N_228,In_1409,In_1262);
and U229 (N_229,In_534,In_1399);
or U230 (N_230,In_281,In_1561);
or U231 (N_231,In_618,In_750);
nand U232 (N_232,In_421,In_495);
xnor U233 (N_233,In_154,In_2241);
xnor U234 (N_234,In_1978,In_2112);
and U235 (N_235,In_1753,In_2323);
and U236 (N_236,In_1837,In_1001);
and U237 (N_237,In_1579,In_1922);
or U238 (N_238,In_307,In_1564);
nand U239 (N_239,In_1544,In_494);
xor U240 (N_240,In_1972,In_35);
xor U241 (N_241,In_2318,In_1320);
nand U242 (N_242,In_2044,In_498);
and U243 (N_243,In_2303,In_414);
nor U244 (N_244,In_802,In_2270);
and U245 (N_245,In_951,In_1800);
and U246 (N_246,In_1063,In_438);
xnor U247 (N_247,In_2389,In_2151);
or U248 (N_248,In_1430,In_910);
or U249 (N_249,In_1609,In_58);
or U250 (N_250,In_658,In_703);
nor U251 (N_251,In_1918,In_689);
and U252 (N_252,In_2475,In_1786);
and U253 (N_253,In_1375,In_352);
nand U254 (N_254,In_160,In_927);
and U255 (N_255,In_1502,In_2346);
nand U256 (N_256,In_2100,In_356);
or U257 (N_257,In_465,In_103);
xnor U258 (N_258,In_2485,In_1253);
and U259 (N_259,In_1688,In_1898);
xor U260 (N_260,In_1391,In_379);
nand U261 (N_261,In_2499,In_1308);
nor U262 (N_262,In_280,In_997);
and U263 (N_263,In_454,In_843);
and U264 (N_264,In_1883,In_412);
nor U265 (N_265,In_2360,In_2444);
nand U266 (N_266,In_636,In_1233);
xor U267 (N_267,In_2307,In_860);
nand U268 (N_268,In_321,In_330);
xor U269 (N_269,In_1791,In_1736);
nand U270 (N_270,In_1067,In_436);
xnor U271 (N_271,In_980,In_679);
and U272 (N_272,In_1290,In_1056);
nand U273 (N_273,In_478,In_1600);
or U274 (N_274,In_2157,In_49);
or U275 (N_275,In_2231,In_983);
and U276 (N_276,In_2060,In_714);
or U277 (N_277,In_1131,In_1643);
nor U278 (N_278,In_1053,In_1558);
or U279 (N_279,In_1000,In_2261);
nand U280 (N_280,In_1289,In_994);
nand U281 (N_281,In_524,In_1764);
nand U282 (N_282,In_845,In_1850);
nand U283 (N_283,In_1616,In_555);
nor U284 (N_284,In_2474,In_1367);
nand U285 (N_285,In_2337,In_97);
and U286 (N_286,In_1470,In_786);
xnor U287 (N_287,In_552,In_630);
nand U288 (N_288,In_1662,In_2443);
or U289 (N_289,In_410,In_1129);
nand U290 (N_290,In_965,In_1912);
nor U291 (N_291,In_2242,In_777);
nand U292 (N_292,In_2043,In_2030);
xnor U293 (N_293,In_1878,In_1627);
nor U294 (N_294,In_9,In_2363);
nor U295 (N_295,In_1828,In_2415);
nor U296 (N_296,In_1821,In_1953);
nand U297 (N_297,In_766,In_664);
xor U298 (N_298,In_984,In_1740);
nor U299 (N_299,In_2021,In_2406);
nor U300 (N_300,In_1235,In_633);
nor U301 (N_301,In_1342,In_1457);
or U302 (N_302,In_1845,In_2182);
and U303 (N_303,In_252,In_1154);
and U304 (N_304,In_1410,In_759);
nand U305 (N_305,In_396,In_2322);
or U306 (N_306,In_42,In_276);
nand U307 (N_307,In_1136,In_1757);
xor U308 (N_308,In_1384,In_2198);
or U309 (N_309,In_539,In_1400);
nor U310 (N_310,In_672,In_1829);
and U311 (N_311,In_1322,In_1901);
nand U312 (N_312,In_2297,In_156);
and U313 (N_313,In_1765,In_847);
or U314 (N_314,In_437,In_2294);
nor U315 (N_315,In_1888,In_2487);
nor U316 (N_316,In_164,In_1613);
xnor U317 (N_317,In_1324,In_2333);
nand U318 (N_318,In_1188,In_2174);
or U319 (N_319,In_2358,In_2082);
and U320 (N_320,In_1031,In_765);
nor U321 (N_321,In_2271,In_364);
or U322 (N_322,In_270,In_1292);
or U323 (N_323,In_1639,In_5);
xnor U324 (N_324,In_2210,In_2019);
and U325 (N_325,In_151,In_1164);
xor U326 (N_326,In_76,In_1669);
or U327 (N_327,In_288,In_433);
nand U328 (N_328,In_2018,In_697);
nand U329 (N_329,In_2227,In_2047);
and U330 (N_330,In_1442,In_744);
and U331 (N_331,In_1606,In_2491);
nor U332 (N_332,In_1361,In_1365);
xnor U333 (N_333,In_1346,In_1748);
or U334 (N_334,In_1418,In_929);
and U335 (N_335,In_145,In_477);
and U336 (N_336,In_296,In_1246);
and U337 (N_337,In_1134,In_2014);
nor U338 (N_338,In_1345,In_1515);
nand U339 (N_339,In_1799,In_310);
or U340 (N_340,In_370,In_917);
and U341 (N_341,In_123,In_969);
or U342 (N_342,In_882,In_2117);
xor U343 (N_343,In_1924,In_1396);
or U344 (N_344,In_2440,In_1684);
xor U345 (N_345,In_121,In_367);
and U346 (N_346,In_2445,In_1083);
xnor U347 (N_347,In_1718,In_0);
nand U348 (N_348,In_234,In_1155);
or U349 (N_349,In_585,In_832);
xor U350 (N_350,In_1456,In_822);
and U351 (N_351,In_233,In_1624);
or U352 (N_352,In_398,In_1601);
or U353 (N_353,In_401,In_834);
and U354 (N_354,In_676,In_2001);
nor U355 (N_355,In_27,In_559);
xnor U356 (N_356,In_93,In_466);
xor U357 (N_357,In_575,In_1507);
xor U358 (N_358,In_1498,In_2029);
or U359 (N_359,In_1403,In_1066);
and U360 (N_360,In_683,In_583);
nor U361 (N_361,In_2392,In_255);
xor U362 (N_362,In_2237,In_2416);
xnor U363 (N_363,In_2190,In_211);
xor U364 (N_364,In_1673,In_1840);
and U365 (N_365,In_26,In_1438);
and U366 (N_366,In_286,In_1871);
nand U367 (N_367,In_1145,In_1296);
xnor U368 (N_368,In_870,In_248);
nand U369 (N_369,In_556,In_2448);
nand U370 (N_370,In_1023,In_1424);
and U371 (N_371,In_2250,In_157);
nor U372 (N_372,In_536,In_397);
and U373 (N_373,In_2343,In_251);
or U374 (N_374,In_1334,In_138);
and U375 (N_375,In_915,In_701);
nand U376 (N_376,In_2288,In_2245);
nor U377 (N_377,In_1036,In_1731);
xor U378 (N_378,In_1958,In_2140);
nand U379 (N_379,In_2170,In_2161);
nor U380 (N_380,In_1693,In_1304);
xnor U381 (N_381,In_1819,In_747);
xor U382 (N_382,In_1274,In_133);
nor U383 (N_383,In_1044,In_1387);
nand U384 (N_384,In_615,In_1419);
nor U385 (N_385,In_804,In_2193);
and U386 (N_386,In_1264,In_2202);
or U387 (N_387,In_338,In_2330);
xor U388 (N_388,In_381,In_1439);
or U389 (N_389,In_877,In_89);
and U390 (N_390,In_36,In_496);
nand U391 (N_391,In_643,In_434);
xnor U392 (N_392,In_197,In_3);
xor U393 (N_393,In_571,In_1116);
xor U394 (N_394,In_1027,In_640);
and U395 (N_395,In_277,In_1998);
xor U396 (N_396,In_1771,In_957);
nand U397 (N_397,In_933,In_181);
xor U398 (N_398,In_1221,In_2012);
and U399 (N_399,In_456,In_511);
or U400 (N_400,In_54,In_998);
nor U401 (N_401,In_723,In_449);
or U402 (N_402,In_223,In_378);
or U403 (N_403,In_725,In_2159);
and U404 (N_404,In_196,In_1061);
and U405 (N_405,In_287,In_970);
or U406 (N_406,In_1697,In_704);
and U407 (N_407,In_1478,In_662);
xor U408 (N_408,In_2379,In_480);
or U409 (N_409,In_2489,In_1923);
or U410 (N_410,In_789,In_1014);
nand U411 (N_411,In_1077,In_1687);
nor U412 (N_412,In_1415,In_1497);
or U413 (N_413,In_900,In_2111);
or U414 (N_414,In_1886,In_582);
nand U415 (N_415,In_848,In_2424);
xor U416 (N_416,In_1943,In_2065);
xor U417 (N_417,In_2192,In_172);
nor U418 (N_418,In_141,In_394);
nor U419 (N_419,In_2274,In_886);
nor U420 (N_420,In_746,In_1040);
nor U421 (N_421,In_2409,In_654);
nand U422 (N_422,In_1032,In_1178);
nor U423 (N_423,In_635,In_220);
nor U424 (N_424,In_1947,In_663);
or U425 (N_425,In_2135,In_366);
nor U426 (N_426,In_788,In_1789);
xnor U427 (N_427,In_1711,In_611);
or U428 (N_428,In_203,In_2441);
nor U429 (N_429,In_185,In_648);
and U430 (N_430,In_432,In_1576);
nand U431 (N_431,In_1117,In_2116);
and U432 (N_432,In_652,In_690);
xor U433 (N_433,In_451,In_2078);
nand U434 (N_434,In_319,In_721);
xor U435 (N_435,In_369,In_1747);
xnor U436 (N_436,In_1976,In_2071);
and U437 (N_437,In_2311,In_2365);
or U438 (N_438,In_815,In_792);
nor U439 (N_439,In_1371,In_1197);
nand U440 (N_440,In_318,In_372);
nor U441 (N_441,In_1065,In_481);
nor U442 (N_442,In_1146,In_985);
nor U443 (N_443,In_260,In_230);
and U444 (N_444,In_320,In_1523);
and U445 (N_445,In_538,In_1681);
or U446 (N_446,In_1509,In_1635);
or U447 (N_447,In_256,In_1665);
nor U448 (N_448,In_638,In_317);
xnor U449 (N_449,In_1677,In_1604);
and U450 (N_450,In_1352,In_1565);
nand U451 (N_451,In_2434,In_1803);
xor U452 (N_452,In_1670,In_1511);
nand U453 (N_453,In_1247,In_13);
or U454 (N_454,In_1584,In_482);
and U455 (N_455,In_623,In_2467);
or U456 (N_456,In_2306,In_2331);
nand U457 (N_457,In_599,In_1967);
or U458 (N_458,In_1311,In_1239);
and U459 (N_459,In_1055,In_1386);
nand U460 (N_460,In_134,In_284);
and U461 (N_461,In_1229,In_40);
nand U462 (N_462,In_2027,In_245);
and U463 (N_463,In_1554,In_1876);
nand U464 (N_464,In_1816,In_149);
nand U465 (N_465,In_681,In_961);
nand U466 (N_466,In_2470,In_1303);
or U467 (N_467,In_1744,In_2070);
or U468 (N_468,In_1012,In_439);
xor U469 (N_469,In_981,In_1148);
or U470 (N_470,In_2497,In_628);
nor U471 (N_471,In_1022,In_1128);
and U472 (N_472,In_894,In_2232);
nor U473 (N_473,In_227,In_1524);
xnor U474 (N_474,In_1842,In_383);
xnor U475 (N_475,In_531,In_892);
or U476 (N_476,In_1865,In_1914);
nand U477 (N_477,In_1339,In_1426);
xnor U478 (N_478,In_2305,In_2171);
and U479 (N_479,In_752,In_1660);
and U480 (N_480,In_2457,In_950);
nor U481 (N_481,In_952,In_447);
nor U482 (N_482,In_978,In_490);
or U483 (N_483,In_1421,In_1179);
nor U484 (N_484,In_1638,In_1784);
and U485 (N_485,In_1795,In_1629);
nand U486 (N_486,In_1152,In_1450);
or U487 (N_487,In_2048,In_987);
xor U488 (N_488,In_2423,In_2498);
nor U489 (N_489,In_485,In_2299);
xor U490 (N_490,In_1500,In_799);
or U491 (N_491,In_1489,In_472);
xnor U492 (N_492,In_1935,In_1156);
and U493 (N_493,In_99,In_1714);
or U494 (N_494,In_316,In_1370);
nor U495 (N_495,In_812,In_2278);
nand U496 (N_496,In_2196,In_520);
nor U497 (N_497,In_2176,In_642);
nand U498 (N_498,In_2430,In_170);
or U499 (N_499,In_116,In_2054);
nand U500 (N_500,N_301,N_229);
nand U501 (N_501,In_1005,In_1196);
xor U502 (N_502,In_2222,In_290);
xor U503 (N_503,In_717,In_809);
xor U504 (N_504,N_329,N_350);
xnor U505 (N_505,N_53,N_209);
nand U506 (N_506,In_1223,In_976);
or U507 (N_507,In_1172,N_470);
xnor U508 (N_508,N_175,In_1811);
or U509 (N_509,In_2393,In_947);
and U510 (N_510,In_1504,In_1255);
and U511 (N_511,In_1864,In_350);
xnor U512 (N_512,In_2298,N_174);
nor U513 (N_513,N_187,In_1260);
xor U514 (N_514,In_1856,In_813);
and U515 (N_515,In_1505,In_308);
or U516 (N_516,In_2032,In_565);
nor U517 (N_517,N_132,In_1773);
or U518 (N_518,N_87,In_1043);
nor U519 (N_519,N_447,In_332);
nand U520 (N_520,In_2258,In_1338);
nand U521 (N_521,In_2239,In_1350);
and U522 (N_522,In_2229,N_114);
or U523 (N_523,In_459,In_1162);
and U524 (N_524,In_314,In_574);
and U525 (N_525,In_2059,In_702);
nor U526 (N_526,In_1204,N_69);
nand U527 (N_527,In_250,In_2328);
and U528 (N_528,In_371,N_88);
nand U529 (N_529,N_497,N_208);
nor U530 (N_530,In_795,In_1648);
and U531 (N_531,N_319,In_1118);
xor U532 (N_532,In_2281,In_2077);
or U533 (N_533,In_1427,In_1143);
nor U534 (N_534,In_174,In_657);
or U535 (N_535,N_281,In_1161);
or U536 (N_536,In_2132,N_346);
nor U537 (N_537,In_2468,In_2180);
nand U538 (N_538,In_2169,In_1533);
or U539 (N_539,In_1492,In_1009);
or U540 (N_540,In_1678,In_1177);
xor U541 (N_541,In_674,In_2428);
nor U542 (N_542,In_844,In_2272);
nand U543 (N_543,In_1335,N_372);
nor U544 (N_544,In_186,In_2041);
and U545 (N_545,In_1356,In_853);
and U546 (N_546,In_1202,In_1380);
xnor U547 (N_547,N_476,In_1054);
nor U548 (N_548,In_699,In_41);
and U549 (N_549,N_60,In_218);
nand U550 (N_550,N_177,In_2126);
nor U551 (N_551,In_1163,In_1211);
and U552 (N_552,In_1611,In_1389);
nand U553 (N_553,In_169,In_1990);
nand U554 (N_554,In_1904,In_1675);
or U555 (N_555,N_58,In_1899);
or U556 (N_556,In_1425,N_420);
or U557 (N_557,N_324,In_139);
and U558 (N_558,In_2486,In_1360);
and U559 (N_559,In_2183,In_32);
or U560 (N_560,N_273,In_1588);
xnor U561 (N_561,In_861,In_358);
nor U562 (N_562,N_486,In_1090);
nand U563 (N_563,In_1169,N_295);
or U564 (N_564,In_967,In_1318);
xor U565 (N_565,In_1157,In_543);
or U566 (N_566,In_988,In_1170);
xor U567 (N_567,N_272,In_413);
nand U568 (N_568,In_1358,In_713);
or U569 (N_569,N_115,In_706);
nor U570 (N_570,In_1215,In_2436);
xor U571 (N_571,In_2081,In_2265);
nor U572 (N_572,N_164,In_242);
nand U573 (N_573,In_964,In_2315);
xor U574 (N_574,N_376,N_413);
nor U575 (N_575,In_1295,In_2439);
nand U576 (N_576,In_2349,In_2215);
or U577 (N_577,N_439,In_1254);
and U578 (N_578,N_392,In_2102);
nand U579 (N_579,In_1885,In_866);
and U580 (N_580,N_330,In_1905);
xor U581 (N_581,In_1710,N_354);
nand U582 (N_582,In_353,In_724);
and U583 (N_583,N_154,In_1988);
xnor U584 (N_584,N_391,In_2429);
nand U585 (N_585,In_707,In_199);
or U586 (N_586,In_2205,In_587);
nand U587 (N_587,In_1862,In_1977);
or U588 (N_588,N_336,In_1966);
or U589 (N_589,In_1226,In_1741);
nor U590 (N_590,In_523,N_304);
and U591 (N_591,In_1720,In_948);
nor U592 (N_592,N_121,In_39);
and U593 (N_593,In_2332,In_1151);
nor U594 (N_594,N_448,In_1694);
xnor U595 (N_595,In_1567,In_2413);
xnor U596 (N_596,In_194,In_1218);
or U597 (N_597,In_118,N_370);
nand U598 (N_598,In_144,In_904);
nand U599 (N_599,In_1950,In_1622);
or U600 (N_600,In_105,In_1187);
xor U601 (N_601,In_2249,In_695);
xnor U602 (N_602,In_1250,In_1854);
nor U603 (N_603,N_279,In_2284);
nor U604 (N_604,In_142,In_899);
or U605 (N_605,In_2089,In_59);
xor U606 (N_606,In_720,N_463);
nor U607 (N_607,In_1717,N_394);
or U608 (N_608,In_168,In_1343);
or U609 (N_609,In_584,N_130);
nand U610 (N_610,In_1776,In_2207);
xnor U611 (N_611,In_1702,In_2267);
nand U612 (N_612,N_479,N_134);
nor U613 (N_613,In_1522,In_1402);
nor U614 (N_614,In_1249,In_1686);
and U615 (N_615,In_2455,In_60);
nor U616 (N_616,In_709,In_856);
xnor U617 (N_617,In_2053,N_126);
or U618 (N_618,In_954,In_2394);
and U619 (N_619,In_1602,In_1631);
and U620 (N_620,In_1406,N_80);
or U621 (N_621,N_477,In_1275);
nand U622 (N_622,In_1276,In_820);
or U623 (N_623,N_180,In_2402);
xor U624 (N_624,In_2252,In_2149);
nor U625 (N_625,N_458,In_1108);
or U626 (N_626,N_117,N_485);
xor U627 (N_627,In_561,N_438);
xor U628 (N_628,In_1192,In_1111);
or U629 (N_629,In_268,N_79);
and U630 (N_630,In_1499,In_924);
nor U631 (N_631,In_2260,In_1762);
nand U632 (N_632,In_2471,In_1149);
and U633 (N_633,N_75,N_160);
nor U634 (N_634,In_1999,In_1647);
xor U635 (N_635,In_513,N_430);
nor U636 (N_636,In_165,In_206);
nor U637 (N_637,In_1927,In_1288);
or U638 (N_638,In_1549,In_1732);
or U639 (N_639,N_323,In_601);
xnor U640 (N_640,N_298,In_148);
or U641 (N_641,In_249,N_63);
nor U642 (N_642,In_751,In_389);
xnor U643 (N_643,N_242,In_1394);
nand U644 (N_644,In_841,In_254);
nand U645 (N_645,In_463,In_1462);
or U646 (N_646,N_99,In_124);
or U647 (N_647,In_269,In_1759);
and U648 (N_648,In_1769,In_1167);
nand U649 (N_649,In_2391,In_1881);
xnor U650 (N_650,N_373,In_1395);
xnor U651 (N_651,In_1168,N_116);
and U652 (N_652,N_406,N_37);
or U653 (N_653,In_272,N_148);
nand U654 (N_654,In_1230,N_265);
nor U655 (N_655,In_1366,N_19);
nor U656 (N_656,In_794,N_153);
or U657 (N_657,In_1671,In_549);
and U658 (N_658,In_632,In_2128);
xor U659 (N_659,N_136,In_1228);
and U660 (N_660,In_1746,In_1995);
nand U661 (N_661,In_1294,In_850);
and U662 (N_662,In_620,In_991);
nor U663 (N_663,N_400,In_854);
or U664 (N_664,In_1033,In_1775);
nand U665 (N_665,In_2219,In_542);
nor U666 (N_666,In_1102,In_527);
nor U667 (N_667,N_493,In_1130);
nand U668 (N_668,In_487,N_149);
xor U669 (N_669,In_1362,N_290);
nand U670 (N_670,In_639,In_1213);
nor U671 (N_671,In_226,In_283);
nor U672 (N_672,In_1018,N_364);
and U673 (N_673,In_1047,N_328);
and U674 (N_674,In_1546,In_442);
nor U675 (N_675,In_544,In_112);
nor U676 (N_676,In_790,N_473);
and U677 (N_677,In_1293,In_1580);
nand U678 (N_678,In_1449,N_291);
and U679 (N_679,In_2329,In_859);
nand U680 (N_680,In_1448,In_593);
xnor U681 (N_681,In_2387,N_47);
or U682 (N_682,In_64,In_2129);
xnor U683 (N_683,In_85,In_1628);
nand U684 (N_684,In_1214,In_1004);
and U685 (N_685,In_440,In_728);
and U686 (N_686,N_286,In_147);
xnor U687 (N_687,In_572,In_1039);
or U688 (N_688,In_1658,In_1974);
or U689 (N_689,In_129,N_197);
nor U690 (N_690,N_288,In_2462);
xnor U691 (N_691,In_1454,In_908);
nand U692 (N_692,N_12,In_92);
or U693 (N_693,In_1987,N_239);
xor U694 (N_694,In_1024,N_292);
xnor U695 (N_695,N_256,In_2259);
xnor U696 (N_696,In_1607,In_1195);
nand U697 (N_697,In_935,In_1050);
nor U698 (N_698,In_1068,In_2251);
and U699 (N_699,In_1132,In_1997);
xor U700 (N_700,In_1139,N_305);
or U701 (N_701,N_166,In_1946);
nor U702 (N_702,N_122,In_2055);
xnor U703 (N_703,In_407,In_417);
nor U704 (N_704,In_876,N_244);
nand U705 (N_705,In_2312,N_332);
and U706 (N_706,In_2277,In_1642);
xnor U707 (N_707,N_15,In_2452);
or U708 (N_708,In_491,In_2046);
and U709 (N_709,N_310,In_1525);
xor U710 (N_710,In_1932,N_235);
or U711 (N_711,In_852,N_409);
and U712 (N_712,In_301,N_358);
nor U713 (N_713,N_216,In_2408);
xor U714 (N_714,In_1123,In_989);
and U715 (N_715,In_1312,In_2039);
nor U716 (N_716,In_1550,In_1980);
nor U717 (N_717,In_1733,In_1364);
nor U718 (N_718,In_2377,In_1695);
nor U719 (N_719,In_2446,In_2137);
nor U720 (N_720,In_1225,N_386);
and U721 (N_721,In_1257,N_210);
xnor U722 (N_722,In_77,N_200);
nor U723 (N_723,N_314,In_1431);
and U724 (N_724,N_431,In_1158);
and U725 (N_725,N_128,In_362);
and U726 (N_726,In_846,N_383);
xnor U727 (N_727,N_64,In_1783);
nand U728 (N_728,In_1843,In_6);
nand U729 (N_729,In_767,In_2496);
or U730 (N_730,In_388,In_903);
and U731 (N_731,In_738,In_873);
nand U732 (N_732,In_2092,In_1379);
nand U733 (N_733,In_1761,In_675);
or U734 (N_734,N_139,In_1827);
nand U735 (N_735,In_16,In_224);
and U736 (N_736,In_1605,N_155);
and U737 (N_737,In_188,In_926);
or U738 (N_738,N_365,In_435);
nand U739 (N_739,In_1532,In_2179);
xor U740 (N_740,N_107,In_1703);
nand U741 (N_741,In_98,N_313);
nor U742 (N_742,In_1902,In_1237);
and U743 (N_743,N_33,N_20);
nor U744 (N_744,In_578,In_1970);
xor U745 (N_745,In_209,In_1689);
nand U746 (N_746,In_1378,N_261);
xor U747 (N_747,N_196,N_315);
nor U748 (N_748,In_1894,In_2316);
nand U749 (N_749,In_2147,In_132);
xnor U750 (N_750,N_59,In_501);
nand U751 (N_751,In_2106,N_102);
and U752 (N_752,N_73,N_232);
and U753 (N_753,In_883,In_1556);
nand U754 (N_754,N_480,In_1859);
xnor U755 (N_755,In_923,In_1519);
nand U756 (N_756,In_564,In_1382);
nor U757 (N_757,In_1787,N_201);
nand U758 (N_758,In_2033,N_49);
nor U759 (N_759,In_1428,N_389);
xor U760 (N_760,In_1420,N_41);
nor U761 (N_761,In_801,In_415);
or U762 (N_762,N_90,N_226);
and U763 (N_763,In_1818,In_2453);
xor U764 (N_764,In_614,In_1185);
xor U765 (N_765,In_213,In_2123);
nand U766 (N_766,In_1236,In_2287);
or U767 (N_767,In_1529,N_255);
and U768 (N_768,In_1916,In_1326);
and U769 (N_769,N_396,In_334);
and U770 (N_770,In_641,In_1739);
nor U771 (N_771,In_1724,N_35);
or U772 (N_772,In_475,N_455);
and U773 (N_773,N_260,In_514);
or U774 (N_774,N_417,In_219);
nor U775 (N_775,In_1712,In_627);
and U776 (N_776,In_1650,In_1279);
or U777 (N_777,In_1730,In_617);
nor U778 (N_778,In_2372,N_67);
xnor U779 (N_779,In_610,In_1224);
nor U780 (N_780,In_2145,In_1625);
nor U781 (N_781,In_1251,In_687);
nor U782 (N_782,In_865,In_1915);
xnor U783 (N_783,In_143,In_1432);
and U784 (N_784,In_1592,In_31);
or U785 (N_785,In_2273,N_459);
nand U786 (N_786,In_1141,In_1879);
nor U787 (N_787,In_1903,In_1282);
or U788 (N_788,In_2080,In_857);
nand U789 (N_789,In_1698,In_936);
nand U790 (N_790,In_1986,In_266);
and U791 (N_791,N_95,In_889);
or U792 (N_792,In_1513,In_1944);
or U793 (N_793,In_1302,N_92);
nor U794 (N_794,N_26,N_297);
nand U795 (N_795,In_1474,In_430);
and U796 (N_796,In_1548,In_2473);
and U797 (N_797,In_22,In_2233);
and U798 (N_798,N_56,In_2178);
nand U799 (N_799,In_1463,In_1472);
nand U800 (N_800,In_1572,N_380);
nand U801 (N_801,N_425,In_1715);
xnor U802 (N_802,In_956,N_393);
nor U803 (N_803,In_15,In_303);
nand U804 (N_804,In_2398,In_295);
or U805 (N_805,In_1137,In_1283);
nand U806 (N_806,In_2189,N_264);
xor U807 (N_807,In_1212,N_2);
nor U808 (N_808,In_2008,In_505);
nand U809 (N_809,N_247,In_1781);
or U810 (N_810,In_38,In_2327);
and U811 (N_811,N_198,In_225);
nand U812 (N_812,In_399,In_560);
xor U813 (N_813,In_2040,In_1306);
nand U814 (N_814,In_2093,In_931);
nand U815 (N_815,N_320,In_380);
xnor U816 (N_816,N_408,In_562);
xor U817 (N_817,In_315,In_2028);
xor U818 (N_818,In_595,In_971);
nand U819 (N_819,In_1094,N_252);
or U820 (N_820,In_1086,In_840);
nor U821 (N_821,In_1256,In_2276);
or U822 (N_822,In_1802,In_2253);
xor U823 (N_823,In_29,N_460);
and U824 (N_824,N_169,In_1655);
nand U825 (N_825,In_1794,In_1103);
or U826 (N_826,In_2268,In_300);
xor U827 (N_827,In_1777,In_619);
or U828 (N_828,In_2289,In_2020);
nor U829 (N_829,In_1193,In_1124);
nor U830 (N_830,N_483,In_2366);
and U831 (N_831,In_624,In_1002);
and U832 (N_832,In_999,In_368);
or U833 (N_833,N_140,In_881);
nor U834 (N_834,In_830,In_1416);
xor U835 (N_835,In_609,In_56);
nand U836 (N_836,N_474,In_2005);
xor U837 (N_837,In_357,In_152);
nand U838 (N_838,N_398,In_1298);
and U839 (N_839,N_374,N_259);
xor U840 (N_840,N_97,N_105);
nor U841 (N_841,In_667,N_111);
or U842 (N_842,N_275,In_741);
and U843 (N_843,N_211,In_2442);
nor U844 (N_844,In_868,In_1183);
nor U845 (N_845,N_206,In_1440);
nand U846 (N_846,In_2130,In_2417);
or U847 (N_847,N_326,In_1708);
nand U848 (N_848,In_1330,In_1436);
nand U849 (N_849,In_2296,In_2479);
and U850 (N_850,In_2321,N_327);
xor U851 (N_851,In_155,In_192);
or U852 (N_852,In_30,In_1098);
and U853 (N_853,In_175,In_644);
nor U854 (N_854,In_411,N_359);
and U855 (N_855,N_465,N_9);
xor U856 (N_856,In_120,In_84);
nand U857 (N_857,In_1206,In_2286);
and U858 (N_858,In_1107,In_1199);
nand U859 (N_859,In_849,In_202);
nand U860 (N_860,In_778,In_416);
xnor U861 (N_861,In_1664,N_48);
xor U862 (N_862,In_1836,In_1184);
xnor U863 (N_863,In_1459,N_404);
xor U864 (N_864,In_753,N_270);
or U865 (N_865,In_1429,In_1017);
or U866 (N_866,In_829,In_1052);
xor U867 (N_867,N_171,In_1401);
and U868 (N_868,In_887,In_21);
nor U869 (N_869,In_1956,In_354);
nand U870 (N_870,In_2195,In_682);
nor U871 (N_871,In_1369,In_580);
nor U872 (N_872,In_404,In_1070);
nand U873 (N_873,N_258,In_94);
and U874 (N_874,In_774,In_1991);
xnor U875 (N_875,In_1144,In_1855);
nand U876 (N_876,In_2465,In_1443);
nand U877 (N_877,N_31,In_2072);
or U878 (N_878,N_311,In_1963);
nand U879 (N_879,In_2188,In_756);
nor U880 (N_880,In_1833,N_189);
and U881 (N_881,N_11,In_1176);
or U882 (N_882,In_2244,In_1268);
and U883 (N_883,In_2133,In_1860);
and U884 (N_884,N_250,In_512);
xnor U885 (N_885,In_2464,In_760);
nor U886 (N_886,In_453,In_214);
and U887 (N_887,In_2280,In_304);
or U888 (N_888,In_1543,In_2007);
and U889 (N_889,N_101,N_257);
nor U890 (N_890,In_783,In_782);
or U891 (N_891,N_195,In_2025);
nor U892 (N_892,In_2246,In_1553);
nand U893 (N_893,In_1960,In_2375);
or U894 (N_894,In_244,In_1704);
nand U895 (N_895,N_113,In_107);
nand U896 (N_896,N_168,In_91);
or U897 (N_897,N_362,N_86);
xor U898 (N_898,In_1939,N_45);
or U899 (N_899,In_787,N_462);
and U900 (N_900,In_1277,N_55);
nor U901 (N_901,N_451,In_1314);
and U902 (N_902,In_1486,In_591);
nand U903 (N_903,In_1516,In_2045);
or U904 (N_904,In_1174,N_6);
nand U905 (N_905,In_2370,In_1807);
nand U906 (N_906,In_1779,In_551);
or U907 (N_907,In_1363,N_468);
nand U908 (N_908,In_1612,In_1207);
or U909 (N_909,In_2127,In_292);
or U910 (N_910,In_912,In_1541);
nand U911 (N_911,In_1397,In_548);
nand U912 (N_912,In_1810,In_1417);
xor U913 (N_913,In_541,In_1911);
and U914 (N_914,In_1874,N_340);
nor U915 (N_915,N_494,In_2396);
nand U916 (N_916,In_963,In_291);
xor U917 (N_917,In_385,In_348);
nor U918 (N_918,In_2304,In_52);
xor U919 (N_919,In_1615,In_622);
or U920 (N_920,In_1585,N_384);
xor U921 (N_921,In_1349,In_522);
and U922 (N_922,In_835,N_93);
or U923 (N_923,N_23,In_158);
nor U924 (N_924,In_1931,N_156);
nor U925 (N_925,In_313,In_570);
nand U926 (N_926,In_102,N_82);
xor U927 (N_927,N_410,In_1587);
or U928 (N_928,In_2079,N_120);
nor U929 (N_929,In_1166,In_361);
nor U930 (N_930,In_173,In_2262);
nor U931 (N_931,N_124,In_247);
and U932 (N_932,In_1287,In_336);
or U933 (N_933,In_72,In_761);
xor U934 (N_934,In_625,N_317);
xor U935 (N_935,In_1909,In_1517);
xnor U936 (N_936,In_1337,In_1064);
nand U937 (N_937,In_2407,In_1659);
nor U938 (N_938,In_1645,In_208);
and U939 (N_939,In_468,In_1305);
nor U940 (N_940,In_888,In_1266);
nor U941 (N_941,N_492,In_974);
nor U942 (N_942,N_366,In_1248);
nand U943 (N_943,In_53,In_530);
and U944 (N_944,N_3,In_2087);
and U945 (N_945,In_518,In_1652);
or U946 (N_946,In_62,In_1113);
and U947 (N_947,In_1617,In_1954);
nor U948 (N_948,In_515,In_995);
nand U949 (N_949,In_1820,N_377);
xor U950 (N_950,In_1460,N_495);
and U951 (N_951,In_1962,In_1480);
or U952 (N_952,In_1081,N_98);
or U953 (N_953,In_329,In_1806);
nand U954 (N_954,N_233,N_21);
and U955 (N_955,N_306,N_246);
and U956 (N_956,N_484,In_1608);
xnor U957 (N_957,In_891,N_489);
nand U958 (N_958,In_1933,In_1993);
nand U959 (N_959,In_212,In_2435);
nor U960 (N_960,N_32,N_144);
xor U961 (N_961,In_2184,N_161);
nand U962 (N_962,N_221,In_1392);
and U963 (N_963,In_637,In_996);
nand U964 (N_964,In_191,In_1321);
xor U965 (N_965,In_896,In_2301);
or U966 (N_966,N_76,In_508);
nor U967 (N_967,In_1453,In_1634);
and U968 (N_968,In_2114,In_1555);
or U969 (N_969,In_1038,In_1007);
xnor U970 (N_970,In_2383,In_1618);
xnor U971 (N_971,N_1,In_33);
or U972 (N_972,In_605,N_27);
and U973 (N_973,In_718,In_2013);
nor U974 (N_974,N_338,In_2248);
and U975 (N_975,In_1035,In_2362);
and U976 (N_976,In_742,In_360);
or U977 (N_977,In_600,In_2103);
and U978 (N_978,In_1666,In_1728);
xnor U979 (N_979,In_2052,In_1705);
and U980 (N_980,In_833,In_1722);
xnor U981 (N_981,In_913,In_939);
or U982 (N_982,In_2490,In_1667);
nor U983 (N_983,N_38,In_653);
xor U984 (N_984,In_2104,In_2122);
xor U985 (N_985,In_429,In_1381);
xnor U986 (N_986,In_730,In_2279);
nor U987 (N_987,In_2004,In_331);
nand U988 (N_988,In_533,In_1896);
or U989 (N_989,In_1284,In_1355);
and U990 (N_990,In_1147,In_82);
xor U991 (N_991,N_488,In_51);
nand U992 (N_992,In_754,N_203);
or U993 (N_993,In_2380,In_2234);
nand U994 (N_994,In_87,In_1969);
nor U995 (N_995,N_18,N_222);
nand U996 (N_996,In_71,In_2451);
nor U997 (N_997,In_1844,In_1341);
or U998 (N_998,In_2154,In_2206);
xnor U999 (N_999,In_2164,In_2091);
or U1000 (N_1000,N_307,In_1273);
and U1001 (N_1001,In_824,N_791);
and U1002 (N_1002,N_24,In_1046);
xnor U1003 (N_1003,N_985,In_2488);
nor U1004 (N_1004,In_1640,In_1661);
and U1005 (N_1005,In_1281,In_73);
nand U1006 (N_1006,N_170,In_1301);
xor U1007 (N_1007,In_1025,N_342);
nand U1008 (N_1008,In_1200,N_243);
nor U1009 (N_1009,N_312,N_641);
nand U1010 (N_1010,In_402,In_1537);
xor U1011 (N_1011,In_666,N_756);
nand U1012 (N_1012,N_925,In_1059);
and U1013 (N_1013,N_402,N_441);
nor U1014 (N_1014,N_989,In_684);
and U1015 (N_1015,In_1841,In_88);
xor U1016 (N_1016,N_768,N_536);
and U1017 (N_1017,In_2308,In_2419);
xnor U1018 (N_1018,N_77,N_773);
nor U1019 (N_1019,N_496,N_68);
and U1020 (N_1020,In_1539,In_1227);
or U1021 (N_1021,In_217,In_1957);
nand U1022 (N_1022,In_1853,N_869);
or U1023 (N_1023,In_128,N_916);
nand U1024 (N_1024,N_975,N_505);
or U1025 (N_1025,N_717,In_770);
nand U1026 (N_1026,N_433,In_2168);
or U1027 (N_1027,In_8,N_71);
nand U1028 (N_1028,In_2472,In_1393);
or U1029 (N_1029,In_1122,In_2386);
xor U1030 (N_1030,In_1630,N_520);
xor U1031 (N_1031,N_737,In_749);
nand U1032 (N_1032,In_2421,N_499);
xnor U1033 (N_1033,In_365,N_825);
or U1034 (N_1034,N_787,N_705);
and U1035 (N_1035,In_1713,N_8);
nor U1036 (N_1036,N_900,In_1676);
or U1037 (N_1037,In_2314,In_1900);
nand U1038 (N_1038,In_1049,N_104);
or U1039 (N_1039,In_590,N_274);
and U1040 (N_1040,N_576,N_933);
nor U1041 (N_1041,In_83,In_2384);
nor U1042 (N_1042,N_159,N_193);
nand U1043 (N_1043,In_210,In_2016);
nor U1044 (N_1044,In_940,In_231);
nor U1045 (N_1045,In_137,N_131);
xor U1046 (N_1046,N_735,N_356);
or U1047 (N_1047,In_1333,N_603);
nor U1048 (N_1048,In_780,N_478);
or U1049 (N_1049,In_2002,In_1015);
or U1050 (N_1050,In_629,In_311);
or U1051 (N_1051,In_1857,In_1578);
nand U1052 (N_1052,In_1870,N_248);
or U1053 (N_1053,In_1873,N_904);
nand U1054 (N_1054,In_1832,N_85);
nor U1055 (N_1055,In_1309,In_2290);
and U1056 (N_1056,N_861,N_815);
or U1057 (N_1057,In_100,In_909);
nand U1058 (N_1058,In_1020,In_2447);
xnor U1059 (N_1059,In_239,N_929);
nand U1060 (N_1060,In_2035,In_686);
and U1061 (N_1061,In_798,N_249);
nand U1062 (N_1062,N_530,N_631);
nand U1063 (N_1063,N_840,N_626);
or U1064 (N_1064,N_924,N_845);
or U1065 (N_1065,N_357,N_137);
and U1066 (N_1066,In_902,N_578);
or U1067 (N_1067,In_2003,In_114);
and U1068 (N_1068,In_1267,N_723);
or U1069 (N_1069,N_809,N_881);
nor U1070 (N_1070,N_509,In_1272);
xor U1071 (N_1071,In_198,N_979);
nor U1072 (N_1072,In_698,N_469);
or U1073 (N_1073,N_990,In_1913);
or U1074 (N_1074,N_456,N_558);
xor U1075 (N_1075,In_1701,In_1809);
nand U1076 (N_1076,N_343,In_297);
or U1077 (N_1077,N_868,N_780);
or U1078 (N_1078,N_800,N_575);
xnor U1079 (N_1079,N_884,In_61);
nor U1080 (N_1080,In_2425,N_403);
nor U1081 (N_1081,N_656,In_715);
nand U1082 (N_1082,In_669,In_566);
nand U1083 (N_1083,In_2197,In_2418);
or U1084 (N_1084,In_959,In_1551);
or U1085 (N_1085,In_11,In_545);
nand U1086 (N_1086,N_930,In_2217);
nand U1087 (N_1087,N_587,In_1755);
xor U1088 (N_1088,N_797,In_222);
xor U1089 (N_1089,In_200,In_2414);
nand U1090 (N_1090,N_219,In_554);
and U1091 (N_1091,N_988,In_1825);
nor U1092 (N_1092,In_46,In_1636);
nor U1093 (N_1093,N_50,In_2107);
nand U1094 (N_1094,In_2432,In_1760);
nand U1095 (N_1095,In_424,In_2320);
or U1096 (N_1096,N_864,N_801);
or U1097 (N_1097,N_710,N_795);
nor U1098 (N_1098,In_274,N_498);
and U1099 (N_1099,In_586,N_263);
or U1100 (N_1100,In_2254,N_836);
nor U1101 (N_1101,In_1985,In_265);
nor U1102 (N_1102,In_659,In_400);
or U1103 (N_1103,N_349,N_810);
or U1104 (N_1104,In_497,N_573);
xor U1105 (N_1105,In_540,N_224);
nand U1106 (N_1106,In_634,In_2075);
nand U1107 (N_1107,N_907,In_1461);
or U1108 (N_1108,In_616,N_194);
or U1109 (N_1109,N_204,N_908);
and U1110 (N_1110,In_1388,In_1646);
or U1111 (N_1111,In_1926,In_1300);
xor U1112 (N_1112,In_1093,N_738);
nor U1113 (N_1113,N_464,In_958);
nand U1114 (N_1114,In_1877,N_610);
nor U1115 (N_1115,N_701,In_1258);
nand U1116 (N_1116,N_230,N_839);
xnor U1117 (N_1117,In_10,N_950);
nand U1118 (N_1118,N_207,N_412);
and U1119 (N_1119,In_1907,N_158);
nand U1120 (N_1120,N_331,In_1593);
nand U1121 (N_1121,N_572,N_147);
and U1122 (N_1122,In_1340,N_666);
nor U1123 (N_1123,N_630,N_684);
xnor U1124 (N_1124,In_1793,In_253);
xor U1125 (N_1125,In_80,N_108);
xor U1126 (N_1126,N_541,In_474);
nand U1127 (N_1127,N_849,N_808);
xnor U1128 (N_1128,In_461,N_52);
or U1129 (N_1129,N_143,N_596);
and U1130 (N_1130,In_797,In_1569);
or U1131 (N_1131,N_680,N_672);
xnor U1132 (N_1132,N_724,N_677);
or U1133 (N_1133,In_2347,N_886);
and U1134 (N_1134,N_866,In_1934);
nor U1135 (N_1135,N_619,N_769);
nor U1136 (N_1136,N_972,N_678);
and U1137 (N_1137,In_1808,In_464);
nor U1138 (N_1138,N_212,In_1891);
nand U1139 (N_1139,In_2221,In_2138);
or U1140 (N_1140,N_696,N_585);
nor U1141 (N_1141,In_1003,N_646);
or U1142 (N_1142,N_535,N_141);
and U1143 (N_1143,N_501,In_2118);
or U1144 (N_1144,In_1045,N_679);
or U1145 (N_1145,N_0,N_987);
nand U1146 (N_1146,N_561,N_759);
or U1147 (N_1147,In_2293,In_2438);
nor U1148 (N_1148,In_1165,N_435);
nand U1149 (N_1149,In_2011,N_191);
nand U1150 (N_1150,In_2469,In_20);
nand U1151 (N_1151,N_466,In_748);
and U1152 (N_1152,N_17,N_612);
nor U1153 (N_1153,In_1234,N_816);
or U1154 (N_1154,N_580,In_1220);
nand U1155 (N_1155,In_1804,N_841);
xor U1156 (N_1156,N_387,N_481);
and U1157 (N_1157,N_942,N_34);
nor U1158 (N_1158,N_309,In_2108);
nor U1159 (N_1159,In_1190,In_1796);
nor U1160 (N_1160,In_1127,N_517);
nand U1161 (N_1161,N_78,N_931);
xnor U1162 (N_1162,N_289,In_1085);
xor U1163 (N_1163,In_1994,N_16);
nand U1164 (N_1164,In_2036,In_2098);
and U1165 (N_1165,N_471,N_223);
xnor U1166 (N_1166,In_1868,N_318);
nand U1167 (N_1167,In_63,In_568);
nor U1168 (N_1168,In_325,In_500);
nor U1169 (N_1169,N_711,In_2144);
or U1170 (N_1170,N_846,In_734);
nand U1171 (N_1171,In_229,In_1357);
and U1172 (N_1172,N_316,In_2404);
xnor U1173 (N_1173,In_355,In_117);
xor U1174 (N_1174,In_2034,In_2437);
xnor U1175 (N_1175,In_1846,N_682);
xor U1176 (N_1176,In_67,In_1323);
or U1177 (N_1177,In_1271,In_1880);
and U1178 (N_1178,In_113,In_343);
or U1179 (N_1179,N_245,In_205);
and U1180 (N_1180,In_838,N_794);
nor U1181 (N_1181,N_745,N_921);
xnor U1182 (N_1182,In_166,In_898);
nand U1183 (N_1183,N_640,N_771);
xnor U1184 (N_1184,In_178,In_1691);
xor U1185 (N_1185,In_2141,In_922);
or U1186 (N_1186,In_573,N_664);
nand U1187 (N_1187,In_2422,N_57);
or U1188 (N_1188,In_2083,In_925);
nand U1189 (N_1189,In_1413,In_14);
and U1190 (N_1190,N_39,In_2356);
or U1191 (N_1191,In_2354,N_986);
or U1192 (N_1192,N_758,N_238);
and U1193 (N_1193,In_2449,In_1955);
xnor U1194 (N_1194,N_653,N_681);
or U1195 (N_1195,N_415,In_1307);
and U1196 (N_1196,In_729,N_225);
xor U1197 (N_1197,In_1945,N_729);
and U1198 (N_1198,In_982,In_722);
or U1199 (N_1199,In_1482,In_2216);
or U1200 (N_1200,N_788,In_1996);
and U1201 (N_1201,N_870,N_867);
or U1202 (N_1202,N_635,In_2160);
nand U1203 (N_1203,In_1813,In_1735);
nor U1204 (N_1204,N_534,N_667);
and U1205 (N_1205,In_2143,In_1435);
nand U1206 (N_1206,In_1778,N_704);
and U1207 (N_1207,In_2101,N_693);
or U1208 (N_1208,In_1331,In_1632);
and U1209 (N_1209,In_2390,N_736);
and U1210 (N_1210,In_1201,N_790);
nand U1211 (N_1211,In_1908,N_457);
or U1212 (N_1212,N_109,In_2152);
and U1213 (N_1213,N_982,In_1770);
nor U1214 (N_1214,In_1772,In_119);
or U1215 (N_1215,In_755,In_493);
xor U1216 (N_1216,N_568,In_550);
xnor U1217 (N_1217,N_686,N_707);
nor U1218 (N_1218,N_70,N_418);
xor U1219 (N_1219,N_636,In_135);
and U1220 (N_1220,N_388,In_1245);
xor U1221 (N_1221,N_142,In_2342);
nor U1222 (N_1222,N_66,N_938);
and U1223 (N_1223,N_368,N_948);
xnor U1224 (N_1224,N_529,N_962);
nand U1225 (N_1225,N_29,In_221);
or U1226 (N_1226,In_1,In_406);
nand U1227 (N_1227,In_1297,In_479);
xnor U1228 (N_1228,In_2460,In_1458);
nor U1229 (N_1229,In_694,N_752);
nor U1230 (N_1230,N_969,N_963);
and U1231 (N_1231,N_36,N_826);
nor U1232 (N_1232,N_453,N_83);
xor U1233 (N_1233,In_1114,N_865);
nand U1234 (N_1234,N_749,N_569);
nor U1235 (N_1235,N_586,N_740);
nand U1236 (N_1236,N_973,In_2397);
or U1237 (N_1237,N_814,In_426);
xor U1238 (N_1238,N_302,N_296);
or U1239 (N_1239,In_685,N_624);
nor U1240 (N_1240,In_678,In_2458);
nor U1241 (N_1241,N_172,N_882);
nor U1242 (N_1242,In_1942,N_943);
nor U1243 (N_1243,In_1329,N_591);
and U1244 (N_1244,N_685,N_760);
nand U1245 (N_1245,N_981,N_213);
xor U1246 (N_1246,N_363,In_1452);
nand U1247 (N_1247,N_401,N_721);
nor U1248 (N_1248,N_910,N_663);
or U1249 (N_1249,In_693,N_511);
nor U1250 (N_1250,N_325,N_236);
xor U1251 (N_1251,In_2142,In_966);
nand U1252 (N_1252,In_1491,N_926);
nor U1253 (N_1253,In_1084,In_96);
or U1254 (N_1254,N_588,N_658);
or U1255 (N_1255,In_503,N_675);
nor U1256 (N_1256,N_436,In_2);
nor U1257 (N_1257,N_61,N_673);
xnor U1258 (N_1258,In_55,In_1042);
or U1259 (N_1259,In_1487,N_633);
nor U1260 (N_1260,N_905,In_793);
nand U1261 (N_1261,In_1189,N_842);
nor U1262 (N_1262,N_227,In_2282);
or U1263 (N_1263,N_783,In_1510);
nand U1264 (N_1264,In_1069,In_1866);
xnor U1265 (N_1265,N_700,In_943);
xnor U1266 (N_1266,In_183,N_932);
xnor U1267 (N_1267,In_1494,N_713);
xor U1268 (N_1268,In_825,In_1709);
and U1269 (N_1269,In_1153,N_628);
or U1270 (N_1270,In_309,N_784);
xnor U1271 (N_1271,N_722,N_351);
xor U1272 (N_1272,N_598,N_54);
and U1273 (N_1273,In_2484,N_730);
or U1274 (N_1274,N_583,N_731);
xnor U1275 (N_1275,In_445,In_19);
xnor U1276 (N_1276,N_548,N_454);
xnor U1277 (N_1277,N_577,N_824);
nand U1278 (N_1278,In_2056,N_838);
nand U1279 (N_1279,In_2146,In_1407);
and U1280 (N_1280,N_657,N_461);
or U1281 (N_1281,N_602,In_2009);
nand U1282 (N_1282,In_1805,N_549);
or U1283 (N_1283,In_182,In_781);
nand U1284 (N_1284,N_774,In_1028);
or U1285 (N_1285,N_947,In_806);
nand U1286 (N_1286,In_1668,In_1466);
nand U1287 (N_1287,In_836,In_278);
nor U1288 (N_1288,In_553,In_1547);
nand U1289 (N_1289,In_796,N_763);
xnor U1290 (N_1290,N_831,In_2134);
and U1291 (N_1291,In_95,N_694);
nand U1292 (N_1292,N_835,N_789);
and U1293 (N_1293,N_516,In_1858);
nand U1294 (N_1294,N_594,In_342);
nor U1295 (N_1295,N_638,In_2350);
xnor U1296 (N_1296,In_1080,N_964);
nor U1297 (N_1297,In_973,N_959);
xor U1298 (N_1298,N_579,N_876);
xnor U1299 (N_1299,N_30,N_823);
and U1300 (N_1300,In_1716,N_874);
or U1301 (N_1301,N_891,N_135);
nor U1302 (N_1302,N_51,In_1351);
or U1303 (N_1303,In_2309,In_37);
xnor U1304 (N_1304,In_1445,In_1089);
nand U1305 (N_1305,In_190,In_671);
nand U1306 (N_1306,In_1198,In_1723);
nor U1307 (N_1307,In_163,N_555);
and U1308 (N_1308,N_424,In_1374);
xnor U1309 (N_1309,N_819,In_2208);
xor U1310 (N_1310,In_115,In_2158);
or U1311 (N_1311,In_193,N_178);
nand U1312 (N_1312,In_1095,In_1621);
and U1313 (N_1313,In_2385,N_632);
or U1314 (N_1314,In_1514,In_1422);
nand U1315 (N_1315,N_411,N_165);
nor U1316 (N_1316,In_719,In_606);
and U1317 (N_1317,In_1573,N_118);
or U1318 (N_1318,N_850,N_651);
nand U1319 (N_1319,N_621,N_940);
xnor U1320 (N_1320,N_62,N_703);
or U1321 (N_1321,In_1726,N_652);
nor U1322 (N_1322,N_262,In_171);
nand U1323 (N_1323,In_1383,In_1614);
xor U1324 (N_1324,In_2120,In_1872);
nor U1325 (N_1325,N_100,In_1875);
xor U1326 (N_1326,In_2214,In_563);
nand U1327 (N_1327,In_1768,In_1619);
xnor U1328 (N_1328,N_138,In_581);
and U1329 (N_1329,In_349,N_582);
xor U1330 (N_1330,In_519,N_605);
nor U1331 (N_1331,In_1037,N_977);
or U1332 (N_1332,N_936,N_855);
xor U1333 (N_1333,N_778,In_2110);
or U1334 (N_1334,N_277,N_44);
and U1335 (N_1335,N_995,N_880);
nor U1336 (N_1336,In_726,N_563);
nor U1337 (N_1337,N_779,N_72);
xor U1338 (N_1338,In_2476,In_1560);
xnor U1339 (N_1339,In_2201,In_2482);
and U1340 (N_1340,N_899,In_246);
nor U1341 (N_1341,In_597,In_1721);
xor U1342 (N_1342,N_851,In_1021);
or U1343 (N_1343,N_944,In_1863);
nor U1344 (N_1344,In_1637,N_743);
and U1345 (N_1345,In_1690,In_2022);
xnor U1346 (N_1346,In_403,N_381);
and U1347 (N_1347,N_515,In_2230);
xnor U1348 (N_1348,N_152,In_1542);
nor U1349 (N_1349,N_793,In_1682);
nor U1350 (N_1350,In_1780,In_878);
nand U1351 (N_1351,In_159,N_371);
xnor U1352 (N_1352,N_719,In_469);
xor U1353 (N_1353,N_237,N_806);
and U1354 (N_1354,N_898,In_928);
xor U1355 (N_1355,In_125,In_1848);
and U1356 (N_1356,In_2334,In_488);
or U1357 (N_1357,In_1752,N_94);
or U1358 (N_1358,In_1171,In_968);
or U1359 (N_1359,N_294,N_127);
xnor U1360 (N_1360,In_867,N_807);
nor U1361 (N_1361,In_1133,N_545);
and U1362 (N_1362,In_384,N_599);
or U1363 (N_1363,In_492,N_606);
or U1364 (N_1364,N_837,N_367);
nor U1365 (N_1365,In_2353,In_1575);
xnor U1366 (N_1366,N_966,N_571);
nor U1367 (N_1367,N_643,N_546);
and U1368 (N_1368,N_22,N_967);
xnor U1369 (N_1369,In_1030,In_423);
xnor U1370 (N_1370,N_951,In_275);
xor U1371 (N_1371,N_957,In_1325);
or U1372 (N_1372,N_877,N_220);
nand U1373 (N_1373,N_10,In_201);
nor U1374 (N_1374,In_328,In_2094);
or U1375 (N_1375,In_1501,In_1299);
xor U1376 (N_1376,N_89,N_714);
nand U1377 (N_1377,In_1599,N_525);
or U1378 (N_1378,In_731,In_743);
and U1379 (N_1379,N_554,In_23);
nor U1380 (N_1380,N_560,N_74);
nand U1381 (N_1381,N_629,In_1072);
nand U1382 (N_1382,N_452,In_34);
nor U1383 (N_1383,In_1920,N_798);
nand U1384 (N_1384,In_826,In_2344);
and U1385 (N_1385,In_2235,In_2136);
and U1386 (N_1386,In_920,N_726);
and U1387 (N_1387,N_915,In_108);
nand U1388 (N_1388,N_25,In_2388);
and U1389 (N_1389,N_716,In_2348);
or U1390 (N_1390,N_970,In_1936);
and U1391 (N_1391,In_938,In_914);
nor U1392 (N_1392,In_462,N_542);
or U1393 (N_1393,N_968,In_2163);
or U1394 (N_1394,N_341,N_217);
or U1395 (N_1395,In_446,N_514);
nor U1396 (N_1396,N_544,In_2194);
nand U1397 (N_1397,N_81,N_422);
nand U1398 (N_1398,In_1412,In_763);
or U1399 (N_1399,N_518,N_176);
or U1400 (N_1400,N_234,In_863);
xor U1401 (N_1401,In_444,In_1347);
or U1402 (N_1402,In_1241,N_978);
nand U1403 (N_1403,N_818,In_1707);
xor U1404 (N_1404,In_1743,N_269);
nand U1405 (N_1405,In_1906,N_537);
nor U1406 (N_1406,N_570,N_927);
xor U1407 (N_1407,In_1469,In_577);
xnor U1408 (N_1408,N_482,In_1073);
nor U1409 (N_1409,In_1506,N_490);
xnor U1410 (N_1410,N_355,In_1313);
nor U1411 (N_1411,N_475,In_344);
nand U1412 (N_1412,In_1952,In_932);
xnor U1413 (N_1413,N_283,In_374);
and U1414 (N_1414,In_2368,In_2341);
and U1415 (N_1415,N_875,In_1327);
xor U1416 (N_1416,N_584,In_306);
or U1417 (N_1417,N_361,In_762);
or U1418 (N_1418,N_84,In_919);
and U1419 (N_1419,N_510,In_1651);
nor U1420 (N_1420,In_680,N_556);
nor U1421 (N_1421,N_895,In_2378);
xor U1422 (N_1422,N_872,N_993);
and U1423 (N_1423,N_613,In_740);
xnor U1424 (N_1424,In_1812,In_176);
xnor U1425 (N_1425,In_655,N_702);
xnor U1426 (N_1426,N_335,In_1581);
xnor U1427 (N_1427,N_375,In_1041);
nor U1428 (N_1428,In_240,N_862);
nor U1429 (N_1429,N_956,In_645);
nor U1430 (N_1430,In_484,In_4);
xor U1431 (N_1431,N_669,In_1110);
or U1432 (N_1432,N_953,In_800);
nor U1433 (N_1433,In_187,N_668);
or U1434 (N_1434,In_1240,In_1261);
and U1435 (N_1435,In_289,N_133);
nor U1436 (N_1436,In_1447,N_890);
nand U1437 (N_1437,In_1792,N_378);
and U1438 (N_1438,In_1826,N_285);
xnor U1439 (N_1439,N_856,N_46);
xnor U1440 (N_1440,In_890,N_28);
and U1441 (N_1441,In_44,In_1767);
and U1442 (N_1442,In_2412,In_391);
and U1443 (N_1443,In_944,N_215);
nand U1444 (N_1444,In_337,N_708);
nor U1445 (N_1445,N_999,N_205);
and U1446 (N_1446,N_443,In_1563);
or U1447 (N_1447,N_939,In_823);
or U1448 (N_1448,In_1536,N_321);
xnor U1449 (N_1449,N_954,In_2238);
and U1450 (N_1450,In_457,N_893);
and U1451 (N_1451,In_1538,N_506);
xnor U1452 (N_1452,N_106,N_733);
nand U1453 (N_1453,N_4,In_419);
nor U1454 (N_1454,N_532,N_960);
nor U1455 (N_1455,In_86,In_375);
nor U1456 (N_1456,In_2292,N_828);
and U1457 (N_1457,In_1526,In_1839);
nor U1458 (N_1458,N_946,In_1545);
nand U1459 (N_1459,N_813,N_421);
xnor U1460 (N_1460,N_600,N_192);
nor U1461 (N_1461,N_186,N_589);
and U1462 (N_1462,N_267,N_805);
xor U1463 (N_1463,N_625,In_1992);
and U1464 (N_1464,In_2400,In_207);
nand U1465 (N_1465,In_2494,N_648);
and U1466 (N_1466,N_190,In_241);
and U1467 (N_1467,N_983,N_199);
or U1468 (N_1468,In_993,In_1528);
or U1469 (N_1469,In_131,N_559);
and U1470 (N_1470,In_1278,N_848);
nor U1471 (N_1471,N_414,In_839);
or U1472 (N_1472,N_802,N_920);
and U1473 (N_1473,N_339,N_597);
and U1474 (N_1474,In_811,N_634);
nand U1475 (N_1475,N_369,N_173);
nand U1476 (N_1476,N_732,N_379);
xor U1477 (N_1477,In_816,N_614);
nor U1478 (N_1478,In_140,In_1376);
and U1479 (N_1479,In_69,In_2295);
or U1480 (N_1480,N_14,In_2364);
nand U1481 (N_1481,N_695,N_595);
and U1482 (N_1482,N_526,In_282);
or U1483 (N_1483,N_670,N_853);
nor U1484 (N_1484,N_655,N_557);
or U1485 (N_1485,In_2263,N_429);
and U1486 (N_1486,In_869,N_416);
or U1487 (N_1487,In_567,In_1586);
and U1488 (N_1488,N_775,N_622);
nor U1489 (N_1489,N_254,N_399);
and U1490 (N_1490,N_615,In_1243);
xnor U1491 (N_1491,In_104,N_937);
or U1492 (N_1492,N_691,In_2006);
xnor U1493 (N_1493,In_807,In_1034);
or U1494 (N_1494,N_776,N_689);
nand U1495 (N_1495,N_698,N_502);
nand U1496 (N_1496,In_1265,N_734);
and U1497 (N_1497,N_889,In_470);
nor U1498 (N_1498,N_935,N_639);
xnor U1499 (N_1499,N_533,In_2204);
xor U1500 (N_1500,N_1049,N_608);
and U1501 (N_1501,N_1405,N_1075);
or U1502 (N_1502,N_1178,N_266);
nor U1503 (N_1503,In_2357,N_1264);
and U1504 (N_1504,In_65,In_819);
or U1505 (N_1505,N_1058,N_1209);
nor U1506 (N_1506,N_1092,N_843);
nor U1507 (N_1507,In_180,N_1488);
or U1508 (N_1508,N_1274,N_1008);
or U1509 (N_1509,N_607,In_893);
or U1510 (N_1510,In_1851,N_637);
and U1511 (N_1511,In_2015,In_602);
and U1512 (N_1512,N_1116,N_1187);
or U1513 (N_1513,In_1348,N_1216);
nand U1514 (N_1514,N_581,N_1007);
and U1515 (N_1515,N_1341,In_1434);
xor U1516 (N_1516,N_1230,N_1380);
nor U1517 (N_1517,N_1284,N_1223);
or U1518 (N_1518,N_1250,N_1111);
xor U1519 (N_1519,N_1466,N_1252);
or U1520 (N_1520,In_90,N_1379);
and U1521 (N_1521,N_1248,N_1081);
nand U1522 (N_1522,N_654,N_1040);
nand U1523 (N_1523,N_971,N_1027);
or U1524 (N_1524,N_1154,In_764);
nand U1525 (N_1525,In_1692,N_1325);
nor U1526 (N_1526,N_1445,N_1393);
nand U1527 (N_1527,In_1706,In_452);
nand U1528 (N_1528,N_426,In_294);
xor U1529 (N_1529,In_1830,N_1382);
and U1530 (N_1530,N_1061,In_916);
and U1531 (N_1531,N_1469,N_1195);
or U1532 (N_1532,N_538,N_524);
nor U1533 (N_1533,N_1074,N_699);
nand U1534 (N_1534,In_2175,N_1104);
nor U1535 (N_1535,In_2317,N_1210);
or U1536 (N_1536,N_1304,N_1428);
or U1537 (N_1537,N_1189,N_833);
xnor U1538 (N_1538,N_1055,N_887);
or U1539 (N_1539,N_1366,N_1381);
nor U1540 (N_1540,N_620,N_1109);
and U1541 (N_1541,In_408,In_2247);
nor U1542 (N_1542,N_706,N_1121);
xnor U1543 (N_1543,N_945,In_1175);
or U1544 (N_1544,N_1408,N_543);
or U1545 (N_1545,N_1082,N_1181);
and U1546 (N_1546,N_42,N_1482);
nand U1547 (N_1547,N_857,N_1174);
nor U1548 (N_1548,N_1011,N_1450);
nand U1549 (N_1549,In_458,In_1490);
xor U1550 (N_1550,N_1120,N_1468);
or U1551 (N_1551,N_1493,In_1263);
nor U1552 (N_1552,N_718,N_1254);
nand U1553 (N_1553,In_1861,N_1371);
and U1554 (N_1554,N_1140,In_2433);
xor U1555 (N_1555,N_1346,N_1460);
xnor U1556 (N_1556,N_1395,N_1378);
or U1557 (N_1557,In_1087,In_608);
nor U1558 (N_1558,N_1161,N_1387);
nand U1559 (N_1559,N_1278,N_352);
nand U1560 (N_1560,In_1242,In_773);
nor U1561 (N_1561,In_613,In_1527);
nor U1562 (N_1562,N_649,N_1012);
xnor U1563 (N_1563,In_2367,N_1283);
or U1564 (N_1564,N_1227,N_1037);
or U1565 (N_1565,In_557,N_1164);
or U1566 (N_1566,N_43,N_1159);
nand U1567 (N_1567,N_692,N_1041);
and U1568 (N_1568,N_347,N_888);
and U1569 (N_1569,N_1355,In_1160);
and U1570 (N_1570,N_1280,N_991);
and U1571 (N_1571,N_547,In_2213);
or U1572 (N_1572,In_333,N_1090);
xnor U1573 (N_1573,N_961,In_189);
nor U1574 (N_1574,N_1259,N_1184);
nand U1575 (N_1575,N_1310,N_746);
and U1576 (N_1576,N_551,N_1483);
or U1577 (N_1577,N_1130,N_1175);
xnor U1578 (N_1578,N_767,N_419);
or U1579 (N_1579,N_1461,N_781);
nor U1580 (N_1580,N_829,N_1391);
xnor U1581 (N_1581,N_1351,N_1155);
or U1582 (N_1582,N_1067,N_1420);
nor U1583 (N_1583,In_1680,N_770);
and U1584 (N_1584,N_593,N_293);
or U1585 (N_1585,N_1449,N_1125);
or U1586 (N_1586,N_1267,N_873);
and U1587 (N_1587,N_1233,N_1349);
or U1588 (N_1588,N_1285,N_522);
xnor U1589 (N_1589,N_659,N_110);
nand U1590 (N_1590,N_1415,N_1403);
xor U1591 (N_1591,N_1261,N_1481);
or U1592 (N_1592,N_1098,N_923);
or U1593 (N_1593,N_1451,N_1052);
xor U1594 (N_1594,N_941,N_1272);
and U1595 (N_1595,N_1242,N_741);
nor U1596 (N_1596,N_1103,N_1432);
nor U1597 (N_1597,N_765,N_1214);
xor U1598 (N_1598,N_1473,N_1047);
nor U1599 (N_1599,N_268,N_112);
or U1600 (N_1600,N_671,N_507);
or U1601 (N_1601,N_1462,N_688);
xnor U1602 (N_1602,N_592,In_1822);
xnor U1603 (N_1603,In_2369,In_1835);
xnor U1604 (N_1604,N_1013,N_1228);
nor U1605 (N_1605,N_1307,In_901);
and U1606 (N_1606,N_623,N_811);
and U1607 (N_1607,N_739,N_1335);
xor U1608 (N_1608,In_776,N_1484);
or U1609 (N_1609,N_1263,In_1961);
and U1610 (N_1610,N_847,N_1376);
and U1611 (N_1611,N_1016,In_1984);
xor U1612 (N_1612,N_1245,N_1309);
nand U1613 (N_1613,In_2085,N_446);
and U1614 (N_1614,N_753,N_1028);
nor U1615 (N_1615,N_1394,N_1035);
nand U1616 (N_1616,N_1367,N_1162);
nand U1617 (N_1617,N_1318,N_1324);
xnor U1618 (N_1618,N_1319,N_1200);
or U1619 (N_1619,In_1633,N_119);
nand U1620 (N_1620,In_1437,N_1066);
xor U1621 (N_1621,N_1235,In_1074);
xor U1622 (N_1622,N_1133,N_1072);
and U1623 (N_1623,In_130,N_528);
and U1624 (N_1624,N_1176,N_1206);
and U1625 (N_1625,N_1357,N_1426);
and U1626 (N_1626,N_1207,In_1738);
nor U1627 (N_1627,N_1490,In_785);
nor U1628 (N_1628,In_1464,In_2119);
nor U1629 (N_1629,N_998,N_1330);
xor U1630 (N_1630,In_1867,N_1157);
nor U1631 (N_1631,N_552,N_1265);
or U1632 (N_1632,N_897,N_504);
xor U1633 (N_1633,In_1238,In_2076);
and U1634 (N_1634,N_1089,In_895);
xnor U1635 (N_1635,N_333,N_300);
nand U1636 (N_1636,N_992,N_150);
nand U1637 (N_1637,N_1277,In_1317);
nand U1638 (N_1638,In_1485,In_1595);
nand U1639 (N_1639,N_442,N_40);
or U1640 (N_1640,N_1059,In_1471);
xor U1641 (N_1641,N_650,N_662);
nor U1642 (N_1642,In_2339,In_2459);
or U1643 (N_1643,N_1279,In_621);
nand U1644 (N_1644,N_1053,N_531);
nand U1645 (N_1645,N_96,N_1193);
nor U1646 (N_1646,N_449,In_2185);
xnor U1647 (N_1647,N_764,N_1105);
nor U1648 (N_1648,In_326,N_1459);
nand U1649 (N_1649,In_1359,N_444);
nand U1650 (N_1650,N_683,In_228);
xnor U1651 (N_1651,N_830,N_1316);
nand U1652 (N_1652,N_1220,N_1009);
nand U1653 (N_1653,N_1196,In_1488);
nand U1654 (N_1654,N_1056,In_28);
and U1655 (N_1655,N_757,N_906);
or U1656 (N_1656,N_1485,N_1418);
nor U1657 (N_1657,N_231,N_1491);
nor U1658 (N_1658,N_1317,N_852);
nor U1659 (N_1659,N_1088,N_500);
nor U1660 (N_1660,N_467,In_872);
or U1661 (N_1661,In_1191,N_1084);
or U1662 (N_1662,In_2024,N_1326);
nor U1663 (N_1663,In_2426,N_1114);
xor U1664 (N_1664,N_1253,N_1434);
or U1665 (N_1665,N_1477,N_202);
or U1666 (N_1666,In_1925,N_1298);
nand U1667 (N_1667,N_562,In_235);
or U1668 (N_1668,N_1118,N_527);
nor U1669 (N_1669,In_509,N_1457);
xnor U1670 (N_1670,In_2236,N_1410);
and U1671 (N_1671,N_1444,N_1303);
nand U1672 (N_1672,N_1249,In_489);
nor U1673 (N_1673,N_508,N_1127);
or U1674 (N_1674,N_214,N_863);
nand U1675 (N_1675,In_814,N_280);
nor U1676 (N_1676,In_1577,N_405);
or U1677 (N_1677,N_397,In_2325);
xnor U1678 (N_1678,In_1610,N_1475);
or U1679 (N_1679,N_1026,N_1365);
and U1680 (N_1680,In_1930,In_1109);
xor U1681 (N_1681,N_1050,N_1476);
nand U1682 (N_1682,N_218,N_1023);
nor U1683 (N_1683,In_2477,N_1498);
and U1684 (N_1684,N_1168,N_1244);
xor U1685 (N_1685,N_820,In_1941);
or U1686 (N_1686,N_761,In_2300);
xor U1687 (N_1687,N_1054,N_1268);
nor U1688 (N_1688,N_949,N_1229);
nand U1689 (N_1689,N_997,In_1441);
xnor U1690 (N_1690,In_2199,N_883);
and U1691 (N_1691,N_1455,N_1375);
nand U1692 (N_1692,N_1302,N_1281);
and U1693 (N_1693,N_1290,N_146);
or U1694 (N_1694,N_450,N_1204);
and U1695 (N_1695,In_864,N_980);
xnor U1696 (N_1696,N_821,N_1062);
nor U1697 (N_1697,N_184,N_1078);
xnor U1698 (N_1698,N_1386,N_1292);
nor U1699 (N_1699,In_1259,N_1332);
xnor U1700 (N_1700,N_1407,N_1427);
nor U1701 (N_1701,N_1400,N_1000);
and U1702 (N_1702,N_1003,N_574);
nor U1703 (N_1703,N_125,In_1411);
and U1704 (N_1704,N_1138,N_1406);
or U1705 (N_1705,N_871,In_1674);
or U1706 (N_1706,N_382,N_1010);
or U1707 (N_1707,In_2359,In_884);
or U1708 (N_1708,In_2338,In_2493);
nor U1709 (N_1709,In_2187,In_1209);
nor U1710 (N_1710,N_1313,In_1882);
nand U1711 (N_1711,N_550,N_1496);
nand U1712 (N_1712,In_735,N_1487);
nor U1713 (N_1713,In_2310,N_1306);
nor U1714 (N_1714,N_1396,N_647);
nand U1715 (N_1715,In_2131,N_1424);
or U1716 (N_1716,N_859,N_123);
nand U1717 (N_1717,N_1238,N_1399);
nor U1718 (N_1718,N_644,N_253);
nand U1719 (N_1719,In_1101,N_1201);
nand U1720 (N_1720,In_537,N_1100);
nor U1721 (N_1721,N_65,In_716);
nand U1722 (N_1722,N_1364,N_1107);
nand U1723 (N_1723,In_150,N_1431);
and U1724 (N_1724,N_434,N_1173);
nand U1725 (N_1725,In_677,N_1202);
and U1726 (N_1726,In_521,N_241);
and U1727 (N_1727,N_1094,In_528);
nor U1728 (N_1728,N_762,N_1308);
nand U1729 (N_1729,In_1583,N_1147);
nand U1730 (N_1730,N_928,N_1288);
xnor U1731 (N_1731,N_1015,In_2420);
xor U1732 (N_1732,In_127,In_2051);
nand U1733 (N_1733,N_1160,In_2243);
nand U1734 (N_1734,N_1441,N_1240);
nand U1735 (N_1735,N_1042,N_1231);
nor U1736 (N_1736,N_690,N_427);
or U1737 (N_1737,In_81,N_1260);
nor U1738 (N_1738,N_1255,N_1199);
nor U1739 (N_1739,N_1102,In_341);
or U1740 (N_1740,N_728,N_1036);
nand U1741 (N_1741,N_1137,N_1348);
or U1742 (N_1742,N_720,N_1124);
and U1743 (N_1743,N_1063,N_179);
nand U1744 (N_1744,N_284,N_183);
nand U1745 (N_1745,N_1002,N_1232);
and U1746 (N_1746,N_1217,N_1142);
nor U1747 (N_1747,N_742,N_715);
xnor U1748 (N_1748,N_1091,In_1451);
and U1749 (N_1749,N_1043,N_1294);
or U1750 (N_1750,N_1024,N_1225);
nor U1751 (N_1751,In_603,In_1455);
or U1752 (N_1752,N_1397,N_1270);
xor U1753 (N_1753,N_1392,N_1384);
or U1754 (N_1754,N_1243,N_1293);
or U1755 (N_1755,N_1276,N_1197);
xor U1756 (N_1756,N_642,N_1369);
nor U1757 (N_1757,In_650,N_167);
and U1758 (N_1758,In_858,N_299);
or U1759 (N_1759,N_1005,N_282);
or U1760 (N_1760,N_1186,N_1320);
or U1761 (N_1761,N_984,N_1172);
nand U1762 (N_1762,N_1134,N_1033);
or U1763 (N_1763,N_958,N_922);
nand U1764 (N_1764,In_1968,N_1354);
or U1765 (N_1765,N_1422,N_271);
or U1766 (N_1766,N_1385,In_1919);
and U1767 (N_1767,In_2351,N_1323);
and U1768 (N_1768,In_2209,N_601);
nor U1769 (N_1769,N_1071,N_423);
nand U1770 (N_1770,N_1312,In_1890);
nand U1771 (N_1771,N_1438,N_1014);
nor U1772 (N_1772,N_322,In_2049);
xor U1773 (N_1773,N_1039,In_1817);
xor U1774 (N_1774,N_1131,N_1425);
nand U1775 (N_1775,N_860,In_2283);
and U1776 (N_1776,In_1656,N_1203);
nand U1777 (N_1777,In_1216,N_1353);
nand U1778 (N_1778,In_2373,In_2172);
xnor U1779 (N_1779,N_834,N_1358);
nor U1780 (N_1780,N_1336,N_1372);
or U1781 (N_1781,N_1239,N_151);
and U1782 (N_1782,N_519,In_1222);
and U1783 (N_1783,N_1343,N_1170);
nor U1784 (N_1784,N_1416,In_1971);
nor U1785 (N_1785,N_1271,N_1262);
nor U1786 (N_1786,N_1144,N_1087);
xnor U1787 (N_1787,N_1322,N_1374);
xor U1788 (N_1788,N_1106,N_566);
and U1789 (N_1789,In_579,N_1057);
or U1790 (N_1790,N_385,N_1241);
nor U1791 (N_1791,In_1940,N_1083);
xor U1792 (N_1792,N_1388,N_1031);
or U1793 (N_1793,N_1183,In_885);
nand U1794 (N_1794,N_858,N_1212);
xnor U1795 (N_1795,In_262,N_1177);
nor U1796 (N_1796,N_348,N_917);
and U1797 (N_1797,N_395,N_1305);
xor U1798 (N_1798,N_1299,N_1219);
and U1799 (N_1799,In_12,N_1373);
nand U1800 (N_1800,N_822,In_1135);
nor U1801 (N_1801,N_725,N_1167);
or U1802 (N_1802,N_1065,N_565);
or U1803 (N_1803,N_712,N_1234);
or U1804 (N_1804,N_1287,N_616);
xor U1805 (N_1805,N_1115,N_1070);
or U1806 (N_1806,N_1096,N_1086);
or U1807 (N_1807,N_627,N_390);
or U1808 (N_1808,N_1421,N_1150);
and U1809 (N_1809,N_503,N_345);
nor U1810 (N_1810,N_1205,N_676);
xor U1811 (N_1811,N_674,In_2324);
and U1812 (N_1812,N_976,N_523);
or U1813 (N_1813,In_1217,In_955);
or U1814 (N_1814,N_432,In_1082);
nand U1815 (N_1815,In_805,N_1030);
xor U1816 (N_1816,N_308,N_902);
nand U1817 (N_1817,N_1339,N_185);
and U1818 (N_1818,N_1158,N_1472);
or U1819 (N_1819,N_912,N_744);
and U1820 (N_1820,N_1480,N_1337);
nand U1821 (N_1821,N_1051,N_617);
and U1822 (N_1822,In_803,N_1165);
nand U1823 (N_1823,In_1750,N_1085);
or U1824 (N_1824,N_344,N_1101);
xor U1825 (N_1825,N_251,N_1236);
nand U1826 (N_1826,N_1218,In_2000);
or U1827 (N_1827,N_1029,In_942);
and U1828 (N_1828,N_181,N_665);
xor U1829 (N_1829,N_1006,N_1034);
or U1830 (N_1830,N_1300,In_232);
nor U1831 (N_1831,N_772,In_1852);
and U1832 (N_1832,In_626,N_1297);
and U1833 (N_1833,N_1163,N_1079);
nand U1834 (N_1834,N_1060,N_1368);
or U1835 (N_1835,N_1439,In_2162);
xnor U1836 (N_1836,N_1409,N_1153);
and U1837 (N_1837,In_1597,N_303);
or U1838 (N_1838,N_748,N_1479);
and U1839 (N_1839,In_47,In_177);
xnor U1840 (N_1840,N_1414,N_1443);
xnor U1841 (N_1841,In_2181,N_1191);
and U1842 (N_1842,In_1280,In_810);
and U1843 (N_1843,In_386,N_1383);
nand U1844 (N_1844,N_129,N_1334);
nor U1845 (N_1845,In_1446,N_1093);
and U1846 (N_1846,N_1152,N_1464);
nand U1847 (N_1847,N_1110,N_337);
xor U1848 (N_1848,In_660,N_1256);
and U1849 (N_1849,N_1447,N_1494);
and U1850 (N_1850,N_1311,N_854);
xor U1851 (N_1851,N_1327,N_1301);
and U1852 (N_1852,N_799,N_567);
and U1853 (N_1853,N_1440,N_1430);
nor U1854 (N_1854,N_918,N_1136);
nor U1855 (N_1855,N_1126,N_832);
or U1856 (N_1856,N_1448,N_1021);
xnor U1857 (N_1857,N_1269,N_934);
or U1858 (N_1858,N_1143,N_1251);
and U1859 (N_1859,N_896,N_1001);
and U1860 (N_1860,N_1452,N_1429);
and U1861 (N_1861,N_1370,N_1446);
xor U1862 (N_1862,N_1486,N_955);
nand U1863 (N_1863,In_1503,N_1454);
nand U1864 (N_1864,N_1069,N_1046);
xor U1865 (N_1865,N_513,In_594);
xor U1866 (N_1866,N_1129,N_697);
nor U1867 (N_1867,In_1291,In_1749);
nor U1868 (N_1868,N_1453,N_1179);
nor U1869 (N_1869,N_1321,N_1291);
or U1870 (N_1870,N_1123,N_909);
and U1871 (N_1871,N_145,N_1224);
nand U1872 (N_1872,N_188,N_1470);
or U1873 (N_1873,N_645,N_1025);
or U1874 (N_1874,N_1442,N_1344);
nor U1875 (N_1875,In_2291,N_1108);
and U1876 (N_1876,N_437,In_293);
and U1877 (N_1877,N_901,N_1073);
nor U1878 (N_1878,N_1474,N_428);
and U1879 (N_1879,N_1185,N_885);
nor U1880 (N_1880,In_1467,N_1352);
nand U1881 (N_1881,In_347,N_1350);
nor U1882 (N_1882,N_1171,N_1020);
nand U1883 (N_1883,N_803,N_1314);
xnor U1884 (N_1884,N_564,N_1182);
nand U1885 (N_1885,In_2165,N_1356);
xor U1886 (N_1886,N_1017,N_1032);
nor U1887 (N_1887,N_1417,N_1390);
and U1888 (N_1888,In_1566,N_1149);
nand U1889 (N_1889,N_1169,In_101);
nor U1890 (N_1890,N_1347,In_1594);
nand U1891 (N_1891,N_1492,N_1331);
and U1892 (N_1892,N_812,In_1535);
nand U1893 (N_1893,In_1838,N_553);
nand U1894 (N_1894,In_1672,N_1226);
nand U1895 (N_1895,N_491,In_1788);
xor U1896 (N_1896,N_796,N_1359);
xor U1897 (N_1897,N_1045,N_1389);
xor U1898 (N_1898,N_1151,N_1213);
nor U1899 (N_1899,In_612,N_952);
xnor U1900 (N_1900,N_1465,N_1489);
and U1901 (N_1901,N_750,N_1192);
and U1902 (N_1902,N_1019,N_1194);
nor U1903 (N_1903,In_1286,N_472);
nand U1904 (N_1904,N_1295,In_1078);
nand U1905 (N_1905,N_1478,N_1132);
nor U1906 (N_1906,In_471,N_777);
xor U1907 (N_1907,In_460,N_754);
or U1908 (N_1908,In_322,N_276);
nor U1909 (N_1909,N_804,N_914);
xor U1910 (N_1910,N_5,N_1436);
and U1911 (N_1911,N_1404,N_1044);
nor U1912 (N_1912,In_305,N_1258);
xnor U1913 (N_1913,In_1026,N_1068);
nand U1914 (N_1914,N_407,N_1208);
and U1915 (N_1915,In_2167,In_547);
xor U1916 (N_1916,N_1433,In_327);
nand U1917 (N_1917,N_792,N_157);
xor U1918 (N_1918,N_487,N_1128);
and U1919 (N_1919,N_1471,N_1139);
xor U1920 (N_1920,N_1296,N_590);
or U1921 (N_1921,N_1221,In_392);
or U1922 (N_1922,N_1048,N_91);
or U1923 (N_1923,N_440,In_1700);
and U1924 (N_1924,N_1190,N_1437);
xnor U1925 (N_1925,N_540,N_994);
and U1926 (N_1926,N_1113,N_1342);
and U1927 (N_1927,N_1340,N_240);
or U1928 (N_1928,In_1895,N_1247);
nor U1929 (N_1929,N_163,In_772);
xor U1930 (N_1930,N_1135,In_2226);
nor U1931 (N_1931,N_7,N_1423);
and U1932 (N_1932,N_878,In_126);
and U1933 (N_1933,N_1333,N_709);
and U1934 (N_1934,N_996,In_661);
nor U1935 (N_1935,N_1211,N_965);
nor U1936 (N_1936,N_1289,N_445);
nor U1937 (N_1937,In_2084,N_1119);
nand U1938 (N_1938,N_1141,N_1095);
and U1939 (N_1939,N_1275,N_1156);
or U1940 (N_1940,N_1148,N_1362);
or U1941 (N_1941,N_1345,N_334);
xor U1942 (N_1942,In_700,In_818);
xor U1943 (N_1943,N_1499,N_1180);
nor U1944 (N_1944,In_2057,N_1329);
nor U1945 (N_1945,N_1038,N_913);
or U1946 (N_1946,In_2456,In_1620);
and U1947 (N_1947,In_153,N_1456);
nand U1948 (N_1948,N_892,N_786);
and U1949 (N_1949,In_1203,N_1286);
xor U1950 (N_1950,N_894,N_1401);
and U1951 (N_1951,N_618,N_1077);
xnor U1952 (N_1952,N_1222,N_521);
xnor U1953 (N_1953,N_879,N_182);
nor U1954 (N_1954,N_661,N_1463);
and U1955 (N_1955,In_1071,N_1363);
nor U1956 (N_1956,N_911,In_2492);
nand U1957 (N_1957,N_1411,N_1215);
and U1958 (N_1958,N_1377,N_1257);
xor U1959 (N_1959,In_74,N_766);
nand U1960 (N_1960,N_1112,N_1360);
nor U1961 (N_1961,N_1467,N_1064);
and U1962 (N_1962,N_1495,N_1076);
xnor U1963 (N_1963,N_13,N_287);
and U1964 (N_1964,N_747,N_817);
xnor U1965 (N_1965,N_1413,In_2109);
or U1966 (N_1966,N_353,In_1814);
nand U1967 (N_1967,In_1508,In_1315);
nand U1968 (N_1968,In_2212,N_1273);
xnor U1969 (N_1969,N_1402,N_1419);
nand U1970 (N_1970,N_1097,N_162);
xnor U1971 (N_1971,N_1266,In_425);
xor U1972 (N_1972,N_782,N_539);
and U1973 (N_1973,N_1282,N_1458);
nor U1974 (N_1974,N_1497,N_1080);
or U1975 (N_1975,N_1328,N_903);
or U1976 (N_1976,N_660,In_2399);
and U1977 (N_1977,In_2095,In_1405);
or U1978 (N_1978,N_755,N_751);
and U1979 (N_1979,N_278,In_975);
xnor U1980 (N_1980,N_727,N_360);
xnor U1981 (N_1981,N_512,N_1099);
nor U1982 (N_1982,N_103,N_1237);
xor U1983 (N_1983,N_827,N_919);
or U1984 (N_1984,In_1270,N_611);
xnor U1985 (N_1985,N_1435,In_941);
nor U1986 (N_1986,N_1117,In_1252);
xor U1987 (N_1987,N_1338,N_1398);
nand U1988 (N_1988,N_1166,In_1115);
and U1989 (N_1989,N_785,N_1188);
nand U1990 (N_1990,N_1315,N_1018);
nor U1991 (N_1991,N_974,N_1361);
xnor U1992 (N_1992,N_228,N_1004);
and U1993 (N_1993,N_1146,N_1122);
nor U1994 (N_1994,N_604,In_237);
nor U1995 (N_1995,In_486,N_609);
or U1996 (N_1996,N_844,N_1145);
nor U1997 (N_1997,N_1412,N_1198);
nand U1998 (N_1998,In_607,N_687);
nor U1999 (N_1999,N_1022,N_1246);
nor U2000 (N_2000,N_1887,N_1779);
xor U2001 (N_2001,N_1738,N_1908);
nand U2002 (N_2002,N_1625,N_1856);
xnor U2003 (N_2003,N_1673,N_1726);
and U2004 (N_2004,N_1796,N_1747);
nor U2005 (N_2005,N_1700,N_1722);
xor U2006 (N_2006,N_1966,N_1637);
and U2007 (N_2007,N_1566,N_1527);
or U2008 (N_2008,N_1716,N_1585);
nand U2009 (N_2009,N_1969,N_1704);
or U2010 (N_2010,N_1827,N_1951);
nand U2011 (N_2011,N_1762,N_1727);
nand U2012 (N_2012,N_1741,N_1694);
or U2013 (N_2013,N_1583,N_1822);
and U2014 (N_2014,N_1780,N_1599);
nor U2015 (N_2015,N_1772,N_1659);
nand U2016 (N_2016,N_1664,N_1981);
nand U2017 (N_2017,N_1924,N_1562);
and U2018 (N_2018,N_1650,N_1874);
or U2019 (N_2019,N_1885,N_1658);
nand U2020 (N_2020,N_1946,N_1857);
xnor U2021 (N_2021,N_1720,N_1802);
xor U2022 (N_2022,N_1701,N_1627);
or U2023 (N_2023,N_1941,N_1850);
or U2024 (N_2024,N_1555,N_1537);
xnor U2025 (N_2025,N_1972,N_1757);
nand U2026 (N_2026,N_1823,N_1524);
xor U2027 (N_2027,N_1962,N_1809);
nand U2028 (N_2028,N_1753,N_1554);
and U2029 (N_2029,N_1645,N_1513);
xnor U2030 (N_2030,N_1996,N_1713);
xor U2031 (N_2031,N_1628,N_1521);
nor U2032 (N_2032,N_1845,N_1774);
xor U2033 (N_2033,N_1884,N_1761);
nor U2034 (N_2034,N_1516,N_1967);
xnor U2035 (N_2035,N_1731,N_1897);
nor U2036 (N_2036,N_1510,N_1913);
nand U2037 (N_2037,N_1719,N_1667);
nor U2038 (N_2038,N_1843,N_1905);
nor U2039 (N_2039,N_1580,N_1935);
xor U2040 (N_2040,N_1961,N_1503);
nor U2041 (N_2041,N_1984,N_1877);
nor U2042 (N_2042,N_1528,N_1564);
nor U2043 (N_2043,N_1797,N_1609);
nor U2044 (N_2044,N_1514,N_1759);
nand U2045 (N_2045,N_1690,N_1640);
or U2046 (N_2046,N_1711,N_1811);
or U2047 (N_2047,N_1771,N_1932);
nand U2048 (N_2048,N_1954,N_1501);
nand U2049 (N_2049,N_1532,N_1922);
xnor U2050 (N_2050,N_1557,N_1600);
nor U2051 (N_2051,N_1914,N_1841);
nor U2052 (N_2052,N_1575,N_1839);
and U2053 (N_2053,N_1910,N_1688);
or U2054 (N_2054,N_1590,N_1512);
or U2055 (N_2055,N_1824,N_1815);
nand U2056 (N_2056,N_1859,N_1565);
and U2057 (N_2057,N_1619,N_1522);
nand U2058 (N_2058,N_1749,N_1531);
or U2059 (N_2059,N_1923,N_1970);
or U2060 (N_2060,N_1876,N_1927);
nor U2061 (N_2061,N_1602,N_1952);
or U2062 (N_2062,N_1587,N_1601);
nor U2063 (N_2063,N_1813,N_1872);
or U2064 (N_2064,N_1655,N_1743);
nand U2065 (N_2065,N_1579,N_1933);
or U2066 (N_2066,N_1681,N_1568);
or U2067 (N_2067,N_1679,N_1612);
nor U2068 (N_2068,N_1763,N_1570);
nor U2069 (N_2069,N_1957,N_1960);
xnor U2070 (N_2070,N_1735,N_1816);
xor U2071 (N_2071,N_1808,N_1789);
nand U2072 (N_2072,N_1948,N_1838);
xnor U2073 (N_2073,N_1896,N_1620);
xnor U2074 (N_2074,N_1770,N_1670);
and U2075 (N_2075,N_1803,N_1760);
or U2076 (N_2076,N_1548,N_1929);
and U2077 (N_2077,N_1710,N_1975);
nand U2078 (N_2078,N_1608,N_1756);
and U2079 (N_2079,N_1781,N_1915);
nand U2080 (N_2080,N_1810,N_1976);
or U2081 (N_2081,N_1665,N_1672);
and U2082 (N_2082,N_1545,N_1862);
nor U2083 (N_2083,N_1663,N_1551);
nor U2084 (N_2084,N_1560,N_1638);
nand U2085 (N_2085,N_1748,N_1881);
xor U2086 (N_2086,N_1733,N_1536);
nor U2087 (N_2087,N_1549,N_1807);
or U2088 (N_2088,N_1798,N_1626);
xnor U2089 (N_2089,N_1879,N_1574);
nor U2090 (N_2090,N_1709,N_1840);
and U2091 (N_2091,N_1993,N_1820);
nor U2092 (N_2092,N_1944,N_1745);
nor U2093 (N_2093,N_1868,N_1692);
xor U2094 (N_2094,N_1894,N_1677);
or U2095 (N_2095,N_1994,N_1606);
nor U2096 (N_2096,N_1805,N_1530);
nand U2097 (N_2097,N_1919,N_1603);
nand U2098 (N_2098,N_1523,N_1624);
nor U2099 (N_2099,N_1890,N_1682);
nor U2100 (N_2100,N_1893,N_1651);
nand U2101 (N_2101,N_1926,N_1949);
nand U2102 (N_2102,N_1518,N_1561);
nor U2103 (N_2103,N_1596,N_1703);
xor U2104 (N_2104,N_1559,N_1942);
nand U2105 (N_2105,N_1552,N_1892);
nor U2106 (N_2106,N_1730,N_1533);
and U2107 (N_2107,N_1714,N_1764);
nand U2108 (N_2108,N_1633,N_1715);
or U2109 (N_2109,N_1988,N_1794);
or U2110 (N_2110,N_1754,N_1869);
and U2111 (N_2111,N_1854,N_1502);
xnor U2112 (N_2112,N_1832,N_1964);
xnor U2113 (N_2113,N_1834,N_1610);
nor U2114 (N_2114,N_1687,N_1669);
and U2115 (N_2115,N_1765,N_1739);
nand U2116 (N_2116,N_1540,N_1736);
nor U2117 (N_2117,N_1595,N_1729);
xnor U2118 (N_2118,N_1649,N_1812);
or U2119 (N_2119,N_1848,N_1788);
nand U2120 (N_2120,N_1911,N_1578);
nand U2121 (N_2121,N_1744,N_1934);
xor U2122 (N_2122,N_1734,N_1642);
and U2123 (N_2123,N_1526,N_1543);
and U2124 (N_2124,N_1630,N_1547);
and U2125 (N_2125,N_1755,N_1577);
nand U2126 (N_2126,N_1616,N_1717);
nor U2127 (N_2127,N_1963,N_1746);
xnor U2128 (N_2128,N_1691,N_1844);
or U2129 (N_2129,N_1953,N_1696);
nor U2130 (N_2130,N_1998,N_1582);
and U2131 (N_2131,N_1978,N_1706);
or U2132 (N_2132,N_1835,N_1847);
and U2133 (N_2133,N_1855,N_1852);
nand U2134 (N_2134,N_1724,N_1842);
or U2135 (N_2135,N_1657,N_1790);
nor U2136 (N_2136,N_1973,N_1916);
nand U2137 (N_2137,N_1680,N_1758);
nand U2138 (N_2138,N_1666,N_1904);
xnor U2139 (N_2139,N_1883,N_1785);
nor U2140 (N_2140,N_1831,N_1992);
and U2141 (N_2141,N_1684,N_1662);
xnor U2142 (N_2142,N_1539,N_1786);
or U2143 (N_2143,N_1907,N_1742);
nor U2144 (N_2144,N_1632,N_1573);
or U2145 (N_2145,N_1817,N_1500);
and U2146 (N_2146,N_1768,N_1902);
and U2147 (N_2147,N_1699,N_1928);
and U2148 (N_2148,N_1604,N_1751);
nor U2149 (N_2149,N_1977,N_1611);
nand U2150 (N_2150,N_1938,N_1886);
xnor U2151 (N_2151,N_1851,N_1593);
xnor U2152 (N_2152,N_1586,N_1517);
nand U2153 (N_2153,N_1828,N_1945);
xnor U2154 (N_2154,N_1678,N_1931);
xor U2155 (N_2155,N_1674,N_1631);
and U2156 (N_2156,N_1728,N_1889);
nor U2157 (N_2157,N_1986,N_1939);
xnor U2158 (N_2158,N_1698,N_1689);
nand U2159 (N_2159,N_1592,N_1507);
nor U2160 (N_2160,N_1544,N_1776);
and U2161 (N_2161,N_1903,N_1656);
and U2162 (N_2162,N_1775,N_1635);
and U2163 (N_2163,N_1778,N_1825);
nor U2164 (N_2164,N_1870,N_1576);
nor U2165 (N_2165,N_1871,N_1535);
xor U2166 (N_2166,N_1980,N_1818);
or U2167 (N_2167,N_1918,N_1792);
and U2168 (N_2168,N_1833,N_1648);
nor U2169 (N_2169,N_1708,N_1959);
nor U2170 (N_2170,N_1519,N_1653);
xnor U2171 (N_2171,N_1644,N_1880);
xor U2172 (N_2172,N_1793,N_1636);
nor U2173 (N_2173,N_1829,N_1861);
and U2174 (N_2174,N_1750,N_1806);
or U2175 (N_2175,N_1605,N_1506);
or U2176 (N_2176,N_1509,N_1542);
nand U2177 (N_2177,N_1752,N_1661);
nor U2178 (N_2178,N_1849,N_1995);
or U2179 (N_2179,N_1652,N_1901);
and U2180 (N_2180,N_1646,N_1925);
nand U2181 (N_2181,N_1623,N_1643);
nor U2182 (N_2182,N_1660,N_1990);
or U2183 (N_2183,N_1511,N_1584);
or U2184 (N_2184,N_1906,N_1801);
or U2185 (N_2185,N_1997,N_1826);
nor U2186 (N_2186,N_1538,N_1529);
xnor U2187 (N_2187,N_1597,N_1819);
xnor U2188 (N_2188,N_1937,N_1615);
and U2189 (N_2189,N_1550,N_1766);
nor U2190 (N_2190,N_1799,N_1899);
nand U2191 (N_2191,N_1891,N_1777);
xnor U2192 (N_2192,N_1675,N_1991);
nor U2193 (N_2193,N_1769,N_1968);
or U2194 (N_2194,N_1863,N_1618);
or U2195 (N_2195,N_1987,N_1591);
and U2196 (N_2196,N_1955,N_1634);
or U2197 (N_2197,N_1846,N_1821);
and U2198 (N_2198,N_1858,N_1695);
nand U2199 (N_2199,N_1940,N_1702);
nand U2200 (N_2200,N_1697,N_1830);
xor U2201 (N_2201,N_1614,N_1740);
nor U2202 (N_2202,N_1971,N_1965);
and U2203 (N_2203,N_1909,N_1685);
xnor U2204 (N_2204,N_1737,N_1718);
and U2205 (N_2205,N_1725,N_1647);
nor U2206 (N_2206,N_1917,N_1804);
and U2207 (N_2207,N_1705,N_1676);
nand U2208 (N_2208,N_1784,N_1505);
xnor U2209 (N_2209,N_1873,N_1867);
nand U2210 (N_2210,N_1882,N_1800);
nor U2211 (N_2211,N_1732,N_1520);
xor U2212 (N_2212,N_1598,N_1629);
or U2213 (N_2213,N_1723,N_1581);
or U2214 (N_2214,N_1693,N_1989);
xor U2215 (N_2215,N_1571,N_1654);
or U2216 (N_2216,N_1546,N_1569);
and U2217 (N_2217,N_1837,N_1508);
or U2218 (N_2218,N_1721,N_1791);
nand U2219 (N_2219,N_1895,N_1920);
or U2220 (N_2220,N_1974,N_1556);
and U2221 (N_2221,N_1898,N_1947);
nor U2222 (N_2222,N_1783,N_1686);
and U2223 (N_2223,N_1567,N_1795);
nor U2224 (N_2224,N_1541,N_1594);
and U2225 (N_2225,N_1588,N_1639);
or U2226 (N_2226,N_1707,N_1860);
or U2227 (N_2227,N_1641,N_1787);
xor U2228 (N_2228,N_1553,N_1558);
nor U2229 (N_2229,N_1982,N_1912);
and U2230 (N_2230,N_1525,N_1613);
xor U2231 (N_2231,N_1875,N_1671);
nand U2232 (N_2232,N_1866,N_1943);
xor U2233 (N_2233,N_1572,N_1683);
xor U2234 (N_2234,N_1864,N_1836);
xor U2235 (N_2235,N_1668,N_1999);
nor U2236 (N_2236,N_1979,N_1563);
and U2237 (N_2237,N_1814,N_1589);
nand U2238 (N_2238,N_1534,N_1956);
and U2239 (N_2239,N_1888,N_1622);
nor U2240 (N_2240,N_1773,N_1930);
and U2241 (N_2241,N_1878,N_1515);
or U2242 (N_2242,N_1617,N_1983);
nor U2243 (N_2243,N_1985,N_1767);
nand U2244 (N_2244,N_1621,N_1865);
or U2245 (N_2245,N_1504,N_1782);
and U2246 (N_2246,N_1712,N_1853);
nand U2247 (N_2247,N_1607,N_1921);
nand U2248 (N_2248,N_1936,N_1958);
nor U2249 (N_2249,N_1950,N_1900);
nor U2250 (N_2250,N_1828,N_1884);
or U2251 (N_2251,N_1612,N_1752);
xor U2252 (N_2252,N_1950,N_1963);
xor U2253 (N_2253,N_1944,N_1833);
and U2254 (N_2254,N_1871,N_1815);
nand U2255 (N_2255,N_1514,N_1590);
nor U2256 (N_2256,N_1898,N_1895);
and U2257 (N_2257,N_1630,N_1791);
nand U2258 (N_2258,N_1873,N_1578);
xnor U2259 (N_2259,N_1811,N_1911);
nand U2260 (N_2260,N_1706,N_1947);
or U2261 (N_2261,N_1501,N_1991);
or U2262 (N_2262,N_1559,N_1563);
and U2263 (N_2263,N_1912,N_1653);
and U2264 (N_2264,N_1508,N_1615);
or U2265 (N_2265,N_1669,N_1570);
nand U2266 (N_2266,N_1740,N_1771);
nor U2267 (N_2267,N_1553,N_1752);
nor U2268 (N_2268,N_1543,N_1688);
nor U2269 (N_2269,N_1576,N_1842);
nand U2270 (N_2270,N_1720,N_1796);
nor U2271 (N_2271,N_1610,N_1813);
or U2272 (N_2272,N_1737,N_1806);
xor U2273 (N_2273,N_1523,N_1659);
nand U2274 (N_2274,N_1929,N_1958);
and U2275 (N_2275,N_1594,N_1648);
nand U2276 (N_2276,N_1685,N_1786);
nor U2277 (N_2277,N_1647,N_1861);
and U2278 (N_2278,N_1818,N_1759);
or U2279 (N_2279,N_1530,N_1794);
nor U2280 (N_2280,N_1666,N_1777);
nand U2281 (N_2281,N_1946,N_1929);
nor U2282 (N_2282,N_1978,N_1872);
or U2283 (N_2283,N_1534,N_1866);
nand U2284 (N_2284,N_1541,N_1960);
or U2285 (N_2285,N_1847,N_1790);
or U2286 (N_2286,N_1929,N_1507);
or U2287 (N_2287,N_1820,N_1575);
xnor U2288 (N_2288,N_1781,N_1965);
or U2289 (N_2289,N_1939,N_1754);
or U2290 (N_2290,N_1719,N_1608);
nand U2291 (N_2291,N_1726,N_1507);
or U2292 (N_2292,N_1524,N_1726);
xnor U2293 (N_2293,N_1677,N_1935);
and U2294 (N_2294,N_1578,N_1614);
xnor U2295 (N_2295,N_1513,N_1516);
xnor U2296 (N_2296,N_1869,N_1993);
or U2297 (N_2297,N_1664,N_1635);
xnor U2298 (N_2298,N_1508,N_1521);
or U2299 (N_2299,N_1767,N_1569);
and U2300 (N_2300,N_1577,N_1588);
or U2301 (N_2301,N_1644,N_1830);
xor U2302 (N_2302,N_1531,N_1796);
and U2303 (N_2303,N_1691,N_1780);
and U2304 (N_2304,N_1693,N_1567);
and U2305 (N_2305,N_1612,N_1843);
and U2306 (N_2306,N_1801,N_1900);
nor U2307 (N_2307,N_1859,N_1879);
nand U2308 (N_2308,N_1503,N_1893);
nor U2309 (N_2309,N_1592,N_1698);
or U2310 (N_2310,N_1581,N_1871);
nand U2311 (N_2311,N_1811,N_1844);
nand U2312 (N_2312,N_1652,N_1640);
and U2313 (N_2313,N_1727,N_1527);
nand U2314 (N_2314,N_1885,N_1863);
and U2315 (N_2315,N_1788,N_1673);
nand U2316 (N_2316,N_1860,N_1561);
or U2317 (N_2317,N_1763,N_1591);
nor U2318 (N_2318,N_1555,N_1530);
nand U2319 (N_2319,N_1987,N_1699);
and U2320 (N_2320,N_1535,N_1916);
and U2321 (N_2321,N_1528,N_1730);
nand U2322 (N_2322,N_1674,N_1679);
and U2323 (N_2323,N_1527,N_1825);
or U2324 (N_2324,N_1798,N_1964);
and U2325 (N_2325,N_1661,N_1743);
nor U2326 (N_2326,N_1912,N_1504);
xor U2327 (N_2327,N_1844,N_1723);
nand U2328 (N_2328,N_1591,N_1854);
nor U2329 (N_2329,N_1688,N_1735);
xor U2330 (N_2330,N_1592,N_1912);
or U2331 (N_2331,N_1822,N_1917);
nor U2332 (N_2332,N_1672,N_1832);
or U2333 (N_2333,N_1876,N_1829);
or U2334 (N_2334,N_1555,N_1698);
nor U2335 (N_2335,N_1656,N_1786);
nand U2336 (N_2336,N_1748,N_1927);
or U2337 (N_2337,N_1901,N_1621);
nor U2338 (N_2338,N_1596,N_1542);
nor U2339 (N_2339,N_1962,N_1966);
nor U2340 (N_2340,N_1876,N_1500);
nor U2341 (N_2341,N_1824,N_1938);
xor U2342 (N_2342,N_1782,N_1764);
nand U2343 (N_2343,N_1717,N_1555);
nor U2344 (N_2344,N_1963,N_1908);
nor U2345 (N_2345,N_1954,N_1883);
nor U2346 (N_2346,N_1667,N_1584);
and U2347 (N_2347,N_1697,N_1840);
or U2348 (N_2348,N_1597,N_1853);
nor U2349 (N_2349,N_1823,N_1626);
nand U2350 (N_2350,N_1766,N_1504);
nor U2351 (N_2351,N_1946,N_1602);
nor U2352 (N_2352,N_1847,N_1763);
and U2353 (N_2353,N_1949,N_1821);
xor U2354 (N_2354,N_1934,N_1817);
or U2355 (N_2355,N_1585,N_1817);
or U2356 (N_2356,N_1950,N_1572);
nor U2357 (N_2357,N_1960,N_1756);
or U2358 (N_2358,N_1685,N_1956);
nand U2359 (N_2359,N_1687,N_1604);
nand U2360 (N_2360,N_1678,N_1764);
nor U2361 (N_2361,N_1885,N_1721);
nand U2362 (N_2362,N_1907,N_1947);
and U2363 (N_2363,N_1523,N_1662);
or U2364 (N_2364,N_1863,N_1802);
and U2365 (N_2365,N_1900,N_1645);
or U2366 (N_2366,N_1637,N_1810);
nor U2367 (N_2367,N_1814,N_1894);
xor U2368 (N_2368,N_1855,N_1547);
and U2369 (N_2369,N_1834,N_1613);
nor U2370 (N_2370,N_1580,N_1572);
nand U2371 (N_2371,N_1758,N_1767);
and U2372 (N_2372,N_1785,N_1803);
nor U2373 (N_2373,N_1771,N_1668);
nor U2374 (N_2374,N_1865,N_1822);
nor U2375 (N_2375,N_1812,N_1834);
or U2376 (N_2376,N_1917,N_1552);
or U2377 (N_2377,N_1848,N_1636);
nor U2378 (N_2378,N_1726,N_1976);
xor U2379 (N_2379,N_1505,N_1773);
xnor U2380 (N_2380,N_1646,N_1946);
or U2381 (N_2381,N_1941,N_1558);
xnor U2382 (N_2382,N_1986,N_1896);
nor U2383 (N_2383,N_1874,N_1638);
and U2384 (N_2384,N_1790,N_1528);
and U2385 (N_2385,N_1661,N_1719);
nor U2386 (N_2386,N_1625,N_1671);
nor U2387 (N_2387,N_1620,N_1553);
xnor U2388 (N_2388,N_1550,N_1966);
and U2389 (N_2389,N_1950,N_1665);
and U2390 (N_2390,N_1926,N_1804);
and U2391 (N_2391,N_1774,N_1513);
nand U2392 (N_2392,N_1647,N_1790);
nand U2393 (N_2393,N_1876,N_1722);
nor U2394 (N_2394,N_1526,N_1885);
nor U2395 (N_2395,N_1555,N_1878);
and U2396 (N_2396,N_1793,N_1770);
xor U2397 (N_2397,N_1667,N_1983);
xnor U2398 (N_2398,N_1669,N_1774);
nor U2399 (N_2399,N_1953,N_1750);
nor U2400 (N_2400,N_1860,N_1542);
nand U2401 (N_2401,N_1540,N_1801);
nand U2402 (N_2402,N_1750,N_1898);
and U2403 (N_2403,N_1805,N_1840);
nor U2404 (N_2404,N_1761,N_1741);
nand U2405 (N_2405,N_1973,N_1997);
xor U2406 (N_2406,N_1596,N_1898);
and U2407 (N_2407,N_1539,N_1908);
xor U2408 (N_2408,N_1588,N_1859);
nor U2409 (N_2409,N_1687,N_1652);
nor U2410 (N_2410,N_1808,N_1625);
xnor U2411 (N_2411,N_1558,N_1696);
nand U2412 (N_2412,N_1623,N_1734);
xor U2413 (N_2413,N_1954,N_1600);
nand U2414 (N_2414,N_1719,N_1834);
nand U2415 (N_2415,N_1844,N_1721);
and U2416 (N_2416,N_1822,N_1963);
and U2417 (N_2417,N_1930,N_1909);
xor U2418 (N_2418,N_1504,N_1922);
nor U2419 (N_2419,N_1771,N_1515);
or U2420 (N_2420,N_1669,N_1620);
or U2421 (N_2421,N_1789,N_1675);
and U2422 (N_2422,N_1910,N_1587);
nand U2423 (N_2423,N_1651,N_1889);
or U2424 (N_2424,N_1533,N_1680);
nand U2425 (N_2425,N_1725,N_1573);
xnor U2426 (N_2426,N_1744,N_1899);
xor U2427 (N_2427,N_1932,N_1968);
nor U2428 (N_2428,N_1828,N_1535);
and U2429 (N_2429,N_1877,N_1966);
xnor U2430 (N_2430,N_1783,N_1794);
nor U2431 (N_2431,N_1782,N_1556);
nor U2432 (N_2432,N_1860,N_1778);
or U2433 (N_2433,N_1525,N_1841);
nor U2434 (N_2434,N_1609,N_1545);
or U2435 (N_2435,N_1869,N_1516);
xor U2436 (N_2436,N_1544,N_1966);
nand U2437 (N_2437,N_1617,N_1549);
and U2438 (N_2438,N_1672,N_1820);
nor U2439 (N_2439,N_1515,N_1840);
xnor U2440 (N_2440,N_1830,N_1801);
xor U2441 (N_2441,N_1951,N_1576);
xnor U2442 (N_2442,N_1882,N_1959);
xnor U2443 (N_2443,N_1734,N_1603);
nor U2444 (N_2444,N_1796,N_1763);
nand U2445 (N_2445,N_1505,N_1781);
nand U2446 (N_2446,N_1677,N_1682);
nand U2447 (N_2447,N_1736,N_1643);
nand U2448 (N_2448,N_1876,N_1891);
nor U2449 (N_2449,N_1941,N_1931);
nand U2450 (N_2450,N_1639,N_1695);
nand U2451 (N_2451,N_1613,N_1510);
xnor U2452 (N_2452,N_1841,N_1876);
xor U2453 (N_2453,N_1994,N_1827);
nor U2454 (N_2454,N_1781,N_1702);
or U2455 (N_2455,N_1550,N_1514);
or U2456 (N_2456,N_1627,N_1940);
nor U2457 (N_2457,N_1739,N_1915);
or U2458 (N_2458,N_1844,N_1898);
nor U2459 (N_2459,N_1704,N_1594);
and U2460 (N_2460,N_1941,N_1731);
and U2461 (N_2461,N_1620,N_1684);
and U2462 (N_2462,N_1617,N_1901);
nand U2463 (N_2463,N_1514,N_1679);
and U2464 (N_2464,N_1731,N_1931);
nor U2465 (N_2465,N_1549,N_1978);
nor U2466 (N_2466,N_1649,N_1655);
xor U2467 (N_2467,N_1701,N_1835);
and U2468 (N_2468,N_1811,N_1895);
nor U2469 (N_2469,N_1956,N_1968);
or U2470 (N_2470,N_1560,N_1915);
xnor U2471 (N_2471,N_1613,N_1859);
and U2472 (N_2472,N_1802,N_1938);
nand U2473 (N_2473,N_1518,N_1754);
xor U2474 (N_2474,N_1505,N_1539);
and U2475 (N_2475,N_1849,N_1639);
or U2476 (N_2476,N_1706,N_1920);
and U2477 (N_2477,N_1534,N_1575);
xnor U2478 (N_2478,N_1942,N_1685);
nor U2479 (N_2479,N_1753,N_1905);
or U2480 (N_2480,N_1510,N_1869);
nor U2481 (N_2481,N_1661,N_1924);
or U2482 (N_2482,N_1594,N_1582);
xnor U2483 (N_2483,N_1605,N_1569);
and U2484 (N_2484,N_1932,N_1500);
and U2485 (N_2485,N_1620,N_1895);
or U2486 (N_2486,N_1918,N_1687);
and U2487 (N_2487,N_1652,N_1917);
and U2488 (N_2488,N_1780,N_1581);
and U2489 (N_2489,N_1743,N_1644);
xnor U2490 (N_2490,N_1715,N_1570);
and U2491 (N_2491,N_1825,N_1523);
nand U2492 (N_2492,N_1723,N_1727);
nand U2493 (N_2493,N_1640,N_1880);
and U2494 (N_2494,N_1826,N_1597);
nor U2495 (N_2495,N_1617,N_1896);
xnor U2496 (N_2496,N_1654,N_1916);
nor U2497 (N_2497,N_1518,N_1683);
xnor U2498 (N_2498,N_1600,N_1689);
xnor U2499 (N_2499,N_1845,N_1638);
nor U2500 (N_2500,N_2163,N_2195);
nand U2501 (N_2501,N_2090,N_2248);
xnor U2502 (N_2502,N_2370,N_2039);
xnor U2503 (N_2503,N_2217,N_2473);
xor U2504 (N_2504,N_2397,N_2491);
nor U2505 (N_2505,N_2308,N_2227);
or U2506 (N_2506,N_2395,N_2459);
and U2507 (N_2507,N_2445,N_2382);
and U2508 (N_2508,N_2185,N_2030);
or U2509 (N_2509,N_2375,N_2447);
nor U2510 (N_2510,N_2086,N_2475);
or U2511 (N_2511,N_2009,N_2012);
nand U2512 (N_2512,N_2063,N_2453);
xor U2513 (N_2513,N_2340,N_2174);
and U2514 (N_2514,N_2189,N_2207);
and U2515 (N_2515,N_2401,N_2178);
or U2516 (N_2516,N_2411,N_2094);
and U2517 (N_2517,N_2436,N_2321);
and U2518 (N_2518,N_2320,N_2241);
nor U2519 (N_2519,N_2372,N_2474);
xor U2520 (N_2520,N_2179,N_2425);
xor U2521 (N_2521,N_2098,N_2097);
or U2522 (N_2522,N_2266,N_2113);
nand U2523 (N_2523,N_2138,N_2298);
and U2524 (N_2524,N_2047,N_2344);
nand U2525 (N_2525,N_2381,N_2256);
and U2526 (N_2526,N_2084,N_2343);
or U2527 (N_2527,N_2018,N_2019);
xnor U2528 (N_2528,N_2299,N_2306);
xnor U2529 (N_2529,N_2017,N_2457);
xor U2530 (N_2530,N_2048,N_2158);
or U2531 (N_2531,N_2262,N_2389);
nor U2532 (N_2532,N_2114,N_2077);
nor U2533 (N_2533,N_2118,N_2192);
or U2534 (N_2534,N_2140,N_2136);
nand U2535 (N_2535,N_2383,N_2269);
nand U2536 (N_2536,N_2250,N_2267);
nand U2537 (N_2537,N_2460,N_2424);
or U2538 (N_2538,N_2186,N_2371);
nor U2539 (N_2539,N_2487,N_2222);
xor U2540 (N_2540,N_2232,N_2280);
and U2541 (N_2541,N_2496,N_2480);
or U2542 (N_2542,N_2304,N_2398);
and U2543 (N_2543,N_2464,N_2007);
and U2544 (N_2544,N_2235,N_2111);
nor U2545 (N_2545,N_2409,N_2127);
nand U2546 (N_2546,N_2323,N_2023);
and U2547 (N_2547,N_2479,N_2054);
nand U2548 (N_2548,N_2287,N_2257);
or U2549 (N_2549,N_2223,N_2025);
nand U2550 (N_2550,N_2446,N_2301);
or U2551 (N_2551,N_2106,N_2384);
nand U2552 (N_2552,N_2218,N_2184);
nor U2553 (N_2553,N_2003,N_2302);
xnor U2554 (N_2554,N_2075,N_2008);
nor U2555 (N_2555,N_2245,N_2193);
or U2556 (N_2556,N_2366,N_2190);
and U2557 (N_2557,N_2043,N_2049);
nand U2558 (N_2558,N_2420,N_2044);
and U2559 (N_2559,N_2000,N_2427);
and U2560 (N_2560,N_2078,N_2388);
nand U2561 (N_2561,N_2068,N_2338);
nand U2562 (N_2562,N_2105,N_2221);
xor U2563 (N_2563,N_2350,N_2351);
nor U2564 (N_2564,N_2021,N_2310);
nor U2565 (N_2565,N_2264,N_2139);
nor U2566 (N_2566,N_2279,N_2191);
nor U2567 (N_2567,N_2405,N_2212);
nor U2568 (N_2568,N_2166,N_2087);
xor U2569 (N_2569,N_2470,N_2426);
xor U2570 (N_2570,N_2334,N_2100);
and U2571 (N_2571,N_2415,N_2249);
xnor U2572 (N_2572,N_2283,N_2064);
nor U2573 (N_2573,N_2325,N_2327);
nor U2574 (N_2574,N_2135,N_2471);
xnor U2575 (N_2575,N_2160,N_2339);
nor U2576 (N_2576,N_2385,N_2169);
or U2577 (N_2577,N_2103,N_2305);
xnor U2578 (N_2578,N_2294,N_2130);
nor U2579 (N_2579,N_2242,N_2418);
nor U2580 (N_2580,N_2159,N_2434);
and U2581 (N_2581,N_2176,N_2076);
and U2582 (N_2582,N_2246,N_2208);
nand U2583 (N_2583,N_2324,N_2499);
nand U2584 (N_2584,N_2380,N_2002);
xor U2585 (N_2585,N_2187,N_2233);
or U2586 (N_2586,N_2303,N_2155);
nand U2587 (N_2587,N_2034,N_2108);
or U2588 (N_2588,N_2161,N_2011);
nand U2589 (N_2589,N_2081,N_2296);
nand U2590 (N_2590,N_2051,N_2033);
or U2591 (N_2591,N_2465,N_2188);
nor U2592 (N_2592,N_2288,N_2326);
xnor U2593 (N_2593,N_2046,N_2229);
or U2594 (N_2594,N_2364,N_2202);
xor U2595 (N_2595,N_2252,N_2337);
xnor U2596 (N_2596,N_2123,N_2069);
xnor U2597 (N_2597,N_2414,N_2170);
nand U2598 (N_2598,N_2201,N_2031);
or U2599 (N_2599,N_2365,N_2316);
nor U2600 (N_2600,N_2148,N_2005);
nor U2601 (N_2601,N_2346,N_2154);
xor U2602 (N_2602,N_2199,N_2482);
nor U2603 (N_2603,N_2276,N_2055);
and U2604 (N_2604,N_2037,N_2092);
nand U2605 (N_2605,N_2416,N_2125);
and U2606 (N_2606,N_2115,N_2029);
xor U2607 (N_2607,N_2355,N_2421);
nor U2608 (N_2608,N_2342,N_2236);
and U2609 (N_2609,N_2374,N_2282);
nand U2610 (N_2610,N_2260,N_2490);
and U2611 (N_2611,N_2444,N_2319);
nand U2612 (N_2612,N_2407,N_2433);
xnor U2613 (N_2613,N_2121,N_2492);
and U2614 (N_2614,N_2391,N_2356);
xor U2615 (N_2615,N_2329,N_2162);
or U2616 (N_2616,N_2057,N_2435);
or U2617 (N_2617,N_2157,N_2335);
and U2618 (N_2618,N_2152,N_2362);
nor U2619 (N_2619,N_2423,N_2172);
and U2620 (N_2620,N_2014,N_2358);
and U2621 (N_2621,N_2165,N_2095);
and U2622 (N_2622,N_2052,N_2476);
xnor U2623 (N_2623,N_2050,N_2110);
or U2624 (N_2624,N_2101,N_2203);
or U2625 (N_2625,N_2104,N_2291);
or U2626 (N_2626,N_2429,N_2489);
or U2627 (N_2627,N_2484,N_2290);
nor U2628 (N_2628,N_2142,N_2378);
or U2629 (N_2629,N_2073,N_2026);
and U2630 (N_2630,N_2001,N_2438);
xor U2631 (N_2631,N_2451,N_2183);
or U2632 (N_2632,N_2058,N_2373);
and U2633 (N_2633,N_2336,N_2137);
nand U2634 (N_2634,N_2428,N_2450);
xnor U2635 (N_2635,N_2454,N_2219);
xor U2636 (N_2636,N_2146,N_2144);
and U2637 (N_2637,N_2281,N_2495);
xnor U2638 (N_2638,N_2419,N_2156);
or U2639 (N_2639,N_2124,N_2486);
nor U2640 (N_2640,N_2056,N_2059);
and U2641 (N_2641,N_2349,N_2079);
nor U2642 (N_2642,N_2348,N_2224);
nor U2643 (N_2643,N_2390,N_2333);
or U2644 (N_2644,N_2175,N_2117);
nand U2645 (N_2645,N_2015,N_2353);
nor U2646 (N_2646,N_2231,N_2149);
xor U2647 (N_2647,N_2237,N_2053);
and U2648 (N_2648,N_2116,N_2258);
nor U2649 (N_2649,N_2399,N_2247);
nor U2650 (N_2650,N_2196,N_2284);
or U2651 (N_2651,N_2234,N_2006);
and U2652 (N_2652,N_2197,N_2387);
nand U2653 (N_2653,N_2147,N_2198);
and U2654 (N_2654,N_2109,N_2472);
or U2655 (N_2655,N_2220,N_2074);
nor U2656 (N_2656,N_2028,N_2261);
nand U2657 (N_2657,N_2107,N_2413);
nor U2658 (N_2658,N_2347,N_2168);
or U2659 (N_2659,N_2263,N_2143);
or U2660 (N_2660,N_2400,N_2455);
nand U2661 (N_2661,N_2060,N_2270);
xnor U2662 (N_2662,N_2027,N_2456);
nor U2663 (N_2663,N_2369,N_2225);
and U2664 (N_2664,N_2357,N_2331);
nor U2665 (N_2665,N_2341,N_2200);
nand U2666 (N_2666,N_2312,N_2478);
and U2667 (N_2667,N_2255,N_2022);
xnor U2668 (N_2668,N_2368,N_2093);
and U2669 (N_2669,N_2412,N_2209);
nor U2670 (N_2670,N_2004,N_2354);
nor U2671 (N_2671,N_2352,N_2439);
and U2672 (N_2672,N_2293,N_2403);
and U2673 (N_2673,N_2361,N_2265);
nand U2674 (N_2674,N_2317,N_2497);
nor U2675 (N_2675,N_2315,N_2036);
and U2676 (N_2676,N_2216,N_2182);
and U2677 (N_2677,N_2448,N_2061);
xor U2678 (N_2678,N_2275,N_2181);
nand U2679 (N_2679,N_2253,N_2286);
nand U2680 (N_2680,N_2089,N_2311);
or U2681 (N_2681,N_2129,N_2243);
and U2682 (N_2682,N_2040,N_2483);
or U2683 (N_2683,N_2498,N_2443);
xnor U2684 (N_2684,N_2430,N_2133);
and U2685 (N_2685,N_2307,N_2041);
and U2686 (N_2686,N_2035,N_2469);
xnor U2687 (N_2687,N_2240,N_2322);
xnor U2688 (N_2688,N_2239,N_2013);
nor U2689 (N_2689,N_2481,N_2145);
xor U2690 (N_2690,N_2102,N_2406);
xnor U2691 (N_2691,N_2259,N_2112);
nor U2692 (N_2692,N_2488,N_2016);
or U2693 (N_2693,N_2210,N_2462);
nand U2694 (N_2694,N_2230,N_2062);
and U2695 (N_2695,N_2318,N_2494);
nor U2696 (N_2696,N_2177,N_2164);
or U2697 (N_2697,N_2379,N_2211);
and U2698 (N_2698,N_2300,N_2330);
nand U2699 (N_2699,N_2417,N_2440);
or U2700 (N_2700,N_2431,N_2134);
and U2701 (N_2701,N_2180,N_2466);
nand U2702 (N_2702,N_2404,N_2402);
and U2703 (N_2703,N_2437,N_2080);
or U2704 (N_2704,N_2238,N_2332);
nor U2705 (N_2705,N_2151,N_2126);
and U2706 (N_2706,N_2070,N_2214);
nor U2707 (N_2707,N_2360,N_2205);
nor U2708 (N_2708,N_2461,N_2032);
nand U2709 (N_2709,N_2268,N_2408);
xor U2710 (N_2710,N_2442,N_2458);
and U2711 (N_2711,N_2167,N_2376);
nand U2712 (N_2712,N_2278,N_2493);
xor U2713 (N_2713,N_2066,N_2432);
nand U2714 (N_2714,N_2010,N_2132);
nand U2715 (N_2715,N_2410,N_2272);
xor U2716 (N_2716,N_2099,N_2254);
nor U2717 (N_2717,N_2083,N_2277);
or U2718 (N_2718,N_2082,N_2122);
and U2719 (N_2719,N_2153,N_2065);
nand U2720 (N_2720,N_2194,N_2273);
nand U2721 (N_2721,N_2088,N_2020);
xnor U2722 (N_2722,N_2314,N_2345);
nand U2723 (N_2723,N_2367,N_2213);
nand U2724 (N_2724,N_2141,N_2422);
nor U2725 (N_2725,N_2071,N_2120);
nand U2726 (N_2726,N_2226,N_2452);
xnor U2727 (N_2727,N_2392,N_2128);
nor U2728 (N_2728,N_2386,N_2171);
nor U2729 (N_2729,N_2441,N_2468);
nor U2730 (N_2730,N_2309,N_2085);
or U2731 (N_2731,N_2067,N_2091);
nand U2732 (N_2732,N_2072,N_2150);
and U2733 (N_2733,N_2215,N_2173);
xnor U2734 (N_2734,N_2024,N_2285);
and U2735 (N_2735,N_2485,N_2449);
and U2736 (N_2736,N_2377,N_2363);
nor U2737 (N_2737,N_2289,N_2396);
or U2738 (N_2738,N_2463,N_2119);
xor U2739 (N_2739,N_2394,N_2477);
nor U2740 (N_2740,N_2131,N_2271);
nor U2741 (N_2741,N_2328,N_2393);
xnor U2742 (N_2742,N_2313,N_2206);
nor U2743 (N_2743,N_2297,N_2045);
nand U2744 (N_2744,N_2467,N_2292);
nand U2745 (N_2745,N_2228,N_2295);
xor U2746 (N_2746,N_2244,N_2096);
nor U2747 (N_2747,N_2042,N_2274);
and U2748 (N_2748,N_2251,N_2359);
or U2749 (N_2749,N_2204,N_2038);
nand U2750 (N_2750,N_2118,N_2046);
xnor U2751 (N_2751,N_2276,N_2250);
nor U2752 (N_2752,N_2249,N_2456);
nor U2753 (N_2753,N_2464,N_2499);
xor U2754 (N_2754,N_2085,N_2452);
or U2755 (N_2755,N_2096,N_2169);
nand U2756 (N_2756,N_2052,N_2283);
or U2757 (N_2757,N_2062,N_2004);
and U2758 (N_2758,N_2035,N_2233);
nand U2759 (N_2759,N_2481,N_2465);
nand U2760 (N_2760,N_2387,N_2093);
xnor U2761 (N_2761,N_2039,N_2223);
or U2762 (N_2762,N_2306,N_2104);
or U2763 (N_2763,N_2252,N_2313);
xor U2764 (N_2764,N_2094,N_2288);
nand U2765 (N_2765,N_2494,N_2224);
or U2766 (N_2766,N_2353,N_2431);
or U2767 (N_2767,N_2309,N_2354);
nor U2768 (N_2768,N_2262,N_2477);
xnor U2769 (N_2769,N_2023,N_2227);
and U2770 (N_2770,N_2170,N_2459);
xor U2771 (N_2771,N_2435,N_2490);
nor U2772 (N_2772,N_2174,N_2484);
nor U2773 (N_2773,N_2095,N_2046);
nor U2774 (N_2774,N_2118,N_2036);
nor U2775 (N_2775,N_2356,N_2378);
or U2776 (N_2776,N_2336,N_2442);
and U2777 (N_2777,N_2262,N_2186);
xnor U2778 (N_2778,N_2455,N_2492);
xor U2779 (N_2779,N_2345,N_2253);
nand U2780 (N_2780,N_2388,N_2246);
nor U2781 (N_2781,N_2092,N_2031);
and U2782 (N_2782,N_2073,N_2362);
nor U2783 (N_2783,N_2101,N_2238);
xnor U2784 (N_2784,N_2017,N_2104);
nor U2785 (N_2785,N_2347,N_2025);
nor U2786 (N_2786,N_2136,N_2155);
or U2787 (N_2787,N_2268,N_2020);
or U2788 (N_2788,N_2420,N_2148);
and U2789 (N_2789,N_2333,N_2164);
nor U2790 (N_2790,N_2254,N_2298);
and U2791 (N_2791,N_2358,N_2003);
and U2792 (N_2792,N_2141,N_2135);
nand U2793 (N_2793,N_2113,N_2224);
nor U2794 (N_2794,N_2149,N_2395);
nand U2795 (N_2795,N_2324,N_2217);
nand U2796 (N_2796,N_2187,N_2455);
xor U2797 (N_2797,N_2338,N_2412);
or U2798 (N_2798,N_2359,N_2265);
and U2799 (N_2799,N_2240,N_2479);
nand U2800 (N_2800,N_2152,N_2183);
nor U2801 (N_2801,N_2247,N_2302);
nand U2802 (N_2802,N_2006,N_2305);
and U2803 (N_2803,N_2307,N_2344);
xnor U2804 (N_2804,N_2447,N_2413);
nand U2805 (N_2805,N_2354,N_2188);
and U2806 (N_2806,N_2062,N_2121);
xor U2807 (N_2807,N_2060,N_2012);
nor U2808 (N_2808,N_2266,N_2156);
nand U2809 (N_2809,N_2324,N_2475);
or U2810 (N_2810,N_2031,N_2246);
nand U2811 (N_2811,N_2176,N_2207);
nand U2812 (N_2812,N_2256,N_2239);
and U2813 (N_2813,N_2333,N_2076);
nor U2814 (N_2814,N_2430,N_2062);
and U2815 (N_2815,N_2121,N_2497);
or U2816 (N_2816,N_2181,N_2425);
nand U2817 (N_2817,N_2218,N_2390);
and U2818 (N_2818,N_2080,N_2367);
and U2819 (N_2819,N_2172,N_2171);
and U2820 (N_2820,N_2288,N_2307);
and U2821 (N_2821,N_2127,N_2174);
nor U2822 (N_2822,N_2310,N_2325);
nor U2823 (N_2823,N_2068,N_2049);
nand U2824 (N_2824,N_2363,N_2093);
xor U2825 (N_2825,N_2289,N_2130);
xor U2826 (N_2826,N_2371,N_2263);
nor U2827 (N_2827,N_2323,N_2146);
and U2828 (N_2828,N_2023,N_2112);
or U2829 (N_2829,N_2304,N_2208);
and U2830 (N_2830,N_2468,N_2137);
nand U2831 (N_2831,N_2208,N_2213);
or U2832 (N_2832,N_2122,N_2226);
nand U2833 (N_2833,N_2216,N_2070);
or U2834 (N_2834,N_2236,N_2426);
nand U2835 (N_2835,N_2308,N_2148);
and U2836 (N_2836,N_2116,N_2056);
and U2837 (N_2837,N_2148,N_2413);
or U2838 (N_2838,N_2007,N_2000);
and U2839 (N_2839,N_2100,N_2476);
or U2840 (N_2840,N_2105,N_2007);
nor U2841 (N_2841,N_2455,N_2134);
xnor U2842 (N_2842,N_2363,N_2025);
and U2843 (N_2843,N_2182,N_2490);
nand U2844 (N_2844,N_2015,N_2074);
and U2845 (N_2845,N_2419,N_2159);
and U2846 (N_2846,N_2396,N_2204);
or U2847 (N_2847,N_2024,N_2461);
and U2848 (N_2848,N_2379,N_2186);
and U2849 (N_2849,N_2067,N_2312);
and U2850 (N_2850,N_2180,N_2283);
nor U2851 (N_2851,N_2015,N_2318);
xor U2852 (N_2852,N_2331,N_2339);
and U2853 (N_2853,N_2458,N_2227);
nand U2854 (N_2854,N_2029,N_2445);
nor U2855 (N_2855,N_2204,N_2343);
xor U2856 (N_2856,N_2060,N_2281);
or U2857 (N_2857,N_2486,N_2079);
and U2858 (N_2858,N_2373,N_2127);
xor U2859 (N_2859,N_2049,N_2066);
nand U2860 (N_2860,N_2015,N_2021);
nor U2861 (N_2861,N_2323,N_2471);
xnor U2862 (N_2862,N_2402,N_2420);
xor U2863 (N_2863,N_2147,N_2010);
xnor U2864 (N_2864,N_2339,N_2002);
nor U2865 (N_2865,N_2085,N_2199);
nor U2866 (N_2866,N_2198,N_2321);
nor U2867 (N_2867,N_2463,N_2054);
xor U2868 (N_2868,N_2186,N_2239);
nand U2869 (N_2869,N_2272,N_2201);
or U2870 (N_2870,N_2385,N_2490);
or U2871 (N_2871,N_2437,N_2146);
or U2872 (N_2872,N_2484,N_2073);
xor U2873 (N_2873,N_2335,N_2099);
or U2874 (N_2874,N_2014,N_2210);
nand U2875 (N_2875,N_2000,N_2155);
or U2876 (N_2876,N_2139,N_2117);
nor U2877 (N_2877,N_2490,N_2068);
nand U2878 (N_2878,N_2060,N_2131);
xor U2879 (N_2879,N_2312,N_2329);
nand U2880 (N_2880,N_2082,N_2274);
and U2881 (N_2881,N_2155,N_2024);
and U2882 (N_2882,N_2493,N_2033);
and U2883 (N_2883,N_2330,N_2413);
nor U2884 (N_2884,N_2184,N_2204);
xnor U2885 (N_2885,N_2288,N_2049);
xnor U2886 (N_2886,N_2229,N_2303);
nand U2887 (N_2887,N_2474,N_2196);
nand U2888 (N_2888,N_2305,N_2208);
nor U2889 (N_2889,N_2461,N_2156);
and U2890 (N_2890,N_2326,N_2307);
nor U2891 (N_2891,N_2473,N_2218);
or U2892 (N_2892,N_2309,N_2326);
xor U2893 (N_2893,N_2493,N_2473);
nand U2894 (N_2894,N_2289,N_2117);
or U2895 (N_2895,N_2010,N_2211);
xor U2896 (N_2896,N_2109,N_2436);
nor U2897 (N_2897,N_2234,N_2241);
and U2898 (N_2898,N_2067,N_2471);
or U2899 (N_2899,N_2119,N_2187);
nor U2900 (N_2900,N_2000,N_2297);
and U2901 (N_2901,N_2430,N_2456);
or U2902 (N_2902,N_2341,N_2040);
xnor U2903 (N_2903,N_2290,N_2494);
or U2904 (N_2904,N_2392,N_2466);
nor U2905 (N_2905,N_2457,N_2319);
nor U2906 (N_2906,N_2108,N_2291);
or U2907 (N_2907,N_2330,N_2087);
or U2908 (N_2908,N_2345,N_2139);
or U2909 (N_2909,N_2187,N_2321);
nand U2910 (N_2910,N_2394,N_2149);
xor U2911 (N_2911,N_2060,N_2102);
nand U2912 (N_2912,N_2454,N_2076);
or U2913 (N_2913,N_2139,N_2002);
nor U2914 (N_2914,N_2266,N_2200);
nand U2915 (N_2915,N_2345,N_2260);
and U2916 (N_2916,N_2288,N_2140);
or U2917 (N_2917,N_2109,N_2473);
nand U2918 (N_2918,N_2440,N_2262);
and U2919 (N_2919,N_2083,N_2299);
xnor U2920 (N_2920,N_2444,N_2391);
nor U2921 (N_2921,N_2467,N_2146);
xor U2922 (N_2922,N_2366,N_2187);
nand U2923 (N_2923,N_2429,N_2030);
and U2924 (N_2924,N_2269,N_2400);
xnor U2925 (N_2925,N_2301,N_2089);
and U2926 (N_2926,N_2252,N_2069);
nor U2927 (N_2927,N_2205,N_2311);
nor U2928 (N_2928,N_2420,N_2434);
xor U2929 (N_2929,N_2110,N_2207);
or U2930 (N_2930,N_2026,N_2219);
and U2931 (N_2931,N_2207,N_2024);
nor U2932 (N_2932,N_2335,N_2254);
xor U2933 (N_2933,N_2465,N_2020);
or U2934 (N_2934,N_2152,N_2030);
nand U2935 (N_2935,N_2044,N_2482);
nand U2936 (N_2936,N_2106,N_2471);
nand U2937 (N_2937,N_2347,N_2366);
and U2938 (N_2938,N_2405,N_2480);
and U2939 (N_2939,N_2308,N_2000);
nor U2940 (N_2940,N_2094,N_2342);
or U2941 (N_2941,N_2341,N_2143);
or U2942 (N_2942,N_2476,N_2480);
xnor U2943 (N_2943,N_2324,N_2207);
nor U2944 (N_2944,N_2312,N_2148);
nor U2945 (N_2945,N_2409,N_2367);
or U2946 (N_2946,N_2477,N_2000);
or U2947 (N_2947,N_2057,N_2254);
nand U2948 (N_2948,N_2172,N_2206);
or U2949 (N_2949,N_2051,N_2345);
nand U2950 (N_2950,N_2063,N_2373);
nand U2951 (N_2951,N_2062,N_2244);
nor U2952 (N_2952,N_2096,N_2466);
xor U2953 (N_2953,N_2208,N_2228);
xnor U2954 (N_2954,N_2424,N_2094);
and U2955 (N_2955,N_2344,N_2168);
or U2956 (N_2956,N_2372,N_2406);
nand U2957 (N_2957,N_2440,N_2236);
xor U2958 (N_2958,N_2475,N_2299);
or U2959 (N_2959,N_2245,N_2053);
xor U2960 (N_2960,N_2192,N_2441);
nand U2961 (N_2961,N_2133,N_2041);
or U2962 (N_2962,N_2374,N_2010);
and U2963 (N_2963,N_2102,N_2139);
nor U2964 (N_2964,N_2388,N_2223);
nand U2965 (N_2965,N_2099,N_2077);
nand U2966 (N_2966,N_2463,N_2313);
nand U2967 (N_2967,N_2006,N_2358);
nand U2968 (N_2968,N_2264,N_2175);
nand U2969 (N_2969,N_2269,N_2167);
nand U2970 (N_2970,N_2346,N_2258);
xor U2971 (N_2971,N_2344,N_2113);
and U2972 (N_2972,N_2467,N_2340);
nand U2973 (N_2973,N_2350,N_2302);
nor U2974 (N_2974,N_2418,N_2054);
nor U2975 (N_2975,N_2165,N_2378);
nor U2976 (N_2976,N_2329,N_2441);
nor U2977 (N_2977,N_2138,N_2398);
or U2978 (N_2978,N_2401,N_2447);
or U2979 (N_2979,N_2300,N_2161);
xnor U2980 (N_2980,N_2372,N_2117);
xor U2981 (N_2981,N_2364,N_2023);
or U2982 (N_2982,N_2264,N_2052);
xor U2983 (N_2983,N_2493,N_2108);
nand U2984 (N_2984,N_2475,N_2270);
xor U2985 (N_2985,N_2055,N_2243);
or U2986 (N_2986,N_2234,N_2438);
or U2987 (N_2987,N_2146,N_2264);
nand U2988 (N_2988,N_2048,N_2357);
nand U2989 (N_2989,N_2280,N_2097);
and U2990 (N_2990,N_2175,N_2054);
and U2991 (N_2991,N_2226,N_2323);
xnor U2992 (N_2992,N_2459,N_2499);
nor U2993 (N_2993,N_2196,N_2433);
nand U2994 (N_2994,N_2478,N_2071);
nor U2995 (N_2995,N_2018,N_2408);
and U2996 (N_2996,N_2061,N_2144);
or U2997 (N_2997,N_2444,N_2288);
or U2998 (N_2998,N_2265,N_2398);
xnor U2999 (N_2999,N_2096,N_2463);
nor U3000 (N_3000,N_2800,N_2538);
xor U3001 (N_3001,N_2631,N_2524);
and U3002 (N_3002,N_2956,N_2887);
xor U3003 (N_3003,N_2544,N_2862);
xor U3004 (N_3004,N_2643,N_2733);
or U3005 (N_3005,N_2965,N_2689);
nand U3006 (N_3006,N_2658,N_2760);
and U3007 (N_3007,N_2575,N_2685);
nand U3008 (N_3008,N_2703,N_2645);
or U3009 (N_3009,N_2619,N_2755);
nand U3010 (N_3010,N_2845,N_2701);
and U3011 (N_3011,N_2963,N_2940);
nand U3012 (N_3012,N_2667,N_2769);
nand U3013 (N_3013,N_2780,N_2641);
xor U3014 (N_3014,N_2736,N_2856);
nand U3015 (N_3015,N_2825,N_2992);
and U3016 (N_3016,N_2787,N_2717);
and U3017 (N_3017,N_2713,N_2712);
and U3018 (N_3018,N_2605,N_2706);
nor U3019 (N_3019,N_2982,N_2718);
or U3020 (N_3020,N_2593,N_2743);
nand U3021 (N_3021,N_2900,N_2528);
nor U3022 (N_3022,N_2796,N_2813);
nand U3023 (N_3023,N_2836,N_2700);
or U3024 (N_3024,N_2579,N_2727);
nor U3025 (N_3025,N_2967,N_2596);
xor U3026 (N_3026,N_2625,N_2566);
xor U3027 (N_3027,N_2832,N_2642);
nand U3028 (N_3028,N_2680,N_2971);
or U3029 (N_3029,N_2931,N_2547);
or U3030 (N_3030,N_2920,N_2728);
nand U3031 (N_3031,N_2790,N_2635);
and U3032 (N_3032,N_2895,N_2758);
or U3033 (N_3033,N_2879,N_2565);
or U3034 (N_3034,N_2501,N_2710);
nand U3035 (N_3035,N_2716,N_2788);
nand U3036 (N_3036,N_2721,N_2617);
nand U3037 (N_3037,N_2610,N_2725);
and U3038 (N_3038,N_2823,N_2724);
and U3039 (N_3039,N_2909,N_2919);
xnor U3040 (N_3040,N_2898,N_2863);
xor U3041 (N_3041,N_2936,N_2673);
xnor U3042 (N_3042,N_2616,N_2866);
nand U3043 (N_3043,N_2508,N_2629);
nand U3044 (N_3044,N_2542,N_2814);
xor U3045 (N_3045,N_2607,N_2562);
nor U3046 (N_3046,N_2976,N_2918);
xnor U3047 (N_3047,N_2742,N_2648);
or U3048 (N_3048,N_2774,N_2653);
nor U3049 (N_3049,N_2821,N_2762);
nand U3050 (N_3050,N_2699,N_2798);
and U3051 (N_3051,N_2763,N_2860);
nor U3052 (N_3052,N_2666,N_2595);
and U3053 (N_3053,N_2938,N_2600);
xor U3054 (N_3054,N_2684,N_2877);
nand U3055 (N_3055,N_2513,N_2626);
nand U3056 (N_3056,N_2922,N_2584);
nor U3057 (N_3057,N_2585,N_2882);
nand U3058 (N_3058,N_2531,N_2805);
and U3059 (N_3059,N_2750,N_2886);
nor U3060 (N_3060,N_2812,N_2880);
nor U3061 (N_3061,N_2915,N_2799);
or U3062 (N_3062,N_2789,N_2709);
xor U3063 (N_3063,N_2687,N_2551);
and U3064 (N_3064,N_2896,N_2606);
nand U3065 (N_3065,N_2988,N_2776);
nand U3066 (N_3066,N_2857,N_2534);
nor U3067 (N_3067,N_2502,N_2654);
nor U3068 (N_3068,N_2615,N_2694);
nor U3069 (N_3069,N_2775,N_2591);
or U3070 (N_3070,N_2794,N_2726);
nor U3071 (N_3071,N_2949,N_2783);
and U3072 (N_3072,N_2809,N_2644);
and U3073 (N_3073,N_2894,N_2671);
xnor U3074 (N_3074,N_2791,N_2878);
nand U3075 (N_3075,N_2681,N_2530);
nor U3076 (N_3076,N_2737,N_2628);
nor U3077 (N_3077,N_2603,N_2852);
xor U3078 (N_3078,N_2969,N_2651);
nor U3079 (N_3079,N_2580,N_2601);
and U3080 (N_3080,N_2810,N_2808);
nor U3081 (N_3081,N_2933,N_2636);
nand U3082 (N_3082,N_2831,N_2885);
nor U3083 (N_3083,N_2686,N_2868);
and U3084 (N_3084,N_2911,N_2980);
and U3085 (N_3085,N_2883,N_2512);
nand U3086 (N_3086,N_2589,N_2568);
xor U3087 (N_3087,N_2577,N_2683);
nand U3088 (N_3088,N_2989,N_2582);
nor U3089 (N_3089,N_2830,N_2874);
and U3090 (N_3090,N_2731,N_2545);
and U3091 (N_3091,N_2520,N_2848);
xnor U3092 (N_3092,N_2509,N_2739);
and U3093 (N_3093,N_2676,N_2663);
xor U3094 (N_3094,N_2650,N_2637);
xnor U3095 (N_3095,N_2844,N_2792);
nor U3096 (N_3096,N_2897,N_2881);
nor U3097 (N_3097,N_2732,N_2981);
nor U3098 (N_3098,N_2914,N_2952);
nor U3099 (N_3099,N_2795,N_2533);
nand U3100 (N_3100,N_2899,N_2510);
xor U3101 (N_3101,N_2839,N_2818);
or U3102 (N_3102,N_2957,N_2893);
or U3103 (N_3103,N_2801,N_2527);
or U3104 (N_3104,N_2536,N_2675);
nor U3105 (N_3105,N_2782,N_2829);
nand U3106 (N_3106,N_2926,N_2850);
nor U3107 (N_3107,N_2745,N_2738);
nand U3108 (N_3108,N_2872,N_2968);
nand U3109 (N_3109,N_2962,N_2656);
xor U3110 (N_3110,N_2778,N_2958);
nand U3111 (N_3111,N_2554,N_2855);
nand U3112 (N_3112,N_2708,N_2902);
nand U3113 (N_3113,N_2715,N_2768);
or U3114 (N_3114,N_2630,N_2993);
and U3115 (N_3115,N_2835,N_2574);
and U3116 (N_3116,N_2678,N_2822);
or U3117 (N_3117,N_2741,N_2537);
and U3118 (N_3118,N_2837,N_2867);
xor U3119 (N_3119,N_2834,N_2945);
and U3120 (N_3120,N_2854,N_2532);
or U3121 (N_3121,N_2786,N_2655);
xor U3122 (N_3122,N_2811,N_2983);
nand U3123 (N_3123,N_2702,N_2613);
nand U3124 (N_3124,N_2623,N_2500);
xnor U3125 (N_3125,N_2652,N_2638);
nor U3126 (N_3126,N_2588,N_2679);
nand U3127 (N_3127,N_2779,N_2908);
nor U3128 (N_3128,N_2549,N_2657);
and U3129 (N_3129,N_2759,N_2573);
xor U3130 (N_3130,N_2592,N_2870);
nor U3131 (N_3131,N_2504,N_2752);
xor U3132 (N_3132,N_2590,N_2930);
xor U3133 (N_3133,N_2696,N_2548);
and U3134 (N_3134,N_2747,N_2973);
and U3135 (N_3135,N_2987,N_2569);
xnor U3136 (N_3136,N_2546,N_2691);
nand U3137 (N_3137,N_2515,N_2978);
and U3138 (N_3138,N_2711,N_2541);
or U3139 (N_3139,N_2797,N_2729);
nor U3140 (N_3140,N_2744,N_2633);
or U3141 (N_3141,N_2612,N_2517);
and U3142 (N_3142,N_2511,N_2543);
nand U3143 (N_3143,N_2570,N_2556);
or U3144 (N_3144,N_2889,N_2979);
nand U3145 (N_3145,N_2851,N_2820);
or U3146 (N_3146,N_2806,N_2526);
or U3147 (N_3147,N_2984,N_2888);
or U3148 (N_3148,N_2925,N_2996);
or U3149 (N_3149,N_2853,N_2514);
or U3150 (N_3150,N_2695,N_2561);
and U3151 (N_3151,N_2507,N_2660);
xor U3152 (N_3152,N_2819,N_2905);
or U3153 (N_3153,N_2998,N_2773);
nor U3154 (N_3154,N_2505,N_2519);
xnor U3155 (N_3155,N_2594,N_2757);
nand U3156 (N_3156,N_2999,N_2772);
or U3157 (N_3157,N_2917,N_2661);
nor U3158 (N_3158,N_2581,N_2597);
xor U3159 (N_3159,N_2693,N_2720);
nor U3160 (N_3160,N_2766,N_2559);
xor U3161 (N_3161,N_2910,N_2884);
xor U3162 (N_3162,N_2698,N_2781);
nand U3163 (N_3163,N_2913,N_2751);
nand U3164 (N_3164,N_2664,N_2826);
xnor U3165 (N_3165,N_2934,N_2506);
xnor U3166 (N_3166,N_2640,N_2639);
nand U3167 (N_3167,N_2662,N_2578);
and U3168 (N_3168,N_2932,N_2690);
xor U3169 (N_3169,N_2997,N_2903);
and U3170 (N_3170,N_2525,N_2959);
nand U3171 (N_3171,N_2828,N_2955);
and U3172 (N_3172,N_2602,N_2954);
and U3173 (N_3173,N_2682,N_2785);
and U3174 (N_3174,N_2516,N_2555);
and U3175 (N_3175,N_2618,N_2622);
nor U3176 (N_3176,N_2912,N_2847);
and U3177 (N_3177,N_2807,N_2771);
nor U3178 (N_3178,N_2608,N_2924);
or U3179 (N_3179,N_2990,N_2707);
and U3180 (N_3180,N_2539,N_2767);
xor U3181 (N_3181,N_2859,N_2705);
nor U3182 (N_3182,N_2535,N_2986);
xor U3183 (N_3183,N_2649,N_2817);
nor U3184 (N_3184,N_2598,N_2892);
nor U3185 (N_3185,N_2827,N_2632);
nor U3186 (N_3186,N_2740,N_2951);
xnor U3187 (N_3187,N_2599,N_2974);
or U3188 (N_3188,N_2558,N_2761);
and U3189 (N_3189,N_2961,N_2670);
nand U3190 (N_3190,N_2692,N_2947);
xor U3191 (N_3191,N_2704,N_2864);
nand U3192 (N_3192,N_2875,N_2935);
and U3193 (N_3193,N_2975,N_2735);
and U3194 (N_3194,N_2557,N_2804);
or U3195 (N_3195,N_2677,N_2904);
and U3196 (N_3196,N_2521,N_2972);
xnor U3197 (N_3197,N_2764,N_2722);
xor U3198 (N_3198,N_2672,N_2846);
nor U3199 (N_3199,N_2901,N_2995);
nor U3200 (N_3200,N_2560,N_2966);
nand U3201 (N_3201,N_2991,N_2576);
xor U3202 (N_3202,N_2503,N_2833);
nor U3203 (N_3203,N_2840,N_2553);
nor U3204 (N_3204,N_2939,N_2550);
xnor U3205 (N_3205,N_2907,N_2937);
and U3206 (N_3206,N_2540,N_2611);
xor U3207 (N_3207,N_2838,N_2841);
and U3208 (N_3208,N_2803,N_2923);
and U3209 (N_3209,N_2770,N_2953);
or U3210 (N_3210,N_2964,N_2793);
and U3211 (N_3211,N_2994,N_2890);
xnor U3212 (N_3212,N_2824,N_2858);
nand U3213 (N_3213,N_2753,N_2916);
nor U3214 (N_3214,N_2564,N_2624);
nand U3215 (N_3215,N_2604,N_2518);
xnor U3216 (N_3216,N_2950,N_2929);
or U3217 (N_3217,N_2960,N_2620);
nor U3218 (N_3218,N_2688,N_2567);
and U3219 (N_3219,N_2843,N_2665);
nand U3220 (N_3220,N_2754,N_2849);
xor U3221 (N_3221,N_2946,N_2944);
xnor U3222 (N_3222,N_2869,N_2861);
nand U3223 (N_3223,N_2719,N_2765);
and U3224 (N_3224,N_2627,N_2668);
and U3225 (N_3225,N_2523,N_2777);
or U3226 (N_3226,N_2784,N_2746);
or U3227 (N_3227,N_2583,N_2614);
nor U3228 (N_3228,N_2587,N_2977);
and U3229 (N_3229,N_2943,N_2802);
nand U3230 (N_3230,N_2927,N_2646);
and U3231 (N_3231,N_2970,N_2873);
nand U3232 (N_3232,N_2876,N_2669);
xnor U3233 (N_3233,N_2748,N_2723);
nor U3234 (N_3234,N_2634,N_2815);
or U3235 (N_3235,N_2891,N_2871);
and U3236 (N_3236,N_2571,N_2942);
and U3237 (N_3237,N_2697,N_2714);
and U3238 (N_3238,N_2572,N_2609);
nor U3239 (N_3239,N_2659,N_2730);
nand U3240 (N_3240,N_2529,N_2948);
nor U3241 (N_3241,N_2816,N_2941);
or U3242 (N_3242,N_2563,N_2621);
nand U3243 (N_3243,N_2906,N_2749);
nor U3244 (N_3244,N_2647,N_2674);
or U3245 (N_3245,N_2522,N_2985);
nand U3246 (N_3246,N_2921,N_2734);
or U3247 (N_3247,N_2552,N_2586);
xor U3248 (N_3248,N_2842,N_2865);
nand U3249 (N_3249,N_2928,N_2756);
xnor U3250 (N_3250,N_2598,N_2537);
or U3251 (N_3251,N_2912,N_2506);
or U3252 (N_3252,N_2733,N_2911);
nand U3253 (N_3253,N_2512,N_2889);
nor U3254 (N_3254,N_2862,N_2536);
nor U3255 (N_3255,N_2961,N_2885);
xor U3256 (N_3256,N_2513,N_2752);
or U3257 (N_3257,N_2558,N_2534);
nand U3258 (N_3258,N_2884,N_2810);
nor U3259 (N_3259,N_2561,N_2757);
xor U3260 (N_3260,N_2986,N_2601);
xor U3261 (N_3261,N_2586,N_2978);
and U3262 (N_3262,N_2995,N_2822);
xor U3263 (N_3263,N_2746,N_2801);
nand U3264 (N_3264,N_2710,N_2768);
or U3265 (N_3265,N_2733,N_2772);
xor U3266 (N_3266,N_2549,N_2523);
nor U3267 (N_3267,N_2587,N_2963);
and U3268 (N_3268,N_2926,N_2666);
nor U3269 (N_3269,N_2650,N_2516);
and U3270 (N_3270,N_2630,N_2566);
and U3271 (N_3271,N_2565,N_2656);
or U3272 (N_3272,N_2784,N_2843);
nand U3273 (N_3273,N_2978,N_2794);
xor U3274 (N_3274,N_2626,N_2899);
or U3275 (N_3275,N_2822,N_2879);
xnor U3276 (N_3276,N_2526,N_2543);
nand U3277 (N_3277,N_2916,N_2979);
and U3278 (N_3278,N_2629,N_2857);
nor U3279 (N_3279,N_2861,N_2712);
nor U3280 (N_3280,N_2780,N_2516);
xor U3281 (N_3281,N_2847,N_2675);
xor U3282 (N_3282,N_2931,N_2836);
xor U3283 (N_3283,N_2794,N_2981);
and U3284 (N_3284,N_2817,N_2943);
or U3285 (N_3285,N_2637,N_2799);
and U3286 (N_3286,N_2719,N_2747);
nand U3287 (N_3287,N_2998,N_2978);
or U3288 (N_3288,N_2854,N_2689);
and U3289 (N_3289,N_2913,N_2932);
or U3290 (N_3290,N_2519,N_2897);
and U3291 (N_3291,N_2643,N_2655);
nand U3292 (N_3292,N_2527,N_2867);
or U3293 (N_3293,N_2862,N_2817);
or U3294 (N_3294,N_2574,N_2637);
and U3295 (N_3295,N_2881,N_2813);
nor U3296 (N_3296,N_2771,N_2975);
nand U3297 (N_3297,N_2603,N_2740);
nand U3298 (N_3298,N_2729,N_2553);
or U3299 (N_3299,N_2700,N_2707);
or U3300 (N_3300,N_2765,N_2553);
and U3301 (N_3301,N_2707,N_2639);
or U3302 (N_3302,N_2826,N_2769);
xnor U3303 (N_3303,N_2651,N_2662);
nor U3304 (N_3304,N_2604,N_2834);
and U3305 (N_3305,N_2902,N_2985);
and U3306 (N_3306,N_2691,N_2540);
nor U3307 (N_3307,N_2532,N_2585);
nand U3308 (N_3308,N_2824,N_2909);
nand U3309 (N_3309,N_2715,N_2873);
nor U3310 (N_3310,N_2774,N_2792);
xnor U3311 (N_3311,N_2898,N_2793);
and U3312 (N_3312,N_2741,N_2792);
xor U3313 (N_3313,N_2524,N_2853);
nor U3314 (N_3314,N_2913,N_2520);
nor U3315 (N_3315,N_2639,N_2822);
or U3316 (N_3316,N_2851,N_2540);
and U3317 (N_3317,N_2535,N_2769);
nand U3318 (N_3318,N_2806,N_2963);
or U3319 (N_3319,N_2896,N_2628);
nand U3320 (N_3320,N_2743,N_2851);
xor U3321 (N_3321,N_2926,N_2728);
or U3322 (N_3322,N_2697,N_2541);
and U3323 (N_3323,N_2909,N_2992);
and U3324 (N_3324,N_2540,N_2863);
nand U3325 (N_3325,N_2678,N_2788);
nand U3326 (N_3326,N_2671,N_2945);
or U3327 (N_3327,N_2906,N_2704);
nor U3328 (N_3328,N_2580,N_2893);
and U3329 (N_3329,N_2512,N_2926);
xor U3330 (N_3330,N_2962,N_2754);
or U3331 (N_3331,N_2999,N_2689);
and U3332 (N_3332,N_2752,N_2881);
or U3333 (N_3333,N_2643,N_2749);
xnor U3334 (N_3334,N_2633,N_2662);
xor U3335 (N_3335,N_2942,N_2509);
nand U3336 (N_3336,N_2515,N_2970);
nor U3337 (N_3337,N_2817,N_2973);
xor U3338 (N_3338,N_2823,N_2976);
and U3339 (N_3339,N_2980,N_2892);
and U3340 (N_3340,N_2796,N_2703);
or U3341 (N_3341,N_2790,N_2598);
and U3342 (N_3342,N_2586,N_2659);
and U3343 (N_3343,N_2539,N_2867);
or U3344 (N_3344,N_2643,N_2806);
and U3345 (N_3345,N_2953,N_2686);
or U3346 (N_3346,N_2526,N_2748);
xnor U3347 (N_3347,N_2566,N_2728);
and U3348 (N_3348,N_2579,N_2836);
xnor U3349 (N_3349,N_2694,N_2738);
and U3350 (N_3350,N_2740,N_2555);
nor U3351 (N_3351,N_2785,N_2930);
nand U3352 (N_3352,N_2595,N_2943);
nand U3353 (N_3353,N_2500,N_2643);
or U3354 (N_3354,N_2677,N_2986);
nor U3355 (N_3355,N_2975,N_2951);
nand U3356 (N_3356,N_2610,N_2809);
and U3357 (N_3357,N_2610,N_2788);
nor U3358 (N_3358,N_2897,N_2899);
and U3359 (N_3359,N_2635,N_2960);
nand U3360 (N_3360,N_2802,N_2593);
and U3361 (N_3361,N_2593,N_2645);
nand U3362 (N_3362,N_2718,N_2880);
nor U3363 (N_3363,N_2990,N_2704);
xnor U3364 (N_3364,N_2761,N_2903);
nor U3365 (N_3365,N_2672,N_2860);
xnor U3366 (N_3366,N_2525,N_2817);
nand U3367 (N_3367,N_2770,N_2650);
or U3368 (N_3368,N_2624,N_2859);
and U3369 (N_3369,N_2544,N_2692);
nor U3370 (N_3370,N_2964,N_2828);
nor U3371 (N_3371,N_2908,N_2853);
xor U3372 (N_3372,N_2990,N_2538);
nor U3373 (N_3373,N_2739,N_2850);
or U3374 (N_3374,N_2939,N_2779);
and U3375 (N_3375,N_2799,N_2508);
nor U3376 (N_3376,N_2728,N_2895);
xnor U3377 (N_3377,N_2997,N_2768);
nor U3378 (N_3378,N_2822,N_2938);
nand U3379 (N_3379,N_2875,N_2909);
nand U3380 (N_3380,N_2585,N_2806);
xor U3381 (N_3381,N_2650,N_2929);
or U3382 (N_3382,N_2753,N_2996);
xnor U3383 (N_3383,N_2617,N_2946);
nor U3384 (N_3384,N_2954,N_2653);
nand U3385 (N_3385,N_2678,N_2863);
or U3386 (N_3386,N_2572,N_2684);
nand U3387 (N_3387,N_2842,N_2731);
xor U3388 (N_3388,N_2867,N_2519);
or U3389 (N_3389,N_2689,N_2840);
or U3390 (N_3390,N_2974,N_2546);
and U3391 (N_3391,N_2608,N_2826);
xor U3392 (N_3392,N_2712,N_2826);
nand U3393 (N_3393,N_2994,N_2522);
or U3394 (N_3394,N_2581,N_2867);
and U3395 (N_3395,N_2520,N_2700);
nor U3396 (N_3396,N_2951,N_2513);
or U3397 (N_3397,N_2734,N_2747);
nand U3398 (N_3398,N_2781,N_2533);
or U3399 (N_3399,N_2554,N_2965);
and U3400 (N_3400,N_2510,N_2839);
nor U3401 (N_3401,N_2807,N_2911);
and U3402 (N_3402,N_2950,N_2775);
nor U3403 (N_3403,N_2994,N_2746);
or U3404 (N_3404,N_2612,N_2939);
nor U3405 (N_3405,N_2725,N_2593);
nor U3406 (N_3406,N_2902,N_2516);
nand U3407 (N_3407,N_2591,N_2615);
xor U3408 (N_3408,N_2924,N_2516);
xor U3409 (N_3409,N_2543,N_2704);
nand U3410 (N_3410,N_2877,N_2553);
nand U3411 (N_3411,N_2604,N_2944);
and U3412 (N_3412,N_2874,N_2666);
or U3413 (N_3413,N_2739,N_2875);
xor U3414 (N_3414,N_2518,N_2749);
xnor U3415 (N_3415,N_2678,N_2587);
or U3416 (N_3416,N_2720,N_2800);
nand U3417 (N_3417,N_2768,N_2572);
nand U3418 (N_3418,N_2763,N_2983);
nand U3419 (N_3419,N_2542,N_2571);
nand U3420 (N_3420,N_2881,N_2747);
xor U3421 (N_3421,N_2537,N_2965);
nor U3422 (N_3422,N_2843,N_2934);
nand U3423 (N_3423,N_2844,N_2527);
or U3424 (N_3424,N_2850,N_2833);
nor U3425 (N_3425,N_2792,N_2672);
nor U3426 (N_3426,N_2786,N_2903);
or U3427 (N_3427,N_2894,N_2561);
xnor U3428 (N_3428,N_2558,N_2798);
or U3429 (N_3429,N_2876,N_2832);
xnor U3430 (N_3430,N_2976,N_2705);
or U3431 (N_3431,N_2600,N_2994);
nand U3432 (N_3432,N_2887,N_2550);
or U3433 (N_3433,N_2656,N_2529);
or U3434 (N_3434,N_2997,N_2731);
nand U3435 (N_3435,N_2583,N_2565);
nor U3436 (N_3436,N_2977,N_2785);
nand U3437 (N_3437,N_2548,N_2898);
or U3438 (N_3438,N_2991,N_2727);
xor U3439 (N_3439,N_2724,N_2754);
nor U3440 (N_3440,N_2660,N_2662);
and U3441 (N_3441,N_2795,N_2742);
nor U3442 (N_3442,N_2787,N_2558);
and U3443 (N_3443,N_2715,N_2799);
nand U3444 (N_3444,N_2524,N_2620);
or U3445 (N_3445,N_2796,N_2525);
xnor U3446 (N_3446,N_2515,N_2911);
and U3447 (N_3447,N_2794,N_2995);
and U3448 (N_3448,N_2950,N_2919);
and U3449 (N_3449,N_2781,N_2830);
xnor U3450 (N_3450,N_2676,N_2731);
nor U3451 (N_3451,N_2972,N_2894);
xnor U3452 (N_3452,N_2624,N_2690);
or U3453 (N_3453,N_2545,N_2751);
or U3454 (N_3454,N_2710,N_2953);
or U3455 (N_3455,N_2976,N_2586);
and U3456 (N_3456,N_2559,N_2792);
nand U3457 (N_3457,N_2852,N_2961);
or U3458 (N_3458,N_2783,N_2799);
xor U3459 (N_3459,N_2995,N_2725);
nand U3460 (N_3460,N_2558,N_2692);
or U3461 (N_3461,N_2964,N_2977);
xnor U3462 (N_3462,N_2568,N_2577);
and U3463 (N_3463,N_2751,N_2645);
and U3464 (N_3464,N_2671,N_2939);
and U3465 (N_3465,N_2797,N_2842);
and U3466 (N_3466,N_2579,N_2707);
and U3467 (N_3467,N_2897,N_2590);
or U3468 (N_3468,N_2770,N_2977);
and U3469 (N_3469,N_2916,N_2840);
or U3470 (N_3470,N_2671,N_2804);
nand U3471 (N_3471,N_2547,N_2558);
nand U3472 (N_3472,N_2502,N_2632);
or U3473 (N_3473,N_2971,N_2796);
or U3474 (N_3474,N_2651,N_2881);
or U3475 (N_3475,N_2895,N_2518);
xnor U3476 (N_3476,N_2656,N_2954);
and U3477 (N_3477,N_2776,N_2882);
nor U3478 (N_3478,N_2898,N_2769);
nand U3479 (N_3479,N_2611,N_2727);
or U3480 (N_3480,N_2910,N_2902);
nor U3481 (N_3481,N_2731,N_2736);
and U3482 (N_3482,N_2633,N_2947);
and U3483 (N_3483,N_2610,N_2915);
or U3484 (N_3484,N_2721,N_2818);
xnor U3485 (N_3485,N_2621,N_2737);
nand U3486 (N_3486,N_2883,N_2854);
and U3487 (N_3487,N_2758,N_2662);
and U3488 (N_3488,N_2660,N_2519);
xnor U3489 (N_3489,N_2894,N_2793);
nor U3490 (N_3490,N_2538,N_2654);
nor U3491 (N_3491,N_2698,N_2510);
nor U3492 (N_3492,N_2538,N_2680);
xor U3493 (N_3493,N_2663,N_2730);
nor U3494 (N_3494,N_2858,N_2655);
xor U3495 (N_3495,N_2939,N_2512);
nor U3496 (N_3496,N_2670,N_2561);
and U3497 (N_3497,N_2946,N_2805);
or U3498 (N_3498,N_2874,N_2536);
or U3499 (N_3499,N_2553,N_2761);
xor U3500 (N_3500,N_3444,N_3240);
xnor U3501 (N_3501,N_3489,N_3291);
and U3502 (N_3502,N_3411,N_3137);
and U3503 (N_3503,N_3148,N_3025);
or U3504 (N_3504,N_3062,N_3490);
and U3505 (N_3505,N_3275,N_3453);
or U3506 (N_3506,N_3386,N_3316);
nor U3507 (N_3507,N_3263,N_3242);
nor U3508 (N_3508,N_3072,N_3269);
xnor U3509 (N_3509,N_3175,N_3041);
nor U3510 (N_3510,N_3116,N_3117);
nor U3511 (N_3511,N_3216,N_3380);
nor U3512 (N_3512,N_3225,N_3480);
xor U3513 (N_3513,N_3479,N_3324);
nand U3514 (N_3514,N_3382,N_3421);
nor U3515 (N_3515,N_3146,N_3425);
or U3516 (N_3516,N_3337,N_3310);
nand U3517 (N_3517,N_3153,N_3052);
and U3518 (N_3518,N_3270,N_3300);
xor U3519 (N_3519,N_3473,N_3363);
nor U3520 (N_3520,N_3404,N_3155);
or U3521 (N_3521,N_3235,N_3027);
nand U3522 (N_3522,N_3390,N_3230);
and U3523 (N_3523,N_3481,N_3384);
xor U3524 (N_3524,N_3004,N_3198);
and U3525 (N_3525,N_3405,N_3152);
xor U3526 (N_3526,N_3200,N_3005);
nand U3527 (N_3527,N_3008,N_3399);
or U3528 (N_3528,N_3340,N_3351);
and U3529 (N_3529,N_3167,N_3371);
or U3530 (N_3530,N_3123,N_3112);
or U3531 (N_3531,N_3187,N_3082);
and U3532 (N_3532,N_3066,N_3206);
nor U3533 (N_3533,N_3199,N_3410);
nand U3534 (N_3534,N_3438,N_3189);
nand U3535 (N_3535,N_3303,N_3249);
nand U3536 (N_3536,N_3472,N_3477);
xnor U3537 (N_3537,N_3201,N_3318);
or U3538 (N_3538,N_3369,N_3276);
nor U3539 (N_3539,N_3036,N_3252);
and U3540 (N_3540,N_3427,N_3184);
xnor U3541 (N_3541,N_3344,N_3026);
and U3542 (N_3542,N_3075,N_3045);
or U3543 (N_3543,N_3032,N_3266);
nor U3544 (N_3544,N_3284,N_3120);
xor U3545 (N_3545,N_3057,N_3499);
xnor U3546 (N_3546,N_3233,N_3278);
or U3547 (N_3547,N_3035,N_3089);
nor U3548 (N_3548,N_3437,N_3214);
nor U3549 (N_3549,N_3277,N_3389);
or U3550 (N_3550,N_3166,N_3090);
or U3551 (N_3551,N_3494,N_3271);
nand U3552 (N_3552,N_3431,N_3194);
or U3553 (N_3553,N_3244,N_3209);
and U3554 (N_3554,N_3498,N_3013);
xnor U3555 (N_3555,N_3264,N_3442);
or U3556 (N_3556,N_3463,N_3295);
xnor U3557 (N_3557,N_3367,N_3335);
nand U3558 (N_3558,N_3033,N_3238);
nand U3559 (N_3559,N_3468,N_3406);
xor U3560 (N_3560,N_3417,N_3109);
nand U3561 (N_3561,N_3193,N_3448);
or U3562 (N_3562,N_3403,N_3077);
xor U3563 (N_3563,N_3345,N_3034);
xnor U3564 (N_3564,N_3359,N_3086);
nor U3565 (N_3565,N_3044,N_3160);
nand U3566 (N_3566,N_3038,N_3069);
nor U3567 (N_3567,N_3451,N_3322);
xnor U3568 (N_3568,N_3311,N_3113);
or U3569 (N_3569,N_3255,N_3177);
nor U3570 (N_3570,N_3248,N_3128);
nor U3571 (N_3571,N_3450,N_3495);
nor U3572 (N_3572,N_3228,N_3434);
nand U3573 (N_3573,N_3063,N_3105);
nor U3574 (N_3574,N_3222,N_3354);
nand U3575 (N_3575,N_3119,N_3039);
or U3576 (N_3576,N_3169,N_3445);
xnor U3577 (N_3577,N_3124,N_3423);
xnor U3578 (N_3578,N_3383,N_3205);
nand U3579 (N_3579,N_3118,N_3400);
xnor U3580 (N_3580,N_3338,N_3103);
xnor U3581 (N_3581,N_3285,N_3084);
and U3582 (N_3582,N_3211,N_3164);
and U3583 (N_3583,N_3002,N_3458);
nor U3584 (N_3584,N_3001,N_3165);
xnor U3585 (N_3585,N_3296,N_3061);
nand U3586 (N_3586,N_3098,N_3293);
xnor U3587 (N_3587,N_3433,N_3179);
nor U3588 (N_3588,N_3254,N_3262);
nand U3589 (N_3589,N_3079,N_3343);
xor U3590 (N_3590,N_3016,N_3297);
or U3591 (N_3591,N_3029,N_3265);
and U3592 (N_3592,N_3286,N_3290);
nand U3593 (N_3593,N_3304,N_3009);
and U3594 (N_3594,N_3243,N_3455);
nand U3595 (N_3595,N_3274,N_3456);
nor U3596 (N_3596,N_3136,N_3110);
or U3597 (N_3597,N_3462,N_3190);
or U3598 (N_3598,N_3356,N_3172);
or U3599 (N_3599,N_3100,N_3215);
xor U3600 (N_3600,N_3102,N_3101);
or U3601 (N_3601,N_3111,N_3047);
and U3602 (N_3602,N_3070,N_3131);
nand U3603 (N_3603,N_3010,N_3186);
and U3604 (N_3604,N_3454,N_3094);
xnor U3605 (N_3605,N_3336,N_3125);
nor U3606 (N_3606,N_3093,N_3373);
and U3607 (N_3607,N_3151,N_3129);
nor U3608 (N_3608,N_3048,N_3461);
nand U3609 (N_3609,N_3145,N_3159);
nand U3610 (N_3610,N_3268,N_3099);
nor U3611 (N_3611,N_3173,N_3191);
nor U3612 (N_3612,N_3245,N_3358);
and U3613 (N_3613,N_3327,N_3301);
or U3614 (N_3614,N_3246,N_3402);
xnor U3615 (N_3615,N_3334,N_3071);
and U3616 (N_3616,N_3452,N_3279);
nand U3617 (N_3617,N_3024,N_3178);
or U3618 (N_3618,N_3317,N_3256);
nand U3619 (N_3619,N_3483,N_3493);
or U3620 (N_3620,N_3127,N_3474);
or U3621 (N_3621,N_3368,N_3023);
nor U3622 (N_3622,N_3292,N_3212);
nand U3623 (N_3623,N_3015,N_3306);
xnor U3624 (N_3624,N_3106,N_3046);
nand U3625 (N_3625,N_3372,N_3007);
and U3626 (N_3626,N_3022,N_3207);
nor U3627 (N_3627,N_3260,N_3298);
xnor U3628 (N_3628,N_3312,N_3294);
xor U3629 (N_3629,N_3006,N_3067);
nand U3630 (N_3630,N_3060,N_3439);
xnor U3631 (N_3631,N_3122,N_3229);
or U3632 (N_3632,N_3171,N_3435);
nor U3633 (N_3633,N_3357,N_3219);
nand U3634 (N_3634,N_3349,N_3174);
and U3635 (N_3635,N_3043,N_3388);
nor U3636 (N_3636,N_3287,N_3302);
or U3637 (N_3637,N_3227,N_3050);
xnor U3638 (N_3638,N_3202,N_3289);
and U3639 (N_3639,N_3428,N_3104);
xnor U3640 (N_3640,N_3154,N_3339);
xor U3641 (N_3641,N_3429,N_3486);
nor U3642 (N_3642,N_3261,N_3475);
xor U3643 (N_3643,N_3144,N_3091);
nand U3644 (N_3644,N_3299,N_3347);
nor U3645 (N_3645,N_3393,N_3096);
or U3646 (N_3646,N_3247,N_3234);
nor U3647 (N_3647,N_3196,N_3250);
nor U3648 (N_3648,N_3326,N_3440);
nor U3649 (N_3649,N_3012,N_3447);
and U3650 (N_3650,N_3134,N_3204);
and U3651 (N_3651,N_3115,N_3321);
nand U3652 (N_3652,N_3040,N_3288);
nor U3653 (N_3653,N_3073,N_3385);
xnor U3654 (N_3654,N_3253,N_3408);
or U3655 (N_3655,N_3487,N_3330);
and U3656 (N_3656,N_3161,N_3471);
nand U3657 (N_3657,N_3095,N_3181);
nor U3658 (N_3658,N_3000,N_3464);
or U3659 (N_3659,N_3350,N_3436);
or U3660 (N_3660,N_3381,N_3315);
nor U3661 (N_3661,N_3221,N_3192);
nor U3662 (N_3662,N_3108,N_3366);
nand U3663 (N_3663,N_3396,N_3195);
and U3664 (N_3664,N_3011,N_3259);
nor U3665 (N_3665,N_3018,N_3126);
xor U3666 (N_3666,N_3051,N_3037);
xor U3667 (N_3667,N_3021,N_3348);
nor U3668 (N_3668,N_3378,N_3485);
nand U3669 (N_3669,N_3355,N_3017);
nor U3670 (N_3670,N_3319,N_3149);
or U3671 (N_3671,N_3163,N_3398);
xor U3672 (N_3672,N_3394,N_3346);
nand U3673 (N_3673,N_3183,N_3375);
xor U3674 (N_3674,N_3076,N_3496);
nand U3675 (N_3675,N_3132,N_3059);
xor U3676 (N_3676,N_3432,N_3443);
and U3677 (N_3677,N_3391,N_3465);
or U3678 (N_3678,N_3370,N_3459);
or U3679 (N_3679,N_3413,N_3203);
xnor U3680 (N_3680,N_3401,N_3135);
and U3681 (N_3681,N_3491,N_3208);
nor U3682 (N_3682,N_3220,N_3068);
and U3683 (N_3683,N_3308,N_3283);
nor U3684 (N_3684,N_3441,N_3418);
nor U3685 (N_3685,N_3087,N_3130);
nor U3686 (N_3686,N_3049,N_3446);
nand U3687 (N_3687,N_3139,N_3085);
and U3688 (N_3688,N_3042,N_3114);
nand U3689 (N_3689,N_3313,N_3064);
nand U3690 (N_3690,N_3223,N_3392);
nor U3691 (N_3691,N_3231,N_3232);
nor U3692 (N_3692,N_3088,N_3158);
xnor U3693 (N_3693,N_3210,N_3014);
xor U3694 (N_3694,N_3218,N_3150);
nor U3695 (N_3695,N_3281,N_3328);
and U3696 (N_3696,N_3476,N_3314);
nand U3697 (N_3697,N_3156,N_3267);
nor U3698 (N_3698,N_3019,N_3185);
nor U3699 (N_3699,N_3412,N_3056);
nor U3700 (N_3700,N_3168,N_3020);
nor U3701 (N_3701,N_3377,N_3031);
or U3702 (N_3702,N_3416,N_3467);
nor U3703 (N_3703,N_3466,N_3449);
nand U3704 (N_3704,N_3469,N_3419);
nand U3705 (N_3705,N_3141,N_3307);
nor U3706 (N_3706,N_3217,N_3420);
nor U3707 (N_3707,N_3182,N_3080);
or U3708 (N_3708,N_3083,N_3365);
nor U3709 (N_3709,N_3147,N_3360);
nor U3710 (N_3710,N_3379,N_3376);
nor U3711 (N_3711,N_3305,N_3342);
and U3712 (N_3712,N_3197,N_3488);
nor U3713 (N_3713,N_3341,N_3460);
nor U3714 (N_3714,N_3484,N_3457);
and U3715 (N_3715,N_3092,N_3236);
or U3716 (N_3716,N_3188,N_3239);
nand U3717 (N_3717,N_3309,N_3078);
or U3718 (N_3718,N_3251,N_3180);
nand U3719 (N_3719,N_3140,N_3362);
nor U3720 (N_3720,N_3387,N_3329);
nand U3721 (N_3721,N_3224,N_3422);
nor U3722 (N_3722,N_3353,N_3097);
xor U3723 (N_3723,N_3055,N_3054);
xor U3724 (N_3724,N_3352,N_3374);
nor U3725 (N_3725,N_3320,N_3325);
xor U3726 (N_3726,N_3323,N_3282);
nor U3727 (N_3727,N_3395,N_3053);
nand U3728 (N_3728,N_3492,N_3482);
or U3729 (N_3729,N_3058,N_3121);
nand U3730 (N_3730,N_3258,N_3397);
nand U3731 (N_3731,N_3143,N_3333);
xnor U3732 (N_3732,N_3407,N_3241);
xnor U3733 (N_3733,N_3237,N_3081);
nand U3734 (N_3734,N_3273,N_3138);
xnor U3735 (N_3735,N_3107,N_3272);
nor U3736 (N_3736,N_3170,N_3157);
or U3737 (N_3737,N_3332,N_3331);
or U3738 (N_3738,N_3426,N_3176);
or U3739 (N_3739,N_3030,N_3213);
or U3740 (N_3740,N_3257,N_3424);
nand U3741 (N_3741,N_3409,N_3470);
xnor U3742 (N_3742,N_3361,N_3028);
nand U3743 (N_3743,N_3074,N_3414);
or U3744 (N_3744,N_3478,N_3415);
or U3745 (N_3745,N_3133,N_3226);
nand U3746 (N_3746,N_3162,N_3003);
nor U3747 (N_3747,N_3142,N_3364);
nor U3748 (N_3748,N_3065,N_3280);
nand U3749 (N_3749,N_3497,N_3430);
and U3750 (N_3750,N_3485,N_3156);
and U3751 (N_3751,N_3192,N_3468);
nor U3752 (N_3752,N_3285,N_3251);
and U3753 (N_3753,N_3338,N_3405);
or U3754 (N_3754,N_3253,N_3053);
or U3755 (N_3755,N_3101,N_3364);
nor U3756 (N_3756,N_3487,N_3052);
or U3757 (N_3757,N_3157,N_3055);
xor U3758 (N_3758,N_3235,N_3360);
or U3759 (N_3759,N_3474,N_3498);
nor U3760 (N_3760,N_3440,N_3287);
and U3761 (N_3761,N_3445,N_3408);
and U3762 (N_3762,N_3201,N_3438);
and U3763 (N_3763,N_3042,N_3022);
or U3764 (N_3764,N_3031,N_3326);
nand U3765 (N_3765,N_3497,N_3288);
xor U3766 (N_3766,N_3038,N_3031);
xnor U3767 (N_3767,N_3081,N_3341);
nor U3768 (N_3768,N_3370,N_3030);
or U3769 (N_3769,N_3433,N_3043);
or U3770 (N_3770,N_3243,N_3184);
or U3771 (N_3771,N_3356,N_3295);
nor U3772 (N_3772,N_3097,N_3219);
or U3773 (N_3773,N_3222,N_3253);
nand U3774 (N_3774,N_3296,N_3027);
and U3775 (N_3775,N_3455,N_3459);
nand U3776 (N_3776,N_3470,N_3052);
nor U3777 (N_3777,N_3143,N_3162);
or U3778 (N_3778,N_3022,N_3487);
nor U3779 (N_3779,N_3429,N_3409);
or U3780 (N_3780,N_3110,N_3215);
nor U3781 (N_3781,N_3275,N_3140);
xor U3782 (N_3782,N_3304,N_3174);
nor U3783 (N_3783,N_3200,N_3206);
or U3784 (N_3784,N_3429,N_3216);
nor U3785 (N_3785,N_3021,N_3380);
nand U3786 (N_3786,N_3119,N_3496);
or U3787 (N_3787,N_3434,N_3045);
xor U3788 (N_3788,N_3362,N_3366);
xor U3789 (N_3789,N_3047,N_3156);
nand U3790 (N_3790,N_3000,N_3289);
nand U3791 (N_3791,N_3018,N_3080);
and U3792 (N_3792,N_3419,N_3162);
and U3793 (N_3793,N_3487,N_3114);
and U3794 (N_3794,N_3162,N_3133);
xnor U3795 (N_3795,N_3156,N_3163);
nand U3796 (N_3796,N_3405,N_3279);
nor U3797 (N_3797,N_3476,N_3284);
and U3798 (N_3798,N_3288,N_3445);
xor U3799 (N_3799,N_3340,N_3475);
xor U3800 (N_3800,N_3492,N_3322);
xor U3801 (N_3801,N_3437,N_3132);
nand U3802 (N_3802,N_3185,N_3124);
nand U3803 (N_3803,N_3347,N_3459);
or U3804 (N_3804,N_3271,N_3008);
xor U3805 (N_3805,N_3213,N_3419);
or U3806 (N_3806,N_3450,N_3339);
nand U3807 (N_3807,N_3220,N_3294);
or U3808 (N_3808,N_3017,N_3323);
and U3809 (N_3809,N_3236,N_3251);
nor U3810 (N_3810,N_3325,N_3095);
and U3811 (N_3811,N_3225,N_3344);
and U3812 (N_3812,N_3058,N_3364);
nand U3813 (N_3813,N_3030,N_3204);
or U3814 (N_3814,N_3037,N_3038);
nand U3815 (N_3815,N_3149,N_3265);
xor U3816 (N_3816,N_3348,N_3095);
xnor U3817 (N_3817,N_3356,N_3062);
nor U3818 (N_3818,N_3025,N_3105);
nand U3819 (N_3819,N_3015,N_3227);
nor U3820 (N_3820,N_3230,N_3232);
nor U3821 (N_3821,N_3194,N_3273);
and U3822 (N_3822,N_3157,N_3295);
or U3823 (N_3823,N_3439,N_3036);
nand U3824 (N_3824,N_3082,N_3437);
and U3825 (N_3825,N_3026,N_3324);
or U3826 (N_3826,N_3294,N_3378);
or U3827 (N_3827,N_3122,N_3293);
nor U3828 (N_3828,N_3119,N_3499);
or U3829 (N_3829,N_3080,N_3369);
xor U3830 (N_3830,N_3399,N_3031);
xor U3831 (N_3831,N_3101,N_3308);
nand U3832 (N_3832,N_3390,N_3494);
nand U3833 (N_3833,N_3474,N_3178);
nand U3834 (N_3834,N_3240,N_3293);
xnor U3835 (N_3835,N_3244,N_3323);
or U3836 (N_3836,N_3423,N_3182);
and U3837 (N_3837,N_3492,N_3196);
or U3838 (N_3838,N_3188,N_3459);
xor U3839 (N_3839,N_3236,N_3482);
nand U3840 (N_3840,N_3011,N_3073);
and U3841 (N_3841,N_3251,N_3357);
nand U3842 (N_3842,N_3054,N_3003);
nor U3843 (N_3843,N_3247,N_3453);
nand U3844 (N_3844,N_3356,N_3202);
and U3845 (N_3845,N_3467,N_3492);
xor U3846 (N_3846,N_3268,N_3303);
and U3847 (N_3847,N_3079,N_3325);
nand U3848 (N_3848,N_3373,N_3276);
and U3849 (N_3849,N_3225,N_3309);
nand U3850 (N_3850,N_3404,N_3000);
xnor U3851 (N_3851,N_3189,N_3442);
xnor U3852 (N_3852,N_3021,N_3430);
nor U3853 (N_3853,N_3017,N_3467);
or U3854 (N_3854,N_3062,N_3233);
nand U3855 (N_3855,N_3327,N_3159);
nor U3856 (N_3856,N_3131,N_3197);
or U3857 (N_3857,N_3111,N_3430);
nor U3858 (N_3858,N_3382,N_3462);
or U3859 (N_3859,N_3084,N_3265);
xor U3860 (N_3860,N_3108,N_3394);
or U3861 (N_3861,N_3274,N_3206);
and U3862 (N_3862,N_3135,N_3076);
xor U3863 (N_3863,N_3121,N_3188);
xor U3864 (N_3864,N_3304,N_3267);
nor U3865 (N_3865,N_3029,N_3156);
nand U3866 (N_3866,N_3152,N_3111);
or U3867 (N_3867,N_3081,N_3152);
nand U3868 (N_3868,N_3484,N_3306);
or U3869 (N_3869,N_3012,N_3454);
or U3870 (N_3870,N_3241,N_3005);
nor U3871 (N_3871,N_3160,N_3446);
xnor U3872 (N_3872,N_3006,N_3001);
and U3873 (N_3873,N_3146,N_3245);
xnor U3874 (N_3874,N_3251,N_3264);
nor U3875 (N_3875,N_3460,N_3024);
nand U3876 (N_3876,N_3305,N_3439);
xor U3877 (N_3877,N_3221,N_3185);
xnor U3878 (N_3878,N_3367,N_3179);
xnor U3879 (N_3879,N_3038,N_3398);
or U3880 (N_3880,N_3224,N_3200);
or U3881 (N_3881,N_3472,N_3393);
nor U3882 (N_3882,N_3073,N_3090);
nor U3883 (N_3883,N_3030,N_3120);
or U3884 (N_3884,N_3453,N_3480);
or U3885 (N_3885,N_3436,N_3262);
xnor U3886 (N_3886,N_3492,N_3224);
or U3887 (N_3887,N_3303,N_3071);
xor U3888 (N_3888,N_3367,N_3302);
and U3889 (N_3889,N_3171,N_3080);
xor U3890 (N_3890,N_3368,N_3277);
xor U3891 (N_3891,N_3243,N_3208);
nor U3892 (N_3892,N_3197,N_3492);
xor U3893 (N_3893,N_3080,N_3424);
or U3894 (N_3894,N_3068,N_3354);
nor U3895 (N_3895,N_3302,N_3498);
nand U3896 (N_3896,N_3214,N_3183);
and U3897 (N_3897,N_3181,N_3051);
nor U3898 (N_3898,N_3296,N_3059);
and U3899 (N_3899,N_3194,N_3345);
or U3900 (N_3900,N_3092,N_3078);
and U3901 (N_3901,N_3198,N_3034);
nor U3902 (N_3902,N_3298,N_3405);
nand U3903 (N_3903,N_3306,N_3039);
or U3904 (N_3904,N_3276,N_3347);
xnor U3905 (N_3905,N_3071,N_3494);
nand U3906 (N_3906,N_3392,N_3335);
nand U3907 (N_3907,N_3072,N_3147);
nand U3908 (N_3908,N_3081,N_3499);
or U3909 (N_3909,N_3189,N_3045);
and U3910 (N_3910,N_3153,N_3232);
nand U3911 (N_3911,N_3433,N_3155);
or U3912 (N_3912,N_3148,N_3233);
and U3913 (N_3913,N_3100,N_3341);
or U3914 (N_3914,N_3382,N_3201);
nor U3915 (N_3915,N_3341,N_3361);
nor U3916 (N_3916,N_3014,N_3450);
xor U3917 (N_3917,N_3310,N_3322);
xor U3918 (N_3918,N_3148,N_3264);
and U3919 (N_3919,N_3189,N_3089);
nand U3920 (N_3920,N_3468,N_3024);
or U3921 (N_3921,N_3440,N_3161);
nor U3922 (N_3922,N_3399,N_3113);
and U3923 (N_3923,N_3233,N_3472);
xor U3924 (N_3924,N_3371,N_3204);
or U3925 (N_3925,N_3469,N_3324);
or U3926 (N_3926,N_3319,N_3401);
nor U3927 (N_3927,N_3243,N_3446);
or U3928 (N_3928,N_3178,N_3207);
nor U3929 (N_3929,N_3095,N_3480);
and U3930 (N_3930,N_3426,N_3076);
xor U3931 (N_3931,N_3486,N_3474);
and U3932 (N_3932,N_3023,N_3199);
xor U3933 (N_3933,N_3390,N_3409);
and U3934 (N_3934,N_3230,N_3421);
nor U3935 (N_3935,N_3312,N_3307);
nand U3936 (N_3936,N_3007,N_3498);
and U3937 (N_3937,N_3282,N_3265);
and U3938 (N_3938,N_3287,N_3493);
and U3939 (N_3939,N_3256,N_3259);
xor U3940 (N_3940,N_3400,N_3344);
or U3941 (N_3941,N_3285,N_3164);
nand U3942 (N_3942,N_3186,N_3130);
xnor U3943 (N_3943,N_3468,N_3288);
xor U3944 (N_3944,N_3257,N_3421);
and U3945 (N_3945,N_3185,N_3345);
nand U3946 (N_3946,N_3256,N_3445);
nand U3947 (N_3947,N_3448,N_3442);
or U3948 (N_3948,N_3103,N_3173);
or U3949 (N_3949,N_3126,N_3113);
nor U3950 (N_3950,N_3188,N_3483);
and U3951 (N_3951,N_3206,N_3273);
nand U3952 (N_3952,N_3373,N_3286);
nor U3953 (N_3953,N_3065,N_3357);
or U3954 (N_3954,N_3476,N_3455);
nor U3955 (N_3955,N_3080,N_3073);
or U3956 (N_3956,N_3115,N_3237);
xor U3957 (N_3957,N_3479,N_3199);
and U3958 (N_3958,N_3273,N_3344);
and U3959 (N_3959,N_3471,N_3076);
nand U3960 (N_3960,N_3104,N_3299);
and U3961 (N_3961,N_3323,N_3054);
nor U3962 (N_3962,N_3434,N_3235);
nor U3963 (N_3963,N_3028,N_3457);
nor U3964 (N_3964,N_3279,N_3393);
nand U3965 (N_3965,N_3496,N_3137);
and U3966 (N_3966,N_3285,N_3119);
nand U3967 (N_3967,N_3419,N_3452);
and U3968 (N_3968,N_3471,N_3483);
nor U3969 (N_3969,N_3392,N_3372);
xor U3970 (N_3970,N_3099,N_3236);
or U3971 (N_3971,N_3258,N_3029);
xor U3972 (N_3972,N_3015,N_3221);
nor U3973 (N_3973,N_3359,N_3286);
xnor U3974 (N_3974,N_3036,N_3484);
nor U3975 (N_3975,N_3367,N_3443);
or U3976 (N_3976,N_3419,N_3047);
nor U3977 (N_3977,N_3169,N_3209);
nor U3978 (N_3978,N_3186,N_3251);
xor U3979 (N_3979,N_3048,N_3167);
nand U3980 (N_3980,N_3294,N_3400);
and U3981 (N_3981,N_3012,N_3355);
or U3982 (N_3982,N_3180,N_3438);
nor U3983 (N_3983,N_3021,N_3400);
and U3984 (N_3984,N_3285,N_3121);
or U3985 (N_3985,N_3315,N_3053);
nor U3986 (N_3986,N_3124,N_3374);
and U3987 (N_3987,N_3035,N_3124);
xor U3988 (N_3988,N_3033,N_3282);
xor U3989 (N_3989,N_3144,N_3350);
xnor U3990 (N_3990,N_3387,N_3070);
and U3991 (N_3991,N_3044,N_3247);
nor U3992 (N_3992,N_3408,N_3050);
and U3993 (N_3993,N_3383,N_3349);
or U3994 (N_3994,N_3316,N_3097);
xnor U3995 (N_3995,N_3033,N_3060);
xor U3996 (N_3996,N_3045,N_3123);
nand U3997 (N_3997,N_3366,N_3197);
and U3998 (N_3998,N_3167,N_3201);
xnor U3999 (N_3999,N_3159,N_3101);
or U4000 (N_4000,N_3874,N_3640);
nor U4001 (N_4001,N_3747,N_3942);
nand U4002 (N_4002,N_3614,N_3579);
nor U4003 (N_4003,N_3604,N_3516);
xnor U4004 (N_4004,N_3897,N_3683);
and U4005 (N_4005,N_3616,N_3500);
nand U4006 (N_4006,N_3847,N_3755);
and U4007 (N_4007,N_3827,N_3704);
and U4008 (N_4008,N_3896,N_3633);
nand U4009 (N_4009,N_3799,N_3679);
and U4010 (N_4010,N_3694,N_3963);
or U4011 (N_4011,N_3918,N_3900);
and U4012 (N_4012,N_3526,N_3651);
nand U4013 (N_4013,N_3591,N_3710);
nor U4014 (N_4014,N_3842,N_3766);
xor U4015 (N_4015,N_3939,N_3811);
nor U4016 (N_4016,N_3760,N_3693);
nor U4017 (N_4017,N_3719,N_3666);
nand U4018 (N_4018,N_3731,N_3586);
xor U4019 (N_4019,N_3739,N_3785);
and U4020 (N_4020,N_3905,N_3836);
and U4021 (N_4021,N_3853,N_3922);
xnor U4022 (N_4022,N_3517,N_3549);
and U4023 (N_4023,N_3955,N_3953);
and U4024 (N_4024,N_3854,N_3912);
or U4025 (N_4025,N_3891,N_3584);
nor U4026 (N_4026,N_3966,N_3792);
nand U4027 (N_4027,N_3934,N_3818);
nand U4028 (N_4028,N_3665,N_3743);
and U4029 (N_4029,N_3813,N_3736);
xnor U4030 (N_4030,N_3916,N_3812);
nand U4031 (N_4031,N_3833,N_3636);
xor U4032 (N_4032,N_3835,N_3932);
nand U4033 (N_4033,N_3995,N_3774);
nand U4034 (N_4034,N_3856,N_3938);
xnor U4035 (N_4035,N_3940,N_3978);
nand U4036 (N_4036,N_3879,N_3554);
nand U4037 (N_4037,N_3696,N_3546);
and U4038 (N_4038,N_3864,N_3589);
and U4039 (N_4039,N_3937,N_3750);
nand U4040 (N_4040,N_3634,N_3730);
nor U4041 (N_4041,N_3506,N_3684);
nand U4042 (N_4042,N_3569,N_3822);
nand U4043 (N_4043,N_3594,N_3674);
nand U4044 (N_4044,N_3769,N_3678);
and U4045 (N_4045,N_3565,N_3954);
nand U4046 (N_4046,N_3968,N_3789);
and U4047 (N_4047,N_3949,N_3510);
or U4048 (N_4048,N_3598,N_3733);
nor U4049 (N_4049,N_3685,N_3712);
nor U4050 (N_4050,N_3592,N_3946);
or U4051 (N_4051,N_3858,N_3837);
xnor U4052 (N_4052,N_3692,N_3987);
nor U4053 (N_4053,N_3819,N_3863);
nor U4054 (N_4054,N_3568,N_3791);
xnor U4055 (N_4055,N_3534,N_3843);
or U4056 (N_4056,N_3642,N_3512);
and U4057 (N_4057,N_3830,N_3699);
xor U4058 (N_4058,N_3825,N_3556);
nor U4059 (N_4059,N_3862,N_3804);
and U4060 (N_4060,N_3979,N_3670);
and U4061 (N_4061,N_3610,N_3869);
nand U4062 (N_4062,N_3522,N_3521);
and U4063 (N_4063,N_3971,N_3680);
xnor U4064 (N_4064,N_3548,N_3664);
or U4065 (N_4065,N_3880,N_3926);
nand U4066 (N_4066,N_3723,N_3682);
and U4067 (N_4067,N_3524,N_3761);
nand U4068 (N_4068,N_3889,N_3502);
and U4069 (N_4069,N_3732,N_3801);
xor U4070 (N_4070,N_3657,N_3991);
and U4071 (N_4071,N_3803,N_3841);
or U4072 (N_4072,N_3722,N_3566);
and U4073 (N_4073,N_3536,N_3740);
and U4074 (N_4074,N_3532,N_3550);
nor U4075 (N_4075,N_3805,N_3538);
xor U4076 (N_4076,N_3845,N_3824);
nand U4077 (N_4077,N_3686,N_3910);
nand U4078 (N_4078,N_3840,N_3793);
nor U4079 (N_4079,N_3823,N_3697);
and U4080 (N_4080,N_3795,N_3871);
or U4081 (N_4081,N_3742,N_3802);
or U4082 (N_4082,N_3588,N_3878);
and U4083 (N_4083,N_3915,N_3571);
or U4084 (N_4084,N_3936,N_3706);
or U4085 (N_4085,N_3558,N_3515);
nor U4086 (N_4086,N_3903,N_3709);
nor U4087 (N_4087,N_3893,N_3529);
xnor U4088 (N_4088,N_3638,N_3757);
nor U4089 (N_4089,N_3875,N_3773);
nand U4090 (N_4090,N_3668,N_3528);
and U4091 (N_4091,N_3615,N_3831);
nand U4092 (N_4092,N_3846,N_3844);
and U4093 (N_4093,N_3715,N_3655);
and U4094 (N_4094,N_3980,N_3751);
xnor U4095 (N_4095,N_3876,N_3624);
xnor U4096 (N_4096,N_3577,N_3720);
or U4097 (N_4097,N_3572,N_3783);
or U4098 (N_4098,N_3794,N_3718);
nand U4099 (N_4099,N_3930,N_3676);
xnor U4100 (N_4100,N_3659,N_3698);
and U4101 (N_4101,N_3859,N_3919);
and U4102 (N_4102,N_3713,N_3611);
xnor U4103 (N_4103,N_3628,N_3920);
nand U4104 (N_4104,N_3944,N_3618);
or U4105 (N_4105,N_3931,N_3660);
or U4106 (N_4106,N_3906,N_3927);
nand U4107 (N_4107,N_3653,N_3737);
nand U4108 (N_4108,N_3977,N_3644);
xor U4109 (N_4109,N_3511,N_3990);
or U4110 (N_4110,N_3902,N_3575);
nand U4111 (N_4111,N_3834,N_3892);
and U4112 (N_4112,N_3951,N_3559);
nor U4113 (N_4113,N_3625,N_3908);
nor U4114 (N_4114,N_3508,N_3829);
nand U4115 (N_4115,N_3907,N_3580);
nand U4116 (N_4116,N_3525,N_3754);
nor U4117 (N_4117,N_3778,N_3999);
nor U4118 (N_4118,N_3551,N_3917);
nand U4119 (N_4119,N_3620,N_3563);
nand U4120 (N_4120,N_3816,N_3702);
nor U4121 (N_4121,N_3690,N_3958);
nor U4122 (N_4122,N_3535,N_3721);
xnor U4123 (N_4123,N_3839,N_3590);
or U4124 (N_4124,N_3701,N_3643);
or U4125 (N_4125,N_3639,N_3882);
nand U4126 (N_4126,N_3852,N_3790);
nor U4127 (N_4127,N_3972,N_3581);
or U4128 (N_4128,N_3585,N_3714);
nor U4129 (N_4129,N_3541,N_3545);
xnor U4130 (N_4130,N_3716,N_3641);
xnor U4131 (N_4131,N_3923,N_3602);
nor U4132 (N_4132,N_3850,N_3899);
nand U4133 (N_4133,N_3725,N_3543);
or U4134 (N_4134,N_3505,N_3531);
nor U4135 (N_4135,N_3888,N_3994);
and U4136 (N_4136,N_3860,N_3851);
nor U4137 (N_4137,N_3998,N_3989);
or U4138 (N_4138,N_3738,N_3996);
xor U4139 (N_4139,N_3870,N_3983);
nor U4140 (N_4140,N_3909,N_3654);
and U4141 (N_4141,N_3509,N_3895);
nand U4142 (N_4142,N_3914,N_3782);
nand U4143 (N_4143,N_3962,N_3630);
or U4144 (N_4144,N_3970,N_3735);
nand U4145 (N_4145,N_3700,N_3943);
nor U4146 (N_4146,N_3941,N_3560);
and U4147 (N_4147,N_3788,N_3992);
or U4148 (N_4148,N_3729,N_3796);
nor U4149 (N_4149,N_3768,N_3599);
or U4150 (N_4150,N_3724,N_3973);
nor U4151 (N_4151,N_3646,N_3520);
and U4152 (N_4152,N_3772,N_3519);
and U4153 (N_4153,N_3688,N_3775);
and U4154 (N_4154,N_3652,N_3985);
and U4155 (N_4155,N_3911,N_3540);
xor U4156 (N_4156,N_3925,N_3626);
nand U4157 (N_4157,N_3607,N_3935);
nand U4158 (N_4158,N_3514,N_3527);
nor U4159 (N_4159,N_3809,N_3798);
and U4160 (N_4160,N_3663,N_3650);
and U4161 (N_4161,N_3595,N_3838);
and U4162 (N_4162,N_3726,N_3956);
nor U4163 (N_4163,N_3649,N_3617);
and U4164 (N_4164,N_3993,N_3627);
and U4165 (N_4165,N_3632,N_3763);
xnor U4166 (N_4166,N_3921,N_3501);
xnor U4167 (N_4167,N_3518,N_3848);
nor U4168 (N_4168,N_3821,N_3557);
nand U4169 (N_4169,N_3564,N_3744);
or U4170 (N_4170,N_3997,N_3904);
and U4171 (N_4171,N_3597,N_3562);
and U4172 (N_4172,N_3658,N_3779);
nand U4173 (N_4173,N_3807,N_3894);
nand U4174 (N_4174,N_3887,N_3984);
nand U4175 (N_4175,N_3947,N_3814);
and U4176 (N_4176,N_3857,N_3877);
nand U4177 (N_4177,N_3787,N_3734);
nor U4178 (N_4178,N_3695,N_3758);
or U4179 (N_4179,N_3924,N_3583);
or U4180 (N_4180,N_3800,N_3974);
and U4181 (N_4181,N_3537,N_3884);
nand U4182 (N_4182,N_3945,N_3960);
nand U4183 (N_4183,N_3952,N_3645);
or U4184 (N_4184,N_3544,N_3605);
and U4185 (N_4185,N_3703,N_3957);
or U4186 (N_4186,N_3752,N_3913);
or U4187 (N_4187,N_3865,N_3885);
and U4188 (N_4188,N_3507,N_3759);
and U4189 (N_4189,N_3777,N_3687);
nand U4190 (N_4190,N_3959,N_3832);
nand U4191 (N_4191,N_3728,N_3622);
and U4192 (N_4192,N_3547,N_3975);
xnor U4193 (N_4193,N_3948,N_3770);
and U4194 (N_4194,N_3672,N_3555);
nor U4195 (N_4195,N_3866,N_3629);
and U4196 (N_4196,N_3553,N_3867);
nand U4197 (N_4197,N_3705,N_3587);
or U4198 (N_4198,N_3606,N_3868);
xnor U4199 (N_4199,N_3808,N_3886);
or U4200 (N_4200,N_3741,N_3901);
nor U4201 (N_4201,N_3817,N_3609);
xnor U4202 (N_4202,N_3573,N_3539);
or U4203 (N_4203,N_3561,N_3708);
nor U4204 (N_4204,N_3745,N_3771);
and U4205 (N_4205,N_3756,N_3523);
and U4206 (N_4206,N_3542,N_3578);
xnor U4207 (N_4207,N_3574,N_3872);
xnor U4208 (N_4208,N_3890,N_3593);
and U4209 (N_4209,N_3675,N_3621);
and U4210 (N_4210,N_3691,N_3567);
or U4211 (N_4211,N_3810,N_3619);
and U4212 (N_4212,N_3603,N_3883);
xnor U4213 (N_4213,N_3797,N_3647);
nor U4214 (N_4214,N_3828,N_3671);
or U4215 (N_4215,N_3806,N_3503);
xnor U4216 (N_4216,N_3533,N_3929);
nand U4217 (N_4217,N_3784,N_3707);
nand U4218 (N_4218,N_3570,N_3513);
or U4219 (N_4219,N_3855,N_3964);
and U4220 (N_4220,N_3669,N_3982);
nand U4221 (N_4221,N_3965,N_3849);
nand U4222 (N_4222,N_3820,N_3746);
xor U4223 (N_4223,N_3976,N_3600);
or U4224 (N_4224,N_3612,N_3780);
or U4225 (N_4225,N_3764,N_3933);
xnor U4226 (N_4226,N_3631,N_3762);
nor U4227 (N_4227,N_3661,N_3988);
nand U4228 (N_4228,N_3689,N_3673);
nand U4229 (N_4229,N_3881,N_3748);
or U4230 (N_4230,N_3530,N_3861);
or U4231 (N_4231,N_3786,N_3648);
nand U4232 (N_4232,N_3753,N_3767);
and U4233 (N_4233,N_3717,N_3898);
and U4234 (N_4234,N_3981,N_3781);
nor U4235 (N_4235,N_3969,N_3635);
nand U4236 (N_4236,N_3576,N_3986);
and U4237 (N_4237,N_3656,N_3623);
and U4238 (N_4238,N_3826,N_3608);
nor U4239 (N_4239,N_3596,N_3727);
nor U4240 (N_4240,N_3928,N_3667);
nor U4241 (N_4241,N_3815,N_3601);
nor U4242 (N_4242,N_3582,N_3776);
and U4243 (N_4243,N_3662,N_3681);
xnor U4244 (N_4244,N_3873,N_3950);
xnor U4245 (N_4245,N_3765,N_3967);
and U4246 (N_4246,N_3749,N_3504);
xor U4247 (N_4247,N_3552,N_3637);
or U4248 (N_4248,N_3677,N_3711);
or U4249 (N_4249,N_3961,N_3613);
or U4250 (N_4250,N_3506,N_3551);
nand U4251 (N_4251,N_3735,N_3687);
nor U4252 (N_4252,N_3561,N_3601);
or U4253 (N_4253,N_3566,N_3527);
and U4254 (N_4254,N_3661,N_3767);
and U4255 (N_4255,N_3994,N_3581);
nand U4256 (N_4256,N_3554,N_3660);
and U4257 (N_4257,N_3555,N_3631);
or U4258 (N_4258,N_3540,N_3904);
or U4259 (N_4259,N_3610,N_3578);
nor U4260 (N_4260,N_3806,N_3979);
nor U4261 (N_4261,N_3705,N_3583);
and U4262 (N_4262,N_3568,N_3528);
xor U4263 (N_4263,N_3505,N_3665);
and U4264 (N_4264,N_3693,N_3956);
xor U4265 (N_4265,N_3596,N_3547);
nor U4266 (N_4266,N_3890,N_3585);
xnor U4267 (N_4267,N_3547,N_3796);
nand U4268 (N_4268,N_3860,N_3595);
and U4269 (N_4269,N_3936,N_3787);
or U4270 (N_4270,N_3789,N_3622);
nand U4271 (N_4271,N_3575,N_3761);
xnor U4272 (N_4272,N_3879,N_3713);
or U4273 (N_4273,N_3706,N_3647);
nor U4274 (N_4274,N_3982,N_3945);
xnor U4275 (N_4275,N_3533,N_3816);
nor U4276 (N_4276,N_3665,N_3681);
or U4277 (N_4277,N_3716,N_3619);
and U4278 (N_4278,N_3803,N_3668);
nand U4279 (N_4279,N_3826,N_3778);
and U4280 (N_4280,N_3803,N_3787);
nand U4281 (N_4281,N_3638,N_3601);
nor U4282 (N_4282,N_3909,N_3605);
xor U4283 (N_4283,N_3935,N_3556);
or U4284 (N_4284,N_3518,N_3954);
nor U4285 (N_4285,N_3507,N_3932);
and U4286 (N_4286,N_3746,N_3513);
or U4287 (N_4287,N_3704,N_3549);
nor U4288 (N_4288,N_3520,N_3669);
and U4289 (N_4289,N_3526,N_3548);
nor U4290 (N_4290,N_3651,N_3720);
nand U4291 (N_4291,N_3785,N_3775);
xor U4292 (N_4292,N_3706,N_3639);
or U4293 (N_4293,N_3588,N_3962);
nor U4294 (N_4294,N_3982,N_3793);
xnor U4295 (N_4295,N_3874,N_3782);
and U4296 (N_4296,N_3788,N_3916);
or U4297 (N_4297,N_3826,N_3632);
nand U4298 (N_4298,N_3523,N_3505);
xor U4299 (N_4299,N_3831,N_3588);
xnor U4300 (N_4300,N_3916,N_3732);
nand U4301 (N_4301,N_3923,N_3796);
nand U4302 (N_4302,N_3632,N_3891);
xnor U4303 (N_4303,N_3643,N_3812);
or U4304 (N_4304,N_3717,N_3991);
xor U4305 (N_4305,N_3656,N_3580);
and U4306 (N_4306,N_3834,N_3888);
nand U4307 (N_4307,N_3849,N_3596);
nand U4308 (N_4308,N_3926,N_3656);
nor U4309 (N_4309,N_3722,N_3535);
and U4310 (N_4310,N_3567,N_3528);
xnor U4311 (N_4311,N_3663,N_3774);
nand U4312 (N_4312,N_3869,N_3809);
xor U4313 (N_4313,N_3843,N_3825);
nand U4314 (N_4314,N_3887,N_3670);
or U4315 (N_4315,N_3943,N_3831);
nor U4316 (N_4316,N_3721,N_3545);
xor U4317 (N_4317,N_3910,N_3515);
or U4318 (N_4318,N_3704,N_3570);
nor U4319 (N_4319,N_3865,N_3965);
xor U4320 (N_4320,N_3652,N_3736);
xor U4321 (N_4321,N_3804,N_3632);
and U4322 (N_4322,N_3746,N_3575);
nor U4323 (N_4323,N_3958,N_3515);
xnor U4324 (N_4324,N_3598,N_3615);
or U4325 (N_4325,N_3910,N_3672);
nor U4326 (N_4326,N_3892,N_3546);
and U4327 (N_4327,N_3775,N_3984);
nand U4328 (N_4328,N_3649,N_3776);
nand U4329 (N_4329,N_3516,N_3550);
nand U4330 (N_4330,N_3878,N_3809);
or U4331 (N_4331,N_3976,N_3979);
xor U4332 (N_4332,N_3875,N_3604);
nor U4333 (N_4333,N_3836,N_3922);
nor U4334 (N_4334,N_3531,N_3524);
or U4335 (N_4335,N_3667,N_3688);
or U4336 (N_4336,N_3955,N_3599);
and U4337 (N_4337,N_3819,N_3973);
xor U4338 (N_4338,N_3719,N_3820);
nand U4339 (N_4339,N_3952,N_3894);
and U4340 (N_4340,N_3556,N_3706);
and U4341 (N_4341,N_3738,N_3875);
or U4342 (N_4342,N_3811,N_3534);
or U4343 (N_4343,N_3723,N_3920);
nand U4344 (N_4344,N_3647,N_3826);
nand U4345 (N_4345,N_3895,N_3514);
nand U4346 (N_4346,N_3766,N_3536);
nor U4347 (N_4347,N_3897,N_3526);
or U4348 (N_4348,N_3684,N_3687);
nand U4349 (N_4349,N_3702,N_3747);
xnor U4350 (N_4350,N_3804,N_3763);
nor U4351 (N_4351,N_3904,N_3550);
xor U4352 (N_4352,N_3655,N_3804);
and U4353 (N_4353,N_3943,N_3578);
nor U4354 (N_4354,N_3735,N_3555);
and U4355 (N_4355,N_3728,N_3930);
nor U4356 (N_4356,N_3583,N_3606);
and U4357 (N_4357,N_3856,N_3538);
or U4358 (N_4358,N_3940,N_3786);
xnor U4359 (N_4359,N_3713,N_3835);
and U4360 (N_4360,N_3634,N_3562);
or U4361 (N_4361,N_3581,N_3757);
or U4362 (N_4362,N_3830,N_3839);
nor U4363 (N_4363,N_3690,N_3901);
or U4364 (N_4364,N_3598,N_3800);
or U4365 (N_4365,N_3795,N_3926);
xor U4366 (N_4366,N_3979,N_3557);
nor U4367 (N_4367,N_3909,N_3602);
nor U4368 (N_4368,N_3622,N_3919);
nand U4369 (N_4369,N_3943,N_3947);
and U4370 (N_4370,N_3744,N_3920);
or U4371 (N_4371,N_3702,N_3822);
and U4372 (N_4372,N_3952,N_3935);
nor U4373 (N_4373,N_3564,N_3850);
xor U4374 (N_4374,N_3940,N_3953);
xnor U4375 (N_4375,N_3918,N_3994);
or U4376 (N_4376,N_3593,N_3742);
xor U4377 (N_4377,N_3885,N_3591);
and U4378 (N_4378,N_3539,N_3645);
nand U4379 (N_4379,N_3933,N_3666);
or U4380 (N_4380,N_3652,N_3752);
and U4381 (N_4381,N_3819,N_3506);
and U4382 (N_4382,N_3869,N_3905);
nor U4383 (N_4383,N_3730,N_3525);
nor U4384 (N_4384,N_3819,N_3730);
nand U4385 (N_4385,N_3507,N_3680);
nor U4386 (N_4386,N_3623,N_3908);
or U4387 (N_4387,N_3635,N_3962);
or U4388 (N_4388,N_3704,N_3667);
or U4389 (N_4389,N_3815,N_3529);
or U4390 (N_4390,N_3891,N_3734);
xnor U4391 (N_4391,N_3545,N_3689);
or U4392 (N_4392,N_3737,N_3772);
and U4393 (N_4393,N_3933,N_3835);
nand U4394 (N_4394,N_3565,N_3889);
and U4395 (N_4395,N_3768,N_3682);
nand U4396 (N_4396,N_3786,N_3922);
xnor U4397 (N_4397,N_3662,N_3779);
nor U4398 (N_4398,N_3546,N_3907);
xnor U4399 (N_4399,N_3801,N_3589);
xnor U4400 (N_4400,N_3877,N_3643);
nand U4401 (N_4401,N_3744,N_3531);
nand U4402 (N_4402,N_3772,N_3822);
nand U4403 (N_4403,N_3537,N_3751);
nor U4404 (N_4404,N_3874,N_3542);
and U4405 (N_4405,N_3746,N_3628);
xnor U4406 (N_4406,N_3548,N_3510);
or U4407 (N_4407,N_3853,N_3750);
xor U4408 (N_4408,N_3551,N_3614);
nor U4409 (N_4409,N_3946,N_3725);
nand U4410 (N_4410,N_3568,N_3808);
nor U4411 (N_4411,N_3801,N_3595);
or U4412 (N_4412,N_3954,N_3647);
or U4413 (N_4413,N_3783,N_3951);
nand U4414 (N_4414,N_3747,N_3555);
xor U4415 (N_4415,N_3791,N_3509);
and U4416 (N_4416,N_3977,N_3780);
or U4417 (N_4417,N_3653,N_3961);
nand U4418 (N_4418,N_3998,N_3926);
or U4419 (N_4419,N_3604,N_3730);
xnor U4420 (N_4420,N_3922,N_3562);
or U4421 (N_4421,N_3881,N_3592);
nor U4422 (N_4422,N_3844,N_3800);
xor U4423 (N_4423,N_3577,N_3830);
xor U4424 (N_4424,N_3519,N_3692);
and U4425 (N_4425,N_3992,N_3898);
or U4426 (N_4426,N_3559,N_3558);
and U4427 (N_4427,N_3862,N_3781);
nor U4428 (N_4428,N_3798,N_3722);
or U4429 (N_4429,N_3863,N_3519);
or U4430 (N_4430,N_3892,N_3749);
and U4431 (N_4431,N_3602,N_3571);
or U4432 (N_4432,N_3779,N_3892);
nor U4433 (N_4433,N_3930,N_3694);
and U4434 (N_4434,N_3829,N_3766);
or U4435 (N_4435,N_3753,N_3709);
nor U4436 (N_4436,N_3682,N_3905);
nor U4437 (N_4437,N_3720,N_3919);
nand U4438 (N_4438,N_3639,N_3606);
or U4439 (N_4439,N_3630,N_3858);
nand U4440 (N_4440,N_3666,N_3964);
and U4441 (N_4441,N_3998,N_3584);
xnor U4442 (N_4442,N_3825,N_3643);
or U4443 (N_4443,N_3972,N_3642);
and U4444 (N_4444,N_3686,N_3753);
xor U4445 (N_4445,N_3880,N_3773);
nor U4446 (N_4446,N_3869,N_3648);
xnor U4447 (N_4447,N_3815,N_3767);
or U4448 (N_4448,N_3551,N_3647);
nand U4449 (N_4449,N_3764,N_3590);
xor U4450 (N_4450,N_3911,N_3904);
xor U4451 (N_4451,N_3610,N_3597);
or U4452 (N_4452,N_3699,N_3587);
xor U4453 (N_4453,N_3737,N_3932);
nor U4454 (N_4454,N_3833,N_3660);
nor U4455 (N_4455,N_3623,N_3712);
xor U4456 (N_4456,N_3596,N_3594);
nand U4457 (N_4457,N_3703,N_3900);
and U4458 (N_4458,N_3827,N_3644);
nor U4459 (N_4459,N_3710,N_3991);
and U4460 (N_4460,N_3526,N_3555);
nand U4461 (N_4461,N_3859,N_3944);
and U4462 (N_4462,N_3522,N_3783);
nand U4463 (N_4463,N_3571,N_3878);
nand U4464 (N_4464,N_3564,N_3585);
nor U4465 (N_4465,N_3686,N_3504);
and U4466 (N_4466,N_3905,N_3692);
or U4467 (N_4467,N_3854,N_3919);
nand U4468 (N_4468,N_3691,N_3611);
and U4469 (N_4469,N_3562,N_3665);
xor U4470 (N_4470,N_3574,N_3610);
or U4471 (N_4471,N_3639,N_3527);
xor U4472 (N_4472,N_3944,N_3567);
or U4473 (N_4473,N_3660,N_3663);
or U4474 (N_4474,N_3813,N_3892);
and U4475 (N_4475,N_3634,N_3959);
and U4476 (N_4476,N_3644,N_3915);
or U4477 (N_4477,N_3807,N_3684);
xor U4478 (N_4478,N_3753,N_3557);
xnor U4479 (N_4479,N_3856,N_3767);
nor U4480 (N_4480,N_3898,N_3583);
nand U4481 (N_4481,N_3751,N_3513);
xnor U4482 (N_4482,N_3860,N_3933);
or U4483 (N_4483,N_3765,N_3746);
nand U4484 (N_4484,N_3987,N_3922);
xnor U4485 (N_4485,N_3549,N_3814);
nand U4486 (N_4486,N_3826,N_3566);
nand U4487 (N_4487,N_3896,N_3566);
or U4488 (N_4488,N_3826,N_3657);
xnor U4489 (N_4489,N_3744,N_3542);
nand U4490 (N_4490,N_3984,N_3565);
xnor U4491 (N_4491,N_3520,N_3734);
and U4492 (N_4492,N_3970,N_3503);
and U4493 (N_4493,N_3724,N_3983);
xnor U4494 (N_4494,N_3563,N_3864);
xnor U4495 (N_4495,N_3736,N_3620);
xor U4496 (N_4496,N_3535,N_3820);
or U4497 (N_4497,N_3703,N_3596);
nor U4498 (N_4498,N_3949,N_3728);
xnor U4499 (N_4499,N_3500,N_3604);
and U4500 (N_4500,N_4219,N_4325);
xnor U4501 (N_4501,N_4155,N_4279);
xor U4502 (N_4502,N_4093,N_4403);
and U4503 (N_4503,N_4020,N_4426);
and U4504 (N_4504,N_4493,N_4223);
or U4505 (N_4505,N_4470,N_4035);
nand U4506 (N_4506,N_4287,N_4388);
nor U4507 (N_4507,N_4006,N_4289);
xor U4508 (N_4508,N_4113,N_4324);
and U4509 (N_4509,N_4402,N_4045);
nor U4510 (N_4510,N_4248,N_4183);
xnor U4511 (N_4511,N_4476,N_4356);
nand U4512 (N_4512,N_4185,N_4122);
nand U4513 (N_4513,N_4283,N_4420);
and U4514 (N_4514,N_4036,N_4332);
nor U4515 (N_4515,N_4226,N_4267);
xnor U4516 (N_4516,N_4444,N_4489);
xnor U4517 (N_4517,N_4172,N_4018);
and U4518 (N_4518,N_4451,N_4186);
or U4519 (N_4519,N_4319,N_4256);
and U4520 (N_4520,N_4382,N_4178);
nor U4521 (N_4521,N_4247,N_4021);
and U4522 (N_4522,N_4378,N_4288);
nor U4523 (N_4523,N_4410,N_4061);
nor U4524 (N_4524,N_4038,N_4480);
nand U4525 (N_4525,N_4238,N_4157);
nand U4526 (N_4526,N_4235,N_4386);
nor U4527 (N_4527,N_4384,N_4204);
and U4528 (N_4528,N_4068,N_4056);
xor U4529 (N_4529,N_4145,N_4102);
nor U4530 (N_4530,N_4422,N_4269);
or U4531 (N_4531,N_4387,N_4337);
nor U4532 (N_4532,N_4177,N_4207);
nor U4533 (N_4533,N_4486,N_4270);
and U4534 (N_4534,N_4435,N_4355);
nor U4535 (N_4535,N_4492,N_4290);
xor U4536 (N_4536,N_4174,N_4187);
or U4537 (N_4537,N_4499,N_4465);
nor U4538 (N_4538,N_4014,N_4459);
nand U4539 (N_4539,N_4165,N_4398);
nand U4540 (N_4540,N_4468,N_4220);
xnor U4541 (N_4541,N_4043,N_4010);
or U4542 (N_4542,N_4280,N_4066);
nand U4543 (N_4543,N_4253,N_4329);
or U4544 (N_4544,N_4494,N_4141);
xnor U4545 (N_4545,N_4005,N_4277);
and U4546 (N_4546,N_4026,N_4338);
or U4547 (N_4547,N_4193,N_4362);
nand U4548 (N_4548,N_4110,N_4379);
xor U4549 (N_4549,N_4366,N_4104);
nor U4550 (N_4550,N_4404,N_4222);
or U4551 (N_4551,N_4063,N_4371);
xor U4552 (N_4552,N_4128,N_4351);
nand U4553 (N_4553,N_4027,N_4249);
nor U4554 (N_4554,N_4022,N_4159);
nor U4555 (N_4555,N_4138,N_4368);
nand U4556 (N_4556,N_4042,N_4450);
and U4557 (N_4557,N_4359,N_4051);
nor U4558 (N_4558,N_4413,N_4312);
and U4559 (N_4559,N_4437,N_4100);
or U4560 (N_4560,N_4472,N_4019);
or U4561 (N_4561,N_4184,N_4111);
nor U4562 (N_4562,N_4481,N_4206);
nand U4563 (N_4563,N_4408,N_4461);
and U4564 (N_4564,N_4399,N_4152);
nor U4565 (N_4565,N_4372,N_4103);
or U4566 (N_4566,N_4041,N_4254);
or U4567 (N_4567,N_4430,N_4439);
nand U4568 (N_4568,N_4134,N_4080);
or U4569 (N_4569,N_4455,N_4300);
and U4570 (N_4570,N_4032,N_4101);
and U4571 (N_4571,N_4213,N_4483);
or U4572 (N_4572,N_4030,N_4394);
nand U4573 (N_4573,N_4214,N_4092);
nand U4574 (N_4574,N_4469,N_4234);
and U4575 (N_4575,N_4487,N_4322);
nand U4576 (N_4576,N_4278,N_4129);
and U4577 (N_4577,N_4390,N_4286);
nor U4578 (N_4578,N_4175,N_4268);
or U4579 (N_4579,N_4428,N_4391);
and U4580 (N_4580,N_4471,N_4393);
nor U4581 (N_4581,N_4447,N_4331);
xnor U4582 (N_4582,N_4415,N_4085);
or U4583 (N_4583,N_4004,N_4306);
xor U4584 (N_4584,N_4054,N_4373);
nand U4585 (N_4585,N_4064,N_4297);
nand U4586 (N_4586,N_4412,N_4317);
and U4587 (N_4587,N_4293,N_4143);
xnor U4588 (N_4588,N_4230,N_4243);
nor U4589 (N_4589,N_4257,N_4370);
xnor U4590 (N_4590,N_4115,N_4137);
nor U4591 (N_4591,N_4473,N_4136);
nor U4592 (N_4592,N_4154,N_4215);
or U4593 (N_4593,N_4160,N_4442);
nand U4594 (N_4594,N_4158,N_4212);
or U4595 (N_4595,N_4191,N_4417);
and U4596 (N_4596,N_4485,N_4446);
nand U4597 (N_4597,N_4496,N_4484);
nand U4598 (N_4598,N_4203,N_4292);
or U4599 (N_4599,N_4168,N_4491);
xnor U4600 (N_4600,N_4281,N_4360);
or U4601 (N_4601,N_4313,N_4327);
or U4602 (N_4602,N_4139,N_4350);
and U4603 (N_4603,N_4199,N_4252);
nand U4604 (N_4604,N_4424,N_4082);
nor U4605 (N_4605,N_4105,N_4315);
and U4606 (N_4606,N_4448,N_4088);
xnor U4607 (N_4607,N_4369,N_4376);
or U4608 (N_4608,N_4016,N_4255);
nor U4609 (N_4609,N_4169,N_4040);
xnor U4610 (N_4610,N_4309,N_4414);
and U4611 (N_4611,N_4416,N_4049);
xor U4612 (N_4612,N_4344,N_4340);
xnor U4613 (N_4613,N_4326,N_4334);
or U4614 (N_4614,N_4454,N_4335);
nor U4615 (N_4615,N_4000,N_4140);
nor U4616 (N_4616,N_4072,N_4003);
and U4617 (N_4617,N_4098,N_4339);
or U4618 (N_4618,N_4440,N_4421);
nand U4619 (N_4619,N_4071,N_4303);
and U4620 (N_4620,N_4112,N_4478);
xor U4621 (N_4621,N_4001,N_4374);
and U4622 (N_4622,N_4272,N_4176);
or U4623 (N_4623,N_4017,N_4050);
or U4624 (N_4624,N_4179,N_4405);
or U4625 (N_4625,N_4271,N_4125);
xor U4626 (N_4626,N_4198,N_4133);
nand U4627 (N_4627,N_4062,N_4084);
nor U4628 (N_4628,N_4224,N_4182);
and U4629 (N_4629,N_4298,N_4342);
xnor U4630 (N_4630,N_4095,N_4047);
nor U4631 (N_4631,N_4314,N_4434);
nor U4632 (N_4632,N_4096,N_4411);
or U4633 (N_4633,N_4089,N_4211);
xor U4634 (N_4634,N_4239,N_4033);
and U4635 (N_4635,N_4012,N_4029);
or U4636 (N_4636,N_4008,N_4353);
and U4637 (N_4637,N_4090,N_4246);
and U4638 (N_4638,N_4094,N_4304);
nand U4639 (N_4639,N_4131,N_4354);
and U4640 (N_4640,N_4261,N_4273);
nor U4641 (N_4641,N_4197,N_4087);
xor U4642 (N_4642,N_4341,N_4052);
nor U4643 (N_4643,N_4463,N_4449);
nand U4644 (N_4644,N_4119,N_4190);
nand U4645 (N_4645,N_4395,N_4156);
and U4646 (N_4646,N_4400,N_4218);
and U4647 (N_4647,N_4167,N_4381);
and U4648 (N_4648,N_4189,N_4299);
xor U4649 (N_4649,N_4423,N_4196);
or U4650 (N_4650,N_4295,N_4144);
or U4651 (N_4651,N_4067,N_4282);
and U4652 (N_4652,N_4039,N_4228);
xnor U4653 (N_4653,N_4466,N_4409);
xnor U4654 (N_4654,N_4028,N_4233);
nand U4655 (N_4655,N_4429,N_4251);
xor U4656 (N_4656,N_4109,N_4148);
nor U4657 (N_4657,N_4241,N_4240);
and U4658 (N_4658,N_4146,N_4121);
or U4659 (N_4659,N_4445,N_4441);
and U4660 (N_4660,N_4229,N_4117);
or U4661 (N_4661,N_4132,N_4227);
xor U4662 (N_4662,N_4107,N_4361);
nand U4663 (N_4663,N_4192,N_4275);
nor U4664 (N_4664,N_4392,N_4310);
nor U4665 (N_4665,N_4364,N_4209);
nor U4666 (N_4666,N_4078,N_4232);
nor U4667 (N_4667,N_4116,N_4336);
nor U4668 (N_4668,N_4318,N_4173);
nor U4669 (N_4669,N_4023,N_4285);
nand U4670 (N_4670,N_4163,N_4320);
and U4671 (N_4671,N_4210,N_4118);
or U4672 (N_4672,N_4407,N_4086);
nor U4673 (N_4673,N_4345,N_4477);
nor U4674 (N_4674,N_4301,N_4180);
xor U4675 (N_4675,N_4365,N_4266);
and U4676 (N_4676,N_4059,N_4048);
or U4677 (N_4677,N_4436,N_4377);
nand U4678 (N_4678,N_4108,N_4343);
or U4679 (N_4679,N_4161,N_4076);
and U4680 (N_4680,N_4147,N_4221);
nor U4681 (N_4681,N_4053,N_4151);
or U4682 (N_4682,N_4188,N_4242);
nor U4683 (N_4683,N_4034,N_4075);
xor U4684 (N_4684,N_4205,N_4396);
and U4685 (N_4685,N_4262,N_4367);
xnor U4686 (N_4686,N_4120,N_4024);
nand U4687 (N_4687,N_4316,N_4418);
or U4688 (N_4688,N_4419,N_4467);
xor U4689 (N_4689,N_4091,N_4401);
xor U4690 (N_4690,N_4258,N_4456);
nor U4691 (N_4691,N_4291,N_4225);
xnor U4692 (N_4692,N_4311,N_4495);
and U4693 (N_4693,N_4244,N_4352);
or U4694 (N_4694,N_4263,N_4305);
nor U4695 (N_4695,N_4202,N_4328);
xor U4696 (N_4696,N_4363,N_4060);
xnor U4697 (N_4697,N_4259,N_4482);
or U4698 (N_4698,N_4046,N_4025);
and U4699 (N_4699,N_4069,N_4260);
and U4700 (N_4700,N_4201,N_4479);
nand U4701 (N_4701,N_4077,N_4217);
and U4702 (N_4702,N_4250,N_4181);
nand U4703 (N_4703,N_4037,N_4127);
xnor U4704 (N_4704,N_4498,N_4427);
and U4705 (N_4705,N_4323,N_4079);
or U4706 (N_4706,N_4044,N_4149);
nor U4707 (N_4707,N_4081,N_4106);
or U4708 (N_4708,N_4015,N_4236);
nor U4709 (N_4709,N_4380,N_4057);
or U4710 (N_4710,N_4308,N_4284);
and U4711 (N_4711,N_4490,N_4142);
xor U4712 (N_4712,N_4348,N_4457);
nand U4713 (N_4713,N_4074,N_4123);
and U4714 (N_4714,N_4274,N_4452);
nand U4715 (N_4715,N_4130,N_4083);
nor U4716 (N_4716,N_4296,N_4265);
nand U4717 (N_4717,N_4432,N_4302);
nand U4718 (N_4718,N_4195,N_4347);
xor U4719 (N_4719,N_4200,N_4099);
nor U4720 (N_4720,N_4346,N_4124);
xor U4721 (N_4721,N_4497,N_4488);
xor U4722 (N_4722,N_4358,N_4031);
or U4723 (N_4723,N_4126,N_4065);
xor U4724 (N_4724,N_4164,N_4460);
or U4725 (N_4725,N_4475,N_4002);
nor U4726 (N_4726,N_4433,N_4166);
and U4727 (N_4727,N_4055,N_4194);
nor U4728 (N_4728,N_4385,N_4438);
xor U4729 (N_4729,N_4237,N_4389);
nor U4730 (N_4730,N_4458,N_4231);
and U4731 (N_4731,N_4208,N_4330);
nor U4732 (N_4732,N_4307,N_4153);
xnor U4733 (N_4733,N_4150,N_4333);
nor U4734 (N_4734,N_4349,N_4464);
nand U4735 (N_4735,N_4058,N_4114);
and U4736 (N_4736,N_4245,N_4135);
nand U4737 (N_4737,N_4425,N_4443);
or U4738 (N_4738,N_4357,N_4294);
and U4739 (N_4739,N_4397,N_4073);
xnor U4740 (N_4740,N_4070,N_4162);
xnor U4741 (N_4741,N_4431,N_4171);
and U4742 (N_4742,N_4383,N_4264);
nor U4743 (N_4743,N_4216,N_4474);
and U4744 (N_4744,N_4276,N_4009);
xnor U4745 (N_4745,N_4453,N_4013);
and U4746 (N_4746,N_4097,N_4321);
or U4747 (N_4747,N_4406,N_4007);
nor U4748 (N_4748,N_4462,N_4375);
or U4749 (N_4749,N_4011,N_4170);
nand U4750 (N_4750,N_4266,N_4135);
xor U4751 (N_4751,N_4365,N_4475);
xnor U4752 (N_4752,N_4226,N_4308);
and U4753 (N_4753,N_4466,N_4172);
nand U4754 (N_4754,N_4025,N_4121);
nand U4755 (N_4755,N_4334,N_4032);
nor U4756 (N_4756,N_4331,N_4126);
or U4757 (N_4757,N_4388,N_4190);
nand U4758 (N_4758,N_4309,N_4480);
xor U4759 (N_4759,N_4228,N_4478);
or U4760 (N_4760,N_4063,N_4293);
nand U4761 (N_4761,N_4499,N_4444);
nor U4762 (N_4762,N_4079,N_4452);
and U4763 (N_4763,N_4240,N_4041);
xnor U4764 (N_4764,N_4093,N_4156);
nand U4765 (N_4765,N_4435,N_4275);
or U4766 (N_4766,N_4092,N_4240);
or U4767 (N_4767,N_4340,N_4213);
and U4768 (N_4768,N_4347,N_4198);
nor U4769 (N_4769,N_4176,N_4086);
nor U4770 (N_4770,N_4238,N_4462);
nand U4771 (N_4771,N_4030,N_4371);
nand U4772 (N_4772,N_4428,N_4197);
nand U4773 (N_4773,N_4046,N_4094);
and U4774 (N_4774,N_4331,N_4335);
xor U4775 (N_4775,N_4233,N_4311);
or U4776 (N_4776,N_4256,N_4405);
xnor U4777 (N_4777,N_4188,N_4169);
nand U4778 (N_4778,N_4184,N_4087);
xor U4779 (N_4779,N_4053,N_4285);
nand U4780 (N_4780,N_4411,N_4480);
nor U4781 (N_4781,N_4077,N_4043);
nand U4782 (N_4782,N_4295,N_4263);
nand U4783 (N_4783,N_4460,N_4154);
xnor U4784 (N_4784,N_4304,N_4019);
and U4785 (N_4785,N_4396,N_4416);
nor U4786 (N_4786,N_4293,N_4065);
nand U4787 (N_4787,N_4272,N_4300);
nor U4788 (N_4788,N_4232,N_4309);
xnor U4789 (N_4789,N_4377,N_4223);
nor U4790 (N_4790,N_4415,N_4438);
nand U4791 (N_4791,N_4135,N_4214);
and U4792 (N_4792,N_4076,N_4140);
nor U4793 (N_4793,N_4238,N_4095);
nor U4794 (N_4794,N_4055,N_4298);
nand U4795 (N_4795,N_4443,N_4347);
xor U4796 (N_4796,N_4053,N_4166);
and U4797 (N_4797,N_4297,N_4149);
and U4798 (N_4798,N_4029,N_4065);
xor U4799 (N_4799,N_4129,N_4176);
nor U4800 (N_4800,N_4312,N_4218);
nand U4801 (N_4801,N_4226,N_4313);
xnor U4802 (N_4802,N_4103,N_4434);
nand U4803 (N_4803,N_4430,N_4425);
and U4804 (N_4804,N_4251,N_4098);
and U4805 (N_4805,N_4011,N_4248);
nor U4806 (N_4806,N_4299,N_4013);
or U4807 (N_4807,N_4337,N_4183);
nor U4808 (N_4808,N_4236,N_4270);
or U4809 (N_4809,N_4413,N_4292);
or U4810 (N_4810,N_4031,N_4199);
xor U4811 (N_4811,N_4494,N_4264);
xor U4812 (N_4812,N_4070,N_4172);
nor U4813 (N_4813,N_4273,N_4383);
nor U4814 (N_4814,N_4034,N_4021);
nor U4815 (N_4815,N_4492,N_4326);
nand U4816 (N_4816,N_4103,N_4257);
nand U4817 (N_4817,N_4311,N_4005);
xnor U4818 (N_4818,N_4215,N_4392);
xnor U4819 (N_4819,N_4384,N_4398);
or U4820 (N_4820,N_4306,N_4057);
nor U4821 (N_4821,N_4047,N_4466);
xnor U4822 (N_4822,N_4397,N_4036);
nand U4823 (N_4823,N_4062,N_4066);
and U4824 (N_4824,N_4205,N_4157);
nor U4825 (N_4825,N_4233,N_4001);
nand U4826 (N_4826,N_4063,N_4081);
nor U4827 (N_4827,N_4482,N_4144);
or U4828 (N_4828,N_4301,N_4195);
nor U4829 (N_4829,N_4487,N_4277);
or U4830 (N_4830,N_4068,N_4305);
or U4831 (N_4831,N_4095,N_4044);
nor U4832 (N_4832,N_4213,N_4444);
xor U4833 (N_4833,N_4236,N_4383);
or U4834 (N_4834,N_4137,N_4100);
xor U4835 (N_4835,N_4439,N_4383);
xnor U4836 (N_4836,N_4375,N_4279);
nor U4837 (N_4837,N_4488,N_4376);
nand U4838 (N_4838,N_4315,N_4342);
or U4839 (N_4839,N_4414,N_4044);
nand U4840 (N_4840,N_4284,N_4295);
nand U4841 (N_4841,N_4005,N_4376);
and U4842 (N_4842,N_4078,N_4007);
xnor U4843 (N_4843,N_4466,N_4414);
nor U4844 (N_4844,N_4429,N_4205);
nand U4845 (N_4845,N_4258,N_4312);
xnor U4846 (N_4846,N_4022,N_4497);
or U4847 (N_4847,N_4039,N_4266);
or U4848 (N_4848,N_4034,N_4096);
nor U4849 (N_4849,N_4335,N_4017);
nor U4850 (N_4850,N_4403,N_4165);
nand U4851 (N_4851,N_4255,N_4454);
xnor U4852 (N_4852,N_4003,N_4134);
nor U4853 (N_4853,N_4005,N_4295);
xnor U4854 (N_4854,N_4093,N_4062);
nor U4855 (N_4855,N_4145,N_4472);
or U4856 (N_4856,N_4134,N_4107);
or U4857 (N_4857,N_4106,N_4300);
and U4858 (N_4858,N_4127,N_4120);
nor U4859 (N_4859,N_4011,N_4196);
or U4860 (N_4860,N_4149,N_4306);
nor U4861 (N_4861,N_4353,N_4285);
nand U4862 (N_4862,N_4109,N_4448);
nor U4863 (N_4863,N_4254,N_4361);
or U4864 (N_4864,N_4339,N_4470);
nor U4865 (N_4865,N_4193,N_4059);
xor U4866 (N_4866,N_4209,N_4311);
and U4867 (N_4867,N_4341,N_4263);
and U4868 (N_4868,N_4061,N_4322);
xor U4869 (N_4869,N_4272,N_4271);
nand U4870 (N_4870,N_4022,N_4089);
xor U4871 (N_4871,N_4143,N_4313);
or U4872 (N_4872,N_4246,N_4140);
nor U4873 (N_4873,N_4284,N_4418);
or U4874 (N_4874,N_4212,N_4054);
nor U4875 (N_4875,N_4033,N_4224);
or U4876 (N_4876,N_4210,N_4326);
nor U4877 (N_4877,N_4370,N_4209);
or U4878 (N_4878,N_4485,N_4124);
xnor U4879 (N_4879,N_4469,N_4075);
nor U4880 (N_4880,N_4192,N_4326);
or U4881 (N_4881,N_4187,N_4374);
xnor U4882 (N_4882,N_4394,N_4029);
xnor U4883 (N_4883,N_4435,N_4196);
or U4884 (N_4884,N_4232,N_4425);
xor U4885 (N_4885,N_4156,N_4396);
nand U4886 (N_4886,N_4244,N_4399);
nand U4887 (N_4887,N_4270,N_4362);
and U4888 (N_4888,N_4281,N_4182);
nand U4889 (N_4889,N_4043,N_4273);
nor U4890 (N_4890,N_4053,N_4002);
nand U4891 (N_4891,N_4413,N_4237);
nor U4892 (N_4892,N_4038,N_4011);
or U4893 (N_4893,N_4487,N_4111);
xor U4894 (N_4894,N_4089,N_4213);
nand U4895 (N_4895,N_4253,N_4219);
nand U4896 (N_4896,N_4125,N_4378);
nor U4897 (N_4897,N_4187,N_4331);
xnor U4898 (N_4898,N_4416,N_4369);
nand U4899 (N_4899,N_4152,N_4096);
nand U4900 (N_4900,N_4349,N_4144);
or U4901 (N_4901,N_4273,N_4473);
nor U4902 (N_4902,N_4124,N_4437);
and U4903 (N_4903,N_4337,N_4381);
xnor U4904 (N_4904,N_4205,N_4446);
nand U4905 (N_4905,N_4089,N_4084);
nor U4906 (N_4906,N_4326,N_4124);
nand U4907 (N_4907,N_4181,N_4347);
or U4908 (N_4908,N_4367,N_4310);
and U4909 (N_4909,N_4275,N_4323);
nand U4910 (N_4910,N_4104,N_4286);
or U4911 (N_4911,N_4386,N_4304);
and U4912 (N_4912,N_4474,N_4159);
and U4913 (N_4913,N_4405,N_4065);
xor U4914 (N_4914,N_4133,N_4058);
or U4915 (N_4915,N_4494,N_4244);
or U4916 (N_4916,N_4325,N_4361);
xnor U4917 (N_4917,N_4336,N_4361);
and U4918 (N_4918,N_4134,N_4377);
or U4919 (N_4919,N_4023,N_4109);
xnor U4920 (N_4920,N_4389,N_4010);
nor U4921 (N_4921,N_4174,N_4274);
xnor U4922 (N_4922,N_4165,N_4383);
nand U4923 (N_4923,N_4284,N_4484);
nor U4924 (N_4924,N_4493,N_4338);
nand U4925 (N_4925,N_4151,N_4483);
or U4926 (N_4926,N_4356,N_4248);
nor U4927 (N_4927,N_4374,N_4040);
xnor U4928 (N_4928,N_4095,N_4066);
or U4929 (N_4929,N_4350,N_4279);
or U4930 (N_4930,N_4191,N_4437);
and U4931 (N_4931,N_4255,N_4432);
or U4932 (N_4932,N_4330,N_4289);
or U4933 (N_4933,N_4142,N_4263);
nor U4934 (N_4934,N_4354,N_4469);
nor U4935 (N_4935,N_4284,N_4270);
or U4936 (N_4936,N_4264,N_4291);
nand U4937 (N_4937,N_4138,N_4373);
nor U4938 (N_4938,N_4466,N_4343);
nor U4939 (N_4939,N_4208,N_4422);
nand U4940 (N_4940,N_4197,N_4129);
nand U4941 (N_4941,N_4143,N_4418);
nor U4942 (N_4942,N_4356,N_4354);
or U4943 (N_4943,N_4000,N_4247);
nor U4944 (N_4944,N_4239,N_4214);
nor U4945 (N_4945,N_4230,N_4251);
nand U4946 (N_4946,N_4371,N_4142);
and U4947 (N_4947,N_4459,N_4062);
nand U4948 (N_4948,N_4226,N_4297);
nor U4949 (N_4949,N_4100,N_4099);
nand U4950 (N_4950,N_4388,N_4259);
nand U4951 (N_4951,N_4356,N_4153);
nor U4952 (N_4952,N_4251,N_4250);
nand U4953 (N_4953,N_4010,N_4111);
xor U4954 (N_4954,N_4222,N_4376);
or U4955 (N_4955,N_4056,N_4454);
nor U4956 (N_4956,N_4047,N_4492);
xnor U4957 (N_4957,N_4181,N_4066);
nand U4958 (N_4958,N_4375,N_4355);
and U4959 (N_4959,N_4457,N_4188);
nor U4960 (N_4960,N_4207,N_4156);
and U4961 (N_4961,N_4362,N_4363);
and U4962 (N_4962,N_4009,N_4363);
xor U4963 (N_4963,N_4082,N_4426);
xor U4964 (N_4964,N_4089,N_4251);
and U4965 (N_4965,N_4276,N_4449);
xor U4966 (N_4966,N_4377,N_4251);
xor U4967 (N_4967,N_4248,N_4450);
or U4968 (N_4968,N_4459,N_4306);
nand U4969 (N_4969,N_4111,N_4433);
and U4970 (N_4970,N_4194,N_4276);
nand U4971 (N_4971,N_4094,N_4344);
and U4972 (N_4972,N_4016,N_4126);
nand U4973 (N_4973,N_4311,N_4111);
and U4974 (N_4974,N_4425,N_4012);
xnor U4975 (N_4975,N_4016,N_4420);
or U4976 (N_4976,N_4108,N_4258);
and U4977 (N_4977,N_4498,N_4095);
nor U4978 (N_4978,N_4158,N_4243);
or U4979 (N_4979,N_4189,N_4043);
nor U4980 (N_4980,N_4117,N_4137);
nand U4981 (N_4981,N_4112,N_4028);
xnor U4982 (N_4982,N_4002,N_4473);
xor U4983 (N_4983,N_4326,N_4378);
xnor U4984 (N_4984,N_4018,N_4015);
xor U4985 (N_4985,N_4070,N_4313);
nand U4986 (N_4986,N_4261,N_4366);
nor U4987 (N_4987,N_4445,N_4211);
and U4988 (N_4988,N_4467,N_4133);
nand U4989 (N_4989,N_4006,N_4103);
xnor U4990 (N_4990,N_4104,N_4257);
and U4991 (N_4991,N_4334,N_4499);
nand U4992 (N_4992,N_4141,N_4149);
nand U4993 (N_4993,N_4425,N_4356);
xnor U4994 (N_4994,N_4385,N_4041);
xor U4995 (N_4995,N_4358,N_4205);
xor U4996 (N_4996,N_4454,N_4127);
nor U4997 (N_4997,N_4010,N_4174);
or U4998 (N_4998,N_4292,N_4012);
nor U4999 (N_4999,N_4130,N_4200);
or U5000 (N_5000,N_4625,N_4647);
or U5001 (N_5001,N_4990,N_4862);
xnor U5002 (N_5002,N_4919,N_4787);
and U5003 (N_5003,N_4558,N_4732);
nor U5004 (N_5004,N_4772,N_4511);
nand U5005 (N_5005,N_4945,N_4950);
nand U5006 (N_5006,N_4626,N_4559);
nand U5007 (N_5007,N_4624,N_4810);
or U5008 (N_5008,N_4578,N_4582);
xor U5009 (N_5009,N_4649,N_4727);
nor U5010 (N_5010,N_4673,N_4991);
nand U5011 (N_5011,N_4640,N_4526);
nor U5012 (N_5012,N_4946,N_4937);
and U5013 (N_5013,N_4980,N_4829);
and U5014 (N_5014,N_4885,N_4634);
nor U5015 (N_5015,N_4739,N_4948);
nor U5016 (N_5016,N_4508,N_4910);
xor U5017 (N_5017,N_4738,N_4823);
nand U5018 (N_5018,N_4963,N_4541);
and U5019 (N_5019,N_4944,N_4675);
xnor U5020 (N_5020,N_4602,N_4960);
and U5021 (N_5021,N_4533,N_4549);
xor U5022 (N_5022,N_4590,N_4763);
xor U5023 (N_5023,N_4598,N_4712);
nor U5024 (N_5024,N_4908,N_4722);
nor U5025 (N_5025,N_4537,N_4695);
nand U5026 (N_5026,N_4627,N_4791);
nor U5027 (N_5027,N_4755,N_4706);
and U5028 (N_5028,N_4663,N_4502);
nand U5029 (N_5029,N_4790,N_4825);
or U5030 (N_5030,N_4971,N_4645);
nor U5031 (N_5031,N_4633,N_4788);
or U5032 (N_5032,N_4740,N_4761);
or U5033 (N_5033,N_4674,N_4561);
or U5034 (N_5034,N_4799,N_4857);
and U5035 (N_5035,N_4691,N_4892);
or U5036 (N_5036,N_4643,N_4547);
or U5037 (N_5037,N_4539,N_4966);
or U5038 (N_5038,N_4701,N_4782);
or U5039 (N_5039,N_4965,N_4891);
nand U5040 (N_5040,N_4655,N_4893);
nand U5041 (N_5041,N_4976,N_4784);
nor U5042 (N_5042,N_4979,N_4583);
nand U5043 (N_5043,N_4593,N_4835);
xor U5044 (N_5044,N_4959,N_4708);
and U5045 (N_5045,N_4619,N_4653);
nand U5046 (N_5046,N_4664,N_4877);
nor U5047 (N_5047,N_4756,N_4843);
nand U5048 (N_5048,N_4913,N_4770);
nand U5049 (N_5049,N_4571,N_4716);
xor U5050 (N_5050,N_4630,N_4592);
and U5051 (N_5051,N_4648,N_4978);
and U5052 (N_5052,N_4639,N_4748);
xor U5053 (N_5053,N_4972,N_4607);
and U5054 (N_5054,N_4641,N_4928);
and U5055 (N_5055,N_4860,N_4753);
and U5056 (N_5056,N_4830,N_4730);
and U5057 (N_5057,N_4528,N_4514);
nand U5058 (N_5058,N_4994,N_4702);
or U5059 (N_5059,N_4737,N_4551);
nand U5060 (N_5060,N_4831,N_4882);
nor U5061 (N_5061,N_4520,N_4690);
and U5062 (N_5062,N_4769,N_4778);
and U5063 (N_5063,N_4905,N_4609);
or U5064 (N_5064,N_4826,N_4524);
xnor U5065 (N_5065,N_4926,N_4855);
and U5066 (N_5066,N_4838,N_4713);
or U5067 (N_5067,N_4970,N_4934);
xnor U5068 (N_5068,N_4556,N_4767);
or U5069 (N_5069,N_4909,N_4768);
xor U5070 (N_5070,N_4506,N_4509);
and U5071 (N_5071,N_4554,N_4816);
and U5072 (N_5072,N_4523,N_4588);
and U5073 (N_5073,N_4985,N_4989);
nand U5074 (N_5074,N_4773,N_4765);
nand U5075 (N_5075,N_4600,N_4747);
or U5076 (N_5076,N_4605,N_4819);
nand U5077 (N_5077,N_4595,N_4660);
nor U5078 (N_5078,N_4557,N_4513);
and U5079 (N_5079,N_4760,N_4943);
or U5080 (N_5080,N_4570,N_4845);
nor U5081 (N_5081,N_4581,N_4572);
nand U5082 (N_5082,N_4591,N_4646);
or U5083 (N_5083,N_4589,N_4642);
and U5084 (N_5084,N_4665,N_4846);
nand U5085 (N_5085,N_4775,N_4900);
and U5086 (N_5086,N_4873,N_4552);
xor U5087 (N_5087,N_4711,N_4780);
or U5088 (N_5088,N_4697,N_4656);
or U5089 (N_5089,N_4856,N_4839);
nor U5090 (N_5090,N_4563,N_4543);
nand U5091 (N_5091,N_4682,N_4901);
xor U5092 (N_5092,N_4516,N_4529);
nor U5093 (N_5093,N_4721,N_4569);
or U5094 (N_5094,N_4916,N_4638);
xor U5095 (N_5095,N_4870,N_4661);
and U5096 (N_5096,N_4903,N_4704);
nor U5097 (N_5097,N_4566,N_4568);
nor U5098 (N_5098,N_4872,N_4813);
or U5099 (N_5099,N_4883,N_4923);
and U5100 (N_5100,N_4610,N_4745);
nor U5101 (N_5101,N_4703,N_4612);
nor U5102 (N_5102,N_4844,N_4601);
nand U5103 (N_5103,N_4801,N_4505);
or U5104 (N_5104,N_4623,N_4785);
and U5105 (N_5105,N_4938,N_4743);
nand U5106 (N_5106,N_4837,N_4676);
xnor U5107 (N_5107,N_4951,N_4798);
and U5108 (N_5108,N_4918,N_4658);
nand U5109 (N_5109,N_4876,N_4973);
and U5110 (N_5110,N_4710,N_4828);
and U5111 (N_5111,N_4930,N_4726);
or U5112 (N_5112,N_4820,N_4988);
and U5113 (N_5113,N_4929,N_4954);
nor U5114 (N_5114,N_4977,N_4999);
nor U5115 (N_5115,N_4808,N_4789);
nor U5116 (N_5116,N_4781,N_4847);
nor U5117 (N_5117,N_4874,N_4729);
nor U5118 (N_5118,N_4632,N_4955);
nand U5119 (N_5119,N_4853,N_4672);
nor U5120 (N_5120,N_4577,N_4961);
nand U5121 (N_5121,N_4548,N_4709);
or U5122 (N_5122,N_4987,N_4530);
xnor U5123 (N_5123,N_4503,N_4925);
xnor U5124 (N_5124,N_4636,N_4594);
xnor U5125 (N_5125,N_4869,N_4565);
xor U5126 (N_5126,N_4757,N_4654);
xnor U5127 (N_5127,N_4797,N_4504);
xor U5128 (N_5128,N_4501,N_4817);
and U5129 (N_5129,N_4546,N_4827);
and U5130 (N_5130,N_4993,N_4678);
or U5131 (N_5131,N_4515,N_4628);
nor U5132 (N_5132,N_4604,N_4670);
and U5133 (N_5133,N_4952,N_4814);
or U5134 (N_5134,N_4841,N_4890);
nor U5135 (N_5135,N_4939,N_4544);
nor U5136 (N_5136,N_4957,N_4834);
nor U5137 (N_5137,N_4806,N_4906);
nand U5138 (N_5138,N_4720,N_4824);
nand U5139 (N_5139,N_4807,N_4680);
and U5140 (N_5140,N_4766,N_4519);
xnor U5141 (N_5141,N_4685,N_4983);
nor U5142 (N_5142,N_4956,N_4852);
nand U5143 (N_5143,N_4687,N_4764);
nand U5144 (N_5144,N_4863,N_4736);
nand U5145 (N_5145,N_4881,N_4567);
nor U5146 (N_5146,N_4671,N_4718);
nor U5147 (N_5147,N_4725,N_4811);
nor U5148 (N_5148,N_4586,N_4936);
or U5149 (N_5149,N_4880,N_4611);
xnor U5150 (N_5150,N_4538,N_4606);
xnor U5151 (N_5151,N_4500,N_4620);
nand U5152 (N_5152,N_4861,N_4849);
or U5153 (N_5153,N_4836,N_4894);
or U5154 (N_5154,N_4562,N_4777);
or U5155 (N_5155,N_4662,N_4758);
nor U5156 (N_5156,N_4992,N_4522);
or U5157 (N_5157,N_4545,N_4584);
nor U5158 (N_5158,N_4996,N_4677);
nand U5159 (N_5159,N_4652,N_4599);
nor U5160 (N_5160,N_4684,N_4510);
and U5161 (N_5161,N_4868,N_4746);
and U5162 (N_5162,N_4866,N_4986);
xor U5163 (N_5163,N_4618,N_4962);
xnor U5164 (N_5164,N_4686,N_4527);
nor U5165 (N_5165,N_4832,N_4750);
nand U5166 (N_5166,N_4532,N_4507);
and U5167 (N_5167,N_4560,N_4714);
or U5168 (N_5168,N_4735,N_4724);
xor U5169 (N_5169,N_4783,N_4805);
nand U5170 (N_5170,N_4555,N_4698);
or U5171 (N_5171,N_4617,N_4749);
xor U5172 (N_5172,N_4800,N_4969);
xnor U5173 (N_5173,N_4981,N_4719);
xor U5174 (N_5174,N_4953,N_4603);
xnor U5175 (N_5175,N_4886,N_4637);
xor U5176 (N_5176,N_4751,N_4631);
xnor U5177 (N_5177,N_4580,N_4669);
nor U5178 (N_5178,N_4995,N_4614);
xnor U5179 (N_5179,N_4911,N_4897);
and U5180 (N_5180,N_4942,N_4613);
or U5181 (N_5181,N_4879,N_4967);
or U5182 (N_5182,N_4615,N_4899);
nand U5183 (N_5183,N_4888,N_4786);
or U5184 (N_5184,N_4752,N_4821);
or U5185 (N_5185,N_4848,N_4668);
xnor U5186 (N_5186,N_4809,N_4922);
nor U5187 (N_5187,N_4699,N_4635);
and U5188 (N_5188,N_4622,N_4793);
or U5189 (N_5189,N_4912,N_4689);
nand U5190 (N_5190,N_4576,N_4927);
nor U5191 (N_5191,N_4666,N_4754);
or U5192 (N_5192,N_4688,N_4964);
or U5193 (N_5193,N_4667,N_4812);
nor U5194 (N_5194,N_4958,N_4536);
and U5195 (N_5195,N_4657,N_4982);
or U5196 (N_5196,N_4840,N_4907);
or U5197 (N_5197,N_4728,N_4794);
nand U5198 (N_5198,N_4733,N_4917);
xor U5199 (N_5199,N_4744,N_4621);
nand U5200 (N_5200,N_4629,N_4884);
nor U5201 (N_5201,N_4776,N_4700);
nand U5202 (N_5202,N_4850,N_4898);
nor U5203 (N_5203,N_4596,N_4587);
nand U5204 (N_5204,N_4867,N_4521);
and U5205 (N_5205,N_4920,N_4887);
nand U5206 (N_5206,N_4715,N_4553);
nor U5207 (N_5207,N_4707,N_4651);
and U5208 (N_5208,N_4579,N_4875);
nand U5209 (N_5209,N_4842,N_4889);
nor U5210 (N_5210,N_4692,N_4742);
nand U5211 (N_5211,N_4644,N_4573);
or U5212 (N_5212,N_4535,N_4525);
or U5213 (N_5213,N_4693,N_4731);
xnor U5214 (N_5214,N_4796,N_4795);
and U5215 (N_5215,N_4531,N_4984);
xnor U5216 (N_5216,N_4681,N_4924);
nor U5217 (N_5217,N_4574,N_4914);
xor U5218 (N_5218,N_4803,N_4851);
xor U5219 (N_5219,N_4512,N_4542);
nor U5220 (N_5220,N_4774,N_4997);
nand U5221 (N_5221,N_4833,N_4650);
xnor U5222 (N_5222,N_4904,N_4616);
and U5223 (N_5223,N_4517,N_4815);
or U5224 (N_5224,N_4575,N_4822);
nand U5225 (N_5225,N_4802,N_4818);
nor U5226 (N_5226,N_4858,N_4723);
xor U5227 (N_5227,N_4878,N_4931);
nand U5228 (N_5228,N_4941,N_4871);
xnor U5229 (N_5229,N_4935,N_4968);
nand U5230 (N_5230,N_4659,N_4864);
nor U5231 (N_5231,N_4792,N_4694);
nand U5232 (N_5232,N_4683,N_4998);
or U5233 (N_5233,N_4564,N_4915);
nor U5234 (N_5234,N_4696,N_4585);
nor U5235 (N_5235,N_4902,N_4896);
and U5236 (N_5236,N_4534,N_4705);
and U5237 (N_5237,N_4949,N_4771);
xor U5238 (N_5238,N_4854,N_4741);
or U5239 (N_5239,N_4932,N_4895);
nand U5240 (N_5240,N_4550,N_4762);
xor U5241 (N_5241,N_4608,N_4933);
nor U5242 (N_5242,N_4859,N_4865);
or U5243 (N_5243,N_4540,N_4717);
nor U5244 (N_5244,N_4518,N_4734);
or U5245 (N_5245,N_4947,N_4679);
nand U5246 (N_5246,N_4597,N_4759);
and U5247 (N_5247,N_4940,N_4975);
and U5248 (N_5248,N_4974,N_4804);
and U5249 (N_5249,N_4779,N_4921);
or U5250 (N_5250,N_4739,N_4523);
xnor U5251 (N_5251,N_4926,N_4587);
and U5252 (N_5252,N_4999,N_4982);
or U5253 (N_5253,N_4503,N_4700);
nand U5254 (N_5254,N_4505,N_4895);
or U5255 (N_5255,N_4527,N_4512);
nor U5256 (N_5256,N_4967,N_4688);
or U5257 (N_5257,N_4987,N_4866);
nor U5258 (N_5258,N_4527,N_4638);
nor U5259 (N_5259,N_4889,N_4700);
nor U5260 (N_5260,N_4655,N_4979);
xor U5261 (N_5261,N_4837,N_4644);
xnor U5262 (N_5262,N_4544,N_4612);
nand U5263 (N_5263,N_4877,N_4793);
and U5264 (N_5264,N_4752,N_4662);
nand U5265 (N_5265,N_4907,N_4855);
nand U5266 (N_5266,N_4715,N_4594);
nand U5267 (N_5267,N_4739,N_4841);
and U5268 (N_5268,N_4766,N_4713);
nor U5269 (N_5269,N_4658,N_4753);
xor U5270 (N_5270,N_4748,N_4997);
or U5271 (N_5271,N_4879,N_4650);
and U5272 (N_5272,N_4826,N_4834);
and U5273 (N_5273,N_4989,N_4697);
nand U5274 (N_5274,N_4732,N_4894);
or U5275 (N_5275,N_4920,N_4559);
and U5276 (N_5276,N_4982,N_4580);
and U5277 (N_5277,N_4909,N_4636);
and U5278 (N_5278,N_4886,N_4981);
nand U5279 (N_5279,N_4652,N_4960);
nand U5280 (N_5280,N_4507,N_4917);
xnor U5281 (N_5281,N_4572,N_4708);
or U5282 (N_5282,N_4818,N_4611);
or U5283 (N_5283,N_4722,N_4723);
and U5284 (N_5284,N_4796,N_4500);
or U5285 (N_5285,N_4724,N_4795);
and U5286 (N_5286,N_4762,N_4613);
nand U5287 (N_5287,N_4772,N_4761);
nand U5288 (N_5288,N_4951,N_4934);
xor U5289 (N_5289,N_4822,N_4765);
or U5290 (N_5290,N_4730,N_4925);
and U5291 (N_5291,N_4858,N_4738);
xnor U5292 (N_5292,N_4980,N_4594);
xor U5293 (N_5293,N_4844,N_4599);
and U5294 (N_5294,N_4724,N_4805);
or U5295 (N_5295,N_4600,N_4725);
nand U5296 (N_5296,N_4730,N_4514);
and U5297 (N_5297,N_4832,N_4727);
xor U5298 (N_5298,N_4533,N_4984);
xor U5299 (N_5299,N_4977,N_4817);
or U5300 (N_5300,N_4672,N_4898);
or U5301 (N_5301,N_4631,N_4707);
nor U5302 (N_5302,N_4894,N_4524);
nor U5303 (N_5303,N_4967,N_4710);
and U5304 (N_5304,N_4855,N_4619);
nand U5305 (N_5305,N_4682,N_4956);
and U5306 (N_5306,N_4605,N_4709);
xnor U5307 (N_5307,N_4772,N_4817);
and U5308 (N_5308,N_4820,N_4853);
nor U5309 (N_5309,N_4595,N_4628);
or U5310 (N_5310,N_4627,N_4799);
xnor U5311 (N_5311,N_4806,N_4679);
and U5312 (N_5312,N_4977,N_4594);
or U5313 (N_5313,N_4574,N_4545);
xor U5314 (N_5314,N_4765,N_4914);
or U5315 (N_5315,N_4738,N_4546);
nor U5316 (N_5316,N_4786,N_4666);
nor U5317 (N_5317,N_4765,N_4862);
nor U5318 (N_5318,N_4801,N_4589);
nand U5319 (N_5319,N_4822,N_4563);
xnor U5320 (N_5320,N_4649,N_4956);
nor U5321 (N_5321,N_4652,N_4882);
and U5322 (N_5322,N_4831,N_4802);
nand U5323 (N_5323,N_4645,N_4970);
or U5324 (N_5324,N_4713,N_4562);
nand U5325 (N_5325,N_4579,N_4866);
nor U5326 (N_5326,N_4552,N_4843);
nor U5327 (N_5327,N_4966,N_4880);
nor U5328 (N_5328,N_4846,N_4661);
nor U5329 (N_5329,N_4691,N_4816);
nand U5330 (N_5330,N_4791,N_4530);
and U5331 (N_5331,N_4804,N_4988);
nor U5332 (N_5332,N_4603,N_4967);
nor U5333 (N_5333,N_4793,N_4668);
and U5334 (N_5334,N_4568,N_4778);
and U5335 (N_5335,N_4648,N_4799);
nor U5336 (N_5336,N_4866,N_4620);
or U5337 (N_5337,N_4732,N_4974);
and U5338 (N_5338,N_4934,N_4567);
nand U5339 (N_5339,N_4672,N_4960);
nand U5340 (N_5340,N_4910,N_4674);
and U5341 (N_5341,N_4948,N_4855);
or U5342 (N_5342,N_4596,N_4614);
nor U5343 (N_5343,N_4925,N_4598);
or U5344 (N_5344,N_4894,N_4756);
nand U5345 (N_5345,N_4547,N_4585);
nor U5346 (N_5346,N_4722,N_4670);
nor U5347 (N_5347,N_4550,N_4699);
and U5348 (N_5348,N_4619,N_4891);
xnor U5349 (N_5349,N_4902,N_4965);
nand U5350 (N_5350,N_4889,N_4808);
xnor U5351 (N_5351,N_4938,N_4775);
xnor U5352 (N_5352,N_4855,N_4786);
or U5353 (N_5353,N_4613,N_4976);
nor U5354 (N_5354,N_4903,N_4633);
nand U5355 (N_5355,N_4954,N_4797);
xnor U5356 (N_5356,N_4652,N_4712);
nor U5357 (N_5357,N_4765,N_4582);
xor U5358 (N_5358,N_4924,N_4790);
xor U5359 (N_5359,N_4701,N_4973);
xor U5360 (N_5360,N_4529,N_4511);
nor U5361 (N_5361,N_4572,N_4743);
nand U5362 (N_5362,N_4924,N_4892);
or U5363 (N_5363,N_4619,N_4515);
xor U5364 (N_5364,N_4703,N_4967);
and U5365 (N_5365,N_4905,N_4719);
and U5366 (N_5366,N_4698,N_4504);
and U5367 (N_5367,N_4750,N_4685);
or U5368 (N_5368,N_4942,N_4848);
xor U5369 (N_5369,N_4897,N_4572);
nand U5370 (N_5370,N_4688,N_4817);
xnor U5371 (N_5371,N_4870,N_4664);
nand U5372 (N_5372,N_4949,N_4508);
xnor U5373 (N_5373,N_4871,N_4828);
xor U5374 (N_5374,N_4754,N_4727);
nand U5375 (N_5375,N_4873,N_4979);
xnor U5376 (N_5376,N_4693,N_4522);
nor U5377 (N_5377,N_4662,N_4950);
and U5378 (N_5378,N_4937,N_4653);
nand U5379 (N_5379,N_4762,N_4527);
or U5380 (N_5380,N_4845,N_4675);
nor U5381 (N_5381,N_4575,N_4775);
nor U5382 (N_5382,N_4863,N_4984);
nand U5383 (N_5383,N_4809,N_4951);
or U5384 (N_5384,N_4982,N_4666);
nand U5385 (N_5385,N_4596,N_4510);
and U5386 (N_5386,N_4799,N_4864);
nand U5387 (N_5387,N_4501,N_4914);
nor U5388 (N_5388,N_4621,N_4863);
xnor U5389 (N_5389,N_4887,N_4606);
and U5390 (N_5390,N_4701,N_4562);
nand U5391 (N_5391,N_4813,N_4885);
xor U5392 (N_5392,N_4958,N_4729);
nand U5393 (N_5393,N_4884,N_4945);
or U5394 (N_5394,N_4662,N_4820);
nand U5395 (N_5395,N_4835,N_4758);
or U5396 (N_5396,N_4765,N_4947);
or U5397 (N_5397,N_4937,N_4590);
or U5398 (N_5398,N_4991,N_4743);
and U5399 (N_5399,N_4898,N_4827);
nor U5400 (N_5400,N_4869,N_4529);
nor U5401 (N_5401,N_4979,N_4936);
xor U5402 (N_5402,N_4725,N_4741);
nor U5403 (N_5403,N_4631,N_4581);
nand U5404 (N_5404,N_4535,N_4642);
nand U5405 (N_5405,N_4947,N_4674);
and U5406 (N_5406,N_4501,N_4742);
or U5407 (N_5407,N_4764,N_4685);
and U5408 (N_5408,N_4964,N_4789);
nor U5409 (N_5409,N_4682,N_4953);
and U5410 (N_5410,N_4766,N_4712);
and U5411 (N_5411,N_4938,N_4650);
nand U5412 (N_5412,N_4506,N_4782);
and U5413 (N_5413,N_4945,N_4810);
nor U5414 (N_5414,N_4773,N_4827);
xor U5415 (N_5415,N_4535,N_4657);
or U5416 (N_5416,N_4543,N_4668);
xnor U5417 (N_5417,N_4929,N_4730);
xnor U5418 (N_5418,N_4640,N_4596);
nor U5419 (N_5419,N_4703,N_4898);
nand U5420 (N_5420,N_4505,N_4707);
xnor U5421 (N_5421,N_4818,N_4942);
xor U5422 (N_5422,N_4808,N_4840);
xor U5423 (N_5423,N_4769,N_4734);
xor U5424 (N_5424,N_4693,N_4739);
nand U5425 (N_5425,N_4923,N_4996);
nand U5426 (N_5426,N_4797,N_4728);
and U5427 (N_5427,N_4651,N_4956);
and U5428 (N_5428,N_4726,N_4820);
xnor U5429 (N_5429,N_4754,N_4614);
or U5430 (N_5430,N_4974,N_4536);
or U5431 (N_5431,N_4878,N_4564);
or U5432 (N_5432,N_4722,N_4761);
nor U5433 (N_5433,N_4539,N_4581);
nand U5434 (N_5434,N_4647,N_4853);
nor U5435 (N_5435,N_4906,N_4511);
nor U5436 (N_5436,N_4799,N_4730);
and U5437 (N_5437,N_4693,N_4628);
and U5438 (N_5438,N_4501,N_4677);
and U5439 (N_5439,N_4645,N_4938);
nor U5440 (N_5440,N_4818,N_4575);
and U5441 (N_5441,N_4822,N_4725);
and U5442 (N_5442,N_4577,N_4698);
and U5443 (N_5443,N_4697,N_4634);
nor U5444 (N_5444,N_4627,N_4647);
nand U5445 (N_5445,N_4555,N_4890);
nor U5446 (N_5446,N_4522,N_4949);
nand U5447 (N_5447,N_4930,N_4650);
xor U5448 (N_5448,N_4977,N_4936);
or U5449 (N_5449,N_4598,N_4549);
or U5450 (N_5450,N_4617,N_4896);
or U5451 (N_5451,N_4914,N_4597);
and U5452 (N_5452,N_4531,N_4942);
nand U5453 (N_5453,N_4616,N_4633);
and U5454 (N_5454,N_4651,N_4857);
and U5455 (N_5455,N_4727,N_4523);
and U5456 (N_5456,N_4976,N_4616);
xor U5457 (N_5457,N_4688,N_4649);
nand U5458 (N_5458,N_4853,N_4904);
or U5459 (N_5459,N_4999,N_4718);
or U5460 (N_5460,N_4714,N_4883);
nand U5461 (N_5461,N_4500,N_4994);
nand U5462 (N_5462,N_4842,N_4836);
or U5463 (N_5463,N_4502,N_4735);
or U5464 (N_5464,N_4600,N_4731);
xnor U5465 (N_5465,N_4687,N_4641);
xnor U5466 (N_5466,N_4916,N_4931);
and U5467 (N_5467,N_4771,N_4921);
or U5468 (N_5468,N_4761,N_4852);
and U5469 (N_5469,N_4875,N_4828);
nand U5470 (N_5470,N_4714,N_4678);
or U5471 (N_5471,N_4503,N_4763);
and U5472 (N_5472,N_4795,N_4683);
nand U5473 (N_5473,N_4960,N_4635);
nand U5474 (N_5474,N_4816,N_4536);
nand U5475 (N_5475,N_4683,N_4657);
or U5476 (N_5476,N_4556,N_4793);
xor U5477 (N_5477,N_4996,N_4793);
nand U5478 (N_5478,N_4992,N_4521);
or U5479 (N_5479,N_4596,N_4661);
xor U5480 (N_5480,N_4558,N_4516);
and U5481 (N_5481,N_4971,N_4688);
nor U5482 (N_5482,N_4793,N_4585);
nor U5483 (N_5483,N_4714,N_4615);
and U5484 (N_5484,N_4849,N_4916);
or U5485 (N_5485,N_4858,N_4811);
nor U5486 (N_5486,N_4799,N_4698);
xnor U5487 (N_5487,N_4797,N_4935);
xor U5488 (N_5488,N_4942,N_4815);
and U5489 (N_5489,N_4993,N_4630);
and U5490 (N_5490,N_4741,N_4967);
or U5491 (N_5491,N_4763,N_4891);
or U5492 (N_5492,N_4603,N_4507);
xor U5493 (N_5493,N_4763,N_4655);
or U5494 (N_5494,N_4996,N_4886);
xor U5495 (N_5495,N_4514,N_4571);
or U5496 (N_5496,N_4573,N_4712);
nand U5497 (N_5497,N_4578,N_4922);
nor U5498 (N_5498,N_4577,N_4854);
or U5499 (N_5499,N_4808,N_4914);
xor U5500 (N_5500,N_5007,N_5278);
nand U5501 (N_5501,N_5009,N_5282);
xnor U5502 (N_5502,N_5416,N_5075);
xnor U5503 (N_5503,N_5292,N_5385);
xnor U5504 (N_5504,N_5195,N_5076);
xor U5505 (N_5505,N_5456,N_5143);
or U5506 (N_5506,N_5373,N_5375);
nor U5507 (N_5507,N_5438,N_5115);
xnor U5508 (N_5508,N_5365,N_5372);
nor U5509 (N_5509,N_5175,N_5166);
xnor U5510 (N_5510,N_5199,N_5204);
nand U5511 (N_5511,N_5295,N_5410);
or U5512 (N_5512,N_5350,N_5257);
xnor U5513 (N_5513,N_5086,N_5064);
and U5514 (N_5514,N_5008,N_5481);
xnor U5515 (N_5515,N_5269,N_5145);
or U5516 (N_5516,N_5432,N_5404);
xor U5517 (N_5517,N_5367,N_5260);
nor U5518 (N_5518,N_5408,N_5276);
or U5519 (N_5519,N_5376,N_5133);
or U5520 (N_5520,N_5490,N_5047);
nor U5521 (N_5521,N_5489,N_5381);
nor U5522 (N_5522,N_5400,N_5138);
or U5523 (N_5523,N_5283,N_5461);
nor U5524 (N_5524,N_5111,N_5296);
nand U5525 (N_5525,N_5083,N_5221);
nor U5526 (N_5526,N_5171,N_5273);
and U5527 (N_5527,N_5429,N_5208);
nor U5528 (N_5528,N_5346,N_5314);
nor U5529 (N_5529,N_5493,N_5156);
nand U5530 (N_5530,N_5174,N_5485);
and U5531 (N_5531,N_5182,N_5453);
nand U5532 (N_5532,N_5227,N_5303);
or U5533 (N_5533,N_5205,N_5442);
and U5534 (N_5534,N_5207,N_5304);
nand U5535 (N_5535,N_5417,N_5452);
or U5536 (N_5536,N_5117,N_5271);
nand U5537 (N_5537,N_5266,N_5394);
xor U5538 (N_5538,N_5251,N_5230);
and U5539 (N_5539,N_5027,N_5019);
and U5540 (N_5540,N_5063,N_5164);
or U5541 (N_5541,N_5446,N_5341);
nand U5542 (N_5542,N_5335,N_5060);
or U5543 (N_5543,N_5413,N_5362);
nor U5544 (N_5544,N_5078,N_5387);
and U5545 (N_5545,N_5479,N_5109);
nor U5546 (N_5546,N_5026,N_5356);
xor U5547 (N_5547,N_5361,N_5358);
and U5548 (N_5548,N_5157,N_5401);
nand U5549 (N_5549,N_5349,N_5337);
nand U5550 (N_5550,N_5041,N_5325);
or U5551 (N_5551,N_5353,N_5149);
or U5552 (N_5552,N_5286,N_5105);
nand U5553 (N_5553,N_5395,N_5242);
xnor U5554 (N_5554,N_5137,N_5403);
or U5555 (N_5555,N_5354,N_5077);
xor U5556 (N_5556,N_5448,N_5229);
or U5557 (N_5557,N_5308,N_5285);
nand U5558 (N_5558,N_5213,N_5294);
xor U5559 (N_5559,N_5056,N_5470);
nor U5560 (N_5560,N_5445,N_5084);
or U5561 (N_5561,N_5345,N_5342);
nor U5562 (N_5562,N_5409,N_5024);
or U5563 (N_5563,N_5412,N_5360);
nor U5564 (N_5564,N_5068,N_5211);
nor U5565 (N_5565,N_5033,N_5431);
and U5566 (N_5566,N_5352,N_5180);
nand U5567 (N_5567,N_5324,N_5085);
nand U5568 (N_5568,N_5263,N_5100);
nand U5569 (N_5569,N_5032,N_5359);
and U5570 (N_5570,N_5106,N_5396);
nor U5571 (N_5571,N_5465,N_5318);
or U5572 (N_5572,N_5167,N_5457);
xor U5573 (N_5573,N_5038,N_5247);
and U5574 (N_5574,N_5284,N_5113);
nor U5575 (N_5575,N_5173,N_5151);
and U5576 (N_5576,N_5232,N_5190);
or U5577 (N_5577,N_5206,N_5114);
nand U5578 (N_5578,N_5148,N_5194);
nor U5579 (N_5579,N_5018,N_5246);
and U5580 (N_5580,N_5252,N_5101);
nand U5581 (N_5581,N_5329,N_5338);
nand U5582 (N_5582,N_5398,N_5241);
nand U5583 (N_5583,N_5159,N_5476);
nand U5584 (N_5584,N_5236,N_5288);
nand U5585 (N_5585,N_5186,N_5326);
and U5586 (N_5586,N_5333,N_5424);
nor U5587 (N_5587,N_5193,N_5460);
and U5588 (N_5588,N_5467,N_5189);
nor U5589 (N_5589,N_5067,N_5176);
or U5590 (N_5590,N_5293,N_5081);
nand U5591 (N_5591,N_5274,N_5022);
or U5592 (N_5592,N_5094,N_5216);
and U5593 (N_5593,N_5209,N_5127);
or U5594 (N_5594,N_5317,N_5418);
or U5595 (N_5595,N_5297,N_5158);
nor U5596 (N_5596,N_5444,N_5474);
nand U5597 (N_5597,N_5357,N_5455);
or U5598 (N_5598,N_5374,N_5217);
or U5599 (N_5599,N_5089,N_5484);
nand U5600 (N_5600,N_5421,N_5343);
nor U5601 (N_5601,N_5128,N_5051);
nand U5602 (N_5602,N_5002,N_5183);
or U5603 (N_5603,N_5497,N_5015);
nand U5604 (N_5604,N_5091,N_5003);
nand U5605 (N_5605,N_5146,N_5370);
or U5606 (N_5606,N_5298,N_5426);
nand U5607 (N_5607,N_5264,N_5184);
xor U5608 (N_5608,N_5116,N_5050);
xnor U5609 (N_5609,N_5131,N_5427);
or U5610 (N_5610,N_5316,N_5073);
or U5611 (N_5611,N_5380,N_5055);
and U5612 (N_5612,N_5407,N_5331);
nand U5613 (N_5613,N_5382,N_5119);
nor U5614 (N_5614,N_5126,N_5220);
nor U5615 (N_5615,N_5201,N_5347);
nor U5616 (N_5616,N_5090,N_5098);
nand U5617 (N_5617,N_5035,N_5388);
nand U5618 (N_5618,N_5440,N_5203);
nor U5619 (N_5619,N_5322,N_5499);
nor U5620 (N_5620,N_5462,N_5144);
nand U5621 (N_5621,N_5238,N_5016);
nor U5622 (N_5622,N_5178,N_5468);
nand U5623 (N_5623,N_5177,N_5226);
nor U5624 (N_5624,N_5052,N_5475);
and U5625 (N_5625,N_5267,N_5492);
xnor U5626 (N_5626,N_5219,N_5480);
nand U5627 (N_5627,N_5256,N_5486);
nor U5628 (N_5628,N_5306,N_5253);
xor U5629 (N_5629,N_5430,N_5021);
nand U5630 (N_5630,N_5348,N_5366);
and U5631 (N_5631,N_5469,N_5488);
and U5632 (N_5632,N_5363,N_5272);
xor U5633 (N_5633,N_5312,N_5034);
nor U5634 (N_5634,N_5428,N_5170);
xor U5635 (N_5635,N_5287,N_5054);
and U5636 (N_5636,N_5118,N_5040);
xnor U5637 (N_5637,N_5001,N_5415);
xor U5638 (N_5638,N_5384,N_5327);
nand U5639 (N_5639,N_5344,N_5458);
nand U5640 (N_5640,N_5437,N_5202);
xnor U5641 (N_5641,N_5301,N_5074);
xnor U5642 (N_5642,N_5134,N_5152);
and U5643 (N_5643,N_5459,N_5218);
xnor U5644 (N_5644,N_5025,N_5196);
or U5645 (N_5645,N_5210,N_5061);
nand U5646 (N_5646,N_5255,N_5120);
and U5647 (N_5647,N_5478,N_5393);
nand U5648 (N_5648,N_5261,N_5187);
and U5649 (N_5649,N_5447,N_5332);
xor U5650 (N_5650,N_5179,N_5140);
nand U5651 (N_5651,N_5291,N_5240);
nor U5652 (N_5652,N_5065,N_5223);
or U5653 (N_5653,N_5435,N_5069);
nor U5654 (N_5654,N_5192,N_5270);
nor U5655 (N_5655,N_5235,N_5147);
or U5656 (N_5656,N_5425,N_5124);
or U5657 (N_5657,N_5249,N_5058);
nand U5658 (N_5658,N_5099,N_5150);
nor U5659 (N_5659,N_5129,N_5231);
or U5660 (N_5660,N_5030,N_5154);
xor U5661 (N_5661,N_5057,N_5355);
nor U5662 (N_5662,N_5351,N_5414);
nand U5663 (N_5663,N_5494,N_5244);
nor U5664 (N_5664,N_5095,N_5419);
and U5665 (N_5665,N_5368,N_5228);
nor U5666 (N_5666,N_5265,N_5454);
or U5667 (N_5667,N_5305,N_5315);
and U5668 (N_5668,N_5302,N_5200);
xnor U5669 (N_5669,N_5036,N_5121);
xnor U5670 (N_5670,N_5390,N_5142);
and U5671 (N_5671,N_5254,N_5004);
nand U5672 (N_5672,N_5181,N_5496);
nor U5673 (N_5673,N_5321,N_5371);
or U5674 (N_5674,N_5049,N_5017);
nor U5675 (N_5675,N_5377,N_5320);
and U5676 (N_5676,N_5433,N_5013);
or U5677 (N_5677,N_5139,N_5299);
xnor U5678 (N_5678,N_5309,N_5020);
and U5679 (N_5679,N_5014,N_5102);
xnor U5680 (N_5680,N_5482,N_5044);
and U5681 (N_5681,N_5406,N_5443);
nand U5682 (N_5682,N_5328,N_5439);
nor U5683 (N_5683,N_5012,N_5191);
nor U5684 (N_5684,N_5062,N_5104);
nand U5685 (N_5685,N_5125,N_5498);
xnor U5686 (N_5686,N_5402,N_5392);
nand U5687 (N_5687,N_5472,N_5248);
nand U5688 (N_5688,N_5262,N_5123);
or U5689 (N_5689,N_5028,N_5122);
nand U5690 (N_5690,N_5188,N_5330);
nor U5691 (N_5691,N_5340,N_5059);
nand U5692 (N_5692,N_5023,N_5399);
nand U5693 (N_5693,N_5289,N_5378);
and U5694 (N_5694,N_5082,N_5163);
nand U5695 (N_5695,N_5389,N_5072);
and U5696 (N_5696,N_5491,N_5092);
nand U5697 (N_5697,N_5165,N_5155);
xnor U5698 (N_5698,N_5185,N_5239);
and U5699 (N_5699,N_5112,N_5212);
xor U5700 (N_5700,N_5088,N_5011);
xor U5701 (N_5701,N_5245,N_5096);
xnor U5702 (N_5702,N_5483,N_5471);
nor U5703 (N_5703,N_5463,N_5334);
xnor U5704 (N_5704,N_5449,N_5369);
and U5705 (N_5705,N_5258,N_5215);
and U5706 (N_5706,N_5168,N_5070);
xnor U5707 (N_5707,N_5495,N_5048);
xnor U5708 (N_5708,N_5053,N_5243);
xnor U5709 (N_5709,N_5422,N_5161);
or U5710 (N_5710,N_5259,N_5300);
and U5711 (N_5711,N_5319,N_5110);
xor U5712 (N_5712,N_5234,N_5135);
nand U5713 (N_5713,N_5141,N_5275);
or U5714 (N_5714,N_5268,N_5093);
xor U5715 (N_5715,N_5046,N_5136);
and U5716 (N_5716,N_5420,N_5280);
nand U5717 (N_5717,N_5169,N_5441);
and U5718 (N_5718,N_5310,N_5097);
or U5719 (N_5719,N_5473,N_5225);
and U5720 (N_5720,N_5397,N_5277);
and U5721 (N_5721,N_5079,N_5411);
nor U5722 (N_5722,N_5162,N_5364);
xnor U5723 (N_5723,N_5279,N_5237);
xor U5724 (N_5724,N_5451,N_5042);
or U5725 (N_5725,N_5031,N_5383);
or U5726 (N_5726,N_5233,N_5045);
and U5727 (N_5727,N_5039,N_5250);
and U5728 (N_5728,N_5379,N_5290);
xnor U5729 (N_5729,N_5160,N_5005);
xnor U5730 (N_5730,N_5103,N_5172);
nand U5731 (N_5731,N_5006,N_5222);
nor U5732 (N_5732,N_5307,N_5386);
and U5733 (N_5733,N_5029,N_5130);
xor U5734 (N_5734,N_5434,N_5339);
and U5735 (N_5735,N_5197,N_5311);
and U5736 (N_5736,N_5477,N_5336);
nor U5737 (N_5737,N_5108,N_5000);
or U5738 (N_5738,N_5037,N_5132);
xor U5739 (N_5739,N_5405,N_5323);
nand U5740 (N_5740,N_5080,N_5313);
nand U5741 (N_5741,N_5487,N_5071);
nand U5742 (N_5742,N_5436,N_5464);
nor U5743 (N_5743,N_5087,N_5107);
and U5744 (N_5744,N_5423,N_5391);
or U5745 (N_5745,N_5281,N_5010);
nor U5746 (N_5746,N_5066,N_5043);
xor U5747 (N_5747,N_5153,N_5224);
or U5748 (N_5748,N_5214,N_5466);
nor U5749 (N_5749,N_5450,N_5198);
xor U5750 (N_5750,N_5244,N_5261);
nand U5751 (N_5751,N_5138,N_5237);
xor U5752 (N_5752,N_5370,N_5098);
xnor U5753 (N_5753,N_5149,N_5456);
and U5754 (N_5754,N_5312,N_5308);
or U5755 (N_5755,N_5048,N_5168);
xnor U5756 (N_5756,N_5278,N_5444);
or U5757 (N_5757,N_5408,N_5092);
nand U5758 (N_5758,N_5442,N_5366);
xor U5759 (N_5759,N_5087,N_5489);
nor U5760 (N_5760,N_5320,N_5034);
nand U5761 (N_5761,N_5108,N_5103);
and U5762 (N_5762,N_5279,N_5227);
or U5763 (N_5763,N_5272,N_5089);
nor U5764 (N_5764,N_5187,N_5203);
nor U5765 (N_5765,N_5321,N_5315);
nor U5766 (N_5766,N_5300,N_5446);
xor U5767 (N_5767,N_5286,N_5352);
xor U5768 (N_5768,N_5436,N_5420);
nand U5769 (N_5769,N_5199,N_5059);
nand U5770 (N_5770,N_5306,N_5135);
and U5771 (N_5771,N_5259,N_5264);
and U5772 (N_5772,N_5365,N_5109);
nand U5773 (N_5773,N_5491,N_5471);
and U5774 (N_5774,N_5015,N_5171);
nor U5775 (N_5775,N_5416,N_5184);
nor U5776 (N_5776,N_5046,N_5234);
or U5777 (N_5777,N_5087,N_5452);
xor U5778 (N_5778,N_5269,N_5226);
nor U5779 (N_5779,N_5141,N_5446);
and U5780 (N_5780,N_5185,N_5248);
nand U5781 (N_5781,N_5279,N_5289);
xnor U5782 (N_5782,N_5375,N_5259);
nor U5783 (N_5783,N_5326,N_5040);
or U5784 (N_5784,N_5388,N_5453);
xor U5785 (N_5785,N_5082,N_5360);
or U5786 (N_5786,N_5031,N_5203);
nand U5787 (N_5787,N_5292,N_5240);
nor U5788 (N_5788,N_5007,N_5450);
nor U5789 (N_5789,N_5153,N_5174);
xor U5790 (N_5790,N_5469,N_5169);
and U5791 (N_5791,N_5150,N_5247);
xor U5792 (N_5792,N_5211,N_5166);
or U5793 (N_5793,N_5277,N_5472);
nor U5794 (N_5794,N_5056,N_5223);
nor U5795 (N_5795,N_5096,N_5445);
or U5796 (N_5796,N_5370,N_5439);
or U5797 (N_5797,N_5225,N_5156);
nand U5798 (N_5798,N_5481,N_5421);
nand U5799 (N_5799,N_5306,N_5183);
xnor U5800 (N_5800,N_5120,N_5140);
nand U5801 (N_5801,N_5219,N_5302);
and U5802 (N_5802,N_5058,N_5350);
and U5803 (N_5803,N_5093,N_5236);
or U5804 (N_5804,N_5423,N_5233);
or U5805 (N_5805,N_5006,N_5286);
and U5806 (N_5806,N_5459,N_5022);
and U5807 (N_5807,N_5482,N_5116);
and U5808 (N_5808,N_5436,N_5015);
nor U5809 (N_5809,N_5335,N_5078);
nor U5810 (N_5810,N_5068,N_5017);
xor U5811 (N_5811,N_5431,N_5436);
and U5812 (N_5812,N_5172,N_5453);
xnor U5813 (N_5813,N_5352,N_5372);
nand U5814 (N_5814,N_5453,N_5474);
nor U5815 (N_5815,N_5147,N_5153);
and U5816 (N_5816,N_5079,N_5429);
nor U5817 (N_5817,N_5010,N_5412);
or U5818 (N_5818,N_5491,N_5338);
and U5819 (N_5819,N_5142,N_5213);
nand U5820 (N_5820,N_5099,N_5196);
xnor U5821 (N_5821,N_5278,N_5366);
nand U5822 (N_5822,N_5218,N_5222);
and U5823 (N_5823,N_5091,N_5426);
nor U5824 (N_5824,N_5164,N_5085);
or U5825 (N_5825,N_5329,N_5293);
nor U5826 (N_5826,N_5098,N_5101);
and U5827 (N_5827,N_5015,N_5026);
xor U5828 (N_5828,N_5171,N_5014);
nand U5829 (N_5829,N_5285,N_5230);
and U5830 (N_5830,N_5231,N_5439);
nand U5831 (N_5831,N_5176,N_5273);
nor U5832 (N_5832,N_5339,N_5042);
and U5833 (N_5833,N_5220,N_5038);
nor U5834 (N_5834,N_5077,N_5346);
xor U5835 (N_5835,N_5138,N_5337);
nand U5836 (N_5836,N_5159,N_5490);
nor U5837 (N_5837,N_5310,N_5433);
nand U5838 (N_5838,N_5003,N_5046);
nand U5839 (N_5839,N_5483,N_5229);
or U5840 (N_5840,N_5107,N_5147);
nand U5841 (N_5841,N_5395,N_5398);
xor U5842 (N_5842,N_5144,N_5120);
nor U5843 (N_5843,N_5058,N_5065);
or U5844 (N_5844,N_5104,N_5137);
nor U5845 (N_5845,N_5445,N_5063);
nand U5846 (N_5846,N_5293,N_5020);
xor U5847 (N_5847,N_5275,N_5386);
and U5848 (N_5848,N_5202,N_5146);
or U5849 (N_5849,N_5291,N_5395);
nand U5850 (N_5850,N_5306,N_5422);
nand U5851 (N_5851,N_5079,N_5032);
xnor U5852 (N_5852,N_5424,N_5259);
and U5853 (N_5853,N_5474,N_5245);
nand U5854 (N_5854,N_5084,N_5166);
nand U5855 (N_5855,N_5245,N_5333);
xnor U5856 (N_5856,N_5486,N_5496);
nor U5857 (N_5857,N_5256,N_5115);
xnor U5858 (N_5858,N_5142,N_5299);
nor U5859 (N_5859,N_5106,N_5424);
nand U5860 (N_5860,N_5275,N_5447);
nand U5861 (N_5861,N_5363,N_5226);
or U5862 (N_5862,N_5458,N_5010);
and U5863 (N_5863,N_5147,N_5117);
or U5864 (N_5864,N_5222,N_5330);
xor U5865 (N_5865,N_5401,N_5281);
xor U5866 (N_5866,N_5092,N_5126);
nand U5867 (N_5867,N_5190,N_5150);
nand U5868 (N_5868,N_5074,N_5026);
nor U5869 (N_5869,N_5215,N_5358);
or U5870 (N_5870,N_5067,N_5220);
nand U5871 (N_5871,N_5104,N_5480);
xnor U5872 (N_5872,N_5092,N_5467);
xnor U5873 (N_5873,N_5366,N_5064);
or U5874 (N_5874,N_5391,N_5380);
and U5875 (N_5875,N_5480,N_5085);
and U5876 (N_5876,N_5081,N_5278);
nor U5877 (N_5877,N_5074,N_5212);
or U5878 (N_5878,N_5115,N_5061);
nand U5879 (N_5879,N_5334,N_5093);
or U5880 (N_5880,N_5184,N_5291);
and U5881 (N_5881,N_5419,N_5052);
nand U5882 (N_5882,N_5481,N_5385);
or U5883 (N_5883,N_5132,N_5489);
and U5884 (N_5884,N_5247,N_5393);
and U5885 (N_5885,N_5318,N_5445);
nand U5886 (N_5886,N_5223,N_5399);
or U5887 (N_5887,N_5152,N_5000);
nor U5888 (N_5888,N_5118,N_5031);
or U5889 (N_5889,N_5151,N_5274);
nand U5890 (N_5890,N_5358,N_5446);
or U5891 (N_5891,N_5251,N_5056);
nor U5892 (N_5892,N_5497,N_5244);
and U5893 (N_5893,N_5086,N_5053);
and U5894 (N_5894,N_5247,N_5321);
xnor U5895 (N_5895,N_5330,N_5245);
and U5896 (N_5896,N_5082,N_5246);
or U5897 (N_5897,N_5414,N_5407);
nand U5898 (N_5898,N_5348,N_5193);
nor U5899 (N_5899,N_5234,N_5189);
or U5900 (N_5900,N_5097,N_5391);
and U5901 (N_5901,N_5098,N_5004);
nand U5902 (N_5902,N_5360,N_5329);
xor U5903 (N_5903,N_5212,N_5280);
and U5904 (N_5904,N_5269,N_5072);
and U5905 (N_5905,N_5262,N_5126);
and U5906 (N_5906,N_5089,N_5259);
nand U5907 (N_5907,N_5304,N_5103);
or U5908 (N_5908,N_5222,N_5098);
nand U5909 (N_5909,N_5396,N_5158);
xor U5910 (N_5910,N_5156,N_5126);
nand U5911 (N_5911,N_5016,N_5360);
nand U5912 (N_5912,N_5144,N_5237);
and U5913 (N_5913,N_5233,N_5447);
nand U5914 (N_5914,N_5456,N_5260);
and U5915 (N_5915,N_5088,N_5276);
and U5916 (N_5916,N_5078,N_5161);
nor U5917 (N_5917,N_5451,N_5400);
and U5918 (N_5918,N_5441,N_5035);
xnor U5919 (N_5919,N_5466,N_5406);
or U5920 (N_5920,N_5338,N_5457);
xnor U5921 (N_5921,N_5274,N_5442);
or U5922 (N_5922,N_5176,N_5358);
nand U5923 (N_5923,N_5064,N_5311);
nor U5924 (N_5924,N_5204,N_5270);
and U5925 (N_5925,N_5090,N_5018);
or U5926 (N_5926,N_5268,N_5423);
or U5927 (N_5927,N_5084,N_5125);
nor U5928 (N_5928,N_5459,N_5401);
and U5929 (N_5929,N_5044,N_5499);
and U5930 (N_5930,N_5241,N_5305);
nand U5931 (N_5931,N_5000,N_5460);
nor U5932 (N_5932,N_5154,N_5489);
xnor U5933 (N_5933,N_5440,N_5381);
and U5934 (N_5934,N_5348,N_5085);
nor U5935 (N_5935,N_5089,N_5362);
nor U5936 (N_5936,N_5480,N_5467);
and U5937 (N_5937,N_5208,N_5182);
nor U5938 (N_5938,N_5223,N_5270);
and U5939 (N_5939,N_5248,N_5173);
or U5940 (N_5940,N_5103,N_5372);
xor U5941 (N_5941,N_5431,N_5188);
xnor U5942 (N_5942,N_5381,N_5217);
or U5943 (N_5943,N_5039,N_5034);
or U5944 (N_5944,N_5457,N_5034);
nor U5945 (N_5945,N_5230,N_5256);
and U5946 (N_5946,N_5377,N_5355);
nand U5947 (N_5947,N_5019,N_5048);
xnor U5948 (N_5948,N_5281,N_5329);
and U5949 (N_5949,N_5187,N_5370);
or U5950 (N_5950,N_5118,N_5261);
and U5951 (N_5951,N_5295,N_5070);
or U5952 (N_5952,N_5396,N_5174);
nor U5953 (N_5953,N_5158,N_5102);
nand U5954 (N_5954,N_5433,N_5358);
nand U5955 (N_5955,N_5285,N_5284);
nand U5956 (N_5956,N_5420,N_5411);
xnor U5957 (N_5957,N_5045,N_5133);
nor U5958 (N_5958,N_5142,N_5455);
nand U5959 (N_5959,N_5445,N_5050);
or U5960 (N_5960,N_5093,N_5442);
xnor U5961 (N_5961,N_5444,N_5283);
nand U5962 (N_5962,N_5054,N_5293);
nor U5963 (N_5963,N_5464,N_5331);
nand U5964 (N_5964,N_5190,N_5467);
nand U5965 (N_5965,N_5025,N_5490);
nor U5966 (N_5966,N_5230,N_5002);
xor U5967 (N_5967,N_5329,N_5242);
and U5968 (N_5968,N_5401,N_5320);
nor U5969 (N_5969,N_5447,N_5223);
or U5970 (N_5970,N_5012,N_5333);
and U5971 (N_5971,N_5267,N_5338);
nand U5972 (N_5972,N_5061,N_5139);
xor U5973 (N_5973,N_5435,N_5433);
nand U5974 (N_5974,N_5251,N_5284);
or U5975 (N_5975,N_5330,N_5383);
nand U5976 (N_5976,N_5469,N_5279);
nor U5977 (N_5977,N_5203,N_5144);
nor U5978 (N_5978,N_5369,N_5467);
and U5979 (N_5979,N_5260,N_5210);
xnor U5980 (N_5980,N_5319,N_5489);
xor U5981 (N_5981,N_5307,N_5005);
nor U5982 (N_5982,N_5066,N_5254);
nor U5983 (N_5983,N_5082,N_5499);
and U5984 (N_5984,N_5296,N_5042);
or U5985 (N_5985,N_5095,N_5319);
nor U5986 (N_5986,N_5326,N_5043);
nor U5987 (N_5987,N_5068,N_5148);
nor U5988 (N_5988,N_5360,N_5339);
or U5989 (N_5989,N_5331,N_5355);
nor U5990 (N_5990,N_5387,N_5195);
nor U5991 (N_5991,N_5399,N_5283);
xnor U5992 (N_5992,N_5037,N_5273);
or U5993 (N_5993,N_5331,N_5031);
and U5994 (N_5994,N_5405,N_5488);
nor U5995 (N_5995,N_5360,N_5321);
nor U5996 (N_5996,N_5149,N_5406);
or U5997 (N_5997,N_5060,N_5460);
nand U5998 (N_5998,N_5462,N_5092);
nor U5999 (N_5999,N_5258,N_5330);
nor U6000 (N_6000,N_5727,N_5511);
xor U6001 (N_6001,N_5904,N_5729);
and U6002 (N_6002,N_5857,N_5767);
and U6003 (N_6003,N_5896,N_5733);
xnor U6004 (N_6004,N_5960,N_5812);
nor U6005 (N_6005,N_5654,N_5668);
and U6006 (N_6006,N_5586,N_5585);
xor U6007 (N_6007,N_5545,N_5593);
nand U6008 (N_6008,N_5947,N_5870);
nor U6009 (N_6009,N_5787,N_5666);
xor U6010 (N_6010,N_5644,N_5778);
and U6011 (N_6011,N_5853,N_5661);
and U6012 (N_6012,N_5709,N_5656);
and U6013 (N_6013,N_5951,N_5541);
or U6014 (N_6014,N_5739,N_5935);
nand U6015 (N_6015,N_5682,N_5886);
xor U6016 (N_6016,N_5818,N_5859);
nor U6017 (N_6017,N_5613,N_5548);
nor U6018 (N_6018,N_5702,N_5711);
and U6019 (N_6019,N_5908,N_5755);
nand U6020 (N_6020,N_5544,N_5703);
nor U6021 (N_6021,N_5925,N_5742);
xor U6022 (N_6022,N_5941,N_5653);
and U6023 (N_6023,N_5581,N_5891);
or U6024 (N_6024,N_5512,N_5866);
xnor U6025 (N_6025,N_5754,N_5557);
and U6026 (N_6026,N_5928,N_5704);
and U6027 (N_6027,N_5991,N_5569);
or U6028 (N_6028,N_5751,N_5527);
xor U6029 (N_6029,N_5753,N_5670);
nand U6030 (N_6030,N_5747,N_5628);
nor U6031 (N_6031,N_5678,N_5636);
or U6032 (N_6032,N_5867,N_5529);
nand U6033 (N_6033,N_5697,N_5917);
xor U6034 (N_6034,N_5551,N_5877);
xor U6035 (N_6035,N_5599,N_5530);
and U6036 (N_6036,N_5770,N_5736);
or U6037 (N_6037,N_5642,N_5905);
nand U6038 (N_6038,N_5611,N_5845);
nand U6039 (N_6039,N_5696,N_5679);
nand U6040 (N_6040,N_5554,N_5712);
and U6041 (N_6041,N_5524,N_5836);
or U6042 (N_6042,N_5930,N_5556);
or U6043 (N_6043,N_5617,N_5777);
nand U6044 (N_6044,N_5620,N_5505);
or U6045 (N_6045,N_5789,N_5549);
nor U6046 (N_6046,N_5592,N_5992);
nand U6047 (N_6047,N_5810,N_5623);
or U6048 (N_6048,N_5912,N_5976);
xor U6049 (N_6049,N_5907,N_5748);
nand U6050 (N_6050,N_5906,N_5657);
and U6051 (N_6051,N_5920,N_5966);
xor U6052 (N_6052,N_5987,N_5562);
xor U6053 (N_6053,N_5664,N_5879);
xnor U6054 (N_6054,N_5771,N_5804);
or U6055 (N_6055,N_5680,N_5981);
and U6056 (N_6056,N_5815,N_5852);
and U6057 (N_6057,N_5690,N_5684);
nor U6058 (N_6058,N_5923,N_5990);
or U6059 (N_6059,N_5932,N_5843);
or U6060 (N_6060,N_5766,N_5889);
and U6061 (N_6061,N_5944,N_5788);
xnor U6062 (N_6062,N_5525,N_5571);
and U6063 (N_6063,N_5779,N_5612);
and U6064 (N_6064,N_5794,N_5553);
xor U6065 (N_6065,N_5868,N_5849);
nor U6066 (N_6066,N_5783,N_5775);
nor U6067 (N_6067,N_5560,N_5821);
or U6068 (N_6068,N_5954,N_5791);
and U6069 (N_6069,N_5792,N_5945);
xnor U6070 (N_6070,N_5894,N_5962);
nor U6071 (N_6071,N_5938,N_5558);
nand U6072 (N_6072,N_5692,N_5506);
xnor U6073 (N_6073,N_5567,N_5937);
nand U6074 (N_6074,N_5745,N_5909);
xnor U6075 (N_6075,N_5827,N_5740);
xor U6076 (N_6076,N_5765,N_5933);
and U6077 (N_6077,N_5974,N_5835);
xor U6078 (N_6078,N_5590,N_5832);
nor U6079 (N_6079,N_5959,N_5714);
and U6080 (N_6080,N_5598,N_5501);
xor U6081 (N_6081,N_5893,N_5784);
nand U6082 (N_6082,N_5880,N_5566);
nand U6083 (N_6083,N_5994,N_5662);
xnor U6084 (N_6084,N_5667,N_5830);
nor U6085 (N_6085,N_5717,N_5926);
nand U6086 (N_6086,N_5610,N_5689);
or U6087 (N_6087,N_5762,N_5584);
nor U6088 (N_6088,N_5624,N_5659);
nor U6089 (N_6089,N_5797,N_5722);
nor U6090 (N_6090,N_5802,N_5713);
xor U6091 (N_6091,N_5750,N_5902);
nor U6092 (N_6092,N_5848,N_5672);
nand U6093 (N_6093,N_5681,N_5977);
and U6094 (N_6094,N_5918,N_5693);
or U6095 (N_6095,N_5675,N_5741);
nand U6096 (N_6096,N_5734,N_5996);
nand U6097 (N_6097,N_5516,N_5911);
and U6098 (N_6098,N_5972,N_5686);
nand U6099 (N_6099,N_5842,N_5806);
or U6100 (N_6100,N_5931,N_5744);
or U6101 (N_6101,N_5943,N_5851);
or U6102 (N_6102,N_5723,N_5691);
nor U6103 (N_6103,N_5732,N_5519);
or U6104 (N_6104,N_5860,N_5887);
xnor U6105 (N_6105,N_5865,N_5898);
nand U6106 (N_6106,N_5942,N_5805);
and U6107 (N_6107,N_5616,N_5946);
xor U6108 (N_6108,N_5824,N_5786);
nand U6109 (N_6109,N_5963,N_5706);
or U6110 (N_6110,N_5601,N_5564);
nor U6111 (N_6111,N_5542,N_5629);
and U6112 (N_6112,N_5803,N_5638);
and U6113 (N_6113,N_5989,N_5757);
xnor U6114 (N_6114,N_5705,N_5983);
or U6115 (N_6115,N_5526,N_5885);
nor U6116 (N_6116,N_5998,N_5890);
nor U6117 (N_6117,N_5600,N_5673);
xnor U6118 (N_6118,N_5969,N_5635);
nand U6119 (N_6119,N_5967,N_5630);
nor U6120 (N_6120,N_5874,N_5546);
nand U6121 (N_6121,N_5700,N_5964);
nor U6122 (N_6122,N_5698,N_5708);
nand U6123 (N_6123,N_5694,N_5577);
or U6124 (N_6124,N_5688,N_5716);
and U6125 (N_6125,N_5536,N_5999);
nor U6126 (N_6126,N_5502,N_5822);
or U6127 (N_6127,N_5658,N_5719);
and U6128 (N_6128,N_5764,N_5854);
nor U6129 (N_6129,N_5521,N_5965);
nand U6130 (N_6130,N_5772,N_5720);
and U6131 (N_6131,N_5507,N_5948);
and U6132 (N_6132,N_5825,N_5597);
xor U6133 (N_6133,N_5594,N_5503);
nor U6134 (N_6134,N_5621,N_5847);
or U6135 (N_6135,N_5514,N_5958);
and U6136 (N_6136,N_5820,N_5955);
and U6137 (N_6137,N_5650,N_5715);
nand U6138 (N_6138,N_5919,N_5985);
nor U6139 (N_6139,N_5504,N_5547);
and U6140 (N_6140,N_5768,N_5718);
nand U6141 (N_6141,N_5578,N_5669);
xnor U6142 (N_6142,N_5838,N_5743);
nor U6143 (N_6143,N_5956,N_5574);
nor U6144 (N_6144,N_5528,N_5575);
nand U6145 (N_6145,N_5572,N_5618);
xnor U6146 (N_6146,N_5850,N_5737);
nor U6147 (N_6147,N_5508,N_5565);
nand U6148 (N_6148,N_5625,N_5872);
or U6149 (N_6149,N_5555,N_5807);
xnor U6150 (N_6150,N_5873,N_5677);
nand U6151 (N_6151,N_5995,N_5614);
and U6152 (N_6152,N_5550,N_5588);
nand U6153 (N_6153,N_5813,N_5671);
nor U6154 (N_6154,N_5568,N_5725);
and U6155 (N_6155,N_5814,N_5897);
or U6156 (N_6156,N_5699,N_5760);
or U6157 (N_6157,N_5619,N_5604);
nand U6158 (N_6158,N_5823,N_5731);
or U6159 (N_6159,N_5561,N_5864);
xnor U6160 (N_6160,N_5769,N_5543);
and U6161 (N_6161,N_5583,N_5573);
nand U6162 (N_6162,N_5888,N_5811);
and U6163 (N_6163,N_5915,N_5961);
nand U6164 (N_6164,N_5790,N_5895);
or U6165 (N_6165,N_5622,N_5634);
nor U6166 (N_6166,N_5829,N_5721);
or U6167 (N_6167,N_5640,N_5982);
nand U6168 (N_6168,N_5685,N_5509);
nor U6169 (N_6169,N_5539,N_5582);
nand U6170 (N_6170,N_5834,N_5649);
xnor U6171 (N_6171,N_5676,N_5809);
nor U6172 (N_6172,N_5683,N_5589);
and U6173 (N_6173,N_5631,N_5522);
or U6174 (N_6174,N_5513,N_5984);
and U6175 (N_6175,N_5913,N_5861);
xor U6176 (N_6176,N_5746,N_5665);
nor U6177 (N_6177,N_5552,N_5591);
nor U6178 (N_6178,N_5795,N_5858);
or U6179 (N_6179,N_5800,N_5816);
nand U6180 (N_6180,N_5763,N_5576);
nand U6181 (N_6181,N_5641,N_5639);
xnor U6182 (N_6182,N_5534,N_5626);
and U6183 (N_6183,N_5730,N_5903);
nor U6184 (N_6184,N_5901,N_5602);
nand U6185 (N_6185,N_5537,N_5970);
nand U6186 (N_6186,N_5726,N_5856);
or U6187 (N_6187,N_5510,N_5869);
xnor U6188 (N_6188,N_5988,N_5940);
or U6189 (N_6189,N_5971,N_5761);
nor U6190 (N_6190,N_5876,N_5968);
xor U6191 (N_6191,N_5846,N_5651);
or U6192 (N_6192,N_5538,N_5817);
or U6193 (N_6193,N_5637,N_5841);
or U6194 (N_6194,N_5973,N_5607);
nor U6195 (N_6195,N_5899,N_5780);
xor U6196 (N_6196,N_5532,N_5914);
or U6197 (N_6197,N_5520,N_5863);
and U6198 (N_6198,N_5776,N_5927);
or U6199 (N_6199,N_5871,N_5587);
nor U6200 (N_6200,N_5515,N_5603);
and U6201 (N_6201,N_5922,N_5957);
xnor U6202 (N_6202,N_5862,N_5609);
and U6203 (N_6203,N_5892,N_5660);
xor U6204 (N_6204,N_5826,N_5934);
xor U6205 (N_6205,N_5615,N_5533);
and U6206 (N_6206,N_5606,N_5648);
xnor U6207 (N_6207,N_5828,N_5939);
and U6208 (N_6208,N_5924,N_5563);
nand U6209 (N_6209,N_5540,N_5978);
xor U6210 (N_6210,N_5949,N_5819);
and U6211 (N_6211,N_5921,N_5655);
nand U6212 (N_6212,N_5710,N_5758);
nor U6213 (N_6213,N_5801,N_5756);
xor U6214 (N_6214,N_5579,N_5596);
xor U6215 (N_6215,N_5855,N_5808);
or U6216 (N_6216,N_5883,N_5799);
nor U6217 (N_6217,N_5929,N_5831);
and U6218 (N_6218,N_5500,N_5749);
or U6219 (N_6219,N_5881,N_5580);
and U6220 (N_6220,N_5975,N_5782);
nor U6221 (N_6221,N_5627,N_5798);
nand U6222 (N_6222,N_5735,N_5724);
or U6223 (N_6223,N_5632,N_5900);
xor U6224 (N_6224,N_5953,N_5518);
and U6225 (N_6225,N_5793,N_5837);
or U6226 (N_6226,N_5643,N_5645);
and U6227 (N_6227,N_5950,N_5916);
nor U6228 (N_6228,N_5844,N_5875);
nor U6229 (N_6229,N_5878,N_5738);
nand U6230 (N_6230,N_5595,N_5993);
and U6231 (N_6231,N_5839,N_5952);
nor U6232 (N_6232,N_5605,N_5559);
and U6233 (N_6233,N_5535,N_5647);
nor U6234 (N_6234,N_5701,N_5663);
nor U6235 (N_6235,N_5570,N_5884);
or U6236 (N_6236,N_5796,N_5774);
or U6237 (N_6237,N_5523,N_5695);
and U6238 (N_6238,N_5608,N_5833);
or U6239 (N_6239,N_5728,N_5785);
xor U6240 (N_6240,N_5773,N_5759);
nand U6241 (N_6241,N_5752,N_5687);
xnor U6242 (N_6242,N_5980,N_5840);
nand U6243 (N_6243,N_5707,N_5979);
or U6244 (N_6244,N_5910,N_5517);
xnor U6245 (N_6245,N_5986,N_5997);
and U6246 (N_6246,N_5646,N_5936);
nand U6247 (N_6247,N_5633,N_5652);
xnor U6248 (N_6248,N_5781,N_5882);
xor U6249 (N_6249,N_5674,N_5531);
or U6250 (N_6250,N_5887,N_5600);
xnor U6251 (N_6251,N_5626,N_5743);
xnor U6252 (N_6252,N_5724,N_5719);
nor U6253 (N_6253,N_5948,N_5646);
and U6254 (N_6254,N_5859,N_5999);
and U6255 (N_6255,N_5590,N_5609);
nor U6256 (N_6256,N_5625,N_5532);
nand U6257 (N_6257,N_5749,N_5645);
xnor U6258 (N_6258,N_5777,N_5741);
nand U6259 (N_6259,N_5661,N_5700);
nand U6260 (N_6260,N_5535,N_5568);
or U6261 (N_6261,N_5860,N_5848);
nand U6262 (N_6262,N_5508,N_5848);
nor U6263 (N_6263,N_5690,N_5745);
nor U6264 (N_6264,N_5516,N_5877);
and U6265 (N_6265,N_5610,N_5794);
or U6266 (N_6266,N_5723,N_5841);
nand U6267 (N_6267,N_5543,N_5592);
or U6268 (N_6268,N_5600,N_5550);
and U6269 (N_6269,N_5623,N_5766);
nand U6270 (N_6270,N_5511,N_5505);
and U6271 (N_6271,N_5964,N_5794);
or U6272 (N_6272,N_5999,N_5782);
xnor U6273 (N_6273,N_5782,N_5577);
nor U6274 (N_6274,N_5881,N_5912);
xor U6275 (N_6275,N_5633,N_5770);
and U6276 (N_6276,N_5786,N_5677);
xor U6277 (N_6277,N_5829,N_5963);
xnor U6278 (N_6278,N_5748,N_5546);
xor U6279 (N_6279,N_5947,N_5598);
nand U6280 (N_6280,N_5737,N_5776);
or U6281 (N_6281,N_5930,N_5959);
nand U6282 (N_6282,N_5971,N_5675);
or U6283 (N_6283,N_5577,N_5777);
nor U6284 (N_6284,N_5588,N_5843);
and U6285 (N_6285,N_5954,N_5633);
xor U6286 (N_6286,N_5942,N_5836);
xnor U6287 (N_6287,N_5654,N_5878);
or U6288 (N_6288,N_5619,N_5898);
xor U6289 (N_6289,N_5723,N_5799);
nor U6290 (N_6290,N_5667,N_5837);
and U6291 (N_6291,N_5876,N_5692);
nand U6292 (N_6292,N_5756,N_5989);
and U6293 (N_6293,N_5741,N_5568);
or U6294 (N_6294,N_5728,N_5830);
nand U6295 (N_6295,N_5856,N_5666);
and U6296 (N_6296,N_5849,N_5729);
and U6297 (N_6297,N_5745,N_5679);
and U6298 (N_6298,N_5578,N_5981);
or U6299 (N_6299,N_5857,N_5770);
xnor U6300 (N_6300,N_5657,N_5530);
nand U6301 (N_6301,N_5554,N_5658);
nand U6302 (N_6302,N_5643,N_5998);
and U6303 (N_6303,N_5744,N_5974);
and U6304 (N_6304,N_5928,N_5700);
and U6305 (N_6305,N_5747,N_5533);
and U6306 (N_6306,N_5695,N_5968);
or U6307 (N_6307,N_5640,N_5738);
nor U6308 (N_6308,N_5731,N_5762);
xnor U6309 (N_6309,N_5620,N_5739);
xor U6310 (N_6310,N_5953,N_5554);
nand U6311 (N_6311,N_5512,N_5879);
xor U6312 (N_6312,N_5694,N_5863);
nand U6313 (N_6313,N_5841,N_5638);
nand U6314 (N_6314,N_5682,N_5657);
nor U6315 (N_6315,N_5705,N_5514);
nand U6316 (N_6316,N_5693,N_5537);
or U6317 (N_6317,N_5833,N_5927);
xor U6318 (N_6318,N_5692,N_5987);
nand U6319 (N_6319,N_5648,N_5609);
or U6320 (N_6320,N_5807,N_5558);
nand U6321 (N_6321,N_5767,N_5683);
and U6322 (N_6322,N_5648,N_5861);
and U6323 (N_6323,N_5758,N_5734);
nor U6324 (N_6324,N_5518,N_5740);
or U6325 (N_6325,N_5613,N_5785);
nor U6326 (N_6326,N_5685,N_5861);
and U6327 (N_6327,N_5714,N_5831);
and U6328 (N_6328,N_5548,N_5544);
or U6329 (N_6329,N_5619,N_5591);
nor U6330 (N_6330,N_5775,N_5788);
xor U6331 (N_6331,N_5542,N_5697);
nor U6332 (N_6332,N_5821,N_5787);
xor U6333 (N_6333,N_5585,N_5749);
or U6334 (N_6334,N_5835,N_5507);
nor U6335 (N_6335,N_5718,N_5506);
or U6336 (N_6336,N_5705,N_5801);
nor U6337 (N_6337,N_5922,N_5718);
or U6338 (N_6338,N_5601,N_5990);
and U6339 (N_6339,N_5909,N_5638);
or U6340 (N_6340,N_5935,N_5501);
or U6341 (N_6341,N_5620,N_5690);
xor U6342 (N_6342,N_5760,N_5692);
nand U6343 (N_6343,N_5969,N_5734);
and U6344 (N_6344,N_5606,N_5612);
xnor U6345 (N_6345,N_5813,N_5822);
nand U6346 (N_6346,N_5700,N_5962);
xnor U6347 (N_6347,N_5847,N_5839);
or U6348 (N_6348,N_5699,N_5718);
xnor U6349 (N_6349,N_5573,N_5593);
or U6350 (N_6350,N_5529,N_5860);
nand U6351 (N_6351,N_5702,N_5797);
and U6352 (N_6352,N_5535,N_5511);
or U6353 (N_6353,N_5642,N_5854);
nor U6354 (N_6354,N_5919,N_5513);
nand U6355 (N_6355,N_5884,N_5628);
xnor U6356 (N_6356,N_5630,N_5940);
nand U6357 (N_6357,N_5569,N_5612);
nand U6358 (N_6358,N_5733,N_5654);
xor U6359 (N_6359,N_5835,N_5513);
or U6360 (N_6360,N_5629,N_5901);
xor U6361 (N_6361,N_5781,N_5522);
xor U6362 (N_6362,N_5684,N_5503);
nand U6363 (N_6363,N_5921,N_5503);
nand U6364 (N_6364,N_5660,N_5795);
and U6365 (N_6365,N_5925,N_5621);
nor U6366 (N_6366,N_5931,N_5775);
nand U6367 (N_6367,N_5540,N_5512);
nand U6368 (N_6368,N_5525,N_5509);
or U6369 (N_6369,N_5622,N_5990);
or U6370 (N_6370,N_5699,N_5507);
and U6371 (N_6371,N_5519,N_5689);
xnor U6372 (N_6372,N_5864,N_5558);
xor U6373 (N_6373,N_5632,N_5951);
xnor U6374 (N_6374,N_5536,N_5527);
and U6375 (N_6375,N_5883,N_5877);
xnor U6376 (N_6376,N_5573,N_5536);
and U6377 (N_6377,N_5768,N_5636);
and U6378 (N_6378,N_5981,N_5748);
nor U6379 (N_6379,N_5906,N_5928);
and U6380 (N_6380,N_5543,N_5770);
xor U6381 (N_6381,N_5548,N_5787);
nand U6382 (N_6382,N_5741,N_5975);
xnor U6383 (N_6383,N_5743,N_5797);
or U6384 (N_6384,N_5955,N_5882);
and U6385 (N_6385,N_5653,N_5649);
or U6386 (N_6386,N_5841,N_5893);
and U6387 (N_6387,N_5546,N_5993);
and U6388 (N_6388,N_5504,N_5632);
and U6389 (N_6389,N_5526,N_5852);
and U6390 (N_6390,N_5825,N_5898);
nand U6391 (N_6391,N_5797,N_5822);
nand U6392 (N_6392,N_5571,N_5676);
xor U6393 (N_6393,N_5810,N_5838);
xnor U6394 (N_6394,N_5878,N_5681);
nor U6395 (N_6395,N_5626,N_5823);
nand U6396 (N_6396,N_5994,N_5611);
xor U6397 (N_6397,N_5643,N_5972);
nor U6398 (N_6398,N_5622,N_5853);
or U6399 (N_6399,N_5794,N_5686);
nor U6400 (N_6400,N_5767,N_5625);
and U6401 (N_6401,N_5650,N_5523);
nand U6402 (N_6402,N_5856,N_5756);
nand U6403 (N_6403,N_5950,N_5649);
xor U6404 (N_6404,N_5900,N_5977);
or U6405 (N_6405,N_5898,N_5552);
and U6406 (N_6406,N_5797,N_5796);
and U6407 (N_6407,N_5801,N_5687);
or U6408 (N_6408,N_5579,N_5609);
nand U6409 (N_6409,N_5890,N_5821);
nor U6410 (N_6410,N_5978,N_5760);
nor U6411 (N_6411,N_5983,N_5932);
nand U6412 (N_6412,N_5586,N_5717);
xnor U6413 (N_6413,N_5691,N_5946);
or U6414 (N_6414,N_5868,N_5914);
or U6415 (N_6415,N_5807,N_5817);
and U6416 (N_6416,N_5506,N_5887);
nor U6417 (N_6417,N_5537,N_5771);
nand U6418 (N_6418,N_5998,N_5932);
nor U6419 (N_6419,N_5965,N_5634);
and U6420 (N_6420,N_5971,N_5855);
nor U6421 (N_6421,N_5643,N_5920);
xnor U6422 (N_6422,N_5933,N_5885);
and U6423 (N_6423,N_5542,N_5675);
or U6424 (N_6424,N_5948,N_5849);
nand U6425 (N_6425,N_5500,N_5814);
nor U6426 (N_6426,N_5997,N_5968);
nor U6427 (N_6427,N_5829,N_5618);
xor U6428 (N_6428,N_5561,N_5776);
or U6429 (N_6429,N_5552,N_5945);
nand U6430 (N_6430,N_5916,N_5823);
or U6431 (N_6431,N_5601,N_5789);
or U6432 (N_6432,N_5988,N_5771);
and U6433 (N_6433,N_5920,N_5610);
nor U6434 (N_6434,N_5522,N_5717);
xnor U6435 (N_6435,N_5523,N_5732);
nand U6436 (N_6436,N_5559,N_5707);
xnor U6437 (N_6437,N_5514,N_5981);
nand U6438 (N_6438,N_5516,N_5515);
or U6439 (N_6439,N_5922,N_5768);
and U6440 (N_6440,N_5851,N_5981);
nor U6441 (N_6441,N_5552,N_5987);
nor U6442 (N_6442,N_5924,N_5971);
or U6443 (N_6443,N_5750,N_5753);
and U6444 (N_6444,N_5993,N_5583);
and U6445 (N_6445,N_5963,N_5946);
and U6446 (N_6446,N_5531,N_5794);
xnor U6447 (N_6447,N_5687,N_5700);
xor U6448 (N_6448,N_5665,N_5964);
and U6449 (N_6449,N_5922,N_5621);
and U6450 (N_6450,N_5719,N_5686);
or U6451 (N_6451,N_5711,N_5653);
or U6452 (N_6452,N_5920,N_5642);
xnor U6453 (N_6453,N_5797,N_5798);
or U6454 (N_6454,N_5871,N_5606);
xnor U6455 (N_6455,N_5700,N_5621);
or U6456 (N_6456,N_5525,N_5670);
and U6457 (N_6457,N_5572,N_5802);
nor U6458 (N_6458,N_5727,N_5798);
and U6459 (N_6459,N_5716,N_5879);
xor U6460 (N_6460,N_5822,N_5896);
nor U6461 (N_6461,N_5566,N_5740);
and U6462 (N_6462,N_5708,N_5621);
and U6463 (N_6463,N_5505,N_5965);
or U6464 (N_6464,N_5703,N_5565);
nor U6465 (N_6465,N_5509,N_5693);
xor U6466 (N_6466,N_5841,N_5717);
or U6467 (N_6467,N_5657,N_5872);
or U6468 (N_6468,N_5755,N_5597);
nand U6469 (N_6469,N_5518,N_5597);
nand U6470 (N_6470,N_5944,N_5598);
nor U6471 (N_6471,N_5940,N_5681);
nor U6472 (N_6472,N_5949,N_5778);
nor U6473 (N_6473,N_5809,N_5619);
xor U6474 (N_6474,N_5618,N_5852);
or U6475 (N_6475,N_5901,N_5793);
xnor U6476 (N_6476,N_5688,N_5906);
or U6477 (N_6477,N_5732,N_5919);
xor U6478 (N_6478,N_5794,N_5734);
or U6479 (N_6479,N_5565,N_5888);
or U6480 (N_6480,N_5986,N_5954);
or U6481 (N_6481,N_5601,N_5575);
or U6482 (N_6482,N_5629,N_5814);
and U6483 (N_6483,N_5782,N_5621);
or U6484 (N_6484,N_5756,N_5674);
nor U6485 (N_6485,N_5986,N_5516);
and U6486 (N_6486,N_5548,N_5686);
nand U6487 (N_6487,N_5875,N_5763);
xnor U6488 (N_6488,N_5819,N_5636);
or U6489 (N_6489,N_5583,N_5727);
xnor U6490 (N_6490,N_5799,N_5662);
nor U6491 (N_6491,N_5946,N_5752);
nor U6492 (N_6492,N_5530,N_5791);
or U6493 (N_6493,N_5762,N_5715);
and U6494 (N_6494,N_5646,N_5680);
and U6495 (N_6495,N_5692,N_5512);
nor U6496 (N_6496,N_5874,N_5958);
xnor U6497 (N_6497,N_5941,N_5659);
or U6498 (N_6498,N_5932,N_5611);
or U6499 (N_6499,N_5817,N_5912);
or U6500 (N_6500,N_6211,N_6061);
nand U6501 (N_6501,N_6271,N_6177);
or U6502 (N_6502,N_6282,N_6070);
nand U6503 (N_6503,N_6472,N_6010);
nand U6504 (N_6504,N_6214,N_6000);
or U6505 (N_6505,N_6264,N_6315);
or U6506 (N_6506,N_6456,N_6018);
or U6507 (N_6507,N_6170,N_6189);
and U6508 (N_6508,N_6122,N_6247);
nor U6509 (N_6509,N_6188,N_6308);
or U6510 (N_6510,N_6489,N_6168);
xor U6511 (N_6511,N_6408,N_6280);
nor U6512 (N_6512,N_6059,N_6160);
or U6513 (N_6513,N_6394,N_6399);
nor U6514 (N_6514,N_6361,N_6058);
or U6515 (N_6515,N_6080,N_6116);
xor U6516 (N_6516,N_6413,N_6419);
nor U6517 (N_6517,N_6192,N_6292);
and U6518 (N_6518,N_6143,N_6216);
nor U6519 (N_6519,N_6106,N_6141);
xor U6520 (N_6520,N_6120,N_6405);
xnor U6521 (N_6521,N_6261,N_6069);
nand U6522 (N_6522,N_6398,N_6378);
nand U6523 (N_6523,N_6017,N_6171);
or U6524 (N_6524,N_6083,N_6291);
and U6525 (N_6525,N_6217,N_6497);
xnor U6526 (N_6526,N_6289,N_6479);
nor U6527 (N_6527,N_6415,N_6397);
and U6528 (N_6528,N_6440,N_6457);
and U6529 (N_6529,N_6037,N_6125);
nor U6530 (N_6530,N_6156,N_6244);
or U6531 (N_6531,N_6387,N_6030);
nand U6532 (N_6532,N_6197,N_6102);
and U6533 (N_6533,N_6429,N_6184);
nor U6534 (N_6534,N_6339,N_6057);
xor U6535 (N_6535,N_6038,N_6130);
nor U6536 (N_6536,N_6180,N_6380);
nand U6537 (N_6537,N_6442,N_6263);
xor U6538 (N_6538,N_6307,N_6224);
xnor U6539 (N_6539,N_6234,N_6402);
xor U6540 (N_6540,N_6097,N_6270);
xnor U6541 (N_6541,N_6368,N_6461);
nor U6542 (N_6542,N_6432,N_6022);
xor U6543 (N_6543,N_6367,N_6464);
and U6544 (N_6544,N_6446,N_6255);
nor U6545 (N_6545,N_6093,N_6275);
nand U6546 (N_6546,N_6135,N_6194);
nor U6547 (N_6547,N_6006,N_6233);
nor U6548 (N_6548,N_6332,N_6101);
and U6549 (N_6549,N_6054,N_6055);
or U6550 (N_6550,N_6240,N_6266);
or U6551 (N_6551,N_6047,N_6203);
and U6552 (N_6552,N_6029,N_6014);
nor U6553 (N_6553,N_6441,N_6322);
and U6554 (N_6554,N_6311,N_6436);
xor U6555 (N_6555,N_6258,N_6334);
nor U6556 (N_6556,N_6366,N_6096);
xnor U6557 (N_6557,N_6024,N_6320);
and U6558 (N_6558,N_6021,N_6046);
or U6559 (N_6559,N_6283,N_6187);
and U6560 (N_6560,N_6483,N_6401);
or U6561 (N_6561,N_6041,N_6357);
xnor U6562 (N_6562,N_6218,N_6068);
nand U6563 (N_6563,N_6081,N_6237);
nor U6564 (N_6564,N_6065,N_6288);
and U6565 (N_6565,N_6485,N_6229);
and U6566 (N_6566,N_6004,N_6133);
or U6567 (N_6567,N_6092,N_6050);
and U6568 (N_6568,N_6467,N_6443);
xnor U6569 (N_6569,N_6012,N_6153);
or U6570 (N_6570,N_6164,N_6369);
and U6571 (N_6571,N_6300,N_6238);
xnor U6572 (N_6572,N_6067,N_6243);
nor U6573 (N_6573,N_6063,N_6294);
nor U6574 (N_6574,N_6466,N_6403);
or U6575 (N_6575,N_6363,N_6144);
nor U6576 (N_6576,N_6202,N_6343);
xor U6577 (N_6577,N_6314,N_6468);
nor U6578 (N_6578,N_6128,N_6252);
or U6579 (N_6579,N_6365,N_6354);
and U6580 (N_6580,N_6213,N_6301);
or U6581 (N_6581,N_6114,N_6349);
or U6582 (N_6582,N_6395,N_6140);
nor U6583 (N_6583,N_6273,N_6094);
or U6584 (N_6584,N_6250,N_6009);
nor U6585 (N_6585,N_6048,N_6480);
or U6586 (N_6586,N_6458,N_6245);
nor U6587 (N_6587,N_6286,N_6195);
nor U6588 (N_6588,N_6073,N_6148);
or U6589 (N_6589,N_6477,N_6089);
and U6590 (N_6590,N_6392,N_6154);
and U6591 (N_6591,N_6227,N_6199);
xnor U6592 (N_6592,N_6269,N_6118);
nor U6593 (N_6593,N_6129,N_6166);
nor U6594 (N_6594,N_6036,N_6391);
nand U6595 (N_6595,N_6103,N_6113);
xor U6596 (N_6596,N_6494,N_6410);
and U6597 (N_6597,N_6345,N_6381);
nor U6598 (N_6598,N_6032,N_6099);
and U6599 (N_6599,N_6033,N_6279);
xor U6600 (N_6600,N_6223,N_6182);
or U6601 (N_6601,N_6191,N_6326);
or U6602 (N_6602,N_6246,N_6299);
xnor U6603 (N_6603,N_6152,N_6277);
nor U6604 (N_6604,N_6469,N_6016);
and U6605 (N_6605,N_6186,N_6151);
nand U6606 (N_6606,N_6404,N_6045);
xnor U6607 (N_6607,N_6475,N_6231);
xor U6608 (N_6608,N_6221,N_6496);
and U6609 (N_6609,N_6344,N_6318);
nand U6610 (N_6610,N_6384,N_6005);
xor U6611 (N_6611,N_6169,N_6139);
nand U6612 (N_6612,N_6178,N_6165);
xor U6613 (N_6613,N_6400,N_6385);
nor U6614 (N_6614,N_6262,N_6420);
nand U6615 (N_6615,N_6185,N_6425);
or U6616 (N_6616,N_6253,N_6312);
nor U6617 (N_6617,N_6064,N_6051);
nand U6618 (N_6618,N_6268,N_6236);
nor U6619 (N_6619,N_6205,N_6181);
nand U6620 (N_6620,N_6082,N_6276);
xnor U6621 (N_6621,N_6444,N_6007);
nor U6622 (N_6622,N_6370,N_6232);
and U6623 (N_6623,N_6119,N_6492);
nand U6624 (N_6624,N_6417,N_6430);
nor U6625 (N_6625,N_6147,N_6281);
and U6626 (N_6626,N_6302,N_6439);
xnor U6627 (N_6627,N_6379,N_6355);
nor U6628 (N_6628,N_6450,N_6060);
nor U6629 (N_6629,N_6137,N_6418);
and U6630 (N_6630,N_6157,N_6407);
xnor U6631 (N_6631,N_6481,N_6452);
nand U6632 (N_6632,N_6179,N_6138);
or U6633 (N_6633,N_6470,N_6115);
or U6634 (N_6634,N_6167,N_6319);
nor U6635 (N_6635,N_6306,N_6206);
xor U6636 (N_6636,N_6110,N_6323);
nand U6637 (N_6637,N_6325,N_6296);
nor U6638 (N_6638,N_6026,N_6331);
xnor U6639 (N_6639,N_6040,N_6098);
or U6640 (N_6640,N_6132,N_6356);
nor U6641 (N_6641,N_6196,N_6267);
nor U6642 (N_6642,N_6136,N_6454);
or U6643 (N_6643,N_6389,N_6134);
or U6644 (N_6644,N_6256,N_6207);
or U6645 (N_6645,N_6412,N_6066);
nor U6646 (N_6646,N_6297,N_6438);
and U6647 (N_6647,N_6215,N_6155);
and U6648 (N_6648,N_6249,N_6053);
xor U6649 (N_6649,N_6117,N_6020);
and U6650 (N_6650,N_6406,N_6085);
xnor U6651 (N_6651,N_6358,N_6107);
xor U6652 (N_6652,N_6304,N_6493);
nand U6653 (N_6653,N_6003,N_6421);
and U6654 (N_6654,N_6422,N_6112);
and U6655 (N_6655,N_6340,N_6044);
or U6656 (N_6656,N_6084,N_6172);
nor U6657 (N_6657,N_6210,N_6198);
or U6658 (N_6658,N_6465,N_6011);
xnor U6659 (N_6659,N_6393,N_6201);
nor U6660 (N_6660,N_6248,N_6149);
nand U6661 (N_6661,N_6478,N_6251);
nor U6662 (N_6662,N_6341,N_6431);
or U6663 (N_6663,N_6150,N_6174);
nand U6664 (N_6664,N_6490,N_6414);
xnor U6665 (N_6665,N_6228,N_6162);
or U6666 (N_6666,N_6337,N_6310);
or U6667 (N_6667,N_6025,N_6290);
or U6668 (N_6668,N_6142,N_6163);
and U6669 (N_6669,N_6409,N_6382);
nand U6670 (N_6670,N_6459,N_6127);
and U6671 (N_6671,N_6056,N_6086);
nand U6672 (N_6672,N_6445,N_6049);
and U6673 (N_6673,N_6293,N_6131);
or U6674 (N_6674,N_6338,N_6390);
and U6675 (N_6675,N_6284,N_6230);
nand U6676 (N_6676,N_6328,N_6287);
or U6677 (N_6677,N_6434,N_6108);
or U6678 (N_6678,N_6019,N_6330);
xnor U6679 (N_6679,N_6274,N_6491);
or U6680 (N_6680,N_6109,N_6352);
nand U6681 (N_6681,N_6145,N_6348);
xor U6682 (N_6682,N_6208,N_6495);
or U6683 (N_6683,N_6462,N_6071);
and U6684 (N_6684,N_6100,N_6242);
or U6685 (N_6685,N_6176,N_6448);
and U6686 (N_6686,N_6427,N_6321);
nand U6687 (N_6687,N_6173,N_6435);
nand U6688 (N_6688,N_6376,N_6200);
xnor U6689 (N_6689,N_6183,N_6476);
nor U6690 (N_6690,N_6002,N_6375);
nand U6691 (N_6691,N_6074,N_6090);
nor U6692 (N_6692,N_6374,N_6034);
nand U6693 (N_6693,N_6272,N_6447);
xor U6694 (N_6694,N_6079,N_6072);
and U6695 (N_6695,N_6031,N_6226);
nor U6696 (N_6696,N_6313,N_6042);
nand U6697 (N_6697,N_6126,N_6499);
xor U6698 (N_6698,N_6416,N_6295);
or U6699 (N_6699,N_6039,N_6222);
and U6700 (N_6700,N_6035,N_6460);
xnor U6701 (N_6701,N_6449,N_6105);
and U6702 (N_6702,N_6335,N_6377);
xor U6703 (N_6703,N_6396,N_6235);
nand U6704 (N_6704,N_6383,N_6124);
or U6705 (N_6705,N_6241,N_6372);
nor U6706 (N_6706,N_6471,N_6316);
or U6707 (N_6707,N_6346,N_6350);
nor U6708 (N_6708,N_6091,N_6209);
nor U6709 (N_6709,N_6161,N_6373);
xor U6710 (N_6710,N_6265,N_6437);
nand U6711 (N_6711,N_6424,N_6062);
or U6712 (N_6712,N_6159,N_6052);
nand U6713 (N_6713,N_6333,N_6305);
or U6714 (N_6714,N_6453,N_6123);
nand U6715 (N_6715,N_6121,N_6342);
or U6716 (N_6716,N_6087,N_6487);
or U6717 (N_6717,N_6474,N_6078);
xnor U6718 (N_6718,N_6254,N_6239);
nor U6719 (N_6719,N_6360,N_6204);
or U6720 (N_6720,N_6455,N_6327);
nor U6721 (N_6721,N_6008,N_6027);
nor U6722 (N_6722,N_6076,N_6353);
and U6723 (N_6723,N_6104,N_6303);
and U6724 (N_6724,N_6219,N_6451);
or U6725 (N_6725,N_6386,N_6193);
nor U6726 (N_6726,N_6488,N_6146);
or U6727 (N_6727,N_6023,N_6324);
nand U6728 (N_6728,N_6362,N_6175);
or U6729 (N_6729,N_6388,N_6482);
nor U6730 (N_6730,N_6001,N_6309);
nand U6731 (N_6731,N_6317,N_6463);
xor U6732 (N_6732,N_6095,N_6111);
xnor U6733 (N_6733,N_6498,N_6473);
nor U6734 (N_6734,N_6075,N_6329);
nand U6735 (N_6735,N_6433,N_6077);
xnor U6736 (N_6736,N_6484,N_6088);
nor U6737 (N_6737,N_6260,N_6043);
nand U6738 (N_6738,N_6351,N_6259);
xnor U6739 (N_6739,N_6285,N_6426);
and U6740 (N_6740,N_6013,N_6347);
nand U6741 (N_6741,N_6359,N_6212);
nor U6742 (N_6742,N_6428,N_6423);
or U6743 (N_6743,N_6158,N_6336);
nand U6744 (N_6744,N_6225,N_6298);
nor U6745 (N_6745,N_6015,N_6190);
and U6746 (N_6746,N_6278,N_6486);
and U6747 (N_6747,N_6028,N_6220);
nand U6748 (N_6748,N_6411,N_6257);
and U6749 (N_6749,N_6371,N_6364);
or U6750 (N_6750,N_6084,N_6117);
and U6751 (N_6751,N_6060,N_6058);
and U6752 (N_6752,N_6033,N_6168);
or U6753 (N_6753,N_6346,N_6254);
xnor U6754 (N_6754,N_6060,N_6353);
or U6755 (N_6755,N_6001,N_6483);
and U6756 (N_6756,N_6226,N_6369);
nor U6757 (N_6757,N_6181,N_6402);
nor U6758 (N_6758,N_6010,N_6350);
nand U6759 (N_6759,N_6292,N_6354);
and U6760 (N_6760,N_6039,N_6298);
or U6761 (N_6761,N_6403,N_6258);
or U6762 (N_6762,N_6419,N_6038);
xor U6763 (N_6763,N_6300,N_6419);
nand U6764 (N_6764,N_6451,N_6192);
nand U6765 (N_6765,N_6468,N_6033);
xor U6766 (N_6766,N_6045,N_6418);
xnor U6767 (N_6767,N_6358,N_6340);
or U6768 (N_6768,N_6410,N_6135);
nand U6769 (N_6769,N_6333,N_6278);
nand U6770 (N_6770,N_6477,N_6279);
and U6771 (N_6771,N_6213,N_6054);
nand U6772 (N_6772,N_6295,N_6074);
and U6773 (N_6773,N_6029,N_6438);
and U6774 (N_6774,N_6237,N_6350);
xor U6775 (N_6775,N_6047,N_6315);
or U6776 (N_6776,N_6213,N_6165);
xor U6777 (N_6777,N_6237,N_6003);
nor U6778 (N_6778,N_6071,N_6023);
nand U6779 (N_6779,N_6189,N_6448);
and U6780 (N_6780,N_6226,N_6423);
or U6781 (N_6781,N_6185,N_6342);
xor U6782 (N_6782,N_6479,N_6193);
or U6783 (N_6783,N_6346,N_6005);
nor U6784 (N_6784,N_6485,N_6216);
xnor U6785 (N_6785,N_6093,N_6071);
nor U6786 (N_6786,N_6367,N_6096);
xor U6787 (N_6787,N_6241,N_6265);
xor U6788 (N_6788,N_6172,N_6111);
xnor U6789 (N_6789,N_6220,N_6052);
or U6790 (N_6790,N_6267,N_6164);
and U6791 (N_6791,N_6227,N_6482);
xor U6792 (N_6792,N_6003,N_6446);
or U6793 (N_6793,N_6484,N_6011);
nor U6794 (N_6794,N_6005,N_6031);
xnor U6795 (N_6795,N_6069,N_6349);
or U6796 (N_6796,N_6370,N_6259);
xor U6797 (N_6797,N_6112,N_6158);
nor U6798 (N_6798,N_6100,N_6072);
nor U6799 (N_6799,N_6067,N_6499);
nand U6800 (N_6800,N_6265,N_6185);
or U6801 (N_6801,N_6059,N_6126);
xor U6802 (N_6802,N_6018,N_6448);
or U6803 (N_6803,N_6140,N_6114);
nor U6804 (N_6804,N_6032,N_6324);
or U6805 (N_6805,N_6243,N_6392);
nor U6806 (N_6806,N_6274,N_6208);
nand U6807 (N_6807,N_6400,N_6006);
or U6808 (N_6808,N_6016,N_6305);
and U6809 (N_6809,N_6203,N_6073);
or U6810 (N_6810,N_6170,N_6283);
nand U6811 (N_6811,N_6333,N_6029);
nand U6812 (N_6812,N_6095,N_6213);
and U6813 (N_6813,N_6190,N_6235);
xnor U6814 (N_6814,N_6355,N_6094);
and U6815 (N_6815,N_6420,N_6135);
or U6816 (N_6816,N_6073,N_6305);
and U6817 (N_6817,N_6029,N_6107);
xnor U6818 (N_6818,N_6254,N_6127);
and U6819 (N_6819,N_6460,N_6407);
xor U6820 (N_6820,N_6306,N_6203);
xnor U6821 (N_6821,N_6180,N_6162);
xnor U6822 (N_6822,N_6181,N_6167);
nand U6823 (N_6823,N_6255,N_6182);
xnor U6824 (N_6824,N_6436,N_6046);
xnor U6825 (N_6825,N_6165,N_6224);
nand U6826 (N_6826,N_6046,N_6282);
or U6827 (N_6827,N_6040,N_6416);
nand U6828 (N_6828,N_6182,N_6032);
nor U6829 (N_6829,N_6304,N_6156);
nor U6830 (N_6830,N_6266,N_6142);
or U6831 (N_6831,N_6073,N_6420);
nor U6832 (N_6832,N_6286,N_6148);
xor U6833 (N_6833,N_6436,N_6403);
nor U6834 (N_6834,N_6152,N_6363);
and U6835 (N_6835,N_6485,N_6243);
nand U6836 (N_6836,N_6413,N_6225);
and U6837 (N_6837,N_6373,N_6478);
or U6838 (N_6838,N_6449,N_6192);
and U6839 (N_6839,N_6169,N_6216);
nor U6840 (N_6840,N_6149,N_6306);
nand U6841 (N_6841,N_6374,N_6288);
xor U6842 (N_6842,N_6080,N_6391);
xnor U6843 (N_6843,N_6196,N_6025);
nor U6844 (N_6844,N_6136,N_6332);
or U6845 (N_6845,N_6323,N_6223);
or U6846 (N_6846,N_6074,N_6113);
and U6847 (N_6847,N_6436,N_6438);
nand U6848 (N_6848,N_6086,N_6178);
and U6849 (N_6849,N_6040,N_6034);
nor U6850 (N_6850,N_6493,N_6408);
nor U6851 (N_6851,N_6482,N_6099);
nor U6852 (N_6852,N_6116,N_6377);
or U6853 (N_6853,N_6269,N_6061);
or U6854 (N_6854,N_6100,N_6458);
nor U6855 (N_6855,N_6117,N_6208);
nor U6856 (N_6856,N_6142,N_6062);
or U6857 (N_6857,N_6367,N_6048);
or U6858 (N_6858,N_6413,N_6183);
or U6859 (N_6859,N_6375,N_6160);
nand U6860 (N_6860,N_6469,N_6280);
nor U6861 (N_6861,N_6329,N_6465);
nand U6862 (N_6862,N_6244,N_6133);
xnor U6863 (N_6863,N_6142,N_6394);
xnor U6864 (N_6864,N_6413,N_6493);
nor U6865 (N_6865,N_6386,N_6350);
or U6866 (N_6866,N_6460,N_6322);
or U6867 (N_6867,N_6163,N_6202);
or U6868 (N_6868,N_6370,N_6154);
nor U6869 (N_6869,N_6477,N_6169);
nand U6870 (N_6870,N_6054,N_6152);
or U6871 (N_6871,N_6412,N_6020);
xnor U6872 (N_6872,N_6306,N_6148);
nand U6873 (N_6873,N_6362,N_6046);
nor U6874 (N_6874,N_6379,N_6046);
nor U6875 (N_6875,N_6113,N_6062);
nor U6876 (N_6876,N_6194,N_6174);
or U6877 (N_6877,N_6454,N_6448);
nand U6878 (N_6878,N_6369,N_6038);
xor U6879 (N_6879,N_6444,N_6179);
or U6880 (N_6880,N_6390,N_6352);
xor U6881 (N_6881,N_6479,N_6414);
and U6882 (N_6882,N_6071,N_6322);
or U6883 (N_6883,N_6326,N_6173);
and U6884 (N_6884,N_6401,N_6284);
or U6885 (N_6885,N_6411,N_6046);
and U6886 (N_6886,N_6280,N_6438);
and U6887 (N_6887,N_6393,N_6350);
or U6888 (N_6888,N_6323,N_6084);
and U6889 (N_6889,N_6040,N_6095);
nor U6890 (N_6890,N_6468,N_6209);
and U6891 (N_6891,N_6163,N_6151);
xnor U6892 (N_6892,N_6132,N_6142);
nand U6893 (N_6893,N_6397,N_6396);
nor U6894 (N_6894,N_6410,N_6237);
nand U6895 (N_6895,N_6449,N_6244);
or U6896 (N_6896,N_6335,N_6459);
nor U6897 (N_6897,N_6472,N_6169);
nand U6898 (N_6898,N_6044,N_6321);
nor U6899 (N_6899,N_6085,N_6478);
nand U6900 (N_6900,N_6412,N_6470);
nor U6901 (N_6901,N_6228,N_6232);
nor U6902 (N_6902,N_6064,N_6475);
xor U6903 (N_6903,N_6232,N_6151);
nor U6904 (N_6904,N_6308,N_6477);
xnor U6905 (N_6905,N_6216,N_6449);
and U6906 (N_6906,N_6103,N_6223);
nor U6907 (N_6907,N_6435,N_6177);
nand U6908 (N_6908,N_6287,N_6257);
xnor U6909 (N_6909,N_6269,N_6369);
nand U6910 (N_6910,N_6188,N_6199);
nor U6911 (N_6911,N_6271,N_6348);
and U6912 (N_6912,N_6241,N_6081);
or U6913 (N_6913,N_6445,N_6266);
nand U6914 (N_6914,N_6472,N_6224);
or U6915 (N_6915,N_6114,N_6426);
or U6916 (N_6916,N_6497,N_6139);
xnor U6917 (N_6917,N_6381,N_6162);
or U6918 (N_6918,N_6047,N_6215);
nor U6919 (N_6919,N_6489,N_6459);
nand U6920 (N_6920,N_6279,N_6147);
nand U6921 (N_6921,N_6272,N_6496);
and U6922 (N_6922,N_6121,N_6207);
nand U6923 (N_6923,N_6281,N_6005);
or U6924 (N_6924,N_6067,N_6248);
nor U6925 (N_6925,N_6377,N_6213);
nor U6926 (N_6926,N_6287,N_6146);
and U6927 (N_6927,N_6080,N_6499);
nand U6928 (N_6928,N_6105,N_6231);
nor U6929 (N_6929,N_6228,N_6317);
or U6930 (N_6930,N_6441,N_6398);
nor U6931 (N_6931,N_6308,N_6034);
nor U6932 (N_6932,N_6154,N_6014);
and U6933 (N_6933,N_6228,N_6364);
or U6934 (N_6934,N_6069,N_6463);
nor U6935 (N_6935,N_6209,N_6461);
nor U6936 (N_6936,N_6107,N_6293);
or U6937 (N_6937,N_6345,N_6152);
nand U6938 (N_6938,N_6091,N_6190);
xor U6939 (N_6939,N_6189,N_6288);
or U6940 (N_6940,N_6444,N_6429);
nand U6941 (N_6941,N_6260,N_6367);
nand U6942 (N_6942,N_6498,N_6206);
xor U6943 (N_6943,N_6027,N_6311);
or U6944 (N_6944,N_6013,N_6408);
and U6945 (N_6945,N_6064,N_6479);
xor U6946 (N_6946,N_6008,N_6205);
xor U6947 (N_6947,N_6477,N_6218);
or U6948 (N_6948,N_6349,N_6298);
and U6949 (N_6949,N_6059,N_6102);
nand U6950 (N_6950,N_6137,N_6062);
nor U6951 (N_6951,N_6316,N_6366);
nor U6952 (N_6952,N_6013,N_6314);
nand U6953 (N_6953,N_6452,N_6414);
nor U6954 (N_6954,N_6393,N_6349);
xor U6955 (N_6955,N_6352,N_6111);
and U6956 (N_6956,N_6223,N_6482);
nand U6957 (N_6957,N_6203,N_6384);
nor U6958 (N_6958,N_6305,N_6164);
or U6959 (N_6959,N_6118,N_6137);
or U6960 (N_6960,N_6406,N_6294);
and U6961 (N_6961,N_6376,N_6225);
xnor U6962 (N_6962,N_6107,N_6159);
nand U6963 (N_6963,N_6375,N_6138);
nor U6964 (N_6964,N_6090,N_6449);
xnor U6965 (N_6965,N_6116,N_6048);
nand U6966 (N_6966,N_6085,N_6472);
nand U6967 (N_6967,N_6090,N_6248);
nor U6968 (N_6968,N_6268,N_6289);
nor U6969 (N_6969,N_6472,N_6364);
xor U6970 (N_6970,N_6068,N_6465);
nand U6971 (N_6971,N_6264,N_6167);
nor U6972 (N_6972,N_6001,N_6467);
or U6973 (N_6973,N_6479,N_6254);
or U6974 (N_6974,N_6256,N_6098);
or U6975 (N_6975,N_6157,N_6431);
or U6976 (N_6976,N_6475,N_6078);
and U6977 (N_6977,N_6010,N_6173);
nor U6978 (N_6978,N_6331,N_6103);
and U6979 (N_6979,N_6495,N_6475);
nor U6980 (N_6980,N_6256,N_6365);
and U6981 (N_6981,N_6494,N_6238);
xnor U6982 (N_6982,N_6364,N_6407);
or U6983 (N_6983,N_6488,N_6068);
nand U6984 (N_6984,N_6014,N_6043);
or U6985 (N_6985,N_6177,N_6356);
nand U6986 (N_6986,N_6452,N_6145);
nor U6987 (N_6987,N_6197,N_6208);
or U6988 (N_6988,N_6251,N_6418);
or U6989 (N_6989,N_6412,N_6195);
nor U6990 (N_6990,N_6451,N_6095);
xor U6991 (N_6991,N_6121,N_6115);
and U6992 (N_6992,N_6411,N_6373);
nor U6993 (N_6993,N_6033,N_6406);
nor U6994 (N_6994,N_6415,N_6380);
or U6995 (N_6995,N_6407,N_6443);
or U6996 (N_6996,N_6403,N_6405);
xnor U6997 (N_6997,N_6397,N_6187);
xor U6998 (N_6998,N_6396,N_6086);
nand U6999 (N_6999,N_6233,N_6274);
xnor U7000 (N_7000,N_6764,N_6911);
nand U7001 (N_7001,N_6562,N_6663);
or U7002 (N_7002,N_6728,N_6887);
and U7003 (N_7003,N_6777,N_6950);
xor U7004 (N_7004,N_6673,N_6957);
nor U7005 (N_7005,N_6771,N_6891);
nand U7006 (N_7006,N_6884,N_6714);
or U7007 (N_7007,N_6840,N_6845);
and U7008 (N_7008,N_6551,N_6806);
nand U7009 (N_7009,N_6585,N_6743);
nor U7010 (N_7010,N_6632,N_6984);
nor U7011 (N_7011,N_6883,N_6800);
nor U7012 (N_7012,N_6652,N_6812);
nand U7013 (N_7013,N_6913,N_6974);
nor U7014 (N_7014,N_6726,N_6706);
nor U7015 (N_7015,N_6682,N_6510);
or U7016 (N_7016,N_6745,N_6868);
or U7017 (N_7017,N_6829,N_6857);
or U7018 (N_7018,N_6920,N_6938);
xnor U7019 (N_7019,N_6986,N_6909);
and U7020 (N_7020,N_6634,N_6543);
or U7021 (N_7021,N_6639,N_6659);
nor U7022 (N_7022,N_6539,N_6552);
or U7023 (N_7023,N_6766,N_6860);
nand U7024 (N_7024,N_6589,N_6504);
nand U7025 (N_7025,N_6571,N_6606);
xor U7026 (N_7026,N_6635,N_6624);
nor U7027 (N_7027,N_6574,N_6980);
nor U7028 (N_7028,N_6849,N_6712);
and U7029 (N_7029,N_6626,N_6942);
and U7030 (N_7030,N_6814,N_6691);
nand U7031 (N_7031,N_6828,N_6977);
and U7032 (N_7032,N_6713,N_6961);
and U7033 (N_7033,N_6981,N_6962);
nor U7034 (N_7034,N_6636,N_6765);
xnor U7035 (N_7035,N_6605,N_6525);
or U7036 (N_7036,N_6776,N_6502);
nor U7037 (N_7037,N_6614,N_6867);
nand U7038 (N_7038,N_6902,N_6536);
nand U7039 (N_7039,N_6566,N_6546);
or U7040 (N_7040,N_6751,N_6959);
xor U7041 (N_7041,N_6826,N_6593);
nor U7042 (N_7042,N_6988,N_6903);
nor U7043 (N_7043,N_6523,N_6676);
or U7044 (N_7044,N_6785,N_6956);
and U7045 (N_7045,N_6792,N_6541);
nand U7046 (N_7046,N_6690,N_6607);
nor U7047 (N_7047,N_6565,N_6651);
nor U7048 (N_7048,N_6907,N_6805);
nor U7049 (N_7049,N_6821,N_6963);
or U7050 (N_7050,N_6665,N_6573);
nor U7051 (N_7051,N_6612,N_6945);
or U7052 (N_7052,N_6952,N_6819);
or U7053 (N_7053,N_6707,N_6608);
and U7054 (N_7054,N_6865,N_6784);
nand U7055 (N_7055,N_6811,N_6699);
or U7056 (N_7056,N_6719,N_6710);
or U7057 (N_7057,N_6610,N_6660);
xnor U7058 (N_7058,N_6555,N_6617);
or U7059 (N_7059,N_6640,N_6897);
or U7060 (N_7060,N_6725,N_6599);
nor U7061 (N_7061,N_6904,N_6797);
nand U7062 (N_7062,N_6874,N_6717);
nor U7063 (N_7063,N_6545,N_6732);
and U7064 (N_7064,N_6804,N_6581);
or U7065 (N_7065,N_6519,N_6944);
xor U7066 (N_7066,N_6683,N_6680);
nand U7067 (N_7067,N_6601,N_6994);
nand U7068 (N_7068,N_6684,N_6861);
or U7069 (N_7069,N_6919,N_6816);
nand U7070 (N_7070,N_6677,N_6955);
nand U7071 (N_7071,N_6924,N_6521);
or U7072 (N_7072,N_6838,N_6538);
xnor U7073 (N_7073,N_6524,N_6841);
nand U7074 (N_7074,N_6746,N_6978);
nor U7075 (N_7075,N_6522,N_6619);
or U7076 (N_7076,N_6675,N_6846);
or U7077 (N_7077,N_6548,N_6761);
nor U7078 (N_7078,N_6901,N_6997);
nor U7079 (N_7079,N_6623,N_6936);
nor U7080 (N_7080,N_6900,N_6852);
xnor U7081 (N_7081,N_6759,N_6879);
or U7082 (N_7082,N_6937,N_6508);
xnor U7083 (N_7083,N_6535,N_6720);
and U7084 (N_7084,N_6989,N_6686);
xnor U7085 (N_7085,N_6899,N_6576);
nand U7086 (N_7086,N_6943,N_6629);
nor U7087 (N_7087,N_6558,N_6987);
and U7088 (N_7088,N_6983,N_6832);
and U7089 (N_7089,N_6970,N_6912);
nand U7090 (N_7090,N_6922,N_6733);
or U7091 (N_7091,N_6685,N_6796);
or U7092 (N_7092,N_6995,N_6625);
nand U7093 (N_7093,N_6637,N_6633);
nand U7094 (N_7094,N_6544,N_6622);
and U7095 (N_7095,N_6954,N_6889);
or U7096 (N_7096,N_6808,N_6768);
and U7097 (N_7097,N_6647,N_6895);
or U7098 (N_7098,N_6697,N_6668);
nand U7099 (N_7099,N_6649,N_6905);
and U7100 (N_7100,N_6918,N_6611);
xor U7101 (N_7101,N_6564,N_6722);
or U7102 (N_7102,N_6616,N_6577);
or U7103 (N_7103,N_6859,N_6966);
xnor U7104 (N_7104,N_6597,N_6596);
nor U7105 (N_7105,N_6563,N_6711);
nand U7106 (N_7106,N_6716,N_6778);
and U7107 (N_7107,N_6529,N_6864);
or U7108 (N_7108,N_6654,N_6964);
xnor U7109 (N_7109,N_6603,N_6853);
or U7110 (N_7110,N_6643,N_6579);
and U7111 (N_7111,N_6917,N_6848);
xor U7112 (N_7112,N_6949,N_6658);
xnor U7113 (N_7113,N_6872,N_6906);
and U7114 (N_7114,N_6769,N_6505);
or U7115 (N_7115,N_6650,N_6542);
and U7116 (N_7116,N_6641,N_6547);
or U7117 (N_7117,N_6709,N_6582);
or U7118 (N_7118,N_6878,N_6774);
nor U7119 (N_7119,N_6910,N_6855);
and U7120 (N_7120,N_6951,N_6674);
or U7121 (N_7121,N_6893,N_6742);
nand U7122 (N_7122,N_6817,N_6818);
nand U7123 (N_7123,N_6584,N_6721);
xor U7124 (N_7124,N_6991,N_6935);
xor U7125 (N_7125,N_6530,N_6513);
xnor U7126 (N_7126,N_6661,N_6644);
or U7127 (N_7127,N_6932,N_6933);
nand U7128 (N_7128,N_6518,N_6927);
nand U7129 (N_7129,N_6866,N_6870);
and U7130 (N_7130,N_6876,N_6550);
xnor U7131 (N_7131,N_6727,N_6734);
nor U7132 (N_7132,N_6940,N_6723);
nor U7133 (N_7133,N_6672,N_6982);
nor U7134 (N_7134,N_6820,N_6568);
xnor U7135 (N_7135,N_6561,N_6602);
xnor U7136 (N_7136,N_6556,N_6786);
xor U7137 (N_7137,N_6559,N_6527);
or U7138 (N_7138,N_6688,N_6923);
nand U7139 (N_7139,N_6515,N_6512);
or U7140 (N_7140,N_6873,N_6528);
xor U7141 (N_7141,N_6557,N_6787);
nand U7142 (N_7142,N_6948,N_6835);
or U7143 (N_7143,N_6825,N_6687);
and U7144 (N_7144,N_6503,N_6664);
nor U7145 (N_7145,N_6730,N_6834);
nand U7146 (N_7146,N_6837,N_6507);
and U7147 (N_7147,N_6526,N_6740);
nor U7148 (N_7148,N_6724,N_6969);
xnor U7149 (N_7149,N_6695,N_6780);
nand U7150 (N_7150,N_6705,N_6985);
nand U7151 (N_7151,N_6506,N_6757);
and U7152 (N_7152,N_6516,N_6531);
xnor U7153 (N_7153,N_6803,N_6567);
and U7154 (N_7154,N_6795,N_6754);
or U7155 (N_7155,N_6752,N_6813);
xnor U7156 (N_7156,N_6591,N_6793);
or U7157 (N_7157,N_6517,N_6560);
nor U7158 (N_7158,N_6815,N_6854);
or U7159 (N_7159,N_6908,N_6670);
and U7160 (N_7160,N_6898,N_6600);
or U7161 (N_7161,N_6748,N_6615);
nand U7162 (N_7162,N_6881,N_6655);
xnor U7163 (N_7163,N_6823,N_6931);
xnor U7164 (N_7164,N_6772,N_6968);
and U7165 (N_7165,N_6592,N_6679);
nand U7166 (N_7166,N_6511,N_6996);
xor U7167 (N_7167,N_6807,N_6590);
nor U7168 (N_7168,N_6880,N_6669);
and U7169 (N_7169,N_6738,N_6877);
nor U7170 (N_7170,N_6758,N_6762);
or U7171 (N_7171,N_6775,N_6501);
nor U7172 (N_7172,N_6946,N_6666);
nand U7173 (N_7173,N_6767,N_6892);
nand U7174 (N_7174,N_6790,N_6788);
xor U7175 (N_7175,N_6520,N_6554);
xnor U7176 (N_7176,N_6930,N_6646);
or U7177 (N_7177,N_6509,N_6953);
nand U7178 (N_7178,N_6653,N_6833);
or U7179 (N_7179,N_6929,N_6830);
xor U7180 (N_7180,N_6972,N_6779);
and U7181 (N_7181,N_6575,N_6894);
nor U7182 (N_7182,N_6532,N_6851);
nand U7183 (N_7183,N_6871,N_6747);
nor U7184 (N_7184,N_6896,N_6628);
nor U7185 (N_7185,N_6744,N_6802);
nand U7186 (N_7186,N_6588,N_6965);
nand U7187 (N_7187,N_6609,N_6753);
or U7188 (N_7188,N_6973,N_6856);
nor U7189 (N_7189,N_6831,N_6809);
nand U7190 (N_7190,N_6760,N_6979);
xor U7191 (N_7191,N_6960,N_6843);
nor U7192 (N_7192,N_6549,N_6990);
and U7193 (N_7193,N_6975,N_6801);
xnor U7194 (N_7194,N_6750,N_6941);
xnor U7195 (N_7195,N_6735,N_6578);
and U7196 (N_7196,N_6971,N_6657);
nand U7197 (N_7197,N_6704,N_6645);
xnor U7198 (N_7198,N_6925,N_6613);
nand U7199 (N_7199,N_6844,N_6822);
and U7200 (N_7200,N_6736,N_6749);
or U7201 (N_7201,N_6708,N_6671);
xor U7202 (N_7202,N_6914,N_6667);
xor U7203 (N_7203,N_6621,N_6798);
nand U7204 (N_7204,N_6842,N_6701);
nor U7205 (N_7205,N_6598,N_6882);
or U7206 (N_7206,N_6537,N_6715);
xor U7207 (N_7207,N_6572,N_6500);
nor U7208 (N_7208,N_6638,N_6540);
xor U7209 (N_7209,N_6794,N_6698);
and U7210 (N_7210,N_6692,N_6999);
and U7211 (N_7211,N_6553,N_6694);
and U7212 (N_7212,N_6890,N_6570);
and U7213 (N_7213,N_6998,N_6939);
or U7214 (N_7214,N_6958,N_6702);
xor U7215 (N_7215,N_6739,N_6847);
or U7216 (N_7216,N_6586,N_6915);
and U7217 (N_7217,N_6662,N_6514);
or U7218 (N_7218,N_6718,N_6703);
nand U7219 (N_7219,N_6836,N_6869);
nor U7220 (N_7220,N_6934,N_6885);
or U7221 (N_7221,N_6693,N_6569);
or U7222 (N_7222,N_6993,N_6858);
or U7223 (N_7223,N_6594,N_6630);
and U7224 (N_7224,N_6642,N_6700);
and U7225 (N_7225,N_6604,N_6620);
xnor U7226 (N_7226,N_6755,N_6886);
or U7227 (N_7227,N_6618,N_6533);
and U7228 (N_7228,N_6799,N_6810);
and U7229 (N_7229,N_6782,N_6731);
nand U7230 (N_7230,N_6773,N_6863);
nand U7231 (N_7231,N_6875,N_6926);
and U7232 (N_7232,N_6928,N_6648);
nand U7233 (N_7233,N_6763,N_6947);
nor U7234 (N_7234,N_6627,N_6756);
nor U7235 (N_7235,N_6587,N_6770);
nand U7236 (N_7236,N_6741,N_6534);
nand U7237 (N_7237,N_6824,N_6976);
and U7238 (N_7238,N_6791,N_6921);
xor U7239 (N_7239,N_6916,N_6789);
and U7240 (N_7240,N_6992,N_6681);
xnor U7241 (N_7241,N_6850,N_6583);
xor U7242 (N_7242,N_6737,N_6781);
xor U7243 (N_7243,N_6862,N_6839);
xor U7244 (N_7244,N_6631,N_6729);
or U7245 (N_7245,N_6827,N_6678);
and U7246 (N_7246,N_6656,N_6580);
and U7247 (N_7247,N_6967,N_6696);
or U7248 (N_7248,N_6783,N_6595);
or U7249 (N_7249,N_6888,N_6689);
nor U7250 (N_7250,N_6738,N_6933);
and U7251 (N_7251,N_6801,N_6940);
nor U7252 (N_7252,N_6859,N_6834);
and U7253 (N_7253,N_6975,N_6581);
nor U7254 (N_7254,N_6803,N_6914);
nand U7255 (N_7255,N_6810,N_6798);
xnor U7256 (N_7256,N_6783,N_6990);
nand U7257 (N_7257,N_6593,N_6810);
xnor U7258 (N_7258,N_6824,N_6512);
xor U7259 (N_7259,N_6720,N_6875);
nor U7260 (N_7260,N_6787,N_6865);
or U7261 (N_7261,N_6655,N_6983);
xnor U7262 (N_7262,N_6909,N_6906);
and U7263 (N_7263,N_6738,N_6531);
nor U7264 (N_7264,N_6637,N_6823);
and U7265 (N_7265,N_6593,N_6510);
nor U7266 (N_7266,N_6619,N_6881);
or U7267 (N_7267,N_6846,N_6585);
xor U7268 (N_7268,N_6921,N_6702);
or U7269 (N_7269,N_6573,N_6599);
and U7270 (N_7270,N_6618,N_6693);
nor U7271 (N_7271,N_6951,N_6513);
or U7272 (N_7272,N_6666,N_6753);
nor U7273 (N_7273,N_6974,N_6630);
xor U7274 (N_7274,N_6994,N_6612);
and U7275 (N_7275,N_6513,N_6611);
xnor U7276 (N_7276,N_6581,N_6772);
or U7277 (N_7277,N_6602,N_6542);
and U7278 (N_7278,N_6792,N_6812);
and U7279 (N_7279,N_6899,N_6807);
nor U7280 (N_7280,N_6511,N_6745);
or U7281 (N_7281,N_6900,N_6592);
and U7282 (N_7282,N_6826,N_6715);
nand U7283 (N_7283,N_6726,N_6989);
xor U7284 (N_7284,N_6715,N_6594);
xnor U7285 (N_7285,N_6509,N_6967);
nor U7286 (N_7286,N_6586,N_6941);
nor U7287 (N_7287,N_6729,N_6951);
nor U7288 (N_7288,N_6973,N_6852);
xnor U7289 (N_7289,N_6686,N_6815);
nor U7290 (N_7290,N_6597,N_6594);
or U7291 (N_7291,N_6703,N_6802);
nor U7292 (N_7292,N_6742,N_6871);
or U7293 (N_7293,N_6661,N_6795);
nor U7294 (N_7294,N_6740,N_6635);
and U7295 (N_7295,N_6844,N_6980);
or U7296 (N_7296,N_6947,N_6748);
xnor U7297 (N_7297,N_6510,N_6922);
or U7298 (N_7298,N_6775,N_6709);
xor U7299 (N_7299,N_6540,N_6679);
or U7300 (N_7300,N_6721,N_6874);
nor U7301 (N_7301,N_6946,N_6957);
nand U7302 (N_7302,N_6829,N_6656);
and U7303 (N_7303,N_6860,N_6594);
and U7304 (N_7304,N_6997,N_6613);
or U7305 (N_7305,N_6632,N_6955);
xnor U7306 (N_7306,N_6845,N_6960);
or U7307 (N_7307,N_6714,N_6796);
or U7308 (N_7308,N_6708,N_6612);
nand U7309 (N_7309,N_6907,N_6770);
nor U7310 (N_7310,N_6685,N_6986);
or U7311 (N_7311,N_6587,N_6544);
nor U7312 (N_7312,N_6892,N_6645);
and U7313 (N_7313,N_6659,N_6505);
nand U7314 (N_7314,N_6784,N_6590);
xor U7315 (N_7315,N_6733,N_6874);
nor U7316 (N_7316,N_6515,N_6706);
nor U7317 (N_7317,N_6895,N_6636);
nand U7318 (N_7318,N_6556,N_6903);
nor U7319 (N_7319,N_6503,N_6533);
or U7320 (N_7320,N_6817,N_6838);
xnor U7321 (N_7321,N_6988,N_6748);
xor U7322 (N_7322,N_6992,N_6901);
xor U7323 (N_7323,N_6628,N_6686);
or U7324 (N_7324,N_6622,N_6572);
nand U7325 (N_7325,N_6992,N_6791);
xnor U7326 (N_7326,N_6926,N_6794);
nor U7327 (N_7327,N_6872,N_6576);
nand U7328 (N_7328,N_6692,N_6775);
nor U7329 (N_7329,N_6885,N_6971);
or U7330 (N_7330,N_6608,N_6706);
nand U7331 (N_7331,N_6735,N_6877);
and U7332 (N_7332,N_6875,N_6886);
xor U7333 (N_7333,N_6777,N_6990);
and U7334 (N_7334,N_6689,N_6566);
xnor U7335 (N_7335,N_6604,N_6539);
xor U7336 (N_7336,N_6661,N_6638);
or U7337 (N_7337,N_6980,N_6810);
or U7338 (N_7338,N_6705,N_6543);
nand U7339 (N_7339,N_6661,N_6681);
xor U7340 (N_7340,N_6558,N_6813);
nand U7341 (N_7341,N_6601,N_6623);
nand U7342 (N_7342,N_6502,N_6547);
nor U7343 (N_7343,N_6804,N_6873);
and U7344 (N_7344,N_6807,N_6950);
nand U7345 (N_7345,N_6548,N_6914);
and U7346 (N_7346,N_6751,N_6903);
and U7347 (N_7347,N_6968,N_6733);
nand U7348 (N_7348,N_6571,N_6560);
xnor U7349 (N_7349,N_6810,N_6884);
xor U7350 (N_7350,N_6862,N_6981);
nand U7351 (N_7351,N_6672,N_6912);
nor U7352 (N_7352,N_6540,N_6926);
nor U7353 (N_7353,N_6999,N_6816);
nor U7354 (N_7354,N_6575,N_6979);
or U7355 (N_7355,N_6622,N_6968);
nor U7356 (N_7356,N_6637,N_6735);
xor U7357 (N_7357,N_6773,N_6594);
nand U7358 (N_7358,N_6586,N_6796);
and U7359 (N_7359,N_6642,N_6817);
xor U7360 (N_7360,N_6769,N_6516);
nand U7361 (N_7361,N_6777,N_6859);
and U7362 (N_7362,N_6984,N_6960);
xor U7363 (N_7363,N_6573,N_6862);
nand U7364 (N_7364,N_6874,N_6563);
nor U7365 (N_7365,N_6789,N_6682);
nor U7366 (N_7366,N_6608,N_6571);
xnor U7367 (N_7367,N_6626,N_6559);
nand U7368 (N_7368,N_6624,N_6633);
and U7369 (N_7369,N_6783,N_6848);
nand U7370 (N_7370,N_6561,N_6926);
nand U7371 (N_7371,N_6538,N_6731);
xnor U7372 (N_7372,N_6974,N_6560);
and U7373 (N_7373,N_6908,N_6593);
xnor U7374 (N_7374,N_6936,N_6842);
or U7375 (N_7375,N_6886,N_6591);
xor U7376 (N_7376,N_6541,N_6928);
nand U7377 (N_7377,N_6785,N_6514);
nor U7378 (N_7378,N_6534,N_6756);
nor U7379 (N_7379,N_6771,N_6823);
nor U7380 (N_7380,N_6973,N_6859);
xnor U7381 (N_7381,N_6571,N_6674);
or U7382 (N_7382,N_6827,N_6996);
nand U7383 (N_7383,N_6927,N_6935);
nand U7384 (N_7384,N_6698,N_6781);
nor U7385 (N_7385,N_6711,N_6680);
or U7386 (N_7386,N_6954,N_6593);
nor U7387 (N_7387,N_6568,N_6572);
xor U7388 (N_7388,N_6698,N_6905);
nor U7389 (N_7389,N_6923,N_6623);
or U7390 (N_7390,N_6554,N_6813);
and U7391 (N_7391,N_6529,N_6829);
xnor U7392 (N_7392,N_6552,N_6692);
or U7393 (N_7393,N_6811,N_6586);
nor U7394 (N_7394,N_6623,N_6938);
nand U7395 (N_7395,N_6512,N_6906);
or U7396 (N_7396,N_6542,N_6931);
nand U7397 (N_7397,N_6985,N_6517);
or U7398 (N_7398,N_6506,N_6911);
nor U7399 (N_7399,N_6990,N_6668);
xnor U7400 (N_7400,N_6897,N_6656);
xnor U7401 (N_7401,N_6629,N_6901);
nand U7402 (N_7402,N_6964,N_6740);
xor U7403 (N_7403,N_6841,N_6949);
and U7404 (N_7404,N_6700,N_6777);
xor U7405 (N_7405,N_6880,N_6918);
xor U7406 (N_7406,N_6594,N_6593);
nand U7407 (N_7407,N_6706,N_6883);
and U7408 (N_7408,N_6974,N_6789);
xnor U7409 (N_7409,N_6690,N_6746);
and U7410 (N_7410,N_6975,N_6619);
nor U7411 (N_7411,N_6883,N_6607);
or U7412 (N_7412,N_6724,N_6594);
nor U7413 (N_7413,N_6733,N_6666);
and U7414 (N_7414,N_6760,N_6632);
or U7415 (N_7415,N_6803,N_6535);
nor U7416 (N_7416,N_6992,N_6787);
nor U7417 (N_7417,N_6730,N_6573);
nand U7418 (N_7418,N_6874,N_6734);
and U7419 (N_7419,N_6685,N_6522);
nor U7420 (N_7420,N_6751,N_6892);
nor U7421 (N_7421,N_6884,N_6502);
or U7422 (N_7422,N_6717,N_6579);
nor U7423 (N_7423,N_6735,N_6640);
or U7424 (N_7424,N_6828,N_6785);
or U7425 (N_7425,N_6692,N_6780);
nor U7426 (N_7426,N_6822,N_6736);
and U7427 (N_7427,N_6872,N_6811);
nand U7428 (N_7428,N_6794,N_6768);
and U7429 (N_7429,N_6687,N_6971);
and U7430 (N_7430,N_6843,N_6920);
and U7431 (N_7431,N_6838,N_6638);
and U7432 (N_7432,N_6746,N_6600);
or U7433 (N_7433,N_6976,N_6971);
or U7434 (N_7434,N_6534,N_6890);
or U7435 (N_7435,N_6959,N_6893);
and U7436 (N_7436,N_6616,N_6891);
nand U7437 (N_7437,N_6906,N_6875);
xnor U7438 (N_7438,N_6767,N_6813);
or U7439 (N_7439,N_6584,N_6914);
nand U7440 (N_7440,N_6627,N_6739);
or U7441 (N_7441,N_6868,N_6552);
nor U7442 (N_7442,N_6624,N_6843);
and U7443 (N_7443,N_6529,N_6750);
nand U7444 (N_7444,N_6927,N_6530);
xnor U7445 (N_7445,N_6971,N_6839);
xor U7446 (N_7446,N_6796,N_6907);
xor U7447 (N_7447,N_6628,N_6536);
and U7448 (N_7448,N_6887,N_6792);
and U7449 (N_7449,N_6806,N_6612);
nand U7450 (N_7450,N_6776,N_6894);
and U7451 (N_7451,N_6880,N_6746);
nand U7452 (N_7452,N_6549,N_6694);
nor U7453 (N_7453,N_6632,N_6977);
nand U7454 (N_7454,N_6942,N_6848);
or U7455 (N_7455,N_6607,N_6507);
nor U7456 (N_7456,N_6850,N_6998);
and U7457 (N_7457,N_6967,N_6813);
xor U7458 (N_7458,N_6978,N_6735);
nor U7459 (N_7459,N_6588,N_6743);
xnor U7460 (N_7460,N_6701,N_6599);
or U7461 (N_7461,N_6931,N_6650);
xnor U7462 (N_7462,N_6606,N_6778);
nand U7463 (N_7463,N_6532,N_6742);
nor U7464 (N_7464,N_6855,N_6604);
nor U7465 (N_7465,N_6922,N_6653);
nand U7466 (N_7466,N_6609,N_6601);
or U7467 (N_7467,N_6696,N_6538);
nand U7468 (N_7468,N_6770,N_6850);
xor U7469 (N_7469,N_6764,N_6610);
nand U7470 (N_7470,N_6540,N_6740);
xor U7471 (N_7471,N_6510,N_6853);
nor U7472 (N_7472,N_6559,N_6647);
nand U7473 (N_7473,N_6706,N_6771);
and U7474 (N_7474,N_6921,N_6567);
nand U7475 (N_7475,N_6925,N_6696);
nand U7476 (N_7476,N_6827,N_6893);
xnor U7477 (N_7477,N_6649,N_6828);
and U7478 (N_7478,N_6867,N_6703);
nor U7479 (N_7479,N_6618,N_6822);
nor U7480 (N_7480,N_6532,N_6798);
nand U7481 (N_7481,N_6776,N_6969);
and U7482 (N_7482,N_6576,N_6768);
xnor U7483 (N_7483,N_6543,N_6926);
xor U7484 (N_7484,N_6666,N_6723);
xnor U7485 (N_7485,N_6995,N_6721);
nand U7486 (N_7486,N_6526,N_6986);
nand U7487 (N_7487,N_6753,N_6566);
nand U7488 (N_7488,N_6944,N_6635);
nor U7489 (N_7489,N_6786,N_6803);
xnor U7490 (N_7490,N_6935,N_6784);
nor U7491 (N_7491,N_6630,N_6694);
and U7492 (N_7492,N_6955,N_6813);
nor U7493 (N_7493,N_6686,N_6978);
and U7494 (N_7494,N_6521,N_6716);
nor U7495 (N_7495,N_6702,N_6913);
xnor U7496 (N_7496,N_6713,N_6633);
or U7497 (N_7497,N_6871,N_6971);
xor U7498 (N_7498,N_6846,N_6571);
nand U7499 (N_7499,N_6688,N_6686);
xnor U7500 (N_7500,N_7462,N_7340);
and U7501 (N_7501,N_7028,N_7367);
and U7502 (N_7502,N_7199,N_7143);
xor U7503 (N_7503,N_7147,N_7344);
and U7504 (N_7504,N_7457,N_7097);
and U7505 (N_7505,N_7451,N_7403);
nand U7506 (N_7506,N_7379,N_7357);
xnor U7507 (N_7507,N_7453,N_7419);
nand U7508 (N_7508,N_7378,N_7196);
and U7509 (N_7509,N_7156,N_7209);
and U7510 (N_7510,N_7105,N_7048);
nor U7511 (N_7511,N_7360,N_7382);
or U7512 (N_7512,N_7253,N_7050);
nand U7513 (N_7513,N_7337,N_7391);
nor U7514 (N_7514,N_7164,N_7091);
nand U7515 (N_7515,N_7016,N_7118);
nor U7516 (N_7516,N_7020,N_7065);
nand U7517 (N_7517,N_7287,N_7151);
and U7518 (N_7518,N_7079,N_7015);
and U7519 (N_7519,N_7288,N_7459);
or U7520 (N_7520,N_7131,N_7333);
xnor U7521 (N_7521,N_7042,N_7186);
and U7522 (N_7522,N_7302,N_7141);
nor U7523 (N_7523,N_7178,N_7145);
or U7524 (N_7524,N_7251,N_7124);
or U7525 (N_7525,N_7386,N_7161);
or U7526 (N_7526,N_7283,N_7359);
xor U7527 (N_7527,N_7301,N_7284);
and U7528 (N_7528,N_7444,N_7117);
xor U7529 (N_7529,N_7137,N_7371);
xor U7530 (N_7530,N_7032,N_7109);
nor U7531 (N_7531,N_7342,N_7235);
nand U7532 (N_7532,N_7049,N_7358);
and U7533 (N_7533,N_7361,N_7431);
or U7534 (N_7534,N_7122,N_7428);
or U7535 (N_7535,N_7089,N_7465);
xor U7536 (N_7536,N_7335,N_7121);
nor U7537 (N_7537,N_7472,N_7076);
xor U7538 (N_7538,N_7477,N_7188);
xnor U7539 (N_7539,N_7277,N_7321);
or U7540 (N_7540,N_7018,N_7353);
or U7541 (N_7541,N_7167,N_7255);
and U7542 (N_7542,N_7006,N_7415);
and U7543 (N_7543,N_7139,N_7410);
and U7544 (N_7544,N_7326,N_7179);
or U7545 (N_7545,N_7427,N_7440);
and U7546 (N_7546,N_7423,N_7345);
nand U7547 (N_7547,N_7036,N_7112);
nor U7548 (N_7548,N_7120,N_7000);
nand U7549 (N_7549,N_7177,N_7250);
or U7550 (N_7550,N_7256,N_7327);
and U7551 (N_7551,N_7046,N_7259);
nor U7552 (N_7552,N_7313,N_7456);
xnor U7553 (N_7553,N_7454,N_7364);
and U7554 (N_7554,N_7395,N_7434);
xor U7555 (N_7555,N_7289,N_7486);
nor U7556 (N_7556,N_7396,N_7102);
nor U7557 (N_7557,N_7045,N_7115);
nor U7558 (N_7558,N_7452,N_7494);
or U7559 (N_7559,N_7374,N_7349);
nand U7560 (N_7560,N_7215,N_7392);
nor U7561 (N_7561,N_7170,N_7401);
nand U7562 (N_7562,N_7474,N_7169);
xor U7563 (N_7563,N_7338,N_7491);
or U7564 (N_7564,N_7263,N_7192);
and U7565 (N_7565,N_7060,N_7153);
and U7566 (N_7566,N_7274,N_7101);
nand U7567 (N_7567,N_7308,N_7087);
nand U7568 (N_7568,N_7126,N_7347);
nand U7569 (N_7569,N_7009,N_7174);
and U7570 (N_7570,N_7365,N_7325);
nor U7571 (N_7571,N_7267,N_7224);
or U7572 (N_7572,N_7280,N_7372);
and U7573 (N_7573,N_7125,N_7258);
nand U7574 (N_7574,N_7322,N_7037);
xnor U7575 (N_7575,N_7129,N_7245);
xor U7576 (N_7576,N_7438,N_7080);
nand U7577 (N_7577,N_7019,N_7231);
xor U7578 (N_7578,N_7265,N_7292);
and U7579 (N_7579,N_7166,N_7216);
nor U7580 (N_7580,N_7138,N_7411);
and U7581 (N_7581,N_7466,N_7248);
nand U7582 (N_7582,N_7189,N_7148);
nor U7583 (N_7583,N_7064,N_7158);
xor U7584 (N_7584,N_7082,N_7232);
and U7585 (N_7585,N_7246,N_7044);
or U7586 (N_7586,N_7356,N_7098);
nand U7587 (N_7587,N_7095,N_7233);
xnor U7588 (N_7588,N_7296,N_7268);
nor U7589 (N_7589,N_7104,N_7424);
nor U7590 (N_7590,N_7221,N_7172);
or U7591 (N_7591,N_7084,N_7257);
nor U7592 (N_7592,N_7468,N_7385);
or U7593 (N_7593,N_7014,N_7146);
nand U7594 (N_7594,N_7414,N_7464);
and U7595 (N_7595,N_7489,N_7239);
and U7596 (N_7596,N_7487,N_7348);
xor U7597 (N_7597,N_7165,N_7299);
nand U7598 (N_7598,N_7476,N_7213);
nand U7599 (N_7599,N_7133,N_7157);
xor U7600 (N_7600,N_7181,N_7418);
xor U7601 (N_7601,N_7404,N_7484);
nand U7602 (N_7602,N_7069,N_7416);
and U7603 (N_7603,N_7314,N_7425);
or U7604 (N_7604,N_7407,N_7282);
or U7605 (N_7605,N_7040,N_7219);
nor U7606 (N_7606,N_7171,N_7134);
xor U7607 (N_7607,N_7220,N_7073);
and U7608 (N_7608,N_7390,N_7470);
xor U7609 (N_7609,N_7305,N_7226);
nand U7610 (N_7610,N_7460,N_7066);
nand U7611 (N_7611,N_7446,N_7234);
nand U7612 (N_7612,N_7497,N_7002);
xor U7613 (N_7613,N_7455,N_7200);
or U7614 (N_7614,N_7394,N_7445);
nor U7615 (N_7615,N_7315,N_7400);
nand U7616 (N_7616,N_7490,N_7180);
nand U7617 (N_7617,N_7218,N_7227);
nor U7618 (N_7618,N_7140,N_7270);
nor U7619 (N_7619,N_7247,N_7225);
nor U7620 (N_7620,N_7208,N_7387);
nor U7621 (N_7621,N_7207,N_7242);
xor U7622 (N_7622,N_7317,N_7100);
nand U7623 (N_7623,N_7421,N_7041);
nor U7624 (N_7624,N_7437,N_7482);
or U7625 (N_7625,N_7197,N_7481);
xor U7626 (N_7626,N_7323,N_7116);
nor U7627 (N_7627,N_7350,N_7492);
nand U7628 (N_7628,N_7029,N_7043);
nand U7629 (N_7629,N_7362,N_7306);
nand U7630 (N_7630,N_7191,N_7123);
xnor U7631 (N_7631,N_7311,N_7290);
and U7632 (N_7632,N_7293,N_7261);
xnor U7633 (N_7633,N_7183,N_7389);
and U7634 (N_7634,N_7328,N_7099);
xor U7635 (N_7635,N_7004,N_7271);
nand U7636 (N_7636,N_7294,N_7399);
xnor U7637 (N_7637,N_7011,N_7343);
nor U7638 (N_7638,N_7047,N_7355);
nand U7639 (N_7639,N_7475,N_7429);
xnor U7640 (N_7640,N_7030,N_7149);
and U7641 (N_7641,N_7442,N_7316);
or U7642 (N_7642,N_7262,N_7034);
or U7643 (N_7643,N_7144,N_7229);
and U7644 (N_7644,N_7275,N_7154);
nand U7645 (N_7645,N_7393,N_7071);
or U7646 (N_7646,N_7458,N_7072);
and U7647 (N_7647,N_7111,N_7329);
or U7648 (N_7648,N_7202,N_7269);
or U7649 (N_7649,N_7254,N_7128);
and U7650 (N_7650,N_7312,N_7383);
xnor U7651 (N_7651,N_7057,N_7230);
nand U7652 (N_7652,N_7496,N_7398);
and U7653 (N_7653,N_7384,N_7436);
or U7654 (N_7654,N_7334,N_7435);
nand U7655 (N_7655,N_7408,N_7412);
and U7656 (N_7656,N_7339,N_7211);
or U7657 (N_7657,N_7086,N_7067);
xnor U7658 (N_7658,N_7273,N_7388);
nand U7659 (N_7659,N_7168,N_7204);
or U7660 (N_7660,N_7278,N_7212);
and U7661 (N_7661,N_7023,N_7363);
and U7662 (N_7662,N_7110,N_7495);
and U7663 (N_7663,N_7184,N_7187);
or U7664 (N_7664,N_7370,N_7078);
and U7665 (N_7665,N_7055,N_7176);
xnor U7666 (N_7666,N_7113,N_7285);
and U7667 (N_7667,N_7038,N_7093);
nand U7668 (N_7668,N_7480,N_7001);
nand U7669 (N_7669,N_7381,N_7075);
nor U7670 (N_7670,N_7448,N_7264);
nand U7671 (N_7671,N_7203,N_7155);
or U7672 (N_7672,N_7304,N_7198);
and U7673 (N_7673,N_7332,N_7108);
and U7674 (N_7674,N_7193,N_7035);
nor U7675 (N_7675,N_7026,N_7324);
and U7676 (N_7676,N_7039,N_7479);
nand U7677 (N_7677,N_7373,N_7090);
nand U7678 (N_7678,N_7380,N_7003);
or U7679 (N_7679,N_7307,N_7222);
xor U7680 (N_7680,N_7114,N_7351);
or U7681 (N_7681,N_7053,N_7498);
nand U7682 (N_7682,N_7236,N_7163);
and U7683 (N_7683,N_7162,N_7135);
nor U7684 (N_7684,N_7150,N_7103);
nor U7685 (N_7685,N_7397,N_7286);
or U7686 (N_7686,N_7405,N_7266);
nor U7687 (N_7687,N_7441,N_7058);
or U7688 (N_7688,N_7318,N_7195);
nand U7689 (N_7689,N_7025,N_7031);
nor U7690 (N_7690,N_7008,N_7130);
and U7691 (N_7691,N_7005,N_7228);
nand U7692 (N_7692,N_7013,N_7022);
nand U7693 (N_7693,N_7402,N_7298);
nand U7694 (N_7694,N_7223,N_7422);
xor U7695 (N_7695,N_7488,N_7417);
xnor U7696 (N_7696,N_7303,N_7433);
or U7697 (N_7697,N_7142,N_7061);
nand U7698 (N_7698,N_7406,N_7377);
xnor U7699 (N_7699,N_7243,N_7300);
xnor U7700 (N_7700,N_7214,N_7450);
or U7701 (N_7701,N_7190,N_7136);
nand U7702 (N_7702,N_7182,N_7194);
xnor U7703 (N_7703,N_7106,N_7320);
xnor U7704 (N_7704,N_7483,N_7354);
nor U7705 (N_7705,N_7107,N_7375);
nand U7706 (N_7706,N_7443,N_7201);
xor U7707 (N_7707,N_7096,N_7063);
xnor U7708 (N_7708,N_7074,N_7068);
nor U7709 (N_7709,N_7185,N_7369);
nor U7710 (N_7710,N_7205,N_7092);
xnor U7711 (N_7711,N_7420,N_7432);
or U7712 (N_7712,N_7352,N_7083);
nor U7713 (N_7713,N_7341,N_7152);
xnor U7714 (N_7714,N_7309,N_7430);
and U7715 (N_7715,N_7281,N_7447);
and U7716 (N_7716,N_7252,N_7297);
and U7717 (N_7717,N_7160,N_7119);
and U7718 (N_7718,N_7279,N_7052);
xnor U7719 (N_7719,N_7336,N_7471);
xnor U7720 (N_7720,N_7276,N_7295);
nand U7721 (N_7721,N_7077,N_7244);
nand U7722 (N_7722,N_7033,N_7175);
and U7723 (N_7723,N_7473,N_7081);
xor U7724 (N_7724,N_7249,N_7469);
nand U7725 (N_7725,N_7493,N_7217);
nand U7726 (N_7726,N_7413,N_7062);
and U7727 (N_7727,N_7238,N_7059);
xnor U7728 (N_7728,N_7346,N_7310);
and U7729 (N_7729,N_7127,N_7007);
nor U7730 (N_7730,N_7159,N_7012);
or U7731 (N_7731,N_7499,N_7449);
or U7732 (N_7732,N_7467,N_7240);
nand U7733 (N_7733,N_7330,N_7010);
nor U7734 (N_7734,N_7027,N_7366);
and U7735 (N_7735,N_7024,N_7461);
nor U7736 (N_7736,N_7051,N_7260);
nor U7737 (N_7737,N_7070,N_7241);
nand U7738 (N_7738,N_7376,N_7463);
or U7739 (N_7739,N_7085,N_7017);
or U7740 (N_7740,N_7331,N_7132);
xor U7741 (N_7741,N_7291,N_7478);
nand U7742 (N_7742,N_7319,N_7054);
xor U7743 (N_7743,N_7210,N_7426);
or U7744 (N_7744,N_7368,N_7173);
nand U7745 (N_7745,N_7485,N_7237);
nand U7746 (N_7746,N_7206,N_7021);
or U7747 (N_7747,N_7056,N_7088);
and U7748 (N_7748,N_7439,N_7272);
nor U7749 (N_7749,N_7094,N_7409);
nand U7750 (N_7750,N_7496,N_7486);
or U7751 (N_7751,N_7162,N_7053);
nor U7752 (N_7752,N_7055,N_7243);
or U7753 (N_7753,N_7197,N_7031);
and U7754 (N_7754,N_7472,N_7197);
or U7755 (N_7755,N_7327,N_7148);
nand U7756 (N_7756,N_7434,N_7147);
and U7757 (N_7757,N_7407,N_7228);
or U7758 (N_7758,N_7040,N_7069);
and U7759 (N_7759,N_7493,N_7383);
nor U7760 (N_7760,N_7388,N_7260);
nand U7761 (N_7761,N_7431,N_7239);
nand U7762 (N_7762,N_7050,N_7103);
nand U7763 (N_7763,N_7489,N_7420);
nand U7764 (N_7764,N_7434,N_7384);
nor U7765 (N_7765,N_7310,N_7264);
xor U7766 (N_7766,N_7396,N_7389);
and U7767 (N_7767,N_7208,N_7359);
nand U7768 (N_7768,N_7073,N_7280);
xnor U7769 (N_7769,N_7493,N_7497);
or U7770 (N_7770,N_7415,N_7496);
nand U7771 (N_7771,N_7031,N_7178);
or U7772 (N_7772,N_7215,N_7135);
and U7773 (N_7773,N_7252,N_7198);
and U7774 (N_7774,N_7233,N_7231);
nor U7775 (N_7775,N_7181,N_7017);
xor U7776 (N_7776,N_7333,N_7286);
nand U7777 (N_7777,N_7012,N_7255);
xnor U7778 (N_7778,N_7337,N_7324);
and U7779 (N_7779,N_7404,N_7215);
nand U7780 (N_7780,N_7082,N_7364);
or U7781 (N_7781,N_7199,N_7127);
nand U7782 (N_7782,N_7004,N_7220);
and U7783 (N_7783,N_7010,N_7237);
nand U7784 (N_7784,N_7017,N_7016);
xor U7785 (N_7785,N_7257,N_7340);
nor U7786 (N_7786,N_7174,N_7031);
and U7787 (N_7787,N_7180,N_7006);
and U7788 (N_7788,N_7433,N_7278);
nor U7789 (N_7789,N_7215,N_7331);
and U7790 (N_7790,N_7323,N_7462);
xor U7791 (N_7791,N_7350,N_7222);
xor U7792 (N_7792,N_7306,N_7070);
xor U7793 (N_7793,N_7025,N_7392);
nor U7794 (N_7794,N_7092,N_7108);
nand U7795 (N_7795,N_7367,N_7168);
nor U7796 (N_7796,N_7018,N_7403);
xor U7797 (N_7797,N_7187,N_7350);
or U7798 (N_7798,N_7267,N_7043);
xor U7799 (N_7799,N_7121,N_7214);
and U7800 (N_7800,N_7181,N_7110);
nand U7801 (N_7801,N_7314,N_7378);
or U7802 (N_7802,N_7133,N_7334);
xor U7803 (N_7803,N_7285,N_7303);
or U7804 (N_7804,N_7150,N_7268);
nand U7805 (N_7805,N_7265,N_7228);
nor U7806 (N_7806,N_7120,N_7052);
xor U7807 (N_7807,N_7328,N_7483);
nor U7808 (N_7808,N_7454,N_7016);
nor U7809 (N_7809,N_7245,N_7439);
xnor U7810 (N_7810,N_7227,N_7471);
nor U7811 (N_7811,N_7270,N_7340);
nor U7812 (N_7812,N_7418,N_7177);
or U7813 (N_7813,N_7250,N_7005);
or U7814 (N_7814,N_7013,N_7338);
nand U7815 (N_7815,N_7135,N_7381);
or U7816 (N_7816,N_7428,N_7013);
xor U7817 (N_7817,N_7152,N_7391);
and U7818 (N_7818,N_7125,N_7223);
xor U7819 (N_7819,N_7173,N_7100);
and U7820 (N_7820,N_7161,N_7169);
xor U7821 (N_7821,N_7261,N_7282);
and U7822 (N_7822,N_7026,N_7430);
xor U7823 (N_7823,N_7143,N_7029);
or U7824 (N_7824,N_7218,N_7271);
nor U7825 (N_7825,N_7092,N_7400);
nand U7826 (N_7826,N_7093,N_7223);
and U7827 (N_7827,N_7142,N_7498);
nand U7828 (N_7828,N_7095,N_7112);
or U7829 (N_7829,N_7000,N_7240);
xnor U7830 (N_7830,N_7074,N_7017);
or U7831 (N_7831,N_7229,N_7078);
and U7832 (N_7832,N_7327,N_7168);
nor U7833 (N_7833,N_7412,N_7173);
nand U7834 (N_7834,N_7152,N_7161);
and U7835 (N_7835,N_7494,N_7128);
nor U7836 (N_7836,N_7194,N_7055);
nor U7837 (N_7837,N_7415,N_7088);
nor U7838 (N_7838,N_7266,N_7073);
nor U7839 (N_7839,N_7174,N_7476);
or U7840 (N_7840,N_7328,N_7408);
nand U7841 (N_7841,N_7288,N_7336);
xnor U7842 (N_7842,N_7346,N_7218);
and U7843 (N_7843,N_7440,N_7212);
and U7844 (N_7844,N_7305,N_7240);
nand U7845 (N_7845,N_7349,N_7036);
nor U7846 (N_7846,N_7045,N_7434);
or U7847 (N_7847,N_7099,N_7141);
nand U7848 (N_7848,N_7148,N_7325);
nor U7849 (N_7849,N_7199,N_7208);
xnor U7850 (N_7850,N_7195,N_7045);
or U7851 (N_7851,N_7005,N_7076);
nand U7852 (N_7852,N_7310,N_7384);
and U7853 (N_7853,N_7084,N_7072);
nand U7854 (N_7854,N_7378,N_7012);
or U7855 (N_7855,N_7466,N_7347);
nand U7856 (N_7856,N_7089,N_7483);
xnor U7857 (N_7857,N_7364,N_7303);
or U7858 (N_7858,N_7370,N_7053);
nand U7859 (N_7859,N_7078,N_7186);
nand U7860 (N_7860,N_7103,N_7015);
xor U7861 (N_7861,N_7494,N_7208);
or U7862 (N_7862,N_7328,N_7496);
and U7863 (N_7863,N_7267,N_7117);
nor U7864 (N_7864,N_7354,N_7468);
and U7865 (N_7865,N_7115,N_7211);
nand U7866 (N_7866,N_7132,N_7100);
or U7867 (N_7867,N_7065,N_7231);
nor U7868 (N_7868,N_7455,N_7394);
nor U7869 (N_7869,N_7360,N_7018);
or U7870 (N_7870,N_7092,N_7436);
or U7871 (N_7871,N_7490,N_7037);
or U7872 (N_7872,N_7475,N_7259);
and U7873 (N_7873,N_7217,N_7231);
or U7874 (N_7874,N_7155,N_7244);
and U7875 (N_7875,N_7160,N_7088);
nand U7876 (N_7876,N_7002,N_7232);
nor U7877 (N_7877,N_7201,N_7182);
and U7878 (N_7878,N_7479,N_7428);
nor U7879 (N_7879,N_7067,N_7031);
or U7880 (N_7880,N_7426,N_7171);
xor U7881 (N_7881,N_7073,N_7097);
nand U7882 (N_7882,N_7088,N_7325);
or U7883 (N_7883,N_7417,N_7319);
nor U7884 (N_7884,N_7449,N_7183);
nand U7885 (N_7885,N_7077,N_7116);
or U7886 (N_7886,N_7476,N_7289);
nand U7887 (N_7887,N_7283,N_7067);
nand U7888 (N_7888,N_7497,N_7443);
xnor U7889 (N_7889,N_7184,N_7179);
or U7890 (N_7890,N_7051,N_7249);
nand U7891 (N_7891,N_7488,N_7342);
nand U7892 (N_7892,N_7234,N_7217);
nand U7893 (N_7893,N_7327,N_7227);
or U7894 (N_7894,N_7039,N_7110);
nand U7895 (N_7895,N_7263,N_7246);
xnor U7896 (N_7896,N_7270,N_7215);
xor U7897 (N_7897,N_7021,N_7276);
nor U7898 (N_7898,N_7284,N_7247);
nor U7899 (N_7899,N_7453,N_7135);
nand U7900 (N_7900,N_7465,N_7272);
xnor U7901 (N_7901,N_7021,N_7425);
or U7902 (N_7902,N_7238,N_7434);
nor U7903 (N_7903,N_7038,N_7073);
nor U7904 (N_7904,N_7261,N_7436);
xnor U7905 (N_7905,N_7316,N_7390);
and U7906 (N_7906,N_7442,N_7441);
nor U7907 (N_7907,N_7005,N_7203);
nor U7908 (N_7908,N_7003,N_7491);
and U7909 (N_7909,N_7299,N_7469);
or U7910 (N_7910,N_7348,N_7422);
and U7911 (N_7911,N_7419,N_7493);
nor U7912 (N_7912,N_7429,N_7189);
nor U7913 (N_7913,N_7402,N_7131);
xnor U7914 (N_7914,N_7302,N_7423);
xor U7915 (N_7915,N_7177,N_7147);
and U7916 (N_7916,N_7130,N_7275);
nor U7917 (N_7917,N_7134,N_7212);
nor U7918 (N_7918,N_7350,N_7054);
nor U7919 (N_7919,N_7180,N_7068);
or U7920 (N_7920,N_7252,N_7124);
and U7921 (N_7921,N_7332,N_7188);
xor U7922 (N_7922,N_7420,N_7241);
xor U7923 (N_7923,N_7380,N_7496);
nor U7924 (N_7924,N_7424,N_7059);
xor U7925 (N_7925,N_7308,N_7052);
and U7926 (N_7926,N_7147,N_7078);
nand U7927 (N_7927,N_7252,N_7116);
and U7928 (N_7928,N_7363,N_7231);
xor U7929 (N_7929,N_7402,N_7348);
and U7930 (N_7930,N_7290,N_7262);
nor U7931 (N_7931,N_7116,N_7271);
xor U7932 (N_7932,N_7200,N_7360);
xor U7933 (N_7933,N_7112,N_7198);
and U7934 (N_7934,N_7403,N_7110);
nand U7935 (N_7935,N_7059,N_7285);
nand U7936 (N_7936,N_7333,N_7317);
nand U7937 (N_7937,N_7338,N_7309);
nand U7938 (N_7938,N_7477,N_7244);
and U7939 (N_7939,N_7089,N_7402);
or U7940 (N_7940,N_7065,N_7284);
nor U7941 (N_7941,N_7361,N_7329);
nand U7942 (N_7942,N_7321,N_7371);
xor U7943 (N_7943,N_7412,N_7114);
and U7944 (N_7944,N_7275,N_7213);
nor U7945 (N_7945,N_7481,N_7377);
xnor U7946 (N_7946,N_7342,N_7489);
nor U7947 (N_7947,N_7371,N_7418);
xor U7948 (N_7948,N_7193,N_7297);
and U7949 (N_7949,N_7208,N_7000);
or U7950 (N_7950,N_7209,N_7283);
xor U7951 (N_7951,N_7259,N_7288);
and U7952 (N_7952,N_7468,N_7088);
nor U7953 (N_7953,N_7236,N_7150);
and U7954 (N_7954,N_7464,N_7072);
or U7955 (N_7955,N_7254,N_7219);
nand U7956 (N_7956,N_7387,N_7190);
nor U7957 (N_7957,N_7169,N_7317);
or U7958 (N_7958,N_7246,N_7354);
or U7959 (N_7959,N_7189,N_7431);
nor U7960 (N_7960,N_7244,N_7130);
xnor U7961 (N_7961,N_7456,N_7399);
nor U7962 (N_7962,N_7449,N_7247);
or U7963 (N_7963,N_7461,N_7385);
xor U7964 (N_7964,N_7163,N_7130);
xor U7965 (N_7965,N_7109,N_7012);
and U7966 (N_7966,N_7249,N_7177);
xor U7967 (N_7967,N_7452,N_7302);
nor U7968 (N_7968,N_7226,N_7324);
xor U7969 (N_7969,N_7022,N_7357);
nand U7970 (N_7970,N_7359,N_7279);
xnor U7971 (N_7971,N_7059,N_7053);
nand U7972 (N_7972,N_7263,N_7090);
and U7973 (N_7973,N_7431,N_7074);
and U7974 (N_7974,N_7306,N_7163);
nand U7975 (N_7975,N_7344,N_7420);
or U7976 (N_7976,N_7011,N_7172);
or U7977 (N_7977,N_7069,N_7499);
xnor U7978 (N_7978,N_7068,N_7438);
or U7979 (N_7979,N_7003,N_7395);
nand U7980 (N_7980,N_7485,N_7302);
nor U7981 (N_7981,N_7051,N_7312);
nor U7982 (N_7982,N_7230,N_7361);
nand U7983 (N_7983,N_7242,N_7104);
nand U7984 (N_7984,N_7192,N_7217);
nand U7985 (N_7985,N_7251,N_7289);
and U7986 (N_7986,N_7232,N_7205);
nor U7987 (N_7987,N_7034,N_7496);
xor U7988 (N_7988,N_7186,N_7239);
and U7989 (N_7989,N_7004,N_7125);
xnor U7990 (N_7990,N_7192,N_7317);
or U7991 (N_7991,N_7247,N_7160);
nor U7992 (N_7992,N_7114,N_7419);
nor U7993 (N_7993,N_7102,N_7112);
and U7994 (N_7994,N_7437,N_7011);
nand U7995 (N_7995,N_7173,N_7302);
nand U7996 (N_7996,N_7085,N_7252);
xor U7997 (N_7997,N_7370,N_7267);
nand U7998 (N_7998,N_7136,N_7144);
nand U7999 (N_7999,N_7482,N_7280);
and U8000 (N_8000,N_7567,N_7886);
nor U8001 (N_8001,N_7584,N_7943);
nand U8002 (N_8002,N_7987,N_7551);
nor U8003 (N_8003,N_7509,N_7605);
or U8004 (N_8004,N_7579,N_7778);
nor U8005 (N_8005,N_7718,N_7773);
xor U8006 (N_8006,N_7601,N_7842);
xor U8007 (N_8007,N_7566,N_7595);
nor U8008 (N_8008,N_7911,N_7656);
xnor U8009 (N_8009,N_7699,N_7929);
and U8010 (N_8010,N_7755,N_7615);
xor U8011 (N_8011,N_7946,N_7978);
xnor U8012 (N_8012,N_7874,N_7899);
or U8013 (N_8013,N_7742,N_7514);
nand U8014 (N_8014,N_7997,N_7836);
nor U8015 (N_8015,N_7593,N_7519);
nor U8016 (N_8016,N_7541,N_7734);
nor U8017 (N_8017,N_7511,N_7954);
xor U8018 (N_8018,N_7654,N_7760);
nand U8019 (N_8019,N_7811,N_7746);
nor U8020 (N_8020,N_7591,N_7688);
xnor U8021 (N_8021,N_7833,N_7883);
nand U8022 (N_8022,N_7569,N_7722);
nor U8023 (N_8023,N_7802,N_7730);
xnor U8024 (N_8024,N_7905,N_7828);
nand U8025 (N_8025,N_7914,N_7621);
xnor U8026 (N_8026,N_7814,N_7554);
nand U8027 (N_8027,N_7664,N_7617);
and U8028 (N_8028,N_7646,N_7702);
xor U8029 (N_8029,N_7652,N_7574);
nand U8030 (N_8030,N_7684,N_7602);
and U8031 (N_8031,N_7558,N_7989);
and U8032 (N_8032,N_7651,N_7825);
xor U8033 (N_8033,N_7637,N_7645);
xor U8034 (N_8034,N_7629,N_7687);
nor U8035 (N_8035,N_7932,N_7927);
nand U8036 (N_8036,N_7990,N_7552);
xor U8037 (N_8037,N_7737,N_7852);
and U8038 (N_8038,N_7904,N_7985);
nor U8039 (N_8039,N_7623,N_7859);
nand U8040 (N_8040,N_7690,N_7530);
nor U8041 (N_8041,N_7919,N_7598);
nand U8042 (N_8042,N_7821,N_7830);
nand U8043 (N_8043,N_7662,N_7731);
xor U8044 (N_8044,N_7635,N_7910);
xnor U8045 (N_8045,N_7894,N_7638);
or U8046 (N_8046,N_7580,N_7515);
and U8047 (N_8047,N_7500,N_7780);
or U8048 (N_8048,N_7588,N_7994);
xnor U8049 (N_8049,N_7572,N_7771);
or U8050 (N_8050,N_7517,N_7763);
nor U8051 (N_8051,N_7855,N_7677);
and U8052 (N_8052,N_7784,N_7959);
and U8053 (N_8053,N_7634,N_7544);
or U8054 (N_8054,N_7856,N_7948);
nand U8055 (N_8055,N_7829,N_7800);
nand U8056 (N_8056,N_7626,N_7594);
and U8057 (N_8057,N_7777,N_7834);
or U8058 (N_8058,N_7522,N_7639);
nand U8059 (N_8059,N_7913,N_7736);
and U8060 (N_8060,N_7807,N_7951);
nor U8061 (N_8061,N_7658,N_7747);
nand U8062 (N_8062,N_7758,N_7930);
nand U8063 (N_8063,N_7741,N_7916);
nor U8064 (N_8064,N_7716,N_7901);
and U8065 (N_8065,N_7752,N_7879);
nand U8066 (N_8066,N_7643,N_7720);
nand U8067 (N_8067,N_7964,N_7714);
and U8068 (N_8068,N_7607,N_7738);
nand U8069 (N_8069,N_7912,N_7861);
nand U8070 (N_8070,N_7967,N_7681);
nor U8071 (N_8071,N_7695,N_7556);
nor U8072 (N_8072,N_7612,N_7884);
and U8073 (N_8073,N_7941,N_7765);
or U8074 (N_8074,N_7922,N_7858);
xnor U8075 (N_8075,N_7553,N_7876);
nor U8076 (N_8076,N_7715,N_7844);
nand U8077 (N_8077,N_7581,N_7640);
and U8078 (N_8078,N_7706,N_7957);
nand U8079 (N_8079,N_7586,N_7823);
xnor U8080 (N_8080,N_7863,N_7525);
nand U8081 (N_8081,N_7513,N_7878);
nor U8082 (N_8082,N_7642,N_7686);
and U8083 (N_8083,N_7712,N_7705);
nor U8084 (N_8084,N_7600,N_7794);
xnor U8085 (N_8085,N_7750,N_7512);
nor U8086 (N_8086,N_7669,N_7787);
xor U8087 (N_8087,N_7848,N_7975);
nand U8088 (N_8088,N_7933,N_7887);
xor U8089 (N_8089,N_7727,N_7613);
nor U8090 (N_8090,N_7703,N_7958);
and U8091 (N_8091,N_7641,N_7676);
and U8092 (N_8092,N_7835,N_7650);
xnor U8093 (N_8093,N_7696,N_7685);
and U8094 (N_8094,N_7862,N_7940);
nor U8095 (N_8095,N_7532,N_7824);
xor U8096 (N_8096,N_7620,N_7679);
nand U8097 (N_8097,N_7523,N_7663);
and U8098 (N_8098,N_7799,N_7938);
nor U8099 (N_8099,N_7816,N_7782);
and U8100 (N_8100,N_7575,N_7733);
nor U8101 (N_8101,N_7808,N_7768);
and U8102 (N_8102,N_7528,N_7561);
or U8103 (N_8103,N_7812,N_7762);
nor U8104 (N_8104,N_7896,N_7810);
nand U8105 (N_8105,N_7503,N_7770);
nor U8106 (N_8106,N_7798,N_7838);
or U8107 (N_8107,N_7724,N_7739);
and U8108 (N_8108,N_7991,N_7701);
and U8109 (N_8109,N_7535,N_7589);
or U8110 (N_8110,N_7564,N_7571);
xnor U8111 (N_8111,N_7804,N_7592);
or U8112 (N_8112,N_7890,N_7865);
nand U8113 (N_8113,N_7507,N_7772);
and U8114 (N_8114,N_7597,N_7944);
nor U8115 (N_8115,N_7900,N_7841);
nand U8116 (N_8116,N_7795,N_7850);
xor U8117 (N_8117,N_7960,N_7949);
nor U8118 (N_8118,N_7548,N_7539);
and U8119 (N_8119,N_7644,N_7839);
or U8120 (N_8120,N_7974,N_7536);
and U8121 (N_8121,N_7920,N_7806);
and U8122 (N_8122,N_7853,N_7783);
and U8123 (N_8123,N_7895,N_7757);
and U8124 (N_8124,N_7538,N_7504);
and U8125 (N_8125,N_7797,N_7764);
nand U8126 (N_8126,N_7837,N_7573);
xor U8127 (N_8127,N_7979,N_7700);
nor U8128 (N_8128,N_7533,N_7792);
or U8129 (N_8129,N_7648,N_7608);
and U8130 (N_8130,N_7893,N_7667);
nor U8131 (N_8131,N_7880,N_7546);
or U8132 (N_8132,N_7653,N_7832);
xnor U8133 (N_8133,N_7953,N_7857);
nand U8134 (N_8134,N_7998,N_7534);
and U8135 (N_8135,N_7691,N_7847);
and U8136 (N_8136,N_7756,N_7518);
and U8137 (N_8137,N_7968,N_7921);
or U8138 (N_8138,N_7549,N_7926);
xor U8139 (N_8139,N_7851,N_7871);
or U8140 (N_8140,N_7934,N_7971);
or U8141 (N_8141,N_7596,N_7697);
xor U8142 (N_8142,N_7576,N_7555);
and U8143 (N_8143,N_7945,N_7547);
xnor U8144 (N_8144,N_7729,N_7826);
or U8145 (N_8145,N_7988,N_7559);
nand U8146 (N_8146,N_7753,N_7708);
nor U8147 (N_8147,N_7993,N_7524);
and U8148 (N_8148,N_7976,N_7627);
or U8149 (N_8149,N_7903,N_7819);
and U8150 (N_8150,N_7962,N_7570);
nor U8151 (N_8151,N_7501,N_7585);
nand U8152 (N_8152,N_7508,N_7704);
xor U8153 (N_8153,N_7631,N_7775);
nor U8154 (N_8154,N_7505,N_7965);
nand U8155 (N_8155,N_7557,N_7560);
nand U8156 (N_8156,N_7732,N_7521);
nor U8157 (N_8157,N_7516,N_7952);
nor U8158 (N_8158,N_7693,N_7578);
nor U8159 (N_8159,N_7831,N_7745);
nand U8160 (N_8160,N_7622,N_7721);
or U8161 (N_8161,N_7980,N_7873);
and U8162 (N_8162,N_7633,N_7609);
nor U8163 (N_8163,N_7801,N_7671);
nand U8164 (N_8164,N_7999,N_7680);
xnor U8165 (N_8165,N_7761,N_7563);
nor U8166 (N_8166,N_7744,N_7906);
nor U8167 (N_8167,N_7779,N_7813);
or U8168 (N_8168,N_7809,N_7786);
xnor U8169 (N_8169,N_7907,N_7675);
nor U8170 (N_8170,N_7582,N_7728);
xor U8171 (N_8171,N_7502,N_7923);
nor U8172 (N_8172,N_7942,N_7611);
xnor U8173 (N_8173,N_7817,N_7986);
and U8174 (N_8174,N_7527,N_7628);
and U8175 (N_8175,N_7902,N_7754);
xor U8176 (N_8176,N_7774,N_7599);
or U8177 (N_8177,N_7791,N_7649);
or U8178 (N_8178,N_7776,N_7984);
nand U8179 (N_8179,N_7769,N_7543);
or U8180 (N_8180,N_7616,N_7520);
or U8181 (N_8181,N_7889,N_7694);
or U8182 (N_8182,N_7843,N_7937);
nand U8183 (N_8183,N_7568,N_7789);
xor U8184 (N_8184,N_7868,N_7785);
xnor U8185 (N_8185,N_7526,N_7888);
nor U8186 (N_8186,N_7939,N_7969);
and U8187 (N_8187,N_7881,N_7632);
or U8188 (N_8188,N_7864,N_7678);
nor U8189 (N_8189,N_7961,N_7796);
nand U8190 (N_8190,N_7790,N_7698);
and U8191 (N_8191,N_7542,N_7726);
nand U8192 (N_8192,N_7749,N_7740);
xnor U8193 (N_8193,N_7793,N_7854);
xor U8194 (N_8194,N_7606,N_7610);
and U8195 (N_8195,N_7885,N_7666);
and U8196 (N_8196,N_7689,N_7587);
and U8197 (N_8197,N_7992,N_7846);
and U8198 (N_8198,N_7866,N_7931);
nor U8199 (N_8199,N_7660,N_7565);
nor U8200 (N_8200,N_7966,N_7972);
xnor U8201 (N_8201,N_7877,N_7545);
xnor U8202 (N_8202,N_7709,N_7909);
or U8203 (N_8203,N_7657,N_7583);
xor U8204 (N_8204,N_7636,N_7982);
and U8205 (N_8205,N_7725,N_7537);
and U8206 (N_8206,N_7529,N_7735);
xor U8207 (N_8207,N_7918,N_7647);
xnor U8208 (N_8208,N_7781,N_7766);
nand U8209 (N_8209,N_7803,N_7717);
or U8210 (N_8210,N_7674,N_7743);
nor U8211 (N_8211,N_7867,N_7815);
or U8212 (N_8212,N_7977,N_7935);
nand U8213 (N_8213,N_7860,N_7692);
nand U8214 (N_8214,N_7590,N_7531);
nand U8215 (N_8215,N_7723,N_7875);
and U8216 (N_8216,N_7707,N_7788);
and U8217 (N_8217,N_7882,N_7619);
nor U8218 (N_8218,N_7872,N_7870);
xnor U8219 (N_8219,N_7822,N_7618);
xnor U8220 (N_8220,N_7973,N_7908);
nor U8221 (N_8221,N_7915,N_7947);
and U8222 (N_8222,N_7682,N_7996);
and U8223 (N_8223,N_7683,N_7719);
xnor U8224 (N_8224,N_7759,N_7748);
xnor U8225 (N_8225,N_7661,N_7550);
xor U8226 (N_8226,N_7950,N_7767);
xnor U8227 (N_8227,N_7668,N_7820);
nor U8228 (N_8228,N_7562,N_7655);
and U8229 (N_8229,N_7614,N_7936);
xor U8230 (N_8230,N_7665,N_7577);
or U8231 (N_8231,N_7805,N_7995);
and U8232 (N_8232,N_7928,N_7713);
xnor U8233 (N_8233,N_7827,N_7849);
xnor U8234 (N_8234,N_7540,N_7963);
or U8235 (N_8235,N_7845,N_7891);
and U8236 (N_8236,N_7970,N_7869);
xor U8237 (N_8237,N_7955,N_7630);
or U8238 (N_8238,N_7840,N_7925);
or U8239 (N_8239,N_7917,N_7897);
or U8240 (N_8240,N_7506,N_7956);
or U8241 (N_8241,N_7624,N_7711);
nand U8242 (N_8242,N_7710,N_7898);
or U8243 (N_8243,N_7659,N_7670);
and U8244 (N_8244,N_7625,N_7751);
or U8245 (N_8245,N_7672,N_7510);
and U8246 (N_8246,N_7983,N_7924);
nand U8247 (N_8247,N_7892,N_7603);
or U8248 (N_8248,N_7604,N_7818);
nand U8249 (N_8249,N_7673,N_7981);
nor U8250 (N_8250,N_7638,N_7866);
or U8251 (N_8251,N_7632,N_7528);
nor U8252 (N_8252,N_7668,N_7893);
nand U8253 (N_8253,N_7797,N_7662);
or U8254 (N_8254,N_7628,N_7526);
xnor U8255 (N_8255,N_7942,N_7518);
nor U8256 (N_8256,N_7802,N_7846);
and U8257 (N_8257,N_7913,N_7621);
or U8258 (N_8258,N_7781,N_7812);
xor U8259 (N_8259,N_7624,N_7978);
nor U8260 (N_8260,N_7669,N_7867);
and U8261 (N_8261,N_7624,N_7856);
or U8262 (N_8262,N_7927,N_7965);
xnor U8263 (N_8263,N_7971,N_7715);
nand U8264 (N_8264,N_7986,N_7558);
and U8265 (N_8265,N_7553,N_7593);
xnor U8266 (N_8266,N_7519,N_7582);
or U8267 (N_8267,N_7684,N_7792);
nand U8268 (N_8268,N_7543,N_7767);
nand U8269 (N_8269,N_7965,N_7580);
or U8270 (N_8270,N_7903,N_7884);
or U8271 (N_8271,N_7604,N_7933);
nand U8272 (N_8272,N_7957,N_7977);
nand U8273 (N_8273,N_7867,N_7889);
xnor U8274 (N_8274,N_7762,N_7748);
or U8275 (N_8275,N_7688,N_7987);
nand U8276 (N_8276,N_7820,N_7901);
or U8277 (N_8277,N_7935,N_7851);
nor U8278 (N_8278,N_7682,N_7835);
or U8279 (N_8279,N_7651,N_7709);
nand U8280 (N_8280,N_7930,N_7671);
or U8281 (N_8281,N_7613,N_7800);
nor U8282 (N_8282,N_7575,N_7685);
and U8283 (N_8283,N_7895,N_7946);
or U8284 (N_8284,N_7598,N_7664);
nand U8285 (N_8285,N_7951,N_7881);
and U8286 (N_8286,N_7739,N_7617);
or U8287 (N_8287,N_7987,N_7563);
xnor U8288 (N_8288,N_7865,N_7650);
and U8289 (N_8289,N_7635,N_7628);
or U8290 (N_8290,N_7540,N_7810);
and U8291 (N_8291,N_7858,N_7868);
nor U8292 (N_8292,N_7826,N_7700);
xor U8293 (N_8293,N_7809,N_7826);
or U8294 (N_8294,N_7990,N_7549);
nand U8295 (N_8295,N_7694,N_7923);
nand U8296 (N_8296,N_7765,N_7512);
or U8297 (N_8297,N_7933,N_7954);
nand U8298 (N_8298,N_7803,N_7718);
and U8299 (N_8299,N_7943,N_7698);
nand U8300 (N_8300,N_7590,N_7573);
or U8301 (N_8301,N_7822,N_7684);
nor U8302 (N_8302,N_7682,N_7962);
nor U8303 (N_8303,N_7832,N_7644);
or U8304 (N_8304,N_7870,N_7857);
or U8305 (N_8305,N_7870,N_7862);
and U8306 (N_8306,N_7813,N_7805);
or U8307 (N_8307,N_7752,N_7622);
and U8308 (N_8308,N_7871,N_7905);
xor U8309 (N_8309,N_7608,N_7686);
nand U8310 (N_8310,N_7515,N_7557);
nand U8311 (N_8311,N_7620,N_7861);
xor U8312 (N_8312,N_7668,N_7532);
nor U8313 (N_8313,N_7737,N_7638);
or U8314 (N_8314,N_7729,N_7668);
and U8315 (N_8315,N_7539,N_7705);
nor U8316 (N_8316,N_7772,N_7839);
and U8317 (N_8317,N_7546,N_7938);
xnor U8318 (N_8318,N_7589,N_7906);
nor U8319 (N_8319,N_7551,N_7662);
nor U8320 (N_8320,N_7833,N_7530);
xor U8321 (N_8321,N_7811,N_7545);
nor U8322 (N_8322,N_7633,N_7530);
xor U8323 (N_8323,N_7513,N_7912);
xor U8324 (N_8324,N_7716,N_7768);
or U8325 (N_8325,N_7772,N_7603);
xor U8326 (N_8326,N_7926,N_7536);
and U8327 (N_8327,N_7848,N_7986);
and U8328 (N_8328,N_7756,N_7503);
xor U8329 (N_8329,N_7894,N_7931);
xnor U8330 (N_8330,N_7833,N_7838);
xnor U8331 (N_8331,N_7878,N_7733);
or U8332 (N_8332,N_7774,N_7866);
and U8333 (N_8333,N_7592,N_7648);
nor U8334 (N_8334,N_7857,N_7613);
nand U8335 (N_8335,N_7748,N_7572);
xor U8336 (N_8336,N_7853,N_7531);
xor U8337 (N_8337,N_7772,N_7899);
nand U8338 (N_8338,N_7620,N_7814);
xor U8339 (N_8339,N_7712,N_7991);
xnor U8340 (N_8340,N_7630,N_7852);
xnor U8341 (N_8341,N_7776,N_7931);
nor U8342 (N_8342,N_7704,N_7990);
xnor U8343 (N_8343,N_7985,N_7707);
xor U8344 (N_8344,N_7641,N_7877);
and U8345 (N_8345,N_7948,N_7686);
or U8346 (N_8346,N_7844,N_7703);
nor U8347 (N_8347,N_7695,N_7806);
xnor U8348 (N_8348,N_7607,N_7613);
or U8349 (N_8349,N_7586,N_7690);
or U8350 (N_8350,N_7520,N_7671);
or U8351 (N_8351,N_7915,N_7783);
nand U8352 (N_8352,N_7900,N_7934);
xnor U8353 (N_8353,N_7509,N_7680);
or U8354 (N_8354,N_7507,N_7906);
nor U8355 (N_8355,N_7598,N_7733);
nor U8356 (N_8356,N_7799,N_7926);
nor U8357 (N_8357,N_7771,N_7846);
xor U8358 (N_8358,N_7623,N_7778);
xnor U8359 (N_8359,N_7544,N_7744);
and U8360 (N_8360,N_7512,N_7547);
and U8361 (N_8361,N_7918,N_7887);
nand U8362 (N_8362,N_7819,N_7957);
xor U8363 (N_8363,N_7997,N_7504);
nand U8364 (N_8364,N_7637,N_7930);
nor U8365 (N_8365,N_7847,N_7798);
and U8366 (N_8366,N_7764,N_7922);
or U8367 (N_8367,N_7668,N_7523);
nor U8368 (N_8368,N_7510,N_7770);
or U8369 (N_8369,N_7654,N_7558);
and U8370 (N_8370,N_7523,N_7932);
nand U8371 (N_8371,N_7834,N_7536);
nand U8372 (N_8372,N_7574,N_7821);
nand U8373 (N_8373,N_7662,N_7775);
xnor U8374 (N_8374,N_7756,N_7803);
and U8375 (N_8375,N_7558,N_7552);
or U8376 (N_8376,N_7868,N_7752);
nand U8377 (N_8377,N_7962,N_7657);
nand U8378 (N_8378,N_7668,N_7709);
or U8379 (N_8379,N_7891,N_7548);
nor U8380 (N_8380,N_7765,N_7533);
nor U8381 (N_8381,N_7544,N_7703);
or U8382 (N_8382,N_7530,N_7502);
nand U8383 (N_8383,N_7913,N_7574);
or U8384 (N_8384,N_7987,N_7795);
nor U8385 (N_8385,N_7651,N_7997);
nor U8386 (N_8386,N_7770,N_7793);
nor U8387 (N_8387,N_7581,N_7844);
nand U8388 (N_8388,N_7783,N_7756);
xor U8389 (N_8389,N_7747,N_7947);
xnor U8390 (N_8390,N_7980,N_7730);
or U8391 (N_8391,N_7725,N_7728);
nand U8392 (N_8392,N_7970,N_7595);
and U8393 (N_8393,N_7918,N_7785);
or U8394 (N_8394,N_7685,N_7780);
nor U8395 (N_8395,N_7609,N_7764);
xor U8396 (N_8396,N_7743,N_7967);
nand U8397 (N_8397,N_7549,N_7617);
nand U8398 (N_8398,N_7577,N_7508);
nor U8399 (N_8399,N_7942,N_7695);
or U8400 (N_8400,N_7857,N_7757);
and U8401 (N_8401,N_7775,N_7628);
and U8402 (N_8402,N_7812,N_7571);
nand U8403 (N_8403,N_7870,N_7745);
or U8404 (N_8404,N_7796,N_7511);
nor U8405 (N_8405,N_7552,N_7790);
nor U8406 (N_8406,N_7926,N_7753);
nand U8407 (N_8407,N_7539,N_7866);
xor U8408 (N_8408,N_7502,N_7799);
nand U8409 (N_8409,N_7908,N_7961);
or U8410 (N_8410,N_7666,N_7802);
xor U8411 (N_8411,N_7668,N_7865);
nor U8412 (N_8412,N_7588,N_7516);
nor U8413 (N_8413,N_7957,N_7520);
and U8414 (N_8414,N_7833,N_7873);
nand U8415 (N_8415,N_7838,N_7902);
xor U8416 (N_8416,N_7753,N_7789);
or U8417 (N_8417,N_7844,N_7878);
nor U8418 (N_8418,N_7746,N_7692);
or U8419 (N_8419,N_7623,N_7874);
nor U8420 (N_8420,N_7619,N_7865);
xor U8421 (N_8421,N_7580,N_7673);
nor U8422 (N_8422,N_7988,N_7800);
xor U8423 (N_8423,N_7525,N_7880);
and U8424 (N_8424,N_7839,N_7879);
or U8425 (N_8425,N_7721,N_7990);
or U8426 (N_8426,N_7893,N_7887);
and U8427 (N_8427,N_7725,N_7792);
xor U8428 (N_8428,N_7658,N_7850);
nand U8429 (N_8429,N_7615,N_7660);
nor U8430 (N_8430,N_7721,N_7686);
nor U8431 (N_8431,N_7820,N_7740);
nor U8432 (N_8432,N_7941,N_7591);
nor U8433 (N_8433,N_7814,N_7725);
nand U8434 (N_8434,N_7827,N_7943);
and U8435 (N_8435,N_7920,N_7705);
xor U8436 (N_8436,N_7778,N_7741);
and U8437 (N_8437,N_7616,N_7699);
nor U8438 (N_8438,N_7649,N_7621);
and U8439 (N_8439,N_7602,N_7642);
nand U8440 (N_8440,N_7956,N_7615);
nor U8441 (N_8441,N_7607,N_7913);
or U8442 (N_8442,N_7941,N_7901);
nand U8443 (N_8443,N_7704,N_7987);
nor U8444 (N_8444,N_7879,N_7860);
xor U8445 (N_8445,N_7814,N_7667);
xor U8446 (N_8446,N_7905,N_7568);
or U8447 (N_8447,N_7527,N_7816);
or U8448 (N_8448,N_7956,N_7802);
xnor U8449 (N_8449,N_7844,N_7879);
nor U8450 (N_8450,N_7929,N_7833);
and U8451 (N_8451,N_7580,N_7969);
or U8452 (N_8452,N_7809,N_7865);
or U8453 (N_8453,N_7766,N_7831);
and U8454 (N_8454,N_7777,N_7608);
and U8455 (N_8455,N_7995,N_7531);
or U8456 (N_8456,N_7713,N_7664);
nor U8457 (N_8457,N_7925,N_7568);
nor U8458 (N_8458,N_7732,N_7789);
nor U8459 (N_8459,N_7564,N_7516);
nor U8460 (N_8460,N_7886,N_7569);
nor U8461 (N_8461,N_7596,N_7973);
xnor U8462 (N_8462,N_7650,N_7670);
nor U8463 (N_8463,N_7783,N_7584);
nor U8464 (N_8464,N_7766,N_7650);
nand U8465 (N_8465,N_7859,N_7744);
xor U8466 (N_8466,N_7687,N_7892);
or U8467 (N_8467,N_7800,N_7506);
nor U8468 (N_8468,N_7684,N_7781);
nand U8469 (N_8469,N_7782,N_7667);
nor U8470 (N_8470,N_7988,N_7975);
nor U8471 (N_8471,N_7883,N_7597);
xor U8472 (N_8472,N_7931,N_7591);
nor U8473 (N_8473,N_7981,N_7711);
xnor U8474 (N_8474,N_7823,N_7801);
xor U8475 (N_8475,N_7600,N_7795);
xnor U8476 (N_8476,N_7810,N_7958);
nand U8477 (N_8477,N_7519,N_7579);
nor U8478 (N_8478,N_7794,N_7648);
nor U8479 (N_8479,N_7544,N_7986);
and U8480 (N_8480,N_7643,N_7934);
nor U8481 (N_8481,N_7516,N_7723);
xnor U8482 (N_8482,N_7810,N_7670);
xor U8483 (N_8483,N_7696,N_7722);
nand U8484 (N_8484,N_7751,N_7870);
or U8485 (N_8485,N_7555,N_7671);
xnor U8486 (N_8486,N_7790,N_7704);
xor U8487 (N_8487,N_7735,N_7843);
and U8488 (N_8488,N_7630,N_7873);
and U8489 (N_8489,N_7868,N_7851);
xor U8490 (N_8490,N_7847,N_7501);
nand U8491 (N_8491,N_7920,N_7717);
xor U8492 (N_8492,N_7567,N_7579);
and U8493 (N_8493,N_7836,N_7654);
xor U8494 (N_8494,N_7902,N_7542);
or U8495 (N_8495,N_7600,N_7949);
xnor U8496 (N_8496,N_7609,N_7553);
nor U8497 (N_8497,N_7913,N_7895);
and U8498 (N_8498,N_7654,N_7522);
nand U8499 (N_8499,N_7961,N_7871);
xor U8500 (N_8500,N_8057,N_8191);
and U8501 (N_8501,N_8216,N_8035);
and U8502 (N_8502,N_8165,N_8234);
or U8503 (N_8503,N_8329,N_8443);
nor U8504 (N_8504,N_8101,N_8140);
or U8505 (N_8505,N_8153,N_8463);
or U8506 (N_8506,N_8289,N_8173);
nor U8507 (N_8507,N_8037,N_8498);
nor U8508 (N_8508,N_8435,N_8485);
nor U8509 (N_8509,N_8146,N_8244);
or U8510 (N_8510,N_8398,N_8198);
nor U8511 (N_8511,N_8360,N_8074);
nor U8512 (N_8512,N_8411,N_8260);
nand U8513 (N_8513,N_8069,N_8113);
or U8514 (N_8514,N_8043,N_8431);
nor U8515 (N_8515,N_8039,N_8407);
nand U8516 (N_8516,N_8160,N_8156);
and U8517 (N_8517,N_8137,N_8040);
or U8518 (N_8518,N_8011,N_8305);
nand U8519 (N_8519,N_8449,N_8080);
xnor U8520 (N_8520,N_8051,N_8390);
xor U8521 (N_8521,N_8325,N_8450);
and U8522 (N_8522,N_8214,N_8127);
and U8523 (N_8523,N_8310,N_8161);
xor U8524 (N_8524,N_8048,N_8255);
xor U8525 (N_8525,N_8351,N_8277);
nand U8526 (N_8526,N_8397,N_8099);
and U8527 (N_8527,N_8404,N_8163);
nor U8528 (N_8528,N_8195,N_8418);
nor U8529 (N_8529,N_8287,N_8142);
and U8530 (N_8530,N_8425,N_8299);
or U8531 (N_8531,N_8338,N_8009);
and U8532 (N_8532,N_8433,N_8107);
nand U8533 (N_8533,N_8267,N_8208);
nand U8534 (N_8534,N_8259,N_8291);
or U8535 (N_8535,N_8362,N_8273);
nor U8536 (N_8536,N_8171,N_8236);
and U8537 (N_8537,N_8182,N_8293);
and U8538 (N_8538,N_8085,N_8175);
xor U8539 (N_8539,N_8220,N_8344);
and U8540 (N_8540,N_8081,N_8100);
nor U8541 (N_8541,N_8031,N_8215);
nor U8542 (N_8542,N_8428,N_8205);
nand U8543 (N_8543,N_8477,N_8478);
and U8544 (N_8544,N_8394,N_8123);
and U8545 (N_8545,N_8001,N_8312);
or U8546 (N_8546,N_8370,N_8281);
xnor U8547 (N_8547,N_8251,N_8166);
xnor U8548 (N_8548,N_8484,N_8374);
or U8549 (N_8549,N_8337,N_8377);
nand U8550 (N_8550,N_8445,N_8353);
nor U8551 (N_8551,N_8423,N_8015);
or U8552 (N_8552,N_8188,N_8049);
nand U8553 (N_8553,N_8062,N_8341);
nand U8554 (N_8554,N_8033,N_8415);
and U8555 (N_8555,N_8228,N_8002);
xor U8556 (N_8556,N_8479,N_8438);
or U8557 (N_8557,N_8053,N_8465);
nand U8558 (N_8558,N_8358,N_8087);
and U8559 (N_8559,N_8496,N_8400);
and U8560 (N_8560,N_8439,N_8481);
nor U8561 (N_8561,N_8006,N_8444);
nor U8562 (N_8562,N_8238,N_8242);
or U8563 (N_8563,N_8239,N_8066);
xnor U8564 (N_8564,N_8256,N_8356);
nand U8565 (N_8565,N_8280,N_8336);
nand U8566 (N_8566,N_8168,N_8247);
or U8567 (N_8567,N_8046,N_8417);
nor U8568 (N_8568,N_8311,N_8410);
and U8569 (N_8569,N_8467,N_8275);
xnor U8570 (N_8570,N_8089,N_8401);
and U8571 (N_8571,N_8105,N_8131);
or U8572 (N_8572,N_8207,N_8098);
nor U8573 (N_8573,N_8248,N_8120);
nor U8574 (N_8574,N_8096,N_8427);
nand U8575 (N_8575,N_8308,N_8409);
nor U8576 (N_8576,N_8170,N_8118);
nor U8577 (N_8577,N_8393,N_8441);
or U8578 (N_8578,N_8488,N_8047);
nand U8579 (N_8579,N_8169,N_8257);
nand U8580 (N_8580,N_8422,N_8283);
and U8581 (N_8581,N_8253,N_8451);
and U8582 (N_8582,N_8038,N_8384);
nand U8583 (N_8583,N_8392,N_8133);
and U8584 (N_8584,N_8482,N_8332);
and U8585 (N_8585,N_8212,N_8327);
and U8586 (N_8586,N_8326,N_8104);
nand U8587 (N_8587,N_8174,N_8399);
and U8588 (N_8588,N_8204,N_8284);
xnor U8589 (N_8589,N_8064,N_8029);
or U8590 (N_8590,N_8381,N_8012);
xor U8591 (N_8591,N_8458,N_8333);
nand U8592 (N_8592,N_8167,N_8237);
and U8593 (N_8593,N_8318,N_8402);
xor U8594 (N_8594,N_8265,N_8456);
or U8595 (N_8595,N_8290,N_8246);
nand U8596 (N_8596,N_8487,N_8454);
nor U8597 (N_8597,N_8112,N_8008);
or U8598 (N_8598,N_8288,N_8295);
and U8599 (N_8599,N_8056,N_8187);
xnor U8600 (N_8600,N_8313,N_8494);
and U8601 (N_8601,N_8181,N_8322);
or U8602 (N_8602,N_8403,N_8379);
nand U8603 (N_8603,N_8486,N_8493);
or U8604 (N_8604,N_8152,N_8278);
nor U8605 (N_8605,N_8178,N_8079);
nor U8606 (N_8606,N_8294,N_8206);
nand U8607 (N_8607,N_8339,N_8190);
and U8608 (N_8608,N_8321,N_8391);
xor U8609 (N_8609,N_8061,N_8328);
nand U8610 (N_8610,N_8218,N_8406);
or U8611 (N_8611,N_8395,N_8230);
or U8612 (N_8612,N_8405,N_8106);
nor U8613 (N_8613,N_8297,N_8453);
xor U8614 (N_8614,N_8192,N_8217);
or U8615 (N_8615,N_8309,N_8426);
nor U8616 (N_8616,N_8301,N_8201);
nor U8617 (N_8617,N_8231,N_8082);
or U8618 (N_8618,N_8372,N_8093);
xor U8619 (N_8619,N_8375,N_8014);
xnor U8620 (N_8620,N_8004,N_8462);
or U8621 (N_8621,N_8306,N_8073);
nor U8622 (N_8622,N_8473,N_8382);
nor U8623 (N_8623,N_8314,N_8420);
nand U8624 (N_8624,N_8032,N_8067);
and U8625 (N_8625,N_8235,N_8474);
nor U8626 (N_8626,N_8022,N_8272);
and U8627 (N_8627,N_8357,N_8386);
and U8628 (N_8628,N_8495,N_8119);
and U8629 (N_8629,N_8437,N_8219);
or U8630 (N_8630,N_8472,N_8020);
nor U8631 (N_8631,N_8194,N_8292);
xnor U8632 (N_8632,N_8468,N_8138);
xnor U8633 (N_8633,N_8319,N_8490);
xor U8634 (N_8634,N_8180,N_8497);
nand U8635 (N_8635,N_8111,N_8457);
xor U8636 (N_8636,N_8252,N_8145);
nor U8637 (N_8637,N_8068,N_8050);
nand U8638 (N_8638,N_8072,N_8005);
and U8639 (N_8639,N_8078,N_8134);
nand U8640 (N_8640,N_8058,N_8148);
nand U8641 (N_8641,N_8109,N_8286);
nor U8642 (N_8642,N_8010,N_8210);
nand U8643 (N_8643,N_8116,N_8075);
nor U8644 (N_8644,N_8376,N_8090);
and U8645 (N_8645,N_8203,N_8324);
or U8646 (N_8646,N_8317,N_8027);
nor U8647 (N_8647,N_8373,N_8355);
and U8648 (N_8648,N_8013,N_8026);
or U8649 (N_8649,N_8350,N_8250);
nor U8650 (N_8650,N_8269,N_8440);
or U8651 (N_8651,N_8455,N_8227);
xor U8652 (N_8652,N_8150,N_8019);
xor U8653 (N_8653,N_8475,N_8183);
xor U8654 (N_8654,N_8442,N_8264);
xnor U8655 (N_8655,N_8076,N_8489);
nor U8656 (N_8656,N_8470,N_8366);
nor U8657 (N_8657,N_8364,N_8065);
xnor U8658 (N_8658,N_8108,N_8249);
and U8659 (N_8659,N_8126,N_8385);
nor U8660 (N_8660,N_8320,N_8083);
and U8661 (N_8661,N_8052,N_8266);
or U8662 (N_8662,N_8158,N_8349);
xor U8663 (N_8663,N_8185,N_8361);
and U8664 (N_8664,N_8448,N_8464);
and U8665 (N_8665,N_8279,N_8424);
xor U8666 (N_8666,N_8077,N_8114);
and U8667 (N_8667,N_8121,N_8179);
or U8668 (N_8668,N_8223,N_8492);
nor U8669 (N_8669,N_8304,N_8254);
nor U8670 (N_8670,N_8303,N_8164);
nand U8671 (N_8671,N_8421,N_8177);
nor U8672 (N_8672,N_8446,N_8300);
xor U8673 (N_8673,N_8434,N_8276);
or U8674 (N_8674,N_8141,N_8389);
and U8675 (N_8675,N_8071,N_8323);
xor U8676 (N_8676,N_8232,N_8115);
nor U8677 (N_8677,N_8018,N_8483);
or U8678 (N_8678,N_8193,N_8088);
nor U8679 (N_8679,N_8459,N_8030);
and U8680 (N_8680,N_8091,N_8343);
xor U8681 (N_8681,N_8285,N_8476);
and U8682 (N_8682,N_8388,N_8028);
xnor U8683 (N_8683,N_8136,N_8245);
nand U8684 (N_8684,N_8128,N_8282);
nand U8685 (N_8685,N_8184,N_8176);
and U8686 (N_8686,N_8155,N_8025);
and U8687 (N_8687,N_8086,N_8197);
and U8688 (N_8688,N_8034,N_8396);
nor U8689 (N_8689,N_8414,N_8466);
or U8690 (N_8690,N_8084,N_8130);
nor U8691 (N_8691,N_8240,N_8348);
or U8692 (N_8692,N_8335,N_8042);
or U8693 (N_8693,N_8225,N_8480);
nand U8694 (N_8694,N_8147,N_8094);
and U8695 (N_8695,N_8172,N_8369);
nand U8696 (N_8696,N_8229,N_8261);
xnor U8697 (N_8697,N_8387,N_8471);
nor U8698 (N_8698,N_8157,N_8226);
nand U8699 (N_8699,N_8243,N_8296);
nor U8700 (N_8700,N_8271,N_8059);
xnor U8701 (N_8701,N_8380,N_8044);
nor U8702 (N_8702,N_8202,N_8095);
xor U8703 (N_8703,N_8054,N_8383);
nor U8704 (N_8704,N_8378,N_8149);
nor U8705 (N_8705,N_8346,N_8063);
nor U8706 (N_8706,N_8144,N_8021);
nand U8707 (N_8707,N_8222,N_8200);
and U8708 (N_8708,N_8447,N_8432);
and U8709 (N_8709,N_8302,N_8262);
and U8710 (N_8710,N_8258,N_8003);
and U8711 (N_8711,N_8045,N_8060);
or U8712 (N_8712,N_8122,N_8092);
nand U8713 (N_8713,N_8154,N_8491);
nand U8714 (N_8714,N_8196,N_8365);
nor U8715 (N_8715,N_8347,N_8330);
xor U8716 (N_8716,N_8221,N_8110);
nand U8717 (N_8717,N_8268,N_8016);
and U8718 (N_8718,N_8416,N_8270);
and U8719 (N_8719,N_8316,N_8129);
and U8720 (N_8720,N_8461,N_8460);
nor U8721 (N_8721,N_8340,N_8135);
or U8722 (N_8722,N_8000,N_8367);
nand U8723 (N_8723,N_8359,N_8209);
nand U8724 (N_8724,N_8124,N_8419);
nor U8725 (N_8725,N_8363,N_8159);
nand U8726 (N_8726,N_8070,N_8162);
and U8727 (N_8727,N_8023,N_8274);
nor U8728 (N_8728,N_8017,N_8452);
nor U8729 (N_8729,N_8368,N_8354);
nand U8730 (N_8730,N_8103,N_8413);
xor U8731 (N_8731,N_8211,N_8189);
nor U8732 (N_8732,N_8412,N_8233);
or U8733 (N_8733,N_8430,N_8097);
or U8734 (N_8734,N_8307,N_8224);
xor U8735 (N_8735,N_8186,N_8315);
and U8736 (N_8736,N_8334,N_8429);
nand U8737 (N_8737,N_8241,N_8055);
xnor U8738 (N_8738,N_8408,N_8125);
nand U8739 (N_8739,N_8436,N_8132);
xnor U8740 (N_8740,N_8102,N_8143);
or U8741 (N_8741,N_8151,N_8117);
xnor U8742 (N_8742,N_8041,N_8036);
xnor U8743 (N_8743,N_8139,N_8371);
and U8744 (N_8744,N_8345,N_8213);
or U8745 (N_8745,N_8298,N_8331);
xnor U8746 (N_8746,N_8469,N_8007);
nor U8747 (N_8747,N_8499,N_8024);
or U8748 (N_8748,N_8342,N_8352);
nand U8749 (N_8749,N_8263,N_8199);
or U8750 (N_8750,N_8003,N_8430);
or U8751 (N_8751,N_8149,N_8414);
and U8752 (N_8752,N_8444,N_8348);
and U8753 (N_8753,N_8011,N_8362);
and U8754 (N_8754,N_8307,N_8218);
xor U8755 (N_8755,N_8436,N_8487);
xor U8756 (N_8756,N_8476,N_8465);
and U8757 (N_8757,N_8139,N_8045);
nor U8758 (N_8758,N_8445,N_8491);
nor U8759 (N_8759,N_8105,N_8016);
nand U8760 (N_8760,N_8412,N_8165);
nor U8761 (N_8761,N_8242,N_8345);
nand U8762 (N_8762,N_8428,N_8296);
and U8763 (N_8763,N_8399,N_8486);
nor U8764 (N_8764,N_8082,N_8363);
and U8765 (N_8765,N_8260,N_8156);
or U8766 (N_8766,N_8250,N_8426);
or U8767 (N_8767,N_8334,N_8333);
or U8768 (N_8768,N_8472,N_8056);
nand U8769 (N_8769,N_8489,N_8425);
nor U8770 (N_8770,N_8028,N_8374);
nor U8771 (N_8771,N_8047,N_8212);
or U8772 (N_8772,N_8003,N_8118);
and U8773 (N_8773,N_8206,N_8236);
nand U8774 (N_8774,N_8084,N_8433);
nor U8775 (N_8775,N_8447,N_8146);
nor U8776 (N_8776,N_8109,N_8103);
or U8777 (N_8777,N_8341,N_8290);
and U8778 (N_8778,N_8440,N_8161);
or U8779 (N_8779,N_8062,N_8384);
and U8780 (N_8780,N_8119,N_8404);
nor U8781 (N_8781,N_8340,N_8074);
nor U8782 (N_8782,N_8027,N_8210);
nor U8783 (N_8783,N_8331,N_8191);
or U8784 (N_8784,N_8116,N_8185);
nand U8785 (N_8785,N_8019,N_8060);
and U8786 (N_8786,N_8203,N_8124);
nand U8787 (N_8787,N_8484,N_8200);
xnor U8788 (N_8788,N_8410,N_8208);
and U8789 (N_8789,N_8136,N_8338);
nor U8790 (N_8790,N_8368,N_8387);
or U8791 (N_8791,N_8176,N_8386);
xor U8792 (N_8792,N_8156,N_8422);
xor U8793 (N_8793,N_8312,N_8467);
nor U8794 (N_8794,N_8329,N_8428);
nor U8795 (N_8795,N_8276,N_8459);
xor U8796 (N_8796,N_8083,N_8216);
and U8797 (N_8797,N_8052,N_8008);
nor U8798 (N_8798,N_8210,N_8349);
or U8799 (N_8799,N_8244,N_8140);
or U8800 (N_8800,N_8204,N_8302);
or U8801 (N_8801,N_8093,N_8036);
nor U8802 (N_8802,N_8112,N_8291);
nand U8803 (N_8803,N_8189,N_8434);
and U8804 (N_8804,N_8410,N_8385);
nand U8805 (N_8805,N_8154,N_8340);
nor U8806 (N_8806,N_8096,N_8314);
and U8807 (N_8807,N_8431,N_8420);
nand U8808 (N_8808,N_8208,N_8233);
xnor U8809 (N_8809,N_8365,N_8480);
xor U8810 (N_8810,N_8253,N_8364);
nor U8811 (N_8811,N_8462,N_8315);
or U8812 (N_8812,N_8108,N_8166);
or U8813 (N_8813,N_8079,N_8378);
or U8814 (N_8814,N_8208,N_8323);
or U8815 (N_8815,N_8199,N_8258);
or U8816 (N_8816,N_8179,N_8114);
xnor U8817 (N_8817,N_8258,N_8354);
nand U8818 (N_8818,N_8038,N_8160);
or U8819 (N_8819,N_8059,N_8422);
or U8820 (N_8820,N_8288,N_8410);
nand U8821 (N_8821,N_8263,N_8188);
xnor U8822 (N_8822,N_8164,N_8384);
or U8823 (N_8823,N_8012,N_8415);
xor U8824 (N_8824,N_8278,N_8042);
or U8825 (N_8825,N_8422,N_8034);
and U8826 (N_8826,N_8219,N_8060);
nand U8827 (N_8827,N_8451,N_8470);
nor U8828 (N_8828,N_8369,N_8426);
nor U8829 (N_8829,N_8312,N_8210);
nand U8830 (N_8830,N_8448,N_8248);
or U8831 (N_8831,N_8222,N_8403);
nor U8832 (N_8832,N_8489,N_8055);
nor U8833 (N_8833,N_8145,N_8413);
and U8834 (N_8834,N_8267,N_8300);
or U8835 (N_8835,N_8450,N_8470);
nand U8836 (N_8836,N_8131,N_8073);
and U8837 (N_8837,N_8265,N_8415);
nor U8838 (N_8838,N_8301,N_8105);
xnor U8839 (N_8839,N_8072,N_8194);
xor U8840 (N_8840,N_8372,N_8408);
xnor U8841 (N_8841,N_8443,N_8499);
xor U8842 (N_8842,N_8026,N_8347);
nand U8843 (N_8843,N_8235,N_8408);
and U8844 (N_8844,N_8287,N_8076);
nand U8845 (N_8845,N_8447,N_8478);
xnor U8846 (N_8846,N_8391,N_8313);
xor U8847 (N_8847,N_8400,N_8330);
nor U8848 (N_8848,N_8097,N_8373);
and U8849 (N_8849,N_8417,N_8160);
xnor U8850 (N_8850,N_8390,N_8234);
nand U8851 (N_8851,N_8447,N_8269);
nand U8852 (N_8852,N_8413,N_8381);
xor U8853 (N_8853,N_8002,N_8294);
or U8854 (N_8854,N_8383,N_8259);
nor U8855 (N_8855,N_8482,N_8289);
nand U8856 (N_8856,N_8245,N_8253);
and U8857 (N_8857,N_8084,N_8497);
xor U8858 (N_8858,N_8348,N_8043);
nand U8859 (N_8859,N_8034,N_8401);
nand U8860 (N_8860,N_8059,N_8343);
xnor U8861 (N_8861,N_8148,N_8256);
nor U8862 (N_8862,N_8205,N_8006);
nor U8863 (N_8863,N_8427,N_8003);
and U8864 (N_8864,N_8252,N_8455);
xnor U8865 (N_8865,N_8254,N_8069);
xnor U8866 (N_8866,N_8351,N_8128);
xor U8867 (N_8867,N_8236,N_8273);
nand U8868 (N_8868,N_8493,N_8379);
xnor U8869 (N_8869,N_8188,N_8360);
nand U8870 (N_8870,N_8012,N_8197);
and U8871 (N_8871,N_8392,N_8246);
or U8872 (N_8872,N_8316,N_8190);
xor U8873 (N_8873,N_8087,N_8077);
nand U8874 (N_8874,N_8386,N_8460);
nand U8875 (N_8875,N_8461,N_8138);
xnor U8876 (N_8876,N_8427,N_8483);
nand U8877 (N_8877,N_8186,N_8418);
or U8878 (N_8878,N_8290,N_8329);
or U8879 (N_8879,N_8070,N_8319);
or U8880 (N_8880,N_8030,N_8402);
and U8881 (N_8881,N_8412,N_8433);
nor U8882 (N_8882,N_8431,N_8156);
nand U8883 (N_8883,N_8355,N_8432);
nand U8884 (N_8884,N_8161,N_8238);
nand U8885 (N_8885,N_8290,N_8422);
nand U8886 (N_8886,N_8166,N_8118);
or U8887 (N_8887,N_8007,N_8046);
nand U8888 (N_8888,N_8236,N_8305);
nand U8889 (N_8889,N_8250,N_8044);
and U8890 (N_8890,N_8383,N_8308);
nor U8891 (N_8891,N_8285,N_8316);
or U8892 (N_8892,N_8194,N_8054);
or U8893 (N_8893,N_8204,N_8232);
nor U8894 (N_8894,N_8037,N_8226);
nand U8895 (N_8895,N_8361,N_8196);
nand U8896 (N_8896,N_8387,N_8297);
nor U8897 (N_8897,N_8263,N_8194);
or U8898 (N_8898,N_8131,N_8349);
or U8899 (N_8899,N_8485,N_8255);
nand U8900 (N_8900,N_8156,N_8240);
nand U8901 (N_8901,N_8371,N_8414);
nor U8902 (N_8902,N_8421,N_8245);
or U8903 (N_8903,N_8021,N_8233);
xor U8904 (N_8904,N_8089,N_8019);
and U8905 (N_8905,N_8166,N_8047);
nor U8906 (N_8906,N_8473,N_8067);
xor U8907 (N_8907,N_8206,N_8459);
nor U8908 (N_8908,N_8051,N_8103);
and U8909 (N_8909,N_8429,N_8465);
nand U8910 (N_8910,N_8108,N_8409);
or U8911 (N_8911,N_8019,N_8043);
nor U8912 (N_8912,N_8037,N_8460);
nand U8913 (N_8913,N_8208,N_8068);
and U8914 (N_8914,N_8182,N_8209);
or U8915 (N_8915,N_8434,N_8265);
and U8916 (N_8916,N_8233,N_8388);
xnor U8917 (N_8917,N_8245,N_8312);
nor U8918 (N_8918,N_8465,N_8319);
nand U8919 (N_8919,N_8116,N_8265);
and U8920 (N_8920,N_8426,N_8028);
and U8921 (N_8921,N_8430,N_8087);
nand U8922 (N_8922,N_8349,N_8149);
xor U8923 (N_8923,N_8009,N_8268);
or U8924 (N_8924,N_8211,N_8415);
xnor U8925 (N_8925,N_8338,N_8452);
or U8926 (N_8926,N_8473,N_8261);
or U8927 (N_8927,N_8443,N_8072);
xnor U8928 (N_8928,N_8286,N_8287);
nor U8929 (N_8929,N_8020,N_8302);
and U8930 (N_8930,N_8094,N_8157);
nand U8931 (N_8931,N_8194,N_8398);
nand U8932 (N_8932,N_8108,N_8161);
or U8933 (N_8933,N_8299,N_8237);
nand U8934 (N_8934,N_8340,N_8425);
nor U8935 (N_8935,N_8285,N_8103);
xor U8936 (N_8936,N_8268,N_8262);
xnor U8937 (N_8937,N_8081,N_8457);
and U8938 (N_8938,N_8233,N_8096);
nor U8939 (N_8939,N_8102,N_8053);
or U8940 (N_8940,N_8438,N_8444);
nor U8941 (N_8941,N_8307,N_8131);
nand U8942 (N_8942,N_8468,N_8183);
nor U8943 (N_8943,N_8406,N_8094);
nor U8944 (N_8944,N_8034,N_8440);
or U8945 (N_8945,N_8076,N_8220);
or U8946 (N_8946,N_8343,N_8070);
and U8947 (N_8947,N_8063,N_8118);
or U8948 (N_8948,N_8033,N_8306);
xor U8949 (N_8949,N_8013,N_8106);
nand U8950 (N_8950,N_8044,N_8203);
nand U8951 (N_8951,N_8056,N_8199);
xnor U8952 (N_8952,N_8323,N_8065);
nand U8953 (N_8953,N_8245,N_8138);
and U8954 (N_8954,N_8348,N_8285);
nand U8955 (N_8955,N_8348,N_8006);
nand U8956 (N_8956,N_8272,N_8157);
nand U8957 (N_8957,N_8089,N_8162);
and U8958 (N_8958,N_8040,N_8177);
nor U8959 (N_8959,N_8258,N_8105);
nor U8960 (N_8960,N_8272,N_8388);
nand U8961 (N_8961,N_8393,N_8263);
and U8962 (N_8962,N_8261,N_8209);
xor U8963 (N_8963,N_8297,N_8471);
nor U8964 (N_8964,N_8171,N_8301);
or U8965 (N_8965,N_8304,N_8260);
nand U8966 (N_8966,N_8097,N_8184);
and U8967 (N_8967,N_8294,N_8366);
and U8968 (N_8968,N_8151,N_8094);
nor U8969 (N_8969,N_8011,N_8036);
and U8970 (N_8970,N_8190,N_8389);
nor U8971 (N_8971,N_8041,N_8319);
and U8972 (N_8972,N_8465,N_8004);
or U8973 (N_8973,N_8293,N_8029);
xnor U8974 (N_8974,N_8030,N_8422);
and U8975 (N_8975,N_8205,N_8399);
and U8976 (N_8976,N_8353,N_8199);
and U8977 (N_8977,N_8112,N_8235);
and U8978 (N_8978,N_8498,N_8329);
nor U8979 (N_8979,N_8406,N_8442);
and U8980 (N_8980,N_8336,N_8202);
xnor U8981 (N_8981,N_8096,N_8213);
nor U8982 (N_8982,N_8237,N_8376);
nand U8983 (N_8983,N_8077,N_8150);
nand U8984 (N_8984,N_8489,N_8385);
and U8985 (N_8985,N_8379,N_8434);
xor U8986 (N_8986,N_8007,N_8251);
or U8987 (N_8987,N_8303,N_8013);
and U8988 (N_8988,N_8400,N_8324);
xor U8989 (N_8989,N_8091,N_8152);
xor U8990 (N_8990,N_8088,N_8308);
and U8991 (N_8991,N_8241,N_8083);
and U8992 (N_8992,N_8481,N_8488);
and U8993 (N_8993,N_8355,N_8277);
and U8994 (N_8994,N_8122,N_8090);
xor U8995 (N_8995,N_8100,N_8119);
or U8996 (N_8996,N_8279,N_8099);
and U8997 (N_8997,N_8119,N_8182);
nor U8998 (N_8998,N_8431,N_8177);
nor U8999 (N_8999,N_8184,N_8431);
and U9000 (N_9000,N_8994,N_8958);
xnor U9001 (N_9001,N_8640,N_8893);
nand U9002 (N_9002,N_8954,N_8961);
nor U9003 (N_9003,N_8684,N_8591);
nor U9004 (N_9004,N_8501,N_8826);
and U9005 (N_9005,N_8946,N_8653);
xor U9006 (N_9006,N_8854,N_8538);
and U9007 (N_9007,N_8533,N_8633);
and U9008 (N_9008,N_8770,N_8894);
nor U9009 (N_9009,N_8839,N_8705);
nor U9010 (N_9010,N_8805,N_8786);
xor U9011 (N_9011,N_8742,N_8689);
and U9012 (N_9012,N_8857,N_8852);
nand U9013 (N_9013,N_8644,N_8790);
and U9014 (N_9014,N_8755,N_8808);
nand U9015 (N_9015,N_8882,N_8575);
nand U9016 (N_9016,N_8835,N_8980);
nor U9017 (N_9017,N_8821,N_8645);
xor U9018 (N_9018,N_8841,N_8701);
xnor U9019 (N_9019,N_8616,N_8995);
or U9020 (N_9020,N_8677,N_8666);
nand U9021 (N_9021,N_8508,N_8801);
and U9022 (N_9022,N_8837,N_8972);
nor U9023 (N_9023,N_8756,N_8788);
or U9024 (N_9024,N_8990,N_8588);
or U9025 (N_9025,N_8696,N_8500);
or U9026 (N_9026,N_8606,N_8962);
nor U9027 (N_9027,N_8728,N_8829);
nand U9028 (N_9028,N_8593,N_8943);
nor U9029 (N_9029,N_8559,N_8667);
or U9030 (N_9030,N_8897,N_8938);
and U9031 (N_9031,N_8827,N_8625);
and U9032 (N_9032,N_8881,N_8964);
nor U9033 (N_9033,N_8914,N_8899);
nor U9034 (N_9034,N_8678,N_8642);
or U9035 (N_9035,N_8657,N_8627);
xor U9036 (N_9036,N_8831,N_8598);
nor U9037 (N_9037,N_8860,N_8524);
or U9038 (N_9038,N_8834,N_8630);
or U9039 (N_9039,N_8996,N_8722);
and U9040 (N_9040,N_8898,N_8842);
nor U9041 (N_9041,N_8798,N_8521);
xnor U9042 (N_9042,N_8953,N_8694);
xnor U9043 (N_9043,N_8804,N_8937);
nor U9044 (N_9044,N_8517,N_8942);
nor U9045 (N_9045,N_8879,N_8718);
nor U9046 (N_9046,N_8939,N_8621);
nand U9047 (N_9047,N_8719,N_8558);
xor U9048 (N_9048,N_8512,N_8960);
or U9049 (N_9049,N_8570,N_8869);
and U9050 (N_9050,N_8776,N_8909);
xor U9051 (N_9051,N_8510,N_8844);
xnor U9052 (N_9052,N_8594,N_8795);
or U9053 (N_9053,N_8608,N_8502);
nand U9054 (N_9054,N_8865,N_8766);
nor U9055 (N_9055,N_8850,N_8966);
nor U9056 (N_9056,N_8761,N_8870);
nand U9057 (N_9057,N_8840,N_8582);
and U9058 (N_9058,N_8771,N_8875);
nor U9059 (N_9059,N_8522,N_8927);
and U9060 (N_9060,N_8520,N_8583);
and U9061 (N_9061,N_8529,N_8765);
and U9062 (N_9062,N_8992,N_8622);
and U9063 (N_9063,N_8631,N_8843);
and U9064 (N_9064,N_8934,N_8671);
xor U9065 (N_9065,N_8643,N_8886);
nand U9066 (N_9066,N_8905,N_8572);
or U9067 (N_9067,N_8717,N_8769);
nor U9068 (N_9068,N_8861,N_8910);
xnor U9069 (N_9069,N_8963,N_8562);
or U9070 (N_9070,N_8955,N_8998);
and U9071 (N_9071,N_8849,N_8968);
or U9072 (N_9072,N_8949,N_8789);
and U9073 (N_9073,N_8546,N_8634);
and U9074 (N_9074,N_8820,N_8611);
or U9075 (N_9075,N_8971,N_8679);
xor U9076 (N_9076,N_8977,N_8751);
nor U9077 (N_9077,N_8750,N_8816);
and U9078 (N_9078,N_8668,N_8615);
nand U9079 (N_9079,N_8885,N_8768);
or U9080 (N_9080,N_8950,N_8989);
and U9081 (N_9081,N_8695,N_8815);
xnor U9082 (N_9082,N_8824,N_8604);
and U9083 (N_9083,N_8628,N_8782);
nor U9084 (N_9084,N_8982,N_8764);
nand U9085 (N_9085,N_8889,N_8532);
and U9086 (N_9086,N_8749,N_8930);
nand U9087 (N_9087,N_8708,N_8799);
and U9088 (N_9088,N_8867,N_8896);
and U9089 (N_9089,N_8637,N_8557);
nand U9090 (N_9090,N_8550,N_8760);
xnor U9091 (N_9091,N_8763,N_8754);
or U9092 (N_9092,N_8932,N_8587);
nor U9093 (N_9093,N_8864,N_8757);
nor U9094 (N_9094,N_8721,N_8911);
nor U9095 (N_9095,N_8813,N_8603);
nor U9096 (N_9096,N_8874,N_8748);
or U9097 (N_9097,N_8812,N_8727);
nor U9098 (N_9098,N_8759,N_8856);
nor U9099 (N_9099,N_8887,N_8567);
nand U9100 (N_9100,N_8851,N_8981);
and U9101 (N_9101,N_8568,N_8880);
and U9102 (N_9102,N_8928,N_8553);
nor U9103 (N_9103,N_8706,N_8988);
nor U9104 (N_9104,N_8586,N_8737);
and U9105 (N_9105,N_8515,N_8672);
nand U9106 (N_9106,N_8537,N_8564);
or U9107 (N_9107,N_8818,N_8952);
and U9108 (N_9108,N_8819,N_8514);
and U9109 (N_9109,N_8636,N_8724);
nand U9110 (N_9110,N_8772,N_8528);
xnor U9111 (N_9111,N_8711,N_8944);
nand U9112 (N_9112,N_8703,N_8681);
or U9113 (N_9113,N_8993,N_8647);
nand U9114 (N_9114,N_8872,N_8542);
xor U9115 (N_9115,N_8597,N_8780);
nand U9116 (N_9116,N_8921,N_8693);
xnor U9117 (N_9117,N_8967,N_8891);
xnor U9118 (N_9118,N_8680,N_8596);
nor U9119 (N_9119,N_8560,N_8574);
nor U9120 (N_9120,N_8506,N_8563);
nand U9121 (N_9121,N_8778,N_8983);
or U9122 (N_9122,N_8592,N_8704);
nand U9123 (N_9123,N_8632,N_8986);
or U9124 (N_9124,N_8859,N_8526);
xor U9125 (N_9125,N_8697,N_8720);
nand U9126 (N_9126,N_8975,N_8784);
xor U9127 (N_9127,N_8600,N_8581);
xnor U9128 (N_9128,N_8809,N_8807);
and U9129 (N_9129,N_8979,N_8554);
and U9130 (N_9130,N_8740,N_8913);
xor U9131 (N_9131,N_8973,N_8626);
xor U9132 (N_9132,N_8551,N_8714);
nor U9133 (N_9133,N_8565,N_8716);
xnor U9134 (N_9134,N_8540,N_8907);
nor U9135 (N_9135,N_8900,N_8638);
nor U9136 (N_9136,N_8833,N_8832);
xor U9137 (N_9137,N_8773,N_8661);
xor U9138 (N_9138,N_8906,N_8609);
or U9139 (N_9139,N_8687,N_8741);
xor U9140 (N_9140,N_8917,N_8791);
and U9141 (N_9141,N_8605,N_8576);
and U9142 (N_9142,N_8641,N_8774);
nand U9143 (N_9143,N_8723,N_8904);
xnor U9144 (N_9144,N_8781,N_8692);
or U9145 (N_9145,N_8941,N_8803);
nand U9146 (N_9146,N_8620,N_8876);
nand U9147 (N_9147,N_8511,N_8922);
nand U9148 (N_9148,N_8890,N_8947);
nand U9149 (N_9149,N_8676,N_8855);
or U9150 (N_9150,N_8997,N_8683);
nor U9151 (N_9151,N_8547,N_8505);
and U9152 (N_9152,N_8503,N_8602);
and U9153 (N_9153,N_8531,N_8624);
nor U9154 (N_9154,N_8544,N_8951);
or U9155 (N_9155,N_8639,N_8931);
nor U9156 (N_9156,N_8965,N_8903);
or U9157 (N_9157,N_8664,N_8970);
or U9158 (N_9158,N_8976,N_8797);
and U9159 (N_9159,N_8599,N_8878);
and U9160 (N_9160,N_8652,N_8571);
or U9161 (N_9161,N_8660,N_8823);
or U9162 (N_9162,N_8607,N_8828);
nor U9163 (N_9163,N_8561,N_8733);
nand U9164 (N_9164,N_8873,N_8735);
and U9165 (N_9165,N_8556,N_8974);
or U9166 (N_9166,N_8775,N_8918);
or U9167 (N_9167,N_8656,N_8920);
xnor U9168 (N_9168,N_8673,N_8916);
nand U9169 (N_9169,N_8548,N_8536);
or U9170 (N_9170,N_8926,N_8577);
and U9171 (N_9171,N_8987,N_8698);
and U9172 (N_9172,N_8649,N_8663);
xnor U9173 (N_9173,N_8635,N_8959);
nor U9174 (N_9174,N_8935,N_8545);
and U9175 (N_9175,N_8787,N_8617);
nand U9176 (N_9176,N_8715,N_8802);
nor U9177 (N_9177,N_8822,N_8523);
xor U9178 (N_9178,N_8902,N_8908);
or U9179 (N_9179,N_8655,N_8810);
nand U9180 (N_9180,N_8691,N_8846);
nor U9181 (N_9181,N_8650,N_8901);
nand U9182 (N_9182,N_8731,N_8707);
and U9183 (N_9183,N_8629,N_8669);
or U9184 (N_9184,N_8578,N_8747);
nand U9185 (N_9185,N_8919,N_8978);
nor U9186 (N_9186,N_8702,N_8888);
xnor U9187 (N_9187,N_8590,N_8734);
nor U9188 (N_9188,N_8753,N_8623);
nand U9189 (N_9189,N_8659,N_8513);
or U9190 (N_9190,N_8923,N_8999);
or U9191 (N_9191,N_8585,N_8767);
and U9192 (N_9192,N_8991,N_8710);
nor U9193 (N_9193,N_8682,N_8783);
xnor U9194 (N_9194,N_8984,N_8595);
and U9195 (N_9195,N_8936,N_8948);
xnor U9196 (N_9196,N_8806,N_8912);
nor U9197 (N_9197,N_8884,N_8614);
and U9198 (N_9198,N_8700,N_8929);
nor U9199 (N_9199,N_8758,N_8646);
or U9200 (N_9200,N_8868,N_8712);
nand U9201 (N_9201,N_8743,N_8895);
and U9202 (N_9202,N_8516,N_8555);
or U9203 (N_9203,N_8569,N_8535);
or U9204 (N_9204,N_8730,N_8871);
or U9205 (N_9205,N_8793,N_8862);
or U9206 (N_9206,N_8580,N_8651);
and U9207 (N_9207,N_8648,N_8662);
or U9208 (N_9208,N_8779,N_8985);
nand U9209 (N_9209,N_8738,N_8665);
xnor U9210 (N_9210,N_8744,N_8877);
xor U9211 (N_9211,N_8525,N_8792);
nor U9212 (N_9212,N_8610,N_8863);
and U9213 (N_9213,N_8519,N_8539);
xor U9214 (N_9214,N_8762,N_8853);
or U9215 (N_9215,N_8579,N_8736);
nor U9216 (N_9216,N_8601,N_8811);
nor U9217 (N_9217,N_8549,N_8584);
and U9218 (N_9218,N_8924,N_8925);
nand U9219 (N_9219,N_8507,N_8796);
and U9220 (N_9220,N_8957,N_8933);
nand U9221 (N_9221,N_8726,N_8836);
and U9222 (N_9222,N_8686,N_8618);
nand U9223 (N_9223,N_8518,N_8674);
nand U9224 (N_9224,N_8713,N_8752);
or U9225 (N_9225,N_8817,N_8729);
xnor U9226 (N_9226,N_8541,N_8690);
xnor U9227 (N_9227,N_8969,N_8847);
nor U9228 (N_9228,N_8777,N_8709);
nor U9229 (N_9229,N_8670,N_8945);
and U9230 (N_9230,N_8534,N_8845);
xor U9231 (N_9231,N_8838,N_8619);
or U9232 (N_9232,N_8589,N_8956);
and U9233 (N_9233,N_8800,N_8543);
nor U9234 (N_9234,N_8504,N_8566);
nor U9235 (N_9235,N_8658,N_8527);
nand U9236 (N_9236,N_8654,N_8940);
or U9237 (N_9237,N_8892,N_8915);
xor U9238 (N_9238,N_8530,N_8739);
xnor U9239 (N_9239,N_8725,N_8830);
xnor U9240 (N_9240,N_8866,N_8552);
or U9241 (N_9241,N_8858,N_8825);
or U9242 (N_9242,N_8794,N_8612);
nand U9243 (N_9243,N_8848,N_8509);
nor U9244 (N_9244,N_8785,N_8688);
xnor U9245 (N_9245,N_8685,N_8675);
and U9246 (N_9246,N_8699,N_8814);
nor U9247 (N_9247,N_8746,N_8732);
nor U9248 (N_9248,N_8613,N_8745);
and U9249 (N_9249,N_8883,N_8573);
and U9250 (N_9250,N_8618,N_8601);
nand U9251 (N_9251,N_8887,N_8854);
nor U9252 (N_9252,N_8899,N_8613);
and U9253 (N_9253,N_8719,N_8699);
nor U9254 (N_9254,N_8603,N_8581);
or U9255 (N_9255,N_8603,N_8988);
xor U9256 (N_9256,N_8640,N_8516);
xnor U9257 (N_9257,N_8680,N_8531);
nor U9258 (N_9258,N_8722,N_8860);
and U9259 (N_9259,N_8904,N_8695);
nand U9260 (N_9260,N_8805,N_8713);
or U9261 (N_9261,N_8661,N_8889);
or U9262 (N_9262,N_8662,N_8723);
or U9263 (N_9263,N_8697,N_8522);
xnor U9264 (N_9264,N_8920,N_8548);
and U9265 (N_9265,N_8982,N_8580);
and U9266 (N_9266,N_8721,N_8800);
xnor U9267 (N_9267,N_8859,N_8776);
or U9268 (N_9268,N_8752,N_8701);
or U9269 (N_9269,N_8937,N_8509);
nor U9270 (N_9270,N_8832,N_8607);
nor U9271 (N_9271,N_8669,N_8630);
xnor U9272 (N_9272,N_8849,N_8973);
nand U9273 (N_9273,N_8933,N_8517);
xnor U9274 (N_9274,N_8870,N_8529);
nand U9275 (N_9275,N_8744,N_8819);
nand U9276 (N_9276,N_8530,N_8763);
nor U9277 (N_9277,N_8545,N_8812);
nand U9278 (N_9278,N_8722,N_8790);
nand U9279 (N_9279,N_8582,N_8687);
or U9280 (N_9280,N_8694,N_8955);
nand U9281 (N_9281,N_8613,N_8857);
xnor U9282 (N_9282,N_8869,N_8599);
or U9283 (N_9283,N_8510,N_8621);
nand U9284 (N_9284,N_8803,N_8828);
or U9285 (N_9285,N_8891,N_8608);
and U9286 (N_9286,N_8922,N_8646);
xor U9287 (N_9287,N_8664,N_8859);
and U9288 (N_9288,N_8785,N_8508);
nor U9289 (N_9289,N_8711,N_8508);
nand U9290 (N_9290,N_8688,N_8663);
nand U9291 (N_9291,N_8789,N_8505);
xor U9292 (N_9292,N_8514,N_8751);
and U9293 (N_9293,N_8712,N_8627);
nand U9294 (N_9294,N_8855,N_8568);
nand U9295 (N_9295,N_8946,N_8745);
nor U9296 (N_9296,N_8607,N_8530);
xnor U9297 (N_9297,N_8641,N_8877);
and U9298 (N_9298,N_8632,N_8770);
or U9299 (N_9299,N_8711,N_8651);
or U9300 (N_9300,N_8932,N_8653);
or U9301 (N_9301,N_8578,N_8611);
and U9302 (N_9302,N_8917,N_8832);
nor U9303 (N_9303,N_8927,N_8966);
or U9304 (N_9304,N_8670,N_8791);
xor U9305 (N_9305,N_8827,N_8503);
nand U9306 (N_9306,N_8649,N_8535);
xor U9307 (N_9307,N_8844,N_8580);
and U9308 (N_9308,N_8938,N_8540);
nand U9309 (N_9309,N_8635,N_8506);
nand U9310 (N_9310,N_8981,N_8852);
or U9311 (N_9311,N_8850,N_8721);
nand U9312 (N_9312,N_8657,N_8599);
xnor U9313 (N_9313,N_8699,N_8769);
or U9314 (N_9314,N_8578,N_8518);
or U9315 (N_9315,N_8582,N_8501);
and U9316 (N_9316,N_8997,N_8954);
or U9317 (N_9317,N_8934,N_8636);
nand U9318 (N_9318,N_8551,N_8639);
nor U9319 (N_9319,N_8957,N_8646);
nor U9320 (N_9320,N_8615,N_8567);
nand U9321 (N_9321,N_8772,N_8641);
xnor U9322 (N_9322,N_8990,N_8592);
nand U9323 (N_9323,N_8766,N_8505);
or U9324 (N_9324,N_8979,N_8941);
and U9325 (N_9325,N_8718,N_8534);
xnor U9326 (N_9326,N_8734,N_8522);
or U9327 (N_9327,N_8762,N_8531);
and U9328 (N_9328,N_8692,N_8578);
or U9329 (N_9329,N_8528,N_8650);
or U9330 (N_9330,N_8909,N_8758);
and U9331 (N_9331,N_8577,N_8854);
xor U9332 (N_9332,N_8782,N_8885);
nor U9333 (N_9333,N_8858,N_8616);
nand U9334 (N_9334,N_8565,N_8691);
nor U9335 (N_9335,N_8735,N_8747);
xnor U9336 (N_9336,N_8712,N_8964);
nor U9337 (N_9337,N_8838,N_8690);
or U9338 (N_9338,N_8625,N_8852);
xnor U9339 (N_9339,N_8597,N_8954);
or U9340 (N_9340,N_8521,N_8629);
and U9341 (N_9341,N_8710,N_8603);
or U9342 (N_9342,N_8502,N_8683);
and U9343 (N_9343,N_8523,N_8816);
nor U9344 (N_9344,N_8500,N_8580);
or U9345 (N_9345,N_8626,N_8586);
nor U9346 (N_9346,N_8668,N_8580);
xor U9347 (N_9347,N_8676,N_8766);
nor U9348 (N_9348,N_8851,N_8608);
nand U9349 (N_9349,N_8928,N_8754);
nand U9350 (N_9350,N_8950,N_8972);
nand U9351 (N_9351,N_8650,N_8607);
and U9352 (N_9352,N_8547,N_8822);
xor U9353 (N_9353,N_8825,N_8527);
or U9354 (N_9354,N_8837,N_8697);
nor U9355 (N_9355,N_8829,N_8644);
nor U9356 (N_9356,N_8937,N_8751);
and U9357 (N_9357,N_8765,N_8636);
nor U9358 (N_9358,N_8627,N_8634);
and U9359 (N_9359,N_8598,N_8680);
nand U9360 (N_9360,N_8649,N_8851);
and U9361 (N_9361,N_8947,N_8606);
xnor U9362 (N_9362,N_8506,N_8671);
or U9363 (N_9363,N_8534,N_8795);
and U9364 (N_9364,N_8520,N_8556);
xnor U9365 (N_9365,N_8591,N_8767);
xnor U9366 (N_9366,N_8630,N_8798);
nand U9367 (N_9367,N_8922,N_8972);
or U9368 (N_9368,N_8627,N_8592);
nand U9369 (N_9369,N_8603,N_8973);
xor U9370 (N_9370,N_8636,N_8606);
nand U9371 (N_9371,N_8537,N_8805);
and U9372 (N_9372,N_8979,N_8879);
and U9373 (N_9373,N_8902,N_8736);
and U9374 (N_9374,N_8898,N_8806);
xor U9375 (N_9375,N_8541,N_8564);
and U9376 (N_9376,N_8898,N_8576);
nand U9377 (N_9377,N_8768,N_8765);
and U9378 (N_9378,N_8961,N_8928);
or U9379 (N_9379,N_8717,N_8924);
nand U9380 (N_9380,N_8851,N_8630);
nor U9381 (N_9381,N_8702,N_8900);
nor U9382 (N_9382,N_8987,N_8749);
or U9383 (N_9383,N_8714,N_8778);
nor U9384 (N_9384,N_8599,N_8553);
or U9385 (N_9385,N_8602,N_8950);
nor U9386 (N_9386,N_8970,N_8685);
or U9387 (N_9387,N_8772,N_8764);
and U9388 (N_9388,N_8905,N_8531);
nand U9389 (N_9389,N_8641,N_8795);
or U9390 (N_9390,N_8515,N_8658);
or U9391 (N_9391,N_8550,N_8987);
and U9392 (N_9392,N_8964,N_8737);
nor U9393 (N_9393,N_8838,N_8934);
nand U9394 (N_9394,N_8879,N_8831);
or U9395 (N_9395,N_8842,N_8582);
xnor U9396 (N_9396,N_8706,N_8845);
and U9397 (N_9397,N_8716,N_8880);
nor U9398 (N_9398,N_8838,N_8843);
nand U9399 (N_9399,N_8588,N_8728);
xnor U9400 (N_9400,N_8564,N_8716);
and U9401 (N_9401,N_8822,N_8791);
xor U9402 (N_9402,N_8943,N_8603);
nand U9403 (N_9403,N_8824,N_8760);
or U9404 (N_9404,N_8747,N_8701);
or U9405 (N_9405,N_8782,N_8986);
or U9406 (N_9406,N_8931,N_8581);
and U9407 (N_9407,N_8826,N_8544);
nor U9408 (N_9408,N_8602,N_8676);
and U9409 (N_9409,N_8941,N_8806);
or U9410 (N_9410,N_8826,N_8792);
or U9411 (N_9411,N_8685,N_8763);
and U9412 (N_9412,N_8569,N_8500);
and U9413 (N_9413,N_8809,N_8566);
xnor U9414 (N_9414,N_8952,N_8876);
xnor U9415 (N_9415,N_8525,N_8981);
and U9416 (N_9416,N_8829,N_8903);
and U9417 (N_9417,N_8774,N_8948);
or U9418 (N_9418,N_8971,N_8515);
nand U9419 (N_9419,N_8712,N_8756);
nor U9420 (N_9420,N_8657,N_8574);
nor U9421 (N_9421,N_8832,N_8868);
nor U9422 (N_9422,N_8713,N_8579);
nor U9423 (N_9423,N_8623,N_8605);
or U9424 (N_9424,N_8737,N_8805);
and U9425 (N_9425,N_8643,N_8722);
nor U9426 (N_9426,N_8747,N_8810);
nor U9427 (N_9427,N_8597,N_8708);
or U9428 (N_9428,N_8911,N_8673);
xor U9429 (N_9429,N_8727,N_8958);
and U9430 (N_9430,N_8540,N_8904);
xnor U9431 (N_9431,N_8748,N_8725);
or U9432 (N_9432,N_8868,N_8871);
or U9433 (N_9433,N_8646,N_8530);
xor U9434 (N_9434,N_8787,N_8896);
and U9435 (N_9435,N_8512,N_8922);
or U9436 (N_9436,N_8659,N_8728);
nand U9437 (N_9437,N_8993,N_8686);
and U9438 (N_9438,N_8759,N_8692);
nor U9439 (N_9439,N_8907,N_8519);
nor U9440 (N_9440,N_8541,N_8854);
xnor U9441 (N_9441,N_8650,N_8977);
nand U9442 (N_9442,N_8635,N_8750);
xor U9443 (N_9443,N_8713,N_8764);
nand U9444 (N_9444,N_8835,N_8947);
nor U9445 (N_9445,N_8604,N_8931);
nand U9446 (N_9446,N_8530,N_8621);
nand U9447 (N_9447,N_8581,N_8546);
and U9448 (N_9448,N_8877,N_8779);
and U9449 (N_9449,N_8630,N_8943);
or U9450 (N_9450,N_8965,N_8541);
or U9451 (N_9451,N_8630,N_8706);
nand U9452 (N_9452,N_8609,N_8954);
nand U9453 (N_9453,N_8930,N_8899);
xor U9454 (N_9454,N_8804,N_8840);
xor U9455 (N_9455,N_8890,N_8592);
nand U9456 (N_9456,N_8604,N_8539);
or U9457 (N_9457,N_8967,N_8570);
nand U9458 (N_9458,N_8742,N_8818);
xnor U9459 (N_9459,N_8512,N_8961);
nand U9460 (N_9460,N_8746,N_8999);
and U9461 (N_9461,N_8901,N_8508);
xnor U9462 (N_9462,N_8696,N_8814);
nand U9463 (N_9463,N_8982,N_8578);
nand U9464 (N_9464,N_8756,N_8587);
nand U9465 (N_9465,N_8964,N_8894);
and U9466 (N_9466,N_8649,N_8591);
nand U9467 (N_9467,N_8796,N_8916);
and U9468 (N_9468,N_8977,N_8794);
xnor U9469 (N_9469,N_8697,N_8727);
nand U9470 (N_9470,N_8668,N_8854);
or U9471 (N_9471,N_8718,N_8852);
nand U9472 (N_9472,N_8901,N_8863);
nand U9473 (N_9473,N_8833,N_8917);
nor U9474 (N_9474,N_8636,N_8668);
nand U9475 (N_9475,N_8680,N_8684);
and U9476 (N_9476,N_8719,N_8813);
nor U9477 (N_9477,N_8511,N_8823);
xor U9478 (N_9478,N_8744,N_8850);
nor U9479 (N_9479,N_8881,N_8684);
or U9480 (N_9480,N_8626,N_8763);
xnor U9481 (N_9481,N_8919,N_8917);
xor U9482 (N_9482,N_8851,N_8663);
nand U9483 (N_9483,N_8549,N_8835);
xnor U9484 (N_9484,N_8519,N_8601);
and U9485 (N_9485,N_8790,N_8714);
nor U9486 (N_9486,N_8933,N_8902);
nor U9487 (N_9487,N_8984,N_8961);
nand U9488 (N_9488,N_8558,N_8932);
xor U9489 (N_9489,N_8503,N_8730);
nor U9490 (N_9490,N_8500,N_8598);
or U9491 (N_9491,N_8714,N_8792);
nor U9492 (N_9492,N_8626,N_8854);
nand U9493 (N_9493,N_8763,N_8709);
and U9494 (N_9494,N_8831,N_8843);
or U9495 (N_9495,N_8664,N_8526);
xnor U9496 (N_9496,N_8512,N_8851);
nand U9497 (N_9497,N_8938,N_8720);
and U9498 (N_9498,N_8770,N_8953);
or U9499 (N_9499,N_8949,N_8618);
nand U9500 (N_9500,N_9199,N_9339);
xnor U9501 (N_9501,N_9308,N_9261);
nand U9502 (N_9502,N_9220,N_9324);
nand U9503 (N_9503,N_9163,N_9457);
nor U9504 (N_9504,N_9254,N_9147);
or U9505 (N_9505,N_9104,N_9140);
and U9506 (N_9506,N_9371,N_9159);
or U9507 (N_9507,N_9200,N_9029);
nand U9508 (N_9508,N_9243,N_9436);
xor U9509 (N_9509,N_9479,N_9024);
and U9510 (N_9510,N_9343,N_9111);
nor U9511 (N_9511,N_9284,N_9233);
and U9512 (N_9512,N_9062,N_9287);
nand U9513 (N_9513,N_9161,N_9172);
xor U9514 (N_9514,N_9450,N_9336);
xor U9515 (N_9515,N_9453,N_9196);
nand U9516 (N_9516,N_9474,N_9411);
nand U9517 (N_9517,N_9098,N_9441);
xor U9518 (N_9518,N_9311,N_9244);
nor U9519 (N_9519,N_9019,N_9301);
nor U9520 (N_9520,N_9241,N_9485);
nand U9521 (N_9521,N_9471,N_9025);
nand U9522 (N_9522,N_9362,N_9443);
and U9523 (N_9523,N_9483,N_9387);
nor U9524 (N_9524,N_9177,N_9340);
nor U9525 (N_9525,N_9020,N_9073);
and U9526 (N_9526,N_9419,N_9191);
or U9527 (N_9527,N_9128,N_9089);
nor U9528 (N_9528,N_9169,N_9412);
nor U9529 (N_9529,N_9065,N_9226);
or U9530 (N_9530,N_9344,N_9268);
or U9531 (N_9531,N_9396,N_9469);
or U9532 (N_9532,N_9363,N_9290);
or U9533 (N_9533,N_9366,N_9302);
xnor U9534 (N_9534,N_9101,N_9151);
xor U9535 (N_9535,N_9206,N_9462);
nor U9536 (N_9536,N_9381,N_9224);
or U9537 (N_9537,N_9262,N_9179);
nand U9538 (N_9538,N_9049,N_9145);
or U9539 (N_9539,N_9021,N_9058);
or U9540 (N_9540,N_9251,N_9373);
nand U9541 (N_9541,N_9495,N_9006);
or U9542 (N_9542,N_9463,N_9153);
xor U9543 (N_9543,N_9245,N_9467);
and U9544 (N_9544,N_9274,N_9064);
nor U9545 (N_9545,N_9361,N_9040);
nor U9546 (N_9546,N_9491,N_9292);
xor U9547 (N_9547,N_9442,N_9042);
xnor U9548 (N_9548,N_9368,N_9134);
or U9549 (N_9549,N_9498,N_9273);
nand U9550 (N_9550,N_9236,N_9078);
nor U9551 (N_9551,N_9326,N_9263);
or U9552 (N_9552,N_9090,N_9416);
nor U9553 (N_9553,N_9372,N_9219);
nand U9554 (N_9554,N_9031,N_9212);
and U9555 (N_9555,N_9297,N_9286);
and U9556 (N_9556,N_9332,N_9192);
or U9557 (N_9557,N_9247,N_9097);
xor U9558 (N_9558,N_9223,N_9237);
nor U9559 (N_9559,N_9185,N_9448);
xnor U9560 (N_9560,N_9328,N_9060);
or U9561 (N_9561,N_9231,N_9075);
nand U9562 (N_9562,N_9080,N_9168);
nor U9563 (N_9563,N_9367,N_9335);
nor U9564 (N_9564,N_9385,N_9136);
nand U9565 (N_9565,N_9176,N_9155);
nor U9566 (N_9566,N_9234,N_9208);
or U9567 (N_9567,N_9026,N_9313);
xor U9568 (N_9568,N_9480,N_9316);
xnor U9569 (N_9569,N_9496,N_9468);
nor U9570 (N_9570,N_9053,N_9426);
nand U9571 (N_9571,N_9085,N_9227);
or U9572 (N_9572,N_9482,N_9310);
nand U9573 (N_9573,N_9460,N_9158);
or U9574 (N_9574,N_9207,N_9276);
nand U9575 (N_9575,N_9407,N_9116);
nand U9576 (N_9576,N_9125,N_9280);
and U9577 (N_9577,N_9182,N_9121);
nand U9578 (N_9578,N_9183,N_9391);
and U9579 (N_9579,N_9322,N_9144);
nor U9580 (N_9580,N_9204,N_9214);
and U9581 (N_9581,N_9187,N_9497);
nor U9582 (N_9582,N_9341,N_9492);
nor U9583 (N_9583,N_9392,N_9403);
xnor U9584 (N_9584,N_9431,N_9257);
and U9585 (N_9585,N_9092,N_9052);
and U9586 (N_9586,N_9033,N_9171);
or U9587 (N_9587,N_9410,N_9493);
or U9588 (N_9588,N_9013,N_9478);
and U9589 (N_9589,N_9300,N_9365);
nand U9590 (N_9590,N_9272,N_9386);
and U9591 (N_9591,N_9056,N_9393);
nand U9592 (N_9592,N_9235,N_9432);
xor U9593 (N_9593,N_9279,N_9112);
or U9594 (N_9594,N_9138,N_9150);
nand U9595 (N_9595,N_9399,N_9294);
xor U9596 (N_9596,N_9016,N_9014);
xor U9597 (N_9597,N_9439,N_9041);
and U9598 (N_9598,N_9127,N_9414);
nand U9599 (N_9599,N_9427,N_9059);
xnor U9600 (N_9600,N_9430,N_9417);
xor U9601 (N_9601,N_9380,N_9413);
nand U9602 (N_9602,N_9022,N_9337);
nand U9603 (N_9603,N_9018,N_9260);
xor U9604 (N_9604,N_9131,N_9083);
nand U9605 (N_9605,N_9036,N_9066);
or U9606 (N_9606,N_9353,N_9255);
or U9607 (N_9607,N_9135,N_9312);
nand U9608 (N_9608,N_9259,N_9109);
nor U9609 (N_9609,N_9215,N_9074);
and U9610 (N_9610,N_9338,N_9425);
nand U9611 (N_9611,N_9428,N_9376);
nor U9612 (N_9612,N_9379,N_9293);
nand U9613 (N_9613,N_9253,N_9008);
xor U9614 (N_9614,N_9117,N_9000);
xor U9615 (N_9615,N_9050,N_9331);
and U9616 (N_9616,N_9067,N_9106);
nor U9617 (N_9617,N_9068,N_9299);
or U9618 (N_9618,N_9242,N_9445);
xor U9619 (N_9619,N_9063,N_9461);
nor U9620 (N_9620,N_9222,N_9239);
and U9621 (N_9621,N_9283,N_9473);
xnor U9622 (N_9622,N_9091,N_9354);
and U9623 (N_9623,N_9180,N_9001);
or U9624 (N_9624,N_9270,N_9321);
xnor U9625 (N_9625,N_9046,N_9295);
nand U9626 (N_9626,N_9499,N_9422);
nor U9627 (N_9627,N_9108,N_9434);
and U9628 (N_9628,N_9438,N_9437);
nand U9629 (N_9629,N_9477,N_9099);
and U9630 (N_9630,N_9077,N_9095);
or U9631 (N_9631,N_9384,N_9277);
xor U9632 (N_9632,N_9408,N_9045);
nand U9633 (N_9633,N_9105,N_9079);
and U9634 (N_9634,N_9023,N_9174);
and U9635 (N_9635,N_9015,N_9149);
nor U9636 (N_9636,N_9325,N_9130);
and U9637 (N_9637,N_9012,N_9435);
xor U9638 (N_9638,N_9160,N_9458);
nand U9639 (N_9639,N_9173,N_9210);
nor U9640 (N_9640,N_9446,N_9114);
nand U9641 (N_9641,N_9027,N_9146);
nand U9642 (N_9642,N_9348,N_9143);
and U9643 (N_9643,N_9488,N_9303);
xnor U9644 (N_9644,N_9394,N_9118);
nor U9645 (N_9645,N_9203,N_9329);
and U9646 (N_9646,N_9154,N_9010);
and U9647 (N_9647,N_9288,N_9454);
or U9648 (N_9648,N_9323,N_9047);
nand U9649 (N_9649,N_9070,N_9320);
and U9650 (N_9650,N_9390,N_9489);
xnor U9651 (N_9651,N_9102,N_9017);
nand U9652 (N_9652,N_9175,N_9358);
or U9653 (N_9653,N_9342,N_9370);
and U9654 (N_9654,N_9197,N_9304);
xnor U9655 (N_9655,N_9028,N_9038);
or U9656 (N_9656,N_9406,N_9418);
and U9657 (N_9657,N_9334,N_9123);
or U9658 (N_9658,N_9126,N_9318);
xnor U9659 (N_9659,N_9377,N_9181);
nor U9660 (N_9660,N_9481,N_9347);
nand U9661 (N_9661,N_9039,N_9087);
and U9662 (N_9662,N_9395,N_9195);
or U9663 (N_9663,N_9319,N_9405);
xnor U9664 (N_9664,N_9475,N_9166);
nand U9665 (N_9665,N_9107,N_9375);
nand U9666 (N_9666,N_9397,N_9082);
nor U9667 (N_9667,N_9081,N_9465);
or U9668 (N_9668,N_9148,N_9178);
xor U9669 (N_9669,N_9352,N_9061);
nand U9670 (N_9670,N_9258,N_9186);
xor U9671 (N_9671,N_9267,N_9289);
xor U9672 (N_9672,N_9364,N_9216);
nor U9673 (N_9673,N_9240,N_9249);
nor U9674 (N_9674,N_9421,N_9048);
xor U9675 (N_9675,N_9369,N_9142);
nor U9676 (N_9676,N_9494,N_9137);
or U9677 (N_9677,N_9266,N_9165);
xor U9678 (N_9678,N_9189,N_9346);
and U9679 (N_9679,N_9487,N_9423);
and U9680 (N_9680,N_9198,N_9246);
nor U9681 (N_9681,N_9269,N_9383);
or U9682 (N_9682,N_9472,N_9201);
or U9683 (N_9683,N_9094,N_9409);
nor U9684 (N_9684,N_9456,N_9141);
and U9685 (N_9685,N_9398,N_9072);
xnor U9686 (N_9686,N_9188,N_9205);
nand U9687 (N_9687,N_9429,N_9209);
nor U9688 (N_9688,N_9228,N_9132);
nor U9689 (N_9689,N_9032,N_9184);
xnor U9690 (N_9690,N_9349,N_9330);
or U9691 (N_9691,N_9096,N_9424);
nand U9692 (N_9692,N_9248,N_9011);
nand U9693 (N_9693,N_9167,N_9110);
xor U9694 (N_9694,N_9069,N_9315);
or U9695 (N_9695,N_9221,N_9057);
xnor U9696 (N_9696,N_9129,N_9004);
nor U9697 (N_9697,N_9113,N_9314);
or U9698 (N_9698,N_9005,N_9281);
or U9699 (N_9699,N_9402,N_9256);
and U9700 (N_9700,N_9211,N_9238);
and U9701 (N_9701,N_9415,N_9275);
nor U9702 (N_9702,N_9213,N_9164);
nor U9703 (N_9703,N_9307,N_9030);
nor U9704 (N_9704,N_9282,N_9190);
xor U9705 (N_9705,N_9265,N_9252);
and U9706 (N_9706,N_9007,N_9202);
or U9707 (N_9707,N_9194,N_9250);
nor U9708 (N_9708,N_9037,N_9378);
xor U9709 (N_9709,N_9309,N_9139);
and U9710 (N_9710,N_9088,N_9333);
nand U9711 (N_9711,N_9388,N_9133);
xnor U9712 (N_9712,N_9317,N_9296);
or U9713 (N_9713,N_9447,N_9470);
xor U9714 (N_9714,N_9124,N_9459);
and U9715 (N_9715,N_9420,N_9306);
and U9716 (N_9716,N_9076,N_9476);
nor U9717 (N_9717,N_9484,N_9156);
nor U9718 (N_9718,N_9086,N_9452);
or U9719 (N_9719,N_9400,N_9298);
or U9720 (N_9720,N_9291,N_9103);
nor U9721 (N_9721,N_9119,N_9225);
nor U9722 (N_9722,N_9217,N_9327);
xor U9723 (N_9723,N_9218,N_9451);
xor U9724 (N_9724,N_9389,N_9120);
nand U9725 (N_9725,N_9229,N_9374);
nor U9726 (N_9726,N_9464,N_9486);
xor U9727 (N_9727,N_9271,N_9232);
or U9728 (N_9728,N_9034,N_9264);
nand U9729 (N_9729,N_9044,N_9157);
nor U9730 (N_9730,N_9285,N_9003);
xnor U9731 (N_9731,N_9278,N_9345);
or U9732 (N_9732,N_9404,N_9035);
nand U9733 (N_9733,N_9043,N_9122);
xnor U9734 (N_9734,N_9444,N_9162);
nand U9735 (N_9735,N_9009,N_9359);
xor U9736 (N_9736,N_9152,N_9305);
nand U9737 (N_9737,N_9382,N_9230);
nand U9738 (N_9738,N_9449,N_9055);
and U9739 (N_9739,N_9466,N_9433);
or U9740 (N_9740,N_9360,N_9355);
or U9741 (N_9741,N_9002,N_9401);
and U9742 (N_9742,N_9356,N_9100);
or U9743 (N_9743,N_9093,N_9071);
nand U9744 (N_9744,N_9351,N_9350);
nand U9745 (N_9745,N_9115,N_9357);
xnor U9746 (N_9746,N_9054,N_9051);
nand U9747 (N_9747,N_9170,N_9193);
and U9748 (N_9748,N_9455,N_9440);
nand U9749 (N_9749,N_9490,N_9084);
and U9750 (N_9750,N_9319,N_9221);
or U9751 (N_9751,N_9280,N_9114);
and U9752 (N_9752,N_9446,N_9052);
or U9753 (N_9753,N_9440,N_9412);
or U9754 (N_9754,N_9391,N_9174);
xor U9755 (N_9755,N_9135,N_9072);
or U9756 (N_9756,N_9238,N_9300);
nor U9757 (N_9757,N_9368,N_9132);
nor U9758 (N_9758,N_9007,N_9402);
nor U9759 (N_9759,N_9392,N_9481);
xnor U9760 (N_9760,N_9087,N_9349);
nor U9761 (N_9761,N_9259,N_9473);
and U9762 (N_9762,N_9466,N_9112);
xor U9763 (N_9763,N_9032,N_9079);
nand U9764 (N_9764,N_9169,N_9088);
and U9765 (N_9765,N_9090,N_9420);
or U9766 (N_9766,N_9196,N_9127);
and U9767 (N_9767,N_9013,N_9467);
xor U9768 (N_9768,N_9271,N_9005);
nor U9769 (N_9769,N_9018,N_9001);
nor U9770 (N_9770,N_9116,N_9064);
and U9771 (N_9771,N_9179,N_9494);
nand U9772 (N_9772,N_9009,N_9044);
or U9773 (N_9773,N_9454,N_9250);
nor U9774 (N_9774,N_9230,N_9239);
xnor U9775 (N_9775,N_9099,N_9066);
nand U9776 (N_9776,N_9478,N_9030);
xnor U9777 (N_9777,N_9168,N_9315);
nor U9778 (N_9778,N_9208,N_9056);
nand U9779 (N_9779,N_9456,N_9396);
nand U9780 (N_9780,N_9416,N_9245);
nand U9781 (N_9781,N_9481,N_9273);
nor U9782 (N_9782,N_9156,N_9257);
nand U9783 (N_9783,N_9149,N_9044);
nand U9784 (N_9784,N_9323,N_9108);
and U9785 (N_9785,N_9408,N_9200);
or U9786 (N_9786,N_9207,N_9456);
xnor U9787 (N_9787,N_9121,N_9333);
nand U9788 (N_9788,N_9310,N_9194);
xor U9789 (N_9789,N_9087,N_9460);
and U9790 (N_9790,N_9493,N_9409);
or U9791 (N_9791,N_9383,N_9032);
nor U9792 (N_9792,N_9470,N_9298);
xnor U9793 (N_9793,N_9140,N_9116);
or U9794 (N_9794,N_9350,N_9062);
nor U9795 (N_9795,N_9224,N_9310);
or U9796 (N_9796,N_9454,N_9194);
xor U9797 (N_9797,N_9138,N_9227);
and U9798 (N_9798,N_9025,N_9435);
or U9799 (N_9799,N_9437,N_9026);
or U9800 (N_9800,N_9416,N_9360);
or U9801 (N_9801,N_9156,N_9314);
or U9802 (N_9802,N_9218,N_9421);
and U9803 (N_9803,N_9377,N_9374);
nor U9804 (N_9804,N_9474,N_9214);
nor U9805 (N_9805,N_9221,N_9022);
or U9806 (N_9806,N_9267,N_9217);
or U9807 (N_9807,N_9175,N_9030);
nor U9808 (N_9808,N_9455,N_9436);
or U9809 (N_9809,N_9040,N_9192);
nand U9810 (N_9810,N_9169,N_9462);
nand U9811 (N_9811,N_9170,N_9177);
nand U9812 (N_9812,N_9172,N_9462);
or U9813 (N_9813,N_9041,N_9405);
nand U9814 (N_9814,N_9004,N_9076);
xnor U9815 (N_9815,N_9343,N_9220);
and U9816 (N_9816,N_9290,N_9355);
nand U9817 (N_9817,N_9366,N_9485);
xnor U9818 (N_9818,N_9398,N_9285);
and U9819 (N_9819,N_9224,N_9364);
nor U9820 (N_9820,N_9011,N_9343);
nor U9821 (N_9821,N_9293,N_9455);
nand U9822 (N_9822,N_9436,N_9440);
or U9823 (N_9823,N_9475,N_9171);
and U9824 (N_9824,N_9331,N_9231);
nand U9825 (N_9825,N_9303,N_9410);
nand U9826 (N_9826,N_9210,N_9063);
and U9827 (N_9827,N_9202,N_9424);
or U9828 (N_9828,N_9441,N_9479);
or U9829 (N_9829,N_9147,N_9134);
and U9830 (N_9830,N_9219,N_9350);
nand U9831 (N_9831,N_9423,N_9146);
and U9832 (N_9832,N_9296,N_9262);
or U9833 (N_9833,N_9257,N_9354);
and U9834 (N_9834,N_9185,N_9180);
nand U9835 (N_9835,N_9010,N_9194);
nand U9836 (N_9836,N_9472,N_9058);
xor U9837 (N_9837,N_9343,N_9416);
nand U9838 (N_9838,N_9031,N_9049);
or U9839 (N_9839,N_9314,N_9403);
nor U9840 (N_9840,N_9397,N_9189);
and U9841 (N_9841,N_9136,N_9347);
nor U9842 (N_9842,N_9066,N_9382);
or U9843 (N_9843,N_9100,N_9268);
or U9844 (N_9844,N_9273,N_9085);
and U9845 (N_9845,N_9304,N_9109);
or U9846 (N_9846,N_9006,N_9090);
and U9847 (N_9847,N_9480,N_9210);
nor U9848 (N_9848,N_9223,N_9012);
nor U9849 (N_9849,N_9172,N_9091);
nand U9850 (N_9850,N_9200,N_9285);
xnor U9851 (N_9851,N_9228,N_9315);
nor U9852 (N_9852,N_9342,N_9071);
nand U9853 (N_9853,N_9326,N_9173);
and U9854 (N_9854,N_9087,N_9103);
nor U9855 (N_9855,N_9354,N_9202);
and U9856 (N_9856,N_9423,N_9181);
xnor U9857 (N_9857,N_9188,N_9085);
or U9858 (N_9858,N_9178,N_9288);
nor U9859 (N_9859,N_9058,N_9417);
nor U9860 (N_9860,N_9382,N_9182);
or U9861 (N_9861,N_9121,N_9082);
and U9862 (N_9862,N_9152,N_9344);
xnor U9863 (N_9863,N_9023,N_9216);
and U9864 (N_9864,N_9317,N_9251);
nand U9865 (N_9865,N_9361,N_9310);
xnor U9866 (N_9866,N_9035,N_9349);
nand U9867 (N_9867,N_9006,N_9060);
nand U9868 (N_9868,N_9133,N_9261);
nor U9869 (N_9869,N_9143,N_9474);
nor U9870 (N_9870,N_9186,N_9328);
xor U9871 (N_9871,N_9415,N_9029);
nand U9872 (N_9872,N_9150,N_9145);
nand U9873 (N_9873,N_9297,N_9436);
nor U9874 (N_9874,N_9276,N_9308);
nand U9875 (N_9875,N_9496,N_9032);
nand U9876 (N_9876,N_9139,N_9244);
and U9877 (N_9877,N_9176,N_9346);
nor U9878 (N_9878,N_9337,N_9152);
xor U9879 (N_9879,N_9312,N_9116);
or U9880 (N_9880,N_9472,N_9431);
nand U9881 (N_9881,N_9436,N_9474);
nand U9882 (N_9882,N_9293,N_9172);
nor U9883 (N_9883,N_9172,N_9126);
or U9884 (N_9884,N_9342,N_9114);
nand U9885 (N_9885,N_9016,N_9002);
xor U9886 (N_9886,N_9497,N_9147);
or U9887 (N_9887,N_9111,N_9148);
nor U9888 (N_9888,N_9089,N_9013);
or U9889 (N_9889,N_9327,N_9174);
and U9890 (N_9890,N_9096,N_9213);
nand U9891 (N_9891,N_9347,N_9183);
xnor U9892 (N_9892,N_9409,N_9403);
xor U9893 (N_9893,N_9380,N_9369);
or U9894 (N_9894,N_9291,N_9381);
and U9895 (N_9895,N_9475,N_9117);
xnor U9896 (N_9896,N_9126,N_9419);
nand U9897 (N_9897,N_9395,N_9259);
nor U9898 (N_9898,N_9498,N_9000);
and U9899 (N_9899,N_9256,N_9232);
xor U9900 (N_9900,N_9285,N_9441);
xor U9901 (N_9901,N_9066,N_9037);
nor U9902 (N_9902,N_9472,N_9483);
or U9903 (N_9903,N_9026,N_9363);
nand U9904 (N_9904,N_9465,N_9263);
nand U9905 (N_9905,N_9469,N_9492);
nand U9906 (N_9906,N_9249,N_9436);
or U9907 (N_9907,N_9137,N_9280);
nor U9908 (N_9908,N_9474,N_9180);
nand U9909 (N_9909,N_9244,N_9354);
and U9910 (N_9910,N_9239,N_9313);
nor U9911 (N_9911,N_9052,N_9046);
xnor U9912 (N_9912,N_9421,N_9348);
or U9913 (N_9913,N_9266,N_9399);
nand U9914 (N_9914,N_9464,N_9380);
or U9915 (N_9915,N_9250,N_9247);
nand U9916 (N_9916,N_9433,N_9075);
xnor U9917 (N_9917,N_9181,N_9235);
nand U9918 (N_9918,N_9251,N_9481);
nor U9919 (N_9919,N_9412,N_9076);
nor U9920 (N_9920,N_9393,N_9476);
or U9921 (N_9921,N_9113,N_9016);
or U9922 (N_9922,N_9090,N_9246);
xor U9923 (N_9923,N_9149,N_9217);
xnor U9924 (N_9924,N_9330,N_9177);
nand U9925 (N_9925,N_9144,N_9362);
and U9926 (N_9926,N_9108,N_9079);
nand U9927 (N_9927,N_9123,N_9213);
and U9928 (N_9928,N_9279,N_9153);
nor U9929 (N_9929,N_9431,N_9224);
and U9930 (N_9930,N_9334,N_9130);
xnor U9931 (N_9931,N_9279,N_9045);
nor U9932 (N_9932,N_9265,N_9422);
and U9933 (N_9933,N_9059,N_9242);
or U9934 (N_9934,N_9113,N_9033);
nand U9935 (N_9935,N_9182,N_9343);
and U9936 (N_9936,N_9092,N_9118);
nor U9937 (N_9937,N_9496,N_9491);
nand U9938 (N_9938,N_9132,N_9112);
xor U9939 (N_9939,N_9236,N_9448);
nor U9940 (N_9940,N_9463,N_9115);
and U9941 (N_9941,N_9147,N_9108);
or U9942 (N_9942,N_9439,N_9197);
xnor U9943 (N_9943,N_9278,N_9206);
or U9944 (N_9944,N_9027,N_9283);
or U9945 (N_9945,N_9210,N_9050);
xor U9946 (N_9946,N_9334,N_9396);
or U9947 (N_9947,N_9241,N_9346);
and U9948 (N_9948,N_9491,N_9178);
and U9949 (N_9949,N_9093,N_9419);
or U9950 (N_9950,N_9009,N_9030);
or U9951 (N_9951,N_9371,N_9469);
xnor U9952 (N_9952,N_9376,N_9116);
and U9953 (N_9953,N_9156,N_9472);
and U9954 (N_9954,N_9433,N_9440);
xor U9955 (N_9955,N_9422,N_9089);
or U9956 (N_9956,N_9233,N_9125);
and U9957 (N_9957,N_9246,N_9336);
nor U9958 (N_9958,N_9417,N_9359);
or U9959 (N_9959,N_9386,N_9378);
nor U9960 (N_9960,N_9164,N_9222);
and U9961 (N_9961,N_9088,N_9349);
nand U9962 (N_9962,N_9388,N_9312);
nand U9963 (N_9963,N_9090,N_9192);
nor U9964 (N_9964,N_9289,N_9247);
nor U9965 (N_9965,N_9097,N_9105);
nand U9966 (N_9966,N_9217,N_9015);
and U9967 (N_9967,N_9120,N_9328);
and U9968 (N_9968,N_9046,N_9338);
or U9969 (N_9969,N_9288,N_9378);
nand U9970 (N_9970,N_9051,N_9478);
nor U9971 (N_9971,N_9493,N_9397);
nand U9972 (N_9972,N_9247,N_9251);
xor U9973 (N_9973,N_9374,N_9382);
or U9974 (N_9974,N_9090,N_9285);
xnor U9975 (N_9975,N_9211,N_9323);
or U9976 (N_9976,N_9249,N_9343);
nor U9977 (N_9977,N_9479,N_9373);
xor U9978 (N_9978,N_9053,N_9071);
and U9979 (N_9979,N_9341,N_9371);
xnor U9980 (N_9980,N_9073,N_9498);
nand U9981 (N_9981,N_9451,N_9228);
and U9982 (N_9982,N_9068,N_9198);
nor U9983 (N_9983,N_9283,N_9166);
xnor U9984 (N_9984,N_9173,N_9028);
and U9985 (N_9985,N_9261,N_9293);
nor U9986 (N_9986,N_9452,N_9376);
nor U9987 (N_9987,N_9140,N_9440);
nor U9988 (N_9988,N_9412,N_9285);
nand U9989 (N_9989,N_9188,N_9083);
or U9990 (N_9990,N_9141,N_9304);
xnor U9991 (N_9991,N_9155,N_9086);
and U9992 (N_9992,N_9331,N_9448);
and U9993 (N_9993,N_9231,N_9336);
nand U9994 (N_9994,N_9425,N_9223);
xor U9995 (N_9995,N_9019,N_9452);
or U9996 (N_9996,N_9472,N_9298);
nand U9997 (N_9997,N_9102,N_9444);
xnor U9998 (N_9998,N_9131,N_9493);
or U9999 (N_9999,N_9126,N_9213);
or U10000 (N_10000,N_9948,N_9986);
xor U10001 (N_10001,N_9811,N_9912);
nand U10002 (N_10002,N_9944,N_9776);
and U10003 (N_10003,N_9606,N_9706);
nor U10004 (N_10004,N_9574,N_9862);
or U10005 (N_10005,N_9741,N_9897);
xnor U10006 (N_10006,N_9530,N_9791);
and U10007 (N_10007,N_9712,N_9605);
and U10008 (N_10008,N_9683,N_9586);
or U10009 (N_10009,N_9691,N_9748);
nand U10010 (N_10010,N_9671,N_9810);
nand U10011 (N_10011,N_9511,N_9608);
xor U10012 (N_10012,N_9532,N_9611);
nand U10013 (N_10013,N_9752,N_9803);
nand U10014 (N_10014,N_9731,N_9956);
nand U10015 (N_10015,N_9729,N_9778);
nand U10016 (N_10016,N_9673,N_9755);
nand U10017 (N_10017,N_9554,N_9722);
or U10018 (N_10018,N_9587,N_9728);
nor U10019 (N_10019,N_9837,N_9550);
and U10020 (N_10020,N_9756,N_9704);
xnor U10021 (N_10021,N_9987,N_9854);
nand U10022 (N_10022,N_9982,N_9819);
nand U10023 (N_10023,N_9926,N_9537);
or U10024 (N_10024,N_9512,N_9925);
or U10025 (N_10025,N_9754,N_9820);
nor U10026 (N_10026,N_9928,N_9594);
xnor U10027 (N_10027,N_9962,N_9604);
nor U10028 (N_10028,N_9679,N_9515);
nand U10029 (N_10029,N_9898,N_9996);
xor U10030 (N_10030,N_9724,N_9792);
nor U10031 (N_10031,N_9788,N_9790);
or U10032 (N_10032,N_9868,N_9964);
nor U10033 (N_10033,N_9649,N_9975);
or U10034 (N_10034,N_9760,N_9838);
nand U10035 (N_10035,N_9509,N_9578);
nand U10036 (N_10036,N_9769,N_9805);
or U10037 (N_10037,N_9817,N_9607);
nor U10038 (N_10038,N_9840,N_9937);
xor U10039 (N_10039,N_9814,N_9800);
nor U10040 (N_10040,N_9603,N_9907);
xnor U10041 (N_10041,N_9716,N_9645);
or U10042 (N_10042,N_9892,N_9709);
and U10043 (N_10043,N_9534,N_9832);
nor U10044 (N_10044,N_9634,N_9643);
xnor U10045 (N_10045,N_9547,N_9516);
nor U10046 (N_10046,N_9508,N_9707);
nand U10047 (N_10047,N_9619,N_9886);
or U10048 (N_10048,N_9980,N_9821);
and U10049 (N_10049,N_9524,N_9797);
or U10050 (N_10050,N_9561,N_9599);
and U10051 (N_10051,N_9573,N_9879);
or U10052 (N_10052,N_9917,N_9627);
or U10053 (N_10053,N_9545,N_9654);
and U10054 (N_10054,N_9786,N_9806);
nor U10055 (N_10055,N_9670,N_9872);
nor U10056 (N_10056,N_9610,N_9595);
xor U10057 (N_10057,N_9782,N_9884);
xor U10058 (N_10058,N_9664,N_9885);
nor U10059 (N_10059,N_9585,N_9602);
and U10060 (N_10060,N_9965,N_9826);
and U10061 (N_10061,N_9802,N_9500);
and U10062 (N_10062,N_9580,N_9950);
nand U10063 (N_10063,N_9620,N_9946);
and U10064 (N_10064,N_9686,N_9940);
nand U10065 (N_10065,N_9913,N_9757);
and U10066 (N_10066,N_9902,N_9552);
or U10067 (N_10067,N_9501,N_9582);
nor U10068 (N_10068,N_9998,N_9637);
or U10069 (N_10069,N_9990,N_9702);
xnor U10070 (N_10070,N_9528,N_9967);
nand U10071 (N_10071,N_9676,N_9714);
xnor U10072 (N_10072,N_9531,N_9973);
and U10073 (N_10073,N_9957,N_9644);
xor U10074 (N_10074,N_9718,N_9629);
nand U10075 (N_10075,N_9641,N_9985);
and U10076 (N_10076,N_9939,N_9999);
nand U10077 (N_10077,N_9652,N_9539);
nand U10078 (N_10078,N_9758,N_9992);
nand U10079 (N_10079,N_9529,N_9815);
nor U10080 (N_10080,N_9863,N_9548);
nor U10081 (N_10081,N_9935,N_9688);
nor U10082 (N_10082,N_9768,N_9687);
xor U10083 (N_10083,N_9597,N_9746);
nand U10084 (N_10084,N_9699,N_9504);
xor U10085 (N_10085,N_9659,N_9873);
nor U10086 (N_10086,N_9772,N_9959);
and U10087 (N_10087,N_9572,N_9559);
nand U10088 (N_10088,N_9978,N_9780);
xnor U10089 (N_10089,N_9777,N_9933);
or U10090 (N_10090,N_9989,N_9737);
nand U10091 (N_10091,N_9833,N_9795);
xor U10092 (N_10092,N_9669,N_9653);
nand U10093 (N_10093,N_9765,N_9961);
and U10094 (N_10094,N_9954,N_9853);
nor U10095 (N_10095,N_9824,N_9579);
nor U10096 (N_10096,N_9546,N_9667);
xnor U10097 (N_10097,N_9647,N_9626);
nor U10098 (N_10098,N_9861,N_9541);
nand U10099 (N_10099,N_9934,N_9514);
xor U10100 (N_10100,N_9930,N_9745);
or U10101 (N_10101,N_9801,N_9526);
xnor U10102 (N_10102,N_9571,N_9866);
or U10103 (N_10103,N_9717,N_9905);
nor U10104 (N_10104,N_9600,N_9942);
nand U10105 (N_10105,N_9503,N_9527);
nor U10106 (N_10106,N_9767,N_9834);
nor U10107 (N_10107,N_9614,N_9750);
nand U10108 (N_10108,N_9730,N_9938);
nor U10109 (N_10109,N_9809,N_9979);
nand U10110 (N_10110,N_9677,N_9793);
or U10111 (N_10111,N_9517,N_9556);
xor U10112 (N_10112,N_9825,N_9860);
xnor U10113 (N_10113,N_9506,N_9893);
and U10114 (N_10114,N_9922,N_9900);
nor U10115 (N_10115,N_9520,N_9598);
xnor U10116 (N_10116,N_9710,N_9947);
xor U10117 (N_10117,N_9544,N_9693);
nor U10118 (N_10118,N_9703,N_9855);
or U10119 (N_10119,N_9588,N_9889);
xnor U10120 (N_10120,N_9732,N_9762);
and U10121 (N_10121,N_9949,N_9991);
or U10122 (N_10122,N_9639,N_9918);
nand U10123 (N_10123,N_9770,N_9887);
nand U10124 (N_10124,N_9874,N_9774);
xor U10125 (N_10125,N_9744,N_9592);
or U10126 (N_10126,N_9736,N_9624);
and U10127 (N_10127,N_9618,N_9856);
nand U10128 (N_10128,N_9713,N_9773);
and U10129 (N_10129,N_9914,N_9911);
or U10130 (N_10130,N_9692,N_9830);
nand U10131 (N_10131,N_9636,N_9891);
nand U10132 (N_10132,N_9735,N_9823);
or U10133 (N_10133,N_9799,N_9870);
xor U10134 (N_10134,N_9612,N_9625);
nor U10135 (N_10135,N_9502,N_9551);
nor U10136 (N_10136,N_9658,N_9568);
and U10137 (N_10137,N_9565,N_9734);
and U10138 (N_10138,N_9895,N_9566);
nand U10139 (N_10139,N_9581,N_9738);
nor U10140 (N_10140,N_9540,N_9617);
xor U10141 (N_10141,N_9761,N_9822);
nand U10142 (N_10142,N_9883,N_9705);
xnor U10143 (N_10143,N_9993,N_9969);
nor U10144 (N_10144,N_9642,N_9848);
or U10145 (N_10145,N_9584,N_9543);
and U10146 (N_10146,N_9844,N_9682);
xnor U10147 (N_10147,N_9798,N_9662);
xor U10148 (N_10148,N_9739,N_9951);
xor U10149 (N_10149,N_9994,N_9771);
or U10150 (N_10150,N_9743,N_9747);
and U10151 (N_10151,N_9906,N_9678);
nand U10152 (N_10152,N_9787,N_9763);
xor U10153 (N_10153,N_9726,N_9845);
nor U10154 (N_10154,N_9674,N_9661);
nor U10155 (N_10155,N_9878,N_9689);
nand U10156 (N_10156,N_9711,N_9638);
or U10157 (N_10157,N_9525,N_9518);
nand U10158 (N_10158,N_9591,N_9596);
or U10159 (N_10159,N_9784,N_9953);
or U10160 (N_10160,N_9535,N_9841);
or U10161 (N_10161,N_9523,N_9680);
xor U10162 (N_10162,N_9827,N_9656);
nor U10163 (N_10163,N_9616,N_9849);
and U10164 (N_10164,N_9564,N_9936);
or U10165 (N_10165,N_9997,N_9577);
nor U10166 (N_10166,N_9972,N_9690);
nor U10167 (N_10167,N_9665,N_9764);
or U10168 (N_10168,N_9876,N_9651);
xnor U10169 (N_10169,N_9875,N_9672);
and U10170 (N_10170,N_9613,N_9807);
and U10171 (N_10171,N_9976,N_9813);
xor U10172 (N_10172,N_9557,N_9916);
nand U10173 (N_10173,N_9646,N_9945);
xor U10174 (N_10174,N_9590,N_9984);
and U10175 (N_10175,N_9562,N_9766);
xor U10176 (N_10176,N_9864,N_9971);
nor U10177 (N_10177,N_9881,N_9632);
nand U10178 (N_10178,N_9842,N_9781);
and U10179 (N_10179,N_9921,N_9865);
and U10180 (N_10180,N_9783,N_9666);
and U10181 (N_10181,N_9555,N_9920);
nor U10182 (N_10182,N_9536,N_9818);
and U10183 (N_10183,N_9929,N_9558);
nor U10184 (N_10184,N_9966,N_9589);
nor U10185 (N_10185,N_9675,N_9846);
nor U10186 (N_10186,N_9533,N_9909);
and U10187 (N_10187,N_9899,N_9567);
xnor U10188 (N_10188,N_9727,N_9695);
xnor U10189 (N_10189,N_9850,N_9721);
nand U10190 (N_10190,N_9759,N_9829);
and U10191 (N_10191,N_9901,N_9903);
and U10192 (N_10192,N_9576,N_9648);
nand U10193 (N_10193,N_9919,N_9635);
and U10194 (N_10194,N_9697,N_9742);
xor U10195 (N_10195,N_9839,N_9775);
and U10196 (N_10196,N_9655,N_9621);
or U10197 (N_10197,N_9560,N_9628);
xnor U10198 (N_10198,N_9507,N_9808);
and U10199 (N_10199,N_9740,N_9510);
or U10200 (N_10200,N_9696,N_9977);
nand U10201 (N_10201,N_9753,N_9890);
xnor U10202 (N_10202,N_9812,N_9941);
or U10203 (N_10203,N_9836,N_9796);
xnor U10204 (N_10204,N_9701,N_9749);
or U10205 (N_10205,N_9983,N_9894);
nor U10206 (N_10206,N_9988,N_9981);
nor U10207 (N_10207,N_9549,N_9843);
nand U10208 (N_10208,N_9851,N_9927);
nand U10209 (N_10209,N_9505,N_9751);
xnor U10210 (N_10210,N_9943,N_9896);
or U10211 (N_10211,N_9857,N_9538);
xor U10212 (N_10212,N_9958,N_9601);
nand U10213 (N_10213,N_9955,N_9698);
nor U10214 (N_10214,N_9828,N_9593);
nor U10215 (N_10215,N_9685,N_9908);
or U10216 (N_10216,N_9623,N_9915);
nor U10217 (N_10217,N_9630,N_9888);
nor U10218 (N_10218,N_9904,N_9715);
nor U10219 (N_10219,N_9694,N_9684);
or U10220 (N_10220,N_9615,N_9569);
or U10221 (N_10221,N_9789,N_9970);
or U10222 (N_10222,N_9869,N_9880);
or U10223 (N_10223,N_9583,N_9835);
and U10224 (N_10224,N_9640,N_9725);
nor U10225 (N_10225,N_9952,N_9923);
and U10226 (N_10226,N_9974,N_9877);
xor U10227 (N_10227,N_9910,N_9521);
and U10228 (N_10228,N_9563,N_9733);
or U10229 (N_10229,N_9960,N_9633);
nor U10230 (N_10230,N_9871,N_9660);
xnor U10231 (N_10231,N_9882,N_9650);
nand U10232 (N_10232,N_9859,N_9932);
xor U10233 (N_10233,N_9858,N_9924);
or U10234 (N_10234,N_9816,N_9663);
and U10235 (N_10235,N_9708,N_9785);
and U10236 (N_10236,N_9720,N_9681);
nand U10237 (N_10237,N_9963,N_9867);
xor U10238 (N_10238,N_9804,N_9723);
nor U10239 (N_10239,N_9995,N_9931);
and U10240 (N_10240,N_9622,N_9553);
xnor U10241 (N_10241,N_9847,N_9668);
or U10242 (N_10242,N_9852,N_9719);
xor U10243 (N_10243,N_9968,N_9779);
xnor U10244 (N_10244,N_9570,N_9609);
and U10245 (N_10245,N_9513,N_9657);
and U10246 (N_10246,N_9700,N_9519);
and U10247 (N_10247,N_9575,N_9522);
or U10248 (N_10248,N_9831,N_9631);
or U10249 (N_10249,N_9794,N_9542);
xor U10250 (N_10250,N_9781,N_9603);
and U10251 (N_10251,N_9556,N_9831);
nor U10252 (N_10252,N_9711,N_9517);
xnor U10253 (N_10253,N_9606,N_9536);
xnor U10254 (N_10254,N_9982,N_9839);
and U10255 (N_10255,N_9764,N_9917);
or U10256 (N_10256,N_9868,N_9828);
nand U10257 (N_10257,N_9795,N_9937);
nand U10258 (N_10258,N_9710,N_9790);
xor U10259 (N_10259,N_9864,N_9819);
xnor U10260 (N_10260,N_9916,N_9882);
nor U10261 (N_10261,N_9512,N_9632);
nand U10262 (N_10262,N_9574,N_9693);
xor U10263 (N_10263,N_9615,N_9576);
and U10264 (N_10264,N_9968,N_9639);
nor U10265 (N_10265,N_9874,N_9806);
and U10266 (N_10266,N_9943,N_9973);
or U10267 (N_10267,N_9509,N_9929);
and U10268 (N_10268,N_9878,N_9763);
xor U10269 (N_10269,N_9704,N_9757);
and U10270 (N_10270,N_9927,N_9819);
nor U10271 (N_10271,N_9832,N_9525);
nor U10272 (N_10272,N_9827,N_9526);
nand U10273 (N_10273,N_9917,N_9977);
and U10274 (N_10274,N_9791,N_9614);
nand U10275 (N_10275,N_9642,N_9731);
nor U10276 (N_10276,N_9525,N_9953);
and U10277 (N_10277,N_9878,N_9628);
xnor U10278 (N_10278,N_9606,N_9848);
xor U10279 (N_10279,N_9865,N_9944);
or U10280 (N_10280,N_9940,N_9609);
nor U10281 (N_10281,N_9525,N_9956);
and U10282 (N_10282,N_9617,N_9958);
nor U10283 (N_10283,N_9945,N_9788);
nand U10284 (N_10284,N_9753,N_9750);
nor U10285 (N_10285,N_9686,N_9564);
xnor U10286 (N_10286,N_9519,N_9723);
nor U10287 (N_10287,N_9703,N_9690);
nand U10288 (N_10288,N_9692,N_9968);
and U10289 (N_10289,N_9599,N_9909);
or U10290 (N_10290,N_9643,N_9812);
or U10291 (N_10291,N_9524,N_9676);
nor U10292 (N_10292,N_9526,N_9999);
nand U10293 (N_10293,N_9710,N_9997);
nor U10294 (N_10294,N_9735,N_9797);
or U10295 (N_10295,N_9711,N_9583);
or U10296 (N_10296,N_9575,N_9887);
nor U10297 (N_10297,N_9990,N_9964);
or U10298 (N_10298,N_9726,N_9893);
xor U10299 (N_10299,N_9781,N_9852);
xor U10300 (N_10300,N_9600,N_9597);
xor U10301 (N_10301,N_9729,N_9881);
nor U10302 (N_10302,N_9752,N_9868);
and U10303 (N_10303,N_9753,N_9717);
nor U10304 (N_10304,N_9756,N_9832);
xor U10305 (N_10305,N_9677,N_9589);
and U10306 (N_10306,N_9907,N_9865);
nor U10307 (N_10307,N_9823,N_9798);
or U10308 (N_10308,N_9560,N_9776);
and U10309 (N_10309,N_9510,N_9791);
or U10310 (N_10310,N_9546,N_9991);
or U10311 (N_10311,N_9860,N_9555);
nor U10312 (N_10312,N_9550,N_9583);
xnor U10313 (N_10313,N_9759,N_9682);
nor U10314 (N_10314,N_9978,N_9890);
xor U10315 (N_10315,N_9678,N_9614);
nand U10316 (N_10316,N_9761,N_9898);
or U10317 (N_10317,N_9702,N_9951);
and U10318 (N_10318,N_9951,N_9811);
xnor U10319 (N_10319,N_9505,N_9942);
nor U10320 (N_10320,N_9536,N_9593);
xor U10321 (N_10321,N_9798,N_9971);
nand U10322 (N_10322,N_9555,N_9547);
and U10323 (N_10323,N_9528,N_9773);
nand U10324 (N_10324,N_9996,N_9617);
xor U10325 (N_10325,N_9576,N_9598);
and U10326 (N_10326,N_9660,N_9797);
and U10327 (N_10327,N_9909,N_9928);
nand U10328 (N_10328,N_9939,N_9839);
nor U10329 (N_10329,N_9941,N_9626);
xor U10330 (N_10330,N_9564,N_9940);
xnor U10331 (N_10331,N_9594,N_9969);
or U10332 (N_10332,N_9882,N_9544);
xnor U10333 (N_10333,N_9801,N_9610);
and U10334 (N_10334,N_9556,N_9667);
nor U10335 (N_10335,N_9774,N_9596);
and U10336 (N_10336,N_9948,N_9593);
nor U10337 (N_10337,N_9892,N_9644);
xnor U10338 (N_10338,N_9897,N_9598);
xor U10339 (N_10339,N_9613,N_9745);
nor U10340 (N_10340,N_9542,N_9999);
and U10341 (N_10341,N_9583,N_9563);
nand U10342 (N_10342,N_9774,N_9510);
nor U10343 (N_10343,N_9995,N_9912);
or U10344 (N_10344,N_9517,N_9981);
nor U10345 (N_10345,N_9608,N_9705);
nand U10346 (N_10346,N_9733,N_9699);
or U10347 (N_10347,N_9527,N_9823);
or U10348 (N_10348,N_9633,N_9743);
and U10349 (N_10349,N_9707,N_9600);
nor U10350 (N_10350,N_9675,N_9554);
or U10351 (N_10351,N_9965,N_9666);
nand U10352 (N_10352,N_9549,N_9819);
nor U10353 (N_10353,N_9565,N_9512);
nor U10354 (N_10354,N_9595,N_9728);
and U10355 (N_10355,N_9758,N_9872);
xnor U10356 (N_10356,N_9873,N_9590);
nand U10357 (N_10357,N_9885,N_9590);
xor U10358 (N_10358,N_9559,N_9997);
nand U10359 (N_10359,N_9525,N_9859);
xnor U10360 (N_10360,N_9612,N_9518);
nor U10361 (N_10361,N_9791,N_9733);
or U10362 (N_10362,N_9540,N_9511);
nor U10363 (N_10363,N_9983,N_9887);
and U10364 (N_10364,N_9887,N_9870);
or U10365 (N_10365,N_9725,N_9780);
and U10366 (N_10366,N_9633,N_9689);
or U10367 (N_10367,N_9712,N_9538);
xnor U10368 (N_10368,N_9819,N_9611);
or U10369 (N_10369,N_9991,N_9957);
nand U10370 (N_10370,N_9703,N_9700);
nand U10371 (N_10371,N_9682,N_9791);
or U10372 (N_10372,N_9993,N_9806);
xor U10373 (N_10373,N_9684,N_9701);
nand U10374 (N_10374,N_9733,N_9529);
and U10375 (N_10375,N_9579,N_9747);
or U10376 (N_10376,N_9656,N_9900);
nor U10377 (N_10377,N_9844,N_9782);
nor U10378 (N_10378,N_9600,N_9764);
nand U10379 (N_10379,N_9597,N_9520);
and U10380 (N_10380,N_9785,N_9804);
nand U10381 (N_10381,N_9510,N_9715);
xnor U10382 (N_10382,N_9618,N_9500);
and U10383 (N_10383,N_9884,N_9755);
nor U10384 (N_10384,N_9983,N_9801);
nor U10385 (N_10385,N_9734,N_9808);
nand U10386 (N_10386,N_9899,N_9657);
nor U10387 (N_10387,N_9888,N_9952);
nand U10388 (N_10388,N_9605,N_9614);
nor U10389 (N_10389,N_9740,N_9935);
nand U10390 (N_10390,N_9916,N_9832);
and U10391 (N_10391,N_9888,N_9623);
nand U10392 (N_10392,N_9634,N_9986);
or U10393 (N_10393,N_9839,N_9750);
and U10394 (N_10394,N_9965,N_9698);
xnor U10395 (N_10395,N_9665,N_9765);
nor U10396 (N_10396,N_9558,N_9721);
or U10397 (N_10397,N_9679,N_9695);
and U10398 (N_10398,N_9996,N_9783);
or U10399 (N_10399,N_9544,N_9588);
and U10400 (N_10400,N_9555,N_9525);
nor U10401 (N_10401,N_9591,N_9678);
xor U10402 (N_10402,N_9781,N_9847);
nand U10403 (N_10403,N_9517,N_9695);
xor U10404 (N_10404,N_9538,N_9813);
xnor U10405 (N_10405,N_9906,N_9809);
xor U10406 (N_10406,N_9979,N_9970);
nor U10407 (N_10407,N_9805,N_9919);
or U10408 (N_10408,N_9589,N_9932);
nor U10409 (N_10409,N_9725,N_9684);
or U10410 (N_10410,N_9812,N_9907);
nor U10411 (N_10411,N_9832,N_9705);
and U10412 (N_10412,N_9523,N_9619);
nand U10413 (N_10413,N_9768,N_9900);
nor U10414 (N_10414,N_9610,N_9677);
xnor U10415 (N_10415,N_9999,N_9954);
xnor U10416 (N_10416,N_9738,N_9909);
xnor U10417 (N_10417,N_9886,N_9590);
or U10418 (N_10418,N_9650,N_9833);
nor U10419 (N_10419,N_9601,N_9885);
nand U10420 (N_10420,N_9609,N_9636);
nand U10421 (N_10421,N_9628,N_9793);
xnor U10422 (N_10422,N_9571,N_9920);
nand U10423 (N_10423,N_9812,N_9539);
and U10424 (N_10424,N_9920,N_9533);
nor U10425 (N_10425,N_9976,N_9827);
xor U10426 (N_10426,N_9835,N_9511);
or U10427 (N_10427,N_9900,N_9598);
nor U10428 (N_10428,N_9562,N_9921);
nor U10429 (N_10429,N_9704,N_9618);
nand U10430 (N_10430,N_9573,N_9745);
or U10431 (N_10431,N_9685,N_9703);
or U10432 (N_10432,N_9507,N_9676);
xnor U10433 (N_10433,N_9779,N_9839);
nor U10434 (N_10434,N_9680,N_9781);
and U10435 (N_10435,N_9935,N_9973);
nor U10436 (N_10436,N_9649,N_9818);
and U10437 (N_10437,N_9602,N_9518);
nor U10438 (N_10438,N_9657,N_9690);
nand U10439 (N_10439,N_9903,N_9870);
xor U10440 (N_10440,N_9504,N_9863);
nor U10441 (N_10441,N_9530,N_9633);
xor U10442 (N_10442,N_9717,N_9593);
nor U10443 (N_10443,N_9994,N_9689);
nor U10444 (N_10444,N_9806,N_9712);
or U10445 (N_10445,N_9621,N_9657);
or U10446 (N_10446,N_9864,N_9698);
nand U10447 (N_10447,N_9593,N_9924);
nand U10448 (N_10448,N_9845,N_9989);
xor U10449 (N_10449,N_9545,N_9546);
nor U10450 (N_10450,N_9938,N_9697);
nand U10451 (N_10451,N_9703,N_9763);
or U10452 (N_10452,N_9949,N_9803);
and U10453 (N_10453,N_9621,N_9679);
xnor U10454 (N_10454,N_9575,N_9504);
and U10455 (N_10455,N_9992,N_9867);
nor U10456 (N_10456,N_9758,N_9951);
nor U10457 (N_10457,N_9552,N_9811);
or U10458 (N_10458,N_9595,N_9505);
or U10459 (N_10459,N_9805,N_9524);
xor U10460 (N_10460,N_9928,N_9560);
or U10461 (N_10461,N_9601,N_9884);
and U10462 (N_10462,N_9599,N_9590);
xnor U10463 (N_10463,N_9542,N_9863);
or U10464 (N_10464,N_9860,N_9838);
nor U10465 (N_10465,N_9516,N_9557);
or U10466 (N_10466,N_9683,N_9784);
and U10467 (N_10467,N_9538,N_9549);
or U10468 (N_10468,N_9543,N_9962);
nand U10469 (N_10469,N_9700,N_9782);
xor U10470 (N_10470,N_9993,N_9741);
nand U10471 (N_10471,N_9945,N_9548);
and U10472 (N_10472,N_9624,N_9674);
nor U10473 (N_10473,N_9841,N_9907);
xor U10474 (N_10474,N_9768,N_9600);
nand U10475 (N_10475,N_9908,N_9967);
nor U10476 (N_10476,N_9614,N_9720);
nand U10477 (N_10477,N_9914,N_9981);
or U10478 (N_10478,N_9787,N_9842);
or U10479 (N_10479,N_9584,N_9964);
nor U10480 (N_10480,N_9592,N_9756);
nor U10481 (N_10481,N_9578,N_9978);
or U10482 (N_10482,N_9797,N_9914);
or U10483 (N_10483,N_9736,N_9916);
or U10484 (N_10484,N_9681,N_9948);
nor U10485 (N_10485,N_9873,N_9530);
nor U10486 (N_10486,N_9607,N_9541);
and U10487 (N_10487,N_9619,N_9613);
or U10488 (N_10488,N_9744,N_9791);
or U10489 (N_10489,N_9591,N_9725);
or U10490 (N_10490,N_9814,N_9906);
and U10491 (N_10491,N_9529,N_9650);
nand U10492 (N_10492,N_9904,N_9584);
and U10493 (N_10493,N_9855,N_9698);
nor U10494 (N_10494,N_9793,N_9992);
or U10495 (N_10495,N_9698,N_9852);
xnor U10496 (N_10496,N_9708,N_9637);
xor U10497 (N_10497,N_9941,N_9652);
xnor U10498 (N_10498,N_9987,N_9700);
nand U10499 (N_10499,N_9500,N_9889);
and U10500 (N_10500,N_10168,N_10129);
and U10501 (N_10501,N_10302,N_10043);
or U10502 (N_10502,N_10052,N_10249);
or U10503 (N_10503,N_10425,N_10083);
nand U10504 (N_10504,N_10225,N_10200);
nor U10505 (N_10505,N_10109,N_10223);
xor U10506 (N_10506,N_10299,N_10211);
and U10507 (N_10507,N_10478,N_10330);
or U10508 (N_10508,N_10235,N_10192);
nor U10509 (N_10509,N_10422,N_10405);
nand U10510 (N_10510,N_10306,N_10244);
and U10511 (N_10511,N_10059,N_10335);
nand U10512 (N_10512,N_10466,N_10247);
nor U10513 (N_10513,N_10004,N_10447);
xor U10514 (N_10514,N_10276,N_10137);
nor U10515 (N_10515,N_10414,N_10063);
or U10516 (N_10516,N_10366,N_10490);
nand U10517 (N_10517,N_10240,N_10013);
xor U10518 (N_10518,N_10452,N_10336);
nor U10519 (N_10519,N_10097,N_10324);
xor U10520 (N_10520,N_10162,N_10005);
xnor U10521 (N_10521,N_10309,N_10001);
xor U10522 (N_10522,N_10499,N_10426);
nor U10523 (N_10523,N_10294,N_10160);
or U10524 (N_10524,N_10174,N_10198);
nor U10525 (N_10525,N_10251,N_10081);
xor U10526 (N_10526,N_10238,N_10451);
xor U10527 (N_10527,N_10475,N_10012);
nand U10528 (N_10528,N_10108,N_10494);
and U10529 (N_10529,N_10334,N_10115);
and U10530 (N_10530,N_10224,N_10180);
or U10531 (N_10531,N_10443,N_10088);
nor U10532 (N_10532,N_10188,N_10181);
and U10533 (N_10533,N_10482,N_10374);
nand U10534 (N_10534,N_10460,N_10380);
xor U10535 (N_10535,N_10323,N_10497);
nand U10536 (N_10536,N_10203,N_10357);
nand U10537 (N_10537,N_10364,N_10445);
nand U10538 (N_10538,N_10021,N_10313);
and U10539 (N_10539,N_10411,N_10142);
or U10540 (N_10540,N_10301,N_10123);
nand U10541 (N_10541,N_10328,N_10412);
or U10542 (N_10542,N_10387,N_10427);
or U10543 (N_10543,N_10440,N_10404);
nand U10544 (N_10544,N_10045,N_10477);
and U10545 (N_10545,N_10421,N_10454);
and U10546 (N_10546,N_10161,N_10036);
and U10547 (N_10547,N_10069,N_10316);
xor U10548 (N_10548,N_10250,N_10362);
nor U10549 (N_10549,N_10114,N_10220);
and U10550 (N_10550,N_10228,N_10212);
or U10551 (N_10551,N_10197,N_10070);
or U10552 (N_10552,N_10331,N_10367);
nor U10553 (N_10553,N_10393,N_10020);
nor U10554 (N_10554,N_10435,N_10010);
nor U10555 (N_10555,N_10053,N_10355);
xor U10556 (N_10556,N_10468,N_10448);
or U10557 (N_10557,N_10205,N_10319);
nor U10558 (N_10558,N_10274,N_10107);
xnor U10559 (N_10559,N_10014,N_10345);
xnor U10560 (N_10560,N_10077,N_10480);
and U10561 (N_10561,N_10498,N_10476);
xor U10562 (N_10562,N_10314,N_10450);
and U10563 (N_10563,N_10265,N_10024);
xnor U10564 (N_10564,N_10060,N_10399);
xnor U10565 (N_10565,N_10463,N_10356);
and U10566 (N_10566,N_10491,N_10159);
or U10567 (N_10567,N_10325,N_10076);
and U10568 (N_10568,N_10288,N_10397);
xnor U10569 (N_10569,N_10110,N_10248);
or U10570 (N_10570,N_10230,N_10271);
or U10571 (N_10571,N_10297,N_10116);
nor U10572 (N_10572,N_10103,N_10437);
or U10573 (N_10573,N_10144,N_10227);
nand U10574 (N_10574,N_10474,N_10183);
xnor U10575 (N_10575,N_10255,N_10464);
nor U10576 (N_10576,N_10369,N_10434);
and U10577 (N_10577,N_10204,N_10022);
nand U10578 (N_10578,N_10193,N_10121);
or U10579 (N_10579,N_10016,N_10033);
or U10580 (N_10580,N_10315,N_10312);
or U10581 (N_10581,N_10011,N_10243);
or U10582 (N_10582,N_10195,N_10229);
nor U10583 (N_10583,N_10032,N_10171);
nor U10584 (N_10584,N_10237,N_10322);
nand U10585 (N_10585,N_10000,N_10136);
nand U10586 (N_10586,N_10067,N_10416);
nor U10587 (N_10587,N_10376,N_10140);
xor U10588 (N_10588,N_10038,N_10037);
xor U10589 (N_10589,N_10156,N_10317);
nor U10590 (N_10590,N_10239,N_10175);
xnor U10591 (N_10591,N_10068,N_10101);
and U10592 (N_10592,N_10337,N_10484);
and U10593 (N_10593,N_10326,N_10293);
or U10594 (N_10594,N_10148,N_10072);
and U10595 (N_10595,N_10394,N_10285);
nor U10596 (N_10596,N_10481,N_10157);
nor U10597 (N_10597,N_10260,N_10100);
nand U10598 (N_10598,N_10075,N_10145);
xor U10599 (N_10599,N_10409,N_10209);
nor U10600 (N_10600,N_10358,N_10341);
xor U10601 (N_10601,N_10257,N_10094);
xnor U10602 (N_10602,N_10388,N_10300);
and U10603 (N_10603,N_10365,N_10190);
and U10604 (N_10604,N_10473,N_10007);
xnor U10605 (N_10605,N_10368,N_10402);
nor U10606 (N_10606,N_10206,N_10079);
nand U10607 (N_10607,N_10122,N_10396);
or U10608 (N_10608,N_10270,N_10289);
xnor U10609 (N_10609,N_10361,N_10392);
or U10610 (N_10610,N_10253,N_10058);
nand U10611 (N_10611,N_10329,N_10146);
xor U10612 (N_10612,N_10143,N_10150);
nand U10613 (N_10613,N_10234,N_10026);
or U10614 (N_10614,N_10102,N_10470);
xnor U10615 (N_10615,N_10196,N_10410);
or U10616 (N_10616,N_10166,N_10332);
or U10617 (N_10617,N_10446,N_10495);
nor U10618 (N_10618,N_10210,N_10202);
xor U10619 (N_10619,N_10099,N_10398);
and U10620 (N_10620,N_10370,N_10381);
nor U10621 (N_10621,N_10208,N_10029);
or U10622 (N_10622,N_10308,N_10233);
xor U10623 (N_10623,N_10035,N_10106);
xor U10624 (N_10624,N_10269,N_10456);
nand U10625 (N_10625,N_10406,N_10177);
or U10626 (N_10626,N_10401,N_10111);
nand U10627 (N_10627,N_10483,N_10442);
and U10628 (N_10628,N_10092,N_10453);
xnor U10629 (N_10629,N_10219,N_10382);
xor U10630 (N_10630,N_10119,N_10226);
nor U10631 (N_10631,N_10305,N_10379);
or U10632 (N_10632,N_10173,N_10048);
nor U10633 (N_10633,N_10283,N_10112);
nand U10634 (N_10634,N_10436,N_10429);
xor U10635 (N_10635,N_10178,N_10047);
or U10636 (N_10636,N_10373,N_10261);
or U10637 (N_10637,N_10222,N_10496);
xnor U10638 (N_10638,N_10359,N_10096);
and U10639 (N_10639,N_10182,N_10286);
nand U10640 (N_10640,N_10127,N_10098);
nor U10641 (N_10641,N_10184,N_10236);
nor U10642 (N_10642,N_10384,N_10179);
or U10643 (N_10643,N_10280,N_10041);
or U10644 (N_10644,N_10186,N_10057);
nand U10645 (N_10645,N_10084,N_10438);
nand U10646 (N_10646,N_10458,N_10066);
xor U10647 (N_10647,N_10028,N_10272);
xnor U10648 (N_10648,N_10459,N_10113);
and U10649 (N_10649,N_10167,N_10154);
xnor U10650 (N_10650,N_10488,N_10485);
or U10651 (N_10651,N_10486,N_10055);
and U10652 (N_10652,N_10279,N_10338);
or U10653 (N_10653,N_10034,N_10245);
or U10654 (N_10654,N_10120,N_10147);
and U10655 (N_10655,N_10135,N_10126);
nand U10656 (N_10656,N_10472,N_10489);
xnor U10657 (N_10657,N_10242,N_10377);
and U10658 (N_10658,N_10089,N_10264);
xnor U10659 (N_10659,N_10049,N_10125);
and U10660 (N_10660,N_10131,N_10018);
nand U10661 (N_10661,N_10277,N_10407);
nand U10662 (N_10662,N_10169,N_10064);
nor U10663 (N_10663,N_10130,N_10340);
xnor U10664 (N_10664,N_10295,N_10002);
or U10665 (N_10665,N_10133,N_10441);
nand U10666 (N_10666,N_10093,N_10284);
or U10667 (N_10667,N_10104,N_10263);
nand U10668 (N_10668,N_10006,N_10395);
or U10669 (N_10669,N_10419,N_10351);
nor U10670 (N_10670,N_10085,N_10039);
or U10671 (N_10671,N_10139,N_10372);
and U10672 (N_10672,N_10273,N_10266);
nor U10673 (N_10673,N_10415,N_10389);
nor U10674 (N_10674,N_10417,N_10124);
nand U10675 (N_10675,N_10073,N_10040);
or U10676 (N_10676,N_10354,N_10433);
and U10677 (N_10677,N_10090,N_10091);
or U10678 (N_10678,N_10278,N_10153);
or U10679 (N_10679,N_10462,N_10375);
nor U10680 (N_10680,N_10082,N_10493);
xor U10681 (N_10681,N_10296,N_10194);
nand U10682 (N_10682,N_10025,N_10413);
and U10683 (N_10683,N_10027,N_10042);
nand U10684 (N_10684,N_10391,N_10347);
or U10685 (N_10685,N_10141,N_10214);
or U10686 (N_10686,N_10267,N_10371);
xnor U10687 (N_10687,N_10163,N_10008);
nand U10688 (N_10688,N_10086,N_10439);
xnor U10689 (N_10689,N_10134,N_10282);
nand U10690 (N_10690,N_10221,N_10117);
nand U10691 (N_10691,N_10187,N_10149);
nand U10692 (N_10692,N_10201,N_10138);
nand U10693 (N_10693,N_10465,N_10231);
xor U10694 (N_10694,N_10418,N_10428);
nand U10695 (N_10695,N_10350,N_10449);
or U10696 (N_10696,N_10444,N_10339);
and U10697 (N_10697,N_10333,N_10383);
nand U10698 (N_10698,N_10307,N_10132);
nor U10699 (N_10699,N_10469,N_10065);
and U10700 (N_10700,N_10378,N_10360);
or U10701 (N_10701,N_10246,N_10050);
or U10702 (N_10702,N_10479,N_10430);
and U10703 (N_10703,N_10185,N_10199);
nor U10704 (N_10704,N_10487,N_10281);
nor U10705 (N_10705,N_10087,N_10424);
nor U10706 (N_10706,N_10385,N_10256);
nor U10707 (N_10707,N_10218,N_10054);
nand U10708 (N_10708,N_10348,N_10343);
nor U10709 (N_10709,N_10386,N_10216);
xnor U10710 (N_10710,N_10268,N_10292);
and U10711 (N_10711,N_10342,N_10170);
xnor U10712 (N_10712,N_10363,N_10078);
xor U10713 (N_10713,N_10304,N_10291);
and U10714 (N_10714,N_10031,N_10213);
or U10715 (N_10715,N_10321,N_10262);
xor U10716 (N_10716,N_10017,N_10423);
nor U10717 (N_10717,N_10003,N_10352);
nand U10718 (N_10718,N_10492,N_10056);
or U10719 (N_10719,N_10023,N_10164);
or U10720 (N_10720,N_10431,N_10151);
nor U10721 (N_10721,N_10259,N_10349);
nand U10722 (N_10722,N_10311,N_10457);
nand U10723 (N_10723,N_10118,N_10062);
or U10724 (N_10724,N_10071,N_10320);
and U10725 (N_10725,N_10080,N_10420);
or U10726 (N_10726,N_10400,N_10232);
nand U10727 (N_10727,N_10252,N_10061);
xnor U10728 (N_10728,N_10030,N_10408);
nand U10729 (N_10729,N_10105,N_10471);
nand U10730 (N_10730,N_10074,N_10152);
nor U10731 (N_10731,N_10015,N_10344);
nor U10732 (N_10732,N_10191,N_10128);
nand U10733 (N_10733,N_10290,N_10275);
xor U10734 (N_10734,N_10165,N_10044);
nand U10735 (N_10735,N_10217,N_10403);
xnor U10736 (N_10736,N_10346,N_10298);
or U10737 (N_10737,N_10158,N_10390);
xnor U10738 (N_10738,N_10353,N_10019);
and U10739 (N_10739,N_10318,N_10467);
xor U10740 (N_10740,N_10172,N_10455);
xor U10741 (N_10741,N_10287,N_10051);
xor U10742 (N_10742,N_10310,N_10461);
and U10743 (N_10743,N_10189,N_10432);
and U10744 (N_10744,N_10215,N_10176);
xnor U10745 (N_10745,N_10009,N_10207);
nand U10746 (N_10746,N_10303,N_10046);
xor U10747 (N_10747,N_10254,N_10241);
xnor U10748 (N_10748,N_10095,N_10258);
nor U10749 (N_10749,N_10155,N_10327);
and U10750 (N_10750,N_10387,N_10290);
and U10751 (N_10751,N_10094,N_10013);
nand U10752 (N_10752,N_10024,N_10417);
nand U10753 (N_10753,N_10098,N_10281);
and U10754 (N_10754,N_10376,N_10362);
nand U10755 (N_10755,N_10468,N_10445);
xnor U10756 (N_10756,N_10334,N_10072);
or U10757 (N_10757,N_10410,N_10381);
and U10758 (N_10758,N_10421,N_10085);
or U10759 (N_10759,N_10461,N_10114);
xnor U10760 (N_10760,N_10083,N_10029);
and U10761 (N_10761,N_10024,N_10190);
and U10762 (N_10762,N_10342,N_10334);
and U10763 (N_10763,N_10321,N_10213);
or U10764 (N_10764,N_10101,N_10014);
xnor U10765 (N_10765,N_10010,N_10341);
nor U10766 (N_10766,N_10383,N_10178);
and U10767 (N_10767,N_10387,N_10299);
nor U10768 (N_10768,N_10326,N_10003);
and U10769 (N_10769,N_10498,N_10251);
and U10770 (N_10770,N_10385,N_10012);
nor U10771 (N_10771,N_10051,N_10361);
nor U10772 (N_10772,N_10037,N_10229);
nand U10773 (N_10773,N_10089,N_10358);
and U10774 (N_10774,N_10429,N_10013);
or U10775 (N_10775,N_10313,N_10484);
nand U10776 (N_10776,N_10208,N_10391);
and U10777 (N_10777,N_10147,N_10169);
xor U10778 (N_10778,N_10001,N_10274);
and U10779 (N_10779,N_10132,N_10222);
nand U10780 (N_10780,N_10202,N_10186);
or U10781 (N_10781,N_10246,N_10074);
nor U10782 (N_10782,N_10032,N_10178);
and U10783 (N_10783,N_10068,N_10109);
xor U10784 (N_10784,N_10353,N_10344);
xnor U10785 (N_10785,N_10269,N_10384);
xor U10786 (N_10786,N_10320,N_10438);
nor U10787 (N_10787,N_10084,N_10102);
or U10788 (N_10788,N_10217,N_10058);
or U10789 (N_10789,N_10259,N_10147);
or U10790 (N_10790,N_10274,N_10199);
or U10791 (N_10791,N_10371,N_10320);
or U10792 (N_10792,N_10360,N_10406);
nand U10793 (N_10793,N_10229,N_10124);
nand U10794 (N_10794,N_10171,N_10275);
xnor U10795 (N_10795,N_10007,N_10193);
or U10796 (N_10796,N_10175,N_10479);
nor U10797 (N_10797,N_10138,N_10375);
nor U10798 (N_10798,N_10099,N_10291);
or U10799 (N_10799,N_10035,N_10382);
nand U10800 (N_10800,N_10110,N_10498);
and U10801 (N_10801,N_10230,N_10125);
and U10802 (N_10802,N_10326,N_10448);
and U10803 (N_10803,N_10283,N_10440);
or U10804 (N_10804,N_10223,N_10005);
nor U10805 (N_10805,N_10105,N_10458);
nor U10806 (N_10806,N_10333,N_10331);
or U10807 (N_10807,N_10006,N_10036);
nor U10808 (N_10808,N_10359,N_10308);
and U10809 (N_10809,N_10421,N_10437);
nand U10810 (N_10810,N_10241,N_10215);
and U10811 (N_10811,N_10173,N_10307);
nor U10812 (N_10812,N_10444,N_10187);
nand U10813 (N_10813,N_10236,N_10145);
or U10814 (N_10814,N_10178,N_10466);
nand U10815 (N_10815,N_10193,N_10370);
or U10816 (N_10816,N_10033,N_10090);
nor U10817 (N_10817,N_10313,N_10395);
xor U10818 (N_10818,N_10188,N_10027);
nand U10819 (N_10819,N_10336,N_10129);
nand U10820 (N_10820,N_10082,N_10322);
or U10821 (N_10821,N_10211,N_10156);
xnor U10822 (N_10822,N_10160,N_10277);
nor U10823 (N_10823,N_10226,N_10131);
nand U10824 (N_10824,N_10367,N_10275);
nor U10825 (N_10825,N_10200,N_10047);
xor U10826 (N_10826,N_10038,N_10497);
nor U10827 (N_10827,N_10270,N_10068);
or U10828 (N_10828,N_10129,N_10071);
xor U10829 (N_10829,N_10215,N_10072);
and U10830 (N_10830,N_10063,N_10154);
xnor U10831 (N_10831,N_10282,N_10034);
nand U10832 (N_10832,N_10456,N_10100);
and U10833 (N_10833,N_10372,N_10044);
or U10834 (N_10834,N_10499,N_10070);
or U10835 (N_10835,N_10063,N_10012);
xor U10836 (N_10836,N_10105,N_10020);
and U10837 (N_10837,N_10440,N_10443);
xor U10838 (N_10838,N_10058,N_10178);
nand U10839 (N_10839,N_10312,N_10351);
xnor U10840 (N_10840,N_10100,N_10058);
and U10841 (N_10841,N_10075,N_10353);
or U10842 (N_10842,N_10466,N_10016);
and U10843 (N_10843,N_10201,N_10466);
nand U10844 (N_10844,N_10323,N_10283);
and U10845 (N_10845,N_10326,N_10397);
nand U10846 (N_10846,N_10022,N_10410);
nor U10847 (N_10847,N_10333,N_10052);
and U10848 (N_10848,N_10081,N_10292);
nand U10849 (N_10849,N_10131,N_10039);
nand U10850 (N_10850,N_10453,N_10087);
xor U10851 (N_10851,N_10394,N_10275);
or U10852 (N_10852,N_10265,N_10166);
or U10853 (N_10853,N_10223,N_10370);
or U10854 (N_10854,N_10321,N_10275);
xnor U10855 (N_10855,N_10090,N_10066);
xor U10856 (N_10856,N_10223,N_10081);
nor U10857 (N_10857,N_10438,N_10015);
nand U10858 (N_10858,N_10012,N_10113);
or U10859 (N_10859,N_10382,N_10086);
or U10860 (N_10860,N_10349,N_10253);
nor U10861 (N_10861,N_10298,N_10326);
nand U10862 (N_10862,N_10498,N_10443);
nor U10863 (N_10863,N_10001,N_10042);
nand U10864 (N_10864,N_10425,N_10204);
xor U10865 (N_10865,N_10007,N_10488);
nand U10866 (N_10866,N_10057,N_10322);
and U10867 (N_10867,N_10366,N_10372);
xor U10868 (N_10868,N_10327,N_10159);
xor U10869 (N_10869,N_10321,N_10165);
nand U10870 (N_10870,N_10309,N_10043);
nand U10871 (N_10871,N_10475,N_10416);
xnor U10872 (N_10872,N_10427,N_10484);
nand U10873 (N_10873,N_10142,N_10391);
or U10874 (N_10874,N_10004,N_10337);
or U10875 (N_10875,N_10116,N_10348);
nand U10876 (N_10876,N_10330,N_10247);
nand U10877 (N_10877,N_10145,N_10437);
nand U10878 (N_10878,N_10381,N_10233);
xnor U10879 (N_10879,N_10133,N_10125);
and U10880 (N_10880,N_10242,N_10366);
or U10881 (N_10881,N_10414,N_10232);
nor U10882 (N_10882,N_10393,N_10346);
nor U10883 (N_10883,N_10131,N_10318);
xnor U10884 (N_10884,N_10272,N_10482);
or U10885 (N_10885,N_10132,N_10365);
or U10886 (N_10886,N_10484,N_10083);
nand U10887 (N_10887,N_10288,N_10011);
or U10888 (N_10888,N_10270,N_10442);
nor U10889 (N_10889,N_10004,N_10351);
or U10890 (N_10890,N_10076,N_10204);
nor U10891 (N_10891,N_10463,N_10344);
or U10892 (N_10892,N_10366,N_10315);
and U10893 (N_10893,N_10335,N_10396);
xnor U10894 (N_10894,N_10354,N_10153);
nand U10895 (N_10895,N_10309,N_10198);
xnor U10896 (N_10896,N_10218,N_10177);
or U10897 (N_10897,N_10376,N_10483);
or U10898 (N_10898,N_10276,N_10145);
or U10899 (N_10899,N_10382,N_10212);
xnor U10900 (N_10900,N_10024,N_10045);
or U10901 (N_10901,N_10109,N_10348);
xnor U10902 (N_10902,N_10178,N_10489);
or U10903 (N_10903,N_10323,N_10465);
nor U10904 (N_10904,N_10168,N_10255);
and U10905 (N_10905,N_10469,N_10378);
or U10906 (N_10906,N_10494,N_10358);
xor U10907 (N_10907,N_10211,N_10288);
or U10908 (N_10908,N_10418,N_10477);
or U10909 (N_10909,N_10009,N_10300);
nor U10910 (N_10910,N_10039,N_10345);
and U10911 (N_10911,N_10439,N_10128);
xnor U10912 (N_10912,N_10125,N_10386);
and U10913 (N_10913,N_10496,N_10444);
and U10914 (N_10914,N_10025,N_10448);
nor U10915 (N_10915,N_10488,N_10378);
and U10916 (N_10916,N_10465,N_10070);
nor U10917 (N_10917,N_10430,N_10116);
nor U10918 (N_10918,N_10383,N_10475);
and U10919 (N_10919,N_10116,N_10307);
nor U10920 (N_10920,N_10204,N_10095);
and U10921 (N_10921,N_10252,N_10297);
or U10922 (N_10922,N_10080,N_10269);
and U10923 (N_10923,N_10257,N_10284);
or U10924 (N_10924,N_10496,N_10477);
nor U10925 (N_10925,N_10258,N_10068);
xnor U10926 (N_10926,N_10344,N_10027);
nand U10927 (N_10927,N_10274,N_10095);
and U10928 (N_10928,N_10414,N_10195);
nand U10929 (N_10929,N_10307,N_10105);
xnor U10930 (N_10930,N_10117,N_10439);
xor U10931 (N_10931,N_10339,N_10056);
xnor U10932 (N_10932,N_10192,N_10226);
and U10933 (N_10933,N_10302,N_10291);
nand U10934 (N_10934,N_10280,N_10111);
and U10935 (N_10935,N_10461,N_10490);
and U10936 (N_10936,N_10004,N_10184);
and U10937 (N_10937,N_10442,N_10103);
nand U10938 (N_10938,N_10352,N_10362);
xor U10939 (N_10939,N_10074,N_10465);
and U10940 (N_10940,N_10071,N_10237);
and U10941 (N_10941,N_10342,N_10098);
nor U10942 (N_10942,N_10225,N_10006);
or U10943 (N_10943,N_10273,N_10404);
xor U10944 (N_10944,N_10453,N_10189);
nor U10945 (N_10945,N_10089,N_10473);
nor U10946 (N_10946,N_10082,N_10340);
nand U10947 (N_10947,N_10052,N_10150);
xor U10948 (N_10948,N_10338,N_10383);
or U10949 (N_10949,N_10077,N_10035);
nor U10950 (N_10950,N_10473,N_10023);
and U10951 (N_10951,N_10031,N_10352);
xor U10952 (N_10952,N_10290,N_10447);
and U10953 (N_10953,N_10178,N_10207);
xnor U10954 (N_10954,N_10271,N_10390);
nand U10955 (N_10955,N_10288,N_10476);
or U10956 (N_10956,N_10124,N_10214);
or U10957 (N_10957,N_10083,N_10444);
nor U10958 (N_10958,N_10417,N_10099);
and U10959 (N_10959,N_10082,N_10231);
nor U10960 (N_10960,N_10126,N_10013);
or U10961 (N_10961,N_10229,N_10009);
or U10962 (N_10962,N_10433,N_10298);
xnor U10963 (N_10963,N_10151,N_10395);
nor U10964 (N_10964,N_10466,N_10436);
nand U10965 (N_10965,N_10108,N_10085);
nand U10966 (N_10966,N_10050,N_10482);
and U10967 (N_10967,N_10292,N_10042);
nand U10968 (N_10968,N_10223,N_10419);
and U10969 (N_10969,N_10026,N_10045);
xnor U10970 (N_10970,N_10293,N_10345);
nand U10971 (N_10971,N_10197,N_10151);
nand U10972 (N_10972,N_10090,N_10369);
nor U10973 (N_10973,N_10118,N_10167);
xor U10974 (N_10974,N_10235,N_10227);
xnor U10975 (N_10975,N_10445,N_10262);
nor U10976 (N_10976,N_10081,N_10215);
nand U10977 (N_10977,N_10081,N_10179);
nor U10978 (N_10978,N_10492,N_10142);
and U10979 (N_10979,N_10007,N_10068);
and U10980 (N_10980,N_10146,N_10332);
or U10981 (N_10981,N_10006,N_10459);
nand U10982 (N_10982,N_10113,N_10054);
xnor U10983 (N_10983,N_10152,N_10398);
xor U10984 (N_10984,N_10038,N_10164);
nand U10985 (N_10985,N_10317,N_10180);
nand U10986 (N_10986,N_10365,N_10156);
and U10987 (N_10987,N_10104,N_10440);
nor U10988 (N_10988,N_10442,N_10230);
and U10989 (N_10989,N_10441,N_10153);
or U10990 (N_10990,N_10291,N_10058);
and U10991 (N_10991,N_10361,N_10158);
or U10992 (N_10992,N_10439,N_10431);
or U10993 (N_10993,N_10317,N_10391);
xor U10994 (N_10994,N_10469,N_10460);
nor U10995 (N_10995,N_10445,N_10314);
nand U10996 (N_10996,N_10460,N_10166);
and U10997 (N_10997,N_10297,N_10197);
xor U10998 (N_10998,N_10107,N_10233);
nand U10999 (N_10999,N_10249,N_10446);
xnor U11000 (N_11000,N_10733,N_10589);
or U11001 (N_11001,N_10585,N_10880);
or U11002 (N_11002,N_10685,N_10881);
xnor U11003 (N_11003,N_10853,N_10785);
nand U11004 (N_11004,N_10965,N_10800);
and U11005 (N_11005,N_10550,N_10931);
xnor U11006 (N_11006,N_10503,N_10628);
nand U11007 (N_11007,N_10994,N_10677);
xnor U11008 (N_11008,N_10643,N_10575);
and U11009 (N_11009,N_10809,N_10946);
xor U11010 (N_11010,N_10766,N_10837);
nor U11011 (N_11011,N_10966,N_10990);
nor U11012 (N_11012,N_10744,N_10811);
nand U11013 (N_11013,N_10856,N_10715);
nand U11014 (N_11014,N_10699,N_10875);
xor U11015 (N_11015,N_10641,N_10983);
or U11016 (N_11016,N_10666,N_10908);
xor U11017 (N_11017,N_10708,N_10526);
or U11018 (N_11018,N_10635,N_10629);
and U11019 (N_11019,N_10514,N_10997);
xor U11020 (N_11020,N_10816,N_10841);
nand U11021 (N_11021,N_10764,N_10555);
nor U11022 (N_11022,N_10612,N_10721);
xnor U11023 (N_11023,N_10644,N_10833);
or U11024 (N_11024,N_10515,N_10740);
nor U11025 (N_11025,N_10934,N_10576);
nand U11026 (N_11026,N_10835,N_10971);
and U11027 (N_11027,N_10895,N_10537);
nand U11028 (N_11028,N_10595,N_10977);
or U11029 (N_11029,N_10716,N_10903);
nand U11030 (N_11030,N_10993,N_10639);
or U11031 (N_11031,N_10516,N_10756);
nand U11032 (N_11032,N_10705,N_10664);
nor U11033 (N_11033,N_10673,N_10929);
xnor U11034 (N_11034,N_10519,N_10777);
nand U11035 (N_11035,N_10583,N_10761);
or U11036 (N_11036,N_10548,N_10792);
and U11037 (N_11037,N_10562,N_10989);
or U11038 (N_11038,N_10889,N_10870);
nand U11039 (N_11039,N_10791,N_10571);
xor U11040 (N_11040,N_10649,N_10810);
or U11041 (N_11041,N_10577,N_10963);
xnor U11042 (N_11042,N_10674,N_10836);
and U11043 (N_11043,N_10597,N_10845);
or U11044 (N_11044,N_10572,N_10596);
and U11045 (N_11045,N_10776,N_10787);
nor U11046 (N_11046,N_10942,N_10618);
xnor U11047 (N_11047,N_10857,N_10743);
or U11048 (N_11048,N_10926,N_10952);
nor U11049 (N_11049,N_10688,N_10902);
and U11050 (N_11050,N_10501,N_10788);
nand U11051 (N_11051,N_10861,N_10754);
nor U11052 (N_11052,N_10812,N_10707);
or U11053 (N_11053,N_10603,N_10506);
and U11054 (N_11054,N_10517,N_10502);
and U11055 (N_11055,N_10808,N_10636);
xor U11056 (N_11056,N_10827,N_10591);
nand U11057 (N_11057,N_10654,N_10860);
or U11058 (N_11058,N_10554,N_10710);
nand U11059 (N_11059,N_10752,N_10974);
and U11060 (N_11060,N_10739,N_10694);
xor U11061 (N_11061,N_10704,N_10614);
nand U11062 (N_11062,N_10524,N_10953);
or U11063 (N_11063,N_10558,N_10806);
xnor U11064 (N_11064,N_10862,N_10834);
xnor U11065 (N_11065,N_10540,N_10765);
xor U11066 (N_11066,N_10958,N_10538);
nor U11067 (N_11067,N_10962,N_10858);
or U11068 (N_11068,N_10701,N_10645);
nor U11069 (N_11069,N_10923,N_10536);
nor U11070 (N_11070,N_10927,N_10711);
nand U11071 (N_11071,N_10731,N_10671);
nand U11072 (N_11072,N_10642,N_10770);
or U11073 (N_11073,N_10820,N_10598);
nand U11074 (N_11074,N_10964,N_10905);
nor U11075 (N_11075,N_10867,N_10991);
and U11076 (N_11076,N_10623,N_10657);
nor U11077 (N_11077,N_10753,N_10868);
nand U11078 (N_11078,N_10901,N_10669);
nor U11079 (N_11079,N_10706,N_10850);
nand U11080 (N_11080,N_10987,N_10771);
nand U11081 (N_11081,N_10648,N_10772);
xnor U11082 (N_11082,N_10781,N_10606);
nor U11083 (N_11083,N_10865,N_10702);
nand U11084 (N_11084,N_10522,N_10873);
nand U11085 (N_11085,N_10541,N_10686);
and U11086 (N_11086,N_10794,N_10650);
xnor U11087 (N_11087,N_10566,N_10608);
or U11088 (N_11088,N_10719,N_10610);
and U11089 (N_11089,N_10543,N_10807);
nor U11090 (N_11090,N_10653,N_10802);
and U11091 (N_11091,N_10967,N_10513);
and U11092 (N_11092,N_10814,N_10670);
xnor U11093 (N_11093,N_10924,N_10803);
or U11094 (N_11094,N_10915,N_10945);
nand U11095 (N_11095,N_10823,N_10682);
and U11096 (N_11096,N_10795,N_10604);
xor U11097 (N_11097,N_10976,N_10769);
or U11098 (N_11098,N_10884,N_10528);
nor U11099 (N_11099,N_10930,N_10615);
nand U11100 (N_11100,N_10935,N_10546);
or U11101 (N_11101,N_10779,N_10511);
or U11102 (N_11102,N_10830,N_10844);
or U11103 (N_11103,N_10773,N_10592);
nor U11104 (N_11104,N_10762,N_10869);
nor U11105 (N_11105,N_10892,N_10676);
or U11106 (N_11106,N_10949,N_10832);
or U11107 (N_11107,N_10600,N_10632);
nand U11108 (N_11108,N_10960,N_10819);
nor U11109 (N_11109,N_10980,N_10985);
xnor U11110 (N_11110,N_10605,N_10911);
nand U11111 (N_11111,N_10660,N_10567);
xnor U11112 (N_11112,N_10663,N_10689);
nand U11113 (N_11113,N_10904,N_10638);
nor U11114 (N_11114,N_10594,N_10668);
nand U11115 (N_11115,N_10611,N_10741);
xnor U11116 (N_11116,N_10621,N_10851);
xnor U11117 (N_11117,N_10883,N_10569);
nand U11118 (N_11118,N_10672,N_10864);
or U11119 (N_11119,N_10732,N_10887);
and U11120 (N_11120,N_10920,N_10599);
or U11121 (N_11121,N_10532,N_10886);
nand U11122 (N_11122,N_10975,N_10720);
nand U11123 (N_11123,N_10941,N_10996);
xor U11124 (N_11124,N_10737,N_10692);
nand U11125 (N_11125,N_10619,N_10888);
or U11126 (N_11126,N_10758,N_10718);
and U11127 (N_11127,N_10784,N_10799);
or U11128 (N_11128,N_10972,N_10961);
xor U11129 (N_11129,N_10626,N_10729);
or U11130 (N_11130,N_10969,N_10722);
nand U11131 (N_11131,N_10854,N_10847);
nand U11132 (N_11132,N_10829,N_10896);
and U11133 (N_11133,N_10778,N_10973);
or U11134 (N_11134,N_10796,N_10726);
xor U11135 (N_11135,N_10745,N_10523);
nor U11136 (N_11136,N_10767,N_10917);
nor U11137 (N_11137,N_10981,N_10763);
nand U11138 (N_11138,N_10876,N_10866);
or U11139 (N_11139,N_10932,N_10593);
and U11140 (N_11140,N_10798,N_10700);
and U11141 (N_11141,N_10789,N_10986);
or U11142 (N_11142,N_10564,N_10559);
nand U11143 (N_11143,N_10549,N_10944);
nor U11144 (N_11144,N_10667,N_10534);
or U11145 (N_11145,N_10805,N_10698);
nand U11146 (N_11146,N_10995,N_10938);
or U11147 (N_11147,N_10679,N_10852);
and U11148 (N_11148,N_10992,N_10573);
nor U11149 (N_11149,N_10725,N_10687);
or U11150 (N_11150,N_10912,N_10693);
nand U11151 (N_11151,N_10786,N_10665);
nand U11152 (N_11152,N_10697,N_10813);
nand U11153 (N_11153,N_10557,N_10533);
and U11154 (N_11154,N_10894,N_10797);
xor U11155 (N_11155,N_10630,N_10738);
and U11156 (N_11156,N_10565,N_10936);
nor U11157 (N_11157,N_10957,N_10590);
nand U11158 (N_11158,N_10897,N_10968);
xor U11159 (N_11159,N_10613,N_10882);
and U11160 (N_11160,N_10755,N_10624);
xnor U11161 (N_11161,N_10871,N_10910);
nand U11162 (N_11162,N_10891,N_10510);
nand U11163 (N_11163,N_10955,N_10822);
and U11164 (N_11164,N_10646,N_10742);
xnor U11165 (N_11165,N_10988,N_10916);
nor U11166 (N_11166,N_10821,N_10759);
xnor U11167 (N_11167,N_10574,N_10751);
or U11168 (N_11168,N_10675,N_10757);
or U11169 (N_11169,N_10505,N_10518);
nor U11170 (N_11170,N_10848,N_10748);
nor U11171 (N_11171,N_10586,N_10531);
or U11172 (N_11172,N_10661,N_10504);
nor U11173 (N_11173,N_10839,N_10696);
and U11174 (N_11174,N_10500,N_10793);
or U11175 (N_11175,N_10547,N_10607);
nor U11176 (N_11176,N_10750,N_10999);
xor U11177 (N_11177,N_10817,N_10925);
nand U11178 (N_11178,N_10943,N_10662);
nor U11179 (N_11179,N_10928,N_10855);
nand U11180 (N_11180,N_10900,N_10634);
or U11181 (N_11181,N_10728,N_10937);
nor U11182 (N_11182,N_10940,N_10921);
xor U11183 (N_11183,N_10838,N_10508);
xor U11184 (N_11184,N_10580,N_10530);
and U11185 (N_11185,N_10933,N_10760);
nand U11186 (N_11186,N_10691,N_10651);
nor U11187 (N_11187,N_10749,N_10684);
nor U11188 (N_11188,N_10609,N_10885);
nor U11189 (N_11189,N_10774,N_10951);
or U11190 (N_11190,N_10655,N_10507);
xnor U11191 (N_11191,N_10846,N_10637);
nor U11192 (N_11192,N_10874,N_10631);
or U11193 (N_11193,N_10512,N_10859);
xnor U11194 (N_11194,N_10982,N_10509);
xnor U11195 (N_11195,N_10542,N_10647);
or U11196 (N_11196,N_10890,N_10978);
or U11197 (N_11197,N_10825,N_10747);
nor U11198 (N_11198,N_10909,N_10768);
and U11199 (N_11199,N_10863,N_10736);
and U11200 (N_11200,N_10695,N_10723);
nor U11201 (N_11201,N_10640,N_10842);
xor U11202 (N_11202,N_10579,N_10527);
nand U11203 (N_11203,N_10601,N_10849);
nor U11204 (N_11204,N_10544,N_10713);
or U11205 (N_11205,N_10587,N_10954);
and U11206 (N_11206,N_10843,N_10588);
nor U11207 (N_11207,N_10652,N_10545);
or U11208 (N_11208,N_10570,N_10746);
or U11209 (N_11209,N_10617,N_10535);
and U11210 (N_11210,N_10906,N_10947);
nor U11211 (N_11211,N_10521,N_10893);
nand U11212 (N_11212,N_10556,N_10620);
and U11213 (N_11213,N_10775,N_10551);
and U11214 (N_11214,N_10724,N_10659);
nand U11215 (N_11215,N_10824,N_10520);
nand U11216 (N_11216,N_10907,N_10683);
or U11217 (N_11217,N_10539,N_10563);
or U11218 (N_11218,N_10922,N_10568);
xnor U11219 (N_11219,N_10815,N_10919);
xnor U11220 (N_11220,N_10560,N_10703);
or U11221 (N_11221,N_10582,N_10622);
and U11222 (N_11222,N_10979,N_10948);
and U11223 (N_11223,N_10561,N_10826);
or U11224 (N_11224,N_10780,N_10831);
and U11225 (N_11225,N_10956,N_10602);
nor U11226 (N_11226,N_10690,N_10914);
or U11227 (N_11227,N_10828,N_10801);
xnor U11228 (N_11228,N_10879,N_10804);
and U11229 (N_11229,N_10529,N_10578);
nor U11230 (N_11230,N_10730,N_10984);
nand U11231 (N_11231,N_10616,N_10899);
xor U11232 (N_11232,N_10872,N_10878);
nor U11233 (N_11233,N_10553,N_10970);
or U11234 (N_11234,N_10525,N_10680);
and U11235 (N_11235,N_10783,N_10913);
or U11236 (N_11236,N_10681,N_10950);
or U11237 (N_11237,N_10712,N_10998);
nor U11238 (N_11238,N_10627,N_10714);
nand U11239 (N_11239,N_10918,N_10552);
nor U11240 (N_11240,N_10782,N_10633);
or U11241 (N_11241,N_10818,N_10709);
and U11242 (N_11242,N_10717,N_10625);
nor U11243 (N_11243,N_10959,N_10581);
and U11244 (N_11244,N_10584,N_10790);
and U11245 (N_11245,N_10656,N_10678);
nor U11246 (N_11246,N_10898,N_10658);
xor U11247 (N_11247,N_10939,N_10877);
or U11248 (N_11248,N_10727,N_10735);
nor U11249 (N_11249,N_10734,N_10840);
nor U11250 (N_11250,N_10649,N_10856);
nand U11251 (N_11251,N_10966,N_10948);
nor U11252 (N_11252,N_10885,N_10590);
nor U11253 (N_11253,N_10507,N_10968);
xnor U11254 (N_11254,N_10750,N_10539);
nor U11255 (N_11255,N_10732,N_10627);
nor U11256 (N_11256,N_10870,N_10970);
nand U11257 (N_11257,N_10592,N_10981);
nand U11258 (N_11258,N_10683,N_10894);
nand U11259 (N_11259,N_10918,N_10841);
and U11260 (N_11260,N_10764,N_10694);
xor U11261 (N_11261,N_10592,N_10584);
and U11262 (N_11262,N_10784,N_10547);
or U11263 (N_11263,N_10950,N_10867);
nor U11264 (N_11264,N_10914,N_10942);
and U11265 (N_11265,N_10676,N_10662);
nor U11266 (N_11266,N_10537,N_10921);
nand U11267 (N_11267,N_10788,N_10697);
and U11268 (N_11268,N_10703,N_10908);
nand U11269 (N_11269,N_10987,N_10709);
nand U11270 (N_11270,N_10761,N_10938);
and U11271 (N_11271,N_10907,N_10726);
nor U11272 (N_11272,N_10670,N_10771);
nor U11273 (N_11273,N_10615,N_10956);
nand U11274 (N_11274,N_10807,N_10966);
nor U11275 (N_11275,N_10676,N_10852);
and U11276 (N_11276,N_10911,N_10805);
xor U11277 (N_11277,N_10619,N_10571);
or U11278 (N_11278,N_10925,N_10731);
and U11279 (N_11279,N_10695,N_10538);
nor U11280 (N_11280,N_10583,N_10810);
or U11281 (N_11281,N_10951,N_10917);
and U11282 (N_11282,N_10966,N_10828);
xor U11283 (N_11283,N_10506,N_10817);
nor U11284 (N_11284,N_10996,N_10647);
nand U11285 (N_11285,N_10541,N_10617);
or U11286 (N_11286,N_10554,N_10928);
or U11287 (N_11287,N_10890,N_10530);
nor U11288 (N_11288,N_10788,N_10871);
and U11289 (N_11289,N_10617,N_10722);
nor U11290 (N_11290,N_10512,N_10954);
nand U11291 (N_11291,N_10641,N_10662);
nor U11292 (N_11292,N_10946,N_10595);
nor U11293 (N_11293,N_10515,N_10990);
nor U11294 (N_11294,N_10956,N_10867);
and U11295 (N_11295,N_10677,N_10917);
or U11296 (N_11296,N_10964,N_10612);
or U11297 (N_11297,N_10767,N_10927);
or U11298 (N_11298,N_10544,N_10960);
nor U11299 (N_11299,N_10840,N_10635);
and U11300 (N_11300,N_10686,N_10692);
nor U11301 (N_11301,N_10860,N_10593);
nand U11302 (N_11302,N_10917,N_10681);
nor U11303 (N_11303,N_10633,N_10636);
xnor U11304 (N_11304,N_10912,N_10658);
or U11305 (N_11305,N_10561,N_10713);
xor U11306 (N_11306,N_10668,N_10898);
nand U11307 (N_11307,N_10596,N_10863);
or U11308 (N_11308,N_10530,N_10808);
nand U11309 (N_11309,N_10694,N_10954);
nand U11310 (N_11310,N_10896,N_10993);
and U11311 (N_11311,N_10675,N_10701);
xnor U11312 (N_11312,N_10526,N_10883);
nor U11313 (N_11313,N_10653,N_10678);
or U11314 (N_11314,N_10936,N_10643);
nor U11315 (N_11315,N_10719,N_10736);
or U11316 (N_11316,N_10588,N_10567);
nand U11317 (N_11317,N_10763,N_10537);
and U11318 (N_11318,N_10793,N_10867);
xnor U11319 (N_11319,N_10786,N_10941);
or U11320 (N_11320,N_10650,N_10879);
or U11321 (N_11321,N_10552,N_10713);
nor U11322 (N_11322,N_10697,N_10769);
or U11323 (N_11323,N_10867,N_10662);
nor U11324 (N_11324,N_10661,N_10813);
nand U11325 (N_11325,N_10648,N_10529);
xnor U11326 (N_11326,N_10992,N_10804);
and U11327 (N_11327,N_10704,N_10659);
xnor U11328 (N_11328,N_10704,N_10987);
and U11329 (N_11329,N_10572,N_10584);
nand U11330 (N_11330,N_10626,N_10744);
or U11331 (N_11331,N_10744,N_10977);
or U11332 (N_11332,N_10734,N_10567);
or U11333 (N_11333,N_10563,N_10949);
xor U11334 (N_11334,N_10563,N_10984);
nor U11335 (N_11335,N_10517,N_10555);
xor U11336 (N_11336,N_10550,N_10890);
or U11337 (N_11337,N_10542,N_10986);
or U11338 (N_11338,N_10513,N_10778);
xor U11339 (N_11339,N_10728,N_10657);
xnor U11340 (N_11340,N_10663,N_10901);
nand U11341 (N_11341,N_10759,N_10810);
or U11342 (N_11342,N_10594,N_10603);
and U11343 (N_11343,N_10511,N_10665);
and U11344 (N_11344,N_10808,N_10632);
nand U11345 (N_11345,N_10993,N_10618);
or U11346 (N_11346,N_10686,N_10730);
nand U11347 (N_11347,N_10569,N_10927);
nand U11348 (N_11348,N_10746,N_10623);
nor U11349 (N_11349,N_10573,N_10761);
or U11350 (N_11350,N_10799,N_10806);
and U11351 (N_11351,N_10500,N_10798);
and U11352 (N_11352,N_10959,N_10880);
nand U11353 (N_11353,N_10586,N_10969);
and U11354 (N_11354,N_10549,N_10875);
xnor U11355 (N_11355,N_10841,N_10682);
nand U11356 (N_11356,N_10774,N_10514);
nand U11357 (N_11357,N_10796,N_10763);
nand U11358 (N_11358,N_10898,N_10553);
and U11359 (N_11359,N_10749,N_10960);
nand U11360 (N_11360,N_10559,N_10549);
or U11361 (N_11361,N_10957,N_10620);
xnor U11362 (N_11362,N_10978,N_10832);
and U11363 (N_11363,N_10879,N_10801);
xor U11364 (N_11364,N_10736,N_10505);
nand U11365 (N_11365,N_10709,N_10816);
and U11366 (N_11366,N_10554,N_10924);
and U11367 (N_11367,N_10758,N_10582);
nand U11368 (N_11368,N_10717,N_10605);
nand U11369 (N_11369,N_10973,N_10898);
and U11370 (N_11370,N_10790,N_10710);
nor U11371 (N_11371,N_10930,N_10709);
or U11372 (N_11372,N_10907,N_10858);
or U11373 (N_11373,N_10706,N_10882);
nand U11374 (N_11374,N_10863,N_10769);
and U11375 (N_11375,N_10988,N_10923);
xnor U11376 (N_11376,N_10853,N_10887);
xor U11377 (N_11377,N_10670,N_10891);
nor U11378 (N_11378,N_10515,N_10660);
nand U11379 (N_11379,N_10625,N_10948);
and U11380 (N_11380,N_10649,N_10815);
or U11381 (N_11381,N_10958,N_10542);
xor U11382 (N_11382,N_10683,N_10843);
nand U11383 (N_11383,N_10615,N_10981);
nand U11384 (N_11384,N_10943,N_10960);
or U11385 (N_11385,N_10933,N_10619);
nand U11386 (N_11386,N_10710,N_10984);
nor U11387 (N_11387,N_10843,N_10890);
or U11388 (N_11388,N_10640,N_10894);
xnor U11389 (N_11389,N_10695,N_10543);
xor U11390 (N_11390,N_10998,N_10600);
and U11391 (N_11391,N_10768,N_10855);
or U11392 (N_11392,N_10765,N_10580);
or U11393 (N_11393,N_10584,N_10606);
nand U11394 (N_11394,N_10797,N_10776);
xnor U11395 (N_11395,N_10859,N_10860);
and U11396 (N_11396,N_10747,N_10897);
and U11397 (N_11397,N_10719,N_10975);
nor U11398 (N_11398,N_10985,N_10503);
and U11399 (N_11399,N_10810,N_10937);
and U11400 (N_11400,N_10533,N_10983);
nor U11401 (N_11401,N_10633,N_10537);
xnor U11402 (N_11402,N_10732,N_10689);
xor U11403 (N_11403,N_10661,N_10738);
or U11404 (N_11404,N_10869,N_10542);
nor U11405 (N_11405,N_10986,N_10843);
nand U11406 (N_11406,N_10828,N_10614);
nand U11407 (N_11407,N_10753,N_10811);
or U11408 (N_11408,N_10568,N_10946);
or U11409 (N_11409,N_10978,N_10636);
nand U11410 (N_11410,N_10542,N_10641);
xor U11411 (N_11411,N_10548,N_10751);
and U11412 (N_11412,N_10900,N_10694);
nand U11413 (N_11413,N_10657,N_10981);
and U11414 (N_11414,N_10931,N_10884);
nand U11415 (N_11415,N_10567,N_10634);
or U11416 (N_11416,N_10996,N_10545);
nand U11417 (N_11417,N_10945,N_10612);
nand U11418 (N_11418,N_10979,N_10916);
nor U11419 (N_11419,N_10944,N_10619);
nand U11420 (N_11420,N_10798,N_10843);
xor U11421 (N_11421,N_10549,N_10550);
nand U11422 (N_11422,N_10911,N_10883);
xnor U11423 (N_11423,N_10537,N_10542);
nor U11424 (N_11424,N_10541,N_10675);
xor U11425 (N_11425,N_10651,N_10742);
or U11426 (N_11426,N_10665,N_10625);
nand U11427 (N_11427,N_10743,N_10685);
and U11428 (N_11428,N_10578,N_10716);
nor U11429 (N_11429,N_10864,N_10879);
nor U11430 (N_11430,N_10664,N_10892);
nand U11431 (N_11431,N_10550,N_10518);
and U11432 (N_11432,N_10835,N_10571);
or U11433 (N_11433,N_10909,N_10584);
nand U11434 (N_11434,N_10880,N_10865);
nand U11435 (N_11435,N_10527,N_10808);
nor U11436 (N_11436,N_10523,N_10860);
nor U11437 (N_11437,N_10608,N_10881);
nor U11438 (N_11438,N_10847,N_10749);
nor U11439 (N_11439,N_10890,N_10935);
nor U11440 (N_11440,N_10526,N_10995);
or U11441 (N_11441,N_10591,N_10717);
xnor U11442 (N_11442,N_10671,N_10733);
or U11443 (N_11443,N_10889,N_10797);
xor U11444 (N_11444,N_10969,N_10688);
nand U11445 (N_11445,N_10743,N_10786);
nand U11446 (N_11446,N_10996,N_10837);
nand U11447 (N_11447,N_10962,N_10867);
xnor U11448 (N_11448,N_10942,N_10587);
nand U11449 (N_11449,N_10806,N_10543);
nand U11450 (N_11450,N_10863,N_10917);
and U11451 (N_11451,N_10529,N_10699);
nand U11452 (N_11452,N_10796,N_10786);
nand U11453 (N_11453,N_10910,N_10859);
nor U11454 (N_11454,N_10817,N_10861);
or U11455 (N_11455,N_10627,N_10521);
and U11456 (N_11456,N_10835,N_10906);
xnor U11457 (N_11457,N_10651,N_10980);
nor U11458 (N_11458,N_10680,N_10912);
nor U11459 (N_11459,N_10559,N_10751);
xor U11460 (N_11460,N_10761,N_10675);
xnor U11461 (N_11461,N_10848,N_10977);
and U11462 (N_11462,N_10514,N_10674);
xnor U11463 (N_11463,N_10634,N_10809);
or U11464 (N_11464,N_10620,N_10790);
or U11465 (N_11465,N_10791,N_10862);
nor U11466 (N_11466,N_10914,N_10907);
nand U11467 (N_11467,N_10502,N_10757);
nand U11468 (N_11468,N_10644,N_10540);
xor U11469 (N_11469,N_10840,N_10946);
or U11470 (N_11470,N_10858,N_10558);
or U11471 (N_11471,N_10786,N_10977);
nor U11472 (N_11472,N_10843,N_10620);
xor U11473 (N_11473,N_10704,N_10887);
and U11474 (N_11474,N_10993,N_10539);
nand U11475 (N_11475,N_10739,N_10635);
nand U11476 (N_11476,N_10833,N_10858);
nor U11477 (N_11477,N_10630,N_10572);
nand U11478 (N_11478,N_10845,N_10889);
or U11479 (N_11479,N_10759,N_10954);
nor U11480 (N_11480,N_10863,N_10913);
nand U11481 (N_11481,N_10618,N_10760);
nor U11482 (N_11482,N_10753,N_10799);
nand U11483 (N_11483,N_10712,N_10737);
nor U11484 (N_11484,N_10973,N_10698);
nor U11485 (N_11485,N_10660,N_10874);
nand U11486 (N_11486,N_10983,N_10553);
xor U11487 (N_11487,N_10924,N_10766);
or U11488 (N_11488,N_10889,N_10583);
xnor U11489 (N_11489,N_10682,N_10741);
or U11490 (N_11490,N_10958,N_10885);
or U11491 (N_11491,N_10642,N_10748);
nor U11492 (N_11492,N_10564,N_10960);
nand U11493 (N_11493,N_10701,N_10724);
and U11494 (N_11494,N_10856,N_10633);
xnor U11495 (N_11495,N_10586,N_10901);
nand U11496 (N_11496,N_10552,N_10856);
or U11497 (N_11497,N_10628,N_10514);
or U11498 (N_11498,N_10860,N_10781);
or U11499 (N_11499,N_10530,N_10960);
xor U11500 (N_11500,N_11468,N_11006);
nand U11501 (N_11501,N_11264,N_11139);
nand U11502 (N_11502,N_11229,N_11277);
nor U11503 (N_11503,N_11271,N_11402);
nand U11504 (N_11504,N_11181,N_11392);
or U11505 (N_11505,N_11217,N_11251);
nand U11506 (N_11506,N_11157,N_11457);
or U11507 (N_11507,N_11021,N_11499);
xor U11508 (N_11508,N_11249,N_11494);
nand U11509 (N_11509,N_11484,N_11481);
xor U11510 (N_11510,N_11309,N_11322);
nand U11511 (N_11511,N_11483,N_11199);
and U11512 (N_11512,N_11190,N_11095);
nor U11513 (N_11513,N_11103,N_11474);
xor U11514 (N_11514,N_11220,N_11172);
and U11515 (N_11515,N_11128,N_11147);
or U11516 (N_11516,N_11127,N_11153);
nand U11517 (N_11517,N_11441,N_11071);
or U11518 (N_11518,N_11206,N_11155);
and U11519 (N_11519,N_11299,N_11390);
nand U11520 (N_11520,N_11102,N_11384);
xnor U11521 (N_11521,N_11228,N_11090);
and U11522 (N_11522,N_11209,N_11218);
and U11523 (N_11523,N_11370,N_11182);
nand U11524 (N_11524,N_11412,N_11230);
or U11525 (N_11525,N_11116,N_11174);
xnor U11526 (N_11526,N_11327,N_11288);
xor U11527 (N_11527,N_11242,N_11343);
or U11528 (N_11528,N_11137,N_11238);
and U11529 (N_11529,N_11156,N_11107);
or U11530 (N_11530,N_11247,N_11362);
or U11531 (N_11531,N_11383,N_11083);
and U11532 (N_11532,N_11074,N_11187);
and U11533 (N_11533,N_11145,N_11316);
nand U11534 (N_11534,N_11165,N_11447);
nand U11535 (N_11535,N_11487,N_11196);
and U11536 (N_11536,N_11036,N_11478);
and U11537 (N_11537,N_11120,N_11248);
xor U11538 (N_11538,N_11275,N_11075);
or U11539 (N_11539,N_11476,N_11108);
or U11540 (N_11540,N_11246,N_11261);
or U11541 (N_11541,N_11466,N_11104);
xor U11542 (N_11542,N_11438,N_11212);
nor U11543 (N_11543,N_11378,N_11049);
xnor U11544 (N_11544,N_11197,N_11284);
or U11545 (N_11545,N_11428,N_11141);
nor U11546 (N_11546,N_11078,N_11339);
nand U11547 (N_11547,N_11342,N_11335);
xor U11548 (N_11548,N_11416,N_11471);
nand U11549 (N_11549,N_11365,N_11114);
and U11550 (N_11550,N_11162,N_11056);
and U11551 (N_11551,N_11258,N_11385);
and U11552 (N_11552,N_11082,N_11142);
nor U11553 (N_11553,N_11298,N_11300);
and U11554 (N_11554,N_11255,N_11353);
and U11555 (N_11555,N_11278,N_11051);
xor U11556 (N_11556,N_11057,N_11191);
xor U11557 (N_11557,N_11368,N_11409);
and U11558 (N_11558,N_11444,N_11380);
xor U11559 (N_11559,N_11411,N_11475);
xnor U11560 (N_11560,N_11415,N_11280);
nand U11561 (N_11561,N_11017,N_11164);
nand U11562 (N_11562,N_11241,N_11319);
nor U11563 (N_11563,N_11450,N_11245);
nand U11564 (N_11564,N_11035,N_11010);
nor U11565 (N_11565,N_11138,N_11042);
and U11566 (N_11566,N_11031,N_11143);
and U11567 (N_11567,N_11014,N_11211);
nand U11568 (N_11568,N_11347,N_11038);
and U11569 (N_11569,N_11202,N_11398);
nor U11570 (N_11570,N_11132,N_11223);
nor U11571 (N_11571,N_11427,N_11367);
xnor U11572 (N_11572,N_11391,N_11420);
nor U11573 (N_11573,N_11240,N_11123);
and U11574 (N_11574,N_11019,N_11016);
xnor U11575 (N_11575,N_11344,N_11423);
and U11576 (N_11576,N_11413,N_11281);
or U11577 (N_11577,N_11023,N_11237);
or U11578 (N_11578,N_11158,N_11296);
nor U11579 (N_11579,N_11429,N_11033);
xnor U11580 (N_11580,N_11233,N_11414);
xnor U11581 (N_11581,N_11080,N_11399);
nand U11582 (N_11582,N_11067,N_11331);
nor U11583 (N_11583,N_11363,N_11163);
and U11584 (N_11584,N_11315,N_11183);
xnor U11585 (N_11585,N_11210,N_11109);
nand U11586 (N_11586,N_11081,N_11008);
nor U11587 (N_11587,N_11336,N_11216);
xnor U11588 (N_11588,N_11062,N_11286);
nand U11589 (N_11589,N_11096,N_11348);
xor U11590 (N_11590,N_11394,N_11061);
xor U11591 (N_11591,N_11334,N_11159);
nor U11592 (N_11592,N_11397,N_11152);
and U11593 (N_11593,N_11151,N_11100);
or U11594 (N_11594,N_11352,N_11290);
and U11595 (N_11595,N_11294,N_11040);
nand U11596 (N_11596,N_11333,N_11360);
nor U11597 (N_11597,N_11122,N_11320);
nand U11598 (N_11598,N_11025,N_11207);
nor U11599 (N_11599,N_11028,N_11168);
and U11600 (N_11600,N_11118,N_11171);
xnor U11601 (N_11601,N_11140,N_11452);
nand U11602 (N_11602,N_11305,N_11119);
nor U11603 (N_11603,N_11015,N_11417);
and U11604 (N_11604,N_11454,N_11318);
and U11605 (N_11605,N_11375,N_11192);
or U11606 (N_11606,N_11403,N_11404);
or U11607 (N_11607,N_11401,N_11214);
and U11608 (N_11608,N_11431,N_11054);
nor U11609 (N_11609,N_11213,N_11069);
nand U11610 (N_11610,N_11002,N_11012);
and U11611 (N_11611,N_11027,N_11265);
and U11612 (N_11612,N_11472,N_11451);
nand U11613 (N_11613,N_11045,N_11272);
and U11614 (N_11614,N_11039,N_11072);
xnor U11615 (N_11615,N_11456,N_11092);
nand U11616 (N_11616,N_11359,N_11124);
nor U11617 (N_11617,N_11201,N_11376);
nor U11618 (N_11618,N_11086,N_11449);
or U11619 (N_11619,N_11356,N_11046);
nor U11620 (N_11620,N_11312,N_11382);
xor U11621 (N_11621,N_11204,N_11110);
and U11622 (N_11622,N_11243,N_11059);
and U11623 (N_11623,N_11303,N_11167);
or U11624 (N_11624,N_11032,N_11313);
nor U11625 (N_11625,N_11133,N_11053);
or U11626 (N_11626,N_11077,N_11173);
or U11627 (N_11627,N_11346,N_11371);
and U11628 (N_11628,N_11358,N_11121);
xnor U11629 (N_11629,N_11232,N_11485);
nor U11630 (N_11630,N_11479,N_11462);
nor U11631 (N_11631,N_11144,N_11482);
xnor U11632 (N_11632,N_11470,N_11160);
xnor U11633 (N_11633,N_11259,N_11222);
and U11634 (N_11634,N_11461,N_11337);
xnor U11635 (N_11635,N_11373,N_11282);
or U11636 (N_11636,N_11136,N_11178);
nor U11637 (N_11637,N_11351,N_11226);
and U11638 (N_11638,N_11266,N_11097);
nor U11639 (N_11639,N_11070,N_11361);
nor U11640 (N_11640,N_11345,N_11166);
and U11641 (N_11641,N_11175,N_11007);
xor U11642 (N_11642,N_11186,N_11089);
nand U11643 (N_11643,N_11490,N_11169);
xor U11644 (N_11644,N_11489,N_11099);
or U11645 (N_11645,N_11250,N_11200);
nor U11646 (N_11646,N_11009,N_11325);
nand U11647 (N_11647,N_11003,N_11185);
nor U11648 (N_11648,N_11068,N_11263);
nand U11649 (N_11649,N_11302,N_11203);
or U11650 (N_11650,N_11386,N_11112);
or U11651 (N_11651,N_11270,N_11446);
or U11652 (N_11652,N_11332,N_11443);
or U11653 (N_11653,N_11440,N_11445);
and U11654 (N_11654,N_11338,N_11195);
nand U11655 (N_11655,N_11437,N_11492);
nand U11656 (N_11656,N_11180,N_11341);
nor U11657 (N_11657,N_11126,N_11306);
and U11658 (N_11658,N_11354,N_11469);
nand U11659 (N_11659,N_11011,N_11491);
or U11660 (N_11660,N_11193,N_11418);
or U11661 (N_11661,N_11330,N_11146);
xor U11662 (N_11662,N_11065,N_11131);
xor U11663 (N_11663,N_11150,N_11439);
nand U11664 (N_11664,N_11355,N_11022);
xor U11665 (N_11665,N_11254,N_11430);
xnor U11666 (N_11666,N_11253,N_11340);
nor U11667 (N_11667,N_11396,N_11366);
and U11668 (N_11668,N_11239,N_11455);
xor U11669 (N_11669,N_11276,N_11111);
nor U11670 (N_11670,N_11292,N_11013);
nor U11671 (N_11671,N_11291,N_11154);
or U11672 (N_11672,N_11297,N_11408);
xor U11673 (N_11673,N_11004,N_11426);
and U11674 (N_11674,N_11091,N_11256);
and U11675 (N_11675,N_11477,N_11020);
or U11676 (N_11676,N_11372,N_11129);
nand U11677 (N_11677,N_11029,N_11349);
xnor U11678 (N_11678,N_11026,N_11149);
nor U11679 (N_11679,N_11001,N_11453);
and U11680 (N_11680,N_11084,N_11377);
and U11681 (N_11681,N_11052,N_11219);
or U11682 (N_11682,N_11486,N_11101);
and U11683 (N_11683,N_11395,N_11442);
xnor U11684 (N_11684,N_11369,N_11221);
and U11685 (N_11685,N_11135,N_11227);
or U11686 (N_11686,N_11106,N_11087);
xor U11687 (N_11687,N_11400,N_11194);
or U11688 (N_11688,N_11208,N_11079);
and U11689 (N_11689,N_11374,N_11262);
or U11690 (N_11690,N_11066,N_11093);
nand U11691 (N_11691,N_11324,N_11018);
or U11692 (N_11692,N_11459,N_11434);
nor U11693 (N_11693,N_11424,N_11274);
and U11694 (N_11694,N_11425,N_11498);
xor U11695 (N_11695,N_11048,N_11497);
and U11696 (N_11696,N_11473,N_11000);
or U11697 (N_11697,N_11301,N_11105);
nor U11698 (N_11698,N_11388,N_11117);
nor U11699 (N_11699,N_11433,N_11495);
nor U11700 (N_11700,N_11410,N_11041);
or U11701 (N_11701,N_11064,N_11463);
or U11702 (N_11702,N_11293,N_11005);
and U11703 (N_11703,N_11115,N_11493);
or U11704 (N_11704,N_11205,N_11422);
xor U11705 (N_11705,N_11269,N_11055);
or U11706 (N_11706,N_11448,N_11179);
xnor U11707 (N_11707,N_11357,N_11252);
nand U11708 (N_11708,N_11381,N_11176);
or U11709 (N_11709,N_11060,N_11224);
xor U11710 (N_11710,N_11198,N_11231);
nand U11711 (N_11711,N_11148,N_11465);
nand U11712 (N_11712,N_11257,N_11113);
nand U11713 (N_11713,N_11043,N_11323);
xor U11714 (N_11714,N_11304,N_11387);
and U11715 (N_11715,N_11225,N_11268);
nand U11716 (N_11716,N_11076,N_11044);
nand U11717 (N_11717,N_11406,N_11050);
and U11718 (N_11718,N_11480,N_11350);
nor U11719 (N_11719,N_11405,N_11460);
nand U11720 (N_11720,N_11134,N_11267);
nand U11721 (N_11721,N_11125,N_11189);
xor U11722 (N_11722,N_11279,N_11184);
and U11723 (N_11723,N_11235,N_11435);
and U11724 (N_11724,N_11188,N_11295);
xnor U11725 (N_11725,N_11310,N_11307);
or U11726 (N_11726,N_11037,N_11329);
or U11727 (N_11727,N_11326,N_11030);
nor U11728 (N_11728,N_11432,N_11317);
and U11729 (N_11729,N_11287,N_11436);
nor U11730 (N_11730,N_11215,N_11311);
or U11731 (N_11731,N_11260,N_11458);
or U11732 (N_11732,N_11308,N_11364);
xnor U11733 (N_11733,N_11034,N_11488);
nand U11734 (N_11734,N_11098,N_11177);
and U11735 (N_11735,N_11467,N_11393);
or U11736 (N_11736,N_11063,N_11088);
nand U11737 (N_11737,N_11273,N_11314);
xnor U11738 (N_11738,N_11328,N_11464);
nor U11739 (N_11739,N_11289,N_11389);
or U11740 (N_11740,N_11496,N_11285);
or U11741 (N_11741,N_11407,N_11170);
nand U11742 (N_11742,N_11419,N_11236);
xnor U11743 (N_11743,N_11130,N_11094);
xor U11744 (N_11744,N_11058,N_11379);
nor U11745 (N_11745,N_11073,N_11047);
or U11746 (N_11746,N_11024,N_11234);
and U11747 (N_11747,N_11244,N_11161);
and U11748 (N_11748,N_11085,N_11283);
xnor U11749 (N_11749,N_11321,N_11421);
or U11750 (N_11750,N_11417,N_11381);
and U11751 (N_11751,N_11348,N_11462);
or U11752 (N_11752,N_11332,N_11480);
nand U11753 (N_11753,N_11361,N_11251);
xor U11754 (N_11754,N_11344,N_11370);
xnor U11755 (N_11755,N_11490,N_11461);
nor U11756 (N_11756,N_11062,N_11210);
and U11757 (N_11757,N_11180,N_11060);
nand U11758 (N_11758,N_11071,N_11085);
or U11759 (N_11759,N_11211,N_11445);
and U11760 (N_11760,N_11104,N_11066);
nor U11761 (N_11761,N_11330,N_11009);
nand U11762 (N_11762,N_11321,N_11104);
nand U11763 (N_11763,N_11248,N_11347);
xor U11764 (N_11764,N_11180,N_11136);
or U11765 (N_11765,N_11073,N_11318);
nand U11766 (N_11766,N_11074,N_11112);
or U11767 (N_11767,N_11227,N_11051);
nor U11768 (N_11768,N_11092,N_11331);
and U11769 (N_11769,N_11310,N_11265);
nor U11770 (N_11770,N_11022,N_11172);
nor U11771 (N_11771,N_11223,N_11261);
and U11772 (N_11772,N_11026,N_11444);
xnor U11773 (N_11773,N_11361,N_11261);
or U11774 (N_11774,N_11107,N_11333);
xor U11775 (N_11775,N_11198,N_11453);
nor U11776 (N_11776,N_11265,N_11280);
nand U11777 (N_11777,N_11287,N_11299);
or U11778 (N_11778,N_11472,N_11072);
xnor U11779 (N_11779,N_11210,N_11123);
xor U11780 (N_11780,N_11055,N_11408);
nand U11781 (N_11781,N_11156,N_11325);
and U11782 (N_11782,N_11332,N_11431);
nor U11783 (N_11783,N_11110,N_11318);
nor U11784 (N_11784,N_11478,N_11106);
nand U11785 (N_11785,N_11120,N_11340);
xor U11786 (N_11786,N_11071,N_11476);
nand U11787 (N_11787,N_11243,N_11469);
nand U11788 (N_11788,N_11490,N_11422);
or U11789 (N_11789,N_11315,N_11441);
xor U11790 (N_11790,N_11032,N_11303);
xor U11791 (N_11791,N_11236,N_11087);
or U11792 (N_11792,N_11036,N_11153);
and U11793 (N_11793,N_11285,N_11113);
or U11794 (N_11794,N_11262,N_11297);
nor U11795 (N_11795,N_11221,N_11096);
and U11796 (N_11796,N_11340,N_11424);
nor U11797 (N_11797,N_11164,N_11185);
nand U11798 (N_11798,N_11465,N_11021);
nor U11799 (N_11799,N_11266,N_11148);
and U11800 (N_11800,N_11425,N_11340);
xnor U11801 (N_11801,N_11062,N_11048);
or U11802 (N_11802,N_11451,N_11145);
nor U11803 (N_11803,N_11118,N_11194);
xnor U11804 (N_11804,N_11466,N_11105);
xnor U11805 (N_11805,N_11024,N_11353);
nand U11806 (N_11806,N_11055,N_11292);
xnor U11807 (N_11807,N_11206,N_11348);
nor U11808 (N_11808,N_11311,N_11117);
nor U11809 (N_11809,N_11274,N_11234);
nor U11810 (N_11810,N_11331,N_11172);
xnor U11811 (N_11811,N_11020,N_11284);
or U11812 (N_11812,N_11383,N_11327);
nand U11813 (N_11813,N_11052,N_11338);
and U11814 (N_11814,N_11018,N_11197);
or U11815 (N_11815,N_11455,N_11493);
xnor U11816 (N_11816,N_11015,N_11110);
nand U11817 (N_11817,N_11453,N_11289);
nand U11818 (N_11818,N_11254,N_11255);
xor U11819 (N_11819,N_11247,N_11058);
xnor U11820 (N_11820,N_11161,N_11432);
or U11821 (N_11821,N_11448,N_11427);
xor U11822 (N_11822,N_11144,N_11325);
nand U11823 (N_11823,N_11373,N_11164);
and U11824 (N_11824,N_11137,N_11367);
and U11825 (N_11825,N_11274,N_11235);
or U11826 (N_11826,N_11074,N_11169);
nand U11827 (N_11827,N_11233,N_11431);
and U11828 (N_11828,N_11312,N_11226);
or U11829 (N_11829,N_11234,N_11345);
and U11830 (N_11830,N_11339,N_11199);
and U11831 (N_11831,N_11259,N_11423);
nor U11832 (N_11832,N_11146,N_11038);
and U11833 (N_11833,N_11451,N_11173);
nor U11834 (N_11834,N_11084,N_11130);
or U11835 (N_11835,N_11317,N_11163);
xnor U11836 (N_11836,N_11033,N_11084);
and U11837 (N_11837,N_11306,N_11248);
xor U11838 (N_11838,N_11005,N_11030);
or U11839 (N_11839,N_11033,N_11103);
nor U11840 (N_11840,N_11001,N_11262);
or U11841 (N_11841,N_11033,N_11049);
xnor U11842 (N_11842,N_11029,N_11472);
nand U11843 (N_11843,N_11458,N_11105);
nor U11844 (N_11844,N_11481,N_11344);
xor U11845 (N_11845,N_11271,N_11469);
and U11846 (N_11846,N_11455,N_11260);
xnor U11847 (N_11847,N_11392,N_11060);
and U11848 (N_11848,N_11281,N_11204);
nor U11849 (N_11849,N_11333,N_11270);
nor U11850 (N_11850,N_11455,N_11203);
nand U11851 (N_11851,N_11152,N_11218);
and U11852 (N_11852,N_11493,N_11032);
and U11853 (N_11853,N_11159,N_11384);
or U11854 (N_11854,N_11321,N_11398);
or U11855 (N_11855,N_11363,N_11198);
or U11856 (N_11856,N_11147,N_11202);
nor U11857 (N_11857,N_11475,N_11080);
nor U11858 (N_11858,N_11137,N_11287);
and U11859 (N_11859,N_11211,N_11201);
and U11860 (N_11860,N_11175,N_11301);
nor U11861 (N_11861,N_11410,N_11397);
nand U11862 (N_11862,N_11134,N_11422);
nand U11863 (N_11863,N_11239,N_11048);
nand U11864 (N_11864,N_11015,N_11188);
or U11865 (N_11865,N_11217,N_11407);
nor U11866 (N_11866,N_11098,N_11283);
nand U11867 (N_11867,N_11143,N_11212);
nand U11868 (N_11868,N_11476,N_11495);
nor U11869 (N_11869,N_11010,N_11372);
nor U11870 (N_11870,N_11161,N_11216);
or U11871 (N_11871,N_11082,N_11041);
or U11872 (N_11872,N_11347,N_11237);
nor U11873 (N_11873,N_11054,N_11323);
nand U11874 (N_11874,N_11327,N_11129);
nand U11875 (N_11875,N_11283,N_11199);
xor U11876 (N_11876,N_11306,N_11090);
or U11877 (N_11877,N_11142,N_11448);
nor U11878 (N_11878,N_11154,N_11131);
or U11879 (N_11879,N_11323,N_11264);
nor U11880 (N_11880,N_11192,N_11169);
or U11881 (N_11881,N_11180,N_11333);
xor U11882 (N_11882,N_11321,N_11044);
nand U11883 (N_11883,N_11089,N_11495);
xnor U11884 (N_11884,N_11096,N_11366);
xor U11885 (N_11885,N_11466,N_11297);
xor U11886 (N_11886,N_11347,N_11428);
or U11887 (N_11887,N_11260,N_11281);
xnor U11888 (N_11888,N_11111,N_11399);
nand U11889 (N_11889,N_11493,N_11037);
nor U11890 (N_11890,N_11354,N_11025);
nor U11891 (N_11891,N_11218,N_11090);
and U11892 (N_11892,N_11021,N_11120);
and U11893 (N_11893,N_11298,N_11387);
and U11894 (N_11894,N_11110,N_11042);
and U11895 (N_11895,N_11086,N_11309);
and U11896 (N_11896,N_11024,N_11152);
nand U11897 (N_11897,N_11298,N_11325);
and U11898 (N_11898,N_11129,N_11183);
and U11899 (N_11899,N_11480,N_11346);
and U11900 (N_11900,N_11465,N_11330);
or U11901 (N_11901,N_11254,N_11334);
xnor U11902 (N_11902,N_11474,N_11297);
and U11903 (N_11903,N_11001,N_11145);
and U11904 (N_11904,N_11366,N_11420);
or U11905 (N_11905,N_11367,N_11449);
nor U11906 (N_11906,N_11398,N_11220);
nor U11907 (N_11907,N_11133,N_11315);
nor U11908 (N_11908,N_11132,N_11339);
xnor U11909 (N_11909,N_11103,N_11028);
nor U11910 (N_11910,N_11009,N_11182);
nor U11911 (N_11911,N_11050,N_11288);
nand U11912 (N_11912,N_11349,N_11353);
or U11913 (N_11913,N_11106,N_11421);
and U11914 (N_11914,N_11241,N_11374);
nand U11915 (N_11915,N_11046,N_11088);
or U11916 (N_11916,N_11462,N_11290);
or U11917 (N_11917,N_11259,N_11233);
and U11918 (N_11918,N_11012,N_11440);
nor U11919 (N_11919,N_11189,N_11134);
nand U11920 (N_11920,N_11050,N_11004);
or U11921 (N_11921,N_11283,N_11367);
and U11922 (N_11922,N_11278,N_11012);
and U11923 (N_11923,N_11186,N_11281);
and U11924 (N_11924,N_11353,N_11061);
or U11925 (N_11925,N_11357,N_11058);
xnor U11926 (N_11926,N_11438,N_11432);
nand U11927 (N_11927,N_11215,N_11012);
and U11928 (N_11928,N_11111,N_11059);
xor U11929 (N_11929,N_11012,N_11263);
nor U11930 (N_11930,N_11227,N_11122);
and U11931 (N_11931,N_11052,N_11217);
nor U11932 (N_11932,N_11363,N_11295);
xor U11933 (N_11933,N_11233,N_11012);
and U11934 (N_11934,N_11070,N_11040);
and U11935 (N_11935,N_11279,N_11496);
xnor U11936 (N_11936,N_11279,N_11327);
or U11937 (N_11937,N_11337,N_11472);
nand U11938 (N_11938,N_11228,N_11285);
nand U11939 (N_11939,N_11216,N_11377);
and U11940 (N_11940,N_11341,N_11161);
or U11941 (N_11941,N_11428,N_11025);
xor U11942 (N_11942,N_11253,N_11499);
and U11943 (N_11943,N_11362,N_11054);
nor U11944 (N_11944,N_11298,N_11319);
and U11945 (N_11945,N_11162,N_11270);
nand U11946 (N_11946,N_11383,N_11343);
nand U11947 (N_11947,N_11219,N_11300);
and U11948 (N_11948,N_11323,N_11084);
nand U11949 (N_11949,N_11498,N_11047);
nand U11950 (N_11950,N_11274,N_11386);
nor U11951 (N_11951,N_11383,N_11491);
nand U11952 (N_11952,N_11491,N_11246);
xor U11953 (N_11953,N_11278,N_11201);
nor U11954 (N_11954,N_11163,N_11049);
or U11955 (N_11955,N_11328,N_11252);
nor U11956 (N_11956,N_11381,N_11018);
nor U11957 (N_11957,N_11364,N_11212);
and U11958 (N_11958,N_11068,N_11237);
nand U11959 (N_11959,N_11052,N_11081);
and U11960 (N_11960,N_11206,N_11071);
nand U11961 (N_11961,N_11105,N_11275);
nor U11962 (N_11962,N_11395,N_11116);
nand U11963 (N_11963,N_11276,N_11076);
nand U11964 (N_11964,N_11408,N_11066);
and U11965 (N_11965,N_11486,N_11225);
or U11966 (N_11966,N_11488,N_11461);
nand U11967 (N_11967,N_11492,N_11242);
xnor U11968 (N_11968,N_11268,N_11079);
nand U11969 (N_11969,N_11081,N_11364);
and U11970 (N_11970,N_11154,N_11481);
xor U11971 (N_11971,N_11360,N_11083);
xor U11972 (N_11972,N_11373,N_11470);
nor U11973 (N_11973,N_11305,N_11392);
nand U11974 (N_11974,N_11049,N_11027);
and U11975 (N_11975,N_11389,N_11240);
nand U11976 (N_11976,N_11241,N_11296);
and U11977 (N_11977,N_11377,N_11352);
or U11978 (N_11978,N_11134,N_11314);
nor U11979 (N_11979,N_11062,N_11443);
xnor U11980 (N_11980,N_11050,N_11001);
xor U11981 (N_11981,N_11203,N_11371);
and U11982 (N_11982,N_11464,N_11275);
nor U11983 (N_11983,N_11198,N_11000);
or U11984 (N_11984,N_11259,N_11104);
nor U11985 (N_11985,N_11453,N_11050);
and U11986 (N_11986,N_11382,N_11454);
or U11987 (N_11987,N_11002,N_11231);
and U11988 (N_11988,N_11029,N_11218);
xnor U11989 (N_11989,N_11226,N_11045);
nor U11990 (N_11990,N_11481,N_11128);
xnor U11991 (N_11991,N_11446,N_11298);
xor U11992 (N_11992,N_11315,N_11391);
nor U11993 (N_11993,N_11145,N_11459);
nand U11994 (N_11994,N_11365,N_11130);
and U11995 (N_11995,N_11365,N_11134);
nor U11996 (N_11996,N_11247,N_11293);
xnor U11997 (N_11997,N_11253,N_11114);
and U11998 (N_11998,N_11404,N_11277);
nor U11999 (N_11999,N_11367,N_11291);
and U12000 (N_12000,N_11999,N_11600);
nand U12001 (N_12001,N_11824,N_11865);
and U12002 (N_12002,N_11585,N_11541);
nor U12003 (N_12003,N_11873,N_11722);
nand U12004 (N_12004,N_11870,N_11798);
xor U12005 (N_12005,N_11923,N_11739);
nand U12006 (N_12006,N_11509,N_11614);
nor U12007 (N_12007,N_11639,N_11539);
and U12008 (N_12008,N_11501,N_11975);
nand U12009 (N_12009,N_11616,N_11641);
nand U12010 (N_12010,N_11931,N_11506);
xnor U12011 (N_12011,N_11637,N_11821);
and U12012 (N_12012,N_11591,N_11550);
nand U12013 (N_12013,N_11508,N_11828);
xor U12014 (N_12014,N_11986,N_11933);
xnor U12015 (N_12015,N_11504,N_11738);
or U12016 (N_12016,N_11954,N_11640);
xnor U12017 (N_12017,N_11862,N_11768);
xnor U12018 (N_12018,N_11608,N_11731);
and U12019 (N_12019,N_11645,N_11747);
nor U12020 (N_12020,N_11676,N_11606);
nand U12021 (N_12021,N_11664,N_11932);
nor U12022 (N_12022,N_11609,N_11698);
nor U12023 (N_12023,N_11900,N_11940);
nand U12024 (N_12024,N_11844,N_11612);
xor U12025 (N_12025,N_11813,N_11990);
or U12026 (N_12026,N_11534,N_11961);
xor U12027 (N_12027,N_11989,N_11946);
nor U12028 (N_12028,N_11827,N_11901);
nand U12029 (N_12029,N_11527,N_11959);
xor U12030 (N_12030,N_11835,N_11582);
xnor U12031 (N_12031,N_11950,N_11906);
and U12032 (N_12032,N_11604,N_11719);
nor U12033 (N_12033,N_11708,N_11547);
nand U12034 (N_12034,N_11806,N_11872);
nor U12035 (N_12035,N_11543,N_11701);
or U12036 (N_12036,N_11567,N_11558);
nor U12037 (N_12037,N_11638,N_11973);
nand U12038 (N_12038,N_11800,N_11788);
and U12039 (N_12039,N_11744,N_11758);
or U12040 (N_12040,N_11998,N_11757);
xnor U12041 (N_12041,N_11880,N_11693);
and U12042 (N_12042,N_11847,N_11883);
or U12043 (N_12043,N_11598,N_11692);
nand U12044 (N_12044,N_11575,N_11732);
and U12045 (N_12045,N_11893,N_11678);
or U12046 (N_12046,N_11968,N_11529);
nor U12047 (N_12047,N_11503,N_11790);
nor U12048 (N_12048,N_11659,N_11890);
or U12049 (N_12049,N_11526,N_11636);
nor U12050 (N_12050,N_11648,N_11899);
or U12051 (N_12051,N_11819,N_11624);
and U12052 (N_12052,N_11603,N_11753);
nand U12053 (N_12053,N_11881,N_11670);
or U12054 (N_12054,N_11658,N_11568);
nor U12055 (N_12055,N_11619,N_11628);
and U12056 (N_12056,N_11668,N_11512);
xnor U12057 (N_12057,N_11737,N_11884);
nand U12058 (N_12058,N_11620,N_11796);
nand U12059 (N_12059,N_11680,N_11869);
nand U12060 (N_12060,N_11907,N_11761);
and U12061 (N_12061,N_11660,N_11927);
and U12062 (N_12062,N_11976,N_11977);
xnor U12063 (N_12063,N_11607,N_11948);
or U12064 (N_12064,N_11627,N_11850);
nand U12065 (N_12065,N_11736,N_11833);
or U12066 (N_12066,N_11922,N_11840);
xnor U12067 (N_12067,N_11728,N_11983);
nand U12068 (N_12068,N_11755,N_11661);
xnor U12069 (N_12069,N_11594,N_11588);
and U12070 (N_12070,N_11571,N_11533);
nor U12071 (N_12071,N_11908,N_11854);
or U12072 (N_12072,N_11982,N_11684);
nand U12073 (N_12073,N_11895,N_11666);
nand U12074 (N_12074,N_11832,N_11915);
nand U12075 (N_12075,N_11921,N_11702);
xnor U12076 (N_12076,N_11853,N_11792);
xor U12077 (N_12077,N_11980,N_11584);
nand U12078 (N_12078,N_11803,N_11911);
and U12079 (N_12079,N_11864,N_11958);
nand U12080 (N_12080,N_11694,N_11549);
or U12081 (N_12081,N_11823,N_11793);
nor U12082 (N_12082,N_11651,N_11707);
and U12083 (N_12083,N_11517,N_11996);
nand U12084 (N_12084,N_11733,N_11919);
or U12085 (N_12085,N_11972,N_11595);
xor U12086 (N_12086,N_11689,N_11632);
nand U12087 (N_12087,N_11825,N_11552);
and U12088 (N_12088,N_11776,N_11882);
xnor U12089 (N_12089,N_11841,N_11553);
nand U12090 (N_12090,N_11644,N_11679);
nor U12091 (N_12091,N_11981,N_11804);
or U12092 (N_12092,N_11947,N_11740);
or U12093 (N_12093,N_11723,N_11655);
and U12094 (N_12094,N_11569,N_11889);
and U12095 (N_12095,N_11920,N_11891);
nand U12096 (N_12096,N_11672,N_11576);
xor U12097 (N_12097,N_11978,N_11597);
and U12098 (N_12098,N_11879,N_11530);
or U12099 (N_12099,N_11836,N_11786);
nor U12100 (N_12100,N_11729,N_11918);
nand U12101 (N_12101,N_11617,N_11531);
and U12102 (N_12102,N_11943,N_11802);
and U12103 (N_12103,N_11785,N_11532);
nor U12104 (N_12104,N_11759,N_11580);
and U12105 (N_12105,N_11770,N_11794);
or U12106 (N_12106,N_11671,N_11808);
and U12107 (N_12107,N_11746,N_11626);
xor U12108 (N_12108,N_11867,N_11513);
nor U12109 (N_12109,N_11752,N_11629);
or U12110 (N_12110,N_11683,N_11974);
nor U12111 (N_12111,N_11663,N_11599);
and U12112 (N_12112,N_11767,N_11717);
nor U12113 (N_12113,N_11876,N_11797);
nand U12114 (N_12114,N_11787,N_11713);
or U12115 (N_12115,N_11811,N_11700);
or U12116 (N_12116,N_11763,N_11726);
nor U12117 (N_12117,N_11566,N_11618);
nor U12118 (N_12118,N_11710,N_11749);
and U12119 (N_12119,N_11912,N_11952);
nor U12120 (N_12120,N_11554,N_11938);
and U12121 (N_12121,N_11951,N_11716);
xor U12122 (N_12122,N_11653,N_11818);
xnor U12123 (N_12123,N_11602,N_11985);
nand U12124 (N_12124,N_11748,N_11586);
nor U12125 (N_12125,N_11962,N_11646);
xor U12126 (N_12126,N_11565,N_11557);
xnor U12127 (N_12127,N_11590,N_11681);
or U12128 (N_12128,N_11500,N_11537);
and U12129 (N_12129,N_11855,N_11613);
nand U12130 (N_12130,N_11725,N_11937);
xnor U12131 (N_12131,N_11642,N_11784);
or U12132 (N_12132,N_11874,N_11510);
xnor U12133 (N_12133,N_11942,N_11765);
and U12134 (N_12134,N_11695,N_11944);
or U12135 (N_12135,N_11546,N_11801);
xor U12136 (N_12136,N_11505,N_11631);
nand U12137 (N_12137,N_11718,N_11551);
and U12138 (N_12138,N_11696,N_11789);
or U12139 (N_12139,N_11913,N_11544);
and U12140 (N_12140,N_11542,N_11831);
and U12141 (N_12141,N_11887,N_11894);
nor U12142 (N_12142,N_11814,N_11846);
and U12143 (N_12143,N_11685,N_11745);
or U12144 (N_12144,N_11779,N_11783);
nor U12145 (N_12145,N_11574,N_11843);
nand U12146 (N_12146,N_11605,N_11799);
or U12147 (N_12147,N_11845,N_11878);
or U12148 (N_12148,N_11762,N_11555);
nand U12149 (N_12149,N_11714,N_11967);
xnor U12150 (N_12150,N_11916,N_11564);
and U12151 (N_12151,N_11939,N_11706);
or U12152 (N_12152,N_11704,N_11711);
nor U12153 (N_12153,N_11634,N_11764);
xnor U12154 (N_12154,N_11523,N_11751);
nand U12155 (N_12155,N_11925,N_11610);
and U12156 (N_12156,N_11866,N_11650);
nor U12157 (N_12157,N_11623,N_11992);
or U12158 (N_12158,N_11540,N_11581);
and U12159 (N_12159,N_11817,N_11721);
or U12160 (N_12160,N_11596,N_11511);
and U12161 (N_12161,N_11579,N_11837);
nand U12162 (N_12162,N_11548,N_11720);
and U12163 (N_12163,N_11871,N_11743);
nor U12164 (N_12164,N_11780,N_11697);
or U12165 (N_12165,N_11754,N_11935);
nand U12166 (N_12166,N_11667,N_11652);
or U12167 (N_12167,N_11577,N_11635);
xnor U12168 (N_12168,N_11592,N_11525);
nor U12169 (N_12169,N_11521,N_11795);
and U12170 (N_12170,N_11669,N_11849);
nor U12171 (N_12171,N_11945,N_11934);
xnor U12172 (N_12172,N_11822,N_11910);
nor U12173 (N_12173,N_11699,N_11993);
nand U12174 (N_12174,N_11514,N_11857);
and U12175 (N_12175,N_11677,N_11888);
xor U12176 (N_12176,N_11630,N_11622);
and U12177 (N_12177,N_11791,N_11969);
xnor U12178 (N_12178,N_11987,N_11896);
or U12179 (N_12179,N_11905,N_11649);
nand U12180 (N_12180,N_11928,N_11772);
nand U12181 (N_12181,N_11507,N_11914);
nor U12182 (N_12182,N_11520,N_11665);
and U12183 (N_12183,N_11625,N_11771);
xnor U12184 (N_12184,N_11809,N_11956);
nand U12185 (N_12185,N_11957,N_11675);
nand U12186 (N_12186,N_11522,N_11654);
xnor U12187 (N_12187,N_11774,N_11691);
xor U12188 (N_12188,N_11897,N_11839);
nand U12189 (N_12189,N_11730,N_11593);
xnor U12190 (N_12190,N_11858,N_11656);
or U12191 (N_12191,N_11917,N_11735);
and U12192 (N_12192,N_11515,N_11687);
nand U12193 (N_12193,N_11851,N_11903);
or U12194 (N_12194,N_11615,N_11775);
nand U12195 (N_12195,N_11816,N_11960);
xnor U12196 (N_12196,N_11556,N_11830);
nor U12197 (N_12197,N_11578,N_11773);
and U12198 (N_12198,N_11820,N_11852);
xor U12199 (N_12199,N_11782,N_11705);
or U12200 (N_12200,N_11848,N_11860);
or U12201 (N_12201,N_11561,N_11573);
xor U12202 (N_12202,N_11807,N_11963);
nand U12203 (N_12203,N_11734,N_11984);
xor U12204 (N_12204,N_11750,N_11715);
or U12205 (N_12205,N_11662,N_11904);
nand U12206 (N_12206,N_11861,N_11760);
xor U12207 (N_12207,N_11971,N_11611);
or U12208 (N_12208,N_11995,N_11709);
nor U12209 (N_12209,N_11966,N_11812);
and U12210 (N_12210,N_11842,N_11777);
xnor U12211 (N_12211,N_11815,N_11877);
or U12212 (N_12212,N_11826,N_11587);
nor U12213 (N_12213,N_11875,N_11955);
nand U12214 (N_12214,N_11868,N_11643);
nand U12215 (N_12215,N_11572,N_11930);
xor U12216 (N_12216,N_11781,N_11712);
nand U12217 (N_12217,N_11601,N_11518);
nand U12218 (N_12218,N_11528,N_11657);
xor U12219 (N_12219,N_11892,N_11936);
nand U12220 (N_12220,N_11545,N_11570);
nand U12221 (N_12221,N_11724,N_11756);
nand U12222 (N_12222,N_11991,N_11778);
nand U12223 (N_12223,N_11621,N_11929);
nand U12224 (N_12224,N_11502,N_11965);
nor U12225 (N_12225,N_11562,N_11741);
and U12226 (N_12226,N_11805,N_11536);
xor U12227 (N_12227,N_11810,N_11970);
nor U12228 (N_12228,N_11856,N_11673);
and U12229 (N_12229,N_11690,N_11519);
and U12230 (N_12230,N_11589,N_11703);
and U12231 (N_12231,N_11682,N_11997);
xor U12232 (N_12232,N_11559,N_11516);
xnor U12233 (N_12233,N_11727,N_11898);
or U12234 (N_12234,N_11988,N_11647);
or U12235 (N_12235,N_11885,N_11902);
and U12236 (N_12236,N_11979,N_11538);
and U12237 (N_12237,N_11686,N_11859);
or U12238 (N_12238,N_11834,N_11838);
and U12239 (N_12239,N_11688,N_11886);
nand U12240 (N_12240,N_11964,N_11535);
and U12241 (N_12241,N_11633,N_11829);
and U12242 (N_12242,N_11742,N_11863);
and U12243 (N_12243,N_11994,N_11769);
or U12244 (N_12244,N_11941,N_11583);
nor U12245 (N_12245,N_11524,N_11949);
nand U12246 (N_12246,N_11953,N_11766);
or U12247 (N_12247,N_11563,N_11560);
nand U12248 (N_12248,N_11674,N_11924);
or U12249 (N_12249,N_11909,N_11926);
nand U12250 (N_12250,N_11518,N_11554);
xnor U12251 (N_12251,N_11858,N_11706);
or U12252 (N_12252,N_11785,N_11632);
xnor U12253 (N_12253,N_11905,N_11853);
nor U12254 (N_12254,N_11615,N_11573);
xor U12255 (N_12255,N_11530,N_11877);
nand U12256 (N_12256,N_11637,N_11980);
or U12257 (N_12257,N_11811,N_11736);
xor U12258 (N_12258,N_11667,N_11561);
nor U12259 (N_12259,N_11938,N_11747);
or U12260 (N_12260,N_11771,N_11706);
nor U12261 (N_12261,N_11510,N_11975);
xor U12262 (N_12262,N_11703,N_11895);
xnor U12263 (N_12263,N_11641,N_11760);
and U12264 (N_12264,N_11640,N_11503);
xnor U12265 (N_12265,N_11572,N_11527);
and U12266 (N_12266,N_11512,N_11632);
xnor U12267 (N_12267,N_11553,N_11867);
and U12268 (N_12268,N_11581,N_11924);
or U12269 (N_12269,N_11831,N_11610);
xnor U12270 (N_12270,N_11869,N_11893);
or U12271 (N_12271,N_11849,N_11666);
or U12272 (N_12272,N_11615,N_11822);
nor U12273 (N_12273,N_11514,N_11529);
and U12274 (N_12274,N_11529,N_11789);
or U12275 (N_12275,N_11869,N_11870);
and U12276 (N_12276,N_11958,N_11998);
and U12277 (N_12277,N_11919,N_11712);
or U12278 (N_12278,N_11868,N_11519);
and U12279 (N_12279,N_11738,N_11923);
nor U12280 (N_12280,N_11773,N_11721);
or U12281 (N_12281,N_11698,N_11836);
xor U12282 (N_12282,N_11866,N_11855);
and U12283 (N_12283,N_11637,N_11533);
xor U12284 (N_12284,N_11709,N_11951);
xnor U12285 (N_12285,N_11879,N_11711);
and U12286 (N_12286,N_11785,N_11880);
nor U12287 (N_12287,N_11949,N_11948);
xnor U12288 (N_12288,N_11666,N_11519);
nand U12289 (N_12289,N_11991,N_11527);
nor U12290 (N_12290,N_11989,N_11618);
or U12291 (N_12291,N_11994,N_11773);
nand U12292 (N_12292,N_11628,N_11788);
xor U12293 (N_12293,N_11880,N_11817);
nand U12294 (N_12294,N_11949,N_11988);
and U12295 (N_12295,N_11728,N_11680);
nand U12296 (N_12296,N_11704,N_11675);
nor U12297 (N_12297,N_11764,N_11767);
nand U12298 (N_12298,N_11602,N_11915);
nand U12299 (N_12299,N_11894,N_11839);
nand U12300 (N_12300,N_11623,N_11805);
nand U12301 (N_12301,N_11824,N_11898);
xor U12302 (N_12302,N_11560,N_11584);
and U12303 (N_12303,N_11940,N_11770);
nand U12304 (N_12304,N_11784,N_11662);
xor U12305 (N_12305,N_11510,N_11645);
xor U12306 (N_12306,N_11664,N_11980);
nor U12307 (N_12307,N_11616,N_11983);
nand U12308 (N_12308,N_11646,N_11763);
nor U12309 (N_12309,N_11823,N_11574);
and U12310 (N_12310,N_11573,N_11570);
nor U12311 (N_12311,N_11610,N_11679);
xnor U12312 (N_12312,N_11719,N_11676);
xnor U12313 (N_12313,N_11681,N_11579);
or U12314 (N_12314,N_11719,N_11650);
xor U12315 (N_12315,N_11780,N_11711);
nand U12316 (N_12316,N_11574,N_11775);
nand U12317 (N_12317,N_11603,N_11996);
nor U12318 (N_12318,N_11782,N_11698);
nor U12319 (N_12319,N_11869,N_11906);
nor U12320 (N_12320,N_11854,N_11582);
and U12321 (N_12321,N_11854,N_11627);
xnor U12322 (N_12322,N_11625,N_11627);
and U12323 (N_12323,N_11828,N_11688);
nand U12324 (N_12324,N_11662,N_11836);
nand U12325 (N_12325,N_11992,N_11789);
xnor U12326 (N_12326,N_11908,N_11511);
nor U12327 (N_12327,N_11514,N_11885);
nand U12328 (N_12328,N_11964,N_11781);
nor U12329 (N_12329,N_11535,N_11525);
nand U12330 (N_12330,N_11758,N_11880);
xor U12331 (N_12331,N_11527,N_11882);
xor U12332 (N_12332,N_11848,N_11835);
xor U12333 (N_12333,N_11903,N_11886);
xnor U12334 (N_12334,N_11748,N_11606);
nor U12335 (N_12335,N_11932,N_11606);
or U12336 (N_12336,N_11716,N_11948);
and U12337 (N_12337,N_11619,N_11798);
xnor U12338 (N_12338,N_11590,N_11940);
and U12339 (N_12339,N_11764,N_11865);
nand U12340 (N_12340,N_11854,N_11703);
nand U12341 (N_12341,N_11769,N_11530);
nor U12342 (N_12342,N_11940,N_11896);
nor U12343 (N_12343,N_11667,N_11747);
nor U12344 (N_12344,N_11577,N_11657);
nand U12345 (N_12345,N_11920,N_11780);
xnor U12346 (N_12346,N_11983,N_11784);
and U12347 (N_12347,N_11810,N_11927);
nand U12348 (N_12348,N_11529,N_11677);
nand U12349 (N_12349,N_11598,N_11732);
or U12350 (N_12350,N_11572,N_11517);
or U12351 (N_12351,N_11597,N_11714);
and U12352 (N_12352,N_11774,N_11948);
xor U12353 (N_12353,N_11607,N_11770);
or U12354 (N_12354,N_11682,N_11718);
or U12355 (N_12355,N_11611,N_11912);
nor U12356 (N_12356,N_11768,N_11603);
nand U12357 (N_12357,N_11516,N_11791);
and U12358 (N_12358,N_11575,N_11657);
nor U12359 (N_12359,N_11712,N_11963);
or U12360 (N_12360,N_11677,N_11688);
and U12361 (N_12361,N_11838,N_11832);
or U12362 (N_12362,N_11871,N_11624);
xor U12363 (N_12363,N_11591,N_11918);
nand U12364 (N_12364,N_11922,N_11558);
and U12365 (N_12365,N_11612,N_11833);
nor U12366 (N_12366,N_11784,N_11991);
xnor U12367 (N_12367,N_11882,N_11847);
and U12368 (N_12368,N_11935,N_11850);
and U12369 (N_12369,N_11855,N_11680);
and U12370 (N_12370,N_11839,N_11508);
or U12371 (N_12371,N_11563,N_11802);
nand U12372 (N_12372,N_11801,N_11601);
nand U12373 (N_12373,N_11924,N_11753);
nand U12374 (N_12374,N_11731,N_11745);
xnor U12375 (N_12375,N_11780,N_11839);
and U12376 (N_12376,N_11712,N_11767);
or U12377 (N_12377,N_11762,N_11940);
nand U12378 (N_12378,N_11748,N_11846);
xnor U12379 (N_12379,N_11817,N_11927);
and U12380 (N_12380,N_11931,N_11762);
and U12381 (N_12381,N_11774,N_11778);
nand U12382 (N_12382,N_11875,N_11977);
xor U12383 (N_12383,N_11716,N_11734);
xor U12384 (N_12384,N_11943,N_11623);
xnor U12385 (N_12385,N_11984,N_11814);
xor U12386 (N_12386,N_11911,N_11870);
and U12387 (N_12387,N_11701,N_11532);
nor U12388 (N_12388,N_11738,N_11932);
and U12389 (N_12389,N_11668,N_11994);
or U12390 (N_12390,N_11621,N_11747);
nor U12391 (N_12391,N_11846,N_11793);
or U12392 (N_12392,N_11624,N_11907);
or U12393 (N_12393,N_11734,N_11807);
nor U12394 (N_12394,N_11714,N_11702);
and U12395 (N_12395,N_11517,N_11957);
nand U12396 (N_12396,N_11888,N_11748);
or U12397 (N_12397,N_11985,N_11995);
and U12398 (N_12398,N_11869,N_11730);
xnor U12399 (N_12399,N_11906,N_11538);
xnor U12400 (N_12400,N_11849,N_11727);
and U12401 (N_12401,N_11551,N_11513);
xnor U12402 (N_12402,N_11624,N_11644);
xor U12403 (N_12403,N_11573,N_11807);
or U12404 (N_12404,N_11559,N_11679);
nor U12405 (N_12405,N_11724,N_11975);
xnor U12406 (N_12406,N_11971,N_11506);
and U12407 (N_12407,N_11739,N_11887);
nand U12408 (N_12408,N_11508,N_11533);
xor U12409 (N_12409,N_11842,N_11872);
or U12410 (N_12410,N_11639,N_11829);
nand U12411 (N_12411,N_11619,N_11564);
nand U12412 (N_12412,N_11981,N_11985);
or U12413 (N_12413,N_11854,N_11642);
nand U12414 (N_12414,N_11727,N_11506);
or U12415 (N_12415,N_11553,N_11908);
nor U12416 (N_12416,N_11680,N_11883);
nand U12417 (N_12417,N_11545,N_11573);
nand U12418 (N_12418,N_11776,N_11821);
xnor U12419 (N_12419,N_11546,N_11846);
xnor U12420 (N_12420,N_11532,N_11739);
nand U12421 (N_12421,N_11883,N_11639);
or U12422 (N_12422,N_11675,N_11913);
or U12423 (N_12423,N_11680,N_11875);
or U12424 (N_12424,N_11687,N_11643);
nand U12425 (N_12425,N_11950,N_11851);
xnor U12426 (N_12426,N_11923,N_11840);
xnor U12427 (N_12427,N_11750,N_11604);
and U12428 (N_12428,N_11613,N_11729);
or U12429 (N_12429,N_11567,N_11681);
nor U12430 (N_12430,N_11674,N_11685);
or U12431 (N_12431,N_11953,N_11752);
nand U12432 (N_12432,N_11809,N_11759);
xnor U12433 (N_12433,N_11694,N_11518);
nand U12434 (N_12434,N_11514,N_11852);
and U12435 (N_12435,N_11870,N_11757);
and U12436 (N_12436,N_11887,N_11807);
nor U12437 (N_12437,N_11589,N_11719);
and U12438 (N_12438,N_11621,N_11786);
or U12439 (N_12439,N_11993,N_11674);
nand U12440 (N_12440,N_11618,N_11822);
xnor U12441 (N_12441,N_11796,N_11849);
or U12442 (N_12442,N_11594,N_11875);
or U12443 (N_12443,N_11730,N_11742);
or U12444 (N_12444,N_11801,N_11665);
nand U12445 (N_12445,N_11810,N_11847);
and U12446 (N_12446,N_11782,N_11733);
and U12447 (N_12447,N_11912,N_11907);
nor U12448 (N_12448,N_11826,N_11541);
and U12449 (N_12449,N_11722,N_11743);
nand U12450 (N_12450,N_11955,N_11944);
or U12451 (N_12451,N_11822,N_11938);
nor U12452 (N_12452,N_11554,N_11740);
xor U12453 (N_12453,N_11661,N_11744);
nand U12454 (N_12454,N_11577,N_11643);
nor U12455 (N_12455,N_11724,N_11808);
or U12456 (N_12456,N_11613,N_11662);
xor U12457 (N_12457,N_11920,N_11809);
nor U12458 (N_12458,N_11773,N_11728);
or U12459 (N_12459,N_11776,N_11865);
nor U12460 (N_12460,N_11591,N_11554);
nand U12461 (N_12461,N_11913,N_11596);
xor U12462 (N_12462,N_11911,N_11537);
and U12463 (N_12463,N_11875,N_11846);
or U12464 (N_12464,N_11857,N_11657);
and U12465 (N_12465,N_11633,N_11553);
and U12466 (N_12466,N_11624,N_11929);
or U12467 (N_12467,N_11738,N_11784);
xor U12468 (N_12468,N_11558,N_11755);
and U12469 (N_12469,N_11692,N_11966);
and U12470 (N_12470,N_11521,N_11714);
or U12471 (N_12471,N_11852,N_11585);
nor U12472 (N_12472,N_11667,N_11607);
or U12473 (N_12473,N_11679,N_11948);
nor U12474 (N_12474,N_11598,N_11942);
nor U12475 (N_12475,N_11585,N_11952);
nor U12476 (N_12476,N_11648,N_11767);
nor U12477 (N_12477,N_11949,N_11536);
and U12478 (N_12478,N_11903,N_11899);
nand U12479 (N_12479,N_11585,N_11815);
nor U12480 (N_12480,N_11599,N_11651);
nor U12481 (N_12481,N_11550,N_11528);
nand U12482 (N_12482,N_11770,N_11661);
or U12483 (N_12483,N_11842,N_11806);
nand U12484 (N_12484,N_11931,N_11714);
nor U12485 (N_12485,N_11666,N_11572);
nor U12486 (N_12486,N_11798,N_11662);
xor U12487 (N_12487,N_11796,N_11690);
nand U12488 (N_12488,N_11560,N_11982);
and U12489 (N_12489,N_11918,N_11913);
xnor U12490 (N_12490,N_11848,N_11760);
and U12491 (N_12491,N_11867,N_11583);
nor U12492 (N_12492,N_11647,N_11852);
and U12493 (N_12493,N_11694,N_11522);
or U12494 (N_12494,N_11859,N_11699);
nand U12495 (N_12495,N_11557,N_11515);
xnor U12496 (N_12496,N_11931,N_11755);
xnor U12497 (N_12497,N_11920,N_11707);
nor U12498 (N_12498,N_11890,N_11820);
and U12499 (N_12499,N_11741,N_11583);
xnor U12500 (N_12500,N_12103,N_12251);
nand U12501 (N_12501,N_12126,N_12423);
nor U12502 (N_12502,N_12190,N_12176);
xor U12503 (N_12503,N_12363,N_12014);
nor U12504 (N_12504,N_12340,N_12288);
or U12505 (N_12505,N_12482,N_12321);
or U12506 (N_12506,N_12112,N_12496);
or U12507 (N_12507,N_12428,N_12267);
nand U12508 (N_12508,N_12419,N_12319);
nor U12509 (N_12509,N_12403,N_12488);
nand U12510 (N_12510,N_12392,N_12148);
nor U12511 (N_12511,N_12384,N_12359);
and U12512 (N_12512,N_12373,N_12468);
xor U12513 (N_12513,N_12351,N_12433);
nor U12514 (N_12514,N_12411,N_12413);
nor U12515 (N_12515,N_12466,N_12007);
and U12516 (N_12516,N_12114,N_12202);
nand U12517 (N_12517,N_12388,N_12162);
nor U12518 (N_12518,N_12188,N_12163);
nand U12519 (N_12519,N_12121,N_12110);
or U12520 (N_12520,N_12342,N_12345);
xnor U12521 (N_12521,N_12352,N_12442);
or U12522 (N_12522,N_12375,N_12414);
nor U12523 (N_12523,N_12144,N_12323);
xor U12524 (N_12524,N_12032,N_12383);
xor U12525 (N_12525,N_12369,N_12212);
and U12526 (N_12526,N_12109,N_12254);
nand U12527 (N_12527,N_12074,N_12377);
and U12528 (N_12528,N_12401,N_12235);
xnor U12529 (N_12529,N_12424,N_12196);
xor U12530 (N_12530,N_12037,N_12257);
nand U12531 (N_12531,N_12417,N_12459);
or U12532 (N_12532,N_12472,N_12490);
nor U12533 (N_12533,N_12206,N_12157);
xnor U12534 (N_12534,N_12056,N_12435);
or U12535 (N_12535,N_12180,N_12462);
nor U12536 (N_12536,N_12437,N_12054);
nor U12537 (N_12537,N_12033,N_12486);
nand U12538 (N_12538,N_12222,N_12491);
xor U12539 (N_12539,N_12397,N_12106);
xnor U12540 (N_12540,N_12193,N_12346);
xnor U12541 (N_12541,N_12438,N_12208);
nand U12542 (N_12542,N_12077,N_12365);
or U12543 (N_12543,N_12060,N_12205);
nand U12544 (N_12544,N_12349,N_12400);
nor U12545 (N_12545,N_12451,N_12426);
or U12546 (N_12546,N_12207,N_12443);
or U12547 (N_12547,N_12116,N_12009);
nor U12548 (N_12548,N_12127,N_12296);
xor U12549 (N_12549,N_12250,N_12356);
nand U12550 (N_12550,N_12256,N_12004);
nand U12551 (N_12551,N_12156,N_12456);
nand U12552 (N_12552,N_12260,N_12024);
or U12553 (N_12553,N_12140,N_12063);
or U12554 (N_12554,N_12043,N_12334);
nor U12555 (N_12555,N_12420,N_12436);
xor U12556 (N_12556,N_12463,N_12255);
nor U12557 (N_12557,N_12195,N_12080);
xnor U12558 (N_12558,N_12330,N_12450);
nand U12559 (N_12559,N_12154,N_12278);
nor U12560 (N_12560,N_12380,N_12171);
or U12561 (N_12561,N_12310,N_12481);
or U12562 (N_12562,N_12046,N_12370);
and U12563 (N_12563,N_12371,N_12470);
xnor U12564 (N_12564,N_12059,N_12072);
nand U12565 (N_12565,N_12192,N_12439);
nand U12566 (N_12566,N_12241,N_12282);
or U12567 (N_12567,N_12252,N_12336);
xnor U12568 (N_12568,N_12013,N_12389);
xnor U12569 (N_12569,N_12368,N_12324);
nor U12570 (N_12570,N_12136,N_12402);
nand U12571 (N_12571,N_12233,N_12001);
nor U12572 (N_12572,N_12284,N_12011);
nand U12573 (N_12573,N_12385,N_12227);
xor U12574 (N_12574,N_12115,N_12429);
and U12575 (N_12575,N_12221,N_12134);
nand U12576 (N_12576,N_12259,N_12404);
nor U12577 (N_12577,N_12418,N_12053);
xnor U12578 (N_12578,N_12215,N_12445);
nand U12579 (N_12579,N_12133,N_12066);
or U12580 (N_12580,N_12091,N_12258);
nand U12581 (N_12581,N_12067,N_12304);
or U12582 (N_12582,N_12326,N_12313);
nor U12583 (N_12583,N_12306,N_12360);
nand U12584 (N_12584,N_12494,N_12308);
nor U12585 (N_12585,N_12331,N_12057);
nor U12586 (N_12586,N_12272,N_12027);
and U12587 (N_12587,N_12294,N_12003);
nand U12588 (N_12588,N_12475,N_12016);
and U12589 (N_12589,N_12399,N_12249);
and U12590 (N_12590,N_12076,N_12381);
and U12591 (N_12591,N_12454,N_12303);
and U12592 (N_12592,N_12045,N_12453);
xor U12593 (N_12593,N_12130,N_12030);
xnor U12594 (N_12594,N_12292,N_12293);
xnor U12595 (N_12595,N_12335,N_12409);
xor U12596 (N_12596,N_12253,N_12123);
and U12597 (N_12597,N_12169,N_12317);
nor U12598 (N_12598,N_12231,N_12405);
or U12599 (N_12599,N_12149,N_12350);
xor U12600 (N_12600,N_12230,N_12170);
and U12601 (N_12601,N_12058,N_12497);
xor U12602 (N_12602,N_12085,N_12337);
or U12603 (N_12603,N_12055,N_12108);
or U12604 (N_12604,N_12020,N_12320);
xor U12605 (N_12605,N_12262,N_12042);
xor U12606 (N_12606,N_12487,N_12469);
nand U12607 (N_12607,N_12301,N_12097);
or U12608 (N_12608,N_12309,N_12187);
xnor U12609 (N_12609,N_12299,N_12312);
nand U12610 (N_12610,N_12464,N_12295);
or U12611 (N_12611,N_12019,N_12247);
nand U12612 (N_12612,N_12044,N_12070);
xnor U12613 (N_12613,N_12446,N_12021);
nand U12614 (N_12614,N_12285,N_12372);
or U12615 (N_12615,N_12086,N_12261);
nand U12616 (N_12616,N_12224,N_12201);
and U12617 (N_12617,N_12493,N_12158);
xnor U12618 (N_12618,N_12266,N_12465);
or U12619 (N_12619,N_12364,N_12090);
and U12620 (N_12620,N_12089,N_12248);
or U12621 (N_12621,N_12047,N_12049);
nand U12622 (N_12622,N_12499,N_12209);
nand U12623 (N_12623,N_12084,N_12052);
nor U12624 (N_12624,N_12146,N_12175);
xnor U12625 (N_12625,N_12094,N_12167);
and U12626 (N_12626,N_12025,N_12361);
or U12627 (N_12627,N_12305,N_12172);
nand U12628 (N_12628,N_12141,N_12245);
nor U12629 (N_12629,N_12028,N_12006);
nor U12630 (N_12630,N_12069,N_12166);
xnor U12631 (N_12631,N_12311,N_12159);
nor U12632 (N_12632,N_12122,N_12268);
xor U12633 (N_12633,N_12398,N_12008);
nand U12634 (N_12634,N_12300,N_12150);
xnor U12635 (N_12635,N_12183,N_12449);
or U12636 (N_12636,N_12291,N_12325);
nand U12637 (N_12637,N_12099,N_12165);
nor U12638 (N_12638,N_12218,N_12131);
xnor U12639 (N_12639,N_12104,N_12434);
and U12640 (N_12640,N_12161,N_12480);
xor U12641 (N_12641,N_12395,N_12274);
and U12642 (N_12642,N_12410,N_12279);
nor U12643 (N_12643,N_12137,N_12182);
nand U12644 (N_12644,N_12269,N_12421);
nor U12645 (N_12645,N_12113,N_12005);
xnor U12646 (N_12646,N_12098,N_12366);
nand U12647 (N_12647,N_12302,N_12474);
nor U12648 (N_12648,N_12228,N_12217);
nor U12649 (N_12649,N_12031,N_12026);
xor U12650 (N_12650,N_12328,N_12354);
nand U12651 (N_12651,N_12065,N_12455);
nand U12652 (N_12652,N_12068,N_12275);
nor U12653 (N_12653,N_12064,N_12181);
nor U12654 (N_12654,N_12062,N_12197);
or U12655 (N_12655,N_12393,N_12338);
xor U12656 (N_12656,N_12087,N_12002);
xnor U12657 (N_12657,N_12096,N_12362);
and U12658 (N_12658,N_12347,N_12479);
nand U12659 (N_12659,N_12194,N_12022);
or U12660 (N_12660,N_12394,N_12041);
nand U12661 (N_12661,N_12242,N_12270);
nand U12662 (N_12662,N_12035,N_12498);
nor U12663 (N_12663,N_12151,N_12378);
or U12664 (N_12664,N_12477,N_12236);
nand U12665 (N_12665,N_12117,N_12343);
nor U12666 (N_12666,N_12484,N_12382);
nand U12667 (N_12667,N_12101,N_12124);
or U12668 (N_12668,N_12358,N_12379);
and U12669 (N_12669,N_12322,N_12339);
nor U12670 (N_12670,N_12179,N_12125);
nand U12671 (N_12671,N_12092,N_12286);
xnor U12672 (N_12672,N_12135,N_12489);
and U12673 (N_12673,N_12100,N_12289);
nand U12674 (N_12674,N_12000,N_12229);
nand U12675 (N_12675,N_12147,N_12128);
or U12676 (N_12676,N_12204,N_12203);
or U12677 (N_12677,N_12102,N_12039);
or U12678 (N_12678,N_12376,N_12226);
nand U12679 (N_12679,N_12374,N_12238);
nor U12680 (N_12680,N_12287,N_12199);
and U12681 (N_12681,N_12083,N_12142);
xor U12682 (N_12682,N_12223,N_12214);
nor U12683 (N_12683,N_12120,N_12073);
nand U12684 (N_12684,N_12447,N_12473);
nor U12685 (N_12685,N_12168,N_12457);
xor U12686 (N_12686,N_12119,N_12132);
nand U12687 (N_12687,N_12440,N_12093);
nand U12688 (N_12688,N_12071,N_12153);
and U12689 (N_12689,N_12271,N_12422);
xnor U12690 (N_12690,N_12081,N_12471);
or U12691 (N_12691,N_12152,N_12239);
xor U12692 (N_12692,N_12390,N_12263);
nand U12693 (N_12693,N_12408,N_12186);
nor U12694 (N_12694,N_12430,N_12225);
nand U12695 (N_12695,N_12348,N_12425);
or U12696 (N_12696,N_12210,N_12234);
nor U12697 (N_12697,N_12315,N_12277);
nand U12698 (N_12698,N_12333,N_12177);
nor U12699 (N_12699,N_12452,N_12307);
or U12700 (N_12700,N_12111,N_12495);
nand U12701 (N_12701,N_12211,N_12483);
and U12702 (N_12702,N_12145,N_12220);
nand U12703 (N_12703,N_12174,N_12015);
or U12704 (N_12704,N_12298,N_12184);
xor U12705 (N_12705,N_12018,N_12243);
nand U12706 (N_12706,N_12478,N_12219);
or U12707 (N_12707,N_12427,N_12391);
xor U12708 (N_12708,N_12432,N_12178);
xnor U12709 (N_12709,N_12164,N_12283);
or U12710 (N_12710,N_12412,N_12476);
nand U12711 (N_12711,N_12281,N_12276);
and U12712 (N_12712,N_12441,N_12460);
xor U12713 (N_12713,N_12318,N_12290);
or U12714 (N_12714,N_12118,N_12416);
xnor U12715 (N_12715,N_12316,N_12189);
or U12716 (N_12716,N_12095,N_12012);
or U12717 (N_12717,N_12327,N_12448);
and U12718 (N_12718,N_12036,N_12341);
nor U12719 (N_12719,N_12444,N_12040);
xnor U12720 (N_12720,N_12264,N_12431);
and U12721 (N_12721,N_12160,N_12023);
nand U12722 (N_12722,N_12143,N_12017);
or U12723 (N_12723,N_12244,N_12467);
or U12724 (N_12724,N_12010,N_12265);
and U12725 (N_12725,N_12237,N_12406);
and U12726 (N_12726,N_12485,N_12216);
or U12727 (N_12727,N_12332,N_12139);
xor U12728 (N_12728,N_12173,N_12155);
xnor U12729 (N_12729,N_12082,N_12051);
xnor U12730 (N_12730,N_12387,N_12297);
nor U12731 (N_12731,N_12407,N_12200);
xor U12732 (N_12732,N_12329,N_12240);
nand U12733 (N_12733,N_12355,N_12492);
nor U12734 (N_12734,N_12050,N_12034);
and U12735 (N_12735,N_12314,N_12048);
and U12736 (N_12736,N_12185,N_12088);
xnor U12737 (N_12737,N_12357,N_12280);
nand U12738 (N_12738,N_12075,N_12198);
xor U12739 (N_12739,N_12038,N_12191);
and U12740 (N_12740,N_12246,N_12344);
or U12741 (N_12741,N_12461,N_12386);
xnor U12742 (N_12742,N_12273,N_12107);
and U12743 (N_12743,N_12415,N_12353);
and U12744 (N_12744,N_12061,N_12078);
nor U12745 (N_12745,N_12396,N_12129);
and U12746 (N_12746,N_12458,N_12029);
nand U12747 (N_12747,N_12079,N_12213);
nor U12748 (N_12748,N_12367,N_12105);
xor U12749 (N_12749,N_12138,N_12232);
nor U12750 (N_12750,N_12033,N_12359);
nand U12751 (N_12751,N_12381,N_12285);
or U12752 (N_12752,N_12297,N_12079);
or U12753 (N_12753,N_12298,N_12253);
or U12754 (N_12754,N_12153,N_12381);
and U12755 (N_12755,N_12009,N_12037);
nand U12756 (N_12756,N_12273,N_12099);
nand U12757 (N_12757,N_12485,N_12402);
and U12758 (N_12758,N_12143,N_12316);
and U12759 (N_12759,N_12373,N_12275);
and U12760 (N_12760,N_12410,N_12130);
nand U12761 (N_12761,N_12288,N_12116);
or U12762 (N_12762,N_12190,N_12075);
or U12763 (N_12763,N_12273,N_12218);
xnor U12764 (N_12764,N_12099,N_12299);
xor U12765 (N_12765,N_12320,N_12019);
xor U12766 (N_12766,N_12320,N_12073);
nand U12767 (N_12767,N_12107,N_12219);
or U12768 (N_12768,N_12218,N_12201);
and U12769 (N_12769,N_12014,N_12325);
and U12770 (N_12770,N_12385,N_12132);
nor U12771 (N_12771,N_12015,N_12474);
xor U12772 (N_12772,N_12374,N_12259);
nor U12773 (N_12773,N_12144,N_12492);
or U12774 (N_12774,N_12282,N_12490);
xor U12775 (N_12775,N_12245,N_12372);
nor U12776 (N_12776,N_12163,N_12489);
or U12777 (N_12777,N_12414,N_12480);
and U12778 (N_12778,N_12265,N_12334);
or U12779 (N_12779,N_12237,N_12185);
or U12780 (N_12780,N_12272,N_12002);
and U12781 (N_12781,N_12198,N_12461);
and U12782 (N_12782,N_12493,N_12293);
or U12783 (N_12783,N_12328,N_12405);
nand U12784 (N_12784,N_12428,N_12003);
nand U12785 (N_12785,N_12452,N_12201);
nor U12786 (N_12786,N_12264,N_12212);
or U12787 (N_12787,N_12085,N_12453);
or U12788 (N_12788,N_12357,N_12426);
or U12789 (N_12789,N_12099,N_12120);
or U12790 (N_12790,N_12452,N_12433);
nand U12791 (N_12791,N_12107,N_12062);
and U12792 (N_12792,N_12103,N_12234);
nand U12793 (N_12793,N_12294,N_12439);
and U12794 (N_12794,N_12349,N_12415);
nor U12795 (N_12795,N_12460,N_12358);
nand U12796 (N_12796,N_12077,N_12493);
nor U12797 (N_12797,N_12220,N_12225);
nor U12798 (N_12798,N_12266,N_12117);
and U12799 (N_12799,N_12379,N_12224);
nand U12800 (N_12800,N_12204,N_12085);
nand U12801 (N_12801,N_12404,N_12407);
xor U12802 (N_12802,N_12382,N_12372);
nor U12803 (N_12803,N_12245,N_12403);
nand U12804 (N_12804,N_12018,N_12267);
nor U12805 (N_12805,N_12440,N_12475);
xor U12806 (N_12806,N_12356,N_12434);
nand U12807 (N_12807,N_12424,N_12278);
and U12808 (N_12808,N_12380,N_12423);
nand U12809 (N_12809,N_12451,N_12372);
xnor U12810 (N_12810,N_12042,N_12085);
nor U12811 (N_12811,N_12443,N_12246);
nand U12812 (N_12812,N_12342,N_12378);
and U12813 (N_12813,N_12417,N_12060);
nor U12814 (N_12814,N_12283,N_12145);
and U12815 (N_12815,N_12046,N_12222);
nor U12816 (N_12816,N_12175,N_12192);
nor U12817 (N_12817,N_12340,N_12261);
nor U12818 (N_12818,N_12068,N_12197);
and U12819 (N_12819,N_12443,N_12272);
nor U12820 (N_12820,N_12018,N_12121);
nand U12821 (N_12821,N_12253,N_12480);
or U12822 (N_12822,N_12313,N_12124);
xor U12823 (N_12823,N_12039,N_12422);
xnor U12824 (N_12824,N_12190,N_12228);
and U12825 (N_12825,N_12109,N_12145);
xnor U12826 (N_12826,N_12387,N_12330);
nor U12827 (N_12827,N_12298,N_12388);
nor U12828 (N_12828,N_12315,N_12059);
or U12829 (N_12829,N_12129,N_12419);
or U12830 (N_12830,N_12232,N_12022);
or U12831 (N_12831,N_12227,N_12139);
xnor U12832 (N_12832,N_12432,N_12430);
or U12833 (N_12833,N_12407,N_12347);
nand U12834 (N_12834,N_12206,N_12306);
nor U12835 (N_12835,N_12134,N_12469);
and U12836 (N_12836,N_12138,N_12292);
or U12837 (N_12837,N_12350,N_12093);
nor U12838 (N_12838,N_12231,N_12309);
xnor U12839 (N_12839,N_12262,N_12271);
nand U12840 (N_12840,N_12144,N_12052);
or U12841 (N_12841,N_12076,N_12324);
and U12842 (N_12842,N_12272,N_12282);
xor U12843 (N_12843,N_12252,N_12017);
or U12844 (N_12844,N_12182,N_12177);
nor U12845 (N_12845,N_12307,N_12468);
nor U12846 (N_12846,N_12155,N_12145);
nand U12847 (N_12847,N_12350,N_12212);
or U12848 (N_12848,N_12067,N_12287);
xnor U12849 (N_12849,N_12266,N_12039);
nor U12850 (N_12850,N_12125,N_12312);
xor U12851 (N_12851,N_12146,N_12137);
or U12852 (N_12852,N_12139,N_12274);
and U12853 (N_12853,N_12118,N_12114);
nor U12854 (N_12854,N_12316,N_12252);
nor U12855 (N_12855,N_12214,N_12160);
and U12856 (N_12856,N_12055,N_12338);
and U12857 (N_12857,N_12007,N_12144);
or U12858 (N_12858,N_12088,N_12004);
xnor U12859 (N_12859,N_12179,N_12022);
nand U12860 (N_12860,N_12225,N_12461);
nor U12861 (N_12861,N_12262,N_12048);
or U12862 (N_12862,N_12432,N_12269);
xnor U12863 (N_12863,N_12254,N_12433);
nor U12864 (N_12864,N_12220,N_12387);
nand U12865 (N_12865,N_12021,N_12119);
and U12866 (N_12866,N_12294,N_12344);
xnor U12867 (N_12867,N_12411,N_12051);
and U12868 (N_12868,N_12235,N_12064);
nand U12869 (N_12869,N_12191,N_12041);
nor U12870 (N_12870,N_12215,N_12489);
nor U12871 (N_12871,N_12416,N_12290);
nand U12872 (N_12872,N_12084,N_12470);
nand U12873 (N_12873,N_12332,N_12233);
or U12874 (N_12874,N_12479,N_12269);
or U12875 (N_12875,N_12167,N_12244);
and U12876 (N_12876,N_12107,N_12036);
xnor U12877 (N_12877,N_12400,N_12407);
nand U12878 (N_12878,N_12460,N_12171);
nor U12879 (N_12879,N_12418,N_12097);
and U12880 (N_12880,N_12091,N_12351);
and U12881 (N_12881,N_12274,N_12468);
xnor U12882 (N_12882,N_12327,N_12467);
or U12883 (N_12883,N_12073,N_12448);
or U12884 (N_12884,N_12233,N_12147);
and U12885 (N_12885,N_12485,N_12225);
nor U12886 (N_12886,N_12190,N_12398);
nor U12887 (N_12887,N_12378,N_12217);
and U12888 (N_12888,N_12435,N_12436);
nand U12889 (N_12889,N_12364,N_12300);
nor U12890 (N_12890,N_12348,N_12322);
nand U12891 (N_12891,N_12238,N_12126);
nand U12892 (N_12892,N_12375,N_12311);
xor U12893 (N_12893,N_12424,N_12282);
nor U12894 (N_12894,N_12472,N_12328);
nand U12895 (N_12895,N_12142,N_12120);
nand U12896 (N_12896,N_12421,N_12175);
and U12897 (N_12897,N_12011,N_12327);
or U12898 (N_12898,N_12363,N_12217);
and U12899 (N_12899,N_12138,N_12415);
xor U12900 (N_12900,N_12425,N_12300);
nor U12901 (N_12901,N_12419,N_12402);
xor U12902 (N_12902,N_12246,N_12469);
xor U12903 (N_12903,N_12486,N_12131);
xor U12904 (N_12904,N_12037,N_12493);
nor U12905 (N_12905,N_12195,N_12294);
or U12906 (N_12906,N_12111,N_12460);
and U12907 (N_12907,N_12184,N_12107);
or U12908 (N_12908,N_12009,N_12180);
nand U12909 (N_12909,N_12358,N_12071);
nor U12910 (N_12910,N_12066,N_12429);
and U12911 (N_12911,N_12365,N_12475);
xor U12912 (N_12912,N_12061,N_12348);
or U12913 (N_12913,N_12313,N_12134);
and U12914 (N_12914,N_12337,N_12176);
xnor U12915 (N_12915,N_12380,N_12491);
or U12916 (N_12916,N_12452,N_12464);
nor U12917 (N_12917,N_12064,N_12396);
or U12918 (N_12918,N_12363,N_12366);
and U12919 (N_12919,N_12257,N_12407);
or U12920 (N_12920,N_12265,N_12287);
xor U12921 (N_12921,N_12088,N_12273);
nand U12922 (N_12922,N_12045,N_12460);
xnor U12923 (N_12923,N_12478,N_12119);
and U12924 (N_12924,N_12175,N_12167);
nand U12925 (N_12925,N_12064,N_12186);
or U12926 (N_12926,N_12338,N_12196);
xnor U12927 (N_12927,N_12008,N_12105);
nand U12928 (N_12928,N_12262,N_12498);
and U12929 (N_12929,N_12325,N_12210);
xor U12930 (N_12930,N_12453,N_12171);
nor U12931 (N_12931,N_12189,N_12050);
or U12932 (N_12932,N_12043,N_12425);
or U12933 (N_12933,N_12300,N_12096);
xor U12934 (N_12934,N_12292,N_12196);
xor U12935 (N_12935,N_12174,N_12312);
nor U12936 (N_12936,N_12304,N_12277);
nor U12937 (N_12937,N_12222,N_12442);
and U12938 (N_12938,N_12226,N_12034);
nand U12939 (N_12939,N_12377,N_12335);
or U12940 (N_12940,N_12130,N_12033);
nor U12941 (N_12941,N_12485,N_12181);
nand U12942 (N_12942,N_12486,N_12199);
nand U12943 (N_12943,N_12348,N_12125);
nand U12944 (N_12944,N_12260,N_12119);
and U12945 (N_12945,N_12345,N_12197);
nand U12946 (N_12946,N_12479,N_12445);
or U12947 (N_12947,N_12283,N_12044);
or U12948 (N_12948,N_12072,N_12489);
nor U12949 (N_12949,N_12296,N_12288);
nor U12950 (N_12950,N_12394,N_12093);
and U12951 (N_12951,N_12216,N_12002);
nand U12952 (N_12952,N_12392,N_12340);
xor U12953 (N_12953,N_12235,N_12157);
xor U12954 (N_12954,N_12285,N_12493);
xnor U12955 (N_12955,N_12161,N_12387);
or U12956 (N_12956,N_12394,N_12331);
nand U12957 (N_12957,N_12215,N_12471);
nor U12958 (N_12958,N_12440,N_12128);
xnor U12959 (N_12959,N_12329,N_12113);
xor U12960 (N_12960,N_12182,N_12144);
or U12961 (N_12961,N_12156,N_12343);
nand U12962 (N_12962,N_12066,N_12382);
and U12963 (N_12963,N_12110,N_12307);
or U12964 (N_12964,N_12073,N_12304);
or U12965 (N_12965,N_12414,N_12263);
xor U12966 (N_12966,N_12003,N_12420);
nor U12967 (N_12967,N_12272,N_12053);
and U12968 (N_12968,N_12132,N_12210);
and U12969 (N_12969,N_12040,N_12197);
or U12970 (N_12970,N_12239,N_12286);
nand U12971 (N_12971,N_12158,N_12052);
nor U12972 (N_12972,N_12171,N_12401);
and U12973 (N_12973,N_12223,N_12276);
nand U12974 (N_12974,N_12106,N_12080);
nand U12975 (N_12975,N_12075,N_12068);
nand U12976 (N_12976,N_12176,N_12076);
and U12977 (N_12977,N_12372,N_12237);
nor U12978 (N_12978,N_12037,N_12237);
or U12979 (N_12979,N_12473,N_12030);
nand U12980 (N_12980,N_12438,N_12454);
and U12981 (N_12981,N_12266,N_12350);
and U12982 (N_12982,N_12371,N_12261);
nand U12983 (N_12983,N_12189,N_12497);
nor U12984 (N_12984,N_12247,N_12425);
nand U12985 (N_12985,N_12040,N_12254);
and U12986 (N_12986,N_12131,N_12226);
xor U12987 (N_12987,N_12063,N_12036);
and U12988 (N_12988,N_12274,N_12173);
nand U12989 (N_12989,N_12031,N_12081);
or U12990 (N_12990,N_12451,N_12202);
nand U12991 (N_12991,N_12039,N_12108);
and U12992 (N_12992,N_12020,N_12431);
nand U12993 (N_12993,N_12310,N_12316);
xor U12994 (N_12994,N_12002,N_12388);
and U12995 (N_12995,N_12404,N_12399);
nor U12996 (N_12996,N_12443,N_12059);
xor U12997 (N_12997,N_12234,N_12224);
xor U12998 (N_12998,N_12057,N_12241);
nand U12999 (N_12999,N_12284,N_12319);
or U13000 (N_13000,N_12808,N_12768);
nand U13001 (N_13001,N_12599,N_12774);
or U13002 (N_13002,N_12623,N_12828);
nand U13003 (N_13003,N_12872,N_12817);
nand U13004 (N_13004,N_12593,N_12570);
and U13005 (N_13005,N_12773,N_12647);
and U13006 (N_13006,N_12691,N_12910);
nand U13007 (N_13007,N_12631,N_12884);
nor U13008 (N_13008,N_12710,N_12543);
xor U13009 (N_13009,N_12661,N_12513);
xnor U13010 (N_13010,N_12722,N_12795);
nand U13011 (N_13011,N_12757,N_12527);
and U13012 (N_13012,N_12897,N_12824);
or U13013 (N_13013,N_12696,N_12715);
nor U13014 (N_13014,N_12585,N_12930);
xor U13015 (N_13015,N_12921,N_12770);
and U13016 (N_13016,N_12815,N_12615);
nor U13017 (N_13017,N_12791,N_12765);
nand U13018 (N_13018,N_12880,N_12723);
xnor U13019 (N_13019,N_12727,N_12990);
nand U13020 (N_13020,N_12767,N_12782);
and U13021 (N_13021,N_12684,N_12551);
nand U13022 (N_13022,N_12987,N_12852);
or U13023 (N_13023,N_12946,N_12894);
xor U13024 (N_13024,N_12816,N_12514);
nand U13025 (N_13025,N_12931,N_12706);
nand U13026 (N_13026,N_12885,N_12625);
xnor U13027 (N_13027,N_12827,N_12771);
nor U13028 (N_13028,N_12978,N_12539);
nand U13029 (N_13029,N_12609,N_12976);
xor U13030 (N_13030,N_12833,N_12903);
nor U13031 (N_13031,N_12592,N_12502);
xnor U13032 (N_13032,N_12580,N_12944);
or U13033 (N_13033,N_12656,N_12755);
and U13034 (N_13034,N_12563,N_12558);
nand U13035 (N_13035,N_12888,N_12938);
nor U13036 (N_13036,N_12835,N_12636);
and U13037 (N_13037,N_12581,N_12855);
or U13038 (N_13038,N_12909,N_12531);
and U13039 (N_13039,N_12967,N_12734);
or U13040 (N_13040,N_12686,N_12947);
nor U13041 (N_13041,N_12951,N_12803);
or U13042 (N_13042,N_12801,N_12783);
or U13043 (N_13043,N_12877,N_12793);
nand U13044 (N_13044,N_12736,N_12574);
xnor U13045 (N_13045,N_12640,N_12674);
xor U13046 (N_13046,N_12657,N_12648);
nor U13047 (N_13047,N_12975,N_12848);
nand U13048 (N_13048,N_12557,N_12898);
nand U13049 (N_13049,N_12540,N_12961);
xor U13050 (N_13050,N_12566,N_12890);
and U13051 (N_13051,N_12954,N_12718);
nand U13052 (N_13052,N_12671,N_12673);
nor U13053 (N_13053,N_12821,N_12915);
nand U13054 (N_13054,N_12555,N_12911);
or U13055 (N_13055,N_12918,N_12842);
xnor U13056 (N_13056,N_12567,N_12959);
or U13057 (N_13057,N_12683,N_12814);
nor U13058 (N_13058,N_12829,N_12507);
or U13059 (N_13059,N_12981,N_12618);
xor U13060 (N_13060,N_12526,N_12854);
xnor U13061 (N_13061,N_12995,N_12998);
and U13062 (N_13062,N_12638,N_12874);
or U13063 (N_13063,N_12548,N_12602);
and U13064 (N_13064,N_12650,N_12730);
or U13065 (N_13065,N_12889,N_12545);
nor U13066 (N_13066,N_12639,N_12660);
nor U13067 (N_13067,N_12780,N_12744);
or U13068 (N_13068,N_12572,N_12505);
or U13069 (N_13069,N_12632,N_12860);
xnor U13070 (N_13070,N_12935,N_12969);
or U13071 (N_13071,N_12996,N_12643);
nand U13072 (N_13072,N_12750,N_12784);
xor U13073 (N_13073,N_12823,N_12738);
and U13074 (N_13074,N_12937,N_12832);
nand U13075 (N_13075,N_12948,N_12893);
nor U13076 (N_13076,N_12984,N_12776);
or U13077 (N_13077,N_12943,N_12772);
xnor U13078 (N_13078,N_12622,N_12510);
or U13079 (N_13079,N_12582,N_12693);
xor U13080 (N_13080,N_12861,N_12846);
or U13081 (N_13081,N_12501,N_12752);
nand U13082 (N_13082,N_12927,N_12807);
xnor U13083 (N_13083,N_12663,N_12899);
nand U13084 (N_13084,N_12611,N_12754);
nand U13085 (N_13085,N_12999,N_12741);
nand U13086 (N_13086,N_12716,N_12810);
and U13087 (N_13087,N_12957,N_12595);
and U13088 (N_13088,N_12541,N_12766);
or U13089 (N_13089,N_12552,N_12806);
nor U13090 (N_13090,N_12979,N_12834);
or U13091 (N_13091,N_12728,N_12634);
xnor U13092 (N_13092,N_12924,N_12908);
or U13093 (N_13093,N_12594,N_12952);
nor U13094 (N_13094,N_12778,N_12530);
and U13095 (N_13095,N_12617,N_12624);
nand U13096 (N_13096,N_12579,N_12613);
xor U13097 (N_13097,N_12642,N_12554);
and U13098 (N_13098,N_12515,N_12649);
and U13099 (N_13099,N_12865,N_12840);
nor U13100 (N_13100,N_12608,N_12584);
or U13101 (N_13101,N_12902,N_12553);
nor U13102 (N_13102,N_12779,N_12644);
nand U13103 (N_13103,N_12533,N_12983);
and U13104 (N_13104,N_12794,N_12620);
nand U13105 (N_13105,N_12503,N_12863);
or U13106 (N_13106,N_12812,N_12839);
or U13107 (N_13107,N_12711,N_12912);
or U13108 (N_13108,N_12532,N_12702);
xor U13109 (N_13109,N_12818,N_12601);
nand U13110 (N_13110,N_12883,N_12790);
nor U13111 (N_13111,N_12578,N_12900);
and U13112 (N_13112,N_12964,N_12717);
xnor U13113 (N_13113,N_12798,N_12621);
or U13114 (N_13114,N_12659,N_12701);
xnor U13115 (N_13115,N_12973,N_12788);
and U13116 (N_13116,N_12968,N_12871);
xor U13117 (N_13117,N_12529,N_12887);
nor U13118 (N_13118,N_12596,N_12628);
and U13119 (N_13119,N_12746,N_12799);
or U13120 (N_13120,N_12742,N_12989);
xor U13121 (N_13121,N_12645,N_12785);
nor U13122 (N_13122,N_12837,N_12565);
or U13123 (N_13123,N_12583,N_12637);
nor U13124 (N_13124,N_12925,N_12714);
and U13125 (N_13125,N_12820,N_12651);
nor U13126 (N_13126,N_12690,N_12712);
or U13127 (N_13127,N_12550,N_12993);
and U13128 (N_13128,N_12523,N_12819);
nor U13129 (N_13129,N_12775,N_12685);
nor U13130 (N_13130,N_12980,N_12928);
nor U13131 (N_13131,N_12777,N_12886);
nor U13132 (N_13132,N_12901,N_12597);
and U13133 (N_13133,N_12822,N_12635);
nor U13134 (N_13134,N_12670,N_12627);
and U13135 (N_13135,N_12534,N_12988);
or U13136 (N_13136,N_12956,N_12525);
or U13137 (N_13137,N_12977,N_12753);
and U13138 (N_13138,N_12985,N_12862);
or U13139 (N_13139,N_12869,N_12849);
nor U13140 (N_13140,N_12564,N_12678);
nand U13141 (N_13141,N_12971,N_12986);
and U13142 (N_13142,N_12626,N_12939);
nand U13143 (N_13143,N_12949,N_12926);
and U13144 (N_13144,N_12731,N_12739);
xor U13145 (N_13145,N_12936,N_12546);
nand U13146 (N_13146,N_12518,N_12845);
or U13147 (N_13147,N_12708,N_12720);
nor U13148 (N_13148,N_12809,N_12607);
and U13149 (N_13149,N_12729,N_12748);
and U13150 (N_13150,N_12689,N_12920);
xnor U13151 (N_13151,N_12573,N_12825);
nand U13152 (N_13152,N_12904,N_12916);
nand U13153 (N_13153,N_12917,N_12687);
or U13154 (N_13154,N_12747,N_12856);
or U13155 (N_13155,N_12914,N_12826);
xnor U13156 (N_13156,N_12761,N_12709);
and U13157 (N_13157,N_12652,N_12516);
or U13158 (N_13158,N_12569,N_12830);
and U13159 (N_13159,N_12907,N_12668);
and U13160 (N_13160,N_12796,N_12789);
nand U13161 (N_13161,N_12600,N_12679);
and U13162 (N_13162,N_12974,N_12740);
nand U13163 (N_13163,N_12521,N_12875);
and U13164 (N_13164,N_12882,N_12700);
xor U13165 (N_13165,N_12751,N_12932);
nand U13166 (N_13166,N_12994,N_12726);
xnor U13167 (N_13167,N_12876,N_12559);
nand U13168 (N_13168,N_12655,N_12844);
nor U13169 (N_13169,N_12509,N_12966);
or U13170 (N_13170,N_12811,N_12965);
nor U13171 (N_13171,N_12633,N_12658);
and U13172 (N_13172,N_12853,N_12695);
nor U13173 (N_13173,N_12517,N_12511);
xnor U13174 (N_13174,N_12838,N_12941);
nand U13175 (N_13175,N_12610,N_12732);
nor U13176 (N_13176,N_12571,N_12508);
nor U13177 (N_13177,N_12836,N_12891);
nand U13178 (N_13178,N_12542,N_12577);
or U13179 (N_13179,N_12547,N_12504);
xor U13180 (N_13180,N_12704,N_12619);
nor U13181 (N_13181,N_12867,N_12735);
or U13182 (N_13182,N_12588,N_12682);
and U13183 (N_13183,N_12614,N_12896);
nand U13184 (N_13184,N_12576,N_12970);
and U13185 (N_13185,N_12864,N_12758);
nor U13186 (N_13186,N_12676,N_12528);
nand U13187 (N_13187,N_12512,N_12688);
or U13188 (N_13188,N_12699,N_12698);
nor U13189 (N_13189,N_12950,N_12879);
nand U13190 (N_13190,N_12972,N_12629);
and U13191 (N_13191,N_12707,N_12675);
nor U13192 (N_13192,N_12598,N_12737);
nor U13193 (N_13193,N_12713,N_12681);
or U13194 (N_13194,N_12866,N_12662);
and U13195 (N_13195,N_12560,N_12725);
nand U13196 (N_13196,N_12802,N_12549);
nand U13197 (N_13197,N_12537,N_12850);
nand U13198 (N_13198,N_12697,N_12705);
xor U13199 (N_13199,N_12743,N_12962);
xnor U13200 (N_13200,N_12942,N_12556);
xor U13201 (N_13201,N_12940,N_12666);
xor U13202 (N_13202,N_12847,N_12945);
nor U13203 (N_13203,N_12653,N_12519);
or U13204 (N_13204,N_12544,N_12881);
and U13205 (N_13205,N_12760,N_12960);
or U13206 (N_13206,N_12524,N_12604);
nand U13207 (N_13207,N_12669,N_12538);
nand U13208 (N_13208,N_12756,N_12786);
nand U13209 (N_13209,N_12859,N_12641);
nand U13210 (N_13210,N_12568,N_12745);
nand U13211 (N_13211,N_12992,N_12800);
xnor U13212 (N_13212,N_12805,N_12672);
nand U13213 (N_13213,N_12953,N_12787);
nand U13214 (N_13214,N_12762,N_12535);
or U13215 (N_13215,N_12763,N_12603);
nand U13216 (N_13216,N_12933,N_12851);
and U13217 (N_13217,N_12667,N_12664);
and U13218 (N_13218,N_12878,N_12575);
and U13219 (N_13219,N_12520,N_12922);
nand U13220 (N_13220,N_12843,N_12958);
nor U13221 (N_13221,N_12955,N_12665);
or U13222 (N_13222,N_12982,N_12589);
or U13223 (N_13223,N_12895,N_12913);
nor U13224 (N_13224,N_12906,N_12500);
and U13225 (N_13225,N_12605,N_12749);
nor U13226 (N_13226,N_12590,N_12646);
nand U13227 (N_13227,N_12692,N_12719);
or U13228 (N_13228,N_12870,N_12868);
xor U13229 (N_13229,N_12759,N_12841);
xnor U13230 (N_13230,N_12586,N_12929);
nand U13231 (N_13231,N_12606,N_12587);
or U13232 (N_13232,N_12873,N_12506);
and U13233 (N_13233,N_12733,N_12764);
nand U13234 (N_13234,N_12991,N_12703);
and U13235 (N_13235,N_12769,N_12677);
nand U13236 (N_13236,N_12561,N_12905);
or U13237 (N_13237,N_12654,N_12858);
nor U13238 (N_13238,N_12797,N_12792);
and U13239 (N_13239,N_12630,N_12694);
nand U13240 (N_13240,N_12857,N_12781);
nand U13241 (N_13241,N_12724,N_12892);
or U13242 (N_13242,N_12919,N_12591);
nor U13243 (N_13243,N_12562,N_12831);
or U13244 (N_13244,N_12813,N_12616);
nor U13245 (N_13245,N_12536,N_12923);
or U13246 (N_13246,N_12522,N_12680);
and U13247 (N_13247,N_12721,N_12612);
nor U13248 (N_13248,N_12997,N_12934);
or U13249 (N_13249,N_12963,N_12804);
xor U13250 (N_13250,N_12783,N_12764);
or U13251 (N_13251,N_12783,N_12522);
nor U13252 (N_13252,N_12733,N_12870);
nand U13253 (N_13253,N_12549,N_12670);
nand U13254 (N_13254,N_12708,N_12527);
xnor U13255 (N_13255,N_12519,N_12970);
xor U13256 (N_13256,N_12970,N_12836);
or U13257 (N_13257,N_12718,N_12759);
nor U13258 (N_13258,N_12687,N_12609);
nor U13259 (N_13259,N_12667,N_12703);
or U13260 (N_13260,N_12878,N_12535);
xor U13261 (N_13261,N_12694,N_12861);
and U13262 (N_13262,N_12854,N_12662);
nor U13263 (N_13263,N_12675,N_12531);
nor U13264 (N_13264,N_12746,N_12848);
or U13265 (N_13265,N_12808,N_12764);
nor U13266 (N_13266,N_12524,N_12780);
xor U13267 (N_13267,N_12647,N_12816);
or U13268 (N_13268,N_12712,N_12570);
nor U13269 (N_13269,N_12632,N_12814);
and U13270 (N_13270,N_12910,N_12885);
and U13271 (N_13271,N_12819,N_12875);
nor U13272 (N_13272,N_12974,N_12639);
nand U13273 (N_13273,N_12634,N_12983);
xor U13274 (N_13274,N_12986,N_12864);
nor U13275 (N_13275,N_12692,N_12731);
or U13276 (N_13276,N_12945,N_12529);
or U13277 (N_13277,N_12846,N_12869);
nand U13278 (N_13278,N_12927,N_12756);
nor U13279 (N_13279,N_12870,N_12798);
and U13280 (N_13280,N_12924,N_12659);
and U13281 (N_13281,N_12615,N_12786);
nor U13282 (N_13282,N_12673,N_12835);
nand U13283 (N_13283,N_12765,N_12762);
nand U13284 (N_13284,N_12852,N_12725);
nor U13285 (N_13285,N_12559,N_12665);
or U13286 (N_13286,N_12932,N_12628);
or U13287 (N_13287,N_12531,N_12879);
and U13288 (N_13288,N_12576,N_12836);
nand U13289 (N_13289,N_12518,N_12628);
nand U13290 (N_13290,N_12794,N_12959);
or U13291 (N_13291,N_12914,N_12890);
or U13292 (N_13292,N_12552,N_12971);
xor U13293 (N_13293,N_12574,N_12556);
or U13294 (N_13294,N_12611,N_12613);
and U13295 (N_13295,N_12785,N_12532);
or U13296 (N_13296,N_12789,N_12985);
xnor U13297 (N_13297,N_12565,N_12878);
or U13298 (N_13298,N_12870,N_12579);
or U13299 (N_13299,N_12887,N_12607);
or U13300 (N_13300,N_12523,N_12827);
or U13301 (N_13301,N_12817,N_12678);
and U13302 (N_13302,N_12837,N_12851);
xnor U13303 (N_13303,N_12649,N_12952);
xor U13304 (N_13304,N_12569,N_12667);
and U13305 (N_13305,N_12708,N_12646);
or U13306 (N_13306,N_12825,N_12863);
nand U13307 (N_13307,N_12651,N_12719);
and U13308 (N_13308,N_12689,N_12775);
or U13309 (N_13309,N_12649,N_12799);
xor U13310 (N_13310,N_12643,N_12817);
and U13311 (N_13311,N_12707,N_12920);
nand U13312 (N_13312,N_12612,N_12828);
nand U13313 (N_13313,N_12949,N_12895);
xnor U13314 (N_13314,N_12632,N_12665);
nand U13315 (N_13315,N_12781,N_12576);
or U13316 (N_13316,N_12991,N_12504);
nand U13317 (N_13317,N_12528,N_12572);
nor U13318 (N_13318,N_12805,N_12736);
xor U13319 (N_13319,N_12887,N_12654);
nand U13320 (N_13320,N_12734,N_12964);
nor U13321 (N_13321,N_12688,N_12735);
nor U13322 (N_13322,N_12539,N_12502);
nor U13323 (N_13323,N_12701,N_12700);
nand U13324 (N_13324,N_12660,N_12538);
and U13325 (N_13325,N_12689,N_12715);
xnor U13326 (N_13326,N_12688,N_12659);
nand U13327 (N_13327,N_12870,N_12968);
or U13328 (N_13328,N_12552,N_12961);
xor U13329 (N_13329,N_12794,N_12671);
nand U13330 (N_13330,N_12515,N_12851);
xor U13331 (N_13331,N_12947,N_12704);
nor U13332 (N_13332,N_12829,N_12805);
nand U13333 (N_13333,N_12827,N_12536);
xnor U13334 (N_13334,N_12999,N_12663);
and U13335 (N_13335,N_12720,N_12666);
nand U13336 (N_13336,N_12894,N_12798);
xnor U13337 (N_13337,N_12860,N_12848);
nand U13338 (N_13338,N_12993,N_12562);
or U13339 (N_13339,N_12867,N_12814);
or U13340 (N_13340,N_12562,N_12720);
or U13341 (N_13341,N_12690,N_12893);
nor U13342 (N_13342,N_12666,N_12703);
and U13343 (N_13343,N_12645,N_12802);
xor U13344 (N_13344,N_12983,N_12949);
and U13345 (N_13345,N_12827,N_12930);
nand U13346 (N_13346,N_12689,N_12619);
nand U13347 (N_13347,N_12976,N_12813);
nor U13348 (N_13348,N_12547,N_12952);
and U13349 (N_13349,N_12667,N_12854);
xor U13350 (N_13350,N_12600,N_12647);
or U13351 (N_13351,N_12519,N_12738);
xor U13352 (N_13352,N_12644,N_12708);
and U13353 (N_13353,N_12794,N_12506);
and U13354 (N_13354,N_12904,N_12757);
or U13355 (N_13355,N_12838,N_12670);
xnor U13356 (N_13356,N_12987,N_12980);
xnor U13357 (N_13357,N_12666,N_12641);
nor U13358 (N_13358,N_12705,N_12509);
nand U13359 (N_13359,N_12918,N_12542);
nor U13360 (N_13360,N_12760,N_12764);
or U13361 (N_13361,N_12917,N_12704);
nand U13362 (N_13362,N_12794,N_12695);
or U13363 (N_13363,N_12754,N_12635);
nor U13364 (N_13364,N_12926,N_12504);
xor U13365 (N_13365,N_12763,N_12982);
and U13366 (N_13366,N_12892,N_12911);
xnor U13367 (N_13367,N_12959,N_12730);
or U13368 (N_13368,N_12702,N_12554);
and U13369 (N_13369,N_12899,N_12672);
xor U13370 (N_13370,N_12988,N_12736);
nor U13371 (N_13371,N_12703,N_12819);
or U13372 (N_13372,N_12507,N_12843);
xnor U13373 (N_13373,N_12606,N_12578);
xnor U13374 (N_13374,N_12636,N_12970);
nor U13375 (N_13375,N_12760,N_12852);
xor U13376 (N_13376,N_12825,N_12596);
and U13377 (N_13377,N_12708,N_12567);
and U13378 (N_13378,N_12936,N_12510);
nor U13379 (N_13379,N_12741,N_12722);
or U13380 (N_13380,N_12782,N_12886);
xnor U13381 (N_13381,N_12776,N_12887);
nor U13382 (N_13382,N_12779,N_12672);
xor U13383 (N_13383,N_12925,N_12976);
nor U13384 (N_13384,N_12836,N_12865);
or U13385 (N_13385,N_12507,N_12643);
or U13386 (N_13386,N_12748,N_12786);
xor U13387 (N_13387,N_12575,N_12799);
nand U13388 (N_13388,N_12634,N_12929);
and U13389 (N_13389,N_12812,N_12814);
nor U13390 (N_13390,N_12972,N_12977);
xor U13391 (N_13391,N_12817,N_12563);
xor U13392 (N_13392,N_12882,N_12634);
nor U13393 (N_13393,N_12720,N_12682);
or U13394 (N_13394,N_12820,N_12868);
nand U13395 (N_13395,N_12673,N_12879);
xnor U13396 (N_13396,N_12596,N_12537);
nand U13397 (N_13397,N_12802,N_12971);
xor U13398 (N_13398,N_12536,N_12572);
and U13399 (N_13399,N_12619,N_12684);
xnor U13400 (N_13400,N_12889,N_12923);
xor U13401 (N_13401,N_12564,N_12687);
nand U13402 (N_13402,N_12790,N_12802);
nand U13403 (N_13403,N_12674,N_12862);
nor U13404 (N_13404,N_12823,N_12568);
or U13405 (N_13405,N_12783,N_12520);
nor U13406 (N_13406,N_12586,N_12915);
nor U13407 (N_13407,N_12756,N_12972);
nor U13408 (N_13408,N_12819,N_12938);
or U13409 (N_13409,N_12763,N_12640);
or U13410 (N_13410,N_12726,N_12640);
xor U13411 (N_13411,N_12693,N_12662);
nand U13412 (N_13412,N_12632,N_12695);
and U13413 (N_13413,N_12930,N_12689);
xor U13414 (N_13414,N_12536,N_12916);
and U13415 (N_13415,N_12711,N_12983);
xnor U13416 (N_13416,N_12830,N_12749);
xnor U13417 (N_13417,N_12668,N_12582);
or U13418 (N_13418,N_12695,N_12513);
or U13419 (N_13419,N_12897,N_12957);
and U13420 (N_13420,N_12901,N_12724);
nand U13421 (N_13421,N_12560,N_12964);
xnor U13422 (N_13422,N_12500,N_12930);
or U13423 (N_13423,N_12668,N_12570);
nor U13424 (N_13424,N_12707,N_12818);
nand U13425 (N_13425,N_12917,N_12644);
nor U13426 (N_13426,N_12508,N_12989);
and U13427 (N_13427,N_12777,N_12608);
and U13428 (N_13428,N_12945,N_12763);
or U13429 (N_13429,N_12735,N_12868);
xnor U13430 (N_13430,N_12972,N_12707);
or U13431 (N_13431,N_12561,N_12783);
and U13432 (N_13432,N_12719,N_12519);
nand U13433 (N_13433,N_12818,N_12782);
nor U13434 (N_13434,N_12964,N_12777);
and U13435 (N_13435,N_12595,N_12741);
nor U13436 (N_13436,N_12647,N_12526);
or U13437 (N_13437,N_12694,N_12817);
nor U13438 (N_13438,N_12762,N_12547);
nor U13439 (N_13439,N_12785,N_12943);
nand U13440 (N_13440,N_12762,N_12841);
xor U13441 (N_13441,N_12899,N_12737);
xor U13442 (N_13442,N_12935,N_12835);
or U13443 (N_13443,N_12592,N_12574);
or U13444 (N_13444,N_12790,N_12758);
nor U13445 (N_13445,N_12740,N_12652);
xor U13446 (N_13446,N_12816,N_12757);
nor U13447 (N_13447,N_12933,N_12726);
and U13448 (N_13448,N_12629,N_12793);
nand U13449 (N_13449,N_12756,N_12605);
nor U13450 (N_13450,N_12877,N_12972);
or U13451 (N_13451,N_12846,N_12534);
nand U13452 (N_13452,N_12614,N_12789);
xor U13453 (N_13453,N_12714,N_12871);
or U13454 (N_13454,N_12803,N_12725);
and U13455 (N_13455,N_12819,N_12957);
or U13456 (N_13456,N_12996,N_12986);
nand U13457 (N_13457,N_12757,N_12862);
nand U13458 (N_13458,N_12995,N_12736);
or U13459 (N_13459,N_12828,N_12789);
xnor U13460 (N_13460,N_12580,N_12781);
or U13461 (N_13461,N_12867,N_12588);
nand U13462 (N_13462,N_12570,N_12989);
and U13463 (N_13463,N_12667,N_12997);
nor U13464 (N_13464,N_12799,N_12550);
or U13465 (N_13465,N_12551,N_12789);
and U13466 (N_13466,N_12662,N_12780);
or U13467 (N_13467,N_12675,N_12583);
and U13468 (N_13468,N_12993,N_12507);
xnor U13469 (N_13469,N_12582,N_12572);
nand U13470 (N_13470,N_12670,N_12639);
and U13471 (N_13471,N_12642,N_12822);
nor U13472 (N_13472,N_12557,N_12501);
nand U13473 (N_13473,N_12947,N_12584);
and U13474 (N_13474,N_12881,N_12597);
nand U13475 (N_13475,N_12805,N_12695);
xor U13476 (N_13476,N_12552,N_12749);
xor U13477 (N_13477,N_12949,N_12540);
nand U13478 (N_13478,N_12601,N_12590);
and U13479 (N_13479,N_12969,N_12585);
nor U13480 (N_13480,N_12914,N_12724);
xor U13481 (N_13481,N_12535,N_12680);
xnor U13482 (N_13482,N_12875,N_12888);
or U13483 (N_13483,N_12880,N_12513);
nor U13484 (N_13484,N_12818,N_12848);
xnor U13485 (N_13485,N_12555,N_12641);
xnor U13486 (N_13486,N_12572,N_12800);
xnor U13487 (N_13487,N_12961,N_12712);
nand U13488 (N_13488,N_12791,N_12951);
nand U13489 (N_13489,N_12649,N_12935);
or U13490 (N_13490,N_12966,N_12679);
or U13491 (N_13491,N_12847,N_12628);
and U13492 (N_13492,N_12872,N_12549);
xor U13493 (N_13493,N_12922,N_12641);
nand U13494 (N_13494,N_12690,N_12718);
xor U13495 (N_13495,N_12833,N_12798);
xnor U13496 (N_13496,N_12515,N_12911);
or U13497 (N_13497,N_12891,N_12605);
nand U13498 (N_13498,N_12678,N_12985);
xnor U13499 (N_13499,N_12723,N_12743);
or U13500 (N_13500,N_13245,N_13426);
or U13501 (N_13501,N_13109,N_13266);
nor U13502 (N_13502,N_13022,N_13277);
and U13503 (N_13503,N_13477,N_13211);
nand U13504 (N_13504,N_13081,N_13250);
and U13505 (N_13505,N_13310,N_13028);
nand U13506 (N_13506,N_13382,N_13078);
nand U13507 (N_13507,N_13052,N_13185);
and U13508 (N_13508,N_13229,N_13169);
xnor U13509 (N_13509,N_13137,N_13497);
nand U13510 (N_13510,N_13494,N_13308);
and U13511 (N_13511,N_13369,N_13255);
xor U13512 (N_13512,N_13462,N_13468);
and U13513 (N_13513,N_13150,N_13033);
nand U13514 (N_13514,N_13068,N_13044);
xor U13515 (N_13515,N_13456,N_13241);
or U13516 (N_13516,N_13322,N_13227);
nor U13517 (N_13517,N_13433,N_13180);
and U13518 (N_13518,N_13399,N_13370);
nand U13519 (N_13519,N_13067,N_13305);
xor U13520 (N_13520,N_13298,N_13492);
nor U13521 (N_13521,N_13351,N_13306);
or U13522 (N_13522,N_13095,N_13270);
or U13523 (N_13523,N_13457,N_13034);
xnor U13524 (N_13524,N_13124,N_13316);
or U13525 (N_13525,N_13233,N_13285);
xor U13526 (N_13526,N_13215,N_13410);
nand U13527 (N_13527,N_13222,N_13191);
nand U13528 (N_13528,N_13337,N_13036);
xnor U13529 (N_13529,N_13404,N_13443);
or U13530 (N_13530,N_13471,N_13455);
nand U13531 (N_13531,N_13148,N_13093);
and U13532 (N_13532,N_13321,N_13096);
xnor U13533 (N_13533,N_13166,N_13214);
xnor U13534 (N_13534,N_13323,N_13029);
and U13535 (N_13535,N_13261,N_13007);
nor U13536 (N_13536,N_13393,N_13338);
xor U13537 (N_13537,N_13284,N_13339);
or U13538 (N_13538,N_13098,N_13485);
or U13539 (N_13539,N_13319,N_13289);
nor U13540 (N_13540,N_13445,N_13402);
and U13541 (N_13541,N_13479,N_13063);
and U13542 (N_13542,N_13372,N_13080);
or U13543 (N_13543,N_13307,N_13400);
and U13544 (N_13544,N_13186,N_13299);
nand U13545 (N_13545,N_13210,N_13248);
and U13546 (N_13546,N_13085,N_13315);
xnor U13547 (N_13547,N_13458,N_13171);
or U13548 (N_13548,N_13403,N_13343);
xnor U13549 (N_13549,N_13398,N_13173);
or U13550 (N_13550,N_13160,N_13046);
and U13551 (N_13551,N_13106,N_13431);
xnor U13552 (N_13552,N_13019,N_13149);
nor U13553 (N_13553,N_13060,N_13381);
nor U13554 (N_13554,N_13174,N_13048);
and U13555 (N_13555,N_13206,N_13413);
nor U13556 (N_13556,N_13142,N_13459);
or U13557 (N_13557,N_13450,N_13467);
or U13558 (N_13558,N_13056,N_13444);
xnor U13559 (N_13559,N_13113,N_13355);
nand U13560 (N_13560,N_13010,N_13040);
nand U13561 (N_13561,N_13348,N_13358);
and U13562 (N_13562,N_13179,N_13073);
or U13563 (N_13563,N_13421,N_13001);
and U13564 (N_13564,N_13202,N_13251);
or U13565 (N_13565,N_13053,N_13205);
nand U13566 (N_13566,N_13138,N_13181);
xor U13567 (N_13567,N_13126,N_13201);
or U13568 (N_13568,N_13324,N_13386);
and U13569 (N_13569,N_13216,N_13309);
and U13570 (N_13570,N_13195,N_13000);
or U13571 (N_13571,N_13237,N_13074);
and U13572 (N_13572,N_13139,N_13239);
nor U13573 (N_13573,N_13318,N_13384);
or U13574 (N_13574,N_13268,N_13127);
xor U13575 (N_13575,N_13020,N_13292);
or U13576 (N_13576,N_13466,N_13432);
nand U13577 (N_13577,N_13165,N_13434);
xor U13578 (N_13578,N_13291,N_13273);
xor U13579 (N_13579,N_13389,N_13008);
xor U13580 (N_13580,N_13234,N_13325);
nand U13581 (N_13581,N_13378,N_13226);
nor U13582 (N_13582,N_13184,N_13133);
or U13583 (N_13583,N_13446,N_13035);
and U13584 (N_13584,N_13341,N_13363);
nor U13585 (N_13585,N_13107,N_13484);
nor U13586 (N_13586,N_13177,N_13414);
nor U13587 (N_13587,N_13175,N_13076);
or U13588 (N_13588,N_13481,N_13108);
xnor U13589 (N_13589,N_13367,N_13057);
nor U13590 (N_13590,N_13286,N_13437);
or U13591 (N_13591,N_13061,N_13070);
xnor U13592 (N_13592,N_13238,N_13130);
and U13593 (N_13593,N_13397,N_13167);
nor U13594 (N_13594,N_13087,N_13408);
xor U13595 (N_13595,N_13352,N_13263);
xor U13596 (N_13596,N_13418,N_13474);
or U13597 (N_13597,N_13114,N_13111);
or U13598 (N_13598,N_13366,N_13027);
nand U13599 (N_13599,N_13064,N_13015);
nand U13600 (N_13600,N_13031,N_13193);
nand U13601 (N_13601,N_13331,N_13042);
or U13602 (N_13602,N_13153,N_13496);
xnor U13603 (N_13603,N_13427,N_13281);
nor U13604 (N_13604,N_13303,N_13376);
and U13605 (N_13605,N_13349,N_13272);
xnor U13606 (N_13606,N_13163,N_13041);
or U13607 (N_13607,N_13448,N_13082);
nor U13608 (N_13608,N_13116,N_13221);
and U13609 (N_13609,N_13112,N_13375);
and U13610 (N_13610,N_13212,N_13131);
nand U13611 (N_13611,N_13275,N_13037);
or U13612 (N_13612,N_13145,N_13017);
and U13613 (N_13613,N_13203,N_13065);
and U13614 (N_13614,N_13235,N_13155);
nand U13615 (N_13615,N_13183,N_13430);
or U13616 (N_13616,N_13354,N_13334);
or U13617 (N_13617,N_13220,N_13353);
or U13618 (N_13618,N_13049,N_13092);
nor U13619 (N_13619,N_13194,N_13428);
xor U13620 (N_13620,N_13293,N_13200);
xor U13621 (N_13621,N_13254,N_13151);
and U13622 (N_13622,N_13333,N_13253);
nand U13623 (N_13623,N_13083,N_13192);
and U13624 (N_13624,N_13482,N_13249);
and U13625 (N_13625,N_13438,N_13416);
nor U13626 (N_13626,N_13223,N_13103);
or U13627 (N_13627,N_13209,N_13359);
and U13628 (N_13628,N_13290,N_13328);
xnor U13629 (N_13629,N_13077,N_13391);
and U13630 (N_13630,N_13236,N_13023);
nor U13631 (N_13631,N_13314,N_13213);
nand U13632 (N_13632,N_13217,N_13388);
xnor U13633 (N_13633,N_13276,N_13039);
xor U13634 (N_13634,N_13377,N_13417);
nor U13635 (N_13635,N_13099,N_13486);
xor U13636 (N_13636,N_13360,N_13004);
or U13637 (N_13637,N_13278,N_13009);
nand U13638 (N_13638,N_13154,N_13038);
and U13639 (N_13639,N_13178,N_13346);
and U13640 (N_13640,N_13021,N_13483);
nor U13641 (N_13641,N_13075,N_13495);
or U13642 (N_13642,N_13232,N_13101);
and U13643 (N_13643,N_13461,N_13357);
and U13644 (N_13644,N_13032,N_13062);
or U13645 (N_13645,N_13091,N_13228);
nor U13646 (N_13646,N_13045,N_13287);
and U13647 (N_13647,N_13396,N_13415);
or U13648 (N_13648,N_13409,N_13204);
or U13649 (N_13649,N_13442,N_13014);
and U13650 (N_13650,N_13365,N_13125);
nor U13651 (N_13651,N_13244,N_13240);
nand U13652 (N_13652,N_13487,N_13050);
or U13653 (N_13653,N_13436,N_13447);
or U13654 (N_13654,N_13387,N_13122);
xor U13655 (N_13655,N_13297,N_13419);
nor U13656 (N_13656,N_13412,N_13025);
or U13657 (N_13657,N_13470,N_13347);
nand U13658 (N_13658,N_13401,N_13146);
nand U13659 (N_13659,N_13311,N_13441);
xnor U13660 (N_13660,N_13104,N_13158);
nor U13661 (N_13661,N_13491,N_13439);
or U13662 (N_13662,N_13288,N_13219);
nor U13663 (N_13663,N_13094,N_13243);
or U13664 (N_13664,N_13018,N_13199);
or U13665 (N_13665,N_13498,N_13320);
and U13666 (N_13666,N_13465,N_13383);
xor U13667 (N_13667,N_13252,N_13472);
or U13668 (N_13668,N_13312,N_13089);
xor U13669 (N_13669,N_13463,N_13368);
xor U13670 (N_13670,N_13256,N_13188);
and U13671 (N_13671,N_13043,N_13207);
nor U13672 (N_13672,N_13003,N_13144);
nand U13673 (N_13673,N_13301,N_13120);
xnor U13674 (N_13674,N_13262,N_13069);
xnor U13675 (N_13675,N_13478,N_13411);
nor U13676 (N_13676,N_13128,N_13105);
nand U13677 (N_13677,N_13313,N_13379);
nor U13678 (N_13678,N_13394,N_13016);
and U13679 (N_13679,N_13157,N_13282);
nand U13680 (N_13680,N_13086,N_13344);
xor U13681 (N_13681,N_13161,N_13072);
nand U13682 (N_13682,N_13326,N_13134);
xnor U13683 (N_13683,N_13176,N_13420);
or U13684 (N_13684,N_13265,N_13187);
xnor U13685 (N_13685,N_13279,N_13300);
nand U13686 (N_13686,N_13364,N_13118);
nand U13687 (N_13687,N_13090,N_13168);
nor U13688 (N_13688,N_13147,N_13493);
xor U13689 (N_13689,N_13115,N_13005);
and U13690 (N_13690,N_13373,N_13225);
or U13691 (N_13691,N_13135,N_13395);
nand U13692 (N_13692,N_13159,N_13451);
xnor U13693 (N_13693,N_13058,N_13051);
and U13694 (N_13694,N_13182,N_13336);
xor U13695 (N_13695,N_13264,N_13260);
nand U13696 (N_13696,N_13280,N_13423);
nand U13697 (N_13697,N_13475,N_13361);
and U13698 (N_13698,N_13452,N_13059);
and U13699 (N_13699,N_13390,N_13224);
or U13700 (N_13700,N_13488,N_13231);
nand U13701 (N_13701,N_13121,N_13392);
nor U13702 (N_13702,N_13296,N_13047);
xnor U13703 (N_13703,N_13340,N_13380);
or U13704 (N_13704,N_13164,N_13242);
xor U13705 (N_13705,N_13294,N_13196);
nand U13706 (N_13706,N_13097,N_13117);
and U13707 (N_13707,N_13405,N_13156);
nor U13708 (N_13708,N_13295,N_13317);
xor U13709 (N_13709,N_13274,N_13257);
xor U13710 (N_13710,N_13335,N_13198);
or U13711 (N_13711,N_13464,N_13030);
xnor U13712 (N_13712,N_13102,N_13489);
nor U13713 (N_13713,N_13302,N_13304);
nor U13714 (N_13714,N_13197,N_13271);
nand U13715 (N_13715,N_13269,N_13162);
or U13716 (N_13716,N_13329,N_13327);
and U13717 (N_13717,N_13362,N_13259);
and U13718 (N_13718,N_13371,N_13406);
xor U13719 (N_13719,N_13480,N_13453);
nor U13720 (N_13720,N_13100,N_13189);
nor U13721 (N_13721,N_13267,N_13407);
xnor U13722 (N_13722,N_13345,N_13440);
and U13723 (N_13723,N_13385,N_13476);
nand U13724 (N_13724,N_13071,N_13013);
nor U13725 (N_13725,N_13123,N_13152);
and U13726 (N_13726,N_13119,N_13460);
nor U13727 (N_13727,N_13054,N_13247);
or U13728 (N_13728,N_13429,N_13230);
xnor U13729 (N_13729,N_13258,N_13129);
nand U13730 (N_13730,N_13435,N_13218);
nor U13731 (N_13731,N_13332,N_13011);
xor U13732 (N_13732,N_13141,N_13425);
and U13733 (N_13733,N_13342,N_13374);
nand U13734 (N_13734,N_13110,N_13055);
nand U13735 (N_13735,N_13208,N_13002);
xnor U13736 (N_13736,N_13469,N_13356);
or U13737 (N_13737,N_13490,N_13422);
xnor U13738 (N_13738,N_13026,N_13012);
xor U13739 (N_13739,N_13449,N_13136);
nand U13740 (N_13740,N_13140,N_13283);
xnor U13741 (N_13741,N_13006,N_13350);
and U13742 (N_13742,N_13454,N_13143);
nand U13743 (N_13743,N_13330,N_13084);
or U13744 (N_13744,N_13132,N_13088);
nand U13745 (N_13745,N_13499,N_13424);
or U13746 (N_13746,N_13024,N_13079);
xnor U13747 (N_13747,N_13066,N_13190);
nor U13748 (N_13748,N_13170,N_13172);
nand U13749 (N_13749,N_13473,N_13246);
or U13750 (N_13750,N_13280,N_13326);
and U13751 (N_13751,N_13030,N_13484);
and U13752 (N_13752,N_13090,N_13348);
and U13753 (N_13753,N_13363,N_13159);
nor U13754 (N_13754,N_13052,N_13263);
nand U13755 (N_13755,N_13158,N_13395);
and U13756 (N_13756,N_13205,N_13051);
and U13757 (N_13757,N_13109,N_13218);
nand U13758 (N_13758,N_13145,N_13220);
or U13759 (N_13759,N_13046,N_13307);
nand U13760 (N_13760,N_13110,N_13074);
and U13761 (N_13761,N_13124,N_13058);
nand U13762 (N_13762,N_13074,N_13308);
or U13763 (N_13763,N_13473,N_13013);
or U13764 (N_13764,N_13085,N_13048);
nor U13765 (N_13765,N_13082,N_13268);
nor U13766 (N_13766,N_13233,N_13186);
nor U13767 (N_13767,N_13048,N_13306);
or U13768 (N_13768,N_13042,N_13463);
and U13769 (N_13769,N_13078,N_13196);
and U13770 (N_13770,N_13152,N_13446);
nand U13771 (N_13771,N_13466,N_13137);
nor U13772 (N_13772,N_13311,N_13135);
and U13773 (N_13773,N_13322,N_13037);
or U13774 (N_13774,N_13097,N_13095);
nand U13775 (N_13775,N_13443,N_13070);
or U13776 (N_13776,N_13324,N_13229);
or U13777 (N_13777,N_13348,N_13479);
and U13778 (N_13778,N_13333,N_13442);
xor U13779 (N_13779,N_13492,N_13340);
nand U13780 (N_13780,N_13310,N_13141);
xnor U13781 (N_13781,N_13207,N_13246);
and U13782 (N_13782,N_13140,N_13438);
and U13783 (N_13783,N_13475,N_13075);
and U13784 (N_13784,N_13288,N_13384);
nand U13785 (N_13785,N_13096,N_13437);
nand U13786 (N_13786,N_13286,N_13355);
nand U13787 (N_13787,N_13173,N_13492);
and U13788 (N_13788,N_13043,N_13053);
xnor U13789 (N_13789,N_13190,N_13247);
nand U13790 (N_13790,N_13208,N_13081);
nor U13791 (N_13791,N_13246,N_13371);
nor U13792 (N_13792,N_13425,N_13097);
nor U13793 (N_13793,N_13420,N_13294);
nand U13794 (N_13794,N_13023,N_13096);
nor U13795 (N_13795,N_13298,N_13044);
nor U13796 (N_13796,N_13380,N_13473);
xnor U13797 (N_13797,N_13161,N_13343);
nor U13798 (N_13798,N_13000,N_13277);
or U13799 (N_13799,N_13293,N_13457);
nor U13800 (N_13800,N_13217,N_13393);
nor U13801 (N_13801,N_13063,N_13055);
and U13802 (N_13802,N_13198,N_13484);
nand U13803 (N_13803,N_13231,N_13089);
or U13804 (N_13804,N_13192,N_13146);
nor U13805 (N_13805,N_13064,N_13239);
or U13806 (N_13806,N_13163,N_13119);
nand U13807 (N_13807,N_13216,N_13371);
xnor U13808 (N_13808,N_13245,N_13139);
nand U13809 (N_13809,N_13358,N_13316);
xor U13810 (N_13810,N_13106,N_13409);
nand U13811 (N_13811,N_13111,N_13432);
or U13812 (N_13812,N_13331,N_13029);
nand U13813 (N_13813,N_13433,N_13014);
xor U13814 (N_13814,N_13411,N_13389);
nand U13815 (N_13815,N_13088,N_13363);
nand U13816 (N_13816,N_13206,N_13144);
nand U13817 (N_13817,N_13087,N_13086);
or U13818 (N_13818,N_13313,N_13254);
xor U13819 (N_13819,N_13006,N_13295);
and U13820 (N_13820,N_13046,N_13029);
nand U13821 (N_13821,N_13368,N_13258);
xnor U13822 (N_13822,N_13021,N_13037);
xnor U13823 (N_13823,N_13253,N_13243);
nand U13824 (N_13824,N_13195,N_13244);
nand U13825 (N_13825,N_13057,N_13325);
nor U13826 (N_13826,N_13336,N_13089);
nand U13827 (N_13827,N_13399,N_13449);
nor U13828 (N_13828,N_13398,N_13229);
nor U13829 (N_13829,N_13364,N_13214);
xnor U13830 (N_13830,N_13029,N_13395);
xnor U13831 (N_13831,N_13086,N_13402);
xor U13832 (N_13832,N_13114,N_13444);
and U13833 (N_13833,N_13356,N_13409);
xnor U13834 (N_13834,N_13293,N_13425);
nand U13835 (N_13835,N_13464,N_13119);
xor U13836 (N_13836,N_13457,N_13307);
nor U13837 (N_13837,N_13312,N_13499);
nor U13838 (N_13838,N_13080,N_13265);
xnor U13839 (N_13839,N_13152,N_13363);
xor U13840 (N_13840,N_13217,N_13159);
xnor U13841 (N_13841,N_13181,N_13250);
xor U13842 (N_13842,N_13480,N_13473);
nor U13843 (N_13843,N_13055,N_13147);
and U13844 (N_13844,N_13205,N_13353);
nor U13845 (N_13845,N_13275,N_13309);
and U13846 (N_13846,N_13068,N_13408);
nor U13847 (N_13847,N_13163,N_13030);
nor U13848 (N_13848,N_13078,N_13208);
and U13849 (N_13849,N_13495,N_13077);
xnor U13850 (N_13850,N_13433,N_13050);
and U13851 (N_13851,N_13095,N_13493);
nand U13852 (N_13852,N_13441,N_13240);
nor U13853 (N_13853,N_13431,N_13005);
or U13854 (N_13854,N_13246,N_13189);
nand U13855 (N_13855,N_13003,N_13066);
or U13856 (N_13856,N_13040,N_13493);
nor U13857 (N_13857,N_13268,N_13397);
nand U13858 (N_13858,N_13280,N_13045);
or U13859 (N_13859,N_13101,N_13225);
or U13860 (N_13860,N_13035,N_13110);
and U13861 (N_13861,N_13423,N_13033);
nor U13862 (N_13862,N_13429,N_13051);
or U13863 (N_13863,N_13054,N_13168);
xnor U13864 (N_13864,N_13003,N_13289);
nand U13865 (N_13865,N_13111,N_13188);
nand U13866 (N_13866,N_13116,N_13019);
xnor U13867 (N_13867,N_13054,N_13474);
xor U13868 (N_13868,N_13149,N_13152);
or U13869 (N_13869,N_13385,N_13280);
nand U13870 (N_13870,N_13131,N_13421);
xor U13871 (N_13871,N_13278,N_13160);
nor U13872 (N_13872,N_13056,N_13412);
and U13873 (N_13873,N_13339,N_13217);
xnor U13874 (N_13874,N_13144,N_13232);
and U13875 (N_13875,N_13182,N_13353);
nor U13876 (N_13876,N_13153,N_13228);
xnor U13877 (N_13877,N_13286,N_13393);
nand U13878 (N_13878,N_13314,N_13419);
and U13879 (N_13879,N_13145,N_13294);
or U13880 (N_13880,N_13144,N_13018);
nand U13881 (N_13881,N_13481,N_13475);
xnor U13882 (N_13882,N_13123,N_13026);
or U13883 (N_13883,N_13417,N_13058);
and U13884 (N_13884,N_13162,N_13436);
nand U13885 (N_13885,N_13380,N_13216);
nand U13886 (N_13886,N_13087,N_13456);
xnor U13887 (N_13887,N_13419,N_13406);
nand U13888 (N_13888,N_13165,N_13052);
xnor U13889 (N_13889,N_13216,N_13199);
or U13890 (N_13890,N_13391,N_13050);
nand U13891 (N_13891,N_13021,N_13329);
xor U13892 (N_13892,N_13347,N_13252);
nand U13893 (N_13893,N_13121,N_13475);
nand U13894 (N_13894,N_13487,N_13453);
nor U13895 (N_13895,N_13074,N_13087);
or U13896 (N_13896,N_13377,N_13089);
nor U13897 (N_13897,N_13182,N_13489);
nand U13898 (N_13898,N_13351,N_13330);
nand U13899 (N_13899,N_13064,N_13393);
or U13900 (N_13900,N_13088,N_13080);
or U13901 (N_13901,N_13352,N_13463);
and U13902 (N_13902,N_13010,N_13028);
nand U13903 (N_13903,N_13329,N_13091);
or U13904 (N_13904,N_13082,N_13228);
and U13905 (N_13905,N_13189,N_13096);
or U13906 (N_13906,N_13055,N_13290);
nand U13907 (N_13907,N_13400,N_13473);
or U13908 (N_13908,N_13344,N_13466);
or U13909 (N_13909,N_13205,N_13075);
and U13910 (N_13910,N_13419,N_13251);
nand U13911 (N_13911,N_13301,N_13343);
and U13912 (N_13912,N_13192,N_13338);
nor U13913 (N_13913,N_13328,N_13467);
or U13914 (N_13914,N_13352,N_13367);
and U13915 (N_13915,N_13461,N_13152);
and U13916 (N_13916,N_13291,N_13160);
xor U13917 (N_13917,N_13485,N_13330);
xor U13918 (N_13918,N_13333,N_13117);
xnor U13919 (N_13919,N_13486,N_13180);
nor U13920 (N_13920,N_13182,N_13194);
xnor U13921 (N_13921,N_13115,N_13113);
nand U13922 (N_13922,N_13395,N_13469);
and U13923 (N_13923,N_13320,N_13043);
and U13924 (N_13924,N_13312,N_13084);
and U13925 (N_13925,N_13108,N_13438);
xnor U13926 (N_13926,N_13096,N_13460);
xnor U13927 (N_13927,N_13200,N_13276);
or U13928 (N_13928,N_13060,N_13054);
xnor U13929 (N_13929,N_13133,N_13032);
xnor U13930 (N_13930,N_13249,N_13112);
or U13931 (N_13931,N_13243,N_13465);
nand U13932 (N_13932,N_13132,N_13350);
and U13933 (N_13933,N_13323,N_13182);
nand U13934 (N_13934,N_13442,N_13186);
and U13935 (N_13935,N_13423,N_13135);
xnor U13936 (N_13936,N_13309,N_13355);
and U13937 (N_13937,N_13033,N_13026);
and U13938 (N_13938,N_13424,N_13270);
xnor U13939 (N_13939,N_13138,N_13278);
xor U13940 (N_13940,N_13246,N_13389);
and U13941 (N_13941,N_13440,N_13149);
xnor U13942 (N_13942,N_13029,N_13496);
nand U13943 (N_13943,N_13387,N_13108);
xor U13944 (N_13944,N_13493,N_13261);
and U13945 (N_13945,N_13126,N_13295);
or U13946 (N_13946,N_13119,N_13300);
nand U13947 (N_13947,N_13288,N_13266);
or U13948 (N_13948,N_13137,N_13467);
or U13949 (N_13949,N_13015,N_13088);
xnor U13950 (N_13950,N_13108,N_13279);
nor U13951 (N_13951,N_13179,N_13049);
and U13952 (N_13952,N_13441,N_13445);
nor U13953 (N_13953,N_13000,N_13371);
or U13954 (N_13954,N_13496,N_13185);
nor U13955 (N_13955,N_13406,N_13464);
nand U13956 (N_13956,N_13170,N_13263);
xor U13957 (N_13957,N_13206,N_13492);
or U13958 (N_13958,N_13236,N_13313);
xor U13959 (N_13959,N_13385,N_13151);
nand U13960 (N_13960,N_13202,N_13043);
nand U13961 (N_13961,N_13309,N_13201);
nor U13962 (N_13962,N_13470,N_13434);
and U13963 (N_13963,N_13225,N_13313);
xnor U13964 (N_13964,N_13391,N_13453);
nor U13965 (N_13965,N_13031,N_13146);
nor U13966 (N_13966,N_13450,N_13220);
and U13967 (N_13967,N_13160,N_13154);
xor U13968 (N_13968,N_13190,N_13291);
and U13969 (N_13969,N_13421,N_13334);
and U13970 (N_13970,N_13052,N_13213);
xor U13971 (N_13971,N_13046,N_13202);
nand U13972 (N_13972,N_13174,N_13269);
and U13973 (N_13973,N_13396,N_13315);
nor U13974 (N_13974,N_13376,N_13069);
nand U13975 (N_13975,N_13154,N_13094);
or U13976 (N_13976,N_13182,N_13043);
and U13977 (N_13977,N_13283,N_13442);
nand U13978 (N_13978,N_13046,N_13371);
or U13979 (N_13979,N_13226,N_13407);
nor U13980 (N_13980,N_13046,N_13021);
nand U13981 (N_13981,N_13181,N_13228);
nor U13982 (N_13982,N_13487,N_13028);
and U13983 (N_13983,N_13433,N_13073);
nand U13984 (N_13984,N_13101,N_13201);
xnor U13985 (N_13985,N_13448,N_13061);
nand U13986 (N_13986,N_13416,N_13333);
xnor U13987 (N_13987,N_13289,N_13018);
nor U13988 (N_13988,N_13351,N_13304);
nor U13989 (N_13989,N_13181,N_13170);
nor U13990 (N_13990,N_13401,N_13312);
and U13991 (N_13991,N_13307,N_13362);
nand U13992 (N_13992,N_13062,N_13356);
xnor U13993 (N_13993,N_13124,N_13221);
nor U13994 (N_13994,N_13123,N_13120);
and U13995 (N_13995,N_13364,N_13315);
nand U13996 (N_13996,N_13359,N_13328);
nand U13997 (N_13997,N_13055,N_13214);
and U13998 (N_13998,N_13232,N_13352);
xnor U13999 (N_13999,N_13097,N_13247);
and U14000 (N_14000,N_13614,N_13598);
or U14001 (N_14001,N_13522,N_13834);
xnor U14002 (N_14002,N_13688,N_13521);
nand U14003 (N_14003,N_13991,N_13916);
xor U14004 (N_14004,N_13616,N_13778);
nand U14005 (N_14005,N_13979,N_13730);
xnor U14006 (N_14006,N_13569,N_13534);
and U14007 (N_14007,N_13929,N_13937);
nor U14008 (N_14008,N_13506,N_13726);
xor U14009 (N_14009,N_13513,N_13540);
and U14010 (N_14010,N_13802,N_13610);
xor U14011 (N_14011,N_13580,N_13758);
nor U14012 (N_14012,N_13723,N_13938);
xnor U14013 (N_14013,N_13947,N_13561);
or U14014 (N_14014,N_13539,N_13684);
nor U14015 (N_14015,N_13813,N_13989);
and U14016 (N_14016,N_13967,N_13628);
nor U14017 (N_14017,N_13559,N_13946);
xnor U14018 (N_14018,N_13677,N_13724);
nand U14019 (N_14019,N_13959,N_13860);
xor U14020 (N_14020,N_13533,N_13731);
nand U14021 (N_14021,N_13982,N_13769);
xnor U14022 (N_14022,N_13719,N_13952);
xnor U14023 (N_14023,N_13968,N_13969);
xor U14024 (N_14024,N_13741,N_13836);
xnor U14025 (N_14025,N_13873,N_13557);
nand U14026 (N_14026,N_13538,N_13850);
and U14027 (N_14027,N_13858,N_13592);
nand U14028 (N_14028,N_13918,N_13846);
or U14029 (N_14029,N_13915,N_13823);
nor U14030 (N_14030,N_13795,N_13643);
nor U14031 (N_14031,N_13958,N_13537);
and U14032 (N_14032,N_13923,N_13791);
or U14033 (N_14033,N_13505,N_13953);
nor U14034 (N_14034,N_13543,N_13785);
nand U14035 (N_14035,N_13893,N_13531);
and U14036 (N_14036,N_13949,N_13879);
xnor U14037 (N_14037,N_13922,N_13648);
and U14038 (N_14038,N_13805,N_13831);
or U14039 (N_14039,N_13971,N_13530);
xor U14040 (N_14040,N_13963,N_13514);
and U14041 (N_14041,N_13722,N_13933);
nor U14042 (N_14042,N_13705,N_13735);
and U14043 (N_14043,N_13749,N_13606);
or U14044 (N_14044,N_13931,N_13934);
or U14045 (N_14045,N_13595,N_13596);
xor U14046 (N_14046,N_13733,N_13803);
and U14047 (N_14047,N_13551,N_13859);
or U14048 (N_14048,N_13962,N_13609);
xor U14049 (N_14049,N_13636,N_13626);
or U14050 (N_14050,N_13807,N_13891);
nand U14051 (N_14051,N_13732,N_13972);
and U14052 (N_14052,N_13654,N_13605);
xnor U14053 (N_14053,N_13773,N_13789);
xor U14054 (N_14054,N_13644,N_13585);
nor U14055 (N_14055,N_13544,N_13760);
nand U14056 (N_14056,N_13661,N_13627);
nand U14057 (N_14057,N_13686,N_13720);
or U14058 (N_14058,N_13721,N_13509);
nand U14059 (N_14059,N_13608,N_13886);
nor U14060 (N_14060,N_13623,N_13729);
and U14061 (N_14061,N_13560,N_13620);
and U14062 (N_14062,N_13593,N_13675);
xnor U14063 (N_14063,N_13883,N_13502);
or U14064 (N_14064,N_13871,N_13742);
and U14065 (N_14065,N_13619,N_13553);
and U14066 (N_14066,N_13618,N_13896);
or U14067 (N_14067,N_13699,N_13978);
xnor U14068 (N_14068,N_13518,N_13875);
and U14069 (N_14069,N_13783,N_13840);
nor U14070 (N_14070,N_13510,N_13702);
xor U14071 (N_14071,N_13862,N_13578);
or U14072 (N_14072,N_13861,N_13884);
or U14073 (N_14073,N_13881,N_13695);
xor U14074 (N_14074,N_13913,N_13975);
nand U14075 (N_14075,N_13504,N_13709);
nand U14076 (N_14076,N_13945,N_13713);
and U14077 (N_14077,N_13829,N_13910);
or U14078 (N_14078,N_13828,N_13976);
nor U14079 (N_14079,N_13646,N_13926);
and U14080 (N_14080,N_13507,N_13508);
and U14081 (N_14081,N_13579,N_13716);
nor U14082 (N_14082,N_13650,N_13652);
nand U14083 (N_14083,N_13669,N_13545);
nand U14084 (N_14084,N_13762,N_13615);
xnor U14085 (N_14085,N_13747,N_13667);
and U14086 (N_14086,N_13535,N_13740);
xor U14087 (N_14087,N_13679,N_13872);
nor U14088 (N_14088,N_13685,N_13772);
and U14089 (N_14089,N_13629,N_13529);
nand U14090 (N_14090,N_13792,N_13999);
xor U14091 (N_14091,N_13642,N_13784);
or U14092 (N_14092,N_13894,N_13602);
or U14093 (N_14093,N_13798,N_13683);
nand U14094 (N_14094,N_13941,N_13611);
nor U14095 (N_14095,N_13604,N_13564);
and U14096 (N_14096,N_13710,N_13766);
nor U14097 (N_14097,N_13660,N_13787);
xor U14098 (N_14098,N_13764,N_13672);
and U14099 (N_14099,N_13835,N_13866);
nor U14100 (N_14100,N_13919,N_13811);
nand U14101 (N_14101,N_13512,N_13890);
nand U14102 (N_14102,N_13997,N_13700);
nand U14103 (N_14103,N_13630,N_13547);
nor U14104 (N_14104,N_13693,N_13691);
nor U14105 (N_14105,N_13617,N_13590);
and U14106 (N_14106,N_13757,N_13908);
or U14107 (N_14107,N_13704,N_13622);
and U14108 (N_14108,N_13799,N_13689);
and U14109 (N_14109,N_13759,N_13885);
nor U14110 (N_14110,N_13921,N_13820);
and U14111 (N_14111,N_13567,N_13556);
xor U14112 (N_14112,N_13638,N_13532);
or U14113 (N_14113,N_13992,N_13708);
xnor U14114 (N_14114,N_13867,N_13788);
xnor U14115 (N_14115,N_13847,N_13746);
nand U14116 (N_14116,N_13651,N_13956);
xor U14117 (N_14117,N_13523,N_13848);
xnor U14118 (N_14118,N_13712,N_13780);
nand U14119 (N_14119,N_13878,N_13707);
and U14120 (N_14120,N_13570,N_13500);
xor U14121 (N_14121,N_13576,N_13554);
and U14122 (N_14122,N_13656,N_13822);
and U14123 (N_14123,N_13902,N_13815);
nor U14124 (N_14124,N_13857,N_13601);
nor U14125 (N_14125,N_13624,N_13743);
and U14126 (N_14126,N_13550,N_13821);
xnor U14127 (N_14127,N_13899,N_13898);
xor U14128 (N_14128,N_13583,N_13698);
nand U14129 (N_14129,N_13714,N_13892);
or U14130 (N_14130,N_13613,N_13548);
and U14131 (N_14131,N_13806,N_13680);
nand U14132 (N_14132,N_13765,N_13657);
nand U14133 (N_14133,N_13736,N_13571);
xnor U14134 (N_14134,N_13767,N_13897);
or U14135 (N_14135,N_13673,N_13904);
and U14136 (N_14136,N_13663,N_13911);
or U14137 (N_14137,N_13715,N_13837);
nand U14138 (N_14138,N_13819,N_13817);
xnor U14139 (N_14139,N_13718,N_13986);
or U14140 (N_14140,N_13844,N_13943);
xor U14141 (N_14141,N_13725,N_13944);
nand U14142 (N_14142,N_13935,N_13797);
and U14143 (N_14143,N_13965,N_13870);
nand U14144 (N_14144,N_13800,N_13816);
or U14145 (N_14145,N_13964,N_13668);
nor U14146 (N_14146,N_13637,N_13503);
nor U14147 (N_14147,N_13864,N_13818);
and U14148 (N_14148,N_13701,N_13536);
nor U14149 (N_14149,N_13744,N_13666);
or U14150 (N_14150,N_13696,N_13706);
nor U14151 (N_14151,N_13584,N_13856);
and U14152 (N_14152,N_13841,N_13863);
or U14153 (N_14153,N_13768,N_13659);
nor U14154 (N_14154,N_13594,N_13634);
and U14155 (N_14155,N_13801,N_13843);
xor U14156 (N_14156,N_13516,N_13511);
or U14157 (N_14157,N_13542,N_13901);
or U14158 (N_14158,N_13865,N_13808);
and U14159 (N_14159,N_13955,N_13582);
nand U14160 (N_14160,N_13824,N_13525);
nand U14161 (N_14161,N_13854,N_13939);
xor U14162 (N_14162,N_13761,N_13786);
nor U14163 (N_14163,N_13948,N_13640);
nor U14164 (N_14164,N_13527,N_13703);
and U14165 (N_14165,N_13981,N_13670);
xnor U14166 (N_14166,N_13555,N_13526);
nor U14167 (N_14167,N_13794,N_13565);
nor U14168 (N_14168,N_13960,N_13515);
nor U14169 (N_14169,N_13887,N_13809);
or U14170 (N_14170,N_13826,N_13658);
nor U14171 (N_14171,N_13603,N_13562);
nor U14172 (N_14172,N_13552,N_13751);
xnor U14173 (N_14173,N_13868,N_13664);
nand U14174 (N_14174,N_13671,N_13832);
nand U14175 (N_14175,N_13909,N_13574);
nand U14176 (N_14176,N_13833,N_13690);
and U14177 (N_14177,N_13647,N_13903);
nor U14178 (N_14178,N_13546,N_13914);
nand U14179 (N_14179,N_13812,N_13519);
nand U14180 (N_14180,N_13905,N_13734);
and U14181 (N_14181,N_13825,N_13755);
or U14182 (N_14182,N_13612,N_13845);
nor U14183 (N_14183,N_13572,N_13777);
and U14184 (N_14184,N_13853,N_13880);
or U14185 (N_14185,N_13932,N_13951);
xor U14186 (N_14186,N_13995,N_13739);
xnor U14187 (N_14187,N_13961,N_13830);
xor U14188 (N_14188,N_13838,N_13641);
xor U14189 (N_14189,N_13599,N_13876);
nor U14190 (N_14190,N_13600,N_13589);
nor U14191 (N_14191,N_13973,N_13711);
or U14192 (N_14192,N_13756,N_13874);
nand U14193 (N_14193,N_13839,N_13631);
and U14194 (N_14194,N_13804,N_13907);
nor U14195 (N_14195,N_13925,N_13588);
and U14196 (N_14196,N_13639,N_13814);
xnor U14197 (N_14197,N_13983,N_13697);
and U14198 (N_14198,N_13763,N_13662);
nor U14199 (N_14199,N_13842,N_13586);
or U14200 (N_14200,N_13776,N_13737);
and U14201 (N_14201,N_13682,N_13676);
nand U14202 (N_14202,N_13745,N_13541);
and U14203 (N_14203,N_13970,N_13653);
and U14204 (N_14204,N_13581,N_13649);
nand U14205 (N_14205,N_13524,N_13591);
nand U14206 (N_14206,N_13990,N_13984);
and U14207 (N_14207,N_13573,N_13900);
and U14208 (N_14208,N_13575,N_13549);
nand U14209 (N_14209,N_13954,N_13694);
nor U14210 (N_14210,N_13754,N_13888);
nor U14211 (N_14211,N_13936,N_13940);
or U14212 (N_14212,N_13877,N_13950);
nand U14213 (N_14213,N_13752,N_13738);
nor U14214 (N_14214,N_13692,N_13849);
nand U14215 (N_14215,N_13501,N_13987);
nand U14216 (N_14216,N_13577,N_13748);
nand U14217 (N_14217,N_13889,N_13974);
nand U14218 (N_14218,N_13771,N_13996);
nor U14219 (N_14219,N_13942,N_13993);
and U14220 (N_14220,N_13597,N_13966);
nor U14221 (N_14221,N_13681,N_13655);
xnor U14222 (N_14222,N_13727,N_13645);
or U14223 (N_14223,N_13980,N_13796);
and U14224 (N_14224,N_13810,N_13775);
nor U14225 (N_14225,N_13851,N_13852);
nor U14226 (N_14226,N_13920,N_13753);
xor U14227 (N_14227,N_13632,N_13558);
xnor U14228 (N_14228,N_13779,N_13930);
xnor U14229 (N_14229,N_13621,N_13568);
xor U14230 (N_14230,N_13994,N_13790);
xnor U14231 (N_14231,N_13635,N_13927);
nand U14232 (N_14232,N_13678,N_13770);
nand U14233 (N_14233,N_13633,N_13985);
and U14234 (N_14234,N_13563,N_13924);
xor U14235 (N_14235,N_13665,N_13895);
nand U14236 (N_14236,N_13687,N_13674);
nand U14237 (N_14237,N_13781,N_13928);
xnor U14238 (N_14238,N_13607,N_13520);
or U14239 (N_14239,N_13977,N_13750);
nor U14240 (N_14240,N_13793,N_13528);
nand U14241 (N_14241,N_13517,N_13717);
and U14242 (N_14242,N_13957,N_13869);
and U14243 (N_14243,N_13566,N_13882);
nand U14244 (N_14244,N_13988,N_13855);
and U14245 (N_14245,N_13774,N_13728);
xor U14246 (N_14246,N_13998,N_13906);
xnor U14247 (N_14247,N_13782,N_13827);
and U14248 (N_14248,N_13587,N_13917);
or U14249 (N_14249,N_13625,N_13912);
nand U14250 (N_14250,N_13612,N_13823);
nand U14251 (N_14251,N_13965,N_13596);
nand U14252 (N_14252,N_13581,N_13535);
xnor U14253 (N_14253,N_13786,N_13818);
or U14254 (N_14254,N_13796,N_13886);
and U14255 (N_14255,N_13705,N_13715);
and U14256 (N_14256,N_13897,N_13746);
xnor U14257 (N_14257,N_13507,N_13674);
xnor U14258 (N_14258,N_13573,N_13595);
nor U14259 (N_14259,N_13825,N_13611);
and U14260 (N_14260,N_13501,N_13788);
xor U14261 (N_14261,N_13647,N_13854);
nand U14262 (N_14262,N_13969,N_13709);
and U14263 (N_14263,N_13728,N_13576);
xor U14264 (N_14264,N_13606,N_13750);
nand U14265 (N_14265,N_13950,N_13980);
and U14266 (N_14266,N_13831,N_13524);
and U14267 (N_14267,N_13840,N_13647);
nor U14268 (N_14268,N_13913,N_13940);
nand U14269 (N_14269,N_13692,N_13893);
xor U14270 (N_14270,N_13591,N_13530);
xor U14271 (N_14271,N_13638,N_13642);
xor U14272 (N_14272,N_13690,N_13500);
nand U14273 (N_14273,N_13812,N_13829);
and U14274 (N_14274,N_13753,N_13651);
nand U14275 (N_14275,N_13716,N_13917);
nor U14276 (N_14276,N_13899,N_13650);
nand U14277 (N_14277,N_13770,N_13631);
and U14278 (N_14278,N_13803,N_13911);
xnor U14279 (N_14279,N_13827,N_13709);
and U14280 (N_14280,N_13825,N_13826);
nor U14281 (N_14281,N_13882,N_13902);
xnor U14282 (N_14282,N_13917,N_13775);
nand U14283 (N_14283,N_13593,N_13725);
or U14284 (N_14284,N_13784,N_13686);
nor U14285 (N_14285,N_13829,N_13926);
nand U14286 (N_14286,N_13601,N_13700);
xor U14287 (N_14287,N_13940,N_13851);
xor U14288 (N_14288,N_13762,N_13713);
nand U14289 (N_14289,N_13723,N_13819);
nor U14290 (N_14290,N_13629,N_13811);
and U14291 (N_14291,N_13634,N_13866);
nand U14292 (N_14292,N_13714,N_13854);
or U14293 (N_14293,N_13701,N_13920);
xor U14294 (N_14294,N_13695,N_13694);
xor U14295 (N_14295,N_13905,N_13800);
or U14296 (N_14296,N_13538,N_13758);
xnor U14297 (N_14297,N_13547,N_13600);
nor U14298 (N_14298,N_13999,N_13993);
or U14299 (N_14299,N_13727,N_13987);
and U14300 (N_14300,N_13803,N_13761);
nand U14301 (N_14301,N_13543,N_13708);
or U14302 (N_14302,N_13782,N_13663);
nand U14303 (N_14303,N_13932,N_13551);
nand U14304 (N_14304,N_13787,N_13553);
nor U14305 (N_14305,N_13968,N_13531);
or U14306 (N_14306,N_13811,N_13841);
nand U14307 (N_14307,N_13607,N_13765);
and U14308 (N_14308,N_13620,N_13923);
xor U14309 (N_14309,N_13806,N_13979);
nand U14310 (N_14310,N_13608,N_13961);
and U14311 (N_14311,N_13827,N_13892);
nand U14312 (N_14312,N_13904,N_13828);
or U14313 (N_14313,N_13535,N_13995);
and U14314 (N_14314,N_13692,N_13904);
nor U14315 (N_14315,N_13546,N_13841);
or U14316 (N_14316,N_13604,N_13995);
and U14317 (N_14317,N_13832,N_13926);
nor U14318 (N_14318,N_13986,N_13903);
xnor U14319 (N_14319,N_13961,N_13848);
and U14320 (N_14320,N_13844,N_13571);
xor U14321 (N_14321,N_13590,N_13980);
nand U14322 (N_14322,N_13873,N_13676);
nand U14323 (N_14323,N_13987,N_13943);
or U14324 (N_14324,N_13931,N_13981);
xor U14325 (N_14325,N_13563,N_13594);
xor U14326 (N_14326,N_13994,N_13677);
nor U14327 (N_14327,N_13751,N_13825);
xor U14328 (N_14328,N_13738,N_13500);
nor U14329 (N_14329,N_13775,N_13838);
and U14330 (N_14330,N_13915,N_13800);
or U14331 (N_14331,N_13581,N_13599);
xnor U14332 (N_14332,N_13836,N_13776);
nand U14333 (N_14333,N_13693,N_13656);
or U14334 (N_14334,N_13530,N_13890);
or U14335 (N_14335,N_13730,N_13784);
or U14336 (N_14336,N_13942,N_13865);
xor U14337 (N_14337,N_13783,N_13590);
nor U14338 (N_14338,N_13707,N_13673);
or U14339 (N_14339,N_13847,N_13812);
nor U14340 (N_14340,N_13584,N_13503);
nor U14341 (N_14341,N_13571,N_13982);
nor U14342 (N_14342,N_13677,N_13699);
nor U14343 (N_14343,N_13548,N_13667);
nor U14344 (N_14344,N_13978,N_13850);
nor U14345 (N_14345,N_13731,N_13700);
and U14346 (N_14346,N_13933,N_13790);
or U14347 (N_14347,N_13750,N_13971);
nor U14348 (N_14348,N_13880,N_13652);
xor U14349 (N_14349,N_13535,N_13520);
xor U14350 (N_14350,N_13694,N_13559);
or U14351 (N_14351,N_13645,N_13982);
and U14352 (N_14352,N_13943,N_13805);
nor U14353 (N_14353,N_13951,N_13816);
nand U14354 (N_14354,N_13907,N_13921);
and U14355 (N_14355,N_13832,N_13747);
and U14356 (N_14356,N_13985,N_13710);
and U14357 (N_14357,N_13914,N_13761);
nor U14358 (N_14358,N_13599,N_13610);
xnor U14359 (N_14359,N_13608,N_13760);
and U14360 (N_14360,N_13653,N_13980);
xnor U14361 (N_14361,N_13761,N_13956);
or U14362 (N_14362,N_13877,N_13551);
xor U14363 (N_14363,N_13973,N_13749);
nor U14364 (N_14364,N_13878,N_13950);
or U14365 (N_14365,N_13809,N_13696);
or U14366 (N_14366,N_13658,N_13884);
and U14367 (N_14367,N_13816,N_13755);
xor U14368 (N_14368,N_13543,N_13670);
nand U14369 (N_14369,N_13917,N_13619);
nor U14370 (N_14370,N_13844,N_13815);
nand U14371 (N_14371,N_13541,N_13977);
and U14372 (N_14372,N_13776,N_13515);
xor U14373 (N_14373,N_13772,N_13895);
or U14374 (N_14374,N_13673,N_13744);
and U14375 (N_14375,N_13777,N_13728);
nand U14376 (N_14376,N_13577,N_13721);
and U14377 (N_14377,N_13923,N_13918);
and U14378 (N_14378,N_13836,N_13843);
xnor U14379 (N_14379,N_13613,N_13636);
and U14380 (N_14380,N_13596,N_13900);
nand U14381 (N_14381,N_13714,N_13717);
nor U14382 (N_14382,N_13826,N_13553);
nor U14383 (N_14383,N_13510,N_13922);
and U14384 (N_14384,N_13900,N_13672);
xnor U14385 (N_14385,N_13629,N_13864);
xnor U14386 (N_14386,N_13598,N_13583);
or U14387 (N_14387,N_13639,N_13928);
nand U14388 (N_14388,N_13503,N_13903);
xor U14389 (N_14389,N_13560,N_13944);
xor U14390 (N_14390,N_13737,N_13734);
nor U14391 (N_14391,N_13883,N_13640);
and U14392 (N_14392,N_13516,N_13753);
nor U14393 (N_14393,N_13803,N_13717);
or U14394 (N_14394,N_13787,N_13831);
nand U14395 (N_14395,N_13619,N_13933);
xor U14396 (N_14396,N_13815,N_13929);
or U14397 (N_14397,N_13767,N_13847);
nor U14398 (N_14398,N_13919,N_13595);
nand U14399 (N_14399,N_13717,N_13703);
and U14400 (N_14400,N_13890,N_13617);
xnor U14401 (N_14401,N_13859,N_13637);
nand U14402 (N_14402,N_13561,N_13881);
nor U14403 (N_14403,N_13923,N_13825);
xnor U14404 (N_14404,N_13674,N_13908);
and U14405 (N_14405,N_13908,N_13648);
nand U14406 (N_14406,N_13631,N_13685);
nor U14407 (N_14407,N_13769,N_13669);
nand U14408 (N_14408,N_13504,N_13585);
and U14409 (N_14409,N_13748,N_13623);
or U14410 (N_14410,N_13979,N_13833);
nor U14411 (N_14411,N_13549,N_13655);
and U14412 (N_14412,N_13723,N_13689);
xor U14413 (N_14413,N_13698,N_13887);
nor U14414 (N_14414,N_13850,N_13792);
or U14415 (N_14415,N_13542,N_13668);
and U14416 (N_14416,N_13664,N_13654);
xnor U14417 (N_14417,N_13618,N_13982);
and U14418 (N_14418,N_13636,N_13863);
or U14419 (N_14419,N_13741,N_13508);
and U14420 (N_14420,N_13532,N_13826);
xnor U14421 (N_14421,N_13669,N_13793);
nand U14422 (N_14422,N_13530,N_13547);
and U14423 (N_14423,N_13826,N_13838);
or U14424 (N_14424,N_13645,N_13567);
nor U14425 (N_14425,N_13994,N_13645);
xnor U14426 (N_14426,N_13576,N_13732);
xor U14427 (N_14427,N_13752,N_13807);
nor U14428 (N_14428,N_13792,N_13743);
or U14429 (N_14429,N_13758,N_13895);
xor U14430 (N_14430,N_13824,N_13604);
or U14431 (N_14431,N_13931,N_13974);
or U14432 (N_14432,N_13510,N_13643);
xor U14433 (N_14433,N_13516,N_13771);
nor U14434 (N_14434,N_13646,N_13889);
xnor U14435 (N_14435,N_13771,N_13908);
or U14436 (N_14436,N_13801,N_13675);
nor U14437 (N_14437,N_13571,N_13905);
nor U14438 (N_14438,N_13979,N_13677);
nor U14439 (N_14439,N_13634,N_13549);
or U14440 (N_14440,N_13940,N_13761);
nand U14441 (N_14441,N_13927,N_13851);
nand U14442 (N_14442,N_13756,N_13620);
nand U14443 (N_14443,N_13870,N_13942);
xnor U14444 (N_14444,N_13505,N_13689);
and U14445 (N_14445,N_13716,N_13609);
or U14446 (N_14446,N_13814,N_13644);
nor U14447 (N_14447,N_13637,N_13579);
nand U14448 (N_14448,N_13873,N_13813);
and U14449 (N_14449,N_13786,N_13890);
xnor U14450 (N_14450,N_13605,N_13683);
and U14451 (N_14451,N_13660,N_13844);
or U14452 (N_14452,N_13737,N_13856);
and U14453 (N_14453,N_13595,N_13980);
xor U14454 (N_14454,N_13733,N_13575);
nor U14455 (N_14455,N_13761,N_13662);
and U14456 (N_14456,N_13519,N_13620);
and U14457 (N_14457,N_13959,N_13513);
and U14458 (N_14458,N_13911,N_13677);
xor U14459 (N_14459,N_13878,N_13999);
and U14460 (N_14460,N_13690,N_13711);
nor U14461 (N_14461,N_13508,N_13803);
nand U14462 (N_14462,N_13830,N_13885);
or U14463 (N_14463,N_13516,N_13592);
nor U14464 (N_14464,N_13671,N_13817);
and U14465 (N_14465,N_13862,N_13923);
or U14466 (N_14466,N_13897,N_13820);
nand U14467 (N_14467,N_13511,N_13828);
xnor U14468 (N_14468,N_13662,N_13994);
or U14469 (N_14469,N_13583,N_13767);
xor U14470 (N_14470,N_13890,N_13783);
xor U14471 (N_14471,N_13988,N_13769);
nand U14472 (N_14472,N_13966,N_13586);
nor U14473 (N_14473,N_13972,N_13997);
nor U14474 (N_14474,N_13708,N_13736);
and U14475 (N_14475,N_13657,N_13966);
nor U14476 (N_14476,N_13702,N_13793);
xnor U14477 (N_14477,N_13851,N_13538);
and U14478 (N_14478,N_13619,N_13996);
and U14479 (N_14479,N_13520,N_13701);
or U14480 (N_14480,N_13785,N_13809);
or U14481 (N_14481,N_13976,N_13767);
nor U14482 (N_14482,N_13514,N_13775);
xor U14483 (N_14483,N_13939,N_13937);
nor U14484 (N_14484,N_13530,N_13933);
or U14485 (N_14485,N_13508,N_13942);
or U14486 (N_14486,N_13595,N_13765);
nand U14487 (N_14487,N_13605,N_13906);
and U14488 (N_14488,N_13748,N_13536);
and U14489 (N_14489,N_13985,N_13545);
xor U14490 (N_14490,N_13948,N_13817);
nand U14491 (N_14491,N_13964,N_13503);
nand U14492 (N_14492,N_13972,N_13512);
nand U14493 (N_14493,N_13973,N_13938);
nor U14494 (N_14494,N_13990,N_13825);
and U14495 (N_14495,N_13943,N_13817);
or U14496 (N_14496,N_13814,N_13579);
nand U14497 (N_14497,N_13591,N_13512);
nor U14498 (N_14498,N_13999,N_13877);
nand U14499 (N_14499,N_13852,N_13769);
xnor U14500 (N_14500,N_14141,N_14113);
nor U14501 (N_14501,N_14204,N_14195);
xor U14502 (N_14502,N_14292,N_14360);
nand U14503 (N_14503,N_14110,N_14255);
and U14504 (N_14504,N_14092,N_14352);
xor U14505 (N_14505,N_14398,N_14216);
and U14506 (N_14506,N_14243,N_14032);
and U14507 (N_14507,N_14358,N_14024);
xor U14508 (N_14508,N_14453,N_14047);
nand U14509 (N_14509,N_14248,N_14397);
xor U14510 (N_14510,N_14326,N_14390);
nor U14511 (N_14511,N_14013,N_14038);
or U14512 (N_14512,N_14341,N_14134);
xor U14513 (N_14513,N_14062,N_14056);
or U14514 (N_14514,N_14048,N_14448);
or U14515 (N_14515,N_14432,N_14258);
nand U14516 (N_14516,N_14042,N_14021);
nand U14517 (N_14517,N_14452,N_14127);
xor U14518 (N_14518,N_14040,N_14321);
and U14519 (N_14519,N_14283,N_14100);
xor U14520 (N_14520,N_14218,N_14333);
nand U14521 (N_14521,N_14261,N_14329);
nand U14522 (N_14522,N_14193,N_14354);
xor U14523 (N_14523,N_14391,N_14147);
or U14524 (N_14524,N_14319,N_14177);
nor U14525 (N_14525,N_14137,N_14036);
nor U14526 (N_14526,N_14178,N_14249);
and U14527 (N_14527,N_14470,N_14473);
or U14528 (N_14528,N_14241,N_14280);
or U14529 (N_14529,N_14348,N_14488);
nand U14530 (N_14530,N_14288,N_14160);
or U14531 (N_14531,N_14157,N_14236);
nor U14532 (N_14532,N_14413,N_14079);
nand U14533 (N_14533,N_14221,N_14270);
xnor U14534 (N_14534,N_14217,N_14444);
or U14535 (N_14535,N_14422,N_14054);
and U14536 (N_14536,N_14230,N_14325);
nand U14537 (N_14537,N_14146,N_14463);
nor U14538 (N_14538,N_14046,N_14023);
nand U14539 (N_14539,N_14431,N_14388);
nor U14540 (N_14540,N_14439,N_14459);
or U14541 (N_14541,N_14359,N_14240);
or U14542 (N_14542,N_14294,N_14327);
nand U14543 (N_14543,N_14298,N_14440);
nand U14544 (N_14544,N_14392,N_14133);
nor U14545 (N_14545,N_14365,N_14231);
or U14546 (N_14546,N_14286,N_14197);
nor U14547 (N_14547,N_14315,N_14293);
or U14548 (N_14548,N_14428,N_14165);
xor U14549 (N_14549,N_14033,N_14139);
xor U14550 (N_14550,N_14183,N_14406);
xnor U14551 (N_14551,N_14020,N_14318);
nand U14552 (N_14552,N_14096,N_14087);
xnor U14553 (N_14553,N_14402,N_14170);
and U14554 (N_14554,N_14163,N_14244);
nand U14555 (N_14555,N_14269,N_14091);
nand U14556 (N_14556,N_14200,N_14136);
nand U14557 (N_14557,N_14161,N_14460);
xnor U14558 (N_14558,N_14214,N_14252);
xnor U14559 (N_14559,N_14469,N_14336);
and U14560 (N_14560,N_14149,N_14320);
xor U14561 (N_14561,N_14227,N_14371);
and U14562 (N_14562,N_14456,N_14167);
and U14563 (N_14563,N_14250,N_14380);
xnor U14564 (N_14564,N_14361,N_14089);
nand U14565 (N_14565,N_14454,N_14060);
or U14566 (N_14566,N_14407,N_14445);
or U14567 (N_14567,N_14260,N_14399);
and U14568 (N_14568,N_14052,N_14105);
nand U14569 (N_14569,N_14308,N_14458);
or U14570 (N_14570,N_14478,N_14190);
and U14571 (N_14571,N_14226,N_14345);
nand U14572 (N_14572,N_14233,N_14037);
nand U14573 (N_14573,N_14118,N_14065);
xor U14574 (N_14574,N_14187,N_14479);
nand U14575 (N_14575,N_14242,N_14404);
nand U14576 (N_14576,N_14486,N_14421);
nand U14577 (N_14577,N_14276,N_14061);
nand U14578 (N_14578,N_14259,N_14386);
nor U14579 (N_14579,N_14003,N_14279);
nand U14580 (N_14580,N_14184,N_14416);
and U14581 (N_14581,N_14420,N_14109);
nor U14582 (N_14582,N_14430,N_14115);
nor U14583 (N_14583,N_14011,N_14296);
nand U14584 (N_14584,N_14462,N_14316);
nand U14585 (N_14585,N_14309,N_14496);
and U14586 (N_14586,N_14499,N_14173);
nor U14587 (N_14587,N_14441,N_14271);
xor U14588 (N_14588,N_14497,N_14374);
xor U14589 (N_14589,N_14284,N_14369);
or U14590 (N_14590,N_14239,N_14495);
or U14591 (N_14591,N_14436,N_14073);
nand U14592 (N_14592,N_14395,N_14274);
or U14593 (N_14593,N_14289,N_14229);
nand U14594 (N_14594,N_14340,N_14384);
nor U14595 (N_14595,N_14050,N_14017);
and U14596 (N_14596,N_14306,N_14196);
nand U14597 (N_14597,N_14314,N_14313);
and U14598 (N_14598,N_14297,N_14211);
and U14599 (N_14599,N_14411,N_14121);
xor U14600 (N_14600,N_14034,N_14418);
xor U14601 (N_14601,N_14304,N_14475);
nand U14602 (N_14602,N_14375,N_14387);
and U14603 (N_14603,N_14245,N_14350);
and U14604 (N_14604,N_14049,N_14179);
xor U14605 (N_14605,N_14466,N_14433);
or U14606 (N_14606,N_14086,N_14142);
and U14607 (N_14607,N_14468,N_14031);
nand U14608 (N_14608,N_14373,N_14342);
nor U14609 (N_14609,N_14476,N_14349);
and U14610 (N_14610,N_14074,N_14045);
xor U14611 (N_14611,N_14467,N_14238);
xor U14612 (N_14612,N_14343,N_14188);
and U14613 (N_14613,N_14081,N_14180);
nor U14614 (N_14614,N_14265,N_14446);
nor U14615 (N_14615,N_14264,N_14176);
or U14616 (N_14616,N_14175,N_14493);
or U14617 (N_14617,N_14487,N_14078);
or U14618 (N_14618,N_14094,N_14353);
or U14619 (N_14619,N_14053,N_14266);
and U14620 (N_14620,N_14213,N_14155);
and U14621 (N_14621,N_14067,N_14267);
and U14622 (N_14622,N_14203,N_14080);
xor U14623 (N_14623,N_14123,N_14474);
or U14624 (N_14624,N_14041,N_14337);
and U14625 (N_14625,N_14158,N_14449);
xor U14626 (N_14626,N_14090,N_14290);
xor U14627 (N_14627,N_14205,N_14465);
xor U14628 (N_14628,N_14389,N_14135);
nand U14629 (N_14629,N_14098,N_14209);
and U14630 (N_14630,N_14104,N_14307);
and U14631 (N_14631,N_14299,N_14097);
and U14632 (N_14632,N_14103,N_14346);
or U14633 (N_14633,N_14206,N_14442);
and U14634 (N_14634,N_14084,N_14151);
nand U14635 (N_14635,N_14295,N_14044);
xor U14636 (N_14636,N_14077,N_14490);
nand U14637 (N_14637,N_14181,N_14172);
and U14638 (N_14638,N_14237,N_14491);
nand U14639 (N_14639,N_14351,N_14194);
and U14640 (N_14640,N_14379,N_14481);
or U14641 (N_14641,N_14156,N_14363);
or U14642 (N_14642,N_14117,N_14385);
and U14643 (N_14643,N_14370,N_14305);
nand U14644 (N_14644,N_14272,N_14372);
xnor U14645 (N_14645,N_14191,N_14364);
nor U14646 (N_14646,N_14095,N_14039);
xnor U14647 (N_14647,N_14185,N_14287);
nor U14648 (N_14648,N_14303,N_14107);
or U14649 (N_14649,N_14063,N_14059);
nand U14650 (N_14650,N_14251,N_14457);
nor U14651 (N_14651,N_14152,N_14192);
and U14652 (N_14652,N_14182,N_14247);
and U14653 (N_14653,N_14124,N_14403);
nor U14654 (N_14654,N_14401,N_14410);
xnor U14655 (N_14655,N_14235,N_14027);
nand U14656 (N_14656,N_14291,N_14168);
nor U14657 (N_14657,N_14256,N_14106);
nand U14658 (N_14658,N_14120,N_14008);
nor U14659 (N_14659,N_14064,N_14485);
nor U14660 (N_14660,N_14323,N_14016);
or U14661 (N_14661,N_14035,N_14408);
nand U14662 (N_14662,N_14394,N_14409);
and U14663 (N_14663,N_14451,N_14148);
nor U14664 (N_14664,N_14277,N_14143);
nor U14665 (N_14665,N_14331,N_14234);
xnor U14666 (N_14666,N_14128,N_14186);
or U14667 (N_14667,N_14189,N_14138);
nand U14668 (N_14668,N_14068,N_14414);
nand U14669 (N_14669,N_14026,N_14224);
nor U14670 (N_14670,N_14438,N_14246);
xnor U14671 (N_14671,N_14131,N_14419);
and U14672 (N_14672,N_14262,N_14014);
or U14673 (N_14673,N_14417,N_14119);
xor U14674 (N_14674,N_14332,N_14437);
nor U14675 (N_14675,N_14455,N_14057);
and U14676 (N_14676,N_14393,N_14482);
and U14677 (N_14677,N_14164,N_14085);
nand U14678 (N_14678,N_14066,N_14130);
xnor U14679 (N_14679,N_14344,N_14322);
and U14680 (N_14680,N_14076,N_14025);
xnor U14681 (N_14681,N_14001,N_14166);
or U14682 (N_14682,N_14015,N_14400);
xor U14683 (N_14683,N_14377,N_14043);
and U14684 (N_14684,N_14285,N_14132);
and U14685 (N_14685,N_14405,N_14144);
or U14686 (N_14686,N_14140,N_14254);
and U14687 (N_14687,N_14220,N_14415);
and U14688 (N_14688,N_14301,N_14302);
xnor U14689 (N_14689,N_14228,N_14162);
and U14690 (N_14690,N_14328,N_14088);
and U14691 (N_14691,N_14464,N_14169);
or U14692 (N_14692,N_14347,N_14268);
xor U14693 (N_14693,N_14232,N_14171);
and U14694 (N_14694,N_14202,N_14222);
or U14695 (N_14695,N_14219,N_14435);
xor U14696 (N_14696,N_14082,N_14126);
and U14697 (N_14697,N_14450,N_14311);
xor U14698 (N_14698,N_14075,N_14480);
or U14699 (N_14699,N_14434,N_14198);
nand U14700 (N_14700,N_14116,N_14423);
nand U14701 (N_14701,N_14030,N_14099);
and U14702 (N_14702,N_14355,N_14019);
nand U14703 (N_14703,N_14324,N_14275);
or U14704 (N_14704,N_14058,N_14199);
and U14705 (N_14705,N_14004,N_14207);
nor U14706 (N_14706,N_14472,N_14129);
or U14707 (N_14707,N_14029,N_14253);
nor U14708 (N_14708,N_14396,N_14125);
nand U14709 (N_14709,N_14257,N_14070);
or U14710 (N_14710,N_14083,N_14357);
nand U14711 (N_14711,N_14282,N_14006);
or U14712 (N_14712,N_14362,N_14483);
and U14713 (N_14713,N_14300,N_14071);
or U14714 (N_14714,N_14383,N_14212);
xnor U14715 (N_14715,N_14376,N_14102);
xnor U14716 (N_14716,N_14330,N_14278);
nand U14717 (N_14717,N_14339,N_14010);
nor U14718 (N_14718,N_14427,N_14012);
nand U14719 (N_14719,N_14215,N_14335);
xnor U14720 (N_14720,N_14471,N_14028);
nor U14721 (N_14721,N_14498,N_14201);
and U14722 (N_14722,N_14005,N_14111);
nor U14723 (N_14723,N_14145,N_14461);
or U14724 (N_14724,N_14174,N_14108);
and U14725 (N_14725,N_14273,N_14477);
or U14726 (N_14726,N_14263,N_14072);
nor U14727 (N_14727,N_14382,N_14007);
or U14728 (N_14728,N_14443,N_14069);
nor U14729 (N_14729,N_14424,N_14484);
or U14730 (N_14730,N_14009,N_14338);
or U14731 (N_14731,N_14114,N_14334);
xor U14732 (N_14732,N_14494,N_14159);
and U14733 (N_14733,N_14022,N_14366);
or U14734 (N_14734,N_14000,N_14381);
or U14735 (N_14735,N_14447,N_14093);
xor U14736 (N_14736,N_14150,N_14317);
nand U14737 (N_14737,N_14101,N_14281);
and U14738 (N_14738,N_14225,N_14368);
nand U14739 (N_14739,N_14112,N_14208);
nor U14740 (N_14740,N_14312,N_14367);
and U14741 (N_14741,N_14002,N_14122);
or U14742 (N_14742,N_14378,N_14425);
nor U14743 (N_14743,N_14210,N_14310);
xor U14744 (N_14744,N_14055,N_14492);
and U14745 (N_14745,N_14154,N_14356);
and U14746 (N_14746,N_14018,N_14489);
nand U14747 (N_14747,N_14153,N_14429);
and U14748 (N_14748,N_14223,N_14426);
nand U14749 (N_14749,N_14412,N_14051);
or U14750 (N_14750,N_14377,N_14387);
nor U14751 (N_14751,N_14076,N_14245);
nand U14752 (N_14752,N_14132,N_14417);
nand U14753 (N_14753,N_14033,N_14034);
xor U14754 (N_14754,N_14045,N_14068);
or U14755 (N_14755,N_14185,N_14418);
or U14756 (N_14756,N_14001,N_14470);
or U14757 (N_14757,N_14458,N_14482);
nand U14758 (N_14758,N_14052,N_14022);
nand U14759 (N_14759,N_14330,N_14021);
xor U14760 (N_14760,N_14449,N_14019);
or U14761 (N_14761,N_14094,N_14387);
xor U14762 (N_14762,N_14174,N_14020);
nor U14763 (N_14763,N_14011,N_14099);
and U14764 (N_14764,N_14304,N_14249);
or U14765 (N_14765,N_14053,N_14286);
and U14766 (N_14766,N_14375,N_14357);
nand U14767 (N_14767,N_14216,N_14195);
nand U14768 (N_14768,N_14345,N_14157);
or U14769 (N_14769,N_14248,N_14201);
nor U14770 (N_14770,N_14213,N_14425);
and U14771 (N_14771,N_14062,N_14495);
nand U14772 (N_14772,N_14367,N_14239);
and U14773 (N_14773,N_14331,N_14433);
nor U14774 (N_14774,N_14068,N_14336);
or U14775 (N_14775,N_14401,N_14258);
or U14776 (N_14776,N_14207,N_14157);
nor U14777 (N_14777,N_14073,N_14327);
nand U14778 (N_14778,N_14095,N_14393);
xnor U14779 (N_14779,N_14392,N_14352);
nor U14780 (N_14780,N_14076,N_14444);
and U14781 (N_14781,N_14122,N_14080);
nor U14782 (N_14782,N_14007,N_14204);
and U14783 (N_14783,N_14321,N_14083);
or U14784 (N_14784,N_14346,N_14069);
and U14785 (N_14785,N_14374,N_14368);
or U14786 (N_14786,N_14454,N_14336);
and U14787 (N_14787,N_14173,N_14250);
nor U14788 (N_14788,N_14073,N_14224);
xor U14789 (N_14789,N_14451,N_14388);
and U14790 (N_14790,N_14155,N_14401);
nand U14791 (N_14791,N_14061,N_14026);
and U14792 (N_14792,N_14288,N_14232);
nor U14793 (N_14793,N_14431,N_14217);
or U14794 (N_14794,N_14454,N_14437);
nand U14795 (N_14795,N_14219,N_14075);
nor U14796 (N_14796,N_14104,N_14369);
nand U14797 (N_14797,N_14335,N_14348);
or U14798 (N_14798,N_14432,N_14395);
nor U14799 (N_14799,N_14039,N_14379);
nand U14800 (N_14800,N_14206,N_14235);
nor U14801 (N_14801,N_14405,N_14019);
and U14802 (N_14802,N_14494,N_14246);
nor U14803 (N_14803,N_14242,N_14049);
nand U14804 (N_14804,N_14150,N_14490);
and U14805 (N_14805,N_14352,N_14045);
nand U14806 (N_14806,N_14218,N_14403);
nor U14807 (N_14807,N_14085,N_14100);
nand U14808 (N_14808,N_14160,N_14204);
xor U14809 (N_14809,N_14436,N_14225);
or U14810 (N_14810,N_14022,N_14347);
and U14811 (N_14811,N_14034,N_14064);
or U14812 (N_14812,N_14214,N_14465);
nand U14813 (N_14813,N_14204,N_14189);
xor U14814 (N_14814,N_14248,N_14088);
and U14815 (N_14815,N_14247,N_14251);
or U14816 (N_14816,N_14129,N_14399);
or U14817 (N_14817,N_14346,N_14024);
or U14818 (N_14818,N_14112,N_14243);
and U14819 (N_14819,N_14018,N_14329);
nand U14820 (N_14820,N_14358,N_14402);
or U14821 (N_14821,N_14138,N_14218);
nand U14822 (N_14822,N_14435,N_14475);
or U14823 (N_14823,N_14129,N_14471);
nand U14824 (N_14824,N_14006,N_14159);
or U14825 (N_14825,N_14410,N_14390);
nand U14826 (N_14826,N_14396,N_14372);
nor U14827 (N_14827,N_14300,N_14114);
or U14828 (N_14828,N_14301,N_14187);
or U14829 (N_14829,N_14484,N_14231);
and U14830 (N_14830,N_14457,N_14192);
and U14831 (N_14831,N_14401,N_14187);
xor U14832 (N_14832,N_14396,N_14036);
or U14833 (N_14833,N_14366,N_14310);
nor U14834 (N_14834,N_14249,N_14284);
and U14835 (N_14835,N_14170,N_14373);
and U14836 (N_14836,N_14223,N_14134);
or U14837 (N_14837,N_14362,N_14116);
and U14838 (N_14838,N_14121,N_14241);
nor U14839 (N_14839,N_14307,N_14396);
nand U14840 (N_14840,N_14182,N_14067);
nand U14841 (N_14841,N_14012,N_14489);
nand U14842 (N_14842,N_14169,N_14248);
or U14843 (N_14843,N_14240,N_14289);
nor U14844 (N_14844,N_14377,N_14204);
and U14845 (N_14845,N_14287,N_14079);
nand U14846 (N_14846,N_14085,N_14105);
xor U14847 (N_14847,N_14097,N_14295);
xnor U14848 (N_14848,N_14428,N_14064);
or U14849 (N_14849,N_14182,N_14344);
or U14850 (N_14850,N_14342,N_14444);
and U14851 (N_14851,N_14373,N_14135);
nand U14852 (N_14852,N_14086,N_14414);
nand U14853 (N_14853,N_14101,N_14035);
nand U14854 (N_14854,N_14487,N_14406);
or U14855 (N_14855,N_14008,N_14197);
nand U14856 (N_14856,N_14132,N_14299);
nor U14857 (N_14857,N_14088,N_14407);
nor U14858 (N_14858,N_14110,N_14185);
nand U14859 (N_14859,N_14199,N_14308);
xor U14860 (N_14860,N_14250,N_14112);
and U14861 (N_14861,N_14313,N_14017);
and U14862 (N_14862,N_14094,N_14135);
or U14863 (N_14863,N_14484,N_14373);
xnor U14864 (N_14864,N_14237,N_14142);
and U14865 (N_14865,N_14355,N_14039);
nand U14866 (N_14866,N_14209,N_14358);
nor U14867 (N_14867,N_14076,N_14366);
nor U14868 (N_14868,N_14074,N_14146);
nor U14869 (N_14869,N_14346,N_14065);
and U14870 (N_14870,N_14433,N_14131);
or U14871 (N_14871,N_14288,N_14213);
xor U14872 (N_14872,N_14114,N_14162);
or U14873 (N_14873,N_14132,N_14268);
nand U14874 (N_14874,N_14330,N_14200);
and U14875 (N_14875,N_14486,N_14042);
xor U14876 (N_14876,N_14046,N_14492);
or U14877 (N_14877,N_14292,N_14144);
nor U14878 (N_14878,N_14211,N_14320);
nand U14879 (N_14879,N_14237,N_14357);
nand U14880 (N_14880,N_14245,N_14125);
and U14881 (N_14881,N_14335,N_14270);
and U14882 (N_14882,N_14239,N_14135);
xnor U14883 (N_14883,N_14170,N_14455);
xor U14884 (N_14884,N_14265,N_14115);
xnor U14885 (N_14885,N_14045,N_14412);
xor U14886 (N_14886,N_14438,N_14235);
nor U14887 (N_14887,N_14376,N_14148);
or U14888 (N_14888,N_14357,N_14183);
and U14889 (N_14889,N_14094,N_14489);
nand U14890 (N_14890,N_14117,N_14424);
or U14891 (N_14891,N_14045,N_14470);
nand U14892 (N_14892,N_14076,N_14086);
xnor U14893 (N_14893,N_14051,N_14163);
xor U14894 (N_14894,N_14159,N_14328);
or U14895 (N_14895,N_14395,N_14125);
and U14896 (N_14896,N_14308,N_14201);
nand U14897 (N_14897,N_14137,N_14360);
or U14898 (N_14898,N_14288,N_14461);
nand U14899 (N_14899,N_14225,N_14162);
nand U14900 (N_14900,N_14062,N_14095);
and U14901 (N_14901,N_14135,N_14154);
and U14902 (N_14902,N_14223,N_14244);
or U14903 (N_14903,N_14461,N_14113);
nand U14904 (N_14904,N_14366,N_14323);
and U14905 (N_14905,N_14396,N_14404);
xnor U14906 (N_14906,N_14132,N_14201);
xor U14907 (N_14907,N_14108,N_14489);
nor U14908 (N_14908,N_14415,N_14410);
xnor U14909 (N_14909,N_14396,N_14017);
nor U14910 (N_14910,N_14261,N_14060);
nand U14911 (N_14911,N_14105,N_14444);
nand U14912 (N_14912,N_14118,N_14216);
nand U14913 (N_14913,N_14170,N_14312);
nor U14914 (N_14914,N_14133,N_14396);
and U14915 (N_14915,N_14280,N_14219);
or U14916 (N_14916,N_14368,N_14154);
nand U14917 (N_14917,N_14397,N_14234);
nor U14918 (N_14918,N_14351,N_14206);
nor U14919 (N_14919,N_14050,N_14125);
xnor U14920 (N_14920,N_14175,N_14146);
nor U14921 (N_14921,N_14247,N_14343);
and U14922 (N_14922,N_14116,N_14224);
xnor U14923 (N_14923,N_14384,N_14029);
xor U14924 (N_14924,N_14079,N_14195);
and U14925 (N_14925,N_14390,N_14474);
and U14926 (N_14926,N_14218,N_14413);
nand U14927 (N_14927,N_14108,N_14473);
nand U14928 (N_14928,N_14286,N_14300);
xor U14929 (N_14929,N_14189,N_14236);
nor U14930 (N_14930,N_14361,N_14135);
and U14931 (N_14931,N_14334,N_14411);
and U14932 (N_14932,N_14089,N_14486);
nand U14933 (N_14933,N_14438,N_14434);
and U14934 (N_14934,N_14065,N_14177);
or U14935 (N_14935,N_14484,N_14339);
or U14936 (N_14936,N_14397,N_14189);
xnor U14937 (N_14937,N_14324,N_14273);
xor U14938 (N_14938,N_14449,N_14298);
or U14939 (N_14939,N_14388,N_14154);
and U14940 (N_14940,N_14259,N_14280);
nand U14941 (N_14941,N_14313,N_14189);
or U14942 (N_14942,N_14082,N_14129);
nand U14943 (N_14943,N_14455,N_14358);
xor U14944 (N_14944,N_14315,N_14457);
nand U14945 (N_14945,N_14334,N_14167);
nand U14946 (N_14946,N_14134,N_14486);
xor U14947 (N_14947,N_14413,N_14431);
and U14948 (N_14948,N_14208,N_14374);
nor U14949 (N_14949,N_14436,N_14162);
xnor U14950 (N_14950,N_14376,N_14258);
and U14951 (N_14951,N_14161,N_14376);
and U14952 (N_14952,N_14378,N_14305);
and U14953 (N_14953,N_14318,N_14074);
and U14954 (N_14954,N_14142,N_14133);
nand U14955 (N_14955,N_14332,N_14091);
nor U14956 (N_14956,N_14035,N_14075);
xnor U14957 (N_14957,N_14108,N_14264);
nor U14958 (N_14958,N_14050,N_14448);
and U14959 (N_14959,N_14134,N_14209);
nor U14960 (N_14960,N_14395,N_14025);
and U14961 (N_14961,N_14040,N_14028);
nor U14962 (N_14962,N_14193,N_14319);
and U14963 (N_14963,N_14480,N_14346);
or U14964 (N_14964,N_14166,N_14374);
and U14965 (N_14965,N_14061,N_14250);
or U14966 (N_14966,N_14466,N_14489);
xnor U14967 (N_14967,N_14336,N_14126);
nor U14968 (N_14968,N_14158,N_14317);
nand U14969 (N_14969,N_14383,N_14265);
xor U14970 (N_14970,N_14289,N_14287);
nor U14971 (N_14971,N_14332,N_14472);
nor U14972 (N_14972,N_14308,N_14325);
nor U14973 (N_14973,N_14283,N_14309);
or U14974 (N_14974,N_14355,N_14342);
nand U14975 (N_14975,N_14372,N_14056);
xnor U14976 (N_14976,N_14270,N_14100);
or U14977 (N_14977,N_14384,N_14259);
or U14978 (N_14978,N_14204,N_14411);
xnor U14979 (N_14979,N_14386,N_14092);
and U14980 (N_14980,N_14010,N_14498);
nor U14981 (N_14981,N_14280,N_14167);
or U14982 (N_14982,N_14181,N_14330);
nand U14983 (N_14983,N_14228,N_14346);
or U14984 (N_14984,N_14198,N_14355);
xnor U14985 (N_14985,N_14032,N_14465);
xnor U14986 (N_14986,N_14448,N_14001);
nand U14987 (N_14987,N_14379,N_14080);
or U14988 (N_14988,N_14252,N_14037);
and U14989 (N_14989,N_14395,N_14392);
and U14990 (N_14990,N_14307,N_14442);
or U14991 (N_14991,N_14201,N_14330);
xnor U14992 (N_14992,N_14134,N_14427);
nand U14993 (N_14993,N_14105,N_14330);
and U14994 (N_14994,N_14152,N_14194);
nor U14995 (N_14995,N_14474,N_14156);
nor U14996 (N_14996,N_14083,N_14039);
nor U14997 (N_14997,N_14194,N_14288);
nor U14998 (N_14998,N_14400,N_14027);
nor U14999 (N_14999,N_14444,N_14408);
or U15000 (N_15000,N_14546,N_14761);
nor U15001 (N_15001,N_14783,N_14959);
xnor U15002 (N_15002,N_14826,N_14719);
xor U15003 (N_15003,N_14962,N_14507);
xnor U15004 (N_15004,N_14622,N_14846);
and U15005 (N_15005,N_14829,N_14948);
and U15006 (N_15006,N_14784,N_14729);
xor U15007 (N_15007,N_14712,N_14653);
and U15008 (N_15008,N_14926,N_14991);
or U15009 (N_15009,N_14640,N_14697);
or U15010 (N_15010,N_14616,N_14955);
and U15011 (N_15011,N_14654,N_14781);
nor U15012 (N_15012,N_14588,N_14828);
xnor U15013 (N_15013,N_14850,N_14540);
nor U15014 (N_15014,N_14755,N_14514);
nor U15015 (N_15015,N_14597,N_14513);
nor U15016 (N_15016,N_14964,N_14768);
and U15017 (N_15017,N_14522,N_14575);
and U15018 (N_15018,N_14883,N_14541);
xor U15019 (N_15019,N_14790,N_14786);
nor U15020 (N_15020,N_14657,N_14734);
xor U15021 (N_15021,N_14813,N_14780);
nand U15022 (N_15022,N_14680,N_14576);
xor U15023 (N_15023,N_14689,N_14635);
nor U15024 (N_15024,N_14714,N_14544);
xor U15025 (N_15025,N_14698,N_14905);
xor U15026 (N_15026,N_14767,N_14870);
and U15027 (N_15027,N_14830,N_14563);
and U15028 (N_15028,N_14531,N_14839);
and U15029 (N_15029,N_14766,N_14642);
xor U15030 (N_15030,N_14775,N_14695);
nand U15031 (N_15031,N_14778,N_14765);
nand U15032 (N_15032,N_14505,N_14973);
or U15033 (N_15033,N_14994,N_14532);
xnor U15034 (N_15034,N_14735,N_14951);
or U15035 (N_15035,N_14585,N_14848);
xor U15036 (N_15036,N_14679,N_14818);
nor U15037 (N_15037,N_14615,N_14884);
xnor U15038 (N_15038,N_14752,N_14983);
or U15039 (N_15039,N_14587,N_14675);
nand U15040 (N_15040,N_14992,N_14849);
xnor U15041 (N_15041,N_14866,N_14810);
nor U15042 (N_15042,N_14662,N_14750);
xnor U15043 (N_15043,N_14974,N_14791);
xnor U15044 (N_15044,N_14987,N_14935);
nand U15045 (N_15045,N_14692,N_14812);
and U15046 (N_15046,N_14677,N_14667);
nor U15047 (N_15047,N_14525,N_14627);
xor U15048 (N_15048,N_14931,N_14800);
nor U15049 (N_15049,N_14874,N_14669);
xnor U15050 (N_15050,N_14934,N_14868);
nor U15051 (N_15051,N_14979,N_14739);
xnor U15052 (N_15052,N_14872,N_14708);
and U15053 (N_15053,N_14763,N_14590);
or U15054 (N_15054,N_14998,N_14558);
nor U15055 (N_15055,N_14548,N_14877);
xnor U15056 (N_15056,N_14556,N_14799);
nor U15057 (N_15057,N_14710,N_14891);
nand U15058 (N_15058,N_14501,N_14553);
or U15059 (N_15059,N_14841,N_14996);
xor U15060 (N_15060,N_14727,N_14847);
xnor U15061 (N_15061,N_14936,N_14619);
or U15062 (N_15062,N_14878,N_14528);
and U15063 (N_15063,N_14612,N_14543);
nor U15064 (N_15064,N_14997,N_14875);
nor U15065 (N_15065,N_14795,N_14890);
xor U15066 (N_15066,N_14901,N_14625);
nand U15067 (N_15067,N_14820,N_14603);
or U15068 (N_15068,N_14777,N_14821);
xor U15069 (N_15069,N_14945,N_14937);
or U15070 (N_15070,N_14957,N_14571);
nor U15071 (N_15071,N_14764,N_14960);
xor U15072 (N_15072,N_14771,N_14534);
nor U15073 (N_15073,N_14980,N_14941);
nor U15074 (N_15074,N_14824,N_14794);
nor U15075 (N_15075,N_14745,N_14911);
or U15076 (N_15076,N_14977,N_14817);
nor U15077 (N_15077,N_14664,N_14854);
or U15078 (N_15078,N_14711,N_14740);
nor U15079 (N_15079,N_14920,N_14744);
xor U15080 (N_15080,N_14559,N_14939);
xor U15081 (N_15081,N_14871,N_14759);
or U15082 (N_15082,N_14632,N_14814);
and U15083 (N_15083,N_14753,N_14569);
and U15084 (N_15084,N_14516,N_14852);
nor U15085 (N_15085,N_14801,N_14678);
nor U15086 (N_15086,N_14628,N_14637);
nand U15087 (N_15087,N_14929,N_14726);
nor U15088 (N_15088,N_14730,N_14749);
or U15089 (N_15089,N_14614,N_14825);
xnor U15090 (N_15090,N_14545,N_14668);
nand U15091 (N_15091,N_14906,N_14895);
or U15092 (N_15092,N_14882,N_14972);
or U15093 (N_15093,N_14981,N_14990);
nor U15094 (N_15094,N_14646,N_14836);
and U15095 (N_15095,N_14943,N_14873);
nor U15096 (N_15096,N_14733,N_14721);
or U15097 (N_15097,N_14577,N_14834);
and U15098 (N_15098,N_14968,N_14963);
nor U15099 (N_15099,N_14647,N_14832);
or U15100 (N_15100,N_14944,N_14683);
or U15101 (N_15101,N_14725,N_14774);
and U15102 (N_15102,N_14928,N_14988);
and U15103 (N_15103,N_14584,N_14867);
or U15104 (N_15104,N_14518,N_14701);
nor U15105 (N_15105,N_14655,N_14517);
and U15106 (N_15106,N_14999,N_14737);
xnor U15107 (N_15107,N_14555,N_14819);
nand U15108 (N_15108,N_14658,N_14713);
and U15109 (N_15109,N_14731,N_14760);
or U15110 (N_15110,N_14904,N_14792);
or U15111 (N_15111,N_14530,N_14520);
nor U15112 (N_15112,N_14527,N_14924);
xor U15113 (N_15113,N_14881,N_14918);
xor U15114 (N_15114,N_14823,N_14596);
xnor U15115 (N_15115,N_14633,N_14512);
xnor U15116 (N_15116,N_14862,N_14652);
and U15117 (N_15117,N_14909,N_14676);
or U15118 (N_15118,N_14984,N_14703);
xnor U15119 (N_15119,N_14947,N_14912);
xor U15120 (N_15120,N_14706,N_14586);
nand U15121 (N_15121,N_14691,N_14978);
nor U15122 (N_15122,N_14788,N_14837);
or U15123 (N_15123,N_14644,N_14864);
and U15124 (N_15124,N_14693,N_14899);
xor U15125 (N_15125,N_14772,N_14853);
or U15126 (N_15126,N_14961,N_14938);
nand U15127 (N_15127,N_14670,N_14704);
xor U15128 (N_15128,N_14933,N_14521);
nor U15129 (N_15129,N_14705,N_14666);
nor U15130 (N_15130,N_14511,N_14844);
nand U15131 (N_15131,N_14609,N_14898);
nand U15132 (N_15132,N_14770,N_14568);
and U15133 (N_15133,N_14923,N_14797);
nand U15134 (N_15134,N_14958,N_14769);
xor U15135 (N_15135,N_14573,N_14807);
nor U15136 (N_15136,N_14827,N_14526);
xor U15137 (N_15137,N_14822,N_14932);
or U15138 (N_15138,N_14949,N_14842);
or U15139 (N_15139,N_14835,N_14631);
nand U15140 (N_15140,N_14804,N_14665);
and U15141 (N_15141,N_14723,N_14595);
or U15142 (N_15142,N_14551,N_14611);
and U15143 (N_15143,N_14629,N_14674);
nand U15144 (N_15144,N_14565,N_14536);
and U15145 (N_15145,N_14578,N_14741);
xor U15146 (N_15146,N_14634,N_14623);
nor U15147 (N_15147,N_14989,N_14894);
nor U15148 (N_15148,N_14694,N_14865);
nor U15149 (N_15149,N_14720,N_14715);
or U15150 (N_15150,N_14732,N_14581);
xor U15151 (N_15151,N_14716,N_14779);
and U15152 (N_15152,N_14681,N_14656);
or U15153 (N_15153,N_14940,N_14995);
or U15154 (N_15154,N_14684,N_14643);
or U15155 (N_15155,N_14902,N_14509);
nor U15156 (N_15156,N_14722,N_14638);
or U15157 (N_15157,N_14728,N_14965);
nand U15158 (N_15158,N_14976,N_14886);
xnor U15159 (N_15159,N_14682,N_14607);
nand U15160 (N_15160,N_14956,N_14855);
xor U15161 (N_15161,N_14639,N_14591);
or U15162 (N_15162,N_14688,N_14806);
and U15163 (N_15163,N_14896,N_14966);
and U15164 (N_15164,N_14952,N_14993);
nor U15165 (N_15165,N_14608,N_14748);
nand U15166 (N_15166,N_14773,N_14910);
and U15167 (N_15167,N_14925,N_14537);
xor U15168 (N_15168,N_14803,N_14885);
xor U15169 (N_15169,N_14523,N_14787);
and U15170 (N_15170,N_14907,N_14758);
xnor U15171 (N_15171,N_14808,N_14613);
nor U15172 (N_15172,N_14570,N_14802);
nand U15173 (N_15173,N_14547,N_14851);
or U15174 (N_15174,N_14641,N_14503);
xnor U15175 (N_15175,N_14542,N_14504);
or U15176 (N_15176,N_14580,N_14500);
and U15177 (N_15177,N_14809,N_14663);
or U15178 (N_15178,N_14592,N_14594);
nand U15179 (N_15179,N_14922,N_14967);
xnor U15180 (N_15180,N_14859,N_14696);
or U15181 (N_15181,N_14893,N_14970);
or U15182 (N_15182,N_14707,N_14897);
xnor U15183 (N_15183,N_14757,N_14747);
or U15184 (N_15184,N_14876,N_14687);
and U15185 (N_15185,N_14892,N_14650);
or U15186 (N_15186,N_14660,N_14811);
nand U15187 (N_15187,N_14927,N_14583);
xor U15188 (N_15188,N_14869,N_14510);
xnor U15189 (N_15189,N_14579,N_14900);
or U15190 (N_15190,N_14982,N_14599);
nand U15191 (N_15191,N_14702,N_14610);
and U15192 (N_15192,N_14672,N_14564);
nand U15193 (N_15193,N_14942,N_14582);
and U15194 (N_15194,N_14845,N_14557);
and U15195 (N_15195,N_14838,N_14756);
xor U15196 (N_15196,N_14954,N_14645);
or U15197 (N_15197,N_14524,N_14589);
xor U15198 (N_15198,N_14690,N_14562);
xnor U15199 (N_15199,N_14736,N_14879);
nand U15200 (N_15200,N_14574,N_14685);
or U15201 (N_15201,N_14550,N_14913);
nand U15202 (N_15202,N_14751,N_14843);
and U15203 (N_15203,N_14600,N_14782);
xor U15204 (N_15204,N_14502,N_14593);
nand U15205 (N_15205,N_14554,N_14975);
and U15206 (N_15206,N_14506,N_14796);
nor U15207 (N_15207,N_14598,N_14858);
or U15208 (N_15208,N_14986,N_14930);
nor U15209 (N_15209,N_14985,N_14626);
and U15210 (N_15210,N_14861,N_14601);
nand U15211 (N_15211,N_14617,N_14742);
or U15212 (N_15212,N_14789,N_14762);
nand U15213 (N_15213,N_14539,N_14857);
or U15214 (N_15214,N_14604,N_14648);
xnor U15215 (N_15215,N_14921,N_14620);
or U15216 (N_15216,N_14840,N_14671);
and U15217 (N_15217,N_14919,N_14880);
nand U15218 (N_15218,N_14673,N_14971);
xnor U15219 (N_15219,N_14953,N_14916);
nand U15220 (N_15220,N_14566,N_14793);
and U15221 (N_15221,N_14717,N_14572);
nand U15222 (N_15222,N_14561,N_14776);
or U15223 (N_15223,N_14567,N_14538);
xor U15224 (N_15224,N_14621,N_14950);
or U15225 (N_15225,N_14709,N_14917);
and U15226 (N_15226,N_14649,N_14606);
nor U15227 (N_15227,N_14815,N_14798);
nand U15228 (N_15228,N_14903,N_14831);
xor U15229 (N_15229,N_14915,N_14700);
xor U15230 (N_15230,N_14535,N_14908);
nor U15231 (N_15231,N_14533,N_14686);
nor U15232 (N_15232,N_14860,N_14661);
nand U15233 (N_15233,N_14888,N_14699);
nand U15234 (N_15234,N_14833,N_14508);
nand U15235 (N_15235,N_14946,N_14552);
and U15236 (N_15236,N_14914,N_14605);
nand U15237 (N_15237,N_14630,N_14863);
nor U15238 (N_15238,N_14659,N_14887);
or U15239 (N_15239,N_14856,N_14624);
nor U15240 (N_15240,N_14754,N_14718);
nor U15241 (N_15241,N_14651,N_14549);
nand U15242 (N_15242,N_14560,N_14805);
or U15243 (N_15243,N_14738,N_14969);
nor U15244 (N_15244,N_14618,N_14636);
or U15245 (N_15245,N_14515,N_14743);
xor U15246 (N_15246,N_14724,N_14816);
and U15247 (N_15247,N_14519,N_14602);
nand U15248 (N_15248,N_14529,N_14889);
or U15249 (N_15249,N_14746,N_14785);
nor U15250 (N_15250,N_14818,N_14799);
nand U15251 (N_15251,N_14570,N_14781);
xor U15252 (N_15252,N_14921,N_14834);
nand U15253 (N_15253,N_14973,N_14682);
or U15254 (N_15254,N_14647,N_14943);
and U15255 (N_15255,N_14557,N_14996);
nand U15256 (N_15256,N_14970,N_14676);
and U15257 (N_15257,N_14681,N_14664);
nor U15258 (N_15258,N_14940,N_14783);
or U15259 (N_15259,N_14847,N_14640);
and U15260 (N_15260,N_14789,N_14905);
xnor U15261 (N_15261,N_14876,N_14521);
xor U15262 (N_15262,N_14695,N_14983);
xor U15263 (N_15263,N_14942,N_14829);
or U15264 (N_15264,N_14890,N_14781);
nor U15265 (N_15265,N_14831,N_14953);
and U15266 (N_15266,N_14973,N_14997);
or U15267 (N_15267,N_14862,N_14734);
nor U15268 (N_15268,N_14999,N_14731);
nor U15269 (N_15269,N_14642,N_14629);
xnor U15270 (N_15270,N_14720,N_14659);
nand U15271 (N_15271,N_14778,N_14779);
xor U15272 (N_15272,N_14563,N_14625);
and U15273 (N_15273,N_14794,N_14882);
nand U15274 (N_15274,N_14803,N_14734);
xor U15275 (N_15275,N_14604,N_14630);
nor U15276 (N_15276,N_14936,N_14617);
nor U15277 (N_15277,N_14975,N_14815);
nor U15278 (N_15278,N_14904,N_14925);
nor U15279 (N_15279,N_14671,N_14707);
nand U15280 (N_15280,N_14651,N_14908);
nand U15281 (N_15281,N_14939,N_14710);
nor U15282 (N_15282,N_14878,N_14848);
xnor U15283 (N_15283,N_14605,N_14578);
nand U15284 (N_15284,N_14888,N_14590);
nand U15285 (N_15285,N_14912,N_14584);
or U15286 (N_15286,N_14818,N_14673);
and U15287 (N_15287,N_14508,N_14914);
or U15288 (N_15288,N_14699,N_14970);
xor U15289 (N_15289,N_14807,N_14780);
or U15290 (N_15290,N_14665,N_14988);
or U15291 (N_15291,N_14980,N_14706);
or U15292 (N_15292,N_14648,N_14909);
or U15293 (N_15293,N_14806,N_14647);
nor U15294 (N_15294,N_14807,N_14663);
xnor U15295 (N_15295,N_14933,N_14537);
or U15296 (N_15296,N_14689,N_14930);
or U15297 (N_15297,N_14788,N_14819);
and U15298 (N_15298,N_14971,N_14778);
nor U15299 (N_15299,N_14618,N_14584);
and U15300 (N_15300,N_14875,N_14669);
or U15301 (N_15301,N_14897,N_14513);
nand U15302 (N_15302,N_14915,N_14560);
nand U15303 (N_15303,N_14996,N_14851);
xor U15304 (N_15304,N_14925,N_14611);
or U15305 (N_15305,N_14623,N_14512);
nand U15306 (N_15306,N_14625,N_14742);
nor U15307 (N_15307,N_14874,N_14667);
or U15308 (N_15308,N_14884,N_14540);
and U15309 (N_15309,N_14598,N_14763);
nand U15310 (N_15310,N_14850,N_14520);
nor U15311 (N_15311,N_14802,N_14569);
and U15312 (N_15312,N_14846,N_14886);
and U15313 (N_15313,N_14775,N_14631);
xnor U15314 (N_15314,N_14701,N_14599);
xnor U15315 (N_15315,N_14538,N_14711);
xor U15316 (N_15316,N_14896,N_14774);
xnor U15317 (N_15317,N_14906,N_14604);
nor U15318 (N_15318,N_14679,N_14885);
nand U15319 (N_15319,N_14909,N_14710);
xnor U15320 (N_15320,N_14827,N_14609);
nand U15321 (N_15321,N_14944,N_14690);
xnor U15322 (N_15322,N_14989,N_14855);
nor U15323 (N_15323,N_14695,N_14589);
xor U15324 (N_15324,N_14851,N_14882);
nand U15325 (N_15325,N_14540,N_14956);
and U15326 (N_15326,N_14531,N_14741);
nand U15327 (N_15327,N_14728,N_14540);
or U15328 (N_15328,N_14962,N_14626);
nor U15329 (N_15329,N_14675,N_14663);
nand U15330 (N_15330,N_14993,N_14829);
or U15331 (N_15331,N_14738,N_14919);
or U15332 (N_15332,N_14548,N_14518);
nor U15333 (N_15333,N_14915,N_14707);
nor U15334 (N_15334,N_14878,N_14932);
and U15335 (N_15335,N_14686,N_14769);
and U15336 (N_15336,N_14819,N_14873);
or U15337 (N_15337,N_14865,N_14783);
or U15338 (N_15338,N_14992,N_14896);
xnor U15339 (N_15339,N_14957,N_14792);
and U15340 (N_15340,N_14746,N_14590);
nor U15341 (N_15341,N_14989,N_14629);
nand U15342 (N_15342,N_14880,N_14920);
xnor U15343 (N_15343,N_14687,N_14557);
and U15344 (N_15344,N_14927,N_14846);
and U15345 (N_15345,N_14657,N_14648);
or U15346 (N_15346,N_14789,N_14579);
xnor U15347 (N_15347,N_14600,N_14788);
xor U15348 (N_15348,N_14871,N_14751);
nand U15349 (N_15349,N_14790,N_14745);
xor U15350 (N_15350,N_14904,N_14811);
nor U15351 (N_15351,N_14509,N_14650);
nand U15352 (N_15352,N_14725,N_14505);
or U15353 (N_15353,N_14658,N_14722);
xnor U15354 (N_15354,N_14623,N_14603);
xnor U15355 (N_15355,N_14952,N_14992);
or U15356 (N_15356,N_14501,N_14613);
nor U15357 (N_15357,N_14666,N_14989);
nor U15358 (N_15358,N_14989,N_14509);
or U15359 (N_15359,N_14673,N_14908);
nor U15360 (N_15360,N_14533,N_14955);
and U15361 (N_15361,N_14537,N_14624);
nand U15362 (N_15362,N_14570,N_14964);
nand U15363 (N_15363,N_14888,N_14537);
or U15364 (N_15364,N_14993,N_14945);
and U15365 (N_15365,N_14634,N_14591);
or U15366 (N_15366,N_14922,N_14855);
xor U15367 (N_15367,N_14643,N_14650);
nand U15368 (N_15368,N_14994,N_14727);
nor U15369 (N_15369,N_14706,N_14503);
nor U15370 (N_15370,N_14932,N_14535);
nand U15371 (N_15371,N_14590,N_14643);
nor U15372 (N_15372,N_14948,N_14621);
nor U15373 (N_15373,N_14831,N_14793);
xor U15374 (N_15374,N_14660,N_14651);
or U15375 (N_15375,N_14967,N_14731);
nand U15376 (N_15376,N_14831,N_14517);
and U15377 (N_15377,N_14656,N_14852);
or U15378 (N_15378,N_14636,N_14985);
or U15379 (N_15379,N_14965,N_14817);
xor U15380 (N_15380,N_14500,N_14690);
or U15381 (N_15381,N_14593,N_14775);
xor U15382 (N_15382,N_14980,N_14648);
nand U15383 (N_15383,N_14757,N_14540);
and U15384 (N_15384,N_14654,N_14521);
nand U15385 (N_15385,N_14867,N_14841);
nand U15386 (N_15386,N_14811,N_14841);
nand U15387 (N_15387,N_14512,N_14866);
xor U15388 (N_15388,N_14974,N_14720);
or U15389 (N_15389,N_14708,N_14814);
nand U15390 (N_15390,N_14742,N_14511);
nand U15391 (N_15391,N_14595,N_14736);
nand U15392 (N_15392,N_14740,N_14802);
or U15393 (N_15393,N_14725,N_14783);
nor U15394 (N_15394,N_14509,N_14706);
and U15395 (N_15395,N_14959,N_14670);
nand U15396 (N_15396,N_14933,N_14622);
and U15397 (N_15397,N_14713,N_14686);
xnor U15398 (N_15398,N_14932,N_14904);
nor U15399 (N_15399,N_14708,N_14865);
and U15400 (N_15400,N_14620,N_14700);
and U15401 (N_15401,N_14916,N_14619);
and U15402 (N_15402,N_14830,N_14955);
and U15403 (N_15403,N_14573,N_14858);
and U15404 (N_15404,N_14855,N_14657);
nand U15405 (N_15405,N_14605,N_14504);
nor U15406 (N_15406,N_14518,N_14531);
nand U15407 (N_15407,N_14715,N_14989);
nand U15408 (N_15408,N_14984,N_14727);
or U15409 (N_15409,N_14780,N_14951);
and U15410 (N_15410,N_14540,N_14569);
xor U15411 (N_15411,N_14799,N_14976);
nand U15412 (N_15412,N_14801,N_14765);
or U15413 (N_15413,N_14843,N_14978);
nor U15414 (N_15414,N_14828,N_14637);
xor U15415 (N_15415,N_14954,N_14870);
nor U15416 (N_15416,N_14873,N_14902);
xnor U15417 (N_15417,N_14707,N_14883);
and U15418 (N_15418,N_14595,N_14845);
nor U15419 (N_15419,N_14816,N_14961);
and U15420 (N_15420,N_14996,N_14829);
or U15421 (N_15421,N_14791,N_14855);
or U15422 (N_15422,N_14683,N_14551);
nor U15423 (N_15423,N_14832,N_14954);
and U15424 (N_15424,N_14761,N_14506);
xor U15425 (N_15425,N_14983,N_14762);
or U15426 (N_15426,N_14898,N_14715);
nor U15427 (N_15427,N_14525,N_14925);
xnor U15428 (N_15428,N_14960,N_14580);
nand U15429 (N_15429,N_14966,N_14930);
nand U15430 (N_15430,N_14918,N_14506);
and U15431 (N_15431,N_14773,N_14581);
nor U15432 (N_15432,N_14820,N_14564);
xnor U15433 (N_15433,N_14800,N_14763);
nand U15434 (N_15434,N_14822,N_14976);
nand U15435 (N_15435,N_14587,N_14841);
nand U15436 (N_15436,N_14593,N_14931);
nand U15437 (N_15437,N_14995,N_14818);
or U15438 (N_15438,N_14950,N_14879);
nor U15439 (N_15439,N_14645,N_14710);
xor U15440 (N_15440,N_14713,N_14946);
or U15441 (N_15441,N_14855,N_14741);
or U15442 (N_15442,N_14871,N_14590);
nand U15443 (N_15443,N_14915,N_14903);
or U15444 (N_15444,N_14628,N_14560);
xnor U15445 (N_15445,N_14937,N_14646);
xnor U15446 (N_15446,N_14727,N_14539);
and U15447 (N_15447,N_14939,N_14823);
nor U15448 (N_15448,N_14530,N_14714);
nor U15449 (N_15449,N_14955,N_14683);
nor U15450 (N_15450,N_14622,N_14537);
and U15451 (N_15451,N_14880,N_14873);
nand U15452 (N_15452,N_14936,N_14853);
and U15453 (N_15453,N_14812,N_14993);
nand U15454 (N_15454,N_14731,N_14830);
and U15455 (N_15455,N_14570,N_14641);
or U15456 (N_15456,N_14910,N_14642);
or U15457 (N_15457,N_14606,N_14542);
nand U15458 (N_15458,N_14919,N_14978);
xor U15459 (N_15459,N_14692,N_14587);
and U15460 (N_15460,N_14880,N_14823);
nor U15461 (N_15461,N_14959,N_14726);
xnor U15462 (N_15462,N_14687,N_14717);
nor U15463 (N_15463,N_14717,N_14779);
nor U15464 (N_15464,N_14797,N_14832);
nand U15465 (N_15465,N_14685,N_14668);
nand U15466 (N_15466,N_14850,N_14806);
or U15467 (N_15467,N_14683,N_14735);
xor U15468 (N_15468,N_14684,N_14805);
xor U15469 (N_15469,N_14561,N_14902);
nor U15470 (N_15470,N_14665,N_14616);
xor U15471 (N_15471,N_14926,N_14533);
nor U15472 (N_15472,N_14853,N_14504);
xor U15473 (N_15473,N_14553,N_14610);
xnor U15474 (N_15474,N_14716,N_14839);
nand U15475 (N_15475,N_14567,N_14612);
or U15476 (N_15476,N_14820,N_14727);
nor U15477 (N_15477,N_14513,N_14914);
and U15478 (N_15478,N_14871,N_14677);
xnor U15479 (N_15479,N_14544,N_14974);
nand U15480 (N_15480,N_14547,N_14653);
or U15481 (N_15481,N_14585,N_14907);
or U15482 (N_15482,N_14830,N_14632);
and U15483 (N_15483,N_14989,N_14970);
and U15484 (N_15484,N_14647,N_14503);
nand U15485 (N_15485,N_14950,N_14798);
nor U15486 (N_15486,N_14793,N_14902);
nor U15487 (N_15487,N_14837,N_14955);
xnor U15488 (N_15488,N_14741,N_14541);
nor U15489 (N_15489,N_14930,N_14955);
nor U15490 (N_15490,N_14668,N_14544);
xor U15491 (N_15491,N_14743,N_14994);
and U15492 (N_15492,N_14600,N_14591);
or U15493 (N_15493,N_14680,N_14586);
nor U15494 (N_15494,N_14605,N_14895);
xnor U15495 (N_15495,N_14581,N_14657);
xor U15496 (N_15496,N_14589,N_14885);
nand U15497 (N_15497,N_14712,N_14742);
nand U15498 (N_15498,N_14992,N_14760);
xor U15499 (N_15499,N_14878,N_14642);
and U15500 (N_15500,N_15076,N_15129);
xor U15501 (N_15501,N_15072,N_15061);
nand U15502 (N_15502,N_15402,N_15048);
nor U15503 (N_15503,N_15465,N_15185);
xnor U15504 (N_15504,N_15307,N_15496);
xor U15505 (N_15505,N_15386,N_15232);
or U15506 (N_15506,N_15454,N_15257);
xnor U15507 (N_15507,N_15371,N_15338);
and U15508 (N_15508,N_15119,N_15489);
nand U15509 (N_15509,N_15351,N_15008);
xor U15510 (N_15510,N_15494,N_15152);
nand U15511 (N_15511,N_15258,N_15054);
and U15512 (N_15512,N_15175,N_15233);
and U15513 (N_15513,N_15222,N_15144);
nand U15514 (N_15514,N_15192,N_15332);
xor U15515 (N_15515,N_15116,N_15378);
and U15516 (N_15516,N_15039,N_15177);
nand U15517 (N_15517,N_15238,N_15323);
nor U15518 (N_15518,N_15309,N_15486);
or U15519 (N_15519,N_15182,N_15028);
nor U15520 (N_15520,N_15423,N_15255);
or U15521 (N_15521,N_15349,N_15477);
nor U15522 (N_15522,N_15377,N_15388);
nand U15523 (N_15523,N_15020,N_15416);
nor U15524 (N_15524,N_15073,N_15108);
or U15525 (N_15525,N_15140,N_15114);
nor U15526 (N_15526,N_15223,N_15479);
and U15527 (N_15527,N_15139,N_15480);
xnor U15528 (N_15528,N_15414,N_15424);
xor U15529 (N_15529,N_15069,N_15264);
or U15530 (N_15530,N_15207,N_15126);
nand U15531 (N_15531,N_15085,N_15246);
or U15532 (N_15532,N_15447,N_15154);
nor U15533 (N_15533,N_15426,N_15195);
xnor U15534 (N_15534,N_15280,N_15149);
nand U15535 (N_15535,N_15304,N_15273);
xnor U15536 (N_15536,N_15317,N_15023);
or U15537 (N_15537,N_15103,N_15147);
and U15538 (N_15538,N_15049,N_15375);
and U15539 (N_15539,N_15292,N_15363);
or U15540 (N_15540,N_15176,N_15164);
xor U15541 (N_15541,N_15014,N_15310);
and U15542 (N_15542,N_15427,N_15191);
or U15543 (N_15543,N_15247,N_15383);
nand U15544 (N_15544,N_15022,N_15219);
xor U15545 (N_15545,N_15201,N_15253);
nand U15546 (N_15546,N_15090,N_15422);
or U15547 (N_15547,N_15336,N_15256);
nand U15548 (N_15548,N_15325,N_15180);
and U15549 (N_15549,N_15318,N_15074);
and U15550 (N_15550,N_15391,N_15466);
xor U15551 (N_15551,N_15269,N_15131);
nand U15552 (N_15552,N_15044,N_15112);
or U15553 (N_15553,N_15237,N_15458);
nand U15554 (N_15554,N_15339,N_15240);
nand U15555 (N_15555,N_15184,N_15409);
nand U15556 (N_15556,N_15497,N_15208);
nand U15557 (N_15557,N_15032,N_15010);
nand U15558 (N_15558,N_15300,N_15059);
xor U15559 (N_15559,N_15369,N_15230);
or U15560 (N_15560,N_15060,N_15155);
and U15561 (N_15561,N_15354,N_15102);
nor U15562 (N_15562,N_15346,N_15437);
xor U15563 (N_15563,N_15083,N_15367);
xnor U15564 (N_15564,N_15202,N_15215);
and U15565 (N_15565,N_15158,N_15289);
nand U15566 (N_15566,N_15097,N_15428);
nor U15567 (N_15567,N_15006,N_15401);
nor U15568 (N_15568,N_15334,N_15009);
nor U15569 (N_15569,N_15487,N_15231);
nor U15570 (N_15570,N_15450,N_15050);
xor U15571 (N_15571,N_15400,N_15308);
and U15572 (N_15572,N_15294,N_15104);
xnor U15573 (N_15573,N_15056,N_15355);
xnor U15574 (N_15574,N_15299,N_15169);
nor U15575 (N_15575,N_15322,N_15092);
nand U15576 (N_15576,N_15021,N_15098);
nand U15577 (N_15577,N_15071,N_15019);
or U15578 (N_15578,N_15214,N_15384);
and U15579 (N_15579,N_15088,N_15221);
and U15580 (N_15580,N_15080,N_15467);
nor U15581 (N_15581,N_15261,N_15045);
or U15582 (N_15582,N_15365,N_15203);
and U15583 (N_15583,N_15065,N_15151);
nor U15584 (N_15584,N_15474,N_15041);
nand U15585 (N_15585,N_15243,N_15123);
or U15586 (N_15586,N_15319,N_15209);
nor U15587 (N_15587,N_15418,N_15431);
and U15588 (N_15588,N_15373,N_15348);
or U15589 (N_15589,N_15341,N_15493);
nand U15590 (N_15590,N_15315,N_15031);
xor U15591 (N_15591,N_15482,N_15347);
nor U15592 (N_15592,N_15120,N_15381);
nand U15593 (N_15593,N_15360,N_15271);
xnor U15594 (N_15594,N_15012,N_15143);
nor U15595 (N_15595,N_15456,N_15239);
xor U15596 (N_15596,N_15078,N_15326);
xor U15597 (N_15597,N_15011,N_15089);
nor U15598 (N_15598,N_15166,N_15093);
nor U15599 (N_15599,N_15435,N_15473);
xor U15600 (N_15600,N_15033,N_15190);
nand U15601 (N_15601,N_15035,N_15274);
nor U15602 (N_15602,N_15262,N_15263);
and U15603 (N_15603,N_15141,N_15130);
nor U15604 (N_15604,N_15359,N_15138);
xnor U15605 (N_15605,N_15082,N_15016);
and U15606 (N_15606,N_15442,N_15109);
and U15607 (N_15607,N_15267,N_15121);
nand U15608 (N_15608,N_15254,N_15070);
nand U15609 (N_15609,N_15291,N_15469);
nand U15610 (N_15610,N_15382,N_15042);
xnor U15611 (N_15611,N_15026,N_15063);
nand U15612 (N_15612,N_15249,N_15029);
or U15613 (N_15613,N_15217,N_15106);
and U15614 (N_15614,N_15034,N_15079);
nor U15615 (N_15615,N_15245,N_15444);
nand U15616 (N_15616,N_15405,N_15040);
or U15617 (N_15617,N_15296,N_15398);
or U15618 (N_15618,N_15441,N_15000);
or U15619 (N_15619,N_15173,N_15210);
nor U15620 (N_15620,N_15134,N_15174);
or U15621 (N_15621,N_15260,N_15235);
xnor U15622 (N_15622,N_15314,N_15087);
and U15623 (N_15623,N_15410,N_15394);
nor U15624 (N_15624,N_15358,N_15186);
nand U15625 (N_15625,N_15027,N_15146);
nand U15626 (N_15626,N_15024,N_15091);
nor U15627 (N_15627,N_15161,N_15178);
and U15628 (N_15628,N_15259,N_15290);
and U15629 (N_15629,N_15110,N_15077);
or U15630 (N_15630,N_15013,N_15204);
nor U15631 (N_15631,N_15100,N_15286);
and U15632 (N_15632,N_15471,N_15446);
nand U15633 (N_15633,N_15196,N_15227);
nand U15634 (N_15634,N_15297,N_15162);
nor U15635 (N_15635,N_15099,N_15302);
and U15636 (N_15636,N_15086,N_15443);
and U15637 (N_15637,N_15241,N_15283);
nor U15638 (N_15638,N_15328,N_15150);
and U15639 (N_15639,N_15018,N_15420);
xnor U15640 (N_15640,N_15462,N_15313);
or U15641 (N_15641,N_15419,N_15067);
nor U15642 (N_15642,N_15094,N_15293);
or U15643 (N_15643,N_15403,N_15156);
nor U15644 (N_15644,N_15372,N_15081);
nand U15645 (N_15645,N_15179,N_15183);
and U15646 (N_15646,N_15392,N_15281);
nand U15647 (N_15647,N_15007,N_15331);
and U15648 (N_15648,N_15492,N_15408);
nor U15649 (N_15649,N_15193,N_15376);
nand U15650 (N_15650,N_15270,N_15498);
and U15651 (N_15651,N_15395,N_15213);
nand U15652 (N_15652,N_15451,N_15003);
nor U15653 (N_15653,N_15288,N_15357);
or U15654 (N_15654,N_15449,N_15117);
nand U15655 (N_15655,N_15320,N_15189);
nor U15656 (N_15656,N_15198,N_15368);
and U15657 (N_15657,N_15415,N_15481);
nand U15658 (N_15658,N_15285,N_15224);
and U15659 (N_15659,N_15335,N_15188);
xnor U15660 (N_15660,N_15374,N_15350);
nor U15661 (N_15661,N_15301,N_15390);
nor U15662 (N_15662,N_15490,N_15345);
and U15663 (N_15663,N_15036,N_15316);
and U15664 (N_15664,N_15275,N_15046);
and U15665 (N_15665,N_15062,N_15251);
or U15666 (N_15666,N_15366,N_15413);
and U15667 (N_15667,N_15311,N_15167);
nor U15668 (N_15668,N_15340,N_15160);
nand U15669 (N_15669,N_15303,N_15153);
or U15670 (N_15670,N_15057,N_15284);
xor U15671 (N_15671,N_15132,N_15439);
and U15672 (N_15672,N_15172,N_15084);
xor U15673 (N_15673,N_15266,N_15252);
nand U15674 (N_15674,N_15242,N_15043);
nor U15675 (N_15675,N_15133,N_15030);
and U15676 (N_15676,N_15157,N_15187);
nor U15677 (N_15677,N_15485,N_15344);
xnor U15678 (N_15678,N_15200,N_15206);
or U15679 (N_15679,N_15495,N_15298);
xnor U15680 (N_15680,N_15272,N_15244);
nand U15681 (N_15681,N_15148,N_15370);
nand U15682 (N_15682,N_15434,N_15137);
nand U15683 (N_15683,N_15453,N_15197);
or U15684 (N_15684,N_15225,N_15017);
nor U15685 (N_15685,N_15330,N_15096);
nor U15686 (N_15686,N_15005,N_15181);
or U15687 (N_15687,N_15379,N_15279);
nand U15688 (N_15688,N_15124,N_15324);
or U15689 (N_15689,N_15432,N_15216);
nor U15690 (N_15690,N_15250,N_15066);
nand U15691 (N_15691,N_15075,N_15407);
and U15692 (N_15692,N_15228,N_15356);
and U15693 (N_15693,N_15128,N_15455);
and U15694 (N_15694,N_15364,N_15004);
or U15695 (N_15695,N_15025,N_15305);
or U15696 (N_15696,N_15476,N_15306);
or U15697 (N_15697,N_15058,N_15385);
or U15698 (N_15698,N_15361,N_15135);
and U15699 (N_15699,N_15165,N_15047);
nand U15700 (N_15700,N_15464,N_15429);
or U15701 (N_15701,N_15145,N_15276);
nor U15702 (N_15702,N_15127,N_15282);
xnor U15703 (N_15703,N_15488,N_15115);
nand U15704 (N_15704,N_15052,N_15268);
or U15705 (N_15705,N_15312,N_15105);
xor U15706 (N_15706,N_15122,N_15101);
nand U15707 (N_15707,N_15461,N_15142);
nor U15708 (N_15708,N_15037,N_15470);
xor U15709 (N_15709,N_15265,N_15362);
xor U15710 (N_15710,N_15107,N_15448);
and U15711 (N_15711,N_15211,N_15387);
or U15712 (N_15712,N_15352,N_15171);
and U15713 (N_15713,N_15287,N_15499);
and U15714 (N_15714,N_15353,N_15220);
xnor U15715 (N_15715,N_15295,N_15438);
xor U15716 (N_15716,N_15218,N_15459);
nor U15717 (N_15717,N_15001,N_15484);
or U15718 (N_15718,N_15053,N_15472);
nand U15719 (N_15719,N_15248,N_15068);
and U15720 (N_15720,N_15229,N_15343);
or U15721 (N_15721,N_15321,N_15329);
and U15722 (N_15722,N_15404,N_15095);
or U15723 (N_15723,N_15212,N_15337);
or U15724 (N_15724,N_15170,N_15194);
nor U15725 (N_15725,N_15445,N_15412);
nand U15726 (N_15726,N_15118,N_15342);
nor U15727 (N_15727,N_15475,N_15421);
nor U15728 (N_15728,N_15430,N_15436);
and U15729 (N_15729,N_15051,N_15064);
and U15730 (N_15730,N_15389,N_15483);
xor U15731 (N_15731,N_15277,N_15168);
and U15732 (N_15732,N_15136,N_15397);
nor U15733 (N_15733,N_15411,N_15205);
nor U15734 (N_15734,N_15111,N_15396);
xor U15735 (N_15735,N_15425,N_15038);
xor U15736 (N_15736,N_15491,N_15159);
xnor U15737 (N_15737,N_15399,N_15327);
nand U15738 (N_15738,N_15015,N_15226);
xnor U15739 (N_15739,N_15055,N_15234);
nor U15740 (N_15740,N_15333,N_15478);
xor U15741 (N_15741,N_15457,N_15278);
and U15742 (N_15742,N_15417,N_15406);
xor U15743 (N_15743,N_15433,N_15463);
nor U15744 (N_15744,N_15125,N_15452);
and U15745 (N_15745,N_15163,N_15113);
or U15746 (N_15746,N_15380,N_15440);
and U15747 (N_15747,N_15460,N_15236);
nor U15748 (N_15748,N_15468,N_15002);
xnor U15749 (N_15749,N_15393,N_15199);
and U15750 (N_15750,N_15158,N_15199);
nor U15751 (N_15751,N_15055,N_15238);
or U15752 (N_15752,N_15034,N_15409);
or U15753 (N_15753,N_15307,N_15017);
nand U15754 (N_15754,N_15081,N_15289);
or U15755 (N_15755,N_15282,N_15372);
nor U15756 (N_15756,N_15480,N_15331);
or U15757 (N_15757,N_15345,N_15059);
nand U15758 (N_15758,N_15054,N_15310);
xnor U15759 (N_15759,N_15422,N_15322);
nor U15760 (N_15760,N_15364,N_15220);
xnor U15761 (N_15761,N_15010,N_15046);
xor U15762 (N_15762,N_15435,N_15126);
and U15763 (N_15763,N_15426,N_15368);
xor U15764 (N_15764,N_15005,N_15328);
nand U15765 (N_15765,N_15004,N_15162);
nand U15766 (N_15766,N_15316,N_15302);
nor U15767 (N_15767,N_15403,N_15400);
and U15768 (N_15768,N_15460,N_15380);
or U15769 (N_15769,N_15394,N_15275);
and U15770 (N_15770,N_15195,N_15193);
nand U15771 (N_15771,N_15058,N_15125);
nand U15772 (N_15772,N_15161,N_15014);
nand U15773 (N_15773,N_15273,N_15060);
or U15774 (N_15774,N_15093,N_15286);
or U15775 (N_15775,N_15223,N_15286);
xnor U15776 (N_15776,N_15240,N_15138);
and U15777 (N_15777,N_15391,N_15018);
nor U15778 (N_15778,N_15101,N_15459);
nand U15779 (N_15779,N_15116,N_15250);
or U15780 (N_15780,N_15244,N_15415);
nand U15781 (N_15781,N_15475,N_15297);
nand U15782 (N_15782,N_15072,N_15388);
nand U15783 (N_15783,N_15134,N_15026);
or U15784 (N_15784,N_15075,N_15039);
xor U15785 (N_15785,N_15117,N_15208);
nand U15786 (N_15786,N_15270,N_15211);
and U15787 (N_15787,N_15127,N_15073);
nor U15788 (N_15788,N_15155,N_15071);
and U15789 (N_15789,N_15035,N_15127);
xor U15790 (N_15790,N_15386,N_15396);
or U15791 (N_15791,N_15309,N_15223);
nand U15792 (N_15792,N_15475,N_15273);
and U15793 (N_15793,N_15070,N_15393);
nand U15794 (N_15794,N_15179,N_15038);
and U15795 (N_15795,N_15007,N_15147);
and U15796 (N_15796,N_15373,N_15468);
xor U15797 (N_15797,N_15456,N_15193);
nand U15798 (N_15798,N_15089,N_15457);
nand U15799 (N_15799,N_15163,N_15304);
and U15800 (N_15800,N_15309,N_15472);
nor U15801 (N_15801,N_15423,N_15072);
nand U15802 (N_15802,N_15463,N_15259);
nor U15803 (N_15803,N_15188,N_15223);
or U15804 (N_15804,N_15123,N_15460);
and U15805 (N_15805,N_15224,N_15434);
xnor U15806 (N_15806,N_15089,N_15260);
xor U15807 (N_15807,N_15314,N_15208);
xor U15808 (N_15808,N_15460,N_15108);
xnor U15809 (N_15809,N_15438,N_15255);
or U15810 (N_15810,N_15236,N_15061);
or U15811 (N_15811,N_15426,N_15465);
nor U15812 (N_15812,N_15382,N_15080);
nand U15813 (N_15813,N_15366,N_15374);
or U15814 (N_15814,N_15370,N_15407);
xnor U15815 (N_15815,N_15099,N_15207);
nand U15816 (N_15816,N_15181,N_15411);
nand U15817 (N_15817,N_15151,N_15073);
xor U15818 (N_15818,N_15135,N_15080);
xnor U15819 (N_15819,N_15095,N_15067);
nand U15820 (N_15820,N_15359,N_15432);
and U15821 (N_15821,N_15080,N_15359);
or U15822 (N_15822,N_15299,N_15309);
xor U15823 (N_15823,N_15453,N_15360);
and U15824 (N_15824,N_15167,N_15269);
or U15825 (N_15825,N_15020,N_15240);
xnor U15826 (N_15826,N_15324,N_15204);
and U15827 (N_15827,N_15133,N_15124);
nor U15828 (N_15828,N_15422,N_15269);
nand U15829 (N_15829,N_15382,N_15490);
nand U15830 (N_15830,N_15166,N_15102);
and U15831 (N_15831,N_15044,N_15273);
and U15832 (N_15832,N_15395,N_15185);
xor U15833 (N_15833,N_15279,N_15488);
xor U15834 (N_15834,N_15010,N_15184);
xnor U15835 (N_15835,N_15427,N_15063);
xor U15836 (N_15836,N_15167,N_15372);
nand U15837 (N_15837,N_15352,N_15241);
nor U15838 (N_15838,N_15428,N_15315);
nor U15839 (N_15839,N_15127,N_15498);
xor U15840 (N_15840,N_15287,N_15441);
and U15841 (N_15841,N_15295,N_15427);
or U15842 (N_15842,N_15286,N_15004);
xor U15843 (N_15843,N_15007,N_15392);
and U15844 (N_15844,N_15237,N_15343);
nand U15845 (N_15845,N_15265,N_15316);
xor U15846 (N_15846,N_15269,N_15183);
and U15847 (N_15847,N_15348,N_15050);
nor U15848 (N_15848,N_15343,N_15083);
nand U15849 (N_15849,N_15030,N_15457);
nor U15850 (N_15850,N_15035,N_15394);
or U15851 (N_15851,N_15162,N_15308);
nand U15852 (N_15852,N_15298,N_15004);
or U15853 (N_15853,N_15131,N_15456);
nand U15854 (N_15854,N_15060,N_15438);
xnor U15855 (N_15855,N_15327,N_15201);
nor U15856 (N_15856,N_15032,N_15140);
nand U15857 (N_15857,N_15197,N_15095);
xor U15858 (N_15858,N_15224,N_15362);
nand U15859 (N_15859,N_15326,N_15010);
nand U15860 (N_15860,N_15017,N_15324);
or U15861 (N_15861,N_15213,N_15238);
nor U15862 (N_15862,N_15312,N_15484);
xor U15863 (N_15863,N_15422,N_15414);
and U15864 (N_15864,N_15401,N_15121);
nor U15865 (N_15865,N_15406,N_15173);
nand U15866 (N_15866,N_15251,N_15127);
nand U15867 (N_15867,N_15080,N_15041);
nor U15868 (N_15868,N_15325,N_15132);
xor U15869 (N_15869,N_15390,N_15089);
or U15870 (N_15870,N_15386,N_15440);
nor U15871 (N_15871,N_15002,N_15457);
nor U15872 (N_15872,N_15358,N_15241);
nand U15873 (N_15873,N_15248,N_15106);
xor U15874 (N_15874,N_15271,N_15186);
xnor U15875 (N_15875,N_15026,N_15013);
nand U15876 (N_15876,N_15394,N_15190);
xor U15877 (N_15877,N_15082,N_15194);
or U15878 (N_15878,N_15012,N_15010);
nor U15879 (N_15879,N_15310,N_15023);
nand U15880 (N_15880,N_15217,N_15005);
nand U15881 (N_15881,N_15059,N_15458);
or U15882 (N_15882,N_15367,N_15044);
or U15883 (N_15883,N_15088,N_15334);
and U15884 (N_15884,N_15207,N_15003);
xor U15885 (N_15885,N_15354,N_15334);
or U15886 (N_15886,N_15432,N_15237);
nand U15887 (N_15887,N_15062,N_15441);
or U15888 (N_15888,N_15272,N_15408);
nand U15889 (N_15889,N_15269,N_15001);
nand U15890 (N_15890,N_15458,N_15304);
nor U15891 (N_15891,N_15093,N_15285);
nand U15892 (N_15892,N_15099,N_15268);
nand U15893 (N_15893,N_15273,N_15293);
nand U15894 (N_15894,N_15150,N_15093);
xnor U15895 (N_15895,N_15418,N_15407);
nand U15896 (N_15896,N_15104,N_15159);
nand U15897 (N_15897,N_15233,N_15251);
or U15898 (N_15898,N_15206,N_15464);
and U15899 (N_15899,N_15108,N_15240);
nor U15900 (N_15900,N_15387,N_15402);
or U15901 (N_15901,N_15077,N_15411);
xor U15902 (N_15902,N_15093,N_15066);
and U15903 (N_15903,N_15214,N_15402);
and U15904 (N_15904,N_15445,N_15284);
nand U15905 (N_15905,N_15443,N_15474);
xor U15906 (N_15906,N_15132,N_15011);
xnor U15907 (N_15907,N_15389,N_15180);
xnor U15908 (N_15908,N_15493,N_15116);
xor U15909 (N_15909,N_15001,N_15434);
xnor U15910 (N_15910,N_15371,N_15327);
and U15911 (N_15911,N_15041,N_15208);
nand U15912 (N_15912,N_15259,N_15044);
xnor U15913 (N_15913,N_15308,N_15337);
nand U15914 (N_15914,N_15208,N_15076);
nor U15915 (N_15915,N_15352,N_15278);
or U15916 (N_15916,N_15287,N_15214);
and U15917 (N_15917,N_15287,N_15164);
nor U15918 (N_15918,N_15122,N_15212);
nor U15919 (N_15919,N_15179,N_15012);
nand U15920 (N_15920,N_15385,N_15027);
and U15921 (N_15921,N_15353,N_15125);
nand U15922 (N_15922,N_15317,N_15302);
and U15923 (N_15923,N_15413,N_15409);
nand U15924 (N_15924,N_15472,N_15240);
nor U15925 (N_15925,N_15429,N_15058);
xor U15926 (N_15926,N_15389,N_15187);
or U15927 (N_15927,N_15185,N_15075);
nand U15928 (N_15928,N_15494,N_15353);
nor U15929 (N_15929,N_15465,N_15119);
xnor U15930 (N_15930,N_15105,N_15475);
nor U15931 (N_15931,N_15071,N_15166);
nor U15932 (N_15932,N_15466,N_15197);
or U15933 (N_15933,N_15013,N_15353);
nor U15934 (N_15934,N_15245,N_15456);
nand U15935 (N_15935,N_15175,N_15033);
and U15936 (N_15936,N_15397,N_15238);
xor U15937 (N_15937,N_15195,N_15242);
nor U15938 (N_15938,N_15495,N_15107);
xnor U15939 (N_15939,N_15101,N_15462);
and U15940 (N_15940,N_15221,N_15163);
or U15941 (N_15941,N_15220,N_15248);
xor U15942 (N_15942,N_15393,N_15490);
and U15943 (N_15943,N_15099,N_15293);
nand U15944 (N_15944,N_15343,N_15001);
and U15945 (N_15945,N_15038,N_15037);
and U15946 (N_15946,N_15370,N_15183);
nor U15947 (N_15947,N_15009,N_15286);
or U15948 (N_15948,N_15150,N_15293);
or U15949 (N_15949,N_15305,N_15196);
nand U15950 (N_15950,N_15064,N_15431);
and U15951 (N_15951,N_15368,N_15113);
xor U15952 (N_15952,N_15412,N_15118);
or U15953 (N_15953,N_15107,N_15187);
nor U15954 (N_15954,N_15045,N_15359);
or U15955 (N_15955,N_15344,N_15208);
nor U15956 (N_15956,N_15293,N_15333);
nor U15957 (N_15957,N_15110,N_15466);
xnor U15958 (N_15958,N_15196,N_15182);
nand U15959 (N_15959,N_15381,N_15195);
nand U15960 (N_15960,N_15498,N_15346);
nand U15961 (N_15961,N_15409,N_15092);
or U15962 (N_15962,N_15481,N_15051);
and U15963 (N_15963,N_15247,N_15269);
and U15964 (N_15964,N_15454,N_15187);
xnor U15965 (N_15965,N_15109,N_15474);
and U15966 (N_15966,N_15203,N_15298);
xor U15967 (N_15967,N_15406,N_15064);
nor U15968 (N_15968,N_15140,N_15226);
nand U15969 (N_15969,N_15318,N_15373);
and U15970 (N_15970,N_15187,N_15216);
xor U15971 (N_15971,N_15051,N_15391);
nor U15972 (N_15972,N_15434,N_15019);
nor U15973 (N_15973,N_15077,N_15291);
nor U15974 (N_15974,N_15399,N_15078);
nand U15975 (N_15975,N_15268,N_15103);
or U15976 (N_15976,N_15307,N_15428);
and U15977 (N_15977,N_15382,N_15231);
xor U15978 (N_15978,N_15219,N_15056);
nand U15979 (N_15979,N_15045,N_15337);
or U15980 (N_15980,N_15033,N_15101);
nand U15981 (N_15981,N_15079,N_15140);
or U15982 (N_15982,N_15446,N_15322);
nor U15983 (N_15983,N_15447,N_15135);
and U15984 (N_15984,N_15342,N_15065);
nor U15985 (N_15985,N_15476,N_15347);
xor U15986 (N_15986,N_15043,N_15448);
xnor U15987 (N_15987,N_15354,N_15090);
or U15988 (N_15988,N_15345,N_15120);
nor U15989 (N_15989,N_15333,N_15032);
xor U15990 (N_15990,N_15488,N_15499);
and U15991 (N_15991,N_15062,N_15090);
and U15992 (N_15992,N_15333,N_15354);
or U15993 (N_15993,N_15207,N_15229);
nand U15994 (N_15994,N_15022,N_15347);
nor U15995 (N_15995,N_15280,N_15348);
nand U15996 (N_15996,N_15129,N_15004);
or U15997 (N_15997,N_15281,N_15168);
or U15998 (N_15998,N_15380,N_15262);
nor U15999 (N_15999,N_15497,N_15238);
nand U16000 (N_16000,N_15935,N_15587);
xnor U16001 (N_16001,N_15937,N_15977);
nor U16002 (N_16002,N_15851,N_15578);
xor U16003 (N_16003,N_15774,N_15758);
xor U16004 (N_16004,N_15765,N_15998);
or U16005 (N_16005,N_15622,N_15538);
xor U16006 (N_16006,N_15855,N_15603);
or U16007 (N_16007,N_15834,N_15678);
nand U16008 (N_16008,N_15683,N_15957);
xor U16009 (N_16009,N_15944,N_15575);
and U16010 (N_16010,N_15545,N_15674);
or U16011 (N_16011,N_15731,N_15679);
or U16012 (N_16012,N_15627,N_15671);
or U16013 (N_16013,N_15617,N_15767);
nor U16014 (N_16014,N_15543,N_15755);
xnor U16015 (N_16015,N_15684,N_15754);
and U16016 (N_16016,N_15509,N_15695);
or U16017 (N_16017,N_15879,N_15760);
nor U16018 (N_16018,N_15850,N_15925);
and U16019 (N_16019,N_15635,N_15905);
nor U16020 (N_16020,N_15886,N_15611);
or U16021 (N_16021,N_15697,N_15607);
or U16022 (N_16022,N_15835,N_15649);
nor U16023 (N_16023,N_15838,N_15621);
nor U16024 (N_16024,N_15900,N_15973);
and U16025 (N_16025,N_15849,N_15747);
nor U16026 (N_16026,N_15864,N_15595);
xor U16027 (N_16027,N_15664,N_15796);
nand U16028 (N_16028,N_15689,N_15985);
or U16029 (N_16029,N_15532,N_15544);
nor U16030 (N_16030,N_15797,N_15872);
nand U16031 (N_16031,N_15978,N_15856);
xnor U16032 (N_16032,N_15668,N_15517);
nand U16033 (N_16033,N_15554,N_15746);
or U16034 (N_16034,N_15921,N_15582);
nand U16035 (N_16035,N_15776,N_15688);
xnor U16036 (N_16036,N_15936,N_15637);
xnor U16037 (N_16037,N_15766,N_15564);
nor U16038 (N_16038,N_15772,N_15630);
and U16039 (N_16039,N_15616,N_15934);
or U16040 (N_16040,N_15522,N_15640);
or U16041 (N_16041,N_15682,N_15899);
nand U16042 (N_16042,N_15628,N_15923);
and U16043 (N_16043,N_15953,N_15823);
xor U16044 (N_16044,N_15784,N_15779);
or U16045 (N_16045,N_15503,N_15654);
nor U16046 (N_16046,N_15986,N_15815);
and U16047 (N_16047,N_15642,N_15819);
or U16048 (N_16048,N_15919,N_15818);
and U16049 (N_16049,N_15952,N_15696);
xor U16050 (N_16050,N_15605,N_15547);
nor U16051 (N_16051,N_15824,N_15876);
nand U16052 (N_16052,N_15928,N_15857);
or U16053 (N_16053,N_15887,N_15580);
xnor U16054 (N_16054,N_15918,N_15579);
nand U16055 (N_16055,N_15799,N_15828);
or U16056 (N_16056,N_15782,N_15902);
xor U16057 (N_16057,N_15994,N_15894);
nand U16058 (N_16058,N_15585,N_15559);
nand U16059 (N_16059,N_15787,N_15940);
nor U16060 (N_16060,N_15593,N_15576);
nor U16061 (N_16061,N_15577,N_15993);
and U16062 (N_16062,N_15552,N_15681);
or U16063 (N_16063,N_15891,N_15658);
nor U16064 (N_16064,N_15715,N_15553);
or U16065 (N_16065,N_15996,N_15656);
and U16066 (N_16066,N_15811,N_15609);
xor U16067 (N_16067,N_15941,N_15614);
or U16068 (N_16068,N_15694,N_15631);
and U16069 (N_16069,N_15868,N_15558);
nor U16070 (N_16070,N_15992,N_15969);
or U16071 (N_16071,N_15536,N_15505);
nor U16072 (N_16072,N_15926,N_15676);
nand U16073 (N_16073,N_15967,N_15659);
nor U16074 (N_16074,N_15634,N_15653);
and U16075 (N_16075,N_15865,N_15955);
nor U16076 (N_16076,N_15680,N_15665);
xnor U16077 (N_16077,N_15572,N_15590);
nand U16078 (N_16078,N_15860,N_15743);
xnor U16079 (N_16079,N_15730,N_15963);
nor U16080 (N_16080,N_15862,N_15749);
or U16081 (N_16081,N_15939,N_15852);
nand U16082 (N_16082,N_15541,N_15652);
or U16083 (N_16083,N_15848,N_15639);
xnor U16084 (N_16084,N_15707,N_15521);
nor U16085 (N_16085,N_15817,N_15647);
xor U16086 (N_16086,N_15870,N_15650);
nor U16087 (N_16087,N_15563,N_15720);
nor U16088 (N_16088,N_15685,N_15624);
nor U16089 (N_16089,N_15947,N_15691);
nor U16090 (N_16090,N_15945,N_15657);
xnor U16091 (N_16091,N_15518,N_15507);
and U16092 (N_16092,N_15878,N_15795);
nand U16093 (N_16093,N_15863,N_15924);
nand U16094 (N_16094,N_15913,N_15897);
or U16095 (N_16095,N_15636,N_15798);
xnor U16096 (N_16096,N_15903,N_15775);
or U16097 (N_16097,N_15506,N_15602);
nand U16098 (N_16098,N_15556,N_15980);
nand U16099 (N_16099,N_15740,N_15672);
nor U16100 (N_16100,N_15589,N_15946);
nor U16101 (N_16101,N_15839,N_15723);
nor U16102 (N_16102,N_15845,N_15698);
nand U16103 (N_16103,N_15802,N_15666);
nand U16104 (N_16104,N_15990,N_15830);
or U16105 (N_16105,N_15546,N_15531);
or U16106 (N_16106,N_15927,N_15898);
nand U16107 (N_16107,N_15771,N_15513);
xor U16108 (N_16108,N_15997,N_15904);
or U16109 (N_16109,N_15801,N_15808);
nand U16110 (N_16110,N_15648,N_15738);
and U16111 (N_16111,N_15504,N_15592);
or U16112 (N_16112,N_15523,N_15644);
or U16113 (N_16113,N_15524,N_15822);
or U16114 (N_16114,N_15551,N_15979);
nor U16115 (N_16115,N_15831,N_15560);
nor U16116 (N_16116,N_15951,N_15929);
xnor U16117 (N_16117,N_15833,N_15701);
xor U16118 (N_16118,N_15510,N_15528);
nand U16119 (N_16119,N_15885,N_15999);
nor U16120 (N_16120,N_15972,N_15709);
and U16121 (N_16121,N_15596,N_15514);
and U16122 (N_16122,N_15670,N_15932);
xnor U16123 (N_16123,N_15882,N_15566);
xor U16124 (N_16124,N_15608,N_15805);
nand U16125 (N_16125,N_15873,N_15598);
and U16126 (N_16126,N_15761,N_15511);
and U16127 (N_16127,N_15555,N_15705);
xnor U16128 (N_16128,N_15804,N_15909);
and U16129 (N_16129,N_15539,N_15520);
and U16130 (N_16130,N_15949,N_15610);
nand U16131 (N_16131,N_15700,N_15778);
xor U16132 (N_16132,N_15569,N_15962);
xor U16133 (N_16133,N_15806,N_15821);
nand U16134 (N_16134,N_15906,N_15661);
and U16135 (N_16135,N_15571,N_15807);
nor U16136 (N_16136,N_15599,N_15846);
nor U16137 (N_16137,N_15901,N_15620);
nor U16138 (N_16138,N_15959,N_15515);
nand U16139 (N_16139,N_15537,N_15714);
or U16140 (N_16140,N_15750,N_15525);
and U16141 (N_16141,N_15508,N_15966);
xnor U16142 (N_16142,N_15859,N_15742);
and U16143 (N_16143,N_15867,N_15744);
nor U16144 (N_16144,N_15718,N_15646);
and U16145 (N_16145,N_15764,N_15843);
nor U16146 (N_16146,N_15726,N_15703);
and U16147 (N_16147,N_15727,N_15641);
nor U16148 (N_16148,N_15884,N_15570);
or U16149 (N_16149,N_15548,N_15988);
and U16150 (N_16150,N_15768,N_15791);
or U16151 (N_16151,N_15663,N_15780);
or U16152 (N_16152,N_15721,N_15713);
nor U16153 (N_16153,N_15989,N_15890);
nor U16154 (N_16154,N_15619,N_15875);
nor U16155 (N_16155,N_15888,N_15915);
or U16156 (N_16156,N_15914,N_15974);
nand U16157 (N_16157,N_15583,N_15529);
nor U16158 (N_16158,N_15604,N_15734);
nor U16159 (N_16159,N_15789,N_15662);
and U16160 (N_16160,N_15623,N_15943);
and U16161 (N_16161,N_15550,N_15724);
and U16162 (N_16162,N_15773,N_15748);
or U16163 (N_16163,N_15655,N_15896);
xor U16164 (N_16164,N_15785,N_15594);
nand U16165 (N_16165,N_15983,N_15908);
xor U16166 (N_16166,N_15597,N_15601);
nor U16167 (N_16167,N_15812,N_15675);
and U16168 (N_16168,N_15788,N_15673);
nand U16169 (N_16169,N_15920,N_15892);
and U16170 (N_16170,N_15858,N_15557);
or U16171 (N_16171,N_15710,N_15814);
or U16172 (N_16172,N_15792,N_15618);
xor U16173 (N_16173,N_15954,N_15573);
xnor U16174 (N_16174,N_15816,N_15677);
and U16175 (N_16175,N_15794,N_15752);
nand U16176 (N_16176,N_15991,N_15739);
and U16177 (N_16177,N_15971,N_15519);
nand U16178 (N_16178,N_15753,N_15948);
and U16179 (N_16179,N_15931,N_15736);
nor U16180 (N_16180,N_15567,N_15832);
xor U16181 (N_16181,N_15964,N_15874);
or U16182 (N_16182,N_15600,N_15840);
nand U16183 (N_16183,N_15651,N_15741);
nor U16184 (N_16184,N_15933,N_15910);
nand U16185 (N_16185,N_15629,N_15716);
xnor U16186 (N_16186,N_15712,N_15781);
xor U16187 (N_16187,N_15615,N_15638);
or U16188 (N_16188,N_15693,N_15961);
xnor U16189 (N_16189,N_15893,N_15722);
nor U16190 (N_16190,N_15861,N_15733);
or U16191 (N_16191,N_15632,N_15869);
nand U16192 (N_16192,N_15568,N_15708);
nand U16193 (N_16193,N_15813,N_15692);
and U16194 (N_16194,N_15975,N_15895);
nor U16195 (N_16195,N_15976,N_15699);
nand U16196 (N_16196,N_15820,N_15826);
nor U16197 (N_16197,N_15588,N_15565);
or U16198 (N_16198,N_15725,N_15881);
and U16199 (N_16199,N_15965,N_15633);
nor U16200 (N_16200,N_15917,N_15667);
and U16201 (N_16201,N_15526,N_15759);
or U16202 (N_16202,N_15690,N_15956);
or U16203 (N_16203,N_15502,N_15591);
and U16204 (N_16204,N_15769,N_15916);
xor U16205 (N_16205,N_15732,N_15613);
nor U16206 (N_16206,N_15837,N_15803);
and U16207 (N_16207,N_15880,N_15745);
xnor U16208 (N_16208,N_15540,N_15930);
nand U16209 (N_16209,N_15687,N_15883);
and U16210 (N_16210,N_15729,N_15810);
nand U16211 (N_16211,N_15842,N_15500);
or U16212 (N_16212,N_15853,N_15751);
nand U16213 (N_16213,N_15702,N_15960);
nor U16214 (N_16214,N_15756,N_15660);
or U16215 (N_16215,N_15841,N_15866);
nor U16216 (N_16216,N_15763,N_15786);
nor U16217 (N_16217,N_15827,N_15606);
nor U16218 (N_16218,N_15911,N_15711);
or U16219 (N_16219,N_15790,N_15777);
and U16220 (N_16220,N_15530,N_15871);
nand U16221 (N_16221,N_15501,N_15686);
nand U16222 (N_16222,N_15844,N_15950);
or U16223 (N_16223,N_15829,N_15561);
nor U16224 (N_16224,N_15626,N_15757);
nand U16225 (N_16225,N_15581,N_15527);
xnor U16226 (N_16226,N_15535,N_15669);
nand U16227 (N_16227,N_15562,N_15534);
or U16228 (N_16228,N_15719,N_15889);
and U16229 (N_16229,N_15737,N_15970);
and U16230 (N_16230,N_15982,N_15981);
nor U16231 (N_16231,N_15987,N_15783);
xnor U16232 (N_16232,N_15912,N_15717);
xnor U16233 (N_16233,N_15907,N_15922);
or U16234 (N_16234,N_15728,N_15512);
nor U16235 (N_16235,N_15574,N_15612);
xnor U16236 (N_16236,N_15770,N_15995);
or U16237 (N_16237,N_15938,N_15854);
xnor U16238 (N_16238,N_15516,N_15847);
xor U16239 (N_16239,N_15809,N_15549);
nor U16240 (N_16240,N_15942,N_15533);
nor U16241 (N_16241,N_15542,N_15984);
nor U16242 (N_16242,N_15877,N_15704);
nor U16243 (N_16243,N_15706,N_15625);
nand U16244 (N_16244,N_15793,N_15762);
and U16245 (N_16245,N_15645,N_15735);
nand U16246 (N_16246,N_15958,N_15586);
and U16247 (N_16247,N_15584,N_15825);
nand U16248 (N_16248,N_15968,N_15836);
nand U16249 (N_16249,N_15643,N_15800);
nor U16250 (N_16250,N_15942,N_15787);
nand U16251 (N_16251,N_15504,N_15848);
xnor U16252 (N_16252,N_15694,N_15737);
nor U16253 (N_16253,N_15608,N_15617);
or U16254 (N_16254,N_15874,N_15982);
xnor U16255 (N_16255,N_15748,N_15963);
nor U16256 (N_16256,N_15903,N_15756);
xor U16257 (N_16257,N_15962,N_15835);
and U16258 (N_16258,N_15755,N_15976);
or U16259 (N_16259,N_15524,N_15942);
nor U16260 (N_16260,N_15896,N_15531);
or U16261 (N_16261,N_15562,N_15665);
nor U16262 (N_16262,N_15863,N_15517);
xor U16263 (N_16263,N_15951,N_15639);
or U16264 (N_16264,N_15781,N_15543);
xnor U16265 (N_16265,N_15872,N_15946);
or U16266 (N_16266,N_15968,N_15568);
xnor U16267 (N_16267,N_15651,N_15849);
nor U16268 (N_16268,N_15628,N_15911);
and U16269 (N_16269,N_15627,N_15767);
xor U16270 (N_16270,N_15764,N_15548);
xnor U16271 (N_16271,N_15536,N_15728);
and U16272 (N_16272,N_15654,N_15656);
and U16273 (N_16273,N_15862,N_15641);
nor U16274 (N_16274,N_15701,N_15995);
xnor U16275 (N_16275,N_15836,N_15611);
nor U16276 (N_16276,N_15578,N_15516);
or U16277 (N_16277,N_15590,N_15691);
and U16278 (N_16278,N_15637,N_15777);
xor U16279 (N_16279,N_15561,N_15911);
xnor U16280 (N_16280,N_15897,N_15730);
and U16281 (N_16281,N_15659,N_15703);
nor U16282 (N_16282,N_15511,N_15700);
or U16283 (N_16283,N_15803,N_15611);
and U16284 (N_16284,N_15610,N_15940);
xor U16285 (N_16285,N_15709,N_15904);
xnor U16286 (N_16286,N_15784,N_15958);
or U16287 (N_16287,N_15703,N_15594);
nand U16288 (N_16288,N_15802,N_15663);
and U16289 (N_16289,N_15531,N_15914);
and U16290 (N_16290,N_15736,N_15799);
nor U16291 (N_16291,N_15773,N_15628);
and U16292 (N_16292,N_15832,N_15641);
nor U16293 (N_16293,N_15984,N_15858);
nand U16294 (N_16294,N_15615,N_15855);
nor U16295 (N_16295,N_15696,N_15692);
nor U16296 (N_16296,N_15568,N_15691);
xor U16297 (N_16297,N_15769,N_15782);
and U16298 (N_16298,N_15572,N_15742);
nand U16299 (N_16299,N_15752,N_15875);
nand U16300 (N_16300,N_15536,N_15576);
xnor U16301 (N_16301,N_15747,N_15744);
nor U16302 (N_16302,N_15587,N_15882);
nand U16303 (N_16303,N_15773,N_15596);
nand U16304 (N_16304,N_15809,N_15502);
nand U16305 (N_16305,N_15986,N_15520);
xor U16306 (N_16306,N_15508,N_15908);
xor U16307 (N_16307,N_15628,N_15919);
nand U16308 (N_16308,N_15798,N_15894);
and U16309 (N_16309,N_15925,N_15563);
and U16310 (N_16310,N_15718,N_15592);
or U16311 (N_16311,N_15599,N_15960);
nand U16312 (N_16312,N_15511,N_15685);
and U16313 (N_16313,N_15713,N_15508);
nand U16314 (N_16314,N_15808,N_15702);
xnor U16315 (N_16315,N_15947,N_15897);
xor U16316 (N_16316,N_15639,N_15820);
or U16317 (N_16317,N_15591,N_15815);
or U16318 (N_16318,N_15990,N_15753);
and U16319 (N_16319,N_15738,N_15528);
or U16320 (N_16320,N_15672,N_15617);
and U16321 (N_16321,N_15694,N_15987);
nand U16322 (N_16322,N_15637,N_15606);
nor U16323 (N_16323,N_15617,N_15756);
xor U16324 (N_16324,N_15543,N_15616);
and U16325 (N_16325,N_15543,N_15716);
and U16326 (N_16326,N_15870,N_15568);
or U16327 (N_16327,N_15612,N_15548);
nand U16328 (N_16328,N_15666,N_15905);
and U16329 (N_16329,N_15752,N_15611);
xor U16330 (N_16330,N_15656,N_15883);
nand U16331 (N_16331,N_15678,N_15985);
nand U16332 (N_16332,N_15689,N_15864);
nand U16333 (N_16333,N_15706,N_15539);
nand U16334 (N_16334,N_15752,N_15643);
or U16335 (N_16335,N_15624,N_15826);
and U16336 (N_16336,N_15729,N_15570);
nor U16337 (N_16337,N_15616,N_15963);
and U16338 (N_16338,N_15549,N_15784);
and U16339 (N_16339,N_15917,N_15994);
nand U16340 (N_16340,N_15859,N_15730);
and U16341 (N_16341,N_15735,N_15581);
nand U16342 (N_16342,N_15805,N_15963);
xor U16343 (N_16343,N_15828,N_15933);
or U16344 (N_16344,N_15831,N_15791);
nand U16345 (N_16345,N_15973,N_15839);
nand U16346 (N_16346,N_15987,N_15543);
nor U16347 (N_16347,N_15537,N_15572);
and U16348 (N_16348,N_15848,N_15580);
nand U16349 (N_16349,N_15608,N_15923);
nand U16350 (N_16350,N_15900,N_15667);
xor U16351 (N_16351,N_15579,N_15606);
or U16352 (N_16352,N_15914,N_15676);
nand U16353 (N_16353,N_15716,N_15879);
nand U16354 (N_16354,N_15757,N_15762);
and U16355 (N_16355,N_15682,N_15740);
or U16356 (N_16356,N_15945,N_15822);
or U16357 (N_16357,N_15623,N_15560);
and U16358 (N_16358,N_15824,N_15999);
or U16359 (N_16359,N_15700,N_15674);
xnor U16360 (N_16360,N_15852,N_15523);
nand U16361 (N_16361,N_15596,N_15712);
xor U16362 (N_16362,N_15811,N_15802);
nand U16363 (N_16363,N_15843,N_15863);
xnor U16364 (N_16364,N_15615,N_15889);
xor U16365 (N_16365,N_15716,N_15563);
nand U16366 (N_16366,N_15642,N_15641);
xnor U16367 (N_16367,N_15552,N_15719);
xor U16368 (N_16368,N_15896,N_15764);
xor U16369 (N_16369,N_15787,N_15633);
nand U16370 (N_16370,N_15840,N_15779);
nor U16371 (N_16371,N_15936,N_15806);
nand U16372 (N_16372,N_15558,N_15729);
nand U16373 (N_16373,N_15871,N_15714);
or U16374 (N_16374,N_15545,N_15608);
nor U16375 (N_16375,N_15638,N_15599);
xor U16376 (N_16376,N_15879,N_15693);
and U16377 (N_16377,N_15898,N_15531);
xnor U16378 (N_16378,N_15738,N_15599);
xor U16379 (N_16379,N_15671,N_15778);
xor U16380 (N_16380,N_15661,N_15800);
or U16381 (N_16381,N_15506,N_15597);
nor U16382 (N_16382,N_15698,N_15689);
or U16383 (N_16383,N_15500,N_15859);
nor U16384 (N_16384,N_15529,N_15649);
xor U16385 (N_16385,N_15690,N_15600);
nand U16386 (N_16386,N_15731,N_15765);
nor U16387 (N_16387,N_15579,N_15985);
nand U16388 (N_16388,N_15535,N_15924);
nand U16389 (N_16389,N_15789,N_15829);
and U16390 (N_16390,N_15593,N_15749);
nand U16391 (N_16391,N_15988,N_15610);
nand U16392 (N_16392,N_15903,N_15735);
xnor U16393 (N_16393,N_15901,N_15863);
nand U16394 (N_16394,N_15780,N_15798);
nand U16395 (N_16395,N_15754,N_15767);
nor U16396 (N_16396,N_15601,N_15612);
xnor U16397 (N_16397,N_15986,N_15674);
nand U16398 (N_16398,N_15880,N_15630);
nor U16399 (N_16399,N_15668,N_15770);
and U16400 (N_16400,N_15675,N_15931);
or U16401 (N_16401,N_15839,N_15555);
xor U16402 (N_16402,N_15759,N_15578);
and U16403 (N_16403,N_15713,N_15728);
xor U16404 (N_16404,N_15949,N_15735);
xnor U16405 (N_16405,N_15762,N_15670);
xor U16406 (N_16406,N_15769,N_15940);
nor U16407 (N_16407,N_15764,N_15616);
nand U16408 (N_16408,N_15565,N_15744);
or U16409 (N_16409,N_15984,N_15934);
nand U16410 (N_16410,N_15879,N_15973);
nor U16411 (N_16411,N_15513,N_15989);
or U16412 (N_16412,N_15719,N_15888);
and U16413 (N_16413,N_15948,N_15658);
and U16414 (N_16414,N_15511,N_15525);
nand U16415 (N_16415,N_15726,N_15873);
xnor U16416 (N_16416,N_15514,N_15787);
nand U16417 (N_16417,N_15585,N_15861);
xor U16418 (N_16418,N_15756,N_15506);
nand U16419 (N_16419,N_15578,N_15686);
and U16420 (N_16420,N_15716,N_15576);
nor U16421 (N_16421,N_15888,N_15606);
nand U16422 (N_16422,N_15714,N_15796);
xnor U16423 (N_16423,N_15754,N_15733);
xnor U16424 (N_16424,N_15569,N_15595);
and U16425 (N_16425,N_15534,N_15810);
nand U16426 (N_16426,N_15593,N_15644);
nor U16427 (N_16427,N_15974,N_15718);
nand U16428 (N_16428,N_15555,N_15547);
and U16429 (N_16429,N_15875,N_15739);
nor U16430 (N_16430,N_15663,N_15502);
xor U16431 (N_16431,N_15811,N_15789);
nor U16432 (N_16432,N_15786,N_15561);
nor U16433 (N_16433,N_15823,N_15694);
or U16434 (N_16434,N_15804,N_15888);
or U16435 (N_16435,N_15820,N_15686);
nand U16436 (N_16436,N_15791,N_15803);
and U16437 (N_16437,N_15651,N_15740);
or U16438 (N_16438,N_15841,N_15885);
or U16439 (N_16439,N_15588,N_15632);
xnor U16440 (N_16440,N_15678,N_15627);
nand U16441 (N_16441,N_15762,N_15618);
nor U16442 (N_16442,N_15788,N_15507);
xnor U16443 (N_16443,N_15513,N_15506);
and U16444 (N_16444,N_15676,N_15948);
and U16445 (N_16445,N_15889,N_15835);
xnor U16446 (N_16446,N_15655,N_15890);
and U16447 (N_16447,N_15523,N_15645);
nor U16448 (N_16448,N_15958,N_15549);
nor U16449 (N_16449,N_15520,N_15611);
or U16450 (N_16450,N_15802,N_15723);
and U16451 (N_16451,N_15772,N_15673);
nor U16452 (N_16452,N_15731,N_15650);
nor U16453 (N_16453,N_15888,N_15507);
nand U16454 (N_16454,N_15716,N_15949);
and U16455 (N_16455,N_15931,N_15559);
or U16456 (N_16456,N_15974,N_15518);
nor U16457 (N_16457,N_15837,N_15792);
and U16458 (N_16458,N_15832,N_15679);
or U16459 (N_16459,N_15529,N_15975);
or U16460 (N_16460,N_15503,N_15909);
nand U16461 (N_16461,N_15778,N_15752);
xor U16462 (N_16462,N_15786,N_15737);
nor U16463 (N_16463,N_15938,N_15658);
or U16464 (N_16464,N_15551,N_15665);
nand U16465 (N_16465,N_15702,N_15611);
and U16466 (N_16466,N_15971,N_15514);
and U16467 (N_16467,N_15821,N_15594);
xnor U16468 (N_16468,N_15801,N_15858);
or U16469 (N_16469,N_15647,N_15852);
or U16470 (N_16470,N_15730,N_15711);
nor U16471 (N_16471,N_15643,N_15711);
xnor U16472 (N_16472,N_15753,N_15894);
xnor U16473 (N_16473,N_15580,N_15711);
nand U16474 (N_16474,N_15839,N_15891);
and U16475 (N_16475,N_15630,N_15750);
nand U16476 (N_16476,N_15757,N_15759);
or U16477 (N_16477,N_15816,N_15649);
nand U16478 (N_16478,N_15579,N_15778);
and U16479 (N_16479,N_15638,N_15821);
nand U16480 (N_16480,N_15677,N_15593);
and U16481 (N_16481,N_15650,N_15811);
nand U16482 (N_16482,N_15851,N_15951);
xor U16483 (N_16483,N_15750,N_15899);
xnor U16484 (N_16484,N_15580,N_15586);
and U16485 (N_16485,N_15976,N_15722);
nor U16486 (N_16486,N_15743,N_15990);
xor U16487 (N_16487,N_15921,N_15839);
nor U16488 (N_16488,N_15806,N_15840);
and U16489 (N_16489,N_15743,N_15700);
xnor U16490 (N_16490,N_15879,N_15828);
or U16491 (N_16491,N_15578,N_15981);
and U16492 (N_16492,N_15597,N_15501);
xor U16493 (N_16493,N_15551,N_15836);
nand U16494 (N_16494,N_15651,N_15547);
or U16495 (N_16495,N_15890,N_15665);
or U16496 (N_16496,N_15799,N_15730);
or U16497 (N_16497,N_15725,N_15593);
or U16498 (N_16498,N_15948,N_15597);
or U16499 (N_16499,N_15551,N_15526);
nor U16500 (N_16500,N_16121,N_16248);
nor U16501 (N_16501,N_16162,N_16331);
nand U16502 (N_16502,N_16055,N_16315);
or U16503 (N_16503,N_16283,N_16139);
nand U16504 (N_16504,N_16234,N_16375);
and U16505 (N_16505,N_16175,N_16026);
or U16506 (N_16506,N_16452,N_16423);
nand U16507 (N_16507,N_16108,N_16036);
or U16508 (N_16508,N_16437,N_16485);
nor U16509 (N_16509,N_16345,N_16113);
nor U16510 (N_16510,N_16324,N_16300);
nor U16511 (N_16511,N_16314,N_16313);
xnor U16512 (N_16512,N_16465,N_16075);
nand U16513 (N_16513,N_16052,N_16262);
nand U16514 (N_16514,N_16088,N_16021);
xnor U16515 (N_16515,N_16031,N_16002);
xnor U16516 (N_16516,N_16486,N_16280);
nor U16517 (N_16517,N_16080,N_16260);
xnor U16518 (N_16518,N_16250,N_16096);
nand U16519 (N_16519,N_16196,N_16288);
and U16520 (N_16520,N_16320,N_16076);
and U16521 (N_16521,N_16286,N_16063);
nand U16522 (N_16522,N_16073,N_16064);
xor U16523 (N_16523,N_16398,N_16351);
xor U16524 (N_16524,N_16207,N_16428);
and U16525 (N_16525,N_16455,N_16246);
nand U16526 (N_16526,N_16359,N_16144);
nand U16527 (N_16527,N_16176,N_16179);
nand U16528 (N_16528,N_16391,N_16243);
and U16529 (N_16529,N_16186,N_16125);
nor U16530 (N_16530,N_16174,N_16274);
xnor U16531 (N_16531,N_16124,N_16215);
and U16532 (N_16532,N_16466,N_16082);
or U16533 (N_16533,N_16289,N_16490);
nand U16534 (N_16534,N_16358,N_16384);
nor U16535 (N_16535,N_16028,N_16214);
xnor U16536 (N_16536,N_16464,N_16342);
and U16537 (N_16537,N_16387,N_16161);
nor U16538 (N_16538,N_16221,N_16239);
or U16539 (N_16539,N_16279,N_16419);
and U16540 (N_16540,N_16166,N_16449);
or U16541 (N_16541,N_16010,N_16426);
nand U16542 (N_16542,N_16103,N_16429);
nor U16543 (N_16543,N_16296,N_16399);
xor U16544 (N_16544,N_16090,N_16475);
nor U16545 (N_16545,N_16258,N_16167);
and U16546 (N_16546,N_16456,N_16462);
and U16547 (N_16547,N_16370,N_16406);
or U16548 (N_16548,N_16290,N_16381);
nand U16549 (N_16549,N_16413,N_16295);
and U16550 (N_16550,N_16377,N_16257);
xnor U16551 (N_16551,N_16086,N_16050);
xnor U16552 (N_16552,N_16083,N_16453);
nor U16553 (N_16553,N_16225,N_16172);
and U16554 (N_16554,N_16253,N_16322);
nand U16555 (N_16555,N_16478,N_16200);
and U16556 (N_16556,N_16306,N_16066);
xor U16557 (N_16557,N_16037,N_16034);
and U16558 (N_16558,N_16111,N_16056);
nor U16559 (N_16559,N_16224,N_16302);
nand U16560 (N_16560,N_16079,N_16335);
nand U16561 (N_16561,N_16402,N_16321);
xor U16562 (N_16562,N_16187,N_16035);
xnor U16563 (N_16563,N_16163,N_16140);
and U16564 (N_16564,N_16275,N_16433);
or U16565 (N_16565,N_16077,N_16450);
and U16566 (N_16566,N_16194,N_16198);
xor U16567 (N_16567,N_16460,N_16434);
nor U16568 (N_16568,N_16154,N_16308);
nand U16569 (N_16569,N_16061,N_16444);
and U16570 (N_16570,N_16007,N_16023);
and U16571 (N_16571,N_16164,N_16488);
nor U16572 (N_16572,N_16327,N_16467);
nand U16573 (N_16573,N_16134,N_16087);
nor U16574 (N_16574,N_16411,N_16192);
nand U16575 (N_16575,N_16477,N_16223);
xnor U16576 (N_16576,N_16326,N_16158);
nand U16577 (N_16577,N_16285,N_16364);
nand U16578 (N_16578,N_16059,N_16481);
xnor U16579 (N_16579,N_16143,N_16014);
or U16580 (N_16580,N_16222,N_16123);
nor U16581 (N_16581,N_16118,N_16251);
or U16582 (N_16582,N_16183,N_16040);
nor U16583 (N_16583,N_16092,N_16440);
nor U16584 (N_16584,N_16084,N_16181);
and U16585 (N_16585,N_16003,N_16271);
nand U16586 (N_16586,N_16380,N_16135);
xnor U16587 (N_16587,N_16311,N_16304);
nor U16588 (N_16588,N_16017,N_16393);
and U16589 (N_16589,N_16340,N_16093);
nor U16590 (N_16590,N_16137,N_16138);
and U16591 (N_16591,N_16392,N_16483);
nand U16592 (N_16592,N_16217,N_16469);
nand U16593 (N_16593,N_16305,N_16430);
xor U16594 (N_16594,N_16307,N_16498);
nand U16595 (N_16595,N_16199,N_16471);
xor U16596 (N_16596,N_16045,N_16152);
or U16597 (N_16597,N_16316,N_16266);
nor U16598 (N_16598,N_16474,N_16106);
nor U16599 (N_16599,N_16448,N_16104);
nor U16600 (N_16600,N_16150,N_16357);
xnor U16601 (N_16601,N_16097,N_16493);
xor U16602 (N_16602,N_16165,N_16408);
nand U16603 (N_16603,N_16048,N_16197);
or U16604 (N_16604,N_16227,N_16356);
and U16605 (N_16605,N_16293,N_16382);
xnor U16606 (N_16606,N_16202,N_16427);
nor U16607 (N_16607,N_16168,N_16386);
nand U16608 (N_16608,N_16182,N_16269);
and U16609 (N_16609,N_16332,N_16329);
and U16610 (N_16610,N_16365,N_16057);
nand U16611 (N_16611,N_16233,N_16213);
nand U16612 (N_16612,N_16360,N_16041);
xor U16613 (N_16613,N_16229,N_16114);
nand U16614 (N_16614,N_16424,N_16185);
nand U16615 (N_16615,N_16497,N_16496);
nor U16616 (N_16616,N_16212,N_16336);
and U16617 (N_16617,N_16190,N_16008);
and U16618 (N_16618,N_16015,N_16303);
or U16619 (N_16619,N_16282,N_16383);
and U16620 (N_16620,N_16495,N_16441);
nor U16621 (N_16621,N_16232,N_16339);
or U16622 (N_16622,N_16346,N_16349);
and U16623 (N_16623,N_16030,N_16268);
nor U16624 (N_16624,N_16115,N_16270);
or U16625 (N_16625,N_16344,N_16415);
nand U16626 (N_16626,N_16294,N_16334);
xnor U16627 (N_16627,N_16043,N_16119);
xor U16628 (N_16628,N_16319,N_16065);
xor U16629 (N_16629,N_16219,N_16394);
and U16630 (N_16630,N_16445,N_16407);
nor U16631 (N_16631,N_16470,N_16244);
or U16632 (N_16632,N_16473,N_16206);
and U16633 (N_16633,N_16350,N_16362);
or U16634 (N_16634,N_16401,N_16173);
and U16635 (N_16635,N_16395,N_16371);
nor U16636 (N_16636,N_16278,N_16482);
or U16637 (N_16637,N_16385,N_16019);
nand U16638 (N_16638,N_16341,N_16325);
xnor U16639 (N_16639,N_16001,N_16130);
or U16640 (N_16640,N_16072,N_16128);
nand U16641 (N_16641,N_16204,N_16405);
or U16642 (N_16642,N_16102,N_16238);
xor U16643 (N_16643,N_16029,N_16442);
or U16644 (N_16644,N_16338,N_16403);
xnor U16645 (N_16645,N_16012,N_16425);
and U16646 (N_16646,N_16169,N_16291);
and U16647 (N_16647,N_16309,N_16101);
nor U16648 (N_16648,N_16369,N_16265);
and U16649 (N_16649,N_16074,N_16374);
and U16650 (N_16650,N_16151,N_16112);
nor U16651 (N_16651,N_16027,N_16414);
nor U16652 (N_16652,N_16127,N_16312);
or U16653 (N_16653,N_16256,N_16348);
xnor U16654 (N_16654,N_16170,N_16276);
xor U16655 (N_16655,N_16236,N_16107);
and U16656 (N_16656,N_16211,N_16218);
nor U16657 (N_16657,N_16435,N_16067);
nor U16658 (N_16658,N_16155,N_16390);
xor U16659 (N_16659,N_16353,N_16153);
nand U16660 (N_16660,N_16226,N_16489);
and U16661 (N_16661,N_16432,N_16020);
xnor U16662 (N_16662,N_16228,N_16141);
nand U16663 (N_16663,N_16006,N_16000);
and U16664 (N_16664,N_16171,N_16409);
nand U16665 (N_16665,N_16458,N_16231);
xor U16666 (N_16666,N_16259,N_16355);
nor U16667 (N_16667,N_16318,N_16053);
and U16668 (N_16668,N_16177,N_16047);
nor U16669 (N_16669,N_16272,N_16400);
nand U16670 (N_16670,N_16046,N_16094);
nand U16671 (N_16671,N_16373,N_16039);
xnor U16672 (N_16672,N_16418,N_16343);
nor U16673 (N_16673,N_16195,N_16463);
or U16674 (N_16674,N_16438,N_16044);
xnor U16675 (N_16675,N_16230,N_16347);
nor U16676 (N_16676,N_16476,N_16091);
nand U16677 (N_16677,N_16038,N_16479);
nand U16678 (N_16678,N_16060,N_16443);
nand U16679 (N_16679,N_16252,N_16013);
or U16680 (N_16680,N_16416,N_16264);
nand U16681 (N_16681,N_16049,N_16468);
nand U16682 (N_16682,N_16042,N_16116);
xnor U16683 (N_16683,N_16297,N_16009);
or U16684 (N_16684,N_16454,N_16189);
nor U16685 (N_16685,N_16148,N_16254);
or U16686 (N_16686,N_16068,N_16397);
and U16687 (N_16687,N_16378,N_16491);
nand U16688 (N_16688,N_16210,N_16180);
xor U16689 (N_16689,N_16484,N_16089);
nand U16690 (N_16690,N_16368,N_16298);
nand U16691 (N_16691,N_16142,N_16421);
and U16692 (N_16692,N_16022,N_16147);
and U16693 (N_16693,N_16081,N_16203);
nor U16694 (N_16694,N_16281,N_16354);
xnor U16695 (N_16695,N_16145,N_16051);
nand U16696 (N_16696,N_16299,N_16024);
or U16697 (N_16697,N_16404,N_16191);
nand U16698 (N_16698,N_16494,N_16284);
nor U16699 (N_16699,N_16417,N_16133);
nand U16700 (N_16700,N_16457,N_16372);
or U16701 (N_16701,N_16439,N_16287);
and U16702 (N_16702,N_16267,N_16328);
nand U16703 (N_16703,N_16188,N_16005);
nand U16704 (N_16704,N_16277,N_16241);
nand U16705 (N_16705,N_16160,N_16396);
nor U16706 (N_16706,N_16205,N_16178);
nor U16707 (N_16707,N_16447,N_16480);
nand U16708 (N_16708,N_16184,N_16245);
nor U16709 (N_16709,N_16201,N_16193);
or U16710 (N_16710,N_16011,N_16105);
and U16711 (N_16711,N_16025,N_16157);
and U16712 (N_16712,N_16033,N_16420);
or U16713 (N_16713,N_16255,N_16366);
nand U16714 (N_16714,N_16240,N_16110);
or U16715 (N_16715,N_16099,N_16126);
nand U16716 (N_16716,N_16247,N_16436);
xnor U16717 (N_16717,N_16136,N_16078);
nand U16718 (N_16718,N_16363,N_16209);
nand U16719 (N_16719,N_16451,N_16208);
or U16720 (N_16720,N_16129,N_16410);
or U16721 (N_16721,N_16146,N_16054);
nand U16722 (N_16722,N_16117,N_16098);
nor U16723 (N_16723,N_16412,N_16132);
nand U16724 (N_16724,N_16249,N_16273);
nor U16725 (N_16725,N_16263,N_16085);
or U16726 (N_16726,N_16376,N_16422);
and U16727 (N_16727,N_16310,N_16492);
nor U16728 (N_16728,N_16100,N_16032);
xnor U16729 (N_16729,N_16237,N_16388);
or U16730 (N_16730,N_16018,N_16216);
and U16731 (N_16731,N_16361,N_16109);
nand U16732 (N_16732,N_16337,N_16333);
xor U16733 (N_16733,N_16461,N_16062);
and U16734 (N_16734,N_16242,N_16069);
xnor U16735 (N_16735,N_16235,N_16487);
xor U16736 (N_16736,N_16352,N_16446);
xor U16737 (N_16737,N_16004,N_16016);
nor U16738 (N_16738,N_16431,N_16220);
nand U16739 (N_16739,N_16071,N_16292);
xnor U16740 (N_16740,N_16389,N_16379);
and U16741 (N_16741,N_16301,N_16472);
or U16742 (N_16742,N_16323,N_16122);
nand U16743 (N_16743,N_16159,N_16367);
or U16744 (N_16744,N_16120,N_16058);
nand U16745 (N_16745,N_16317,N_16459);
xor U16746 (N_16746,N_16261,N_16131);
and U16747 (N_16747,N_16149,N_16499);
nand U16748 (N_16748,N_16330,N_16156);
nor U16749 (N_16749,N_16070,N_16095);
nor U16750 (N_16750,N_16082,N_16159);
xor U16751 (N_16751,N_16354,N_16378);
xor U16752 (N_16752,N_16360,N_16450);
or U16753 (N_16753,N_16185,N_16454);
xor U16754 (N_16754,N_16296,N_16152);
and U16755 (N_16755,N_16384,N_16293);
and U16756 (N_16756,N_16333,N_16354);
or U16757 (N_16757,N_16033,N_16032);
nand U16758 (N_16758,N_16033,N_16367);
and U16759 (N_16759,N_16401,N_16111);
nor U16760 (N_16760,N_16443,N_16332);
and U16761 (N_16761,N_16142,N_16244);
and U16762 (N_16762,N_16138,N_16244);
or U16763 (N_16763,N_16151,N_16345);
or U16764 (N_16764,N_16248,N_16272);
and U16765 (N_16765,N_16067,N_16044);
xor U16766 (N_16766,N_16073,N_16188);
xnor U16767 (N_16767,N_16029,N_16344);
nor U16768 (N_16768,N_16278,N_16366);
nor U16769 (N_16769,N_16004,N_16284);
or U16770 (N_16770,N_16294,N_16040);
xnor U16771 (N_16771,N_16032,N_16316);
nand U16772 (N_16772,N_16012,N_16163);
or U16773 (N_16773,N_16161,N_16287);
nand U16774 (N_16774,N_16140,N_16387);
or U16775 (N_16775,N_16081,N_16378);
nor U16776 (N_16776,N_16287,N_16372);
or U16777 (N_16777,N_16360,N_16042);
nand U16778 (N_16778,N_16374,N_16072);
nand U16779 (N_16779,N_16240,N_16212);
nor U16780 (N_16780,N_16316,N_16274);
or U16781 (N_16781,N_16063,N_16427);
and U16782 (N_16782,N_16039,N_16370);
and U16783 (N_16783,N_16087,N_16044);
nor U16784 (N_16784,N_16227,N_16426);
nor U16785 (N_16785,N_16433,N_16426);
or U16786 (N_16786,N_16173,N_16339);
nand U16787 (N_16787,N_16019,N_16445);
nand U16788 (N_16788,N_16325,N_16248);
or U16789 (N_16789,N_16301,N_16277);
xnor U16790 (N_16790,N_16218,N_16050);
and U16791 (N_16791,N_16286,N_16403);
xnor U16792 (N_16792,N_16433,N_16288);
or U16793 (N_16793,N_16157,N_16360);
nor U16794 (N_16794,N_16205,N_16422);
and U16795 (N_16795,N_16148,N_16428);
or U16796 (N_16796,N_16278,N_16022);
nor U16797 (N_16797,N_16399,N_16240);
or U16798 (N_16798,N_16304,N_16052);
or U16799 (N_16799,N_16326,N_16123);
nor U16800 (N_16800,N_16228,N_16481);
nand U16801 (N_16801,N_16146,N_16440);
nor U16802 (N_16802,N_16061,N_16143);
nand U16803 (N_16803,N_16140,N_16385);
and U16804 (N_16804,N_16208,N_16440);
xnor U16805 (N_16805,N_16415,N_16153);
or U16806 (N_16806,N_16039,N_16324);
nor U16807 (N_16807,N_16014,N_16366);
and U16808 (N_16808,N_16313,N_16103);
nor U16809 (N_16809,N_16139,N_16051);
nor U16810 (N_16810,N_16256,N_16266);
and U16811 (N_16811,N_16183,N_16006);
nand U16812 (N_16812,N_16257,N_16168);
xor U16813 (N_16813,N_16199,N_16126);
nand U16814 (N_16814,N_16253,N_16109);
nand U16815 (N_16815,N_16287,N_16058);
nand U16816 (N_16816,N_16282,N_16070);
nand U16817 (N_16817,N_16231,N_16244);
xnor U16818 (N_16818,N_16059,N_16182);
or U16819 (N_16819,N_16206,N_16172);
xnor U16820 (N_16820,N_16167,N_16052);
nor U16821 (N_16821,N_16008,N_16260);
and U16822 (N_16822,N_16401,N_16032);
and U16823 (N_16823,N_16161,N_16308);
or U16824 (N_16824,N_16232,N_16466);
nor U16825 (N_16825,N_16267,N_16301);
nand U16826 (N_16826,N_16276,N_16066);
xnor U16827 (N_16827,N_16433,N_16047);
and U16828 (N_16828,N_16264,N_16405);
and U16829 (N_16829,N_16499,N_16026);
nor U16830 (N_16830,N_16135,N_16278);
nor U16831 (N_16831,N_16410,N_16088);
nand U16832 (N_16832,N_16492,N_16263);
nand U16833 (N_16833,N_16122,N_16482);
or U16834 (N_16834,N_16066,N_16087);
nand U16835 (N_16835,N_16034,N_16019);
nand U16836 (N_16836,N_16244,N_16414);
nand U16837 (N_16837,N_16102,N_16312);
nor U16838 (N_16838,N_16065,N_16326);
or U16839 (N_16839,N_16225,N_16033);
nor U16840 (N_16840,N_16461,N_16064);
nor U16841 (N_16841,N_16155,N_16183);
nor U16842 (N_16842,N_16118,N_16053);
nor U16843 (N_16843,N_16311,N_16180);
or U16844 (N_16844,N_16414,N_16451);
and U16845 (N_16845,N_16472,N_16317);
and U16846 (N_16846,N_16462,N_16066);
and U16847 (N_16847,N_16471,N_16383);
xnor U16848 (N_16848,N_16464,N_16344);
nor U16849 (N_16849,N_16280,N_16387);
and U16850 (N_16850,N_16140,N_16166);
nand U16851 (N_16851,N_16343,N_16194);
or U16852 (N_16852,N_16315,N_16286);
nor U16853 (N_16853,N_16031,N_16072);
or U16854 (N_16854,N_16151,N_16361);
and U16855 (N_16855,N_16465,N_16469);
or U16856 (N_16856,N_16396,N_16164);
and U16857 (N_16857,N_16035,N_16366);
nor U16858 (N_16858,N_16308,N_16397);
or U16859 (N_16859,N_16345,N_16199);
xnor U16860 (N_16860,N_16301,N_16060);
xnor U16861 (N_16861,N_16307,N_16187);
and U16862 (N_16862,N_16430,N_16331);
nand U16863 (N_16863,N_16170,N_16410);
or U16864 (N_16864,N_16292,N_16127);
and U16865 (N_16865,N_16141,N_16221);
nand U16866 (N_16866,N_16309,N_16228);
nor U16867 (N_16867,N_16397,N_16008);
or U16868 (N_16868,N_16041,N_16419);
xor U16869 (N_16869,N_16127,N_16158);
or U16870 (N_16870,N_16272,N_16220);
or U16871 (N_16871,N_16054,N_16213);
nor U16872 (N_16872,N_16483,N_16245);
xnor U16873 (N_16873,N_16210,N_16362);
nand U16874 (N_16874,N_16379,N_16440);
nand U16875 (N_16875,N_16347,N_16416);
xor U16876 (N_16876,N_16161,N_16442);
xor U16877 (N_16877,N_16440,N_16325);
nor U16878 (N_16878,N_16449,N_16198);
and U16879 (N_16879,N_16201,N_16463);
and U16880 (N_16880,N_16229,N_16361);
and U16881 (N_16881,N_16194,N_16192);
and U16882 (N_16882,N_16136,N_16408);
nor U16883 (N_16883,N_16374,N_16339);
nand U16884 (N_16884,N_16019,N_16157);
or U16885 (N_16885,N_16406,N_16324);
nand U16886 (N_16886,N_16473,N_16044);
xnor U16887 (N_16887,N_16321,N_16429);
nand U16888 (N_16888,N_16236,N_16231);
nor U16889 (N_16889,N_16456,N_16032);
nand U16890 (N_16890,N_16032,N_16336);
and U16891 (N_16891,N_16125,N_16407);
nor U16892 (N_16892,N_16197,N_16268);
or U16893 (N_16893,N_16306,N_16030);
xor U16894 (N_16894,N_16166,N_16003);
and U16895 (N_16895,N_16481,N_16016);
nand U16896 (N_16896,N_16406,N_16160);
or U16897 (N_16897,N_16147,N_16058);
and U16898 (N_16898,N_16197,N_16096);
and U16899 (N_16899,N_16039,N_16049);
nand U16900 (N_16900,N_16451,N_16205);
or U16901 (N_16901,N_16392,N_16059);
nand U16902 (N_16902,N_16155,N_16018);
xnor U16903 (N_16903,N_16336,N_16414);
nor U16904 (N_16904,N_16105,N_16270);
nor U16905 (N_16905,N_16123,N_16150);
and U16906 (N_16906,N_16430,N_16204);
nand U16907 (N_16907,N_16388,N_16363);
nor U16908 (N_16908,N_16218,N_16467);
and U16909 (N_16909,N_16083,N_16044);
nor U16910 (N_16910,N_16308,N_16050);
xor U16911 (N_16911,N_16219,N_16056);
nor U16912 (N_16912,N_16346,N_16377);
and U16913 (N_16913,N_16304,N_16144);
or U16914 (N_16914,N_16485,N_16451);
nor U16915 (N_16915,N_16236,N_16106);
or U16916 (N_16916,N_16175,N_16351);
nand U16917 (N_16917,N_16111,N_16166);
nor U16918 (N_16918,N_16314,N_16100);
or U16919 (N_16919,N_16468,N_16186);
xor U16920 (N_16920,N_16150,N_16395);
nor U16921 (N_16921,N_16089,N_16192);
xor U16922 (N_16922,N_16116,N_16180);
or U16923 (N_16923,N_16280,N_16452);
or U16924 (N_16924,N_16011,N_16432);
and U16925 (N_16925,N_16182,N_16262);
and U16926 (N_16926,N_16185,N_16041);
xnor U16927 (N_16927,N_16451,N_16105);
nor U16928 (N_16928,N_16361,N_16421);
or U16929 (N_16929,N_16022,N_16156);
or U16930 (N_16930,N_16238,N_16365);
nand U16931 (N_16931,N_16461,N_16342);
nand U16932 (N_16932,N_16094,N_16476);
xor U16933 (N_16933,N_16153,N_16207);
nand U16934 (N_16934,N_16380,N_16217);
nand U16935 (N_16935,N_16418,N_16298);
xnor U16936 (N_16936,N_16310,N_16338);
nor U16937 (N_16937,N_16031,N_16020);
nand U16938 (N_16938,N_16200,N_16352);
and U16939 (N_16939,N_16099,N_16465);
nand U16940 (N_16940,N_16371,N_16324);
nand U16941 (N_16941,N_16362,N_16048);
nor U16942 (N_16942,N_16237,N_16083);
xnor U16943 (N_16943,N_16471,N_16265);
nand U16944 (N_16944,N_16127,N_16018);
nor U16945 (N_16945,N_16418,N_16237);
nor U16946 (N_16946,N_16267,N_16282);
and U16947 (N_16947,N_16280,N_16300);
nor U16948 (N_16948,N_16419,N_16345);
or U16949 (N_16949,N_16287,N_16131);
and U16950 (N_16950,N_16166,N_16334);
nor U16951 (N_16951,N_16121,N_16216);
or U16952 (N_16952,N_16495,N_16145);
nor U16953 (N_16953,N_16380,N_16020);
nand U16954 (N_16954,N_16253,N_16035);
and U16955 (N_16955,N_16457,N_16185);
and U16956 (N_16956,N_16450,N_16185);
xor U16957 (N_16957,N_16187,N_16009);
nor U16958 (N_16958,N_16104,N_16217);
xor U16959 (N_16959,N_16384,N_16486);
nand U16960 (N_16960,N_16433,N_16137);
xnor U16961 (N_16961,N_16201,N_16017);
nor U16962 (N_16962,N_16043,N_16323);
nand U16963 (N_16963,N_16368,N_16077);
nand U16964 (N_16964,N_16404,N_16245);
xnor U16965 (N_16965,N_16165,N_16036);
nor U16966 (N_16966,N_16428,N_16059);
xor U16967 (N_16967,N_16002,N_16245);
nor U16968 (N_16968,N_16320,N_16156);
and U16969 (N_16969,N_16063,N_16219);
nor U16970 (N_16970,N_16297,N_16262);
and U16971 (N_16971,N_16022,N_16428);
or U16972 (N_16972,N_16056,N_16492);
and U16973 (N_16973,N_16160,N_16072);
or U16974 (N_16974,N_16485,N_16004);
nor U16975 (N_16975,N_16118,N_16009);
or U16976 (N_16976,N_16407,N_16073);
or U16977 (N_16977,N_16368,N_16441);
and U16978 (N_16978,N_16336,N_16299);
or U16979 (N_16979,N_16137,N_16172);
and U16980 (N_16980,N_16425,N_16243);
xor U16981 (N_16981,N_16441,N_16178);
nand U16982 (N_16982,N_16032,N_16125);
xor U16983 (N_16983,N_16182,N_16285);
or U16984 (N_16984,N_16070,N_16002);
or U16985 (N_16985,N_16219,N_16459);
or U16986 (N_16986,N_16152,N_16379);
nor U16987 (N_16987,N_16019,N_16479);
and U16988 (N_16988,N_16486,N_16284);
and U16989 (N_16989,N_16079,N_16152);
or U16990 (N_16990,N_16214,N_16047);
xor U16991 (N_16991,N_16207,N_16267);
nor U16992 (N_16992,N_16235,N_16012);
nor U16993 (N_16993,N_16422,N_16387);
and U16994 (N_16994,N_16407,N_16173);
nand U16995 (N_16995,N_16080,N_16231);
or U16996 (N_16996,N_16218,N_16286);
nand U16997 (N_16997,N_16078,N_16470);
nand U16998 (N_16998,N_16362,N_16255);
or U16999 (N_16999,N_16490,N_16228);
xnor U17000 (N_17000,N_16516,N_16717);
and U17001 (N_17001,N_16513,N_16512);
xnor U17002 (N_17002,N_16703,N_16839);
nor U17003 (N_17003,N_16600,N_16992);
xor U17004 (N_17004,N_16594,N_16850);
and U17005 (N_17005,N_16599,N_16862);
and U17006 (N_17006,N_16515,N_16987);
and U17007 (N_17007,N_16748,N_16627);
nand U17008 (N_17008,N_16571,N_16651);
nand U17009 (N_17009,N_16903,N_16995);
xor U17010 (N_17010,N_16573,N_16674);
xor U17011 (N_17011,N_16920,N_16980);
or U17012 (N_17012,N_16560,N_16940);
or U17013 (N_17013,N_16741,N_16527);
nand U17014 (N_17014,N_16583,N_16590);
and U17015 (N_17015,N_16691,N_16952);
and U17016 (N_17016,N_16774,N_16927);
or U17017 (N_17017,N_16928,N_16668);
nor U17018 (N_17018,N_16563,N_16705);
xor U17019 (N_17019,N_16861,N_16756);
nor U17020 (N_17020,N_16575,N_16738);
and U17021 (N_17021,N_16647,N_16589);
xor U17022 (N_17022,N_16798,N_16742);
and U17023 (N_17023,N_16879,N_16949);
xor U17024 (N_17024,N_16853,N_16823);
or U17025 (N_17025,N_16848,N_16921);
nor U17026 (N_17026,N_16506,N_16947);
xnor U17027 (N_17027,N_16704,N_16818);
and U17028 (N_17028,N_16795,N_16731);
nor U17029 (N_17029,N_16548,N_16523);
nand U17030 (N_17030,N_16669,N_16915);
nor U17031 (N_17031,N_16779,N_16721);
and U17032 (N_17032,N_16865,N_16736);
nand U17033 (N_17033,N_16863,N_16544);
nor U17034 (N_17034,N_16812,N_16733);
nor U17035 (N_17035,N_16874,N_16724);
or U17036 (N_17036,N_16632,N_16664);
xor U17037 (N_17037,N_16752,N_16609);
xnor U17038 (N_17038,N_16744,N_16730);
and U17039 (N_17039,N_16893,N_16936);
and U17040 (N_17040,N_16579,N_16914);
or U17041 (N_17041,N_16830,N_16526);
and U17042 (N_17042,N_16710,N_16518);
xnor U17043 (N_17043,N_16747,N_16755);
xnor U17044 (N_17044,N_16801,N_16842);
or U17045 (N_17045,N_16760,N_16775);
and U17046 (N_17046,N_16826,N_16807);
and U17047 (N_17047,N_16790,N_16846);
xor U17048 (N_17048,N_16750,N_16935);
nor U17049 (N_17049,N_16726,N_16567);
and U17050 (N_17050,N_16532,N_16625);
or U17051 (N_17051,N_16644,N_16765);
xor U17052 (N_17052,N_16581,N_16964);
and U17053 (N_17053,N_16822,N_16725);
nor U17054 (N_17054,N_16708,N_16965);
nand U17055 (N_17055,N_16957,N_16661);
nor U17056 (N_17056,N_16628,N_16656);
nor U17057 (N_17057,N_16783,N_16597);
and U17058 (N_17058,N_16536,N_16706);
or U17059 (N_17059,N_16740,N_16638);
and U17060 (N_17060,N_16714,N_16685);
nand U17061 (N_17061,N_16552,N_16892);
nand U17062 (N_17062,N_16593,N_16819);
nor U17063 (N_17063,N_16547,N_16860);
xor U17064 (N_17064,N_16829,N_16529);
or U17065 (N_17065,N_16806,N_16718);
xnor U17066 (N_17066,N_16524,N_16680);
xnor U17067 (N_17067,N_16663,N_16553);
or U17068 (N_17068,N_16734,N_16886);
and U17069 (N_17069,N_16654,N_16635);
nor U17070 (N_17070,N_16944,N_16859);
and U17071 (N_17071,N_16699,N_16780);
nor U17072 (N_17072,N_16700,N_16771);
and U17073 (N_17073,N_16557,N_16649);
and U17074 (N_17074,N_16981,N_16803);
or U17075 (N_17075,N_16875,N_16993);
and U17076 (N_17076,N_16962,N_16520);
nor U17077 (N_17077,N_16569,N_16809);
xnor U17078 (N_17078,N_16847,N_16891);
xnor U17079 (N_17079,N_16501,N_16813);
xnor U17080 (N_17080,N_16528,N_16757);
nor U17081 (N_17081,N_16802,N_16565);
xnor U17082 (N_17082,N_16785,N_16979);
xnor U17083 (N_17083,N_16507,N_16837);
nor U17084 (N_17084,N_16831,N_16530);
xor U17085 (N_17085,N_16960,N_16838);
xor U17086 (N_17086,N_16881,N_16811);
nand U17087 (N_17087,N_16580,N_16919);
and U17088 (N_17088,N_16642,N_16986);
or U17089 (N_17089,N_16946,N_16677);
nor U17090 (N_17090,N_16727,N_16540);
or U17091 (N_17091,N_16994,N_16671);
nor U17092 (N_17092,N_16998,N_16984);
and U17093 (N_17093,N_16871,N_16667);
or U17094 (N_17094,N_16989,N_16604);
and U17095 (N_17095,N_16963,N_16917);
and U17096 (N_17096,N_16766,N_16894);
nor U17097 (N_17097,N_16522,N_16770);
and U17098 (N_17098,N_16603,N_16923);
nand U17099 (N_17099,N_16617,N_16611);
nand U17100 (N_17100,N_16525,N_16550);
nor U17101 (N_17101,N_16556,N_16999);
nor U17102 (N_17102,N_16519,N_16678);
and U17103 (N_17103,N_16626,N_16559);
and U17104 (N_17104,N_16913,N_16799);
nor U17105 (N_17105,N_16896,N_16841);
nand U17106 (N_17106,N_16679,N_16897);
xor U17107 (N_17107,N_16648,N_16665);
or U17108 (N_17108,N_16856,N_16977);
xor U17109 (N_17109,N_16728,N_16618);
nand U17110 (N_17110,N_16814,N_16932);
and U17111 (N_17111,N_16909,N_16619);
nand U17112 (N_17112,N_16595,N_16773);
and U17113 (N_17113,N_16585,N_16630);
or U17114 (N_17114,N_16890,N_16908);
nand U17115 (N_17115,N_16701,N_16531);
nor U17116 (N_17116,N_16845,N_16514);
xnor U17117 (N_17117,N_16966,N_16997);
xnor U17118 (N_17118,N_16614,N_16953);
nand U17119 (N_17119,N_16810,N_16608);
and U17120 (N_17120,N_16688,N_16554);
xnor U17121 (N_17121,N_16786,N_16695);
or U17122 (N_17122,N_16690,N_16922);
nor U17123 (N_17123,N_16538,N_16500);
or U17124 (N_17124,N_16884,N_16777);
or U17125 (N_17125,N_16869,N_16711);
or U17126 (N_17126,N_16693,N_16729);
xnor U17127 (N_17127,N_16877,N_16954);
nand U17128 (N_17128,N_16645,N_16990);
nand U17129 (N_17129,N_16702,N_16673);
nand U17130 (N_17130,N_16732,N_16503);
nor U17131 (N_17131,N_16942,N_16885);
nor U17132 (N_17132,N_16991,N_16937);
or U17133 (N_17133,N_16696,N_16967);
nand U17134 (N_17134,N_16910,N_16720);
nor U17135 (N_17135,N_16817,N_16776);
xnor U17136 (N_17136,N_16956,N_16623);
or U17137 (N_17137,N_16639,N_16534);
nor U17138 (N_17138,N_16689,N_16598);
or U17139 (N_17139,N_16660,N_16983);
nand U17140 (N_17140,N_16939,N_16912);
nor U17141 (N_17141,N_16542,N_16615);
nor U17142 (N_17142,N_16739,N_16653);
or U17143 (N_17143,N_16607,N_16904);
xor U17144 (N_17144,N_16535,N_16658);
or U17145 (N_17145,N_16588,N_16576);
and U17146 (N_17146,N_16652,N_16521);
xnor U17147 (N_17147,N_16517,N_16873);
or U17148 (N_17148,N_16895,N_16888);
nor U17149 (N_17149,N_16754,N_16722);
or U17150 (N_17150,N_16832,N_16707);
xor U17151 (N_17151,N_16792,N_16577);
xnor U17152 (N_17152,N_16629,N_16950);
nor U17153 (N_17153,N_16636,N_16836);
and U17154 (N_17154,N_16620,N_16541);
xor U17155 (N_17155,N_16545,N_16929);
nand U17156 (N_17156,N_16827,N_16723);
or U17157 (N_17157,N_16948,N_16835);
nand U17158 (N_17158,N_16586,N_16681);
nand U17159 (N_17159,N_16610,N_16650);
and U17160 (N_17160,N_16591,N_16737);
and U17161 (N_17161,N_16602,N_16976);
or U17162 (N_17162,N_16505,N_16854);
nor U17163 (N_17163,N_16851,N_16933);
nand U17164 (N_17164,N_16713,N_16974);
and U17165 (N_17165,N_16684,N_16878);
nor U17166 (N_17166,N_16622,N_16788);
nor U17167 (N_17167,N_16631,N_16924);
nor U17168 (N_17168,N_16662,N_16901);
nand U17169 (N_17169,N_16815,N_16709);
or U17170 (N_17170,N_16975,N_16555);
and U17171 (N_17171,N_16973,N_16943);
xor U17172 (N_17172,N_16772,N_16659);
nand U17173 (N_17173,N_16880,N_16969);
nor U17174 (N_17174,N_16930,N_16504);
nand U17175 (N_17175,N_16562,N_16778);
nand U17176 (N_17176,N_16761,N_16561);
xnor U17177 (N_17177,N_16682,N_16925);
and U17178 (N_17178,N_16820,N_16612);
nor U17179 (N_17179,N_16646,N_16551);
nand U17180 (N_17180,N_16934,N_16511);
nand U17181 (N_17181,N_16574,N_16872);
xnor U17182 (N_17182,N_16749,N_16634);
or U17183 (N_17183,N_16971,N_16857);
or U17184 (N_17184,N_16905,N_16849);
nand U17185 (N_17185,N_16712,N_16697);
or U17186 (N_17186,N_16694,N_16655);
and U17187 (N_17187,N_16794,N_16916);
or U17188 (N_17188,N_16868,N_16791);
or U17189 (N_17189,N_16537,N_16751);
nor U17190 (N_17190,N_16686,N_16633);
or U17191 (N_17191,N_16762,N_16596);
nor U17192 (N_17192,N_16666,N_16787);
nor U17193 (N_17193,N_16675,N_16758);
and U17194 (N_17194,N_16564,N_16978);
xnor U17195 (N_17195,N_16745,N_16808);
xor U17196 (N_17196,N_16961,N_16692);
xnor U17197 (N_17197,N_16796,N_16546);
and U17198 (N_17198,N_16855,N_16870);
nor U17199 (N_17199,N_16889,N_16719);
and U17200 (N_17200,N_16882,N_16907);
xor U17201 (N_17201,N_16698,N_16570);
nor U17202 (N_17202,N_16789,N_16938);
nand U17203 (N_17203,N_16970,N_16784);
and U17204 (N_17204,N_16804,N_16985);
nand U17205 (N_17205,N_16509,N_16670);
xor U17206 (N_17206,N_16828,N_16735);
nor U17207 (N_17207,N_16781,N_16996);
and U17208 (N_17208,N_16605,N_16844);
or U17209 (N_17209,N_16959,N_16683);
nor U17210 (N_17210,N_16763,N_16926);
nor U17211 (N_17211,N_16825,N_16621);
and U17212 (N_17212,N_16899,N_16508);
nand U17213 (N_17213,N_16616,N_16968);
or U17214 (N_17214,N_16782,N_16902);
and U17215 (N_17215,N_16955,N_16867);
and U17216 (N_17216,N_16643,N_16864);
and U17217 (N_17217,N_16941,N_16641);
and U17218 (N_17218,N_16900,N_16833);
or U17219 (N_17219,N_16716,N_16587);
xnor U17220 (N_17220,N_16797,N_16876);
or U17221 (N_17221,N_16906,N_16793);
nor U17222 (N_17222,N_16988,N_16606);
and U17223 (N_17223,N_16840,N_16637);
nand U17224 (N_17224,N_16753,N_16918);
nand U17225 (N_17225,N_16582,N_16613);
xor U17226 (N_17226,N_16805,N_16767);
xor U17227 (N_17227,N_16672,N_16566);
and U17228 (N_17228,N_16768,N_16746);
nand U17229 (N_17229,N_16657,N_16624);
and U17230 (N_17230,N_16800,N_16887);
nor U17231 (N_17231,N_16549,N_16568);
or U17232 (N_17232,N_16982,N_16945);
nor U17233 (N_17233,N_16824,N_16584);
and U17234 (N_17234,N_16502,N_16578);
xor U17235 (N_17235,N_16510,N_16676);
and U17236 (N_17236,N_16866,N_16834);
nor U17237 (N_17237,N_16931,N_16539);
nand U17238 (N_17238,N_16592,N_16715);
nor U17239 (N_17239,N_16543,N_16601);
and U17240 (N_17240,N_16743,N_16951);
or U17241 (N_17241,N_16821,N_16958);
nand U17242 (N_17242,N_16759,N_16858);
nor U17243 (N_17243,N_16572,N_16764);
xor U17244 (N_17244,N_16533,N_16640);
nor U17245 (N_17245,N_16911,N_16972);
or U17246 (N_17246,N_16687,N_16883);
nand U17247 (N_17247,N_16852,N_16898);
nor U17248 (N_17248,N_16558,N_16769);
nor U17249 (N_17249,N_16816,N_16843);
xor U17250 (N_17250,N_16500,N_16530);
or U17251 (N_17251,N_16723,N_16572);
nand U17252 (N_17252,N_16599,N_16559);
nand U17253 (N_17253,N_16523,N_16914);
xor U17254 (N_17254,N_16535,N_16854);
or U17255 (N_17255,N_16893,N_16840);
xnor U17256 (N_17256,N_16971,N_16920);
nand U17257 (N_17257,N_16582,N_16873);
xnor U17258 (N_17258,N_16699,N_16525);
nor U17259 (N_17259,N_16770,N_16500);
nand U17260 (N_17260,N_16619,N_16989);
or U17261 (N_17261,N_16925,N_16647);
nor U17262 (N_17262,N_16634,N_16666);
or U17263 (N_17263,N_16982,N_16709);
and U17264 (N_17264,N_16943,N_16749);
or U17265 (N_17265,N_16609,N_16718);
and U17266 (N_17266,N_16794,N_16686);
nand U17267 (N_17267,N_16982,N_16882);
xor U17268 (N_17268,N_16527,N_16803);
xnor U17269 (N_17269,N_16701,N_16761);
nand U17270 (N_17270,N_16854,N_16718);
nand U17271 (N_17271,N_16745,N_16977);
or U17272 (N_17272,N_16710,N_16771);
and U17273 (N_17273,N_16548,N_16856);
nand U17274 (N_17274,N_16718,N_16735);
nand U17275 (N_17275,N_16661,N_16821);
nor U17276 (N_17276,N_16765,N_16983);
nor U17277 (N_17277,N_16941,N_16517);
or U17278 (N_17278,N_16501,N_16998);
or U17279 (N_17279,N_16676,N_16569);
nand U17280 (N_17280,N_16700,N_16558);
nand U17281 (N_17281,N_16554,N_16972);
or U17282 (N_17282,N_16633,N_16552);
or U17283 (N_17283,N_16708,N_16580);
nand U17284 (N_17284,N_16755,N_16882);
nor U17285 (N_17285,N_16911,N_16770);
or U17286 (N_17286,N_16916,N_16533);
xor U17287 (N_17287,N_16966,N_16836);
or U17288 (N_17288,N_16701,N_16512);
or U17289 (N_17289,N_16781,N_16934);
xor U17290 (N_17290,N_16766,N_16703);
or U17291 (N_17291,N_16619,N_16720);
xor U17292 (N_17292,N_16502,N_16787);
and U17293 (N_17293,N_16571,N_16959);
nor U17294 (N_17294,N_16862,N_16556);
or U17295 (N_17295,N_16665,N_16535);
nand U17296 (N_17296,N_16717,N_16690);
and U17297 (N_17297,N_16795,N_16593);
xnor U17298 (N_17298,N_16873,N_16733);
nor U17299 (N_17299,N_16957,N_16701);
nand U17300 (N_17300,N_16989,N_16739);
xnor U17301 (N_17301,N_16554,N_16609);
nand U17302 (N_17302,N_16623,N_16782);
xnor U17303 (N_17303,N_16627,N_16895);
or U17304 (N_17304,N_16514,N_16743);
nor U17305 (N_17305,N_16661,N_16798);
nor U17306 (N_17306,N_16532,N_16952);
and U17307 (N_17307,N_16655,N_16892);
nor U17308 (N_17308,N_16517,N_16847);
nor U17309 (N_17309,N_16579,N_16939);
nand U17310 (N_17310,N_16713,N_16719);
nor U17311 (N_17311,N_16930,N_16918);
and U17312 (N_17312,N_16570,N_16890);
xnor U17313 (N_17313,N_16972,N_16543);
and U17314 (N_17314,N_16692,N_16899);
or U17315 (N_17315,N_16527,N_16827);
nand U17316 (N_17316,N_16591,N_16943);
xor U17317 (N_17317,N_16535,N_16943);
xnor U17318 (N_17318,N_16943,N_16779);
or U17319 (N_17319,N_16908,N_16677);
nand U17320 (N_17320,N_16965,N_16657);
xor U17321 (N_17321,N_16659,N_16978);
or U17322 (N_17322,N_16766,N_16780);
nor U17323 (N_17323,N_16713,N_16852);
nand U17324 (N_17324,N_16829,N_16790);
and U17325 (N_17325,N_16979,N_16638);
nand U17326 (N_17326,N_16868,N_16758);
nor U17327 (N_17327,N_16530,N_16979);
or U17328 (N_17328,N_16998,N_16806);
nor U17329 (N_17329,N_16978,N_16555);
xnor U17330 (N_17330,N_16928,N_16548);
and U17331 (N_17331,N_16826,N_16975);
xnor U17332 (N_17332,N_16500,N_16667);
xor U17333 (N_17333,N_16879,N_16986);
and U17334 (N_17334,N_16511,N_16532);
or U17335 (N_17335,N_16647,N_16882);
nor U17336 (N_17336,N_16991,N_16883);
and U17337 (N_17337,N_16707,N_16782);
xor U17338 (N_17338,N_16850,N_16730);
nand U17339 (N_17339,N_16825,N_16585);
or U17340 (N_17340,N_16673,N_16796);
xor U17341 (N_17341,N_16760,N_16668);
nand U17342 (N_17342,N_16642,N_16860);
nor U17343 (N_17343,N_16763,N_16876);
or U17344 (N_17344,N_16541,N_16785);
or U17345 (N_17345,N_16658,N_16732);
xor U17346 (N_17346,N_16640,N_16732);
or U17347 (N_17347,N_16893,N_16548);
xnor U17348 (N_17348,N_16565,N_16931);
nor U17349 (N_17349,N_16746,N_16773);
nand U17350 (N_17350,N_16565,N_16870);
and U17351 (N_17351,N_16895,N_16659);
and U17352 (N_17352,N_16965,N_16537);
or U17353 (N_17353,N_16867,N_16670);
nand U17354 (N_17354,N_16565,N_16614);
nor U17355 (N_17355,N_16761,N_16784);
nor U17356 (N_17356,N_16910,N_16968);
or U17357 (N_17357,N_16940,N_16744);
xnor U17358 (N_17358,N_16986,N_16717);
nor U17359 (N_17359,N_16755,N_16647);
or U17360 (N_17360,N_16903,N_16561);
xor U17361 (N_17361,N_16518,N_16804);
or U17362 (N_17362,N_16872,N_16772);
nor U17363 (N_17363,N_16769,N_16544);
xnor U17364 (N_17364,N_16740,N_16672);
and U17365 (N_17365,N_16698,N_16660);
xnor U17366 (N_17366,N_16702,N_16740);
or U17367 (N_17367,N_16644,N_16540);
nand U17368 (N_17368,N_16672,N_16598);
nand U17369 (N_17369,N_16512,N_16807);
or U17370 (N_17370,N_16748,N_16967);
and U17371 (N_17371,N_16852,N_16748);
xnor U17372 (N_17372,N_16936,N_16755);
xor U17373 (N_17373,N_16828,N_16914);
and U17374 (N_17374,N_16812,N_16757);
or U17375 (N_17375,N_16549,N_16636);
xnor U17376 (N_17376,N_16566,N_16645);
xnor U17377 (N_17377,N_16654,N_16988);
nor U17378 (N_17378,N_16872,N_16609);
nand U17379 (N_17379,N_16873,N_16995);
and U17380 (N_17380,N_16950,N_16843);
nand U17381 (N_17381,N_16975,N_16547);
nand U17382 (N_17382,N_16668,N_16639);
nor U17383 (N_17383,N_16578,N_16746);
and U17384 (N_17384,N_16504,N_16597);
nand U17385 (N_17385,N_16560,N_16652);
nand U17386 (N_17386,N_16582,N_16931);
or U17387 (N_17387,N_16974,N_16610);
nor U17388 (N_17388,N_16861,N_16874);
nand U17389 (N_17389,N_16595,N_16548);
or U17390 (N_17390,N_16587,N_16828);
xnor U17391 (N_17391,N_16510,N_16541);
nor U17392 (N_17392,N_16957,N_16729);
or U17393 (N_17393,N_16883,N_16542);
xnor U17394 (N_17394,N_16944,N_16851);
xor U17395 (N_17395,N_16900,N_16981);
nor U17396 (N_17396,N_16972,N_16722);
nand U17397 (N_17397,N_16566,N_16798);
and U17398 (N_17398,N_16928,N_16955);
nand U17399 (N_17399,N_16675,N_16763);
or U17400 (N_17400,N_16512,N_16574);
nand U17401 (N_17401,N_16881,N_16798);
or U17402 (N_17402,N_16568,N_16983);
nor U17403 (N_17403,N_16533,N_16701);
or U17404 (N_17404,N_16842,N_16675);
and U17405 (N_17405,N_16653,N_16957);
xnor U17406 (N_17406,N_16883,N_16696);
and U17407 (N_17407,N_16912,N_16763);
and U17408 (N_17408,N_16580,N_16798);
and U17409 (N_17409,N_16805,N_16525);
and U17410 (N_17410,N_16666,N_16629);
and U17411 (N_17411,N_16685,N_16852);
xor U17412 (N_17412,N_16881,N_16610);
or U17413 (N_17413,N_16811,N_16564);
or U17414 (N_17414,N_16885,N_16894);
nor U17415 (N_17415,N_16606,N_16925);
or U17416 (N_17416,N_16555,N_16657);
nor U17417 (N_17417,N_16556,N_16838);
nand U17418 (N_17418,N_16628,N_16813);
nand U17419 (N_17419,N_16905,N_16688);
xnor U17420 (N_17420,N_16863,N_16859);
xor U17421 (N_17421,N_16896,N_16826);
or U17422 (N_17422,N_16801,N_16522);
nor U17423 (N_17423,N_16762,N_16946);
and U17424 (N_17424,N_16775,N_16705);
xor U17425 (N_17425,N_16941,N_16657);
or U17426 (N_17426,N_16646,N_16979);
xor U17427 (N_17427,N_16652,N_16573);
nand U17428 (N_17428,N_16868,N_16811);
and U17429 (N_17429,N_16674,N_16908);
xnor U17430 (N_17430,N_16735,N_16628);
nand U17431 (N_17431,N_16542,N_16963);
or U17432 (N_17432,N_16591,N_16868);
and U17433 (N_17433,N_16579,N_16892);
or U17434 (N_17434,N_16768,N_16848);
or U17435 (N_17435,N_16926,N_16893);
nand U17436 (N_17436,N_16963,N_16629);
nor U17437 (N_17437,N_16869,N_16873);
nor U17438 (N_17438,N_16890,N_16764);
or U17439 (N_17439,N_16753,N_16681);
nor U17440 (N_17440,N_16952,N_16511);
xnor U17441 (N_17441,N_16693,N_16586);
nor U17442 (N_17442,N_16683,N_16719);
xor U17443 (N_17443,N_16930,N_16605);
or U17444 (N_17444,N_16721,N_16656);
and U17445 (N_17445,N_16937,N_16634);
nor U17446 (N_17446,N_16762,N_16520);
or U17447 (N_17447,N_16889,N_16526);
and U17448 (N_17448,N_16849,N_16755);
and U17449 (N_17449,N_16651,N_16915);
or U17450 (N_17450,N_16865,N_16854);
or U17451 (N_17451,N_16717,N_16736);
nor U17452 (N_17452,N_16773,N_16779);
nor U17453 (N_17453,N_16922,N_16638);
or U17454 (N_17454,N_16972,N_16676);
nor U17455 (N_17455,N_16562,N_16727);
nor U17456 (N_17456,N_16937,N_16528);
nand U17457 (N_17457,N_16677,N_16575);
xnor U17458 (N_17458,N_16566,N_16660);
nand U17459 (N_17459,N_16819,N_16705);
or U17460 (N_17460,N_16712,N_16846);
or U17461 (N_17461,N_16770,N_16607);
xor U17462 (N_17462,N_16523,N_16964);
or U17463 (N_17463,N_16558,N_16762);
or U17464 (N_17464,N_16916,N_16570);
and U17465 (N_17465,N_16839,N_16637);
or U17466 (N_17466,N_16804,N_16919);
or U17467 (N_17467,N_16909,N_16693);
xor U17468 (N_17468,N_16599,N_16631);
and U17469 (N_17469,N_16885,N_16611);
or U17470 (N_17470,N_16834,N_16698);
xor U17471 (N_17471,N_16924,N_16927);
xnor U17472 (N_17472,N_16841,N_16801);
or U17473 (N_17473,N_16683,N_16956);
nand U17474 (N_17474,N_16793,N_16996);
nand U17475 (N_17475,N_16552,N_16538);
and U17476 (N_17476,N_16983,N_16514);
or U17477 (N_17477,N_16939,N_16943);
and U17478 (N_17478,N_16735,N_16507);
xnor U17479 (N_17479,N_16523,N_16640);
nor U17480 (N_17480,N_16590,N_16502);
xnor U17481 (N_17481,N_16917,N_16905);
nor U17482 (N_17482,N_16709,N_16809);
nand U17483 (N_17483,N_16816,N_16565);
nor U17484 (N_17484,N_16619,N_16788);
nor U17485 (N_17485,N_16732,N_16834);
nor U17486 (N_17486,N_16718,N_16900);
and U17487 (N_17487,N_16866,N_16651);
xor U17488 (N_17488,N_16690,N_16839);
nand U17489 (N_17489,N_16656,N_16793);
nand U17490 (N_17490,N_16636,N_16645);
and U17491 (N_17491,N_16702,N_16813);
xor U17492 (N_17492,N_16551,N_16846);
xnor U17493 (N_17493,N_16854,N_16526);
or U17494 (N_17494,N_16620,N_16835);
nand U17495 (N_17495,N_16940,N_16534);
or U17496 (N_17496,N_16511,N_16641);
nor U17497 (N_17497,N_16705,N_16807);
nor U17498 (N_17498,N_16815,N_16929);
nor U17499 (N_17499,N_16767,N_16970);
or U17500 (N_17500,N_17063,N_17113);
xor U17501 (N_17501,N_17313,N_17333);
nor U17502 (N_17502,N_17420,N_17261);
and U17503 (N_17503,N_17152,N_17303);
or U17504 (N_17504,N_17344,N_17453);
nand U17505 (N_17505,N_17112,N_17406);
nor U17506 (N_17506,N_17330,N_17416);
nor U17507 (N_17507,N_17194,N_17157);
and U17508 (N_17508,N_17155,N_17383);
xor U17509 (N_17509,N_17286,N_17297);
nor U17510 (N_17510,N_17396,N_17408);
or U17511 (N_17511,N_17473,N_17296);
nand U17512 (N_17512,N_17096,N_17186);
and U17513 (N_17513,N_17445,N_17026);
xor U17514 (N_17514,N_17211,N_17485);
and U17515 (N_17515,N_17311,N_17031);
nor U17516 (N_17516,N_17334,N_17200);
xor U17517 (N_17517,N_17110,N_17141);
and U17518 (N_17518,N_17381,N_17189);
and U17519 (N_17519,N_17405,N_17162);
nand U17520 (N_17520,N_17387,N_17235);
nand U17521 (N_17521,N_17010,N_17125);
nand U17522 (N_17522,N_17439,N_17429);
and U17523 (N_17523,N_17321,N_17305);
or U17524 (N_17524,N_17496,N_17274);
nand U17525 (N_17525,N_17413,N_17434);
xnor U17526 (N_17526,N_17066,N_17092);
or U17527 (N_17527,N_17053,N_17234);
and U17528 (N_17528,N_17067,N_17227);
xor U17529 (N_17529,N_17102,N_17213);
or U17530 (N_17530,N_17204,N_17124);
or U17531 (N_17531,N_17498,N_17254);
nor U17532 (N_17532,N_17368,N_17298);
and U17533 (N_17533,N_17436,N_17058);
xnor U17534 (N_17534,N_17041,N_17217);
and U17535 (N_17535,N_17414,N_17143);
nor U17536 (N_17536,N_17159,N_17009);
nand U17537 (N_17537,N_17250,N_17246);
xor U17538 (N_17538,N_17499,N_17376);
and U17539 (N_17539,N_17397,N_17410);
nand U17540 (N_17540,N_17449,N_17271);
xnor U17541 (N_17541,N_17139,N_17277);
and U17542 (N_17542,N_17367,N_17335);
and U17543 (N_17543,N_17458,N_17479);
or U17544 (N_17544,N_17299,N_17034);
and U17545 (N_17545,N_17273,N_17431);
nand U17546 (N_17546,N_17459,N_17422);
and U17547 (N_17547,N_17080,N_17384);
nand U17548 (N_17548,N_17400,N_17042);
and U17549 (N_17549,N_17475,N_17267);
and U17550 (N_17550,N_17046,N_17259);
or U17551 (N_17551,N_17021,N_17471);
and U17552 (N_17552,N_17202,N_17360);
and U17553 (N_17553,N_17435,N_17399);
and U17554 (N_17554,N_17131,N_17354);
nand U17555 (N_17555,N_17094,N_17145);
or U17556 (N_17556,N_17364,N_17411);
nor U17557 (N_17557,N_17044,N_17095);
nand U17558 (N_17558,N_17295,N_17476);
or U17559 (N_17559,N_17231,N_17243);
or U17560 (N_17560,N_17291,N_17062);
or U17561 (N_17561,N_17266,N_17276);
nand U17562 (N_17562,N_17222,N_17149);
xor U17563 (N_17563,N_17448,N_17494);
xor U17564 (N_17564,N_17275,N_17389);
or U17565 (N_17565,N_17347,N_17158);
nor U17566 (N_17566,N_17433,N_17392);
nor U17567 (N_17567,N_17385,N_17008);
nand U17568 (N_17568,N_17047,N_17309);
nor U17569 (N_17569,N_17190,N_17412);
and U17570 (N_17570,N_17418,N_17083);
xnor U17571 (N_17571,N_17324,N_17358);
nor U17572 (N_17572,N_17055,N_17417);
nor U17573 (N_17573,N_17051,N_17123);
nor U17574 (N_17574,N_17028,N_17444);
nor U17575 (N_17575,N_17315,N_17178);
or U17576 (N_17576,N_17089,N_17341);
or U17577 (N_17577,N_17151,N_17415);
or U17578 (N_17578,N_17081,N_17164);
nand U17579 (N_17579,N_17279,N_17263);
or U17580 (N_17580,N_17201,N_17161);
nand U17581 (N_17581,N_17441,N_17362);
and U17582 (N_17582,N_17181,N_17015);
nand U17583 (N_17583,N_17116,N_17253);
nand U17584 (N_17584,N_17338,N_17019);
and U17585 (N_17585,N_17280,N_17477);
or U17586 (N_17586,N_17265,N_17101);
nor U17587 (N_17587,N_17233,N_17013);
xnor U17588 (N_17588,N_17097,N_17005);
nor U17589 (N_17589,N_17314,N_17264);
xor U17590 (N_17590,N_17322,N_17136);
and U17591 (N_17591,N_17069,N_17029);
nor U17592 (N_17592,N_17401,N_17229);
xor U17593 (N_17593,N_17350,N_17443);
or U17594 (N_17594,N_17054,N_17483);
nand U17595 (N_17595,N_17481,N_17212);
xnor U17596 (N_17596,N_17147,N_17403);
nor U17597 (N_17597,N_17258,N_17377);
and U17598 (N_17598,N_17017,N_17170);
nor U17599 (N_17599,N_17203,N_17114);
nor U17600 (N_17600,N_17379,N_17004);
and U17601 (N_17601,N_17451,N_17375);
xnor U17602 (N_17602,N_17065,N_17038);
or U17603 (N_17603,N_17390,N_17426);
and U17604 (N_17604,N_17352,N_17006);
xnor U17605 (N_17605,N_17393,N_17127);
nand U17606 (N_17606,N_17196,N_17487);
nor U17607 (N_17607,N_17177,N_17118);
nand U17608 (N_17608,N_17130,N_17000);
nand U17609 (N_17609,N_17450,N_17184);
nor U17610 (N_17610,N_17452,N_17318);
and U17611 (N_17611,N_17302,N_17380);
nand U17612 (N_17612,N_17085,N_17355);
and U17613 (N_17613,N_17016,N_17068);
xor U17614 (N_17614,N_17090,N_17346);
xnor U17615 (N_17615,N_17018,N_17462);
or U17616 (N_17616,N_17183,N_17192);
nor U17617 (N_17617,N_17317,N_17033);
xor U17618 (N_17618,N_17230,N_17251);
nor U17619 (N_17619,N_17084,N_17050);
nor U17620 (N_17620,N_17210,N_17040);
nand U17621 (N_17621,N_17359,N_17199);
xor U17622 (N_17622,N_17301,N_17348);
nor U17623 (N_17623,N_17056,N_17070);
xnor U17624 (N_17624,N_17150,N_17268);
nor U17625 (N_17625,N_17216,N_17398);
xnor U17626 (N_17626,N_17099,N_17146);
nor U17627 (N_17627,N_17156,N_17285);
and U17628 (N_17628,N_17419,N_17312);
nor U17629 (N_17629,N_17421,N_17491);
and U17630 (N_17630,N_17071,N_17014);
and U17631 (N_17631,N_17386,N_17109);
nor U17632 (N_17632,N_17478,N_17304);
or U17633 (N_17633,N_17409,N_17002);
nor U17634 (N_17634,N_17492,N_17369);
xor U17635 (N_17635,N_17219,N_17209);
and U17636 (N_17636,N_17205,N_17427);
xor U17637 (N_17637,N_17339,N_17166);
nor U17638 (N_17638,N_17173,N_17122);
xnor U17639 (N_17639,N_17382,N_17308);
or U17640 (N_17640,N_17134,N_17223);
and U17641 (N_17641,N_17402,N_17460);
nand U17642 (N_17642,N_17336,N_17072);
nand U17643 (N_17643,N_17488,N_17024);
or U17644 (N_17644,N_17490,N_17148);
nand U17645 (N_17645,N_17220,N_17351);
nor U17646 (N_17646,N_17456,N_17168);
and U17647 (N_17647,N_17472,N_17388);
xor U17648 (N_17648,N_17370,N_17023);
and U17649 (N_17649,N_17331,N_17486);
nand U17650 (N_17650,N_17269,N_17292);
nor U17651 (N_17651,N_17180,N_17104);
or U17652 (N_17652,N_17262,N_17365);
and U17653 (N_17653,N_17179,N_17256);
or U17654 (N_17654,N_17128,N_17098);
or U17655 (N_17655,N_17045,N_17329);
nor U17656 (N_17656,N_17153,N_17307);
nor U17657 (N_17657,N_17238,N_17218);
xnor U17658 (N_17658,N_17353,N_17003);
nand U17659 (N_17659,N_17074,N_17105);
xor U17660 (N_17660,N_17455,N_17232);
nor U17661 (N_17661,N_17086,N_17198);
and U17662 (N_17662,N_17437,N_17007);
nor U17663 (N_17663,N_17294,N_17446);
nand U17664 (N_17664,N_17423,N_17154);
nand U17665 (N_17665,N_17465,N_17215);
xnor U17666 (N_17666,N_17049,N_17082);
xnor U17667 (N_17667,N_17103,N_17467);
or U17668 (N_17668,N_17343,N_17120);
xor U17669 (N_17669,N_17225,N_17121);
nand U17670 (N_17670,N_17366,N_17332);
xnor U17671 (N_17671,N_17342,N_17091);
xnor U17672 (N_17672,N_17126,N_17241);
xnor U17673 (N_17673,N_17287,N_17242);
and U17674 (N_17674,N_17228,N_17119);
xor U17675 (N_17675,N_17245,N_17226);
and U17676 (N_17676,N_17428,N_17176);
xnor U17677 (N_17677,N_17470,N_17163);
and U17678 (N_17678,N_17293,N_17244);
nand U17679 (N_17679,N_17195,N_17430);
or U17680 (N_17680,N_17466,N_17039);
nor U17681 (N_17681,N_17175,N_17284);
or U17682 (N_17682,N_17237,N_17001);
nand U17683 (N_17683,N_17345,N_17363);
nand U17684 (N_17684,N_17373,N_17440);
nor U17685 (N_17685,N_17132,N_17060);
xnor U17686 (N_17686,N_17371,N_17357);
nor U17687 (N_17687,N_17239,N_17108);
nor U17688 (N_17688,N_17197,N_17061);
xor U17689 (N_17689,N_17328,N_17325);
or U17690 (N_17690,N_17349,N_17497);
and U17691 (N_17691,N_17117,N_17075);
nand U17692 (N_17692,N_17188,N_17167);
nand U17693 (N_17693,N_17260,N_17012);
nand U17694 (N_17694,N_17438,N_17468);
and U17695 (N_17695,N_17270,N_17037);
xor U17696 (N_17696,N_17495,N_17087);
nand U17697 (N_17697,N_17025,N_17395);
xor U17698 (N_17698,N_17171,N_17316);
nor U17699 (N_17699,N_17073,N_17214);
nand U17700 (N_17700,N_17310,N_17337);
nand U17701 (N_17701,N_17052,N_17323);
xnor U17702 (N_17702,N_17137,N_17480);
and U17703 (N_17703,N_17493,N_17240);
or U17704 (N_17704,N_17474,N_17290);
nor U17705 (N_17705,N_17300,N_17059);
xnor U17706 (N_17706,N_17320,N_17447);
or U17707 (N_17707,N_17361,N_17356);
nor U17708 (N_17708,N_17187,N_17372);
and U17709 (N_17709,N_17288,N_17135);
or U17710 (N_17710,N_17432,N_17207);
nor U17711 (N_17711,N_17255,N_17093);
nand U17712 (N_17712,N_17283,N_17461);
nor U17713 (N_17713,N_17182,N_17169);
and U17714 (N_17714,N_17257,N_17165);
and U17715 (N_17715,N_17394,N_17111);
xnor U17716 (N_17716,N_17463,N_17064);
or U17717 (N_17717,N_17057,N_17469);
nor U17718 (N_17718,N_17208,N_17144);
or U17719 (N_17719,N_17172,N_17160);
nand U17720 (N_17720,N_17442,N_17236);
xor U17721 (N_17721,N_17224,N_17306);
nand U17722 (N_17722,N_17088,N_17282);
nand U17723 (N_17723,N_17249,N_17133);
nor U17724 (N_17724,N_17327,N_17027);
nor U17725 (N_17725,N_17378,N_17326);
nand U17726 (N_17726,N_17424,N_17191);
or U17727 (N_17727,N_17035,N_17020);
and U17728 (N_17728,N_17193,N_17374);
or U17729 (N_17729,N_17076,N_17030);
xor U17730 (N_17730,N_17407,N_17425);
xnor U17731 (N_17731,N_17142,N_17484);
nor U17732 (N_17732,N_17048,N_17482);
and U17733 (N_17733,N_17043,N_17032);
and U17734 (N_17734,N_17248,N_17221);
nand U17735 (N_17735,N_17115,N_17489);
or U17736 (N_17736,N_17140,N_17077);
and U17737 (N_17737,N_17036,N_17272);
nor U17738 (N_17738,N_17252,N_17106);
nor U17739 (N_17739,N_17107,N_17206);
or U17740 (N_17740,N_17174,N_17289);
or U17741 (N_17741,N_17454,N_17185);
nor U17742 (N_17742,N_17079,N_17022);
xor U17743 (N_17743,N_17391,N_17464);
nor U17744 (N_17744,N_17078,N_17340);
or U17745 (N_17745,N_17011,N_17278);
and U17746 (N_17746,N_17404,N_17319);
and U17747 (N_17747,N_17100,N_17281);
xor U17748 (N_17748,N_17247,N_17457);
and U17749 (N_17749,N_17138,N_17129);
nand U17750 (N_17750,N_17097,N_17156);
and U17751 (N_17751,N_17105,N_17073);
nand U17752 (N_17752,N_17162,N_17420);
nand U17753 (N_17753,N_17489,N_17352);
or U17754 (N_17754,N_17034,N_17226);
nand U17755 (N_17755,N_17297,N_17072);
and U17756 (N_17756,N_17250,N_17457);
nor U17757 (N_17757,N_17275,N_17364);
xnor U17758 (N_17758,N_17024,N_17419);
or U17759 (N_17759,N_17305,N_17300);
or U17760 (N_17760,N_17094,N_17293);
or U17761 (N_17761,N_17099,N_17203);
nand U17762 (N_17762,N_17378,N_17145);
nand U17763 (N_17763,N_17003,N_17376);
xor U17764 (N_17764,N_17243,N_17012);
and U17765 (N_17765,N_17486,N_17261);
and U17766 (N_17766,N_17139,N_17160);
or U17767 (N_17767,N_17258,N_17030);
nand U17768 (N_17768,N_17086,N_17096);
or U17769 (N_17769,N_17087,N_17028);
nor U17770 (N_17770,N_17166,N_17381);
xnor U17771 (N_17771,N_17366,N_17405);
and U17772 (N_17772,N_17414,N_17475);
nor U17773 (N_17773,N_17072,N_17130);
nand U17774 (N_17774,N_17246,N_17436);
or U17775 (N_17775,N_17104,N_17354);
nand U17776 (N_17776,N_17277,N_17109);
nor U17777 (N_17777,N_17485,N_17346);
nor U17778 (N_17778,N_17414,N_17298);
xor U17779 (N_17779,N_17207,N_17349);
or U17780 (N_17780,N_17126,N_17203);
and U17781 (N_17781,N_17419,N_17487);
or U17782 (N_17782,N_17278,N_17439);
and U17783 (N_17783,N_17243,N_17051);
nor U17784 (N_17784,N_17340,N_17054);
and U17785 (N_17785,N_17073,N_17144);
xor U17786 (N_17786,N_17375,N_17278);
xor U17787 (N_17787,N_17203,N_17219);
nor U17788 (N_17788,N_17404,N_17048);
or U17789 (N_17789,N_17083,N_17118);
or U17790 (N_17790,N_17310,N_17095);
xor U17791 (N_17791,N_17174,N_17163);
or U17792 (N_17792,N_17341,N_17010);
nand U17793 (N_17793,N_17416,N_17159);
and U17794 (N_17794,N_17140,N_17222);
or U17795 (N_17795,N_17153,N_17399);
nand U17796 (N_17796,N_17092,N_17098);
and U17797 (N_17797,N_17279,N_17344);
and U17798 (N_17798,N_17464,N_17012);
xnor U17799 (N_17799,N_17185,N_17005);
xnor U17800 (N_17800,N_17323,N_17237);
and U17801 (N_17801,N_17110,N_17190);
xor U17802 (N_17802,N_17014,N_17389);
nand U17803 (N_17803,N_17096,N_17304);
and U17804 (N_17804,N_17294,N_17383);
nor U17805 (N_17805,N_17265,N_17172);
or U17806 (N_17806,N_17140,N_17152);
nand U17807 (N_17807,N_17465,N_17027);
or U17808 (N_17808,N_17177,N_17325);
or U17809 (N_17809,N_17271,N_17487);
xor U17810 (N_17810,N_17012,N_17200);
and U17811 (N_17811,N_17328,N_17165);
nand U17812 (N_17812,N_17186,N_17232);
and U17813 (N_17813,N_17437,N_17119);
nand U17814 (N_17814,N_17393,N_17006);
nor U17815 (N_17815,N_17290,N_17356);
and U17816 (N_17816,N_17069,N_17066);
xnor U17817 (N_17817,N_17472,N_17342);
and U17818 (N_17818,N_17139,N_17389);
or U17819 (N_17819,N_17418,N_17359);
or U17820 (N_17820,N_17381,N_17499);
nand U17821 (N_17821,N_17428,N_17098);
nand U17822 (N_17822,N_17125,N_17497);
nor U17823 (N_17823,N_17312,N_17334);
or U17824 (N_17824,N_17431,N_17004);
and U17825 (N_17825,N_17337,N_17184);
or U17826 (N_17826,N_17067,N_17173);
nor U17827 (N_17827,N_17491,N_17078);
nand U17828 (N_17828,N_17372,N_17386);
or U17829 (N_17829,N_17250,N_17206);
nor U17830 (N_17830,N_17361,N_17424);
nor U17831 (N_17831,N_17088,N_17075);
and U17832 (N_17832,N_17189,N_17220);
and U17833 (N_17833,N_17248,N_17117);
nor U17834 (N_17834,N_17379,N_17305);
xor U17835 (N_17835,N_17070,N_17160);
or U17836 (N_17836,N_17370,N_17405);
xnor U17837 (N_17837,N_17030,N_17355);
or U17838 (N_17838,N_17352,N_17179);
and U17839 (N_17839,N_17436,N_17032);
and U17840 (N_17840,N_17430,N_17323);
nor U17841 (N_17841,N_17405,N_17441);
or U17842 (N_17842,N_17022,N_17036);
xor U17843 (N_17843,N_17017,N_17332);
nor U17844 (N_17844,N_17200,N_17146);
and U17845 (N_17845,N_17482,N_17030);
nand U17846 (N_17846,N_17047,N_17157);
xnor U17847 (N_17847,N_17237,N_17386);
nor U17848 (N_17848,N_17457,N_17185);
nor U17849 (N_17849,N_17130,N_17009);
xor U17850 (N_17850,N_17235,N_17325);
xnor U17851 (N_17851,N_17050,N_17308);
nor U17852 (N_17852,N_17062,N_17239);
or U17853 (N_17853,N_17009,N_17486);
nor U17854 (N_17854,N_17145,N_17484);
and U17855 (N_17855,N_17248,N_17341);
and U17856 (N_17856,N_17317,N_17121);
nand U17857 (N_17857,N_17029,N_17377);
xor U17858 (N_17858,N_17269,N_17287);
and U17859 (N_17859,N_17010,N_17226);
or U17860 (N_17860,N_17162,N_17433);
nand U17861 (N_17861,N_17190,N_17396);
or U17862 (N_17862,N_17280,N_17411);
or U17863 (N_17863,N_17420,N_17322);
xnor U17864 (N_17864,N_17129,N_17070);
and U17865 (N_17865,N_17299,N_17220);
nand U17866 (N_17866,N_17193,N_17481);
nor U17867 (N_17867,N_17360,N_17190);
or U17868 (N_17868,N_17055,N_17283);
nor U17869 (N_17869,N_17159,N_17040);
nand U17870 (N_17870,N_17464,N_17335);
xor U17871 (N_17871,N_17050,N_17466);
and U17872 (N_17872,N_17371,N_17310);
xor U17873 (N_17873,N_17211,N_17387);
and U17874 (N_17874,N_17163,N_17319);
xor U17875 (N_17875,N_17279,N_17433);
xor U17876 (N_17876,N_17311,N_17384);
nor U17877 (N_17877,N_17486,N_17264);
and U17878 (N_17878,N_17392,N_17091);
xor U17879 (N_17879,N_17277,N_17003);
and U17880 (N_17880,N_17320,N_17089);
xor U17881 (N_17881,N_17078,N_17069);
and U17882 (N_17882,N_17216,N_17075);
xor U17883 (N_17883,N_17390,N_17154);
and U17884 (N_17884,N_17434,N_17037);
or U17885 (N_17885,N_17402,N_17203);
xnor U17886 (N_17886,N_17293,N_17153);
nand U17887 (N_17887,N_17366,N_17444);
nor U17888 (N_17888,N_17167,N_17202);
and U17889 (N_17889,N_17324,N_17013);
or U17890 (N_17890,N_17200,N_17459);
or U17891 (N_17891,N_17232,N_17211);
and U17892 (N_17892,N_17485,N_17392);
or U17893 (N_17893,N_17338,N_17450);
nor U17894 (N_17894,N_17461,N_17260);
nand U17895 (N_17895,N_17384,N_17120);
or U17896 (N_17896,N_17412,N_17116);
nor U17897 (N_17897,N_17440,N_17028);
xor U17898 (N_17898,N_17492,N_17046);
nor U17899 (N_17899,N_17023,N_17108);
nor U17900 (N_17900,N_17228,N_17340);
and U17901 (N_17901,N_17340,N_17208);
and U17902 (N_17902,N_17153,N_17051);
or U17903 (N_17903,N_17269,N_17178);
or U17904 (N_17904,N_17064,N_17128);
nor U17905 (N_17905,N_17297,N_17001);
nor U17906 (N_17906,N_17454,N_17334);
or U17907 (N_17907,N_17030,N_17100);
or U17908 (N_17908,N_17307,N_17102);
or U17909 (N_17909,N_17052,N_17397);
nand U17910 (N_17910,N_17145,N_17281);
or U17911 (N_17911,N_17177,N_17025);
nor U17912 (N_17912,N_17159,N_17122);
xnor U17913 (N_17913,N_17445,N_17255);
or U17914 (N_17914,N_17027,N_17450);
nand U17915 (N_17915,N_17133,N_17141);
nor U17916 (N_17916,N_17177,N_17426);
xnor U17917 (N_17917,N_17351,N_17071);
nor U17918 (N_17918,N_17480,N_17218);
and U17919 (N_17919,N_17140,N_17326);
and U17920 (N_17920,N_17267,N_17018);
nand U17921 (N_17921,N_17371,N_17466);
nand U17922 (N_17922,N_17211,N_17477);
xnor U17923 (N_17923,N_17052,N_17148);
nand U17924 (N_17924,N_17272,N_17013);
nand U17925 (N_17925,N_17104,N_17078);
and U17926 (N_17926,N_17272,N_17185);
nand U17927 (N_17927,N_17125,N_17493);
or U17928 (N_17928,N_17231,N_17353);
or U17929 (N_17929,N_17040,N_17371);
and U17930 (N_17930,N_17197,N_17284);
or U17931 (N_17931,N_17087,N_17146);
xor U17932 (N_17932,N_17362,N_17339);
nand U17933 (N_17933,N_17209,N_17437);
nand U17934 (N_17934,N_17009,N_17421);
or U17935 (N_17935,N_17023,N_17130);
and U17936 (N_17936,N_17408,N_17221);
nand U17937 (N_17937,N_17486,N_17110);
nand U17938 (N_17938,N_17405,N_17384);
and U17939 (N_17939,N_17318,N_17487);
and U17940 (N_17940,N_17464,N_17153);
nor U17941 (N_17941,N_17332,N_17186);
nor U17942 (N_17942,N_17283,N_17144);
and U17943 (N_17943,N_17456,N_17136);
or U17944 (N_17944,N_17406,N_17211);
xor U17945 (N_17945,N_17451,N_17193);
or U17946 (N_17946,N_17261,N_17024);
xor U17947 (N_17947,N_17144,N_17405);
or U17948 (N_17948,N_17178,N_17140);
xnor U17949 (N_17949,N_17445,N_17240);
xor U17950 (N_17950,N_17041,N_17407);
xnor U17951 (N_17951,N_17248,N_17099);
nor U17952 (N_17952,N_17280,N_17218);
nand U17953 (N_17953,N_17175,N_17247);
xnor U17954 (N_17954,N_17343,N_17280);
xor U17955 (N_17955,N_17277,N_17035);
and U17956 (N_17956,N_17361,N_17078);
and U17957 (N_17957,N_17322,N_17369);
or U17958 (N_17958,N_17081,N_17328);
xnor U17959 (N_17959,N_17450,N_17371);
nand U17960 (N_17960,N_17472,N_17481);
nor U17961 (N_17961,N_17024,N_17209);
nor U17962 (N_17962,N_17167,N_17233);
xor U17963 (N_17963,N_17401,N_17332);
nand U17964 (N_17964,N_17442,N_17459);
nor U17965 (N_17965,N_17004,N_17182);
or U17966 (N_17966,N_17368,N_17488);
xor U17967 (N_17967,N_17219,N_17117);
and U17968 (N_17968,N_17227,N_17114);
or U17969 (N_17969,N_17170,N_17385);
or U17970 (N_17970,N_17473,N_17042);
nor U17971 (N_17971,N_17215,N_17180);
nand U17972 (N_17972,N_17281,N_17248);
nor U17973 (N_17973,N_17152,N_17364);
nand U17974 (N_17974,N_17037,N_17389);
nor U17975 (N_17975,N_17494,N_17128);
and U17976 (N_17976,N_17127,N_17271);
nand U17977 (N_17977,N_17442,N_17283);
or U17978 (N_17978,N_17195,N_17472);
or U17979 (N_17979,N_17351,N_17013);
nand U17980 (N_17980,N_17005,N_17311);
xor U17981 (N_17981,N_17086,N_17296);
nand U17982 (N_17982,N_17064,N_17038);
xnor U17983 (N_17983,N_17105,N_17122);
xor U17984 (N_17984,N_17355,N_17262);
nand U17985 (N_17985,N_17028,N_17117);
and U17986 (N_17986,N_17312,N_17412);
nand U17987 (N_17987,N_17036,N_17194);
and U17988 (N_17988,N_17130,N_17192);
xor U17989 (N_17989,N_17266,N_17353);
or U17990 (N_17990,N_17058,N_17315);
or U17991 (N_17991,N_17350,N_17253);
nand U17992 (N_17992,N_17124,N_17377);
or U17993 (N_17993,N_17454,N_17368);
or U17994 (N_17994,N_17009,N_17212);
xor U17995 (N_17995,N_17289,N_17240);
xnor U17996 (N_17996,N_17125,N_17326);
nor U17997 (N_17997,N_17180,N_17086);
nand U17998 (N_17998,N_17404,N_17367);
and U17999 (N_17999,N_17453,N_17166);
nor U18000 (N_18000,N_17528,N_17561);
nand U18001 (N_18001,N_17869,N_17517);
or U18002 (N_18002,N_17660,N_17673);
and U18003 (N_18003,N_17875,N_17549);
or U18004 (N_18004,N_17831,N_17680);
nand U18005 (N_18005,N_17574,N_17953);
and U18006 (N_18006,N_17519,N_17692);
and U18007 (N_18007,N_17954,N_17551);
xnor U18008 (N_18008,N_17633,N_17868);
nand U18009 (N_18009,N_17809,N_17971);
nand U18010 (N_18010,N_17650,N_17732);
xor U18011 (N_18011,N_17957,N_17911);
nor U18012 (N_18012,N_17717,N_17945);
nand U18013 (N_18013,N_17758,N_17990);
or U18014 (N_18014,N_17573,N_17559);
xnor U18015 (N_18015,N_17966,N_17544);
and U18016 (N_18016,N_17641,N_17931);
xnor U18017 (N_18017,N_17932,N_17593);
nor U18018 (N_18018,N_17623,N_17645);
or U18019 (N_18019,N_17882,N_17504);
nor U18020 (N_18020,N_17605,N_17858);
and U18021 (N_18021,N_17893,N_17782);
nand U18022 (N_18022,N_17901,N_17572);
or U18023 (N_18023,N_17999,N_17897);
and U18024 (N_18024,N_17711,N_17859);
nand U18025 (N_18025,N_17698,N_17838);
and U18026 (N_18026,N_17766,N_17750);
nand U18027 (N_18027,N_17860,N_17806);
nor U18028 (N_18028,N_17777,N_17994);
nor U18029 (N_18029,N_17805,N_17686);
nor U18030 (N_18030,N_17647,N_17915);
nand U18031 (N_18031,N_17667,N_17939);
nand U18032 (N_18032,N_17885,N_17850);
nor U18033 (N_18033,N_17761,N_17719);
nand U18034 (N_18034,N_17889,N_17700);
or U18035 (N_18035,N_17703,N_17886);
or U18036 (N_18036,N_17898,N_17563);
nor U18037 (N_18037,N_17514,N_17756);
and U18038 (N_18038,N_17841,N_17943);
and U18039 (N_18039,N_17852,N_17890);
nand U18040 (N_18040,N_17793,N_17724);
or U18041 (N_18041,N_17798,N_17854);
nor U18042 (N_18042,N_17595,N_17699);
nand U18043 (N_18043,N_17951,N_17861);
nand U18044 (N_18044,N_17853,N_17884);
nand U18045 (N_18045,N_17878,N_17855);
nor U18046 (N_18046,N_17786,N_17701);
xor U18047 (N_18047,N_17708,N_17613);
nor U18048 (N_18048,N_17640,N_17787);
nand U18049 (N_18049,N_17618,N_17586);
nand U18050 (N_18050,N_17876,N_17585);
xor U18051 (N_18051,N_17873,N_17946);
and U18052 (N_18052,N_17888,N_17552);
and U18053 (N_18053,N_17783,N_17626);
and U18054 (N_18054,N_17790,N_17808);
and U18055 (N_18055,N_17933,N_17553);
nor U18056 (N_18056,N_17677,N_17601);
or U18057 (N_18057,N_17863,N_17986);
nand U18058 (N_18058,N_17908,N_17634);
nand U18059 (N_18059,N_17762,N_17527);
nor U18060 (N_18060,N_17813,N_17710);
xnor U18061 (N_18061,N_17952,N_17803);
nor U18062 (N_18062,N_17820,N_17907);
nand U18063 (N_18063,N_17739,N_17529);
or U18064 (N_18064,N_17606,N_17578);
and U18065 (N_18065,N_17515,N_17668);
and U18066 (N_18066,N_17991,N_17695);
and U18067 (N_18067,N_17864,N_17520);
nor U18068 (N_18068,N_17735,N_17902);
xnor U18069 (N_18069,N_17771,N_17877);
and U18070 (N_18070,N_17591,N_17845);
and U18071 (N_18071,N_17510,N_17538);
nand U18072 (N_18072,N_17649,N_17665);
or U18073 (N_18073,N_17922,N_17925);
and U18074 (N_18074,N_17584,N_17643);
nand U18075 (N_18075,N_17899,N_17644);
nor U18076 (N_18076,N_17534,N_17799);
nand U18077 (N_18077,N_17693,N_17705);
nor U18078 (N_18078,N_17507,N_17823);
nand U18079 (N_18079,N_17690,N_17804);
or U18080 (N_18080,N_17955,N_17681);
or U18081 (N_18081,N_17731,N_17826);
xnor U18082 (N_18082,N_17988,N_17958);
or U18083 (N_18083,N_17663,N_17862);
or U18084 (N_18084,N_17879,N_17604);
xor U18085 (N_18085,N_17718,N_17594);
xnor U18086 (N_18086,N_17906,N_17576);
and U18087 (N_18087,N_17967,N_17734);
nand U18088 (N_18088,N_17714,N_17631);
nor U18089 (N_18089,N_17842,N_17749);
and U18090 (N_18090,N_17661,N_17599);
or U18091 (N_18091,N_17941,N_17785);
nand U18092 (N_18092,N_17913,N_17580);
and U18093 (N_18093,N_17506,N_17961);
nor U18094 (N_18094,N_17742,N_17814);
nor U18095 (N_18095,N_17993,N_17942);
and U18096 (N_18096,N_17920,N_17977);
nor U18097 (N_18097,N_17546,N_17726);
nor U18098 (N_18098,N_17759,N_17555);
xor U18099 (N_18099,N_17980,N_17696);
and U18100 (N_18100,N_17533,N_17691);
xor U18101 (N_18101,N_17827,N_17929);
nor U18102 (N_18102,N_17646,N_17664);
xor U18103 (N_18103,N_17652,N_17697);
nor U18104 (N_18104,N_17684,N_17629);
or U18105 (N_18105,N_17795,N_17910);
nor U18106 (N_18106,N_17598,N_17775);
or U18107 (N_18107,N_17588,N_17679);
or U18108 (N_18108,N_17763,N_17753);
or U18109 (N_18109,N_17648,N_17694);
and U18110 (N_18110,N_17887,N_17505);
and U18111 (N_18111,N_17521,N_17938);
and U18112 (N_18112,N_17728,N_17716);
and U18113 (N_18113,N_17924,N_17557);
nand U18114 (N_18114,N_17927,N_17655);
nand U18115 (N_18115,N_17748,N_17675);
nand U18116 (N_18116,N_17669,N_17702);
xnor U18117 (N_18117,N_17627,N_17767);
and U18118 (N_18118,N_17562,N_17656);
or U18119 (N_18119,N_17976,N_17755);
nor U18120 (N_18120,N_17968,N_17712);
and U18121 (N_18121,N_17810,N_17956);
or U18122 (N_18122,N_17676,N_17670);
or U18123 (N_18123,N_17821,N_17733);
xor U18124 (N_18124,N_17754,N_17919);
nor U18125 (N_18125,N_17848,N_17543);
nor U18126 (N_18126,N_17581,N_17843);
and U18127 (N_18127,N_17948,N_17794);
nand U18128 (N_18128,N_17801,N_17531);
and U18129 (N_18129,N_17721,N_17583);
nor U18130 (N_18130,N_17896,N_17727);
xor U18131 (N_18131,N_17545,N_17713);
and U18132 (N_18132,N_17959,N_17964);
xor U18133 (N_18133,N_17788,N_17904);
nor U18134 (N_18134,N_17621,N_17635);
nand U18135 (N_18135,N_17638,N_17797);
and U18136 (N_18136,N_17985,N_17789);
nand U18137 (N_18137,N_17628,N_17530);
xor U18138 (N_18138,N_17921,N_17846);
nor U18139 (N_18139,N_17653,N_17725);
and U18140 (N_18140,N_17688,N_17930);
nand U18141 (N_18141,N_17720,N_17865);
xor U18142 (N_18142,N_17597,N_17508);
nand U18143 (N_18143,N_17824,N_17916);
and U18144 (N_18144,N_17666,N_17589);
nor U18145 (N_18145,N_17949,N_17779);
nor U18146 (N_18146,N_17834,N_17587);
and U18147 (N_18147,N_17730,N_17619);
nor U18148 (N_18148,N_17822,N_17503);
or U18149 (N_18149,N_17825,N_17833);
and U18150 (N_18150,N_17659,N_17770);
nor U18151 (N_18151,N_17513,N_17740);
or U18152 (N_18152,N_17772,N_17526);
xnor U18153 (N_18153,N_17987,N_17685);
nor U18154 (N_18154,N_17654,N_17737);
or U18155 (N_18155,N_17819,N_17516);
and U18156 (N_18156,N_17556,N_17774);
xnor U18157 (N_18157,N_17895,N_17607);
and U18158 (N_18158,N_17998,N_17539);
nor U18159 (N_18159,N_17917,N_17632);
nand U18160 (N_18160,N_17566,N_17729);
xor U18161 (N_18161,N_17651,N_17620);
or U18162 (N_18162,N_17983,N_17751);
nor U18163 (N_18163,N_17624,N_17947);
nor U18164 (N_18164,N_17704,N_17818);
or U18165 (N_18165,N_17856,N_17745);
or U18166 (N_18166,N_17642,N_17744);
xor U18167 (N_18167,N_17963,N_17829);
or U18168 (N_18168,N_17535,N_17903);
xor U18169 (N_18169,N_17760,N_17500);
and U18170 (N_18170,N_17894,N_17537);
nand U18171 (N_18171,N_17611,N_17905);
and U18172 (N_18172,N_17600,N_17791);
and U18173 (N_18173,N_17547,N_17837);
or U18174 (N_18174,N_17674,N_17768);
nand U18175 (N_18175,N_17839,N_17844);
nand U18176 (N_18176,N_17891,N_17511);
or U18177 (N_18177,N_17682,N_17867);
nand U18178 (N_18178,N_17541,N_17757);
or U18179 (N_18179,N_17602,N_17579);
xor U18180 (N_18180,N_17773,N_17914);
nor U18181 (N_18181,N_17715,N_17603);
xor U18182 (N_18182,N_17836,N_17792);
or U18183 (N_18183,N_17592,N_17548);
nand U18184 (N_18184,N_17969,N_17912);
and U18185 (N_18185,N_17923,N_17509);
xor U18186 (N_18186,N_17973,N_17741);
nand U18187 (N_18187,N_17997,N_17512);
nor U18188 (N_18188,N_17784,N_17662);
or U18189 (N_18189,N_17706,N_17870);
and U18190 (N_18190,N_17525,N_17937);
nand U18191 (N_18191,N_17612,N_17637);
and U18192 (N_18192,N_17802,N_17900);
nor U18193 (N_18193,N_17816,N_17746);
nor U18194 (N_18194,N_17769,N_17689);
or U18195 (N_18195,N_17996,N_17830);
and U18196 (N_18196,N_17974,N_17502);
or U18197 (N_18197,N_17934,N_17738);
xor U18198 (N_18198,N_17582,N_17874);
xor U18199 (N_18199,N_17960,N_17892);
nor U18200 (N_18200,N_17965,N_17950);
xnor U18201 (N_18201,N_17847,N_17657);
nor U18202 (N_18202,N_17610,N_17558);
and U18203 (N_18203,N_17722,N_17807);
and U18204 (N_18204,N_17536,N_17880);
and U18205 (N_18205,N_17811,N_17992);
or U18206 (N_18206,N_17560,N_17778);
nor U18207 (N_18207,N_17776,N_17752);
nor U18208 (N_18208,N_17982,N_17926);
or U18209 (N_18209,N_17617,N_17940);
xor U18210 (N_18210,N_17928,N_17564);
xor U18211 (N_18211,N_17989,N_17723);
nor U18212 (N_18212,N_17866,N_17909);
xor U18213 (N_18213,N_17540,N_17849);
nor U18214 (N_18214,N_17709,N_17981);
nor U18215 (N_18215,N_17577,N_17532);
or U18216 (N_18216,N_17569,N_17857);
or U18217 (N_18217,N_17872,N_17796);
nor U18218 (N_18218,N_17736,N_17615);
or U18219 (N_18219,N_17972,N_17678);
or U18220 (N_18220,N_17565,N_17780);
nor U18221 (N_18221,N_17743,N_17764);
xor U18222 (N_18222,N_17658,N_17571);
nor U18223 (N_18223,N_17671,N_17815);
and U18224 (N_18224,N_17962,N_17522);
nand U18225 (N_18225,N_17812,N_17781);
or U18226 (N_18226,N_17616,N_17883);
nor U18227 (N_18227,N_17614,N_17567);
xor U18228 (N_18228,N_17672,N_17979);
or U18229 (N_18229,N_17609,N_17630);
nor U18230 (N_18230,N_17835,N_17984);
nor U18231 (N_18231,N_17608,N_17518);
xnor U18232 (N_18232,N_17944,N_17881);
nor U18233 (N_18233,N_17554,N_17622);
or U18234 (N_18234,N_17550,N_17707);
or U18235 (N_18235,N_17828,N_17590);
or U18236 (N_18236,N_17918,N_17568);
nand U18237 (N_18237,N_17800,N_17978);
nor U18238 (N_18238,N_17625,N_17596);
nand U18239 (N_18239,N_17524,N_17501);
and U18240 (N_18240,N_17636,N_17683);
and U18241 (N_18241,N_17995,N_17975);
and U18242 (N_18242,N_17935,N_17570);
and U18243 (N_18243,N_17936,N_17832);
and U18244 (N_18244,N_17765,N_17575);
nor U18245 (N_18245,N_17542,N_17687);
nor U18246 (N_18246,N_17840,N_17747);
nor U18247 (N_18247,N_17639,N_17523);
or U18248 (N_18248,N_17817,N_17970);
xor U18249 (N_18249,N_17851,N_17871);
and U18250 (N_18250,N_17721,N_17967);
xnor U18251 (N_18251,N_17625,N_17622);
nand U18252 (N_18252,N_17677,N_17878);
and U18253 (N_18253,N_17859,N_17744);
and U18254 (N_18254,N_17708,N_17667);
nand U18255 (N_18255,N_17630,N_17533);
xor U18256 (N_18256,N_17835,N_17765);
and U18257 (N_18257,N_17858,N_17720);
or U18258 (N_18258,N_17765,N_17980);
xnor U18259 (N_18259,N_17882,N_17625);
xnor U18260 (N_18260,N_17817,N_17537);
and U18261 (N_18261,N_17818,N_17524);
xnor U18262 (N_18262,N_17658,N_17932);
and U18263 (N_18263,N_17986,N_17902);
nor U18264 (N_18264,N_17746,N_17861);
or U18265 (N_18265,N_17998,N_17582);
xnor U18266 (N_18266,N_17824,N_17604);
nor U18267 (N_18267,N_17886,N_17789);
nand U18268 (N_18268,N_17759,N_17723);
xor U18269 (N_18269,N_17851,N_17670);
nor U18270 (N_18270,N_17982,N_17680);
xor U18271 (N_18271,N_17670,N_17797);
nor U18272 (N_18272,N_17735,N_17971);
nor U18273 (N_18273,N_17837,N_17588);
nor U18274 (N_18274,N_17844,N_17842);
nor U18275 (N_18275,N_17837,N_17782);
or U18276 (N_18276,N_17722,N_17867);
and U18277 (N_18277,N_17981,N_17572);
and U18278 (N_18278,N_17674,N_17972);
nand U18279 (N_18279,N_17802,N_17588);
nor U18280 (N_18280,N_17558,N_17950);
nand U18281 (N_18281,N_17867,N_17580);
nand U18282 (N_18282,N_17520,N_17813);
xnor U18283 (N_18283,N_17543,N_17540);
nand U18284 (N_18284,N_17543,N_17783);
xor U18285 (N_18285,N_17939,N_17594);
xor U18286 (N_18286,N_17875,N_17784);
nand U18287 (N_18287,N_17893,N_17753);
nand U18288 (N_18288,N_17792,N_17817);
nor U18289 (N_18289,N_17638,N_17959);
nand U18290 (N_18290,N_17953,N_17533);
nor U18291 (N_18291,N_17826,N_17888);
nand U18292 (N_18292,N_17557,N_17746);
nor U18293 (N_18293,N_17863,N_17756);
nand U18294 (N_18294,N_17898,N_17875);
or U18295 (N_18295,N_17542,N_17822);
nand U18296 (N_18296,N_17829,N_17971);
or U18297 (N_18297,N_17785,N_17780);
nand U18298 (N_18298,N_17572,N_17605);
and U18299 (N_18299,N_17825,N_17644);
nand U18300 (N_18300,N_17610,N_17675);
nor U18301 (N_18301,N_17900,N_17664);
nor U18302 (N_18302,N_17663,N_17547);
xor U18303 (N_18303,N_17880,N_17518);
nand U18304 (N_18304,N_17785,N_17836);
or U18305 (N_18305,N_17788,N_17666);
and U18306 (N_18306,N_17638,N_17992);
or U18307 (N_18307,N_17889,N_17583);
xor U18308 (N_18308,N_17975,N_17666);
xor U18309 (N_18309,N_17951,N_17554);
nand U18310 (N_18310,N_17721,N_17504);
nand U18311 (N_18311,N_17583,N_17559);
and U18312 (N_18312,N_17768,N_17679);
xnor U18313 (N_18313,N_17618,N_17769);
xor U18314 (N_18314,N_17973,N_17754);
or U18315 (N_18315,N_17648,N_17704);
nand U18316 (N_18316,N_17599,N_17819);
and U18317 (N_18317,N_17626,N_17729);
nor U18318 (N_18318,N_17610,N_17767);
xnor U18319 (N_18319,N_17861,N_17539);
nand U18320 (N_18320,N_17999,N_17903);
nor U18321 (N_18321,N_17805,N_17628);
and U18322 (N_18322,N_17617,N_17886);
and U18323 (N_18323,N_17520,N_17956);
nand U18324 (N_18324,N_17605,N_17676);
nand U18325 (N_18325,N_17892,N_17587);
or U18326 (N_18326,N_17718,N_17680);
and U18327 (N_18327,N_17643,N_17830);
nand U18328 (N_18328,N_17674,N_17555);
nand U18329 (N_18329,N_17660,N_17824);
xor U18330 (N_18330,N_17812,N_17746);
xor U18331 (N_18331,N_17985,N_17638);
xor U18332 (N_18332,N_17683,N_17629);
or U18333 (N_18333,N_17662,N_17613);
or U18334 (N_18334,N_17555,N_17755);
nand U18335 (N_18335,N_17975,N_17600);
or U18336 (N_18336,N_17546,N_17974);
nor U18337 (N_18337,N_17645,N_17860);
nor U18338 (N_18338,N_17833,N_17780);
xor U18339 (N_18339,N_17804,N_17509);
and U18340 (N_18340,N_17892,N_17963);
or U18341 (N_18341,N_17741,N_17971);
xnor U18342 (N_18342,N_17840,N_17922);
or U18343 (N_18343,N_17586,N_17834);
and U18344 (N_18344,N_17537,N_17851);
nand U18345 (N_18345,N_17838,N_17881);
nor U18346 (N_18346,N_17555,N_17628);
or U18347 (N_18347,N_17950,N_17852);
xnor U18348 (N_18348,N_17878,N_17900);
and U18349 (N_18349,N_17808,N_17509);
xor U18350 (N_18350,N_17677,N_17927);
and U18351 (N_18351,N_17815,N_17883);
nand U18352 (N_18352,N_17753,N_17620);
and U18353 (N_18353,N_17601,N_17814);
xnor U18354 (N_18354,N_17861,N_17554);
nor U18355 (N_18355,N_17858,N_17846);
nand U18356 (N_18356,N_17992,N_17823);
and U18357 (N_18357,N_17962,N_17881);
or U18358 (N_18358,N_17633,N_17938);
nand U18359 (N_18359,N_17872,N_17850);
or U18360 (N_18360,N_17604,N_17955);
xnor U18361 (N_18361,N_17742,N_17776);
nor U18362 (N_18362,N_17800,N_17865);
xor U18363 (N_18363,N_17829,N_17912);
or U18364 (N_18364,N_17862,N_17702);
nand U18365 (N_18365,N_17861,N_17806);
nand U18366 (N_18366,N_17781,N_17661);
and U18367 (N_18367,N_17594,N_17613);
nor U18368 (N_18368,N_17868,N_17862);
and U18369 (N_18369,N_17897,N_17705);
nand U18370 (N_18370,N_17998,N_17791);
or U18371 (N_18371,N_17680,N_17535);
nand U18372 (N_18372,N_17559,N_17504);
nand U18373 (N_18373,N_17806,N_17776);
nand U18374 (N_18374,N_17588,N_17796);
nor U18375 (N_18375,N_17756,N_17673);
nand U18376 (N_18376,N_17913,N_17535);
xnor U18377 (N_18377,N_17855,N_17747);
xor U18378 (N_18378,N_17840,N_17948);
nand U18379 (N_18379,N_17648,N_17976);
or U18380 (N_18380,N_17982,N_17745);
nor U18381 (N_18381,N_17598,N_17961);
and U18382 (N_18382,N_17927,N_17836);
or U18383 (N_18383,N_17531,N_17556);
xor U18384 (N_18384,N_17686,N_17812);
nor U18385 (N_18385,N_17723,N_17803);
and U18386 (N_18386,N_17802,N_17513);
nor U18387 (N_18387,N_17584,N_17796);
or U18388 (N_18388,N_17533,N_17728);
nand U18389 (N_18389,N_17906,N_17907);
nor U18390 (N_18390,N_17827,N_17999);
and U18391 (N_18391,N_17575,N_17993);
or U18392 (N_18392,N_17801,N_17857);
nand U18393 (N_18393,N_17731,N_17520);
nor U18394 (N_18394,N_17525,N_17661);
and U18395 (N_18395,N_17522,N_17743);
or U18396 (N_18396,N_17526,N_17930);
and U18397 (N_18397,N_17817,N_17780);
nand U18398 (N_18398,N_17574,N_17603);
xor U18399 (N_18399,N_17810,N_17722);
and U18400 (N_18400,N_17816,N_17675);
nand U18401 (N_18401,N_17643,N_17884);
nand U18402 (N_18402,N_17906,N_17710);
xor U18403 (N_18403,N_17801,N_17750);
and U18404 (N_18404,N_17871,N_17948);
nor U18405 (N_18405,N_17843,N_17935);
or U18406 (N_18406,N_17931,N_17644);
nand U18407 (N_18407,N_17742,N_17723);
nand U18408 (N_18408,N_17741,N_17989);
and U18409 (N_18409,N_17975,N_17832);
nor U18410 (N_18410,N_17641,N_17610);
xnor U18411 (N_18411,N_17925,N_17536);
and U18412 (N_18412,N_17787,N_17921);
xnor U18413 (N_18413,N_17575,N_17866);
nand U18414 (N_18414,N_17756,N_17901);
xnor U18415 (N_18415,N_17679,N_17675);
and U18416 (N_18416,N_17727,N_17789);
nor U18417 (N_18417,N_17679,N_17805);
and U18418 (N_18418,N_17536,N_17990);
nor U18419 (N_18419,N_17763,N_17681);
nand U18420 (N_18420,N_17718,N_17587);
nor U18421 (N_18421,N_17816,N_17804);
or U18422 (N_18422,N_17729,N_17680);
nand U18423 (N_18423,N_17621,N_17535);
xor U18424 (N_18424,N_17922,N_17792);
xnor U18425 (N_18425,N_17667,N_17504);
and U18426 (N_18426,N_17868,N_17833);
and U18427 (N_18427,N_17636,N_17850);
nand U18428 (N_18428,N_17933,N_17694);
or U18429 (N_18429,N_17751,N_17628);
nor U18430 (N_18430,N_17718,N_17701);
xor U18431 (N_18431,N_17509,N_17915);
nand U18432 (N_18432,N_17579,N_17574);
or U18433 (N_18433,N_17902,N_17961);
xnor U18434 (N_18434,N_17568,N_17534);
nand U18435 (N_18435,N_17623,N_17999);
and U18436 (N_18436,N_17954,N_17505);
nor U18437 (N_18437,N_17992,N_17850);
nor U18438 (N_18438,N_17914,N_17762);
nor U18439 (N_18439,N_17509,N_17943);
nor U18440 (N_18440,N_17813,N_17860);
or U18441 (N_18441,N_17919,N_17976);
and U18442 (N_18442,N_17672,N_17704);
and U18443 (N_18443,N_17997,N_17921);
and U18444 (N_18444,N_17870,N_17885);
or U18445 (N_18445,N_17557,N_17768);
nor U18446 (N_18446,N_17589,N_17967);
xor U18447 (N_18447,N_17781,N_17864);
xor U18448 (N_18448,N_17579,N_17646);
or U18449 (N_18449,N_17682,N_17884);
nor U18450 (N_18450,N_17535,N_17821);
nand U18451 (N_18451,N_17601,N_17639);
or U18452 (N_18452,N_17664,N_17538);
xnor U18453 (N_18453,N_17537,N_17899);
or U18454 (N_18454,N_17752,N_17879);
nor U18455 (N_18455,N_17538,N_17585);
or U18456 (N_18456,N_17695,N_17590);
nor U18457 (N_18457,N_17665,N_17858);
nand U18458 (N_18458,N_17961,N_17812);
nor U18459 (N_18459,N_17513,N_17957);
and U18460 (N_18460,N_17881,N_17542);
and U18461 (N_18461,N_17648,N_17835);
and U18462 (N_18462,N_17800,N_17857);
or U18463 (N_18463,N_17644,N_17615);
nor U18464 (N_18464,N_17556,N_17547);
and U18465 (N_18465,N_17882,N_17911);
nor U18466 (N_18466,N_17836,N_17569);
nand U18467 (N_18467,N_17588,N_17763);
or U18468 (N_18468,N_17675,N_17707);
xnor U18469 (N_18469,N_17762,N_17657);
and U18470 (N_18470,N_17829,N_17726);
xnor U18471 (N_18471,N_17686,N_17504);
nor U18472 (N_18472,N_17927,N_17658);
xor U18473 (N_18473,N_17627,N_17572);
nor U18474 (N_18474,N_17828,N_17849);
nor U18475 (N_18475,N_17640,N_17603);
and U18476 (N_18476,N_17930,N_17615);
nor U18477 (N_18477,N_17916,N_17913);
or U18478 (N_18478,N_17680,N_17610);
xor U18479 (N_18479,N_17637,N_17903);
nand U18480 (N_18480,N_17759,N_17569);
and U18481 (N_18481,N_17616,N_17618);
or U18482 (N_18482,N_17905,N_17815);
nand U18483 (N_18483,N_17714,N_17547);
and U18484 (N_18484,N_17766,N_17775);
nor U18485 (N_18485,N_17560,N_17891);
or U18486 (N_18486,N_17999,N_17984);
xor U18487 (N_18487,N_17634,N_17798);
or U18488 (N_18488,N_17993,N_17679);
nor U18489 (N_18489,N_17927,N_17699);
xor U18490 (N_18490,N_17574,N_17531);
and U18491 (N_18491,N_17712,N_17616);
xnor U18492 (N_18492,N_17612,N_17936);
and U18493 (N_18493,N_17916,N_17828);
xor U18494 (N_18494,N_17968,N_17528);
nor U18495 (N_18495,N_17938,N_17677);
nand U18496 (N_18496,N_17785,N_17910);
nor U18497 (N_18497,N_17724,N_17646);
or U18498 (N_18498,N_17522,N_17580);
and U18499 (N_18499,N_17811,N_17605);
nor U18500 (N_18500,N_18233,N_18479);
nand U18501 (N_18501,N_18168,N_18426);
or U18502 (N_18502,N_18107,N_18259);
and U18503 (N_18503,N_18280,N_18494);
xor U18504 (N_18504,N_18030,N_18279);
nor U18505 (N_18505,N_18047,N_18065);
nand U18506 (N_18506,N_18173,N_18491);
nor U18507 (N_18507,N_18268,N_18048);
nand U18508 (N_18508,N_18131,N_18347);
xnor U18509 (N_18509,N_18123,N_18358);
or U18510 (N_18510,N_18484,N_18196);
nor U18511 (N_18511,N_18006,N_18086);
or U18512 (N_18512,N_18264,N_18341);
or U18513 (N_18513,N_18142,N_18410);
or U18514 (N_18514,N_18012,N_18138);
nor U18515 (N_18515,N_18066,N_18143);
nand U18516 (N_18516,N_18291,N_18482);
nor U18517 (N_18517,N_18325,N_18079);
and U18518 (N_18518,N_18407,N_18275);
nor U18519 (N_18519,N_18191,N_18054);
and U18520 (N_18520,N_18496,N_18492);
and U18521 (N_18521,N_18405,N_18366);
or U18522 (N_18522,N_18369,N_18078);
and U18523 (N_18523,N_18331,N_18056);
and U18524 (N_18524,N_18103,N_18424);
nor U18525 (N_18525,N_18081,N_18292);
and U18526 (N_18526,N_18069,N_18318);
xnor U18527 (N_18527,N_18240,N_18256);
or U18528 (N_18528,N_18155,N_18184);
nand U18529 (N_18529,N_18288,N_18321);
xnor U18530 (N_18530,N_18149,N_18043);
nor U18531 (N_18531,N_18285,N_18283);
xor U18532 (N_18532,N_18017,N_18214);
nand U18533 (N_18533,N_18448,N_18339);
nor U18534 (N_18534,N_18013,N_18216);
and U18535 (N_18535,N_18073,N_18402);
nor U18536 (N_18536,N_18229,N_18174);
or U18537 (N_18537,N_18170,N_18190);
nand U18538 (N_18538,N_18286,N_18238);
nand U18539 (N_18539,N_18476,N_18436);
xor U18540 (N_18540,N_18414,N_18367);
xor U18541 (N_18541,N_18129,N_18175);
nand U18542 (N_18542,N_18092,N_18258);
and U18543 (N_18543,N_18307,N_18437);
or U18544 (N_18544,N_18004,N_18446);
xor U18545 (N_18545,N_18120,N_18154);
nand U18546 (N_18546,N_18209,N_18024);
nor U18547 (N_18547,N_18419,N_18261);
or U18548 (N_18548,N_18421,N_18139);
nor U18549 (N_18549,N_18222,N_18248);
xnor U18550 (N_18550,N_18212,N_18281);
nor U18551 (N_18551,N_18035,N_18376);
or U18552 (N_18552,N_18187,N_18117);
nor U18553 (N_18553,N_18353,N_18311);
and U18554 (N_18554,N_18406,N_18045);
nand U18555 (N_18555,N_18374,N_18062);
and U18556 (N_18556,N_18343,N_18213);
xnor U18557 (N_18557,N_18300,N_18433);
or U18558 (N_18558,N_18228,N_18007);
or U18559 (N_18559,N_18096,N_18443);
and U18560 (N_18560,N_18019,N_18005);
or U18561 (N_18561,N_18093,N_18237);
nand U18562 (N_18562,N_18157,N_18176);
nand U18563 (N_18563,N_18221,N_18127);
xnor U18564 (N_18564,N_18051,N_18461);
xor U18565 (N_18565,N_18322,N_18152);
xnor U18566 (N_18566,N_18392,N_18334);
nand U18567 (N_18567,N_18136,N_18385);
or U18568 (N_18568,N_18317,N_18350);
nand U18569 (N_18569,N_18379,N_18162);
xor U18570 (N_18570,N_18098,N_18113);
nor U18571 (N_18571,N_18408,N_18247);
nand U18572 (N_18572,N_18038,N_18359);
and U18573 (N_18573,N_18297,N_18468);
nand U18574 (N_18574,N_18390,N_18135);
nand U18575 (N_18575,N_18000,N_18373);
or U18576 (N_18576,N_18220,N_18206);
xnor U18577 (N_18577,N_18284,N_18420);
nor U18578 (N_18578,N_18011,N_18119);
nor U18579 (N_18579,N_18395,N_18160);
or U18580 (N_18580,N_18380,N_18074);
or U18581 (N_18581,N_18460,N_18179);
or U18582 (N_18582,N_18046,N_18418);
or U18583 (N_18583,N_18346,N_18106);
nor U18584 (N_18584,N_18486,N_18452);
nand U18585 (N_18585,N_18287,N_18188);
and U18586 (N_18586,N_18391,N_18145);
xnor U18587 (N_18587,N_18198,N_18088);
nand U18588 (N_18588,N_18050,N_18147);
nor U18589 (N_18589,N_18029,N_18208);
nand U18590 (N_18590,N_18203,N_18301);
nor U18591 (N_18591,N_18355,N_18197);
or U18592 (N_18592,N_18032,N_18466);
or U18593 (N_18593,N_18052,N_18267);
xor U18594 (N_18594,N_18072,N_18417);
nor U18595 (N_18595,N_18388,N_18277);
nand U18596 (N_18596,N_18495,N_18332);
or U18597 (N_18597,N_18014,N_18276);
or U18598 (N_18598,N_18403,N_18262);
xnor U18599 (N_18599,N_18485,N_18413);
or U18600 (N_18600,N_18178,N_18025);
xor U18601 (N_18601,N_18348,N_18219);
and U18602 (N_18602,N_18039,N_18167);
xor U18603 (N_18603,N_18001,N_18272);
and U18604 (N_18604,N_18112,N_18368);
and U18605 (N_18605,N_18378,N_18021);
and U18606 (N_18606,N_18450,N_18389);
xor U18607 (N_18607,N_18010,N_18180);
and U18608 (N_18608,N_18067,N_18393);
and U18609 (N_18609,N_18016,N_18440);
nand U18610 (N_18610,N_18303,N_18034);
and U18611 (N_18611,N_18314,N_18161);
nand U18612 (N_18612,N_18090,N_18163);
xnor U18613 (N_18613,N_18200,N_18249);
or U18614 (N_18614,N_18320,N_18058);
or U18615 (N_18615,N_18431,N_18449);
nand U18616 (N_18616,N_18061,N_18333);
or U18617 (N_18617,N_18386,N_18327);
xnor U18618 (N_18618,N_18257,N_18077);
nor U18619 (N_18619,N_18159,N_18422);
nand U18620 (N_18620,N_18454,N_18265);
xor U18621 (N_18621,N_18121,N_18429);
xor U18622 (N_18622,N_18095,N_18171);
and U18623 (N_18623,N_18499,N_18441);
and U18624 (N_18624,N_18101,N_18246);
xnor U18625 (N_18625,N_18250,N_18108);
xnor U18626 (N_18626,N_18289,N_18370);
nand U18627 (N_18627,N_18002,N_18068);
xnor U18628 (N_18628,N_18076,N_18478);
xnor U18629 (N_18629,N_18083,N_18415);
or U18630 (N_18630,N_18362,N_18204);
nor U18631 (N_18631,N_18158,N_18344);
nand U18632 (N_18632,N_18445,N_18111);
or U18633 (N_18633,N_18309,N_18104);
nand U18634 (N_18634,N_18224,N_18266);
or U18635 (N_18635,N_18207,N_18401);
or U18636 (N_18636,N_18472,N_18263);
xnor U18637 (N_18637,N_18412,N_18215);
nor U18638 (N_18638,N_18130,N_18202);
nor U18639 (N_18639,N_18141,N_18126);
nor U18640 (N_18640,N_18185,N_18453);
xor U18641 (N_18641,N_18022,N_18467);
nand U18642 (N_18642,N_18336,N_18470);
nand U18643 (N_18643,N_18447,N_18040);
and U18644 (N_18644,N_18278,N_18352);
or U18645 (N_18645,N_18324,N_18457);
or U18646 (N_18646,N_18244,N_18225);
nor U18647 (N_18647,N_18455,N_18236);
xnor U18648 (N_18648,N_18340,N_18140);
xor U18649 (N_18649,N_18316,N_18269);
nand U18650 (N_18650,N_18243,N_18471);
nor U18651 (N_18651,N_18337,N_18254);
and U18652 (N_18652,N_18381,N_18458);
xor U18653 (N_18653,N_18153,N_18308);
or U18654 (N_18654,N_18349,N_18489);
nand U18655 (N_18655,N_18148,N_18084);
or U18656 (N_18656,N_18335,N_18464);
or U18657 (N_18657,N_18328,N_18293);
xnor U18658 (N_18658,N_18481,N_18399);
and U18659 (N_18659,N_18430,N_18356);
or U18660 (N_18660,N_18432,N_18169);
xor U18661 (N_18661,N_18037,N_18463);
nor U18662 (N_18662,N_18094,N_18082);
nand U18663 (N_18663,N_18384,N_18015);
or U18664 (N_18664,N_18055,N_18306);
xnor U18665 (N_18665,N_18151,N_18313);
and U18666 (N_18666,N_18427,N_18114);
and U18667 (N_18667,N_18326,N_18226);
or U18668 (N_18668,N_18156,N_18128);
and U18669 (N_18669,N_18294,N_18396);
xor U18670 (N_18670,N_18315,N_18211);
and U18671 (N_18671,N_18490,N_18080);
nand U18672 (N_18672,N_18363,N_18473);
nor U18673 (N_18673,N_18387,N_18164);
and U18674 (N_18674,N_18255,N_18053);
nand U18675 (N_18675,N_18118,N_18020);
nor U18676 (N_18676,N_18223,N_18097);
or U18677 (N_18677,N_18439,N_18234);
xor U18678 (N_18678,N_18195,N_18245);
xnor U18679 (N_18679,N_18330,N_18282);
and U18680 (N_18680,N_18230,N_18444);
nand U18681 (N_18681,N_18323,N_18271);
or U18682 (N_18682,N_18239,N_18398);
nor U18683 (N_18683,N_18109,N_18122);
nor U18684 (N_18684,N_18456,N_18009);
nand U18685 (N_18685,N_18205,N_18181);
nand U18686 (N_18686,N_18372,N_18260);
xnor U18687 (N_18687,N_18382,N_18199);
and U18688 (N_18688,N_18302,N_18137);
xor U18689 (N_18689,N_18060,N_18218);
nor U18690 (N_18690,N_18274,N_18342);
or U18691 (N_18691,N_18028,N_18360);
nand U18692 (N_18692,N_18150,N_18089);
and U18693 (N_18693,N_18227,N_18475);
xor U18694 (N_18694,N_18361,N_18134);
nor U18695 (N_18695,N_18428,N_18033);
nand U18696 (N_18696,N_18310,N_18049);
nand U18697 (N_18697,N_18304,N_18469);
or U18698 (N_18698,N_18099,N_18442);
xor U18699 (N_18699,N_18351,N_18183);
nor U18700 (N_18700,N_18085,N_18091);
xnor U18701 (N_18701,N_18100,N_18345);
nand U18702 (N_18702,N_18071,N_18409);
or U18703 (N_18703,N_18493,N_18057);
nand U18704 (N_18704,N_18296,N_18365);
and U18705 (N_18705,N_18319,N_18008);
xnor U18706 (N_18706,N_18115,N_18252);
xor U18707 (N_18707,N_18383,N_18416);
or U18708 (N_18708,N_18299,N_18124);
nor U18709 (N_18709,N_18044,N_18063);
or U18710 (N_18710,N_18498,N_18177);
or U18711 (N_18711,N_18102,N_18474);
xor U18712 (N_18712,N_18193,N_18423);
or U18713 (N_18713,N_18400,N_18210);
xor U18714 (N_18714,N_18394,N_18497);
nor U18715 (N_18715,N_18438,N_18459);
nor U18716 (N_18716,N_18031,N_18480);
xor U18717 (N_18717,N_18251,N_18377);
and U18718 (N_18718,N_18087,N_18338);
nand U18719 (N_18719,N_18003,N_18026);
xor U18720 (N_18720,N_18023,N_18146);
xnor U18721 (N_18721,N_18404,N_18273);
nor U18722 (N_18722,N_18435,N_18477);
or U18723 (N_18723,N_18371,N_18166);
and U18724 (N_18724,N_18242,N_18364);
or U18725 (N_18725,N_18434,N_18192);
or U18726 (N_18726,N_18375,N_18041);
or U18727 (N_18727,N_18465,N_18132);
and U18728 (N_18728,N_18232,N_18305);
or U18729 (N_18729,N_18036,N_18217);
nor U18730 (N_18730,N_18075,N_18064);
and U18731 (N_18731,N_18133,N_18295);
nor U18732 (N_18732,N_18018,N_18165);
and U18733 (N_18733,N_18354,N_18270);
and U18734 (N_18734,N_18290,N_18172);
and U18735 (N_18735,N_18194,N_18487);
nand U18736 (N_18736,N_18027,N_18059);
xor U18737 (N_18737,N_18105,N_18241);
or U18738 (N_18738,N_18425,N_18253);
nand U18739 (N_18739,N_18235,N_18144);
xor U18740 (N_18740,N_18451,N_18070);
nand U18741 (N_18741,N_18110,N_18231);
xnor U18742 (N_18742,N_18182,N_18397);
nand U18743 (N_18743,N_18116,N_18125);
or U18744 (N_18744,N_18298,N_18201);
nor U18745 (N_18745,N_18483,N_18312);
or U18746 (N_18746,N_18186,N_18042);
xor U18747 (N_18747,N_18411,N_18488);
nor U18748 (N_18748,N_18357,N_18462);
nand U18749 (N_18749,N_18329,N_18189);
xnor U18750 (N_18750,N_18145,N_18020);
or U18751 (N_18751,N_18370,N_18025);
nor U18752 (N_18752,N_18356,N_18165);
nand U18753 (N_18753,N_18211,N_18360);
nand U18754 (N_18754,N_18290,N_18198);
and U18755 (N_18755,N_18049,N_18007);
or U18756 (N_18756,N_18464,N_18284);
nand U18757 (N_18757,N_18171,N_18430);
nor U18758 (N_18758,N_18125,N_18103);
nand U18759 (N_18759,N_18379,N_18354);
xnor U18760 (N_18760,N_18016,N_18158);
nand U18761 (N_18761,N_18343,N_18032);
and U18762 (N_18762,N_18389,N_18142);
and U18763 (N_18763,N_18339,N_18220);
nor U18764 (N_18764,N_18383,N_18337);
nand U18765 (N_18765,N_18211,N_18146);
or U18766 (N_18766,N_18314,N_18220);
nand U18767 (N_18767,N_18200,N_18218);
xnor U18768 (N_18768,N_18031,N_18414);
and U18769 (N_18769,N_18228,N_18044);
nor U18770 (N_18770,N_18126,N_18361);
nand U18771 (N_18771,N_18232,N_18494);
or U18772 (N_18772,N_18425,N_18196);
xor U18773 (N_18773,N_18362,N_18469);
xor U18774 (N_18774,N_18356,N_18247);
nor U18775 (N_18775,N_18400,N_18356);
nor U18776 (N_18776,N_18261,N_18334);
and U18777 (N_18777,N_18373,N_18295);
xnor U18778 (N_18778,N_18183,N_18212);
nand U18779 (N_18779,N_18468,N_18475);
xnor U18780 (N_18780,N_18115,N_18297);
and U18781 (N_18781,N_18231,N_18472);
nand U18782 (N_18782,N_18001,N_18193);
and U18783 (N_18783,N_18005,N_18379);
and U18784 (N_18784,N_18369,N_18200);
or U18785 (N_18785,N_18445,N_18259);
nor U18786 (N_18786,N_18016,N_18177);
or U18787 (N_18787,N_18071,N_18162);
nand U18788 (N_18788,N_18333,N_18017);
xnor U18789 (N_18789,N_18177,N_18378);
and U18790 (N_18790,N_18303,N_18329);
nor U18791 (N_18791,N_18178,N_18167);
xor U18792 (N_18792,N_18492,N_18391);
xor U18793 (N_18793,N_18049,N_18020);
nor U18794 (N_18794,N_18082,N_18458);
nor U18795 (N_18795,N_18478,N_18214);
and U18796 (N_18796,N_18116,N_18135);
or U18797 (N_18797,N_18479,N_18413);
nor U18798 (N_18798,N_18342,N_18372);
nand U18799 (N_18799,N_18197,N_18308);
nand U18800 (N_18800,N_18462,N_18018);
and U18801 (N_18801,N_18233,N_18180);
xnor U18802 (N_18802,N_18103,N_18455);
and U18803 (N_18803,N_18303,N_18046);
nor U18804 (N_18804,N_18030,N_18052);
or U18805 (N_18805,N_18420,N_18219);
nand U18806 (N_18806,N_18155,N_18430);
and U18807 (N_18807,N_18222,N_18474);
nor U18808 (N_18808,N_18237,N_18434);
xor U18809 (N_18809,N_18279,N_18352);
and U18810 (N_18810,N_18492,N_18498);
and U18811 (N_18811,N_18238,N_18028);
nor U18812 (N_18812,N_18494,N_18214);
nor U18813 (N_18813,N_18025,N_18005);
xor U18814 (N_18814,N_18123,N_18130);
or U18815 (N_18815,N_18346,N_18495);
nand U18816 (N_18816,N_18022,N_18322);
nor U18817 (N_18817,N_18219,N_18078);
or U18818 (N_18818,N_18054,N_18077);
or U18819 (N_18819,N_18228,N_18085);
or U18820 (N_18820,N_18014,N_18382);
and U18821 (N_18821,N_18218,N_18013);
nand U18822 (N_18822,N_18288,N_18300);
or U18823 (N_18823,N_18300,N_18285);
xor U18824 (N_18824,N_18469,N_18035);
xnor U18825 (N_18825,N_18009,N_18323);
and U18826 (N_18826,N_18125,N_18158);
nand U18827 (N_18827,N_18251,N_18424);
or U18828 (N_18828,N_18450,N_18022);
xor U18829 (N_18829,N_18388,N_18270);
xor U18830 (N_18830,N_18136,N_18474);
nor U18831 (N_18831,N_18040,N_18301);
nand U18832 (N_18832,N_18160,N_18350);
nand U18833 (N_18833,N_18434,N_18251);
nor U18834 (N_18834,N_18140,N_18361);
nand U18835 (N_18835,N_18432,N_18170);
or U18836 (N_18836,N_18484,N_18480);
nor U18837 (N_18837,N_18015,N_18447);
or U18838 (N_18838,N_18349,N_18066);
and U18839 (N_18839,N_18223,N_18177);
nor U18840 (N_18840,N_18168,N_18136);
xnor U18841 (N_18841,N_18489,N_18240);
and U18842 (N_18842,N_18069,N_18209);
or U18843 (N_18843,N_18124,N_18087);
xor U18844 (N_18844,N_18299,N_18459);
xor U18845 (N_18845,N_18280,N_18026);
nor U18846 (N_18846,N_18423,N_18400);
or U18847 (N_18847,N_18138,N_18255);
and U18848 (N_18848,N_18333,N_18055);
nand U18849 (N_18849,N_18295,N_18438);
nor U18850 (N_18850,N_18389,N_18070);
nor U18851 (N_18851,N_18287,N_18215);
and U18852 (N_18852,N_18332,N_18138);
and U18853 (N_18853,N_18442,N_18454);
xnor U18854 (N_18854,N_18151,N_18438);
xor U18855 (N_18855,N_18156,N_18235);
nand U18856 (N_18856,N_18141,N_18312);
nand U18857 (N_18857,N_18343,N_18053);
nor U18858 (N_18858,N_18339,N_18468);
nand U18859 (N_18859,N_18058,N_18443);
and U18860 (N_18860,N_18030,N_18239);
or U18861 (N_18861,N_18448,N_18320);
and U18862 (N_18862,N_18205,N_18116);
and U18863 (N_18863,N_18477,N_18008);
nor U18864 (N_18864,N_18448,N_18442);
nand U18865 (N_18865,N_18024,N_18488);
and U18866 (N_18866,N_18166,N_18161);
nand U18867 (N_18867,N_18297,N_18418);
xnor U18868 (N_18868,N_18117,N_18138);
or U18869 (N_18869,N_18440,N_18297);
and U18870 (N_18870,N_18432,N_18035);
nand U18871 (N_18871,N_18404,N_18480);
nand U18872 (N_18872,N_18331,N_18218);
and U18873 (N_18873,N_18219,N_18473);
nand U18874 (N_18874,N_18145,N_18325);
nand U18875 (N_18875,N_18113,N_18008);
xor U18876 (N_18876,N_18275,N_18054);
and U18877 (N_18877,N_18352,N_18321);
xor U18878 (N_18878,N_18135,N_18250);
nand U18879 (N_18879,N_18182,N_18381);
xor U18880 (N_18880,N_18252,N_18319);
nand U18881 (N_18881,N_18388,N_18356);
nor U18882 (N_18882,N_18367,N_18188);
nand U18883 (N_18883,N_18340,N_18354);
xnor U18884 (N_18884,N_18447,N_18190);
nor U18885 (N_18885,N_18316,N_18285);
nand U18886 (N_18886,N_18358,N_18034);
xnor U18887 (N_18887,N_18032,N_18038);
nand U18888 (N_18888,N_18086,N_18166);
nor U18889 (N_18889,N_18144,N_18320);
or U18890 (N_18890,N_18157,N_18457);
nor U18891 (N_18891,N_18054,N_18237);
nor U18892 (N_18892,N_18155,N_18261);
nand U18893 (N_18893,N_18176,N_18392);
and U18894 (N_18894,N_18311,N_18006);
or U18895 (N_18895,N_18345,N_18244);
xor U18896 (N_18896,N_18143,N_18496);
or U18897 (N_18897,N_18343,N_18323);
or U18898 (N_18898,N_18102,N_18247);
nand U18899 (N_18899,N_18353,N_18113);
or U18900 (N_18900,N_18007,N_18268);
nor U18901 (N_18901,N_18140,N_18407);
nor U18902 (N_18902,N_18375,N_18188);
xor U18903 (N_18903,N_18193,N_18003);
nor U18904 (N_18904,N_18178,N_18416);
nor U18905 (N_18905,N_18085,N_18253);
xnor U18906 (N_18906,N_18427,N_18040);
nand U18907 (N_18907,N_18251,N_18026);
nand U18908 (N_18908,N_18020,N_18414);
xnor U18909 (N_18909,N_18168,N_18120);
and U18910 (N_18910,N_18043,N_18058);
or U18911 (N_18911,N_18225,N_18057);
and U18912 (N_18912,N_18497,N_18218);
xor U18913 (N_18913,N_18405,N_18282);
or U18914 (N_18914,N_18461,N_18124);
nand U18915 (N_18915,N_18348,N_18055);
nand U18916 (N_18916,N_18360,N_18187);
nor U18917 (N_18917,N_18449,N_18022);
and U18918 (N_18918,N_18346,N_18416);
nor U18919 (N_18919,N_18446,N_18000);
or U18920 (N_18920,N_18180,N_18408);
or U18921 (N_18921,N_18441,N_18272);
nor U18922 (N_18922,N_18380,N_18051);
xnor U18923 (N_18923,N_18441,N_18404);
or U18924 (N_18924,N_18013,N_18287);
nor U18925 (N_18925,N_18126,N_18159);
xnor U18926 (N_18926,N_18070,N_18288);
or U18927 (N_18927,N_18380,N_18443);
nor U18928 (N_18928,N_18478,N_18357);
and U18929 (N_18929,N_18250,N_18032);
nand U18930 (N_18930,N_18316,N_18343);
nor U18931 (N_18931,N_18011,N_18455);
nor U18932 (N_18932,N_18479,N_18014);
nor U18933 (N_18933,N_18441,N_18432);
or U18934 (N_18934,N_18421,N_18188);
and U18935 (N_18935,N_18424,N_18066);
or U18936 (N_18936,N_18354,N_18433);
and U18937 (N_18937,N_18465,N_18105);
or U18938 (N_18938,N_18390,N_18258);
nor U18939 (N_18939,N_18196,N_18089);
xnor U18940 (N_18940,N_18355,N_18142);
nor U18941 (N_18941,N_18174,N_18053);
and U18942 (N_18942,N_18229,N_18451);
and U18943 (N_18943,N_18232,N_18173);
nand U18944 (N_18944,N_18088,N_18035);
nor U18945 (N_18945,N_18245,N_18325);
and U18946 (N_18946,N_18349,N_18011);
nor U18947 (N_18947,N_18185,N_18210);
or U18948 (N_18948,N_18417,N_18021);
nand U18949 (N_18949,N_18087,N_18472);
nand U18950 (N_18950,N_18148,N_18437);
and U18951 (N_18951,N_18201,N_18498);
xnor U18952 (N_18952,N_18445,N_18158);
or U18953 (N_18953,N_18457,N_18375);
xor U18954 (N_18954,N_18031,N_18025);
or U18955 (N_18955,N_18075,N_18225);
xnor U18956 (N_18956,N_18028,N_18405);
xor U18957 (N_18957,N_18301,N_18309);
or U18958 (N_18958,N_18464,N_18230);
nand U18959 (N_18959,N_18487,N_18253);
xor U18960 (N_18960,N_18249,N_18269);
xnor U18961 (N_18961,N_18007,N_18328);
or U18962 (N_18962,N_18374,N_18386);
or U18963 (N_18963,N_18178,N_18228);
nand U18964 (N_18964,N_18420,N_18310);
and U18965 (N_18965,N_18362,N_18017);
nor U18966 (N_18966,N_18054,N_18321);
nor U18967 (N_18967,N_18354,N_18457);
xor U18968 (N_18968,N_18432,N_18213);
and U18969 (N_18969,N_18187,N_18241);
or U18970 (N_18970,N_18232,N_18322);
nor U18971 (N_18971,N_18081,N_18334);
or U18972 (N_18972,N_18184,N_18342);
nand U18973 (N_18973,N_18111,N_18243);
xnor U18974 (N_18974,N_18125,N_18292);
or U18975 (N_18975,N_18364,N_18010);
or U18976 (N_18976,N_18152,N_18434);
nand U18977 (N_18977,N_18465,N_18143);
xnor U18978 (N_18978,N_18311,N_18137);
nor U18979 (N_18979,N_18474,N_18081);
and U18980 (N_18980,N_18189,N_18031);
xor U18981 (N_18981,N_18044,N_18031);
nand U18982 (N_18982,N_18316,N_18450);
nand U18983 (N_18983,N_18402,N_18026);
xnor U18984 (N_18984,N_18306,N_18049);
or U18985 (N_18985,N_18399,N_18362);
nor U18986 (N_18986,N_18023,N_18114);
and U18987 (N_18987,N_18020,N_18130);
nand U18988 (N_18988,N_18452,N_18461);
and U18989 (N_18989,N_18356,N_18141);
nand U18990 (N_18990,N_18135,N_18429);
and U18991 (N_18991,N_18200,N_18168);
and U18992 (N_18992,N_18350,N_18109);
and U18993 (N_18993,N_18103,N_18385);
or U18994 (N_18994,N_18188,N_18380);
nand U18995 (N_18995,N_18327,N_18205);
nand U18996 (N_18996,N_18376,N_18246);
nor U18997 (N_18997,N_18235,N_18259);
and U18998 (N_18998,N_18356,N_18464);
nand U18999 (N_18999,N_18464,N_18431);
nand U19000 (N_19000,N_18610,N_18651);
and U19001 (N_19001,N_18933,N_18679);
nand U19002 (N_19002,N_18952,N_18881);
nor U19003 (N_19003,N_18694,N_18924);
and U19004 (N_19004,N_18565,N_18680);
and U19005 (N_19005,N_18577,N_18742);
and U19006 (N_19006,N_18678,N_18847);
or U19007 (N_19007,N_18698,N_18686);
nor U19008 (N_19008,N_18615,N_18510);
or U19009 (N_19009,N_18708,N_18997);
and U19010 (N_19010,N_18937,N_18515);
and U19011 (N_19011,N_18647,N_18544);
and U19012 (N_19012,N_18756,N_18971);
nand U19013 (N_19013,N_18690,N_18799);
and U19014 (N_19014,N_18725,N_18836);
xor U19015 (N_19015,N_18906,N_18913);
or U19016 (N_19016,N_18758,N_18511);
xor U19017 (N_19017,N_18957,N_18660);
nor U19018 (N_19018,N_18806,N_18585);
nor U19019 (N_19019,N_18837,N_18546);
xnor U19020 (N_19020,N_18814,N_18870);
and U19021 (N_19021,N_18523,N_18669);
nand U19022 (N_19022,N_18849,N_18960);
nand U19023 (N_19023,N_18797,N_18783);
nor U19024 (N_19024,N_18788,N_18695);
nor U19025 (N_19025,N_18872,N_18888);
and U19026 (N_19026,N_18662,N_18886);
and U19027 (N_19027,N_18588,N_18781);
nand U19028 (N_19028,N_18874,N_18639);
nand U19029 (N_19029,N_18689,N_18688);
xnor U19030 (N_19030,N_18782,N_18752);
or U19031 (N_19031,N_18699,N_18862);
xnor U19032 (N_19032,N_18999,N_18619);
nor U19033 (N_19033,N_18633,N_18815);
xnor U19034 (N_19034,N_18830,N_18606);
xnor U19035 (N_19035,N_18825,N_18851);
nand U19036 (N_19036,N_18640,N_18941);
or U19037 (N_19037,N_18967,N_18571);
xor U19038 (N_19038,N_18521,N_18779);
or U19039 (N_19039,N_18550,N_18575);
or U19040 (N_19040,N_18831,N_18902);
and U19041 (N_19041,N_18704,N_18900);
xnor U19042 (N_19042,N_18807,N_18744);
nor U19043 (N_19043,N_18921,N_18519);
or U19044 (N_19044,N_18590,N_18876);
and U19045 (N_19045,N_18734,N_18976);
and U19046 (N_19046,N_18987,N_18652);
or U19047 (N_19047,N_18721,N_18594);
nor U19048 (N_19048,N_18727,N_18828);
or U19049 (N_19049,N_18533,N_18580);
or U19050 (N_19050,N_18503,N_18697);
or U19051 (N_19051,N_18770,N_18599);
nand U19052 (N_19052,N_18790,N_18701);
xor U19053 (N_19053,N_18843,N_18848);
or U19054 (N_19054,N_18509,N_18573);
nand U19055 (N_19055,N_18659,N_18951);
nand U19056 (N_19056,N_18592,N_18853);
nor U19057 (N_19057,N_18589,N_18826);
nor U19058 (N_19058,N_18556,N_18930);
or U19059 (N_19059,N_18520,N_18560);
xor U19060 (N_19060,N_18798,N_18707);
nand U19061 (N_19061,N_18969,N_18731);
xnor U19062 (N_19062,N_18935,N_18932);
nor U19063 (N_19063,N_18959,N_18925);
or U19064 (N_19064,N_18526,N_18667);
nand U19065 (N_19065,N_18861,N_18859);
xor U19066 (N_19066,N_18841,N_18992);
nand U19067 (N_19067,N_18896,N_18608);
nor U19068 (N_19068,N_18893,N_18956);
nor U19069 (N_19069,N_18990,N_18961);
or U19070 (N_19070,N_18658,N_18978);
xnor U19071 (N_19071,N_18508,N_18674);
nor U19072 (N_19072,N_18844,N_18916);
and U19073 (N_19073,N_18622,N_18771);
xnor U19074 (N_19074,N_18789,N_18865);
or U19075 (N_19075,N_18739,N_18754);
or U19076 (N_19076,N_18824,N_18684);
and U19077 (N_19077,N_18795,N_18648);
xor U19078 (N_19078,N_18624,N_18671);
nor U19079 (N_19079,N_18703,N_18557);
nor U19080 (N_19080,N_18899,N_18512);
xor U19081 (N_19081,N_18813,N_18994);
nor U19082 (N_19082,N_18621,N_18747);
nand U19083 (N_19083,N_18532,N_18856);
xor U19084 (N_19084,N_18666,N_18551);
and U19085 (N_19085,N_18524,N_18778);
nand U19086 (N_19086,N_18904,N_18939);
nor U19087 (N_19087,N_18623,N_18500);
nand U19088 (N_19088,N_18661,N_18863);
and U19089 (N_19089,N_18953,N_18644);
nand U19090 (N_19090,N_18860,N_18772);
nor U19091 (N_19091,N_18948,N_18791);
xor U19092 (N_19092,N_18562,N_18784);
nor U19093 (N_19093,N_18943,N_18670);
and U19094 (N_19094,N_18794,N_18819);
nand U19095 (N_19095,N_18908,N_18709);
and U19096 (N_19096,N_18879,N_18609);
and U19097 (N_19097,N_18912,N_18922);
or U19098 (N_19098,N_18812,N_18683);
nor U19099 (N_19099,N_18832,N_18838);
nand U19100 (N_19100,N_18964,N_18522);
nor U19101 (N_19101,N_18950,N_18850);
nor U19102 (N_19102,N_18579,N_18940);
or U19103 (N_19103,N_18711,N_18685);
and U19104 (N_19104,N_18857,N_18517);
nor U19105 (N_19105,N_18567,N_18988);
xnor U19106 (N_19106,N_18545,N_18715);
nand U19107 (N_19107,N_18542,N_18883);
or U19108 (N_19108,N_18676,N_18616);
nand U19109 (N_19109,N_18966,N_18602);
or U19110 (N_19110,N_18705,N_18962);
nand U19111 (N_19111,N_18611,N_18975);
xnor U19112 (N_19112,N_18757,N_18586);
and U19113 (N_19113,N_18786,N_18839);
and U19114 (N_19114,N_18985,N_18581);
nand U19115 (N_19115,N_18852,N_18636);
and U19116 (N_19116,N_18563,N_18514);
nand U19117 (N_19117,N_18755,N_18834);
nor U19118 (N_19118,N_18954,N_18597);
or U19119 (N_19119,N_18820,N_18918);
xor U19120 (N_19120,N_18972,N_18726);
or U19121 (N_19121,N_18984,N_18891);
xnor U19122 (N_19122,N_18600,N_18657);
nand U19123 (N_19123,N_18822,N_18818);
nand U19124 (N_19124,N_18714,N_18561);
or U19125 (N_19125,N_18774,N_18958);
xor U19126 (N_19126,N_18808,N_18583);
nand U19127 (N_19127,N_18541,N_18724);
nor U19128 (N_19128,N_18973,N_18816);
xor U19129 (N_19129,N_18629,N_18760);
and U19130 (N_19130,N_18646,N_18869);
nand U19131 (N_19131,N_18693,N_18768);
nor U19132 (N_19132,N_18946,N_18570);
nand U19133 (N_19133,N_18846,N_18905);
or U19134 (N_19134,N_18991,N_18800);
and U19135 (N_19135,N_18549,N_18938);
nor U19136 (N_19136,N_18681,N_18655);
xor U19137 (N_19137,N_18665,N_18890);
or U19138 (N_19138,N_18927,N_18823);
and U19139 (N_19139,N_18894,N_18668);
nand U19140 (N_19140,N_18553,N_18801);
nor U19141 (N_19141,N_18885,N_18977);
nand U19142 (N_19142,N_18785,N_18802);
nand U19143 (N_19143,N_18910,N_18634);
nand U19144 (N_19144,N_18649,N_18735);
or U19145 (N_19145,N_18627,N_18745);
nor U19146 (N_19146,N_18817,N_18866);
and U19147 (N_19147,N_18787,N_18982);
xnor U19148 (N_19148,N_18664,N_18777);
and U19149 (N_19149,N_18793,N_18591);
and U19150 (N_19150,N_18717,N_18539);
nor U19151 (N_19151,N_18730,N_18867);
xor U19152 (N_19152,N_18963,N_18620);
xor U19153 (N_19153,N_18626,N_18687);
nand U19154 (N_19154,N_18568,N_18965);
and U19155 (N_19155,N_18773,N_18766);
nand U19156 (N_19156,N_18759,N_18700);
xnor U19157 (N_19157,N_18871,N_18746);
xor U19158 (N_19158,N_18507,N_18552);
nor U19159 (N_19159,N_18702,N_18617);
or U19160 (N_19160,N_18829,N_18566);
and U19161 (N_19161,N_18716,N_18907);
or U19162 (N_19162,N_18696,N_18897);
or U19163 (N_19163,N_18877,N_18596);
xnor U19164 (N_19164,N_18536,N_18628);
xnor U19165 (N_19165,N_18706,N_18873);
and U19166 (N_19166,N_18564,N_18656);
nor U19167 (N_19167,N_18638,N_18605);
and U19168 (N_19168,N_18672,N_18811);
xnor U19169 (N_19169,N_18543,N_18914);
nor U19170 (N_19170,N_18713,N_18947);
xnor U19171 (N_19171,N_18677,N_18538);
nand U19172 (N_19172,N_18722,N_18569);
nor U19173 (N_19173,N_18981,N_18614);
nor U19174 (N_19174,N_18949,N_18555);
or U19175 (N_19175,N_18574,N_18528);
and U19176 (N_19176,N_18632,N_18810);
xnor U19177 (N_19177,N_18682,N_18736);
nand U19178 (N_19178,N_18955,N_18673);
nor U19179 (N_19179,N_18601,N_18986);
nand U19180 (N_19180,N_18931,N_18898);
nand U19181 (N_19181,N_18740,N_18604);
and U19182 (N_19182,N_18733,N_18753);
nor U19183 (N_19183,N_18767,N_18920);
xnor U19184 (N_19184,N_18548,N_18980);
nor U19185 (N_19185,N_18979,N_18547);
and U19186 (N_19186,N_18710,N_18880);
xor U19187 (N_19187,N_18527,N_18607);
or U19188 (N_19188,N_18554,N_18875);
xor U19189 (N_19189,N_18827,N_18559);
and U19190 (N_19190,N_18926,N_18692);
or U19191 (N_19191,N_18723,N_18804);
nand U19192 (N_19192,N_18720,N_18530);
nor U19193 (N_19193,N_18942,N_18712);
and U19194 (N_19194,N_18765,N_18637);
nor U19195 (N_19195,N_18582,N_18663);
xnor U19196 (N_19196,N_18518,N_18970);
and U19197 (N_19197,N_18803,N_18595);
or U19198 (N_19198,N_18968,N_18641);
or U19199 (N_19199,N_18506,N_18944);
xor U19200 (N_19200,N_18749,N_18780);
nand U19201 (N_19201,N_18809,N_18895);
and U19202 (N_19202,N_18998,N_18558);
xnor U19203 (N_19203,N_18625,N_18855);
xnor U19204 (N_19204,N_18796,N_18501);
nor U19205 (N_19205,N_18993,N_18593);
xnor U19206 (N_19206,N_18928,N_18776);
nor U19207 (N_19207,N_18653,N_18738);
xnor U19208 (N_19208,N_18729,N_18936);
nor U19209 (N_19209,N_18833,N_18761);
xnor U19210 (N_19210,N_18909,N_18917);
or U19211 (N_19211,N_18878,N_18901);
or U19212 (N_19212,N_18635,N_18650);
or U19213 (N_19213,N_18525,N_18540);
xor U19214 (N_19214,N_18882,N_18572);
or U19215 (N_19215,N_18645,N_18630);
and U19216 (N_19216,N_18983,N_18643);
nor U19217 (N_19217,N_18989,N_18613);
nor U19218 (N_19218,N_18743,N_18792);
and U19219 (N_19219,N_18654,N_18762);
nand U19220 (N_19220,N_18864,N_18842);
nor U19221 (N_19221,N_18732,N_18513);
or U19222 (N_19222,N_18889,N_18892);
nor U19223 (N_19223,N_18858,N_18884);
nor U19224 (N_19224,N_18718,N_18576);
nor U19225 (N_19225,N_18868,N_18502);
or U19226 (N_19226,N_18775,N_18835);
or U19227 (N_19227,N_18769,N_18750);
and U19228 (N_19228,N_18763,N_18534);
xnor U19229 (N_19229,N_18911,N_18631);
nand U19230 (N_19230,N_18537,N_18516);
or U19231 (N_19231,N_18691,N_18719);
xor U19232 (N_19232,N_18974,N_18529);
nand U19233 (N_19233,N_18805,N_18505);
nand U19234 (N_19234,N_18603,N_18587);
and U19235 (N_19235,N_18995,N_18531);
xnor U19236 (N_19236,N_18923,N_18612);
xor U19237 (N_19237,N_18929,N_18748);
nor U19238 (N_19238,N_18903,N_18821);
xor U19239 (N_19239,N_18764,N_18578);
nand U19240 (N_19240,N_18741,N_18535);
nor U19241 (N_19241,N_18945,N_18854);
xor U19242 (N_19242,N_18919,N_18737);
nor U19243 (N_19243,N_18584,N_18887);
and U19244 (N_19244,N_18598,N_18996);
xnor U19245 (N_19245,N_18675,N_18934);
nor U19246 (N_19246,N_18504,N_18728);
or U19247 (N_19247,N_18642,N_18751);
and U19248 (N_19248,N_18840,N_18618);
or U19249 (N_19249,N_18845,N_18915);
nand U19250 (N_19250,N_18922,N_18738);
and U19251 (N_19251,N_18937,N_18959);
xnor U19252 (N_19252,N_18629,N_18545);
nor U19253 (N_19253,N_18679,N_18673);
or U19254 (N_19254,N_18997,N_18859);
xor U19255 (N_19255,N_18852,N_18830);
and U19256 (N_19256,N_18801,N_18762);
or U19257 (N_19257,N_18850,N_18984);
nand U19258 (N_19258,N_18873,N_18571);
nor U19259 (N_19259,N_18968,N_18502);
and U19260 (N_19260,N_18686,N_18938);
and U19261 (N_19261,N_18818,N_18756);
or U19262 (N_19262,N_18578,N_18502);
or U19263 (N_19263,N_18858,N_18597);
xor U19264 (N_19264,N_18936,N_18564);
xor U19265 (N_19265,N_18548,N_18703);
xor U19266 (N_19266,N_18706,N_18840);
xor U19267 (N_19267,N_18901,N_18580);
or U19268 (N_19268,N_18699,N_18525);
and U19269 (N_19269,N_18654,N_18897);
xor U19270 (N_19270,N_18823,N_18856);
nand U19271 (N_19271,N_18926,N_18582);
or U19272 (N_19272,N_18589,N_18604);
nand U19273 (N_19273,N_18891,N_18872);
nor U19274 (N_19274,N_18552,N_18533);
nand U19275 (N_19275,N_18796,N_18614);
nand U19276 (N_19276,N_18535,N_18577);
xnor U19277 (N_19277,N_18923,N_18690);
and U19278 (N_19278,N_18900,N_18542);
nand U19279 (N_19279,N_18520,N_18863);
and U19280 (N_19280,N_18819,N_18547);
xor U19281 (N_19281,N_18748,N_18992);
nand U19282 (N_19282,N_18934,N_18702);
and U19283 (N_19283,N_18546,N_18980);
nor U19284 (N_19284,N_18500,N_18710);
or U19285 (N_19285,N_18987,N_18719);
and U19286 (N_19286,N_18627,N_18626);
nor U19287 (N_19287,N_18981,N_18829);
xnor U19288 (N_19288,N_18855,N_18741);
or U19289 (N_19289,N_18592,N_18706);
and U19290 (N_19290,N_18988,N_18512);
or U19291 (N_19291,N_18762,N_18775);
nor U19292 (N_19292,N_18817,N_18659);
and U19293 (N_19293,N_18552,N_18730);
nand U19294 (N_19294,N_18642,N_18860);
or U19295 (N_19295,N_18838,N_18621);
or U19296 (N_19296,N_18815,N_18601);
xnor U19297 (N_19297,N_18733,N_18779);
or U19298 (N_19298,N_18659,N_18935);
nand U19299 (N_19299,N_18733,N_18923);
xor U19300 (N_19300,N_18739,N_18795);
and U19301 (N_19301,N_18522,N_18652);
nor U19302 (N_19302,N_18767,N_18792);
or U19303 (N_19303,N_18649,N_18780);
nor U19304 (N_19304,N_18968,N_18529);
or U19305 (N_19305,N_18630,N_18555);
nor U19306 (N_19306,N_18629,N_18888);
xnor U19307 (N_19307,N_18987,N_18630);
xnor U19308 (N_19308,N_18519,N_18878);
and U19309 (N_19309,N_18550,N_18696);
nand U19310 (N_19310,N_18944,N_18720);
or U19311 (N_19311,N_18642,N_18667);
nand U19312 (N_19312,N_18547,N_18553);
nor U19313 (N_19313,N_18715,N_18790);
xnor U19314 (N_19314,N_18845,N_18631);
nor U19315 (N_19315,N_18968,N_18716);
nand U19316 (N_19316,N_18881,N_18918);
nor U19317 (N_19317,N_18587,N_18636);
xnor U19318 (N_19318,N_18566,N_18826);
and U19319 (N_19319,N_18948,N_18816);
nor U19320 (N_19320,N_18729,N_18976);
or U19321 (N_19321,N_18602,N_18757);
nand U19322 (N_19322,N_18738,N_18659);
or U19323 (N_19323,N_18635,N_18947);
or U19324 (N_19324,N_18524,N_18692);
or U19325 (N_19325,N_18611,N_18893);
xnor U19326 (N_19326,N_18700,N_18572);
nor U19327 (N_19327,N_18993,N_18652);
xor U19328 (N_19328,N_18653,N_18627);
nor U19329 (N_19329,N_18903,N_18886);
nand U19330 (N_19330,N_18704,N_18816);
nor U19331 (N_19331,N_18805,N_18976);
or U19332 (N_19332,N_18920,N_18814);
or U19333 (N_19333,N_18530,N_18704);
nand U19334 (N_19334,N_18764,N_18585);
nor U19335 (N_19335,N_18507,N_18907);
nand U19336 (N_19336,N_18740,N_18760);
xnor U19337 (N_19337,N_18532,N_18978);
or U19338 (N_19338,N_18738,N_18588);
nand U19339 (N_19339,N_18767,N_18633);
xor U19340 (N_19340,N_18627,N_18618);
and U19341 (N_19341,N_18884,N_18714);
nor U19342 (N_19342,N_18591,N_18556);
nor U19343 (N_19343,N_18527,N_18576);
or U19344 (N_19344,N_18595,N_18677);
nor U19345 (N_19345,N_18841,N_18933);
and U19346 (N_19346,N_18758,N_18937);
nand U19347 (N_19347,N_18612,N_18876);
and U19348 (N_19348,N_18567,N_18585);
and U19349 (N_19349,N_18642,N_18604);
or U19350 (N_19350,N_18880,N_18566);
or U19351 (N_19351,N_18701,N_18635);
or U19352 (N_19352,N_18914,N_18803);
and U19353 (N_19353,N_18952,N_18617);
nor U19354 (N_19354,N_18965,N_18870);
nand U19355 (N_19355,N_18891,N_18804);
nand U19356 (N_19356,N_18660,N_18868);
nand U19357 (N_19357,N_18626,N_18595);
nor U19358 (N_19358,N_18542,N_18848);
nand U19359 (N_19359,N_18686,N_18652);
or U19360 (N_19360,N_18502,N_18833);
nand U19361 (N_19361,N_18821,N_18932);
and U19362 (N_19362,N_18831,N_18629);
nand U19363 (N_19363,N_18741,N_18746);
xor U19364 (N_19364,N_18693,N_18668);
nand U19365 (N_19365,N_18979,N_18545);
and U19366 (N_19366,N_18669,N_18843);
nand U19367 (N_19367,N_18702,N_18611);
and U19368 (N_19368,N_18980,N_18902);
nand U19369 (N_19369,N_18530,N_18612);
or U19370 (N_19370,N_18700,N_18914);
or U19371 (N_19371,N_18951,N_18876);
and U19372 (N_19372,N_18554,N_18775);
nor U19373 (N_19373,N_18841,N_18854);
or U19374 (N_19374,N_18877,N_18850);
xor U19375 (N_19375,N_18726,N_18596);
or U19376 (N_19376,N_18773,N_18507);
nor U19377 (N_19377,N_18504,N_18847);
xor U19378 (N_19378,N_18946,N_18714);
xor U19379 (N_19379,N_18715,N_18534);
xor U19380 (N_19380,N_18870,N_18904);
or U19381 (N_19381,N_18676,N_18570);
nand U19382 (N_19382,N_18734,N_18507);
xor U19383 (N_19383,N_18872,N_18542);
and U19384 (N_19384,N_18660,N_18559);
nand U19385 (N_19385,N_18962,N_18975);
or U19386 (N_19386,N_18905,N_18683);
nand U19387 (N_19387,N_18757,N_18892);
and U19388 (N_19388,N_18720,N_18514);
nor U19389 (N_19389,N_18676,N_18983);
nand U19390 (N_19390,N_18530,N_18685);
nor U19391 (N_19391,N_18882,N_18542);
and U19392 (N_19392,N_18552,N_18953);
xor U19393 (N_19393,N_18944,N_18930);
and U19394 (N_19394,N_18828,N_18788);
nand U19395 (N_19395,N_18541,N_18798);
or U19396 (N_19396,N_18636,N_18903);
nand U19397 (N_19397,N_18617,N_18984);
nor U19398 (N_19398,N_18807,N_18504);
and U19399 (N_19399,N_18582,N_18940);
and U19400 (N_19400,N_18889,N_18723);
and U19401 (N_19401,N_18981,N_18574);
or U19402 (N_19402,N_18517,N_18910);
and U19403 (N_19403,N_18673,N_18650);
xnor U19404 (N_19404,N_18713,N_18576);
nor U19405 (N_19405,N_18774,N_18775);
nand U19406 (N_19406,N_18564,N_18766);
nand U19407 (N_19407,N_18700,N_18571);
xor U19408 (N_19408,N_18958,N_18506);
nor U19409 (N_19409,N_18526,N_18709);
nand U19410 (N_19410,N_18703,N_18832);
nor U19411 (N_19411,N_18854,N_18718);
xnor U19412 (N_19412,N_18670,N_18833);
or U19413 (N_19413,N_18519,N_18571);
xor U19414 (N_19414,N_18819,N_18979);
xnor U19415 (N_19415,N_18759,N_18826);
nand U19416 (N_19416,N_18986,N_18569);
nor U19417 (N_19417,N_18890,N_18587);
and U19418 (N_19418,N_18576,N_18908);
nand U19419 (N_19419,N_18864,N_18611);
and U19420 (N_19420,N_18664,N_18765);
nand U19421 (N_19421,N_18846,N_18706);
nand U19422 (N_19422,N_18755,N_18573);
and U19423 (N_19423,N_18801,N_18665);
or U19424 (N_19424,N_18620,N_18817);
nand U19425 (N_19425,N_18963,N_18765);
or U19426 (N_19426,N_18906,N_18787);
nand U19427 (N_19427,N_18648,N_18696);
and U19428 (N_19428,N_18528,N_18684);
nor U19429 (N_19429,N_18803,N_18841);
nor U19430 (N_19430,N_18880,N_18568);
nand U19431 (N_19431,N_18613,N_18766);
nand U19432 (N_19432,N_18693,N_18935);
or U19433 (N_19433,N_18766,N_18847);
and U19434 (N_19434,N_18515,N_18934);
nor U19435 (N_19435,N_18526,N_18985);
nand U19436 (N_19436,N_18856,N_18962);
xor U19437 (N_19437,N_18705,N_18724);
nor U19438 (N_19438,N_18720,N_18965);
nand U19439 (N_19439,N_18743,N_18854);
and U19440 (N_19440,N_18590,N_18798);
nor U19441 (N_19441,N_18697,N_18837);
nand U19442 (N_19442,N_18766,N_18929);
nor U19443 (N_19443,N_18620,N_18692);
nor U19444 (N_19444,N_18827,N_18673);
xor U19445 (N_19445,N_18833,N_18877);
or U19446 (N_19446,N_18643,N_18741);
xor U19447 (N_19447,N_18806,N_18785);
xor U19448 (N_19448,N_18642,N_18992);
and U19449 (N_19449,N_18582,N_18825);
and U19450 (N_19450,N_18523,N_18828);
or U19451 (N_19451,N_18556,N_18735);
nor U19452 (N_19452,N_18583,N_18646);
nor U19453 (N_19453,N_18868,N_18818);
and U19454 (N_19454,N_18881,N_18990);
nand U19455 (N_19455,N_18682,N_18702);
nand U19456 (N_19456,N_18668,N_18872);
nand U19457 (N_19457,N_18601,N_18862);
nor U19458 (N_19458,N_18762,N_18882);
nor U19459 (N_19459,N_18762,N_18637);
xor U19460 (N_19460,N_18630,N_18731);
xnor U19461 (N_19461,N_18710,N_18678);
and U19462 (N_19462,N_18730,N_18602);
nand U19463 (N_19463,N_18593,N_18998);
and U19464 (N_19464,N_18551,N_18516);
nor U19465 (N_19465,N_18834,N_18970);
nor U19466 (N_19466,N_18800,N_18552);
xnor U19467 (N_19467,N_18658,N_18869);
xnor U19468 (N_19468,N_18945,N_18577);
nand U19469 (N_19469,N_18851,N_18909);
or U19470 (N_19470,N_18780,N_18914);
or U19471 (N_19471,N_18904,N_18936);
nand U19472 (N_19472,N_18750,N_18637);
nand U19473 (N_19473,N_18734,N_18859);
nor U19474 (N_19474,N_18795,N_18523);
or U19475 (N_19475,N_18594,N_18585);
nor U19476 (N_19476,N_18671,N_18837);
nor U19477 (N_19477,N_18721,N_18518);
nor U19478 (N_19478,N_18526,N_18965);
xor U19479 (N_19479,N_18672,N_18700);
or U19480 (N_19480,N_18794,N_18526);
and U19481 (N_19481,N_18582,N_18685);
xor U19482 (N_19482,N_18831,N_18820);
xor U19483 (N_19483,N_18991,N_18864);
and U19484 (N_19484,N_18952,N_18727);
and U19485 (N_19485,N_18890,N_18956);
nor U19486 (N_19486,N_18764,N_18654);
or U19487 (N_19487,N_18953,N_18817);
xnor U19488 (N_19488,N_18551,N_18977);
nor U19489 (N_19489,N_18673,N_18924);
and U19490 (N_19490,N_18654,N_18539);
or U19491 (N_19491,N_18951,N_18756);
nor U19492 (N_19492,N_18863,N_18507);
and U19493 (N_19493,N_18723,N_18538);
or U19494 (N_19494,N_18519,N_18596);
xnor U19495 (N_19495,N_18630,N_18642);
or U19496 (N_19496,N_18947,N_18609);
nand U19497 (N_19497,N_18994,N_18560);
nand U19498 (N_19498,N_18739,N_18717);
or U19499 (N_19499,N_18984,N_18843);
nand U19500 (N_19500,N_19300,N_19319);
nand U19501 (N_19501,N_19374,N_19214);
nand U19502 (N_19502,N_19070,N_19478);
and U19503 (N_19503,N_19055,N_19174);
and U19504 (N_19504,N_19182,N_19457);
and U19505 (N_19505,N_19441,N_19459);
and U19506 (N_19506,N_19286,N_19344);
nand U19507 (N_19507,N_19033,N_19267);
nand U19508 (N_19508,N_19050,N_19423);
xnor U19509 (N_19509,N_19173,N_19129);
or U19510 (N_19510,N_19398,N_19155);
nand U19511 (N_19511,N_19453,N_19125);
nand U19512 (N_19512,N_19024,N_19222);
nand U19513 (N_19513,N_19490,N_19351);
xnor U19514 (N_19514,N_19434,N_19106);
or U19515 (N_19515,N_19137,N_19311);
or U19516 (N_19516,N_19204,N_19230);
nand U19517 (N_19517,N_19452,N_19361);
or U19518 (N_19518,N_19194,N_19268);
or U19519 (N_19519,N_19007,N_19199);
nor U19520 (N_19520,N_19027,N_19306);
and U19521 (N_19521,N_19305,N_19010);
xnor U19522 (N_19522,N_19333,N_19176);
xnor U19523 (N_19523,N_19405,N_19186);
or U19524 (N_19524,N_19196,N_19234);
nand U19525 (N_19525,N_19074,N_19087);
nand U19526 (N_19526,N_19396,N_19071);
nor U19527 (N_19527,N_19020,N_19118);
or U19528 (N_19528,N_19245,N_19003);
xnor U19529 (N_19529,N_19075,N_19185);
and U19530 (N_19530,N_19313,N_19322);
nor U19531 (N_19531,N_19330,N_19492);
or U19532 (N_19532,N_19251,N_19206);
xor U19533 (N_19533,N_19015,N_19067);
nor U19534 (N_19534,N_19164,N_19422);
and U19535 (N_19535,N_19140,N_19115);
and U19536 (N_19536,N_19336,N_19179);
and U19537 (N_19537,N_19201,N_19348);
or U19538 (N_19538,N_19209,N_19273);
nand U19539 (N_19539,N_19119,N_19253);
and U19540 (N_19540,N_19408,N_19240);
or U19541 (N_19541,N_19308,N_19445);
and U19542 (N_19542,N_19386,N_19416);
xnor U19543 (N_19543,N_19215,N_19021);
nand U19544 (N_19544,N_19407,N_19011);
nand U19545 (N_19545,N_19304,N_19170);
nand U19546 (N_19546,N_19426,N_19138);
nor U19547 (N_19547,N_19370,N_19032);
nor U19548 (N_19548,N_19147,N_19187);
xor U19549 (N_19549,N_19343,N_19143);
nand U19550 (N_19550,N_19346,N_19145);
nand U19551 (N_19551,N_19358,N_19292);
nor U19552 (N_19552,N_19456,N_19467);
and U19553 (N_19553,N_19122,N_19256);
nor U19554 (N_19554,N_19397,N_19250);
nor U19555 (N_19555,N_19377,N_19382);
xnor U19556 (N_19556,N_19475,N_19041);
nand U19557 (N_19557,N_19167,N_19284);
nand U19558 (N_19558,N_19447,N_19418);
xor U19559 (N_19559,N_19241,N_19270);
or U19560 (N_19560,N_19002,N_19178);
nand U19561 (N_19561,N_19139,N_19365);
or U19562 (N_19562,N_19112,N_19193);
nor U19563 (N_19563,N_19181,N_19442);
xnor U19564 (N_19564,N_19128,N_19328);
and U19565 (N_19565,N_19394,N_19068);
nand U19566 (N_19566,N_19092,N_19297);
xnor U19567 (N_19567,N_19157,N_19172);
nand U19568 (N_19568,N_19436,N_19325);
nand U19569 (N_19569,N_19184,N_19005);
nand U19570 (N_19570,N_19224,N_19360);
xnor U19571 (N_19571,N_19095,N_19229);
nor U19572 (N_19572,N_19168,N_19496);
and U19573 (N_19573,N_19142,N_19469);
or U19574 (N_19574,N_19472,N_19057);
and U19575 (N_19575,N_19347,N_19378);
xnor U19576 (N_19576,N_19123,N_19197);
nor U19577 (N_19577,N_19149,N_19329);
xor U19578 (N_19578,N_19152,N_19470);
nand U19579 (N_19579,N_19486,N_19159);
nand U19580 (N_19580,N_19237,N_19030);
nand U19581 (N_19581,N_19354,N_19047);
xnor U19582 (N_19582,N_19086,N_19189);
and U19583 (N_19583,N_19479,N_19078);
and U19584 (N_19584,N_19077,N_19252);
xor U19585 (N_19585,N_19403,N_19316);
nand U19586 (N_19586,N_19421,N_19044);
or U19587 (N_19587,N_19462,N_19497);
xnor U19588 (N_19588,N_19121,N_19244);
nand U19589 (N_19589,N_19312,N_19389);
and U19590 (N_19590,N_19108,N_19180);
nand U19591 (N_19591,N_19066,N_19272);
nor U19592 (N_19592,N_19171,N_19368);
and U19593 (N_19593,N_19216,N_19221);
nor U19594 (N_19594,N_19165,N_19104);
or U19595 (N_19595,N_19130,N_19051);
xnor U19596 (N_19596,N_19349,N_19009);
and U19597 (N_19597,N_19262,N_19260);
xor U19598 (N_19598,N_19376,N_19175);
nand U19599 (N_19599,N_19025,N_19296);
and U19600 (N_19600,N_19029,N_19105);
or U19601 (N_19601,N_19031,N_19056);
and U19602 (N_19602,N_19072,N_19279);
nor U19603 (N_19603,N_19126,N_19309);
and U19604 (N_19604,N_19191,N_19463);
or U19605 (N_19605,N_19283,N_19081);
and U19606 (N_19606,N_19052,N_19079);
xnor U19607 (N_19607,N_19466,N_19254);
nor U19608 (N_19608,N_19158,N_19385);
and U19609 (N_19609,N_19266,N_19135);
or U19610 (N_19610,N_19134,N_19243);
or U19611 (N_19611,N_19488,N_19271);
nand U19612 (N_19612,N_19303,N_19413);
xor U19613 (N_19613,N_19016,N_19146);
and U19614 (N_19614,N_19287,N_19393);
or U19615 (N_19615,N_19339,N_19188);
nand U19616 (N_19616,N_19217,N_19225);
or U19617 (N_19617,N_19446,N_19285);
xor U19618 (N_19618,N_19498,N_19064);
nand U19619 (N_19619,N_19359,N_19383);
nand U19620 (N_19620,N_19362,N_19246);
nor U19621 (N_19621,N_19449,N_19293);
nor U19622 (N_19622,N_19227,N_19116);
nor U19623 (N_19623,N_19063,N_19249);
nor U19624 (N_19624,N_19012,N_19166);
or U19625 (N_19625,N_19213,N_19094);
nor U19626 (N_19626,N_19248,N_19103);
or U19627 (N_19627,N_19468,N_19353);
and U19628 (N_19628,N_19282,N_19263);
xnor U19629 (N_19629,N_19485,N_19090);
nand U19630 (N_19630,N_19428,N_19192);
nor U19631 (N_19631,N_19277,N_19258);
nand U19632 (N_19632,N_19391,N_19257);
nand U19633 (N_19633,N_19307,N_19113);
xnor U19634 (N_19634,N_19473,N_19076);
nor U19635 (N_19635,N_19454,N_19111);
or U19636 (N_19636,N_19162,N_19489);
and U19637 (N_19637,N_19379,N_19402);
or U19638 (N_19638,N_19439,N_19372);
nor U19639 (N_19639,N_19034,N_19364);
nand U19640 (N_19640,N_19019,N_19054);
nor U19641 (N_19641,N_19480,N_19294);
nand U19642 (N_19642,N_19117,N_19499);
and U19643 (N_19643,N_19491,N_19059);
or U19644 (N_19644,N_19318,N_19226);
nor U19645 (N_19645,N_19210,N_19356);
xnor U19646 (N_19646,N_19085,N_19493);
xor U19647 (N_19647,N_19069,N_19028);
nor U19648 (N_19648,N_19202,N_19004);
and U19649 (N_19649,N_19101,N_19474);
and U19650 (N_19650,N_19443,N_19018);
and U19651 (N_19651,N_19124,N_19430);
xor U19652 (N_19652,N_19476,N_19384);
xor U19653 (N_19653,N_19367,N_19355);
xor U19654 (N_19654,N_19471,N_19281);
nor U19655 (N_19655,N_19429,N_19151);
nor U19656 (N_19656,N_19437,N_19371);
and U19657 (N_19657,N_19156,N_19006);
xor U19658 (N_19658,N_19100,N_19022);
nand U19659 (N_19659,N_19427,N_19302);
nor U19660 (N_19660,N_19131,N_19096);
nor U19661 (N_19661,N_19259,N_19388);
nand U19662 (N_19662,N_19036,N_19017);
and U19663 (N_19663,N_19269,N_19205);
or U19664 (N_19664,N_19410,N_19035);
or U19665 (N_19665,N_19107,N_19045);
or U19666 (N_19666,N_19211,N_19363);
and U19667 (N_19667,N_19053,N_19220);
xnor U19668 (N_19668,N_19265,N_19102);
nor U19669 (N_19669,N_19342,N_19482);
or U19670 (N_19670,N_19484,N_19048);
and U19671 (N_19671,N_19247,N_19208);
or U19672 (N_19672,N_19380,N_19477);
nand U19673 (N_19673,N_19242,N_19337);
xor U19674 (N_19674,N_19401,N_19190);
xnor U19675 (N_19675,N_19327,N_19431);
nor U19676 (N_19676,N_19161,N_19089);
xnor U19677 (N_19677,N_19417,N_19392);
and U19678 (N_19678,N_19177,N_19037);
xor U19679 (N_19679,N_19001,N_19425);
xor U19680 (N_19680,N_19233,N_19212);
nor U19681 (N_19681,N_19198,N_19148);
nand U19682 (N_19682,N_19373,N_19219);
and U19683 (N_19683,N_19314,N_19414);
and U19684 (N_19684,N_19494,N_19203);
or U19685 (N_19685,N_19400,N_19350);
and U19686 (N_19686,N_19049,N_19331);
and U19687 (N_19687,N_19420,N_19099);
nand U19688 (N_19688,N_19338,N_19133);
nor U19689 (N_19689,N_19183,N_19326);
or U19690 (N_19690,N_19357,N_19419);
xor U19691 (N_19691,N_19160,N_19120);
xor U19692 (N_19692,N_19409,N_19404);
or U19693 (N_19693,N_19461,N_19065);
nand U19694 (N_19694,N_19073,N_19411);
or U19695 (N_19695,N_19043,N_19375);
and U19696 (N_19696,N_19039,N_19455);
xnor U19697 (N_19697,N_19058,N_19433);
nand U19698 (N_19698,N_19366,N_19275);
nor U19699 (N_19699,N_19369,N_19238);
nand U19700 (N_19700,N_19114,N_19207);
nor U19701 (N_19701,N_19255,N_19341);
nand U19702 (N_19702,N_19448,N_19390);
nand U19703 (N_19703,N_19239,N_19291);
nand U19704 (N_19704,N_19406,N_19046);
and U19705 (N_19705,N_19141,N_19062);
xor U19706 (N_19706,N_19465,N_19387);
nand U19707 (N_19707,N_19093,N_19060);
or U19708 (N_19708,N_19195,N_19150);
xor U19709 (N_19709,N_19109,N_19345);
and U19710 (N_19710,N_19432,N_19424);
xor U19711 (N_19711,N_19091,N_19228);
nor U19712 (N_19712,N_19014,N_19098);
or U19713 (N_19713,N_19231,N_19320);
nand U19714 (N_19714,N_19236,N_19000);
nand U19715 (N_19715,N_19321,N_19481);
nor U19716 (N_19716,N_19169,N_19335);
and U19717 (N_19717,N_19352,N_19136);
and U19718 (N_19718,N_19084,N_19082);
nand U19719 (N_19719,N_19274,N_19288);
nand U19720 (N_19720,N_19144,N_19132);
xor U19721 (N_19721,N_19080,N_19399);
nor U19722 (N_19722,N_19412,N_19460);
xnor U19723 (N_19723,N_19495,N_19276);
nor U19724 (N_19724,N_19223,N_19110);
nand U19725 (N_19725,N_19088,N_19315);
nor U19726 (N_19726,N_19038,N_19264);
xnor U19727 (N_19727,N_19163,N_19487);
or U19728 (N_19728,N_19040,N_19381);
xnor U19729 (N_19729,N_19310,N_19042);
nor U19730 (N_19730,N_19323,N_19298);
nor U19731 (N_19731,N_19061,N_19289);
xor U19732 (N_19732,N_19097,N_19332);
and U19733 (N_19733,N_19395,N_19295);
nor U19734 (N_19734,N_19261,N_19013);
nand U19735 (N_19735,N_19026,N_19444);
and U19736 (N_19736,N_19317,N_19458);
and U19737 (N_19737,N_19438,N_19324);
or U19738 (N_19738,N_19464,N_19278);
and U19739 (N_19739,N_19218,N_19153);
and U19740 (N_19740,N_19299,N_19200);
or U19741 (N_19741,N_19008,N_19483);
xor U19742 (N_19742,N_19154,N_19290);
nor U19743 (N_19743,N_19440,N_19023);
xor U19744 (N_19744,N_19280,N_19127);
xor U19745 (N_19745,N_19083,N_19415);
xnor U19746 (N_19746,N_19435,N_19232);
or U19747 (N_19747,N_19340,N_19235);
nand U19748 (N_19748,N_19301,N_19334);
nor U19749 (N_19749,N_19451,N_19450);
nand U19750 (N_19750,N_19359,N_19355);
nor U19751 (N_19751,N_19076,N_19075);
and U19752 (N_19752,N_19447,N_19483);
nor U19753 (N_19753,N_19298,N_19259);
nand U19754 (N_19754,N_19495,N_19246);
or U19755 (N_19755,N_19234,N_19399);
and U19756 (N_19756,N_19233,N_19113);
nand U19757 (N_19757,N_19113,N_19104);
or U19758 (N_19758,N_19404,N_19437);
xnor U19759 (N_19759,N_19348,N_19314);
and U19760 (N_19760,N_19121,N_19260);
nor U19761 (N_19761,N_19154,N_19075);
nand U19762 (N_19762,N_19128,N_19450);
nor U19763 (N_19763,N_19354,N_19262);
nor U19764 (N_19764,N_19165,N_19428);
nand U19765 (N_19765,N_19444,N_19370);
xor U19766 (N_19766,N_19179,N_19140);
nand U19767 (N_19767,N_19333,N_19377);
xor U19768 (N_19768,N_19348,N_19302);
nor U19769 (N_19769,N_19404,N_19483);
nor U19770 (N_19770,N_19421,N_19484);
xor U19771 (N_19771,N_19449,N_19200);
and U19772 (N_19772,N_19367,N_19472);
and U19773 (N_19773,N_19233,N_19063);
or U19774 (N_19774,N_19065,N_19353);
or U19775 (N_19775,N_19495,N_19046);
xor U19776 (N_19776,N_19037,N_19487);
nor U19777 (N_19777,N_19356,N_19080);
or U19778 (N_19778,N_19292,N_19193);
xor U19779 (N_19779,N_19274,N_19244);
nor U19780 (N_19780,N_19484,N_19197);
nand U19781 (N_19781,N_19394,N_19207);
nand U19782 (N_19782,N_19226,N_19494);
xor U19783 (N_19783,N_19226,N_19243);
nand U19784 (N_19784,N_19378,N_19337);
nor U19785 (N_19785,N_19376,N_19103);
or U19786 (N_19786,N_19230,N_19224);
and U19787 (N_19787,N_19135,N_19468);
nor U19788 (N_19788,N_19296,N_19099);
nor U19789 (N_19789,N_19493,N_19193);
nor U19790 (N_19790,N_19010,N_19443);
nor U19791 (N_19791,N_19326,N_19427);
xnor U19792 (N_19792,N_19070,N_19228);
xnor U19793 (N_19793,N_19215,N_19372);
or U19794 (N_19794,N_19445,N_19404);
nand U19795 (N_19795,N_19472,N_19442);
or U19796 (N_19796,N_19127,N_19490);
nand U19797 (N_19797,N_19400,N_19055);
and U19798 (N_19798,N_19160,N_19397);
or U19799 (N_19799,N_19219,N_19185);
and U19800 (N_19800,N_19008,N_19045);
xor U19801 (N_19801,N_19012,N_19349);
and U19802 (N_19802,N_19077,N_19465);
or U19803 (N_19803,N_19121,N_19306);
nand U19804 (N_19804,N_19214,N_19225);
or U19805 (N_19805,N_19134,N_19395);
xor U19806 (N_19806,N_19060,N_19458);
or U19807 (N_19807,N_19083,N_19377);
nand U19808 (N_19808,N_19187,N_19030);
nand U19809 (N_19809,N_19114,N_19272);
xor U19810 (N_19810,N_19291,N_19461);
nor U19811 (N_19811,N_19247,N_19060);
xor U19812 (N_19812,N_19462,N_19127);
nor U19813 (N_19813,N_19089,N_19241);
nor U19814 (N_19814,N_19376,N_19495);
and U19815 (N_19815,N_19041,N_19292);
nor U19816 (N_19816,N_19130,N_19356);
xnor U19817 (N_19817,N_19121,N_19219);
nand U19818 (N_19818,N_19141,N_19046);
xnor U19819 (N_19819,N_19085,N_19162);
nand U19820 (N_19820,N_19016,N_19182);
and U19821 (N_19821,N_19112,N_19191);
or U19822 (N_19822,N_19075,N_19393);
nor U19823 (N_19823,N_19095,N_19048);
xnor U19824 (N_19824,N_19042,N_19498);
xor U19825 (N_19825,N_19495,N_19052);
and U19826 (N_19826,N_19052,N_19347);
xnor U19827 (N_19827,N_19069,N_19217);
xor U19828 (N_19828,N_19071,N_19127);
and U19829 (N_19829,N_19008,N_19202);
and U19830 (N_19830,N_19180,N_19303);
or U19831 (N_19831,N_19332,N_19169);
nor U19832 (N_19832,N_19060,N_19119);
nor U19833 (N_19833,N_19174,N_19208);
and U19834 (N_19834,N_19075,N_19173);
xor U19835 (N_19835,N_19292,N_19277);
nand U19836 (N_19836,N_19111,N_19347);
or U19837 (N_19837,N_19403,N_19276);
xnor U19838 (N_19838,N_19181,N_19387);
nor U19839 (N_19839,N_19457,N_19271);
or U19840 (N_19840,N_19018,N_19340);
nor U19841 (N_19841,N_19081,N_19129);
xnor U19842 (N_19842,N_19495,N_19273);
or U19843 (N_19843,N_19201,N_19320);
xnor U19844 (N_19844,N_19178,N_19087);
nand U19845 (N_19845,N_19391,N_19055);
or U19846 (N_19846,N_19057,N_19291);
xor U19847 (N_19847,N_19165,N_19197);
nand U19848 (N_19848,N_19053,N_19106);
xor U19849 (N_19849,N_19306,N_19026);
and U19850 (N_19850,N_19412,N_19178);
nand U19851 (N_19851,N_19360,N_19122);
xor U19852 (N_19852,N_19294,N_19489);
or U19853 (N_19853,N_19175,N_19331);
xor U19854 (N_19854,N_19177,N_19333);
xor U19855 (N_19855,N_19159,N_19422);
nand U19856 (N_19856,N_19140,N_19452);
nor U19857 (N_19857,N_19438,N_19032);
and U19858 (N_19858,N_19430,N_19458);
and U19859 (N_19859,N_19328,N_19387);
and U19860 (N_19860,N_19115,N_19003);
nand U19861 (N_19861,N_19098,N_19158);
xor U19862 (N_19862,N_19427,N_19308);
xnor U19863 (N_19863,N_19032,N_19045);
xnor U19864 (N_19864,N_19412,N_19055);
xor U19865 (N_19865,N_19024,N_19472);
and U19866 (N_19866,N_19300,N_19268);
nand U19867 (N_19867,N_19061,N_19426);
or U19868 (N_19868,N_19040,N_19430);
xnor U19869 (N_19869,N_19392,N_19119);
or U19870 (N_19870,N_19008,N_19495);
xor U19871 (N_19871,N_19053,N_19041);
or U19872 (N_19872,N_19088,N_19456);
xor U19873 (N_19873,N_19455,N_19005);
or U19874 (N_19874,N_19211,N_19342);
and U19875 (N_19875,N_19016,N_19488);
or U19876 (N_19876,N_19111,N_19451);
and U19877 (N_19877,N_19375,N_19385);
xor U19878 (N_19878,N_19404,N_19238);
xor U19879 (N_19879,N_19333,N_19123);
xnor U19880 (N_19880,N_19075,N_19339);
or U19881 (N_19881,N_19278,N_19405);
or U19882 (N_19882,N_19045,N_19199);
or U19883 (N_19883,N_19095,N_19408);
nand U19884 (N_19884,N_19085,N_19223);
and U19885 (N_19885,N_19205,N_19401);
xnor U19886 (N_19886,N_19173,N_19498);
nand U19887 (N_19887,N_19444,N_19375);
xor U19888 (N_19888,N_19140,N_19314);
or U19889 (N_19889,N_19187,N_19232);
xor U19890 (N_19890,N_19119,N_19455);
nand U19891 (N_19891,N_19229,N_19210);
nand U19892 (N_19892,N_19349,N_19243);
or U19893 (N_19893,N_19367,N_19174);
nand U19894 (N_19894,N_19292,N_19407);
nand U19895 (N_19895,N_19025,N_19357);
xor U19896 (N_19896,N_19151,N_19478);
or U19897 (N_19897,N_19125,N_19156);
nand U19898 (N_19898,N_19311,N_19496);
xnor U19899 (N_19899,N_19223,N_19445);
nand U19900 (N_19900,N_19365,N_19368);
nand U19901 (N_19901,N_19228,N_19324);
or U19902 (N_19902,N_19385,N_19088);
nand U19903 (N_19903,N_19183,N_19382);
nand U19904 (N_19904,N_19407,N_19365);
and U19905 (N_19905,N_19342,N_19329);
nand U19906 (N_19906,N_19279,N_19447);
nor U19907 (N_19907,N_19022,N_19264);
and U19908 (N_19908,N_19207,N_19402);
and U19909 (N_19909,N_19195,N_19453);
nand U19910 (N_19910,N_19003,N_19432);
nand U19911 (N_19911,N_19214,N_19159);
and U19912 (N_19912,N_19078,N_19286);
and U19913 (N_19913,N_19287,N_19256);
or U19914 (N_19914,N_19258,N_19225);
xnor U19915 (N_19915,N_19149,N_19385);
nand U19916 (N_19916,N_19426,N_19064);
or U19917 (N_19917,N_19210,N_19476);
and U19918 (N_19918,N_19332,N_19437);
xor U19919 (N_19919,N_19298,N_19029);
and U19920 (N_19920,N_19113,N_19251);
or U19921 (N_19921,N_19392,N_19260);
xnor U19922 (N_19922,N_19478,N_19096);
xnor U19923 (N_19923,N_19021,N_19009);
xor U19924 (N_19924,N_19278,N_19472);
and U19925 (N_19925,N_19212,N_19332);
xnor U19926 (N_19926,N_19281,N_19340);
nor U19927 (N_19927,N_19362,N_19022);
and U19928 (N_19928,N_19214,N_19009);
and U19929 (N_19929,N_19363,N_19136);
nor U19930 (N_19930,N_19426,N_19495);
nor U19931 (N_19931,N_19119,N_19412);
and U19932 (N_19932,N_19444,N_19331);
nor U19933 (N_19933,N_19360,N_19103);
or U19934 (N_19934,N_19275,N_19340);
or U19935 (N_19935,N_19365,N_19025);
nand U19936 (N_19936,N_19225,N_19265);
xnor U19937 (N_19937,N_19301,N_19230);
nand U19938 (N_19938,N_19194,N_19409);
xnor U19939 (N_19939,N_19052,N_19360);
nor U19940 (N_19940,N_19213,N_19036);
xor U19941 (N_19941,N_19445,N_19415);
and U19942 (N_19942,N_19465,N_19378);
nand U19943 (N_19943,N_19439,N_19360);
and U19944 (N_19944,N_19311,N_19204);
and U19945 (N_19945,N_19360,N_19426);
xnor U19946 (N_19946,N_19029,N_19374);
and U19947 (N_19947,N_19254,N_19411);
nor U19948 (N_19948,N_19032,N_19315);
and U19949 (N_19949,N_19147,N_19344);
nor U19950 (N_19950,N_19453,N_19055);
nand U19951 (N_19951,N_19287,N_19258);
or U19952 (N_19952,N_19094,N_19479);
nor U19953 (N_19953,N_19036,N_19232);
nor U19954 (N_19954,N_19177,N_19456);
nand U19955 (N_19955,N_19370,N_19087);
or U19956 (N_19956,N_19225,N_19431);
nand U19957 (N_19957,N_19272,N_19139);
nand U19958 (N_19958,N_19195,N_19421);
nor U19959 (N_19959,N_19211,N_19477);
nor U19960 (N_19960,N_19257,N_19167);
nor U19961 (N_19961,N_19294,N_19498);
nor U19962 (N_19962,N_19450,N_19416);
and U19963 (N_19963,N_19455,N_19273);
xor U19964 (N_19964,N_19294,N_19370);
and U19965 (N_19965,N_19422,N_19332);
and U19966 (N_19966,N_19462,N_19224);
nand U19967 (N_19967,N_19194,N_19384);
nor U19968 (N_19968,N_19414,N_19323);
or U19969 (N_19969,N_19344,N_19413);
xor U19970 (N_19970,N_19004,N_19111);
xor U19971 (N_19971,N_19220,N_19437);
nor U19972 (N_19972,N_19392,N_19421);
xor U19973 (N_19973,N_19421,N_19229);
or U19974 (N_19974,N_19426,N_19353);
or U19975 (N_19975,N_19347,N_19475);
xnor U19976 (N_19976,N_19132,N_19320);
and U19977 (N_19977,N_19226,N_19351);
nor U19978 (N_19978,N_19288,N_19387);
nor U19979 (N_19979,N_19071,N_19103);
or U19980 (N_19980,N_19221,N_19321);
nand U19981 (N_19981,N_19199,N_19395);
nor U19982 (N_19982,N_19465,N_19433);
xor U19983 (N_19983,N_19221,N_19123);
nand U19984 (N_19984,N_19285,N_19346);
or U19985 (N_19985,N_19139,N_19170);
nand U19986 (N_19986,N_19443,N_19310);
nor U19987 (N_19987,N_19114,N_19425);
and U19988 (N_19988,N_19368,N_19022);
nand U19989 (N_19989,N_19112,N_19158);
nand U19990 (N_19990,N_19301,N_19489);
xnor U19991 (N_19991,N_19044,N_19453);
xor U19992 (N_19992,N_19181,N_19382);
nor U19993 (N_19993,N_19483,N_19449);
nand U19994 (N_19994,N_19269,N_19318);
and U19995 (N_19995,N_19095,N_19278);
or U19996 (N_19996,N_19444,N_19256);
nor U19997 (N_19997,N_19296,N_19379);
nand U19998 (N_19998,N_19299,N_19259);
or U19999 (N_19999,N_19033,N_19430);
or U20000 (N_20000,N_19740,N_19664);
nand U20001 (N_20001,N_19829,N_19515);
or U20002 (N_20002,N_19728,N_19623);
nor U20003 (N_20003,N_19517,N_19949);
nor U20004 (N_20004,N_19874,N_19941);
xor U20005 (N_20005,N_19582,N_19886);
or U20006 (N_20006,N_19511,N_19882);
nor U20007 (N_20007,N_19945,N_19572);
nor U20008 (N_20008,N_19574,N_19961);
nand U20009 (N_20009,N_19520,N_19998);
and U20010 (N_20010,N_19779,N_19746);
or U20011 (N_20011,N_19772,N_19605);
xor U20012 (N_20012,N_19830,N_19683);
and U20013 (N_20013,N_19692,N_19719);
nor U20014 (N_20014,N_19584,N_19690);
and U20015 (N_20015,N_19516,N_19781);
and U20016 (N_20016,N_19512,N_19879);
xnor U20017 (N_20017,N_19702,N_19983);
or U20018 (N_20018,N_19845,N_19654);
xor U20019 (N_20019,N_19839,N_19617);
or U20020 (N_20020,N_19645,N_19730);
nor U20021 (N_20021,N_19782,N_19864);
nand U20022 (N_20022,N_19710,N_19614);
nor U20023 (N_20023,N_19704,N_19932);
xor U20024 (N_20024,N_19519,N_19817);
or U20025 (N_20025,N_19569,N_19532);
xor U20026 (N_20026,N_19883,N_19641);
nor U20027 (N_20027,N_19981,N_19666);
nor U20028 (N_20028,N_19863,N_19648);
and U20029 (N_20029,N_19554,N_19593);
nand U20030 (N_20030,N_19884,N_19831);
or U20031 (N_20031,N_19788,N_19608);
nand U20032 (N_20032,N_19852,N_19906);
nor U20033 (N_20033,N_19741,N_19607);
xnor U20034 (N_20034,N_19916,N_19501);
nor U20035 (N_20035,N_19531,N_19634);
nor U20036 (N_20036,N_19663,N_19771);
or U20037 (N_20037,N_19815,N_19962);
nor U20038 (N_20038,N_19715,N_19756);
and U20039 (N_20039,N_19753,N_19801);
and U20040 (N_20040,N_19660,N_19861);
and U20041 (N_20041,N_19679,N_19651);
and U20042 (N_20042,N_19652,N_19576);
or U20043 (N_20043,N_19892,N_19625);
or U20044 (N_20044,N_19917,N_19828);
nand U20045 (N_20045,N_19626,N_19503);
nand U20046 (N_20046,N_19967,N_19673);
nand U20047 (N_20047,N_19972,N_19896);
nor U20048 (N_20048,N_19547,N_19948);
and U20049 (N_20049,N_19853,N_19703);
nand U20050 (N_20050,N_19534,N_19676);
nor U20051 (N_20051,N_19693,N_19527);
or U20052 (N_20052,N_19894,N_19834);
nand U20053 (N_20053,N_19758,N_19787);
and U20054 (N_20054,N_19836,N_19566);
or U20055 (N_20055,N_19548,N_19933);
and U20056 (N_20056,N_19604,N_19632);
or U20057 (N_20057,N_19696,N_19729);
or U20058 (N_20058,N_19814,N_19778);
xnor U20059 (N_20059,N_19550,N_19558);
xor U20060 (N_20060,N_19525,N_19562);
nand U20061 (N_20061,N_19594,N_19549);
or U20062 (N_20062,N_19857,N_19988);
nand U20063 (N_20063,N_19543,N_19585);
xnor U20064 (N_20064,N_19678,N_19529);
and U20065 (N_20065,N_19505,N_19975);
xor U20066 (N_20066,N_19766,N_19510);
or U20067 (N_20067,N_19923,N_19726);
and U20068 (N_20068,N_19871,N_19596);
xnor U20069 (N_20069,N_19720,N_19925);
and U20070 (N_20070,N_19599,N_19540);
xor U20071 (N_20071,N_19905,N_19682);
nor U20072 (N_20072,N_19601,N_19738);
nor U20073 (N_20073,N_19609,N_19731);
nand U20074 (N_20074,N_19705,N_19658);
or U20075 (N_20075,N_19752,N_19826);
xnor U20076 (N_20076,N_19813,N_19717);
nor U20077 (N_20077,N_19976,N_19669);
and U20078 (N_20078,N_19956,N_19765);
nand U20079 (N_20079,N_19947,N_19553);
nand U20080 (N_20080,N_19966,N_19754);
or U20081 (N_20081,N_19768,N_19557);
nor U20082 (N_20082,N_19848,N_19761);
and U20083 (N_20083,N_19806,N_19914);
or U20084 (N_20084,N_19960,N_19524);
or U20085 (N_20085,N_19721,N_19943);
or U20086 (N_20086,N_19670,N_19910);
nand U20087 (N_20087,N_19640,N_19544);
xor U20088 (N_20088,N_19637,N_19902);
nor U20089 (N_20089,N_19631,N_19866);
nand U20090 (N_20090,N_19784,N_19895);
xnor U20091 (N_20091,N_19795,N_19659);
and U20092 (N_20092,N_19823,N_19946);
nor U20093 (N_20093,N_19624,N_19958);
nor U20094 (N_20094,N_19964,N_19698);
nor U20095 (N_20095,N_19764,N_19940);
or U20096 (N_20096,N_19591,N_19994);
or U20097 (N_20097,N_19661,N_19850);
nand U20098 (N_20098,N_19577,N_19602);
nor U20099 (N_20099,N_19565,N_19799);
or U20100 (N_20100,N_19775,N_19837);
or U20101 (N_20101,N_19650,N_19952);
nor U20102 (N_20102,N_19615,N_19633);
and U20103 (N_20103,N_19820,N_19950);
and U20104 (N_20104,N_19545,N_19714);
nand U20105 (N_20105,N_19748,N_19708);
xnor U20106 (N_20106,N_19867,N_19571);
nand U20107 (N_20107,N_19610,N_19984);
xnor U20108 (N_20108,N_19595,N_19928);
xnor U20109 (N_20109,N_19570,N_19987);
and U20110 (N_20110,N_19969,N_19802);
or U20111 (N_20111,N_19957,N_19776);
nor U20112 (N_20112,N_19927,N_19955);
nor U20113 (N_20113,N_19913,N_19757);
nand U20114 (N_20114,N_19800,N_19774);
and U20115 (N_20115,N_19749,N_19942);
xor U20116 (N_20116,N_19797,N_19970);
or U20117 (N_20117,N_19711,N_19810);
nor U20118 (N_20118,N_19860,N_19931);
nor U20119 (N_20119,N_19694,N_19622);
nor U20120 (N_20120,N_19734,N_19851);
or U20121 (N_20121,N_19722,N_19526);
nor U20122 (N_20122,N_19671,N_19662);
nor U20123 (N_20123,N_19838,N_19777);
xnor U20124 (N_20124,N_19513,N_19522);
xnor U20125 (N_20125,N_19996,N_19769);
and U20126 (N_20126,N_19747,N_19959);
and U20127 (N_20127,N_19796,N_19603);
nand U20128 (N_20128,N_19875,N_19900);
xor U20129 (N_20129,N_19793,N_19934);
xor U20130 (N_20130,N_19903,N_19870);
nor U20131 (N_20131,N_19811,N_19999);
or U20132 (N_20132,N_19809,N_19885);
nor U20133 (N_20133,N_19653,N_19681);
nand U20134 (N_20134,N_19689,N_19995);
and U20135 (N_20135,N_19856,N_19898);
or U20136 (N_20136,N_19621,N_19805);
nor U20137 (N_20137,N_19613,N_19798);
and U20138 (N_20138,N_19588,N_19509);
nor U20139 (N_20139,N_19611,N_19675);
nor U20140 (N_20140,N_19835,N_19672);
or U20141 (N_20141,N_19786,N_19979);
and U20142 (N_20142,N_19759,N_19854);
and U20143 (N_20143,N_19745,N_19973);
or U20144 (N_20144,N_19612,N_19921);
or U20145 (N_20145,N_19518,N_19713);
and U20146 (N_20146,N_19929,N_19537);
nand U20147 (N_20147,N_19869,N_19818);
nand U20148 (N_20148,N_19918,N_19767);
nand U20149 (N_20149,N_19579,N_19887);
nor U20150 (N_20150,N_19880,N_19862);
nor U20151 (N_20151,N_19655,N_19739);
nand U20152 (N_20152,N_19706,N_19827);
xnor U20153 (N_20153,N_19858,N_19638);
and U20154 (N_20154,N_19922,N_19523);
and U20155 (N_20155,N_19944,N_19600);
or U20156 (N_20156,N_19978,N_19762);
and U20157 (N_20157,N_19794,N_19742);
nor U20158 (N_20158,N_19735,N_19709);
and U20159 (N_20159,N_19844,N_19954);
or U20160 (N_20160,N_19635,N_19897);
and U20161 (N_20161,N_19568,N_19724);
nand U20162 (N_20162,N_19628,N_19926);
and U20163 (N_20163,N_19812,N_19687);
nor U20164 (N_20164,N_19750,N_19643);
xor U20165 (N_20165,N_19907,N_19546);
nand U20166 (N_20166,N_19790,N_19963);
and U20167 (N_20167,N_19751,N_19500);
and U20168 (N_20168,N_19737,N_19953);
or U20169 (N_20169,N_19564,N_19697);
xor U20170 (N_20170,N_19990,N_19620);
and U20171 (N_20171,N_19807,N_19684);
nand U20172 (N_20172,N_19590,N_19938);
nand U20173 (N_20173,N_19804,N_19618);
or U20174 (N_20174,N_19533,N_19974);
nor U20175 (N_20175,N_19783,N_19674);
xnor U20176 (N_20176,N_19559,N_19589);
or U20177 (N_20177,N_19736,N_19808);
nor U20178 (N_20178,N_19824,N_19733);
and U20179 (N_20179,N_19560,N_19868);
or U20180 (N_20180,N_19699,N_19685);
nand U20181 (N_20181,N_19521,N_19592);
nand U20182 (N_20182,N_19865,N_19563);
and U20183 (N_20183,N_19642,N_19502);
nand U20184 (N_20184,N_19580,N_19597);
nor U20185 (N_20185,N_19567,N_19891);
or U20186 (N_20186,N_19630,N_19819);
nand U20187 (N_20187,N_19575,N_19873);
and U20188 (N_20188,N_19968,N_19578);
and U20189 (N_20189,N_19639,N_19665);
and U20190 (N_20190,N_19732,N_19555);
nor U20191 (N_20191,N_19712,N_19668);
nand U20192 (N_20192,N_19707,N_19770);
xnor U20193 (N_20193,N_19583,N_19951);
xnor U20194 (N_20194,N_19514,N_19760);
xor U20195 (N_20195,N_19780,N_19989);
xor U20196 (N_20196,N_19629,N_19606);
or U20197 (N_20197,N_19821,N_19552);
or U20198 (N_20198,N_19843,N_19657);
nor U20199 (N_20199,N_19727,N_19542);
nand U20200 (N_20200,N_19695,N_19688);
xnor U20201 (N_20201,N_19680,N_19536);
nand U20202 (N_20202,N_19816,N_19911);
or U20203 (N_20203,N_19993,N_19935);
or U20204 (N_20204,N_19877,N_19744);
nor U20205 (N_20205,N_19587,N_19893);
and U20206 (N_20206,N_19647,N_19846);
xnor U20207 (N_20207,N_19723,N_19644);
and U20208 (N_20208,N_19677,N_19985);
nor U20209 (N_20209,N_19997,N_19598);
and U20210 (N_20210,N_19888,N_19833);
xor U20211 (N_20211,N_19636,N_19971);
xnor U20212 (N_20212,N_19878,N_19840);
and U20213 (N_20213,N_19701,N_19841);
xor U20214 (N_20214,N_19507,N_19901);
nand U20215 (N_20215,N_19936,N_19743);
nand U20216 (N_20216,N_19538,N_19686);
nor U20217 (N_20217,N_19939,N_19785);
and U20218 (N_20218,N_19822,N_19791);
nand U20219 (N_20219,N_19876,N_19667);
xor U20220 (N_20220,N_19909,N_19847);
nand U20221 (N_20221,N_19508,N_19528);
or U20222 (N_20222,N_19915,N_19904);
and U20223 (N_20223,N_19937,N_19977);
or U20224 (N_20224,N_19700,N_19755);
xnor U20225 (N_20225,N_19619,N_19991);
nand U20226 (N_20226,N_19859,N_19919);
nand U20227 (N_20227,N_19889,N_19616);
nand U20228 (N_20228,N_19825,N_19773);
or U20229 (N_20229,N_19872,N_19586);
xnor U20230 (N_20230,N_19986,N_19530);
nor U20231 (N_20231,N_19541,N_19982);
xnor U20232 (N_20232,N_19789,N_19539);
xor U20233 (N_20233,N_19855,N_19649);
and U20234 (N_20234,N_19899,N_19627);
xor U20235 (N_20235,N_19930,N_19581);
nand U20236 (N_20236,N_19504,N_19832);
nand U20237 (N_20237,N_19535,N_19920);
and U20238 (N_20238,N_19792,N_19561);
xnor U20239 (N_20239,N_19718,N_19763);
or U20240 (N_20240,N_19890,N_19924);
nand U20241 (N_20241,N_19716,N_19725);
and U20242 (N_20242,N_19556,N_19656);
xnor U20243 (N_20243,N_19849,N_19646);
and U20244 (N_20244,N_19908,N_19803);
xor U20245 (N_20245,N_19842,N_19992);
nand U20246 (N_20246,N_19980,N_19506);
nand U20247 (N_20247,N_19691,N_19912);
xnor U20248 (N_20248,N_19551,N_19573);
and U20249 (N_20249,N_19881,N_19965);
nor U20250 (N_20250,N_19531,N_19905);
nor U20251 (N_20251,N_19924,N_19806);
or U20252 (N_20252,N_19561,N_19512);
nand U20253 (N_20253,N_19980,N_19721);
nor U20254 (N_20254,N_19835,N_19734);
or U20255 (N_20255,N_19703,N_19888);
xor U20256 (N_20256,N_19727,N_19520);
nor U20257 (N_20257,N_19925,N_19583);
and U20258 (N_20258,N_19919,N_19614);
nand U20259 (N_20259,N_19960,N_19679);
nand U20260 (N_20260,N_19500,N_19833);
and U20261 (N_20261,N_19830,N_19724);
xor U20262 (N_20262,N_19957,N_19744);
nor U20263 (N_20263,N_19612,N_19805);
or U20264 (N_20264,N_19528,N_19974);
nor U20265 (N_20265,N_19899,N_19757);
nor U20266 (N_20266,N_19749,N_19562);
nand U20267 (N_20267,N_19509,N_19540);
nand U20268 (N_20268,N_19589,N_19615);
nor U20269 (N_20269,N_19568,N_19617);
nand U20270 (N_20270,N_19883,N_19996);
xor U20271 (N_20271,N_19689,N_19934);
and U20272 (N_20272,N_19992,N_19655);
and U20273 (N_20273,N_19585,N_19824);
xnor U20274 (N_20274,N_19518,N_19818);
and U20275 (N_20275,N_19772,N_19991);
or U20276 (N_20276,N_19826,N_19510);
and U20277 (N_20277,N_19715,N_19898);
nand U20278 (N_20278,N_19551,N_19591);
xnor U20279 (N_20279,N_19519,N_19905);
xnor U20280 (N_20280,N_19834,N_19809);
nor U20281 (N_20281,N_19873,N_19836);
and U20282 (N_20282,N_19743,N_19726);
xor U20283 (N_20283,N_19522,N_19754);
and U20284 (N_20284,N_19583,N_19868);
and U20285 (N_20285,N_19946,N_19991);
nor U20286 (N_20286,N_19929,N_19705);
and U20287 (N_20287,N_19973,N_19701);
or U20288 (N_20288,N_19997,N_19582);
nor U20289 (N_20289,N_19732,N_19872);
and U20290 (N_20290,N_19964,N_19941);
nand U20291 (N_20291,N_19931,N_19974);
or U20292 (N_20292,N_19978,N_19646);
or U20293 (N_20293,N_19919,N_19898);
nor U20294 (N_20294,N_19722,N_19742);
xor U20295 (N_20295,N_19506,N_19901);
or U20296 (N_20296,N_19888,N_19713);
and U20297 (N_20297,N_19648,N_19526);
nand U20298 (N_20298,N_19716,N_19777);
xnor U20299 (N_20299,N_19906,N_19945);
nor U20300 (N_20300,N_19727,N_19975);
and U20301 (N_20301,N_19852,N_19772);
and U20302 (N_20302,N_19701,N_19501);
nand U20303 (N_20303,N_19612,N_19958);
nor U20304 (N_20304,N_19656,N_19622);
or U20305 (N_20305,N_19631,N_19966);
xor U20306 (N_20306,N_19726,N_19599);
nand U20307 (N_20307,N_19750,N_19716);
and U20308 (N_20308,N_19522,N_19701);
xor U20309 (N_20309,N_19980,N_19863);
nor U20310 (N_20310,N_19635,N_19554);
nand U20311 (N_20311,N_19538,N_19600);
xor U20312 (N_20312,N_19942,N_19653);
xor U20313 (N_20313,N_19566,N_19900);
nor U20314 (N_20314,N_19789,N_19947);
xnor U20315 (N_20315,N_19849,N_19812);
nor U20316 (N_20316,N_19784,N_19962);
and U20317 (N_20317,N_19928,N_19814);
nand U20318 (N_20318,N_19531,N_19768);
nor U20319 (N_20319,N_19581,N_19928);
nand U20320 (N_20320,N_19579,N_19817);
nand U20321 (N_20321,N_19738,N_19606);
nor U20322 (N_20322,N_19944,N_19901);
or U20323 (N_20323,N_19952,N_19872);
nand U20324 (N_20324,N_19947,N_19708);
and U20325 (N_20325,N_19748,N_19607);
xor U20326 (N_20326,N_19540,N_19526);
nand U20327 (N_20327,N_19675,N_19657);
nor U20328 (N_20328,N_19945,N_19990);
or U20329 (N_20329,N_19740,N_19869);
and U20330 (N_20330,N_19778,N_19836);
nand U20331 (N_20331,N_19608,N_19672);
xor U20332 (N_20332,N_19663,N_19930);
nand U20333 (N_20333,N_19738,N_19592);
nand U20334 (N_20334,N_19972,N_19870);
or U20335 (N_20335,N_19997,N_19656);
nor U20336 (N_20336,N_19875,N_19654);
and U20337 (N_20337,N_19545,N_19905);
and U20338 (N_20338,N_19905,N_19558);
xnor U20339 (N_20339,N_19956,N_19917);
nand U20340 (N_20340,N_19508,N_19692);
and U20341 (N_20341,N_19906,N_19659);
xor U20342 (N_20342,N_19916,N_19896);
nand U20343 (N_20343,N_19738,N_19889);
or U20344 (N_20344,N_19607,N_19783);
or U20345 (N_20345,N_19627,N_19531);
nor U20346 (N_20346,N_19715,N_19921);
nand U20347 (N_20347,N_19653,N_19991);
or U20348 (N_20348,N_19782,N_19900);
xor U20349 (N_20349,N_19986,N_19871);
or U20350 (N_20350,N_19949,N_19851);
nor U20351 (N_20351,N_19827,N_19972);
and U20352 (N_20352,N_19520,N_19870);
xor U20353 (N_20353,N_19948,N_19565);
nand U20354 (N_20354,N_19557,N_19731);
and U20355 (N_20355,N_19533,N_19772);
xnor U20356 (N_20356,N_19627,N_19720);
or U20357 (N_20357,N_19900,N_19599);
or U20358 (N_20358,N_19739,N_19900);
nand U20359 (N_20359,N_19972,N_19930);
xor U20360 (N_20360,N_19887,N_19797);
or U20361 (N_20361,N_19982,N_19659);
nand U20362 (N_20362,N_19699,N_19766);
or U20363 (N_20363,N_19751,N_19899);
nor U20364 (N_20364,N_19646,N_19650);
xor U20365 (N_20365,N_19684,N_19776);
nand U20366 (N_20366,N_19705,N_19619);
xor U20367 (N_20367,N_19895,N_19806);
and U20368 (N_20368,N_19918,N_19521);
xor U20369 (N_20369,N_19918,N_19976);
and U20370 (N_20370,N_19763,N_19854);
or U20371 (N_20371,N_19826,N_19866);
or U20372 (N_20372,N_19620,N_19639);
nand U20373 (N_20373,N_19812,N_19774);
xor U20374 (N_20374,N_19807,N_19930);
nand U20375 (N_20375,N_19765,N_19508);
or U20376 (N_20376,N_19562,N_19629);
xor U20377 (N_20377,N_19897,N_19525);
nor U20378 (N_20378,N_19896,N_19957);
and U20379 (N_20379,N_19740,N_19816);
or U20380 (N_20380,N_19834,N_19847);
nand U20381 (N_20381,N_19937,N_19779);
nand U20382 (N_20382,N_19919,N_19786);
xor U20383 (N_20383,N_19603,N_19503);
nand U20384 (N_20384,N_19752,N_19761);
nand U20385 (N_20385,N_19812,N_19768);
nand U20386 (N_20386,N_19680,N_19736);
or U20387 (N_20387,N_19805,N_19535);
xnor U20388 (N_20388,N_19779,N_19628);
nand U20389 (N_20389,N_19775,N_19883);
xnor U20390 (N_20390,N_19785,N_19790);
xor U20391 (N_20391,N_19739,N_19719);
nand U20392 (N_20392,N_19815,N_19549);
nor U20393 (N_20393,N_19893,N_19645);
or U20394 (N_20394,N_19963,N_19923);
nor U20395 (N_20395,N_19880,N_19924);
nand U20396 (N_20396,N_19692,N_19783);
nand U20397 (N_20397,N_19966,N_19859);
or U20398 (N_20398,N_19590,N_19877);
or U20399 (N_20399,N_19502,N_19545);
xnor U20400 (N_20400,N_19558,N_19731);
and U20401 (N_20401,N_19960,N_19916);
nor U20402 (N_20402,N_19952,N_19874);
or U20403 (N_20403,N_19874,N_19538);
nor U20404 (N_20404,N_19924,N_19807);
xnor U20405 (N_20405,N_19724,N_19989);
xor U20406 (N_20406,N_19794,N_19939);
or U20407 (N_20407,N_19516,N_19711);
xnor U20408 (N_20408,N_19873,N_19941);
xnor U20409 (N_20409,N_19717,N_19949);
nor U20410 (N_20410,N_19576,N_19559);
or U20411 (N_20411,N_19844,N_19836);
and U20412 (N_20412,N_19659,N_19848);
or U20413 (N_20413,N_19903,N_19789);
or U20414 (N_20414,N_19685,N_19959);
and U20415 (N_20415,N_19850,N_19996);
nand U20416 (N_20416,N_19587,N_19875);
nand U20417 (N_20417,N_19635,N_19738);
nand U20418 (N_20418,N_19564,N_19961);
and U20419 (N_20419,N_19549,N_19629);
or U20420 (N_20420,N_19593,N_19933);
and U20421 (N_20421,N_19794,N_19720);
and U20422 (N_20422,N_19734,N_19752);
and U20423 (N_20423,N_19971,N_19993);
nor U20424 (N_20424,N_19788,N_19957);
nor U20425 (N_20425,N_19522,N_19840);
and U20426 (N_20426,N_19729,N_19513);
and U20427 (N_20427,N_19652,N_19707);
nand U20428 (N_20428,N_19542,N_19905);
nor U20429 (N_20429,N_19759,N_19996);
xor U20430 (N_20430,N_19726,N_19666);
xnor U20431 (N_20431,N_19797,N_19687);
nor U20432 (N_20432,N_19588,N_19546);
xnor U20433 (N_20433,N_19734,N_19583);
nand U20434 (N_20434,N_19709,N_19760);
nor U20435 (N_20435,N_19843,N_19517);
xor U20436 (N_20436,N_19910,N_19812);
xor U20437 (N_20437,N_19704,N_19723);
nor U20438 (N_20438,N_19990,N_19921);
or U20439 (N_20439,N_19765,N_19536);
and U20440 (N_20440,N_19563,N_19723);
and U20441 (N_20441,N_19992,N_19717);
xnor U20442 (N_20442,N_19723,N_19919);
xnor U20443 (N_20443,N_19893,N_19655);
nand U20444 (N_20444,N_19630,N_19925);
or U20445 (N_20445,N_19626,N_19635);
or U20446 (N_20446,N_19516,N_19802);
xor U20447 (N_20447,N_19814,N_19561);
or U20448 (N_20448,N_19610,N_19861);
xor U20449 (N_20449,N_19536,N_19971);
nand U20450 (N_20450,N_19952,N_19844);
and U20451 (N_20451,N_19996,N_19516);
and U20452 (N_20452,N_19634,N_19618);
nand U20453 (N_20453,N_19929,N_19685);
xor U20454 (N_20454,N_19944,N_19659);
xnor U20455 (N_20455,N_19595,N_19625);
or U20456 (N_20456,N_19677,N_19651);
and U20457 (N_20457,N_19854,N_19947);
nor U20458 (N_20458,N_19540,N_19694);
xnor U20459 (N_20459,N_19868,N_19788);
or U20460 (N_20460,N_19675,N_19622);
or U20461 (N_20461,N_19839,N_19852);
nor U20462 (N_20462,N_19643,N_19755);
nand U20463 (N_20463,N_19705,N_19516);
or U20464 (N_20464,N_19849,N_19581);
nor U20465 (N_20465,N_19962,N_19976);
or U20466 (N_20466,N_19652,N_19515);
or U20467 (N_20467,N_19965,N_19846);
and U20468 (N_20468,N_19907,N_19773);
nor U20469 (N_20469,N_19767,N_19677);
nand U20470 (N_20470,N_19977,N_19566);
nor U20471 (N_20471,N_19616,N_19579);
or U20472 (N_20472,N_19815,N_19923);
nand U20473 (N_20473,N_19727,N_19752);
or U20474 (N_20474,N_19787,N_19963);
xnor U20475 (N_20475,N_19786,N_19663);
or U20476 (N_20476,N_19543,N_19515);
nor U20477 (N_20477,N_19647,N_19531);
and U20478 (N_20478,N_19928,N_19665);
nand U20479 (N_20479,N_19713,N_19763);
nand U20480 (N_20480,N_19565,N_19847);
and U20481 (N_20481,N_19841,N_19974);
nor U20482 (N_20482,N_19589,N_19865);
nor U20483 (N_20483,N_19517,N_19645);
nor U20484 (N_20484,N_19835,N_19564);
xor U20485 (N_20485,N_19795,N_19651);
and U20486 (N_20486,N_19834,N_19931);
xnor U20487 (N_20487,N_19949,N_19660);
nand U20488 (N_20488,N_19816,N_19859);
xor U20489 (N_20489,N_19750,N_19601);
and U20490 (N_20490,N_19634,N_19934);
nand U20491 (N_20491,N_19891,N_19889);
and U20492 (N_20492,N_19714,N_19595);
nor U20493 (N_20493,N_19689,N_19965);
xor U20494 (N_20494,N_19581,N_19833);
nand U20495 (N_20495,N_19764,N_19658);
or U20496 (N_20496,N_19912,N_19609);
or U20497 (N_20497,N_19924,N_19960);
or U20498 (N_20498,N_19523,N_19595);
nor U20499 (N_20499,N_19540,N_19889);
xnor U20500 (N_20500,N_20128,N_20354);
or U20501 (N_20501,N_20374,N_20277);
or U20502 (N_20502,N_20425,N_20017);
or U20503 (N_20503,N_20152,N_20148);
nor U20504 (N_20504,N_20295,N_20289);
xnor U20505 (N_20505,N_20081,N_20058);
nand U20506 (N_20506,N_20196,N_20229);
nor U20507 (N_20507,N_20411,N_20257);
nor U20508 (N_20508,N_20134,N_20205);
and U20509 (N_20509,N_20047,N_20497);
xor U20510 (N_20510,N_20048,N_20307);
or U20511 (N_20511,N_20076,N_20139);
and U20512 (N_20512,N_20288,N_20266);
nor U20513 (N_20513,N_20328,N_20493);
nand U20514 (N_20514,N_20223,N_20285);
and U20515 (N_20515,N_20206,N_20075);
nor U20516 (N_20516,N_20440,N_20358);
or U20517 (N_20517,N_20439,N_20167);
xnor U20518 (N_20518,N_20299,N_20218);
nand U20519 (N_20519,N_20261,N_20476);
or U20520 (N_20520,N_20136,N_20451);
nor U20521 (N_20521,N_20038,N_20039);
and U20522 (N_20522,N_20292,N_20077);
xnor U20523 (N_20523,N_20499,N_20453);
and U20524 (N_20524,N_20007,N_20385);
nand U20525 (N_20525,N_20060,N_20030);
nand U20526 (N_20526,N_20464,N_20387);
or U20527 (N_20527,N_20325,N_20129);
nand U20528 (N_20528,N_20384,N_20191);
nor U20529 (N_20529,N_20090,N_20226);
xnor U20530 (N_20530,N_20118,N_20303);
or U20531 (N_20531,N_20062,N_20316);
nor U20532 (N_20532,N_20122,N_20403);
nor U20533 (N_20533,N_20203,N_20079);
nor U20534 (N_20534,N_20146,N_20008);
and U20535 (N_20535,N_20315,N_20236);
and U20536 (N_20536,N_20197,N_20485);
xnor U20537 (N_20537,N_20388,N_20249);
nand U20538 (N_20538,N_20297,N_20116);
xnor U20539 (N_20539,N_20399,N_20138);
nand U20540 (N_20540,N_20482,N_20086);
and U20541 (N_20541,N_20431,N_20341);
nor U20542 (N_20542,N_20174,N_20392);
or U20543 (N_20543,N_20274,N_20020);
xnor U20544 (N_20544,N_20127,N_20145);
or U20545 (N_20545,N_20246,N_20421);
or U20546 (N_20546,N_20481,N_20153);
nor U20547 (N_20547,N_20298,N_20462);
nand U20548 (N_20548,N_20260,N_20262);
nor U20549 (N_20549,N_20071,N_20478);
nand U20550 (N_20550,N_20267,N_20084);
nor U20551 (N_20551,N_20068,N_20106);
and U20552 (N_20552,N_20016,N_20487);
nand U20553 (N_20553,N_20092,N_20245);
or U20554 (N_20554,N_20345,N_20396);
or U20555 (N_20555,N_20404,N_20456);
nor U20556 (N_20556,N_20103,N_20158);
nand U20557 (N_20557,N_20053,N_20067);
nand U20558 (N_20558,N_20009,N_20083);
and U20559 (N_20559,N_20104,N_20415);
and U20560 (N_20560,N_20042,N_20240);
or U20561 (N_20561,N_20323,N_20331);
nor U20562 (N_20562,N_20194,N_20386);
nor U20563 (N_20563,N_20488,N_20368);
or U20564 (N_20564,N_20330,N_20375);
and U20565 (N_20565,N_20013,N_20473);
and U20566 (N_20566,N_20112,N_20034);
xnor U20567 (N_20567,N_20347,N_20044);
nand U20568 (N_20568,N_20426,N_20114);
and U20569 (N_20569,N_20416,N_20449);
or U20570 (N_20570,N_20018,N_20061);
nor U20571 (N_20571,N_20282,N_20454);
and U20572 (N_20572,N_20241,N_20459);
nand U20573 (N_20573,N_20093,N_20147);
xnor U20574 (N_20574,N_20169,N_20010);
and U20575 (N_20575,N_20209,N_20037);
or U20576 (N_20576,N_20438,N_20164);
xor U20577 (N_20577,N_20452,N_20135);
nor U20578 (N_20578,N_20435,N_20317);
nand U20579 (N_20579,N_20235,N_20243);
and U20580 (N_20580,N_20200,N_20064);
xor U20581 (N_20581,N_20367,N_20220);
or U20582 (N_20582,N_20442,N_20265);
nor U20583 (N_20583,N_20309,N_20159);
or U20584 (N_20584,N_20080,N_20052);
nand U20585 (N_20585,N_20172,N_20160);
nor U20586 (N_20586,N_20329,N_20019);
nor U20587 (N_20587,N_20308,N_20176);
xor U20588 (N_20588,N_20322,N_20259);
and U20589 (N_20589,N_20348,N_20162);
nor U20590 (N_20590,N_20085,N_20320);
xor U20591 (N_20591,N_20130,N_20254);
xnor U20592 (N_20592,N_20326,N_20340);
nor U20593 (N_20593,N_20429,N_20377);
xor U20594 (N_20594,N_20324,N_20140);
or U20595 (N_20595,N_20069,N_20380);
xor U20596 (N_20596,N_20394,N_20074);
or U20597 (N_20597,N_20263,N_20110);
nor U20598 (N_20598,N_20496,N_20190);
nor U20599 (N_20599,N_20369,N_20357);
or U20600 (N_20600,N_20175,N_20397);
xor U20601 (N_20601,N_20321,N_20001);
nand U20602 (N_20602,N_20187,N_20359);
or U20603 (N_20603,N_20381,N_20418);
xor U20604 (N_20604,N_20371,N_20410);
and U20605 (N_20605,N_20225,N_20272);
nand U20606 (N_20606,N_20054,N_20212);
nor U20607 (N_20607,N_20228,N_20204);
nand U20608 (N_20608,N_20180,N_20311);
xor U20609 (N_20609,N_20021,N_20268);
and U20610 (N_20610,N_20498,N_20005);
xor U20611 (N_20611,N_20433,N_20012);
xor U20612 (N_20612,N_20355,N_20364);
nor U20613 (N_20613,N_20361,N_20370);
and U20614 (N_20614,N_20287,N_20336);
or U20615 (N_20615,N_20484,N_20255);
xnor U20616 (N_20616,N_20294,N_20366);
xor U20617 (N_20617,N_20281,N_20408);
and U20618 (N_20618,N_20306,N_20201);
nor U20619 (N_20619,N_20003,N_20471);
and U20620 (N_20620,N_20231,N_20000);
nor U20621 (N_20621,N_20419,N_20474);
and U20622 (N_20622,N_20319,N_20137);
xor U20623 (N_20623,N_20372,N_20428);
xor U20624 (N_20624,N_20144,N_20441);
nor U20625 (N_20625,N_20269,N_20273);
nand U20626 (N_20626,N_20099,N_20207);
and U20627 (N_20627,N_20445,N_20495);
and U20628 (N_20628,N_20447,N_20275);
xor U20629 (N_20629,N_20125,N_20035);
and U20630 (N_20630,N_20480,N_20107);
nand U20631 (N_20631,N_20237,N_20105);
or U20632 (N_20632,N_20344,N_20252);
nand U20633 (N_20633,N_20166,N_20465);
or U20634 (N_20634,N_20470,N_20436);
nor U20635 (N_20635,N_20494,N_20171);
xor U20636 (N_20636,N_20216,N_20406);
or U20637 (N_20637,N_20043,N_20089);
nand U20638 (N_20638,N_20333,N_20184);
or U20639 (N_20639,N_20391,N_20072);
nand U20640 (N_20640,N_20490,N_20213);
nor U20641 (N_20641,N_20227,N_20131);
nor U20642 (N_20642,N_20132,N_20041);
or U20643 (N_20643,N_20115,N_20117);
nand U20644 (N_20644,N_20270,N_20221);
or U20645 (N_20645,N_20046,N_20278);
and U20646 (N_20646,N_20430,N_20024);
xor U20647 (N_20647,N_20489,N_20242);
or U20648 (N_20648,N_20455,N_20458);
or U20649 (N_20649,N_20350,N_20014);
xor U20650 (N_20650,N_20383,N_20011);
xor U20651 (N_20651,N_20006,N_20379);
nand U20652 (N_20652,N_20256,N_20168);
or U20653 (N_20653,N_20101,N_20179);
and U20654 (N_20654,N_20432,N_20457);
nor U20655 (N_20655,N_20351,N_20126);
and U20656 (N_20656,N_20025,N_20199);
nor U20657 (N_20657,N_20097,N_20477);
nor U20658 (N_20658,N_20049,N_20078);
nand U20659 (N_20659,N_20423,N_20113);
nor U20660 (N_20660,N_20305,N_20376);
xnor U20661 (N_20661,N_20479,N_20123);
nor U20662 (N_20662,N_20318,N_20405);
or U20663 (N_20663,N_20286,N_20301);
xor U20664 (N_20664,N_20100,N_20182);
or U20665 (N_20665,N_20027,N_20091);
and U20666 (N_20666,N_20239,N_20335);
and U20667 (N_20667,N_20393,N_20193);
nor U20668 (N_20668,N_20198,N_20143);
xnor U20669 (N_20669,N_20181,N_20163);
or U20670 (N_20670,N_20119,N_20082);
and U20671 (N_20671,N_20304,N_20302);
nand U20672 (N_20672,N_20264,N_20310);
and U20673 (N_20673,N_20141,N_20186);
or U20674 (N_20674,N_20469,N_20032);
and U20675 (N_20675,N_20395,N_20155);
and U20676 (N_20676,N_20059,N_20211);
nand U20677 (N_20677,N_20202,N_20483);
nand U20678 (N_20678,N_20422,N_20448);
and U20679 (N_20679,N_20248,N_20356);
nand U20680 (N_20680,N_20300,N_20382);
nand U20681 (N_20681,N_20353,N_20293);
or U20682 (N_20682,N_20258,N_20291);
nor U20683 (N_20683,N_20414,N_20028);
nor U20684 (N_20684,N_20466,N_20444);
or U20685 (N_20685,N_20102,N_20446);
and U20686 (N_20686,N_20398,N_20070);
nor U20687 (N_20687,N_20427,N_20156);
nor U20688 (N_20688,N_20098,N_20029);
nand U20689 (N_20689,N_20151,N_20189);
xnor U20690 (N_20690,N_20271,N_20339);
nand U20691 (N_20691,N_20251,N_20230);
and U20692 (N_20692,N_20343,N_20088);
xnor U20693 (N_20693,N_20023,N_20040);
or U20694 (N_20694,N_20036,N_20349);
xor U20695 (N_20695,N_20360,N_20332);
or U20696 (N_20696,N_20337,N_20002);
nor U20697 (N_20697,N_20121,N_20409);
or U20698 (N_20698,N_20401,N_20362);
nand U20699 (N_20699,N_20033,N_20327);
or U20700 (N_20700,N_20334,N_20051);
nand U20701 (N_20701,N_20420,N_20214);
or U20702 (N_20702,N_20312,N_20283);
and U20703 (N_20703,N_20015,N_20413);
nor U20704 (N_20704,N_20177,N_20234);
or U20705 (N_20705,N_20313,N_20183);
nor U20706 (N_20706,N_20342,N_20279);
nor U20707 (N_20707,N_20486,N_20095);
nor U20708 (N_20708,N_20157,N_20210);
nand U20709 (N_20709,N_20412,N_20450);
nand U20710 (N_20710,N_20276,N_20468);
nor U20711 (N_20711,N_20284,N_20224);
nor U20712 (N_20712,N_20253,N_20378);
nand U20713 (N_20713,N_20232,N_20031);
xor U20714 (N_20714,N_20400,N_20463);
nor U20715 (N_20715,N_20443,N_20004);
nand U20716 (N_20716,N_20154,N_20178);
or U20717 (N_20717,N_20250,N_20390);
xor U20718 (N_20718,N_20461,N_20050);
and U20719 (N_20719,N_20363,N_20402);
and U20720 (N_20720,N_20094,N_20109);
or U20721 (N_20721,N_20238,N_20215);
or U20722 (N_20722,N_20165,N_20407);
nor U20723 (N_20723,N_20045,N_20195);
or U20724 (N_20724,N_20222,N_20108);
or U20725 (N_20725,N_20247,N_20296);
or U20726 (N_20726,N_20149,N_20365);
or U20727 (N_20727,N_20389,N_20056);
xnor U20728 (N_20728,N_20026,N_20492);
nand U20729 (N_20729,N_20022,N_20066);
and U20730 (N_20730,N_20065,N_20472);
nand U20731 (N_20731,N_20133,N_20437);
and U20732 (N_20732,N_20208,N_20073);
nor U20733 (N_20733,N_20290,N_20314);
nor U20734 (N_20734,N_20244,N_20111);
xor U20735 (N_20735,N_20192,N_20417);
or U20736 (N_20736,N_20233,N_20434);
or U20737 (N_20737,N_20063,N_20188);
and U20738 (N_20738,N_20219,N_20170);
or U20739 (N_20739,N_20373,N_20142);
nor U20740 (N_20740,N_20055,N_20338);
and U20741 (N_20741,N_20087,N_20173);
nand U20742 (N_20742,N_20120,N_20185);
xor U20743 (N_20743,N_20096,N_20467);
nor U20744 (N_20744,N_20150,N_20491);
xnor U20745 (N_20745,N_20475,N_20217);
nor U20746 (N_20746,N_20352,N_20124);
nand U20747 (N_20747,N_20460,N_20280);
or U20748 (N_20748,N_20161,N_20424);
nor U20749 (N_20749,N_20346,N_20057);
nand U20750 (N_20750,N_20329,N_20416);
nand U20751 (N_20751,N_20369,N_20395);
and U20752 (N_20752,N_20127,N_20433);
xnor U20753 (N_20753,N_20263,N_20480);
xor U20754 (N_20754,N_20105,N_20297);
nand U20755 (N_20755,N_20270,N_20284);
nand U20756 (N_20756,N_20108,N_20022);
xor U20757 (N_20757,N_20477,N_20391);
xnor U20758 (N_20758,N_20399,N_20265);
xor U20759 (N_20759,N_20181,N_20214);
nand U20760 (N_20760,N_20009,N_20350);
or U20761 (N_20761,N_20313,N_20444);
xnor U20762 (N_20762,N_20154,N_20225);
xnor U20763 (N_20763,N_20053,N_20086);
nand U20764 (N_20764,N_20395,N_20321);
nand U20765 (N_20765,N_20385,N_20034);
or U20766 (N_20766,N_20386,N_20316);
nand U20767 (N_20767,N_20245,N_20084);
nor U20768 (N_20768,N_20379,N_20043);
or U20769 (N_20769,N_20249,N_20268);
and U20770 (N_20770,N_20222,N_20090);
nand U20771 (N_20771,N_20249,N_20286);
and U20772 (N_20772,N_20277,N_20199);
or U20773 (N_20773,N_20208,N_20151);
or U20774 (N_20774,N_20134,N_20160);
or U20775 (N_20775,N_20279,N_20394);
xnor U20776 (N_20776,N_20142,N_20357);
nor U20777 (N_20777,N_20372,N_20033);
nor U20778 (N_20778,N_20359,N_20078);
or U20779 (N_20779,N_20342,N_20095);
nor U20780 (N_20780,N_20268,N_20398);
xor U20781 (N_20781,N_20491,N_20326);
and U20782 (N_20782,N_20305,N_20180);
xor U20783 (N_20783,N_20269,N_20452);
nor U20784 (N_20784,N_20047,N_20480);
or U20785 (N_20785,N_20194,N_20125);
xor U20786 (N_20786,N_20026,N_20183);
or U20787 (N_20787,N_20387,N_20429);
and U20788 (N_20788,N_20479,N_20046);
and U20789 (N_20789,N_20089,N_20037);
nor U20790 (N_20790,N_20093,N_20455);
or U20791 (N_20791,N_20118,N_20310);
xor U20792 (N_20792,N_20182,N_20261);
nand U20793 (N_20793,N_20464,N_20014);
xnor U20794 (N_20794,N_20033,N_20053);
or U20795 (N_20795,N_20454,N_20185);
nand U20796 (N_20796,N_20440,N_20311);
or U20797 (N_20797,N_20281,N_20038);
nand U20798 (N_20798,N_20189,N_20135);
xnor U20799 (N_20799,N_20467,N_20314);
xnor U20800 (N_20800,N_20113,N_20043);
or U20801 (N_20801,N_20108,N_20075);
and U20802 (N_20802,N_20374,N_20455);
or U20803 (N_20803,N_20300,N_20138);
xor U20804 (N_20804,N_20317,N_20162);
or U20805 (N_20805,N_20073,N_20278);
or U20806 (N_20806,N_20433,N_20132);
and U20807 (N_20807,N_20271,N_20020);
nand U20808 (N_20808,N_20326,N_20308);
nand U20809 (N_20809,N_20376,N_20368);
nor U20810 (N_20810,N_20336,N_20054);
xnor U20811 (N_20811,N_20329,N_20352);
nor U20812 (N_20812,N_20318,N_20042);
xnor U20813 (N_20813,N_20441,N_20217);
or U20814 (N_20814,N_20030,N_20360);
xnor U20815 (N_20815,N_20242,N_20101);
and U20816 (N_20816,N_20014,N_20118);
nor U20817 (N_20817,N_20101,N_20349);
nand U20818 (N_20818,N_20420,N_20313);
or U20819 (N_20819,N_20465,N_20494);
nand U20820 (N_20820,N_20100,N_20125);
xnor U20821 (N_20821,N_20177,N_20154);
xor U20822 (N_20822,N_20179,N_20195);
nor U20823 (N_20823,N_20196,N_20096);
nor U20824 (N_20824,N_20438,N_20139);
and U20825 (N_20825,N_20203,N_20336);
nor U20826 (N_20826,N_20235,N_20245);
and U20827 (N_20827,N_20089,N_20173);
nor U20828 (N_20828,N_20472,N_20453);
xor U20829 (N_20829,N_20175,N_20318);
nor U20830 (N_20830,N_20253,N_20455);
or U20831 (N_20831,N_20195,N_20129);
xnor U20832 (N_20832,N_20241,N_20344);
nand U20833 (N_20833,N_20310,N_20366);
xnor U20834 (N_20834,N_20469,N_20160);
or U20835 (N_20835,N_20221,N_20423);
or U20836 (N_20836,N_20374,N_20226);
nor U20837 (N_20837,N_20355,N_20090);
and U20838 (N_20838,N_20475,N_20208);
or U20839 (N_20839,N_20304,N_20456);
or U20840 (N_20840,N_20116,N_20000);
and U20841 (N_20841,N_20079,N_20209);
xnor U20842 (N_20842,N_20168,N_20357);
or U20843 (N_20843,N_20475,N_20216);
nand U20844 (N_20844,N_20009,N_20277);
xor U20845 (N_20845,N_20390,N_20001);
nor U20846 (N_20846,N_20188,N_20129);
or U20847 (N_20847,N_20299,N_20285);
and U20848 (N_20848,N_20046,N_20448);
nor U20849 (N_20849,N_20426,N_20276);
and U20850 (N_20850,N_20305,N_20022);
xor U20851 (N_20851,N_20459,N_20463);
xnor U20852 (N_20852,N_20223,N_20313);
nand U20853 (N_20853,N_20270,N_20095);
and U20854 (N_20854,N_20375,N_20392);
nand U20855 (N_20855,N_20250,N_20441);
nand U20856 (N_20856,N_20429,N_20277);
xnor U20857 (N_20857,N_20185,N_20408);
or U20858 (N_20858,N_20327,N_20252);
and U20859 (N_20859,N_20486,N_20226);
xor U20860 (N_20860,N_20195,N_20299);
xnor U20861 (N_20861,N_20233,N_20360);
nand U20862 (N_20862,N_20478,N_20086);
and U20863 (N_20863,N_20315,N_20131);
xnor U20864 (N_20864,N_20027,N_20490);
and U20865 (N_20865,N_20145,N_20380);
and U20866 (N_20866,N_20155,N_20021);
or U20867 (N_20867,N_20089,N_20244);
nor U20868 (N_20868,N_20353,N_20443);
nand U20869 (N_20869,N_20484,N_20083);
xnor U20870 (N_20870,N_20170,N_20147);
nand U20871 (N_20871,N_20328,N_20374);
nor U20872 (N_20872,N_20397,N_20164);
or U20873 (N_20873,N_20167,N_20070);
or U20874 (N_20874,N_20109,N_20479);
xnor U20875 (N_20875,N_20222,N_20415);
nor U20876 (N_20876,N_20287,N_20011);
xnor U20877 (N_20877,N_20451,N_20062);
nor U20878 (N_20878,N_20465,N_20067);
or U20879 (N_20879,N_20267,N_20375);
and U20880 (N_20880,N_20239,N_20304);
nor U20881 (N_20881,N_20147,N_20278);
nand U20882 (N_20882,N_20408,N_20427);
xnor U20883 (N_20883,N_20221,N_20045);
nand U20884 (N_20884,N_20110,N_20480);
nand U20885 (N_20885,N_20359,N_20392);
xnor U20886 (N_20886,N_20356,N_20155);
nor U20887 (N_20887,N_20006,N_20256);
xor U20888 (N_20888,N_20327,N_20388);
and U20889 (N_20889,N_20113,N_20189);
and U20890 (N_20890,N_20471,N_20202);
nor U20891 (N_20891,N_20158,N_20065);
xor U20892 (N_20892,N_20124,N_20146);
and U20893 (N_20893,N_20033,N_20000);
or U20894 (N_20894,N_20040,N_20453);
and U20895 (N_20895,N_20301,N_20395);
nor U20896 (N_20896,N_20242,N_20024);
nor U20897 (N_20897,N_20482,N_20103);
xnor U20898 (N_20898,N_20421,N_20211);
or U20899 (N_20899,N_20277,N_20385);
or U20900 (N_20900,N_20419,N_20252);
nand U20901 (N_20901,N_20068,N_20432);
and U20902 (N_20902,N_20326,N_20061);
xnor U20903 (N_20903,N_20432,N_20062);
nand U20904 (N_20904,N_20227,N_20021);
nor U20905 (N_20905,N_20063,N_20199);
xnor U20906 (N_20906,N_20350,N_20443);
nand U20907 (N_20907,N_20270,N_20066);
or U20908 (N_20908,N_20204,N_20277);
nand U20909 (N_20909,N_20363,N_20482);
xnor U20910 (N_20910,N_20204,N_20456);
nand U20911 (N_20911,N_20272,N_20086);
or U20912 (N_20912,N_20050,N_20217);
nand U20913 (N_20913,N_20322,N_20087);
nand U20914 (N_20914,N_20133,N_20131);
xnor U20915 (N_20915,N_20238,N_20451);
nand U20916 (N_20916,N_20139,N_20462);
nor U20917 (N_20917,N_20038,N_20465);
xor U20918 (N_20918,N_20254,N_20465);
nand U20919 (N_20919,N_20117,N_20404);
or U20920 (N_20920,N_20447,N_20444);
and U20921 (N_20921,N_20239,N_20369);
nor U20922 (N_20922,N_20340,N_20252);
and U20923 (N_20923,N_20433,N_20453);
xor U20924 (N_20924,N_20396,N_20038);
nand U20925 (N_20925,N_20077,N_20449);
nor U20926 (N_20926,N_20312,N_20402);
xor U20927 (N_20927,N_20492,N_20140);
nor U20928 (N_20928,N_20012,N_20404);
nand U20929 (N_20929,N_20225,N_20310);
xor U20930 (N_20930,N_20127,N_20093);
and U20931 (N_20931,N_20124,N_20226);
nand U20932 (N_20932,N_20052,N_20361);
nor U20933 (N_20933,N_20369,N_20330);
or U20934 (N_20934,N_20042,N_20063);
and U20935 (N_20935,N_20041,N_20225);
or U20936 (N_20936,N_20389,N_20311);
nor U20937 (N_20937,N_20222,N_20186);
nand U20938 (N_20938,N_20308,N_20229);
nand U20939 (N_20939,N_20222,N_20372);
and U20940 (N_20940,N_20213,N_20318);
or U20941 (N_20941,N_20400,N_20410);
nand U20942 (N_20942,N_20140,N_20044);
nand U20943 (N_20943,N_20268,N_20066);
nand U20944 (N_20944,N_20402,N_20435);
or U20945 (N_20945,N_20172,N_20330);
xnor U20946 (N_20946,N_20130,N_20253);
xnor U20947 (N_20947,N_20307,N_20092);
and U20948 (N_20948,N_20144,N_20112);
and U20949 (N_20949,N_20238,N_20199);
xor U20950 (N_20950,N_20342,N_20398);
and U20951 (N_20951,N_20463,N_20032);
or U20952 (N_20952,N_20285,N_20160);
and U20953 (N_20953,N_20318,N_20297);
or U20954 (N_20954,N_20427,N_20041);
nand U20955 (N_20955,N_20350,N_20196);
nand U20956 (N_20956,N_20301,N_20448);
nor U20957 (N_20957,N_20025,N_20340);
or U20958 (N_20958,N_20421,N_20073);
nor U20959 (N_20959,N_20027,N_20290);
or U20960 (N_20960,N_20031,N_20121);
and U20961 (N_20961,N_20446,N_20416);
xnor U20962 (N_20962,N_20038,N_20088);
and U20963 (N_20963,N_20115,N_20449);
xor U20964 (N_20964,N_20254,N_20251);
xnor U20965 (N_20965,N_20250,N_20320);
xor U20966 (N_20966,N_20263,N_20111);
xnor U20967 (N_20967,N_20147,N_20013);
and U20968 (N_20968,N_20396,N_20008);
nor U20969 (N_20969,N_20032,N_20392);
xor U20970 (N_20970,N_20032,N_20386);
and U20971 (N_20971,N_20216,N_20211);
nor U20972 (N_20972,N_20063,N_20372);
xnor U20973 (N_20973,N_20339,N_20421);
nand U20974 (N_20974,N_20342,N_20421);
and U20975 (N_20975,N_20368,N_20342);
nor U20976 (N_20976,N_20399,N_20257);
or U20977 (N_20977,N_20313,N_20226);
nand U20978 (N_20978,N_20381,N_20451);
or U20979 (N_20979,N_20413,N_20189);
and U20980 (N_20980,N_20302,N_20359);
or U20981 (N_20981,N_20342,N_20117);
and U20982 (N_20982,N_20340,N_20201);
or U20983 (N_20983,N_20285,N_20131);
xor U20984 (N_20984,N_20391,N_20262);
nor U20985 (N_20985,N_20388,N_20330);
or U20986 (N_20986,N_20434,N_20219);
or U20987 (N_20987,N_20017,N_20046);
and U20988 (N_20988,N_20101,N_20124);
and U20989 (N_20989,N_20256,N_20423);
nand U20990 (N_20990,N_20316,N_20118);
and U20991 (N_20991,N_20190,N_20019);
and U20992 (N_20992,N_20388,N_20118);
nand U20993 (N_20993,N_20303,N_20081);
nor U20994 (N_20994,N_20303,N_20181);
nor U20995 (N_20995,N_20244,N_20420);
xnor U20996 (N_20996,N_20187,N_20489);
nor U20997 (N_20997,N_20297,N_20398);
xor U20998 (N_20998,N_20454,N_20021);
and U20999 (N_20999,N_20016,N_20344);
or U21000 (N_21000,N_20913,N_20509);
nor U21001 (N_21001,N_20689,N_20653);
or U21002 (N_21002,N_20918,N_20784);
xnor U21003 (N_21003,N_20511,N_20774);
nor U21004 (N_21004,N_20963,N_20856);
xor U21005 (N_21005,N_20522,N_20817);
xor U21006 (N_21006,N_20923,N_20569);
nor U21007 (N_21007,N_20515,N_20897);
or U21008 (N_21008,N_20749,N_20674);
or U21009 (N_21009,N_20872,N_20989);
nand U21010 (N_21010,N_20628,N_20852);
xor U21011 (N_21011,N_20928,N_20639);
nor U21012 (N_21012,N_20627,N_20590);
xnor U21013 (N_21013,N_20781,N_20854);
xor U21014 (N_21014,N_20502,N_20768);
and U21015 (N_21015,N_20765,N_20895);
xor U21016 (N_21016,N_20564,N_20646);
nand U21017 (N_21017,N_20953,N_20952);
and U21018 (N_21018,N_20920,N_20853);
xor U21019 (N_21019,N_20779,N_20876);
nor U21020 (N_21020,N_20926,N_20772);
nand U21021 (N_21021,N_20524,N_20761);
nand U21022 (N_21022,N_20724,N_20655);
nand U21023 (N_21023,N_20911,N_20969);
nor U21024 (N_21024,N_20871,N_20507);
nand U21025 (N_21025,N_20747,N_20946);
and U21026 (N_21026,N_20583,N_20565);
or U21027 (N_21027,N_20543,N_20990);
xnor U21028 (N_21028,N_20540,N_20883);
nand U21029 (N_21029,N_20755,N_20991);
xnor U21030 (N_21030,N_20889,N_20710);
nor U21031 (N_21031,N_20916,N_20695);
nor U21032 (N_21032,N_20822,N_20669);
xnor U21033 (N_21033,N_20944,N_20578);
xnor U21034 (N_21034,N_20932,N_20503);
nor U21035 (N_21035,N_20940,N_20589);
xor U21036 (N_21036,N_20796,N_20754);
xor U21037 (N_21037,N_20780,N_20542);
nand U21038 (N_21038,N_20942,N_20976);
or U21039 (N_21039,N_20984,N_20967);
nor U21040 (N_21040,N_20819,N_20869);
and U21041 (N_21041,N_20767,N_20758);
or U21042 (N_21042,N_20974,N_20592);
nand U21043 (N_21043,N_20892,N_20548);
nor U21044 (N_21044,N_20673,N_20625);
nand U21045 (N_21045,N_20824,N_20864);
and U21046 (N_21046,N_20823,N_20997);
or U21047 (N_21047,N_20818,N_20785);
nor U21048 (N_21048,N_20603,N_20732);
nor U21049 (N_21049,N_20786,N_20721);
nor U21050 (N_21050,N_20850,N_20868);
xnor U21051 (N_21051,N_20679,N_20968);
or U21052 (N_21052,N_20688,N_20863);
nand U21053 (N_21053,N_20901,N_20567);
nand U21054 (N_21054,N_20613,N_20925);
or U21055 (N_21055,N_20921,N_20951);
or U21056 (N_21056,N_20577,N_20593);
xnor U21057 (N_21057,N_20844,N_20987);
xnor U21058 (N_21058,N_20641,N_20720);
nor U21059 (N_21059,N_20960,N_20650);
and U21060 (N_21060,N_20829,N_20741);
or U21061 (N_21061,N_20604,N_20830);
nand U21062 (N_21062,N_20793,N_20759);
xnor U21063 (N_21063,N_20644,N_20513);
and U21064 (N_21064,N_20805,N_20675);
xor U21065 (N_21065,N_20715,N_20594);
xor U21066 (N_21066,N_20722,N_20909);
xnor U21067 (N_21067,N_20668,N_20744);
and U21068 (N_21068,N_20566,N_20531);
nor U21069 (N_21069,N_20530,N_20643);
and U21070 (N_21070,N_20701,N_20843);
and U21071 (N_21071,N_20563,N_20894);
nor U21072 (N_21072,N_20615,N_20683);
nand U21073 (N_21073,N_20685,N_20803);
and U21074 (N_21074,N_20927,N_20654);
nor U21075 (N_21075,N_20882,N_20791);
and U21076 (N_21076,N_20813,N_20560);
or U21077 (N_21077,N_20880,N_20866);
xnor U21078 (N_21078,N_20687,N_20988);
or U21079 (N_21079,N_20705,N_20551);
or U21080 (N_21080,N_20919,N_20649);
nor U21081 (N_21081,N_20506,N_20664);
nand U21082 (N_21082,N_20684,N_20908);
and U21083 (N_21083,N_20900,N_20562);
nor U21084 (N_21084,N_20645,N_20535);
nor U21085 (N_21085,N_20745,N_20660);
xor U21086 (N_21086,N_20519,N_20572);
nor U21087 (N_21087,N_20873,N_20978);
xor U21088 (N_21088,N_20550,N_20626);
and U21089 (N_21089,N_20751,N_20945);
and U21090 (N_21090,N_20526,N_20523);
and U21091 (N_21091,N_20504,N_20956);
or U21092 (N_21092,N_20835,N_20996);
nor U21093 (N_21093,N_20518,N_20832);
nor U21094 (N_21094,N_20712,N_20686);
or U21095 (N_21095,N_20962,N_20561);
nor U21096 (N_21096,N_20777,N_20771);
or U21097 (N_21097,N_20552,N_20579);
and U21098 (N_21098,N_20955,N_20611);
or U21099 (N_21099,N_20616,N_20647);
nand U21100 (N_21100,N_20973,N_20608);
xnor U21101 (N_21101,N_20922,N_20587);
nor U21102 (N_21102,N_20612,N_20861);
or U21103 (N_21103,N_20862,N_20792);
nand U21104 (N_21104,N_20776,N_20640);
nor U21105 (N_21105,N_20949,N_20731);
nand U21106 (N_21106,N_20708,N_20541);
or U21107 (N_21107,N_20762,N_20677);
nor U21108 (N_21108,N_20533,N_20851);
and U21109 (N_21109,N_20521,N_20929);
nand U21110 (N_21110,N_20773,N_20971);
nor U21111 (N_21111,N_20580,N_20651);
nor U21112 (N_21112,N_20727,N_20941);
nor U21113 (N_21113,N_20766,N_20980);
nor U21114 (N_21114,N_20898,N_20828);
nor U21115 (N_21115,N_20778,N_20717);
nor U21116 (N_21116,N_20801,N_20757);
or U21117 (N_21117,N_20847,N_20995);
xor U21118 (N_21118,N_20575,N_20881);
nand U21119 (N_21119,N_20825,N_20618);
xnor U21120 (N_21120,N_20576,N_20623);
or U21121 (N_21121,N_20877,N_20586);
xnor U21122 (N_21122,N_20691,N_20716);
xor U21123 (N_21123,N_20887,N_20948);
nor U21124 (N_21124,N_20875,N_20680);
and U21125 (N_21125,N_20734,N_20811);
nand U21126 (N_21126,N_20624,N_20756);
and U21127 (N_21127,N_20975,N_20657);
or U21128 (N_21128,N_20840,N_20665);
and U21129 (N_21129,N_20516,N_20858);
xor U21130 (N_21130,N_20571,N_20638);
xnor U21131 (N_21131,N_20831,N_20886);
nand U21132 (N_21132,N_20934,N_20808);
or U21133 (N_21133,N_20848,N_20707);
nand U21134 (N_21134,N_20917,N_20525);
xnor U21135 (N_21135,N_20692,N_20888);
nand U21136 (N_21136,N_20555,N_20965);
or U21137 (N_21137,N_20939,N_20821);
or U21138 (N_21138,N_20964,N_20902);
nor U21139 (N_21139,N_20558,N_20702);
nor U21140 (N_21140,N_20750,N_20737);
nand U21141 (N_21141,N_20536,N_20982);
or U21142 (N_21142,N_20999,N_20812);
and U21143 (N_21143,N_20763,N_20826);
nand U21144 (N_21144,N_20528,N_20719);
nand U21145 (N_21145,N_20947,N_20827);
xnor U21146 (N_21146,N_20709,N_20595);
or U21147 (N_21147,N_20936,N_20814);
nand U21148 (N_21148,N_20573,N_20859);
nand U21149 (N_21149,N_20570,N_20910);
nand U21150 (N_21150,N_20954,N_20787);
xor U21151 (N_21151,N_20652,N_20802);
nor U21152 (N_21152,N_20617,N_20568);
nand U21153 (N_21153,N_20879,N_20591);
nor U21154 (N_21154,N_20769,N_20714);
xor U21155 (N_21155,N_20635,N_20725);
or U21156 (N_21156,N_20730,N_20697);
nand U21157 (N_21157,N_20748,N_20820);
nor U21158 (N_21158,N_20998,N_20544);
and U21159 (N_21159,N_20703,N_20678);
xnor U21160 (N_21160,N_20581,N_20743);
nor U21161 (N_21161,N_20903,N_20694);
and U21162 (N_21162,N_20728,N_20662);
and U21163 (N_21163,N_20896,N_20809);
nand U21164 (N_21164,N_20607,N_20596);
nor U21165 (N_21165,N_20621,N_20718);
nor U21166 (N_21166,N_20993,N_20783);
xor U21167 (N_21167,N_20508,N_20532);
nor U21168 (N_21168,N_20642,N_20915);
or U21169 (N_21169,N_20656,N_20981);
or U21170 (N_21170,N_20723,N_20633);
nand U21171 (N_21171,N_20797,N_20752);
or U21172 (N_21172,N_20547,N_20629);
and U21173 (N_21173,N_20670,N_20600);
nor U21174 (N_21174,N_20855,N_20735);
xor U21175 (N_21175,N_20738,N_20514);
or U21176 (N_21176,N_20893,N_20935);
or U21177 (N_21177,N_20800,N_20841);
nor U21178 (N_21178,N_20986,N_20890);
nand U21179 (N_21179,N_20839,N_20693);
or U21180 (N_21180,N_20527,N_20842);
nor U21181 (N_21181,N_20512,N_20943);
nor U21182 (N_21182,N_20764,N_20838);
or U21183 (N_21183,N_20891,N_20584);
or U21184 (N_21184,N_20885,N_20970);
or U21185 (N_21185,N_20557,N_20865);
or U21186 (N_21186,N_20878,N_20549);
or U21187 (N_21187,N_20907,N_20598);
nor U21188 (N_21188,N_20795,N_20912);
nand U21189 (N_21189,N_20609,N_20983);
and U21190 (N_21190,N_20950,N_20667);
and U21191 (N_21191,N_20711,N_20924);
nand U21192 (N_21192,N_20870,N_20770);
xor U21193 (N_21193,N_20704,N_20574);
and U21194 (N_21194,N_20682,N_20790);
nor U21195 (N_21195,N_20726,N_20979);
nand U21196 (N_21196,N_20582,N_20740);
nand U21197 (N_21197,N_20846,N_20985);
and U21198 (N_21198,N_20959,N_20545);
xnor U21199 (N_21199,N_20834,N_20782);
and U21200 (N_21200,N_20599,N_20648);
nor U21201 (N_21201,N_20666,N_20804);
nor U21202 (N_21202,N_20661,N_20739);
xor U21203 (N_21203,N_20815,N_20736);
or U21204 (N_21204,N_20857,N_20874);
or U21205 (N_21205,N_20517,N_20957);
nand U21206 (N_21206,N_20810,N_20698);
xor U21207 (N_21207,N_20753,N_20884);
nor U21208 (N_21208,N_20559,N_20867);
nand U21209 (N_21209,N_20699,N_20837);
xnor U21210 (N_21210,N_20510,N_20610);
xor U21211 (N_21211,N_20537,N_20905);
xor U21212 (N_21212,N_20663,N_20676);
nand U21213 (N_21213,N_20836,N_20733);
or U21214 (N_21214,N_20588,N_20630);
and U21215 (N_21215,N_20972,N_20760);
xor U21216 (N_21216,N_20713,N_20529);
nand U21217 (N_21217,N_20631,N_20681);
xor U21218 (N_21218,N_20696,N_20690);
nor U21219 (N_21219,N_20966,N_20938);
nand U21220 (N_21220,N_20961,N_20742);
or U21221 (N_21221,N_20833,N_20539);
nor U21222 (N_21222,N_20500,N_20930);
or U21223 (N_21223,N_20904,N_20788);
or U21224 (N_21224,N_20849,N_20775);
or U21225 (N_21225,N_20602,N_20931);
or U21226 (N_21226,N_20845,N_20937);
or U21227 (N_21227,N_20622,N_20789);
xor U21228 (N_21228,N_20614,N_20597);
nor U21229 (N_21229,N_20706,N_20958);
nand U21230 (N_21230,N_20798,N_20620);
or U21231 (N_21231,N_20601,N_20994);
nand U21232 (N_21232,N_20860,N_20585);
xor U21233 (N_21233,N_20636,N_20729);
xor U21234 (N_21234,N_20619,N_20637);
or U21235 (N_21235,N_20700,N_20659);
or U21236 (N_21236,N_20899,N_20794);
nor U21237 (N_21237,N_20671,N_20816);
xnor U21238 (N_21238,N_20605,N_20520);
and U21239 (N_21239,N_20746,N_20658);
nand U21240 (N_21240,N_20977,N_20992);
nand U21241 (N_21241,N_20672,N_20505);
and U21242 (N_21242,N_20933,N_20914);
or U21243 (N_21243,N_20632,N_20906);
nor U21244 (N_21244,N_20807,N_20806);
xor U21245 (N_21245,N_20546,N_20538);
nor U21246 (N_21246,N_20606,N_20553);
and U21247 (N_21247,N_20501,N_20534);
nand U21248 (N_21248,N_20556,N_20799);
and U21249 (N_21249,N_20554,N_20634);
and U21250 (N_21250,N_20881,N_20864);
nor U21251 (N_21251,N_20682,N_20958);
or U21252 (N_21252,N_20604,N_20790);
or U21253 (N_21253,N_20782,N_20669);
nor U21254 (N_21254,N_20580,N_20962);
nand U21255 (N_21255,N_20830,N_20965);
nor U21256 (N_21256,N_20810,N_20955);
xor U21257 (N_21257,N_20621,N_20855);
xnor U21258 (N_21258,N_20602,N_20518);
xnor U21259 (N_21259,N_20838,N_20699);
nor U21260 (N_21260,N_20546,N_20990);
nor U21261 (N_21261,N_20900,N_20531);
nand U21262 (N_21262,N_20636,N_20986);
or U21263 (N_21263,N_20764,N_20573);
xnor U21264 (N_21264,N_20903,N_20580);
nand U21265 (N_21265,N_20766,N_20725);
xor U21266 (N_21266,N_20621,N_20735);
and U21267 (N_21267,N_20975,N_20640);
nor U21268 (N_21268,N_20586,N_20544);
nor U21269 (N_21269,N_20569,N_20545);
or U21270 (N_21270,N_20677,N_20691);
and U21271 (N_21271,N_20682,N_20609);
nor U21272 (N_21272,N_20505,N_20857);
or U21273 (N_21273,N_20975,N_20859);
or U21274 (N_21274,N_20904,N_20638);
xor U21275 (N_21275,N_20879,N_20569);
or U21276 (N_21276,N_20921,N_20775);
nand U21277 (N_21277,N_20733,N_20770);
nand U21278 (N_21278,N_20905,N_20899);
or U21279 (N_21279,N_20868,N_20802);
nor U21280 (N_21280,N_20563,N_20964);
or U21281 (N_21281,N_20840,N_20638);
or U21282 (N_21282,N_20615,N_20947);
or U21283 (N_21283,N_20724,N_20644);
nand U21284 (N_21284,N_20514,N_20755);
or U21285 (N_21285,N_20899,N_20834);
xor U21286 (N_21286,N_20878,N_20731);
and U21287 (N_21287,N_20750,N_20822);
nor U21288 (N_21288,N_20734,N_20857);
and U21289 (N_21289,N_20627,N_20594);
xnor U21290 (N_21290,N_20606,N_20853);
xnor U21291 (N_21291,N_20889,N_20947);
xor U21292 (N_21292,N_20705,N_20693);
nand U21293 (N_21293,N_20684,N_20575);
xor U21294 (N_21294,N_20558,N_20735);
xor U21295 (N_21295,N_20836,N_20887);
nand U21296 (N_21296,N_20917,N_20752);
xnor U21297 (N_21297,N_20777,N_20604);
xnor U21298 (N_21298,N_20586,N_20742);
and U21299 (N_21299,N_20789,N_20668);
or U21300 (N_21300,N_20987,N_20529);
or U21301 (N_21301,N_20969,N_20520);
nor U21302 (N_21302,N_20501,N_20766);
nand U21303 (N_21303,N_20931,N_20558);
and U21304 (N_21304,N_20907,N_20708);
nor U21305 (N_21305,N_20698,N_20658);
nand U21306 (N_21306,N_20666,N_20654);
nor U21307 (N_21307,N_20788,N_20529);
or U21308 (N_21308,N_20692,N_20941);
and U21309 (N_21309,N_20674,N_20578);
and U21310 (N_21310,N_20627,N_20788);
xor U21311 (N_21311,N_20545,N_20589);
nand U21312 (N_21312,N_20978,N_20984);
xnor U21313 (N_21313,N_20984,N_20959);
nand U21314 (N_21314,N_20710,N_20803);
or U21315 (N_21315,N_20620,N_20705);
and U21316 (N_21316,N_20866,N_20898);
or U21317 (N_21317,N_20656,N_20805);
xnor U21318 (N_21318,N_20677,N_20865);
nand U21319 (N_21319,N_20909,N_20527);
or U21320 (N_21320,N_20660,N_20864);
and U21321 (N_21321,N_20532,N_20991);
and U21322 (N_21322,N_20670,N_20718);
nand U21323 (N_21323,N_20852,N_20900);
nor U21324 (N_21324,N_20746,N_20972);
and U21325 (N_21325,N_20542,N_20517);
nand U21326 (N_21326,N_20813,N_20506);
nor U21327 (N_21327,N_20909,N_20882);
nor U21328 (N_21328,N_20859,N_20791);
xor U21329 (N_21329,N_20719,N_20942);
nor U21330 (N_21330,N_20500,N_20596);
nand U21331 (N_21331,N_20939,N_20671);
nand U21332 (N_21332,N_20969,N_20528);
or U21333 (N_21333,N_20686,N_20665);
and U21334 (N_21334,N_20517,N_20919);
nand U21335 (N_21335,N_20860,N_20649);
nor U21336 (N_21336,N_20762,N_20703);
nor U21337 (N_21337,N_20957,N_20595);
or U21338 (N_21338,N_20688,N_20661);
xor U21339 (N_21339,N_20693,N_20658);
or U21340 (N_21340,N_20977,N_20536);
nor U21341 (N_21341,N_20709,N_20805);
xor U21342 (N_21342,N_20990,N_20837);
or U21343 (N_21343,N_20574,N_20971);
nor U21344 (N_21344,N_20745,N_20906);
and U21345 (N_21345,N_20874,N_20825);
and U21346 (N_21346,N_20758,N_20646);
nand U21347 (N_21347,N_20763,N_20675);
and U21348 (N_21348,N_20631,N_20694);
nor U21349 (N_21349,N_20557,N_20511);
nand U21350 (N_21350,N_20547,N_20638);
and U21351 (N_21351,N_20717,N_20820);
nor U21352 (N_21352,N_20531,N_20747);
nand U21353 (N_21353,N_20922,N_20726);
nor U21354 (N_21354,N_20731,N_20520);
nor U21355 (N_21355,N_20740,N_20528);
nand U21356 (N_21356,N_20635,N_20684);
nand U21357 (N_21357,N_20746,N_20906);
or U21358 (N_21358,N_20655,N_20810);
nor U21359 (N_21359,N_20844,N_20664);
or U21360 (N_21360,N_20734,N_20666);
nand U21361 (N_21361,N_20597,N_20541);
nand U21362 (N_21362,N_20603,N_20658);
and U21363 (N_21363,N_20766,N_20999);
xor U21364 (N_21364,N_20983,N_20611);
nand U21365 (N_21365,N_20820,N_20659);
nor U21366 (N_21366,N_20582,N_20965);
xor U21367 (N_21367,N_20612,N_20789);
nor U21368 (N_21368,N_20598,N_20638);
nor U21369 (N_21369,N_20582,N_20962);
nand U21370 (N_21370,N_20657,N_20665);
or U21371 (N_21371,N_20537,N_20788);
or U21372 (N_21372,N_20939,N_20797);
nor U21373 (N_21373,N_20532,N_20697);
or U21374 (N_21374,N_20538,N_20521);
nor U21375 (N_21375,N_20978,N_20682);
or U21376 (N_21376,N_20995,N_20699);
nor U21377 (N_21377,N_20866,N_20885);
or U21378 (N_21378,N_20732,N_20719);
nand U21379 (N_21379,N_20932,N_20921);
xor U21380 (N_21380,N_20815,N_20725);
nand U21381 (N_21381,N_20851,N_20776);
nand U21382 (N_21382,N_20700,N_20746);
nor U21383 (N_21383,N_20883,N_20567);
nor U21384 (N_21384,N_20961,N_20708);
or U21385 (N_21385,N_20622,N_20723);
nor U21386 (N_21386,N_20971,N_20983);
xnor U21387 (N_21387,N_20873,N_20521);
and U21388 (N_21388,N_20833,N_20873);
nand U21389 (N_21389,N_20996,N_20561);
nor U21390 (N_21390,N_20792,N_20500);
nor U21391 (N_21391,N_20714,N_20918);
nand U21392 (N_21392,N_20614,N_20876);
nor U21393 (N_21393,N_20681,N_20845);
xor U21394 (N_21394,N_20967,N_20531);
nand U21395 (N_21395,N_20664,N_20538);
nand U21396 (N_21396,N_20853,N_20552);
nor U21397 (N_21397,N_20594,N_20685);
nand U21398 (N_21398,N_20666,N_20561);
nand U21399 (N_21399,N_20886,N_20892);
nor U21400 (N_21400,N_20940,N_20827);
and U21401 (N_21401,N_20976,N_20953);
xor U21402 (N_21402,N_20612,N_20723);
nor U21403 (N_21403,N_20564,N_20707);
or U21404 (N_21404,N_20799,N_20900);
nor U21405 (N_21405,N_20967,N_20912);
nor U21406 (N_21406,N_20631,N_20620);
and U21407 (N_21407,N_20691,N_20679);
nor U21408 (N_21408,N_20597,N_20753);
or U21409 (N_21409,N_20922,N_20549);
nand U21410 (N_21410,N_20581,N_20632);
nand U21411 (N_21411,N_20714,N_20871);
or U21412 (N_21412,N_20910,N_20515);
or U21413 (N_21413,N_20665,N_20723);
and U21414 (N_21414,N_20556,N_20668);
or U21415 (N_21415,N_20896,N_20916);
nand U21416 (N_21416,N_20965,N_20539);
nor U21417 (N_21417,N_20913,N_20821);
or U21418 (N_21418,N_20839,N_20926);
or U21419 (N_21419,N_20585,N_20810);
xor U21420 (N_21420,N_20991,N_20957);
nand U21421 (N_21421,N_20644,N_20923);
nor U21422 (N_21422,N_20913,N_20903);
nand U21423 (N_21423,N_20684,N_20549);
nor U21424 (N_21424,N_20697,N_20879);
or U21425 (N_21425,N_20915,N_20938);
xnor U21426 (N_21426,N_20849,N_20687);
or U21427 (N_21427,N_20857,N_20751);
and U21428 (N_21428,N_20776,N_20723);
nor U21429 (N_21429,N_20904,N_20767);
nor U21430 (N_21430,N_20904,N_20553);
nand U21431 (N_21431,N_20906,N_20583);
xor U21432 (N_21432,N_20818,N_20658);
nand U21433 (N_21433,N_20807,N_20661);
nor U21434 (N_21434,N_20838,N_20984);
or U21435 (N_21435,N_20502,N_20992);
nand U21436 (N_21436,N_20888,N_20606);
and U21437 (N_21437,N_20900,N_20868);
and U21438 (N_21438,N_20606,N_20692);
or U21439 (N_21439,N_20724,N_20800);
xor U21440 (N_21440,N_20540,N_20978);
xnor U21441 (N_21441,N_20647,N_20764);
or U21442 (N_21442,N_20990,N_20805);
or U21443 (N_21443,N_20702,N_20917);
or U21444 (N_21444,N_20745,N_20628);
xnor U21445 (N_21445,N_20542,N_20834);
xnor U21446 (N_21446,N_20874,N_20606);
or U21447 (N_21447,N_20979,N_20544);
or U21448 (N_21448,N_20868,N_20977);
or U21449 (N_21449,N_20931,N_20546);
or U21450 (N_21450,N_20578,N_20992);
nor U21451 (N_21451,N_20876,N_20742);
xor U21452 (N_21452,N_20611,N_20951);
nor U21453 (N_21453,N_20577,N_20958);
xnor U21454 (N_21454,N_20925,N_20977);
or U21455 (N_21455,N_20985,N_20583);
and U21456 (N_21456,N_20645,N_20672);
or U21457 (N_21457,N_20785,N_20723);
nand U21458 (N_21458,N_20797,N_20695);
and U21459 (N_21459,N_20750,N_20833);
and U21460 (N_21460,N_20706,N_20586);
or U21461 (N_21461,N_20575,N_20864);
or U21462 (N_21462,N_20812,N_20545);
nor U21463 (N_21463,N_20614,N_20587);
and U21464 (N_21464,N_20749,N_20824);
xnor U21465 (N_21465,N_20625,N_20924);
xor U21466 (N_21466,N_20841,N_20805);
and U21467 (N_21467,N_20825,N_20763);
or U21468 (N_21468,N_20942,N_20527);
or U21469 (N_21469,N_20508,N_20760);
nor U21470 (N_21470,N_20851,N_20612);
or U21471 (N_21471,N_20945,N_20755);
or U21472 (N_21472,N_20891,N_20865);
nor U21473 (N_21473,N_20882,N_20942);
or U21474 (N_21474,N_20709,N_20771);
and U21475 (N_21475,N_20598,N_20686);
and U21476 (N_21476,N_20949,N_20813);
xnor U21477 (N_21477,N_20810,N_20799);
nor U21478 (N_21478,N_20730,N_20986);
xnor U21479 (N_21479,N_20603,N_20671);
or U21480 (N_21480,N_20636,N_20960);
xor U21481 (N_21481,N_20898,N_20957);
and U21482 (N_21482,N_20516,N_20555);
nor U21483 (N_21483,N_20993,N_20698);
and U21484 (N_21484,N_20797,N_20645);
nor U21485 (N_21485,N_20971,N_20703);
nand U21486 (N_21486,N_20656,N_20878);
nor U21487 (N_21487,N_20811,N_20669);
nor U21488 (N_21488,N_20980,N_20928);
xnor U21489 (N_21489,N_20990,N_20946);
or U21490 (N_21490,N_20902,N_20967);
xor U21491 (N_21491,N_20646,N_20512);
nor U21492 (N_21492,N_20927,N_20712);
xnor U21493 (N_21493,N_20517,N_20985);
or U21494 (N_21494,N_20831,N_20769);
nor U21495 (N_21495,N_20802,N_20737);
and U21496 (N_21496,N_20669,N_20807);
xor U21497 (N_21497,N_20649,N_20678);
xor U21498 (N_21498,N_20679,N_20948);
xnor U21499 (N_21499,N_20702,N_20586);
or U21500 (N_21500,N_21350,N_21469);
and U21501 (N_21501,N_21272,N_21089);
xor U21502 (N_21502,N_21387,N_21107);
nor U21503 (N_21503,N_21054,N_21266);
and U21504 (N_21504,N_21023,N_21396);
and U21505 (N_21505,N_21182,N_21376);
xor U21506 (N_21506,N_21132,N_21454);
nor U21507 (N_21507,N_21434,N_21496);
xor U21508 (N_21508,N_21220,N_21276);
or U21509 (N_21509,N_21101,N_21022);
nor U21510 (N_21510,N_21395,N_21018);
nand U21511 (N_21511,N_21056,N_21439);
or U21512 (N_21512,N_21058,N_21317);
and U21513 (N_21513,N_21455,N_21142);
nand U21514 (N_21514,N_21074,N_21229);
nand U21515 (N_21515,N_21131,N_21195);
and U21516 (N_21516,N_21051,N_21086);
and U21517 (N_21517,N_21192,N_21473);
and U21518 (N_21518,N_21451,N_21255);
nor U21519 (N_21519,N_21166,N_21232);
or U21520 (N_21520,N_21362,N_21053);
and U21521 (N_21521,N_21369,N_21010);
nor U21522 (N_21522,N_21334,N_21055);
nor U21523 (N_21523,N_21354,N_21287);
or U21524 (N_21524,N_21380,N_21288);
and U21525 (N_21525,N_21321,N_21363);
nor U21526 (N_21526,N_21459,N_21147);
and U21527 (N_21527,N_21412,N_21206);
and U21528 (N_21528,N_21249,N_21320);
xnor U21529 (N_21529,N_21092,N_21433);
nor U21530 (N_21530,N_21477,N_21224);
and U21531 (N_21531,N_21063,N_21417);
and U21532 (N_21532,N_21355,N_21031);
xor U21533 (N_21533,N_21444,N_21036);
xor U21534 (N_21534,N_21318,N_21271);
and U21535 (N_21535,N_21385,N_21401);
xnor U21536 (N_21536,N_21169,N_21392);
nand U21537 (N_21537,N_21083,N_21091);
nor U21538 (N_21538,N_21311,N_21157);
and U21539 (N_21539,N_21352,N_21331);
and U21540 (N_21540,N_21277,N_21114);
nand U21541 (N_21541,N_21274,N_21218);
xor U21542 (N_21542,N_21445,N_21360);
or U21543 (N_21543,N_21052,N_21134);
nand U21544 (N_21544,N_21047,N_21426);
nand U21545 (N_21545,N_21365,N_21170);
or U21546 (N_21546,N_21269,N_21012);
nor U21547 (N_21547,N_21216,N_21165);
nor U21548 (N_21548,N_21492,N_21208);
xnor U21549 (N_21549,N_21103,N_21239);
nand U21550 (N_21550,N_21286,N_21187);
and U21551 (N_21551,N_21210,N_21476);
or U21552 (N_21552,N_21094,N_21222);
nor U21553 (N_21553,N_21203,N_21160);
xnor U21554 (N_21554,N_21213,N_21389);
nor U21555 (N_21555,N_21440,N_21339);
nand U21556 (N_21556,N_21209,N_21338);
and U21557 (N_21557,N_21005,N_21375);
xor U21558 (N_21558,N_21357,N_21015);
xor U21559 (N_21559,N_21207,N_21489);
xnor U21560 (N_21560,N_21278,N_21102);
or U21561 (N_21561,N_21151,N_21144);
and U21562 (N_21562,N_21124,N_21240);
nor U21563 (N_21563,N_21198,N_21406);
nor U21564 (N_21564,N_21145,N_21066);
nor U21565 (N_21565,N_21322,N_21291);
or U21566 (N_21566,N_21499,N_21378);
and U21567 (N_21567,N_21487,N_21482);
and U21568 (N_21568,N_21327,N_21409);
nor U21569 (N_21569,N_21027,N_21028);
or U21570 (N_21570,N_21410,N_21494);
and U21571 (N_21571,N_21404,N_21221);
xor U21572 (N_21572,N_21405,N_21128);
and U21573 (N_21573,N_21133,N_21100);
nand U21574 (N_21574,N_21457,N_21326);
and U21575 (N_21575,N_21243,N_21423);
and U21576 (N_21576,N_21356,N_21470);
xnor U21577 (N_21577,N_21214,N_21143);
xnor U21578 (N_21578,N_21035,N_21425);
nor U21579 (N_21579,N_21468,N_21267);
nor U21580 (N_21580,N_21110,N_21155);
nand U21581 (N_21581,N_21138,N_21140);
or U21582 (N_21582,N_21186,N_21418);
xor U21583 (N_21583,N_21179,N_21244);
nand U21584 (N_21584,N_21148,N_21032);
nand U21585 (N_21585,N_21093,N_21167);
nor U21586 (N_21586,N_21087,N_21122);
or U21587 (N_21587,N_21004,N_21464);
or U21588 (N_21588,N_21310,N_21493);
nor U21589 (N_21589,N_21258,N_21259);
and U21590 (N_21590,N_21485,N_21163);
and U21591 (N_21591,N_21049,N_21264);
and U21592 (N_21592,N_21011,N_21319);
or U21593 (N_21593,N_21115,N_21307);
xor U21594 (N_21594,N_21484,N_21337);
and U21595 (N_21595,N_21466,N_21429);
and U21596 (N_21596,N_21064,N_21325);
nand U21597 (N_21597,N_21490,N_21449);
and U21598 (N_21598,N_21082,N_21105);
nand U21599 (N_21599,N_21297,N_21177);
xor U21600 (N_21600,N_21399,N_21181);
or U21601 (N_21601,N_21040,N_21121);
nor U21602 (N_21602,N_21296,N_21437);
or U21603 (N_21603,N_21290,N_21106);
and U21604 (N_21604,N_21193,N_21127);
or U21605 (N_21605,N_21479,N_21189);
nor U21606 (N_21606,N_21039,N_21137);
or U21607 (N_21607,N_21029,N_21231);
nor U21608 (N_21608,N_21046,N_21332);
xnor U21609 (N_21609,N_21480,N_21368);
xnor U21610 (N_21610,N_21026,N_21085);
xor U21611 (N_21611,N_21314,N_21384);
or U21612 (N_21612,N_21359,N_21374);
xor U21613 (N_21613,N_21430,N_21071);
nand U21614 (N_21614,N_21045,N_21097);
and U21615 (N_21615,N_21235,N_21308);
xnor U21616 (N_21616,N_21201,N_21377);
or U21617 (N_21617,N_21498,N_21261);
nand U21618 (N_21618,N_21042,N_21164);
nand U21619 (N_21619,N_21407,N_21371);
or U21620 (N_21620,N_21293,N_21073);
xor U21621 (N_21621,N_21495,N_21335);
nand U21622 (N_21622,N_21370,N_21302);
xnor U21623 (N_21623,N_21003,N_21057);
xnor U21624 (N_21624,N_21388,N_21347);
or U21625 (N_21625,N_21095,N_21041);
nor U21626 (N_21626,N_21014,N_21372);
xor U21627 (N_21627,N_21353,N_21006);
or U21628 (N_21628,N_21292,N_21162);
xnor U21629 (N_21629,N_21265,N_21149);
xor U21630 (N_21630,N_21394,N_21204);
and U21631 (N_21631,N_21402,N_21116);
xnor U21632 (N_21632,N_21438,N_21060);
xnor U21633 (N_21633,N_21098,N_21223);
nor U21634 (N_21634,N_21460,N_21129);
or U21635 (N_21635,N_21176,N_21393);
nand U21636 (N_21636,N_21323,N_21196);
xnor U21637 (N_21637,N_21070,N_21159);
or U21638 (N_21638,N_21458,N_21270);
xor U21639 (N_21639,N_21242,N_21237);
or U21640 (N_21640,N_21475,N_21191);
and U21641 (N_21641,N_21034,N_21397);
xnor U21642 (N_21642,N_21481,N_21108);
or U21643 (N_21643,N_21130,N_21065);
nand U21644 (N_21644,N_21497,N_21431);
or U21645 (N_21645,N_21309,N_21341);
and U21646 (N_21646,N_21299,N_21076);
xnor U21647 (N_21647,N_21456,N_21488);
or U21648 (N_21648,N_21281,N_21180);
and U21649 (N_21649,N_21183,N_21421);
nor U21650 (N_21650,N_21398,N_21135);
xnor U21651 (N_21651,N_21025,N_21062);
and U21652 (N_21652,N_21117,N_21283);
xnor U21653 (N_21653,N_21263,N_21465);
xnor U21654 (N_21654,N_21452,N_21215);
nand U21655 (N_21655,N_21119,N_21079);
xnor U21656 (N_21656,N_21342,N_21205);
and U21657 (N_21657,N_21125,N_21017);
nor U21658 (N_21658,N_21351,N_21268);
nand U21659 (N_21659,N_21247,N_21059);
nor U21660 (N_21660,N_21348,N_21386);
and U21661 (N_21661,N_21383,N_21020);
or U21662 (N_21662,N_21251,N_21413);
nand U21663 (N_21663,N_21037,N_21178);
or U21664 (N_21664,N_21194,N_21099);
xor U21665 (N_21665,N_21254,N_21432);
nand U21666 (N_21666,N_21419,N_21185);
and U21667 (N_21667,N_21345,N_21217);
nand U21668 (N_21668,N_21379,N_21013);
or U21669 (N_21669,N_21346,N_21048);
nor U21670 (N_21670,N_21226,N_21021);
or U21671 (N_21671,N_21228,N_21126);
or U21672 (N_21672,N_21343,N_21315);
nand U21673 (N_21673,N_21202,N_21390);
nor U21674 (N_21674,N_21068,N_21486);
and U21675 (N_21675,N_21289,N_21118);
and U21676 (N_21676,N_21078,N_21447);
nand U21677 (N_21677,N_21442,N_21088);
nor U21678 (N_21678,N_21403,N_21256);
xor U21679 (N_21679,N_21472,N_21260);
nand U21680 (N_21680,N_21330,N_21096);
nand U21681 (N_21681,N_21483,N_21146);
or U21682 (N_21682,N_21415,N_21435);
and U21683 (N_21683,N_21227,N_21411);
or U21684 (N_21684,N_21467,N_21211);
nand U21685 (N_21685,N_21112,N_21414);
xor U21686 (N_21686,N_21427,N_21312);
and U21687 (N_21687,N_21241,N_21295);
and U21688 (N_21688,N_21174,N_21252);
nand U21689 (N_21689,N_21367,N_21188);
nand U21690 (N_21690,N_21038,N_21253);
nand U21691 (N_21691,N_21024,N_21084);
and U21692 (N_21692,N_21190,N_21453);
nor U21693 (N_21693,N_21236,N_21285);
and U21694 (N_21694,N_21349,N_21450);
and U21695 (N_21695,N_21043,N_21333);
nor U21696 (N_21696,N_21184,N_21111);
nor U21697 (N_21697,N_21009,N_21303);
nand U21698 (N_21698,N_21158,N_21382);
and U21699 (N_21699,N_21422,N_21200);
and U21700 (N_21700,N_21069,N_21007);
or U21701 (N_21701,N_21171,N_21462);
nand U21702 (N_21702,N_21080,N_21300);
nand U21703 (N_21703,N_21219,N_21361);
and U21704 (N_21704,N_21441,N_21197);
nor U21705 (N_21705,N_21001,N_21446);
nor U21706 (N_21706,N_21400,N_21336);
or U21707 (N_21707,N_21324,N_21298);
nand U21708 (N_21708,N_21340,N_21358);
and U21709 (N_21709,N_21316,N_21420);
xor U21710 (N_21710,N_21152,N_21233);
and U21711 (N_21711,N_21245,N_21067);
nor U21712 (N_21712,N_21275,N_21478);
and U21713 (N_21713,N_21424,N_21123);
nand U21714 (N_21714,N_21373,N_21120);
nand U21715 (N_21715,N_21175,N_21168);
and U21716 (N_21716,N_21257,N_21075);
nand U21717 (N_21717,N_21461,N_21282);
xor U21718 (N_21718,N_21008,N_21161);
and U21719 (N_21719,N_21284,N_21474);
nand U21720 (N_21720,N_21153,N_21016);
xor U21721 (N_21721,N_21280,N_21173);
nand U21722 (N_21722,N_21491,N_21225);
and U21723 (N_21723,N_21156,N_21033);
and U21724 (N_21724,N_21436,N_21081);
and U21725 (N_21725,N_21328,N_21408);
xnor U21726 (N_21726,N_21381,N_21002);
or U21727 (N_21727,N_21443,N_21136);
nor U21728 (N_21728,N_21113,N_21154);
or U21729 (N_21729,N_21305,N_21273);
nand U21730 (N_21730,N_21077,N_21250);
and U21731 (N_21731,N_21030,N_21061);
nand U21732 (N_21732,N_21448,N_21246);
and U21733 (N_21733,N_21019,N_21344);
nand U21734 (N_21734,N_21044,N_21416);
and U21735 (N_21735,N_21139,N_21090);
nand U21736 (N_21736,N_21391,N_21301);
nor U21737 (N_21737,N_21248,N_21364);
nor U21738 (N_21738,N_21262,N_21234);
xor U21739 (N_21739,N_21306,N_21050);
nand U21740 (N_21740,N_21471,N_21428);
nor U21741 (N_21741,N_21463,N_21199);
or U21742 (N_21742,N_21172,N_21366);
nor U21743 (N_21743,N_21279,N_21230);
nand U21744 (N_21744,N_21212,N_21104);
or U21745 (N_21745,N_21141,N_21072);
nor U21746 (N_21746,N_21238,N_21329);
and U21747 (N_21747,N_21313,N_21150);
nor U21748 (N_21748,N_21304,N_21000);
xnor U21749 (N_21749,N_21294,N_21109);
nor U21750 (N_21750,N_21446,N_21088);
nand U21751 (N_21751,N_21047,N_21479);
xor U21752 (N_21752,N_21380,N_21200);
or U21753 (N_21753,N_21179,N_21082);
nand U21754 (N_21754,N_21278,N_21483);
nand U21755 (N_21755,N_21430,N_21078);
nor U21756 (N_21756,N_21138,N_21444);
or U21757 (N_21757,N_21279,N_21201);
or U21758 (N_21758,N_21328,N_21039);
nand U21759 (N_21759,N_21035,N_21305);
nand U21760 (N_21760,N_21423,N_21316);
and U21761 (N_21761,N_21256,N_21347);
and U21762 (N_21762,N_21137,N_21421);
xor U21763 (N_21763,N_21092,N_21387);
nor U21764 (N_21764,N_21321,N_21349);
and U21765 (N_21765,N_21401,N_21428);
nor U21766 (N_21766,N_21017,N_21357);
nand U21767 (N_21767,N_21245,N_21008);
or U21768 (N_21768,N_21070,N_21447);
and U21769 (N_21769,N_21377,N_21441);
nor U21770 (N_21770,N_21446,N_21023);
nor U21771 (N_21771,N_21161,N_21345);
or U21772 (N_21772,N_21482,N_21201);
and U21773 (N_21773,N_21024,N_21082);
nand U21774 (N_21774,N_21195,N_21281);
and U21775 (N_21775,N_21268,N_21238);
nand U21776 (N_21776,N_21450,N_21113);
or U21777 (N_21777,N_21287,N_21027);
xor U21778 (N_21778,N_21357,N_21297);
and U21779 (N_21779,N_21248,N_21098);
nor U21780 (N_21780,N_21371,N_21040);
nor U21781 (N_21781,N_21459,N_21332);
and U21782 (N_21782,N_21461,N_21137);
and U21783 (N_21783,N_21368,N_21148);
nor U21784 (N_21784,N_21078,N_21468);
nand U21785 (N_21785,N_21200,N_21092);
or U21786 (N_21786,N_21310,N_21385);
nor U21787 (N_21787,N_21085,N_21285);
and U21788 (N_21788,N_21134,N_21467);
or U21789 (N_21789,N_21499,N_21040);
nand U21790 (N_21790,N_21106,N_21402);
or U21791 (N_21791,N_21131,N_21025);
or U21792 (N_21792,N_21220,N_21427);
xor U21793 (N_21793,N_21288,N_21454);
nor U21794 (N_21794,N_21140,N_21063);
nor U21795 (N_21795,N_21329,N_21197);
or U21796 (N_21796,N_21112,N_21317);
and U21797 (N_21797,N_21491,N_21335);
nand U21798 (N_21798,N_21338,N_21281);
nor U21799 (N_21799,N_21156,N_21184);
nor U21800 (N_21800,N_21492,N_21341);
nor U21801 (N_21801,N_21444,N_21061);
or U21802 (N_21802,N_21407,N_21047);
nand U21803 (N_21803,N_21160,N_21007);
nor U21804 (N_21804,N_21051,N_21204);
and U21805 (N_21805,N_21277,N_21412);
nor U21806 (N_21806,N_21151,N_21438);
and U21807 (N_21807,N_21477,N_21274);
nor U21808 (N_21808,N_21305,N_21429);
or U21809 (N_21809,N_21073,N_21143);
or U21810 (N_21810,N_21266,N_21008);
xnor U21811 (N_21811,N_21405,N_21199);
or U21812 (N_21812,N_21076,N_21111);
or U21813 (N_21813,N_21071,N_21136);
or U21814 (N_21814,N_21088,N_21341);
or U21815 (N_21815,N_21079,N_21205);
nand U21816 (N_21816,N_21434,N_21349);
xor U21817 (N_21817,N_21073,N_21154);
nand U21818 (N_21818,N_21210,N_21247);
and U21819 (N_21819,N_21374,N_21137);
nand U21820 (N_21820,N_21311,N_21244);
xor U21821 (N_21821,N_21476,N_21322);
xnor U21822 (N_21822,N_21248,N_21232);
nand U21823 (N_21823,N_21306,N_21008);
nand U21824 (N_21824,N_21063,N_21124);
or U21825 (N_21825,N_21116,N_21162);
or U21826 (N_21826,N_21478,N_21302);
nand U21827 (N_21827,N_21469,N_21152);
xnor U21828 (N_21828,N_21063,N_21413);
xnor U21829 (N_21829,N_21148,N_21496);
and U21830 (N_21830,N_21093,N_21476);
or U21831 (N_21831,N_21231,N_21222);
nand U21832 (N_21832,N_21324,N_21169);
or U21833 (N_21833,N_21261,N_21238);
or U21834 (N_21834,N_21157,N_21326);
xnor U21835 (N_21835,N_21287,N_21280);
xnor U21836 (N_21836,N_21269,N_21286);
and U21837 (N_21837,N_21072,N_21413);
xor U21838 (N_21838,N_21109,N_21439);
and U21839 (N_21839,N_21147,N_21029);
and U21840 (N_21840,N_21423,N_21057);
nor U21841 (N_21841,N_21233,N_21011);
or U21842 (N_21842,N_21316,N_21233);
nand U21843 (N_21843,N_21491,N_21216);
nor U21844 (N_21844,N_21063,N_21471);
and U21845 (N_21845,N_21465,N_21456);
or U21846 (N_21846,N_21042,N_21312);
or U21847 (N_21847,N_21324,N_21253);
xor U21848 (N_21848,N_21291,N_21455);
nor U21849 (N_21849,N_21185,N_21065);
or U21850 (N_21850,N_21105,N_21430);
nand U21851 (N_21851,N_21381,N_21251);
nand U21852 (N_21852,N_21371,N_21257);
or U21853 (N_21853,N_21227,N_21474);
nand U21854 (N_21854,N_21202,N_21224);
and U21855 (N_21855,N_21009,N_21048);
nor U21856 (N_21856,N_21014,N_21191);
or U21857 (N_21857,N_21323,N_21260);
and U21858 (N_21858,N_21403,N_21467);
xnor U21859 (N_21859,N_21206,N_21170);
nor U21860 (N_21860,N_21245,N_21364);
nand U21861 (N_21861,N_21490,N_21380);
nor U21862 (N_21862,N_21121,N_21460);
nor U21863 (N_21863,N_21023,N_21146);
or U21864 (N_21864,N_21009,N_21163);
nor U21865 (N_21865,N_21495,N_21232);
and U21866 (N_21866,N_21158,N_21460);
xor U21867 (N_21867,N_21443,N_21177);
xor U21868 (N_21868,N_21146,N_21039);
nor U21869 (N_21869,N_21131,N_21074);
nor U21870 (N_21870,N_21253,N_21146);
xor U21871 (N_21871,N_21217,N_21306);
or U21872 (N_21872,N_21189,N_21394);
nor U21873 (N_21873,N_21447,N_21223);
or U21874 (N_21874,N_21031,N_21425);
nand U21875 (N_21875,N_21469,N_21478);
nor U21876 (N_21876,N_21202,N_21388);
nor U21877 (N_21877,N_21243,N_21076);
or U21878 (N_21878,N_21228,N_21265);
xnor U21879 (N_21879,N_21322,N_21191);
nor U21880 (N_21880,N_21427,N_21171);
or U21881 (N_21881,N_21340,N_21332);
and U21882 (N_21882,N_21107,N_21094);
nor U21883 (N_21883,N_21483,N_21202);
xor U21884 (N_21884,N_21298,N_21432);
xnor U21885 (N_21885,N_21492,N_21226);
or U21886 (N_21886,N_21085,N_21209);
nor U21887 (N_21887,N_21340,N_21405);
and U21888 (N_21888,N_21169,N_21311);
or U21889 (N_21889,N_21252,N_21308);
nand U21890 (N_21890,N_21213,N_21305);
nor U21891 (N_21891,N_21198,N_21061);
nor U21892 (N_21892,N_21346,N_21088);
nand U21893 (N_21893,N_21038,N_21313);
and U21894 (N_21894,N_21444,N_21083);
and U21895 (N_21895,N_21290,N_21257);
and U21896 (N_21896,N_21454,N_21266);
or U21897 (N_21897,N_21114,N_21000);
nor U21898 (N_21898,N_21170,N_21131);
nor U21899 (N_21899,N_21325,N_21226);
nand U21900 (N_21900,N_21308,N_21364);
nor U21901 (N_21901,N_21149,N_21045);
or U21902 (N_21902,N_21159,N_21001);
xor U21903 (N_21903,N_21381,N_21331);
and U21904 (N_21904,N_21127,N_21368);
nand U21905 (N_21905,N_21399,N_21077);
nor U21906 (N_21906,N_21106,N_21107);
or U21907 (N_21907,N_21498,N_21187);
and U21908 (N_21908,N_21106,N_21345);
or U21909 (N_21909,N_21301,N_21298);
nand U21910 (N_21910,N_21067,N_21427);
xnor U21911 (N_21911,N_21384,N_21298);
or U21912 (N_21912,N_21262,N_21350);
or U21913 (N_21913,N_21423,N_21245);
nor U21914 (N_21914,N_21431,N_21379);
nor U21915 (N_21915,N_21020,N_21165);
or U21916 (N_21916,N_21167,N_21289);
xnor U21917 (N_21917,N_21410,N_21038);
and U21918 (N_21918,N_21362,N_21218);
and U21919 (N_21919,N_21069,N_21163);
xor U21920 (N_21920,N_21156,N_21475);
nor U21921 (N_21921,N_21084,N_21126);
nand U21922 (N_21922,N_21441,N_21153);
xor U21923 (N_21923,N_21069,N_21061);
xor U21924 (N_21924,N_21004,N_21102);
xnor U21925 (N_21925,N_21393,N_21069);
nand U21926 (N_21926,N_21073,N_21254);
and U21927 (N_21927,N_21406,N_21167);
xnor U21928 (N_21928,N_21019,N_21169);
nor U21929 (N_21929,N_21478,N_21067);
or U21930 (N_21930,N_21034,N_21420);
nor U21931 (N_21931,N_21295,N_21347);
and U21932 (N_21932,N_21063,N_21265);
xor U21933 (N_21933,N_21272,N_21156);
nor U21934 (N_21934,N_21241,N_21360);
nand U21935 (N_21935,N_21104,N_21351);
nor U21936 (N_21936,N_21475,N_21299);
nand U21937 (N_21937,N_21423,N_21119);
xor U21938 (N_21938,N_21261,N_21496);
nor U21939 (N_21939,N_21438,N_21441);
and U21940 (N_21940,N_21045,N_21361);
xor U21941 (N_21941,N_21275,N_21361);
nor U21942 (N_21942,N_21328,N_21124);
nand U21943 (N_21943,N_21203,N_21270);
nor U21944 (N_21944,N_21367,N_21109);
xnor U21945 (N_21945,N_21280,N_21035);
nor U21946 (N_21946,N_21167,N_21284);
xor U21947 (N_21947,N_21280,N_21027);
nand U21948 (N_21948,N_21299,N_21208);
nor U21949 (N_21949,N_21070,N_21235);
and U21950 (N_21950,N_21048,N_21412);
and U21951 (N_21951,N_21128,N_21191);
and U21952 (N_21952,N_21437,N_21471);
and U21953 (N_21953,N_21113,N_21221);
nand U21954 (N_21954,N_21420,N_21196);
or U21955 (N_21955,N_21141,N_21279);
xor U21956 (N_21956,N_21108,N_21473);
nand U21957 (N_21957,N_21025,N_21350);
nor U21958 (N_21958,N_21396,N_21382);
nor U21959 (N_21959,N_21207,N_21335);
and U21960 (N_21960,N_21003,N_21341);
xor U21961 (N_21961,N_21164,N_21079);
xnor U21962 (N_21962,N_21205,N_21276);
xnor U21963 (N_21963,N_21439,N_21287);
nand U21964 (N_21964,N_21046,N_21274);
nand U21965 (N_21965,N_21301,N_21225);
xor U21966 (N_21966,N_21315,N_21009);
and U21967 (N_21967,N_21118,N_21023);
and U21968 (N_21968,N_21356,N_21101);
or U21969 (N_21969,N_21458,N_21238);
nor U21970 (N_21970,N_21108,N_21276);
xnor U21971 (N_21971,N_21247,N_21180);
and U21972 (N_21972,N_21327,N_21492);
and U21973 (N_21973,N_21230,N_21473);
xnor U21974 (N_21974,N_21414,N_21256);
nand U21975 (N_21975,N_21004,N_21449);
and U21976 (N_21976,N_21056,N_21318);
nand U21977 (N_21977,N_21141,N_21263);
nor U21978 (N_21978,N_21092,N_21145);
xor U21979 (N_21979,N_21172,N_21050);
nor U21980 (N_21980,N_21239,N_21295);
nor U21981 (N_21981,N_21107,N_21144);
nor U21982 (N_21982,N_21369,N_21098);
and U21983 (N_21983,N_21160,N_21190);
or U21984 (N_21984,N_21430,N_21183);
nand U21985 (N_21985,N_21263,N_21072);
nand U21986 (N_21986,N_21376,N_21381);
nor U21987 (N_21987,N_21327,N_21349);
nor U21988 (N_21988,N_21234,N_21191);
nor U21989 (N_21989,N_21176,N_21395);
nor U21990 (N_21990,N_21226,N_21057);
nor U21991 (N_21991,N_21148,N_21116);
nand U21992 (N_21992,N_21017,N_21069);
or U21993 (N_21993,N_21161,N_21473);
or U21994 (N_21994,N_21473,N_21030);
nand U21995 (N_21995,N_21157,N_21148);
nand U21996 (N_21996,N_21029,N_21461);
nand U21997 (N_21997,N_21013,N_21435);
xor U21998 (N_21998,N_21369,N_21494);
and U21999 (N_21999,N_21493,N_21366);
and U22000 (N_22000,N_21918,N_21572);
nor U22001 (N_22001,N_21672,N_21798);
or U22002 (N_22002,N_21971,N_21737);
xnor U22003 (N_22003,N_21696,N_21986);
and U22004 (N_22004,N_21608,N_21771);
or U22005 (N_22005,N_21834,N_21704);
or U22006 (N_22006,N_21648,N_21613);
xor U22007 (N_22007,N_21679,N_21831);
or U22008 (N_22008,N_21855,N_21970);
or U22009 (N_22009,N_21732,N_21892);
nand U22010 (N_22010,N_21684,N_21615);
xnor U22011 (N_22011,N_21954,N_21898);
or U22012 (N_22012,N_21962,N_21693);
nand U22013 (N_22013,N_21724,N_21899);
nor U22014 (N_22014,N_21797,N_21826);
or U22015 (N_22015,N_21707,N_21754);
and U22016 (N_22016,N_21645,N_21744);
and U22017 (N_22017,N_21625,N_21966);
nand U22018 (N_22018,N_21669,N_21836);
nor U22019 (N_22019,N_21505,N_21759);
xnor U22020 (N_22020,N_21775,N_21843);
or U22021 (N_22021,N_21832,N_21916);
or U22022 (N_22022,N_21589,N_21752);
xor U22023 (N_22023,N_21884,N_21886);
and U22024 (N_22024,N_21622,N_21805);
and U22025 (N_22025,N_21793,N_21766);
nor U22026 (N_22026,N_21659,N_21717);
or U22027 (N_22027,N_21537,N_21506);
and U22028 (N_22028,N_21840,N_21879);
or U22029 (N_22029,N_21746,N_21644);
xnor U22030 (N_22030,N_21747,N_21510);
xor U22031 (N_22031,N_21927,N_21567);
and U22032 (N_22032,N_21583,N_21887);
nor U22033 (N_22033,N_21846,N_21847);
nand U22034 (N_22034,N_21690,N_21849);
nand U22035 (N_22035,N_21786,N_21687);
or U22036 (N_22036,N_21921,N_21607);
or U22037 (N_22037,N_21726,N_21545);
xnor U22038 (N_22038,N_21864,N_21725);
or U22039 (N_22039,N_21518,N_21663);
nor U22040 (N_22040,N_21995,N_21857);
or U22041 (N_22041,N_21770,N_21783);
xnor U22042 (N_22042,N_21817,N_21689);
nor U22043 (N_22043,N_21616,N_21891);
and U22044 (N_22044,N_21603,N_21982);
nand U22045 (N_22045,N_21941,N_21757);
and U22046 (N_22046,N_21636,N_21959);
xor U22047 (N_22047,N_21915,N_21623);
xnor U22048 (N_22048,N_21552,N_21697);
nand U22049 (N_22049,N_21952,N_21527);
or U22050 (N_22050,N_21781,N_21534);
xnor U22051 (N_22051,N_21674,N_21595);
nor U22052 (N_22052,N_21610,N_21548);
xor U22053 (N_22053,N_21845,N_21994);
xnor U22054 (N_22054,N_21525,N_21833);
xor U22055 (N_22055,N_21889,N_21722);
or U22056 (N_22056,N_21656,N_21714);
and U22057 (N_22057,N_21695,N_21815);
nor U22058 (N_22058,N_21897,N_21516);
nor U22059 (N_22059,N_21773,N_21555);
and U22060 (N_22060,N_21984,N_21960);
nand U22061 (N_22061,N_21677,N_21578);
or U22062 (N_22062,N_21540,N_21713);
nand U22063 (N_22063,N_21675,N_21647);
nor U22064 (N_22064,N_21967,N_21803);
nor U22065 (N_22065,N_21838,N_21626);
and U22066 (N_22066,N_21908,N_21926);
nand U22067 (N_22067,N_21730,N_21627);
nor U22068 (N_22068,N_21900,N_21731);
xnor U22069 (N_22069,N_21600,N_21522);
xnor U22070 (N_22070,N_21762,N_21706);
nor U22071 (N_22071,N_21923,N_21652);
nor U22072 (N_22072,N_21575,N_21500);
xor U22073 (N_22073,N_21646,N_21951);
nor U22074 (N_22074,N_21563,N_21564);
nand U22075 (N_22075,N_21619,N_21877);
xor U22076 (N_22076,N_21523,N_21880);
or U22077 (N_22077,N_21816,N_21728);
or U22078 (N_22078,N_21894,N_21520);
xor U22079 (N_22079,N_21676,N_21742);
xnor U22080 (N_22080,N_21776,N_21761);
nor U22081 (N_22081,N_21878,N_21691);
or U22082 (N_22082,N_21807,N_21528);
xnor U22083 (N_22083,N_21765,N_21686);
nor U22084 (N_22084,N_21968,N_21869);
and U22085 (N_22085,N_21565,N_21931);
and U22086 (N_22086,N_21907,N_21733);
or U22087 (N_22087,N_21748,N_21649);
and U22088 (N_22088,N_21692,N_21678);
and U22089 (N_22089,N_21827,N_21810);
nand U22090 (N_22090,N_21683,N_21862);
nand U22091 (N_22091,N_21597,N_21939);
or U22092 (N_22092,N_21541,N_21774);
nand U22093 (N_22093,N_21670,N_21850);
and U22094 (N_22094,N_21870,N_21633);
nand U22095 (N_22095,N_21550,N_21976);
nor U22096 (N_22096,N_21573,N_21949);
and U22097 (N_22097,N_21930,N_21789);
and U22098 (N_22098,N_21716,N_21584);
xnor U22099 (N_22099,N_21688,N_21859);
xnor U22100 (N_22100,N_21632,N_21602);
xnor U22101 (N_22101,N_21612,N_21991);
or U22102 (N_22102,N_21576,N_21779);
and U22103 (N_22103,N_21953,N_21928);
xor U22104 (N_22104,N_21574,N_21957);
or U22105 (N_22105,N_21769,N_21973);
and U22106 (N_22106,N_21539,N_21721);
and U22107 (N_22107,N_21943,N_21557);
or U22108 (N_22108,N_21710,N_21547);
nand U22109 (N_22109,N_21658,N_21503);
or U22110 (N_22110,N_21938,N_21609);
and U22111 (N_22111,N_21950,N_21784);
or U22112 (N_22112,N_21796,N_21822);
nand U22113 (N_22113,N_21996,N_21972);
or U22114 (N_22114,N_21740,N_21620);
or U22115 (N_22115,N_21738,N_21910);
or U22116 (N_22116,N_21749,N_21806);
or U22117 (N_22117,N_21685,N_21919);
and U22118 (N_22118,N_21579,N_21587);
xor U22119 (N_22119,N_21912,N_21768);
and U22120 (N_22120,N_21700,N_21566);
or U22121 (N_22121,N_21666,N_21662);
xor U22122 (N_22122,N_21665,N_21818);
or U22123 (N_22123,N_21830,N_21979);
nor U22124 (N_22124,N_21533,N_21514);
and U22125 (N_22125,N_21544,N_21756);
nand U22126 (N_22126,N_21913,N_21551);
or U22127 (N_22127,N_21785,N_21708);
xnor U22128 (N_22128,N_21961,N_21825);
or U22129 (N_22129,N_21881,N_21509);
and U22130 (N_22130,N_21529,N_21701);
or U22131 (N_22131,N_21535,N_21532);
nor U22132 (N_22132,N_21654,N_21592);
or U22133 (N_22133,N_21999,N_21624);
xnor U22134 (N_22134,N_21974,N_21702);
xor U22135 (N_22135,N_21611,N_21804);
nor U22136 (N_22136,N_21842,N_21703);
nor U22137 (N_22137,N_21824,N_21723);
or U22138 (N_22138,N_21504,N_21837);
xor U22139 (N_22139,N_21628,N_21718);
or U22140 (N_22140,N_21865,N_21852);
and U22141 (N_22141,N_21591,N_21874);
nor U22142 (N_22142,N_21811,N_21987);
nand U22143 (N_22143,N_21641,N_21945);
and U22144 (N_22144,N_21629,N_21614);
nand U22145 (N_22145,N_21667,N_21820);
xnor U22146 (N_22146,N_21856,N_21809);
or U22147 (N_22147,N_21604,N_21858);
or U22148 (N_22148,N_21990,N_21942);
and U22149 (N_22149,N_21712,N_21515);
or U22150 (N_22150,N_21998,N_21782);
or U22151 (N_22151,N_21988,N_21517);
xnor U22152 (N_22152,N_21637,N_21935);
and U22153 (N_22153,N_21876,N_21882);
nor U22154 (N_22154,N_21904,N_21888);
and U22155 (N_22155,N_21598,N_21905);
xnor U22156 (N_22156,N_21875,N_21531);
or U22157 (N_22157,N_21940,N_21720);
nand U22158 (N_22158,N_21585,N_21705);
xnor U22159 (N_22159,N_21507,N_21790);
xnor U22160 (N_22160,N_21751,N_21735);
or U22161 (N_22161,N_21958,N_21743);
xnor U22162 (N_22162,N_21902,N_21868);
nand U22163 (N_22163,N_21699,N_21835);
or U22164 (N_22164,N_21668,N_21823);
or U22165 (N_22165,N_21556,N_21767);
nor U22166 (N_22166,N_21821,N_21588);
nor U22167 (N_22167,N_21872,N_21828);
or U22168 (N_22168,N_21562,N_21777);
and U22169 (N_22169,N_21634,N_21521);
nor U22170 (N_22170,N_21524,N_21911);
nor U22171 (N_22171,N_21933,N_21946);
and U22172 (N_22172,N_21922,N_21863);
or U22173 (N_22173,N_21975,N_21594);
and U22174 (N_22174,N_21841,N_21772);
xor U22175 (N_22175,N_21630,N_21727);
xnor U22176 (N_22176,N_21596,N_21558);
nor U22177 (N_22177,N_21794,N_21739);
or U22178 (N_22178,N_21501,N_21801);
and U22179 (N_22179,N_21920,N_21640);
and U22180 (N_22180,N_21839,N_21778);
or U22181 (N_22181,N_21764,N_21681);
and U22182 (N_22182,N_21680,N_21788);
and U22183 (N_22183,N_21711,N_21799);
or U22184 (N_22184,N_21929,N_21980);
or U22185 (N_22185,N_21906,N_21792);
nor U22186 (N_22186,N_21639,N_21715);
nor U22187 (N_22187,N_21992,N_21601);
nor U22188 (N_22188,N_21808,N_21851);
and U22189 (N_22189,N_21568,N_21653);
nand U22190 (N_22190,N_21914,N_21925);
or U22191 (N_22191,N_21526,N_21917);
nand U22192 (N_22192,N_21755,N_21736);
and U22193 (N_22193,N_21924,N_21854);
or U22194 (N_22194,N_21553,N_21955);
or U22195 (N_22195,N_21895,N_21885);
nand U22196 (N_22196,N_21513,N_21848);
nand U22197 (N_22197,N_21661,N_21989);
xor U22198 (N_22198,N_21763,N_21618);
and U22199 (N_22199,N_21549,N_21944);
and U22200 (N_22200,N_21964,N_21536);
nor U22201 (N_22201,N_21936,N_21621);
or U22202 (N_22202,N_21519,N_21948);
nor U22203 (N_22203,N_21969,N_21580);
xnor U22204 (N_22204,N_21590,N_21978);
xnor U22205 (N_22205,N_21750,N_21932);
or U22206 (N_22206,N_21617,N_21934);
and U22207 (N_22207,N_21963,N_21682);
or U22208 (N_22208,N_21593,N_21791);
nor U22209 (N_22209,N_21511,N_21734);
and U22210 (N_22210,N_21543,N_21651);
nand U22211 (N_22211,N_21673,N_21909);
and U22212 (N_22212,N_21586,N_21508);
and U22213 (N_22213,N_21698,N_21861);
xnor U22214 (N_22214,N_21577,N_21570);
or U22215 (N_22215,N_21997,N_21582);
xor U22216 (N_22216,N_21502,N_21903);
nor U22217 (N_22217,N_21829,N_21729);
nand U22218 (N_22218,N_21977,N_21694);
xor U22219 (N_22219,N_21802,N_21635);
xor U22220 (N_22220,N_21871,N_21813);
or U22221 (N_22221,N_21780,N_21800);
nand U22222 (N_22222,N_21671,N_21819);
or U22223 (N_22223,N_21561,N_21745);
nand U22224 (N_22224,N_21642,N_21993);
and U22225 (N_22225,N_21760,N_21709);
xor U22226 (N_22226,N_21542,N_21569);
nand U22227 (N_22227,N_21812,N_21853);
or U22228 (N_22228,N_21560,N_21883);
or U22229 (N_22229,N_21546,N_21599);
nor U22230 (N_22230,N_21983,N_21956);
and U22231 (N_22231,N_21758,N_21650);
and U22232 (N_22232,N_21571,N_21893);
xnor U22233 (N_22233,N_21657,N_21787);
nor U22234 (N_22234,N_21985,N_21965);
nor U22235 (N_22235,N_21866,N_21741);
xor U22236 (N_22236,N_21530,N_21814);
and U22237 (N_22237,N_21605,N_21538);
nor U22238 (N_22238,N_21901,N_21896);
and U22239 (N_22239,N_21795,N_21753);
xor U22240 (N_22240,N_21660,N_21581);
or U22241 (N_22241,N_21643,N_21554);
nand U22242 (N_22242,N_21947,N_21867);
or U22243 (N_22243,N_21719,N_21981);
nand U22244 (N_22244,N_21655,N_21937);
xor U22245 (N_22245,N_21890,N_21664);
xor U22246 (N_22246,N_21559,N_21512);
nand U22247 (N_22247,N_21638,N_21631);
or U22248 (N_22248,N_21860,N_21844);
nor U22249 (N_22249,N_21873,N_21606);
nand U22250 (N_22250,N_21551,N_21722);
nand U22251 (N_22251,N_21536,N_21810);
and U22252 (N_22252,N_21985,N_21529);
and U22253 (N_22253,N_21574,N_21523);
or U22254 (N_22254,N_21959,N_21907);
and U22255 (N_22255,N_21595,N_21829);
or U22256 (N_22256,N_21607,N_21708);
xor U22257 (N_22257,N_21536,N_21796);
or U22258 (N_22258,N_21775,N_21773);
nor U22259 (N_22259,N_21705,N_21720);
nand U22260 (N_22260,N_21994,N_21550);
nand U22261 (N_22261,N_21955,N_21615);
or U22262 (N_22262,N_21856,N_21883);
or U22263 (N_22263,N_21885,N_21517);
nor U22264 (N_22264,N_21998,N_21980);
xor U22265 (N_22265,N_21563,N_21573);
nand U22266 (N_22266,N_21989,N_21671);
nor U22267 (N_22267,N_21807,N_21862);
xnor U22268 (N_22268,N_21785,N_21891);
xor U22269 (N_22269,N_21619,N_21729);
and U22270 (N_22270,N_21668,N_21963);
xnor U22271 (N_22271,N_21654,N_21751);
and U22272 (N_22272,N_21711,N_21864);
nand U22273 (N_22273,N_21602,N_21515);
xor U22274 (N_22274,N_21898,N_21987);
and U22275 (N_22275,N_21932,N_21524);
nand U22276 (N_22276,N_21705,N_21984);
nor U22277 (N_22277,N_21663,N_21793);
xnor U22278 (N_22278,N_21522,N_21816);
or U22279 (N_22279,N_21512,N_21970);
nor U22280 (N_22280,N_21621,N_21811);
nand U22281 (N_22281,N_21912,N_21745);
xnor U22282 (N_22282,N_21851,N_21514);
nor U22283 (N_22283,N_21854,N_21554);
nand U22284 (N_22284,N_21696,N_21560);
or U22285 (N_22285,N_21514,N_21526);
nand U22286 (N_22286,N_21590,N_21909);
and U22287 (N_22287,N_21864,N_21524);
or U22288 (N_22288,N_21584,N_21711);
and U22289 (N_22289,N_21745,N_21511);
or U22290 (N_22290,N_21545,N_21504);
and U22291 (N_22291,N_21849,N_21973);
nor U22292 (N_22292,N_21788,N_21567);
nand U22293 (N_22293,N_21651,N_21579);
or U22294 (N_22294,N_21643,N_21510);
nand U22295 (N_22295,N_21749,N_21995);
nand U22296 (N_22296,N_21988,N_21813);
and U22297 (N_22297,N_21957,N_21883);
and U22298 (N_22298,N_21916,N_21980);
nor U22299 (N_22299,N_21786,N_21697);
xor U22300 (N_22300,N_21641,N_21696);
xnor U22301 (N_22301,N_21837,N_21508);
nand U22302 (N_22302,N_21722,N_21916);
xor U22303 (N_22303,N_21691,N_21831);
or U22304 (N_22304,N_21797,N_21777);
nand U22305 (N_22305,N_21918,N_21989);
xor U22306 (N_22306,N_21782,N_21627);
nand U22307 (N_22307,N_21656,N_21947);
and U22308 (N_22308,N_21702,N_21748);
nor U22309 (N_22309,N_21577,N_21662);
nand U22310 (N_22310,N_21883,N_21763);
and U22311 (N_22311,N_21933,N_21775);
nand U22312 (N_22312,N_21807,N_21676);
nor U22313 (N_22313,N_21821,N_21828);
nor U22314 (N_22314,N_21577,N_21636);
or U22315 (N_22315,N_21859,N_21993);
and U22316 (N_22316,N_21684,N_21934);
and U22317 (N_22317,N_21655,N_21998);
nand U22318 (N_22318,N_21986,N_21577);
and U22319 (N_22319,N_21879,N_21889);
nor U22320 (N_22320,N_21642,N_21708);
and U22321 (N_22321,N_21617,N_21716);
or U22322 (N_22322,N_21630,N_21516);
or U22323 (N_22323,N_21595,N_21821);
nand U22324 (N_22324,N_21635,N_21930);
nand U22325 (N_22325,N_21660,N_21866);
or U22326 (N_22326,N_21813,N_21629);
and U22327 (N_22327,N_21906,N_21886);
and U22328 (N_22328,N_21814,N_21890);
or U22329 (N_22329,N_21835,N_21545);
or U22330 (N_22330,N_21876,N_21951);
and U22331 (N_22331,N_21503,N_21714);
xor U22332 (N_22332,N_21956,N_21916);
xnor U22333 (N_22333,N_21657,N_21581);
nand U22334 (N_22334,N_21729,N_21789);
or U22335 (N_22335,N_21761,N_21783);
and U22336 (N_22336,N_21803,N_21895);
or U22337 (N_22337,N_21731,N_21814);
xnor U22338 (N_22338,N_21815,N_21745);
and U22339 (N_22339,N_21916,N_21633);
xor U22340 (N_22340,N_21658,N_21861);
nor U22341 (N_22341,N_21647,N_21569);
and U22342 (N_22342,N_21857,N_21824);
nor U22343 (N_22343,N_21585,N_21808);
nor U22344 (N_22344,N_21672,N_21709);
xnor U22345 (N_22345,N_21674,N_21785);
and U22346 (N_22346,N_21609,N_21859);
xor U22347 (N_22347,N_21854,N_21897);
or U22348 (N_22348,N_21809,N_21763);
nand U22349 (N_22349,N_21556,N_21968);
nand U22350 (N_22350,N_21614,N_21540);
or U22351 (N_22351,N_21847,N_21656);
and U22352 (N_22352,N_21929,N_21733);
or U22353 (N_22353,N_21622,N_21856);
xnor U22354 (N_22354,N_21663,N_21545);
or U22355 (N_22355,N_21692,N_21517);
and U22356 (N_22356,N_21663,N_21973);
or U22357 (N_22357,N_21646,N_21721);
or U22358 (N_22358,N_21964,N_21996);
nand U22359 (N_22359,N_21575,N_21568);
and U22360 (N_22360,N_21540,N_21926);
nor U22361 (N_22361,N_21754,N_21968);
xor U22362 (N_22362,N_21950,N_21635);
xnor U22363 (N_22363,N_21557,N_21868);
nand U22364 (N_22364,N_21958,N_21929);
or U22365 (N_22365,N_21745,N_21581);
and U22366 (N_22366,N_21627,N_21563);
or U22367 (N_22367,N_21643,N_21723);
and U22368 (N_22368,N_21796,N_21597);
nor U22369 (N_22369,N_21649,N_21586);
or U22370 (N_22370,N_21792,N_21707);
or U22371 (N_22371,N_21654,N_21799);
nand U22372 (N_22372,N_21675,N_21538);
nand U22373 (N_22373,N_21518,N_21714);
nor U22374 (N_22374,N_21774,N_21675);
nand U22375 (N_22375,N_21622,N_21748);
nand U22376 (N_22376,N_21545,N_21922);
xnor U22377 (N_22377,N_21810,N_21794);
and U22378 (N_22378,N_21693,N_21892);
and U22379 (N_22379,N_21595,N_21570);
xnor U22380 (N_22380,N_21519,N_21768);
xnor U22381 (N_22381,N_21599,N_21940);
nand U22382 (N_22382,N_21813,N_21994);
and U22383 (N_22383,N_21794,N_21741);
and U22384 (N_22384,N_21828,N_21692);
and U22385 (N_22385,N_21957,N_21851);
or U22386 (N_22386,N_21707,N_21988);
nand U22387 (N_22387,N_21941,N_21891);
nor U22388 (N_22388,N_21750,N_21550);
or U22389 (N_22389,N_21902,N_21761);
nand U22390 (N_22390,N_21948,N_21876);
and U22391 (N_22391,N_21544,N_21715);
nor U22392 (N_22392,N_21797,N_21726);
nor U22393 (N_22393,N_21685,N_21711);
xnor U22394 (N_22394,N_21815,N_21733);
xor U22395 (N_22395,N_21892,N_21755);
nor U22396 (N_22396,N_21875,N_21739);
nor U22397 (N_22397,N_21654,N_21825);
and U22398 (N_22398,N_21895,N_21605);
or U22399 (N_22399,N_21888,N_21935);
nor U22400 (N_22400,N_21837,N_21558);
or U22401 (N_22401,N_21638,N_21500);
xnor U22402 (N_22402,N_21704,N_21876);
nand U22403 (N_22403,N_21919,N_21931);
and U22404 (N_22404,N_21578,N_21808);
nand U22405 (N_22405,N_21926,N_21687);
xor U22406 (N_22406,N_21878,N_21765);
or U22407 (N_22407,N_21933,N_21628);
or U22408 (N_22408,N_21663,N_21877);
nor U22409 (N_22409,N_21781,N_21518);
xor U22410 (N_22410,N_21880,N_21658);
and U22411 (N_22411,N_21790,N_21657);
nor U22412 (N_22412,N_21739,N_21640);
or U22413 (N_22413,N_21982,N_21769);
xor U22414 (N_22414,N_21525,N_21722);
and U22415 (N_22415,N_21843,N_21630);
nor U22416 (N_22416,N_21769,N_21541);
xor U22417 (N_22417,N_21755,N_21858);
nand U22418 (N_22418,N_21670,N_21609);
or U22419 (N_22419,N_21743,N_21528);
nor U22420 (N_22420,N_21880,N_21886);
or U22421 (N_22421,N_21641,N_21868);
xor U22422 (N_22422,N_21630,N_21909);
xnor U22423 (N_22423,N_21504,N_21826);
nand U22424 (N_22424,N_21976,N_21857);
nand U22425 (N_22425,N_21742,N_21975);
and U22426 (N_22426,N_21947,N_21950);
nand U22427 (N_22427,N_21577,N_21624);
nand U22428 (N_22428,N_21511,N_21807);
nand U22429 (N_22429,N_21824,N_21887);
and U22430 (N_22430,N_21701,N_21914);
nand U22431 (N_22431,N_21780,N_21979);
xnor U22432 (N_22432,N_21683,N_21524);
xnor U22433 (N_22433,N_21860,N_21542);
nand U22434 (N_22434,N_21736,N_21622);
nor U22435 (N_22435,N_21751,N_21816);
nor U22436 (N_22436,N_21822,N_21590);
xnor U22437 (N_22437,N_21871,N_21502);
nand U22438 (N_22438,N_21785,N_21653);
or U22439 (N_22439,N_21922,N_21784);
nand U22440 (N_22440,N_21572,N_21679);
or U22441 (N_22441,N_21939,N_21544);
or U22442 (N_22442,N_21706,N_21626);
nand U22443 (N_22443,N_21632,N_21615);
nor U22444 (N_22444,N_21553,N_21811);
and U22445 (N_22445,N_21522,N_21644);
nor U22446 (N_22446,N_21859,N_21928);
nor U22447 (N_22447,N_21686,N_21619);
nor U22448 (N_22448,N_21822,N_21605);
nor U22449 (N_22449,N_21633,N_21786);
nor U22450 (N_22450,N_21957,N_21524);
xor U22451 (N_22451,N_21650,N_21763);
or U22452 (N_22452,N_21704,N_21809);
xor U22453 (N_22453,N_21869,N_21604);
nand U22454 (N_22454,N_21525,N_21885);
xnor U22455 (N_22455,N_21995,N_21607);
xnor U22456 (N_22456,N_21577,N_21880);
and U22457 (N_22457,N_21742,N_21570);
nand U22458 (N_22458,N_21714,N_21682);
and U22459 (N_22459,N_21785,N_21741);
nand U22460 (N_22460,N_21583,N_21573);
or U22461 (N_22461,N_21716,N_21648);
and U22462 (N_22462,N_21999,N_21705);
nand U22463 (N_22463,N_21880,N_21756);
or U22464 (N_22464,N_21955,N_21658);
and U22465 (N_22465,N_21504,N_21937);
nor U22466 (N_22466,N_21931,N_21858);
nand U22467 (N_22467,N_21685,N_21576);
xor U22468 (N_22468,N_21730,N_21898);
or U22469 (N_22469,N_21926,N_21873);
nand U22470 (N_22470,N_21686,N_21699);
xor U22471 (N_22471,N_21936,N_21672);
and U22472 (N_22472,N_21949,N_21889);
nand U22473 (N_22473,N_21752,N_21728);
or U22474 (N_22474,N_21705,N_21578);
xnor U22475 (N_22475,N_21973,N_21564);
and U22476 (N_22476,N_21677,N_21743);
nor U22477 (N_22477,N_21562,N_21798);
or U22478 (N_22478,N_21589,N_21781);
and U22479 (N_22479,N_21558,N_21633);
xor U22480 (N_22480,N_21942,N_21720);
or U22481 (N_22481,N_21558,N_21587);
nor U22482 (N_22482,N_21808,N_21909);
xnor U22483 (N_22483,N_21777,N_21816);
nor U22484 (N_22484,N_21531,N_21822);
and U22485 (N_22485,N_21560,N_21656);
and U22486 (N_22486,N_21883,N_21675);
nand U22487 (N_22487,N_21778,N_21892);
xor U22488 (N_22488,N_21719,N_21766);
xor U22489 (N_22489,N_21876,N_21946);
or U22490 (N_22490,N_21882,N_21516);
xnor U22491 (N_22491,N_21541,N_21848);
nand U22492 (N_22492,N_21801,N_21781);
nor U22493 (N_22493,N_21566,N_21966);
xnor U22494 (N_22494,N_21790,N_21586);
or U22495 (N_22495,N_21677,N_21789);
and U22496 (N_22496,N_21952,N_21570);
nand U22497 (N_22497,N_21931,N_21884);
xnor U22498 (N_22498,N_21533,N_21701);
nor U22499 (N_22499,N_21560,N_21603);
nor U22500 (N_22500,N_22199,N_22185);
or U22501 (N_22501,N_22278,N_22114);
xnor U22502 (N_22502,N_22090,N_22388);
xnor U22503 (N_22503,N_22397,N_22365);
nand U22504 (N_22504,N_22154,N_22441);
nand U22505 (N_22505,N_22314,N_22073);
or U22506 (N_22506,N_22000,N_22145);
and U22507 (N_22507,N_22172,N_22244);
nand U22508 (N_22508,N_22336,N_22434);
and U22509 (N_22509,N_22206,N_22093);
nor U22510 (N_22510,N_22236,N_22381);
and U22511 (N_22511,N_22173,N_22363);
or U22512 (N_22512,N_22055,N_22061);
xnor U22513 (N_22513,N_22404,N_22062);
xor U22514 (N_22514,N_22100,N_22376);
nand U22515 (N_22515,N_22182,N_22439);
and U22516 (N_22516,N_22402,N_22086);
nand U22517 (N_22517,N_22006,N_22264);
and U22518 (N_22518,N_22281,N_22470);
nor U22519 (N_22519,N_22495,N_22306);
xnor U22520 (N_22520,N_22010,N_22189);
nor U22521 (N_22521,N_22327,N_22462);
nor U22522 (N_22522,N_22208,N_22083);
nor U22523 (N_22523,N_22337,N_22013);
nor U22524 (N_22524,N_22022,N_22012);
nor U22525 (N_22525,N_22028,N_22394);
xor U22526 (N_22526,N_22467,N_22478);
xor U22527 (N_22527,N_22225,N_22252);
xor U22528 (N_22528,N_22274,N_22096);
and U22529 (N_22529,N_22226,N_22435);
and U22530 (N_22530,N_22285,N_22333);
nand U22531 (N_22531,N_22111,N_22192);
nor U22532 (N_22532,N_22380,N_22047);
xor U22533 (N_22533,N_22157,N_22117);
xor U22534 (N_22534,N_22347,N_22104);
and U22535 (N_22535,N_22403,N_22009);
xor U22536 (N_22536,N_22190,N_22140);
and U22537 (N_22537,N_22254,N_22448);
and U22538 (N_22538,N_22310,N_22019);
or U22539 (N_22539,N_22094,N_22121);
or U22540 (N_22540,N_22427,N_22144);
nor U22541 (N_22541,N_22084,N_22491);
nand U22542 (N_22542,N_22414,N_22210);
nand U22543 (N_22543,N_22110,N_22128);
nor U22544 (N_22544,N_22302,N_22422);
xnor U22545 (N_22545,N_22139,N_22450);
nand U22546 (N_22546,N_22361,N_22123);
nor U22547 (N_22547,N_22358,N_22266);
nand U22548 (N_22548,N_22048,N_22168);
xor U22549 (N_22549,N_22290,N_22250);
and U22550 (N_22550,N_22288,N_22178);
and U22551 (N_22551,N_22202,N_22359);
nand U22552 (N_22552,N_22300,N_22280);
nor U22553 (N_22553,N_22227,N_22391);
nor U22554 (N_22554,N_22315,N_22143);
and U22555 (N_22555,N_22122,N_22112);
nor U22556 (N_22556,N_22166,N_22078);
xor U22557 (N_22557,N_22444,N_22385);
xnor U22558 (N_22558,N_22364,N_22423);
nor U22559 (N_22559,N_22301,N_22432);
or U22560 (N_22560,N_22241,N_22308);
nor U22561 (N_22561,N_22375,N_22187);
xor U22562 (N_22562,N_22490,N_22238);
or U22563 (N_22563,N_22319,N_22344);
nor U22564 (N_22564,N_22455,N_22255);
or U22565 (N_22565,N_22379,N_22102);
nor U22566 (N_22566,N_22029,N_22142);
nand U22567 (N_22567,N_22007,N_22454);
and U22568 (N_22568,N_22179,N_22366);
nor U22569 (N_22569,N_22485,N_22223);
xor U22570 (N_22570,N_22228,N_22392);
and U22571 (N_22571,N_22311,N_22080);
or U22572 (N_22572,N_22198,N_22235);
nor U22573 (N_22573,N_22175,N_22204);
or U22574 (N_22574,N_22445,N_22463);
or U22575 (N_22575,N_22262,N_22234);
nand U22576 (N_22576,N_22430,N_22025);
and U22577 (N_22577,N_22256,N_22098);
and U22578 (N_22578,N_22353,N_22473);
nand U22579 (N_22579,N_22351,N_22369);
or U22580 (N_22580,N_22307,N_22471);
nand U22581 (N_22581,N_22127,N_22109);
or U22582 (N_22582,N_22410,N_22312);
nor U22583 (N_22583,N_22212,N_22095);
nor U22584 (N_22584,N_22418,N_22405);
or U22585 (N_22585,N_22461,N_22395);
xnor U22586 (N_22586,N_22220,N_22267);
and U22587 (N_22587,N_22457,N_22494);
nor U22588 (N_22588,N_22456,N_22085);
xnor U22589 (N_22589,N_22041,N_22106);
xnor U22590 (N_22590,N_22331,N_22177);
nand U22591 (N_22591,N_22350,N_22245);
nor U22592 (N_22592,N_22211,N_22174);
xnor U22593 (N_22593,N_22037,N_22477);
xnor U22594 (N_22594,N_22289,N_22400);
or U22595 (N_22595,N_22149,N_22341);
nor U22596 (N_22596,N_22039,N_22035);
or U22597 (N_22597,N_22387,N_22453);
nand U22598 (N_22598,N_22357,N_22382);
nand U22599 (N_22599,N_22325,N_22378);
nor U22600 (N_22600,N_22401,N_22326);
xor U22601 (N_22601,N_22188,N_22354);
nand U22602 (N_22602,N_22156,N_22346);
or U22603 (N_22603,N_22134,N_22042);
and U22604 (N_22604,N_22167,N_22097);
nand U22605 (N_22605,N_22129,N_22051);
and U22606 (N_22606,N_22087,N_22329);
nor U22607 (N_22607,N_22322,N_22049);
nor U22608 (N_22608,N_22053,N_22474);
nor U22609 (N_22609,N_22396,N_22024);
or U22610 (N_22610,N_22089,N_22120);
or U22611 (N_22611,N_22092,N_22304);
nor U22612 (N_22612,N_22483,N_22480);
and U22613 (N_22613,N_22340,N_22355);
nand U22614 (N_22614,N_22107,N_22272);
xnor U22615 (N_22615,N_22437,N_22240);
or U22616 (N_22616,N_22413,N_22031);
or U22617 (N_22617,N_22260,N_22181);
and U22618 (N_22618,N_22425,N_22229);
xnor U22619 (N_22619,N_22348,N_22020);
nor U22620 (N_22620,N_22384,N_22158);
or U22621 (N_22621,N_22066,N_22076);
or U22622 (N_22622,N_22215,N_22295);
nand U22623 (N_22623,N_22360,N_22472);
nand U22624 (N_22624,N_22390,N_22148);
xor U22625 (N_22625,N_22277,N_22044);
and U22626 (N_22626,N_22194,N_22151);
or U22627 (N_22627,N_22313,N_22023);
xnor U22628 (N_22628,N_22057,N_22014);
and U22629 (N_22629,N_22032,N_22299);
nand U22630 (N_22630,N_22040,N_22291);
and U22631 (N_22631,N_22161,N_22294);
nand U22632 (N_22632,N_22251,N_22270);
nand U22633 (N_22633,N_22216,N_22071);
xor U22634 (N_22634,N_22214,N_22424);
or U22635 (N_22635,N_22072,N_22003);
and U22636 (N_22636,N_22162,N_22004);
nor U22637 (N_22637,N_22408,N_22159);
or U22638 (N_22638,N_22372,N_22033);
xor U22639 (N_22639,N_22409,N_22452);
and U22640 (N_22640,N_22116,N_22059);
or U22641 (N_22641,N_22416,N_22165);
or U22642 (N_22642,N_22428,N_22303);
and U22643 (N_22643,N_22339,N_22016);
nor U22644 (N_22644,N_22176,N_22253);
or U22645 (N_22645,N_22328,N_22497);
or U22646 (N_22646,N_22034,N_22440);
or U22647 (N_22647,N_22222,N_22335);
and U22648 (N_22648,N_22421,N_22065);
nand U22649 (N_22649,N_22015,N_22449);
nand U22650 (N_22650,N_22183,N_22332);
or U22651 (N_22651,N_22130,N_22398);
nor U22652 (N_22652,N_22153,N_22077);
and U22653 (N_22653,N_22163,N_22258);
or U22654 (N_22654,N_22242,N_22276);
xor U22655 (N_22655,N_22233,N_22002);
and U22656 (N_22656,N_22433,N_22481);
xor U22657 (N_22657,N_22321,N_22263);
nor U22658 (N_22658,N_22476,N_22133);
nor U22659 (N_22659,N_22279,N_22058);
nor U22660 (N_22660,N_22468,N_22492);
nor U22661 (N_22661,N_22108,N_22249);
xor U22662 (N_22662,N_22067,N_22498);
or U22663 (N_22663,N_22323,N_22011);
and U22664 (N_22664,N_22487,N_22054);
and U22665 (N_22665,N_22493,N_22486);
nor U22666 (N_22666,N_22237,N_22091);
nor U22667 (N_22667,N_22406,N_22197);
nor U22668 (N_22668,N_22268,N_22180);
nor U22669 (N_22669,N_22038,N_22451);
xor U22670 (N_22670,N_22368,N_22287);
or U22671 (N_22671,N_22207,N_22259);
nor U22672 (N_22672,N_22027,N_22146);
nand U22673 (N_22673,N_22105,N_22407);
nor U22674 (N_22674,N_22217,N_22005);
nand U22675 (N_22675,N_22412,N_22115);
xor U22676 (N_22676,N_22273,N_22431);
or U22677 (N_22677,N_22152,N_22318);
and U22678 (N_22678,N_22160,N_22209);
and U22679 (N_22679,N_22320,N_22283);
nor U22680 (N_22680,N_22482,N_22317);
nand U22681 (N_22681,N_22219,N_22488);
or U22682 (N_22682,N_22045,N_22246);
or U22683 (N_22683,N_22309,N_22021);
nand U22684 (N_22684,N_22442,N_22284);
nor U22685 (N_22685,N_22196,N_22371);
xor U22686 (N_22686,N_22075,N_22298);
xor U22687 (N_22687,N_22186,N_22411);
nor U22688 (N_22688,N_22138,N_22113);
and U22689 (N_22689,N_22374,N_22184);
or U22690 (N_22690,N_22213,N_22074);
nand U22691 (N_22691,N_22218,N_22099);
or U22692 (N_22692,N_22417,N_22201);
nand U22693 (N_22693,N_22271,N_22356);
and U22694 (N_22694,N_22008,N_22286);
and U22695 (N_22695,N_22060,N_22224);
nand U22696 (N_22696,N_22275,N_22484);
xnor U22697 (N_22697,N_22499,N_22131);
or U22698 (N_22698,N_22293,N_22338);
nor U22699 (N_22699,N_22330,N_22050);
nor U22700 (N_22700,N_22026,N_22458);
nor U22701 (N_22701,N_22393,N_22030);
xnor U22702 (N_22702,N_22324,N_22269);
and U22703 (N_22703,N_22261,N_22043);
nor U22704 (N_22704,N_22386,N_22118);
xor U22705 (N_22705,N_22170,N_22248);
nor U22706 (N_22706,N_22345,N_22082);
xnor U22707 (N_22707,N_22136,N_22389);
nor U22708 (N_22708,N_22081,N_22195);
nand U22709 (N_22709,N_22446,N_22069);
xor U22710 (N_22710,N_22377,N_22230);
nand U22711 (N_22711,N_22475,N_22018);
nor U22712 (N_22712,N_22046,N_22367);
and U22713 (N_22713,N_22334,N_22342);
xnor U22714 (N_22714,N_22017,N_22126);
and U22715 (N_22715,N_22362,N_22466);
or U22716 (N_22716,N_22150,N_22103);
xnor U22717 (N_22717,N_22079,N_22420);
xnor U22718 (N_22718,N_22419,N_22088);
xor U22719 (N_22719,N_22068,N_22489);
and U22720 (N_22720,N_22155,N_22265);
nand U22721 (N_22721,N_22171,N_22459);
nand U22722 (N_22722,N_22137,N_22429);
nand U22723 (N_22723,N_22436,N_22247);
nand U22724 (N_22724,N_22231,N_22232);
and U22725 (N_22725,N_22239,N_22001);
and U22726 (N_22726,N_22169,N_22305);
nor U22727 (N_22727,N_22205,N_22316);
xnor U22728 (N_22728,N_22056,N_22052);
or U22729 (N_22729,N_22124,N_22297);
and U22730 (N_22730,N_22464,N_22221);
nor U22731 (N_22731,N_22063,N_22141);
nand U22732 (N_22732,N_22438,N_22164);
and U22733 (N_22733,N_22292,N_22399);
and U22734 (N_22734,N_22479,N_22147);
xnor U22735 (N_22735,N_22193,N_22349);
nor U22736 (N_22736,N_22036,N_22373);
and U22737 (N_22737,N_22352,N_22426);
xnor U22738 (N_22738,N_22465,N_22343);
or U22739 (N_22739,N_22125,N_22191);
and U22740 (N_22740,N_22070,N_22383);
xor U22741 (N_22741,N_22064,N_22119);
nand U22742 (N_22742,N_22200,N_22296);
or U22743 (N_22743,N_22257,N_22282);
xnor U22744 (N_22744,N_22203,N_22447);
nand U22745 (N_22745,N_22135,N_22101);
xnor U22746 (N_22746,N_22415,N_22370);
or U22747 (N_22747,N_22132,N_22460);
nor U22748 (N_22748,N_22443,N_22496);
xnor U22749 (N_22749,N_22243,N_22469);
nor U22750 (N_22750,N_22176,N_22242);
or U22751 (N_22751,N_22302,N_22036);
or U22752 (N_22752,N_22489,N_22113);
nand U22753 (N_22753,N_22307,N_22108);
nand U22754 (N_22754,N_22020,N_22442);
or U22755 (N_22755,N_22332,N_22336);
or U22756 (N_22756,N_22485,N_22170);
or U22757 (N_22757,N_22096,N_22207);
or U22758 (N_22758,N_22234,N_22096);
or U22759 (N_22759,N_22435,N_22365);
and U22760 (N_22760,N_22091,N_22491);
nor U22761 (N_22761,N_22269,N_22004);
nand U22762 (N_22762,N_22418,N_22119);
nand U22763 (N_22763,N_22210,N_22147);
nor U22764 (N_22764,N_22096,N_22108);
nand U22765 (N_22765,N_22030,N_22398);
nand U22766 (N_22766,N_22408,N_22326);
or U22767 (N_22767,N_22103,N_22446);
nand U22768 (N_22768,N_22038,N_22323);
nand U22769 (N_22769,N_22066,N_22361);
and U22770 (N_22770,N_22136,N_22461);
and U22771 (N_22771,N_22307,N_22188);
xnor U22772 (N_22772,N_22190,N_22463);
or U22773 (N_22773,N_22236,N_22122);
nand U22774 (N_22774,N_22067,N_22034);
nor U22775 (N_22775,N_22292,N_22483);
xnor U22776 (N_22776,N_22102,N_22338);
and U22777 (N_22777,N_22465,N_22034);
xnor U22778 (N_22778,N_22393,N_22048);
and U22779 (N_22779,N_22417,N_22270);
nor U22780 (N_22780,N_22048,N_22008);
or U22781 (N_22781,N_22149,N_22296);
and U22782 (N_22782,N_22125,N_22268);
xnor U22783 (N_22783,N_22383,N_22312);
nor U22784 (N_22784,N_22088,N_22321);
nor U22785 (N_22785,N_22185,N_22097);
and U22786 (N_22786,N_22324,N_22434);
nor U22787 (N_22787,N_22430,N_22313);
or U22788 (N_22788,N_22177,N_22164);
and U22789 (N_22789,N_22465,N_22009);
or U22790 (N_22790,N_22222,N_22026);
nor U22791 (N_22791,N_22326,N_22342);
xnor U22792 (N_22792,N_22249,N_22091);
or U22793 (N_22793,N_22246,N_22253);
or U22794 (N_22794,N_22098,N_22332);
nand U22795 (N_22795,N_22215,N_22007);
and U22796 (N_22796,N_22472,N_22044);
or U22797 (N_22797,N_22437,N_22058);
nor U22798 (N_22798,N_22420,N_22327);
or U22799 (N_22799,N_22319,N_22288);
xor U22800 (N_22800,N_22496,N_22228);
nand U22801 (N_22801,N_22334,N_22434);
xor U22802 (N_22802,N_22370,N_22156);
nor U22803 (N_22803,N_22207,N_22106);
or U22804 (N_22804,N_22336,N_22085);
xnor U22805 (N_22805,N_22484,N_22340);
xnor U22806 (N_22806,N_22089,N_22487);
nand U22807 (N_22807,N_22092,N_22123);
xor U22808 (N_22808,N_22363,N_22440);
nand U22809 (N_22809,N_22078,N_22324);
nand U22810 (N_22810,N_22215,N_22120);
and U22811 (N_22811,N_22372,N_22258);
nor U22812 (N_22812,N_22361,N_22401);
nor U22813 (N_22813,N_22487,N_22301);
and U22814 (N_22814,N_22459,N_22389);
nor U22815 (N_22815,N_22229,N_22078);
and U22816 (N_22816,N_22105,N_22246);
and U22817 (N_22817,N_22055,N_22150);
nor U22818 (N_22818,N_22411,N_22071);
nor U22819 (N_22819,N_22150,N_22177);
xor U22820 (N_22820,N_22410,N_22496);
nand U22821 (N_22821,N_22333,N_22420);
nor U22822 (N_22822,N_22336,N_22283);
nor U22823 (N_22823,N_22219,N_22187);
or U22824 (N_22824,N_22213,N_22484);
xnor U22825 (N_22825,N_22497,N_22072);
xor U22826 (N_22826,N_22289,N_22238);
or U22827 (N_22827,N_22319,N_22132);
and U22828 (N_22828,N_22025,N_22066);
xor U22829 (N_22829,N_22394,N_22456);
xor U22830 (N_22830,N_22052,N_22468);
nor U22831 (N_22831,N_22391,N_22275);
nor U22832 (N_22832,N_22003,N_22477);
and U22833 (N_22833,N_22104,N_22276);
nor U22834 (N_22834,N_22272,N_22473);
nand U22835 (N_22835,N_22051,N_22055);
or U22836 (N_22836,N_22061,N_22212);
nand U22837 (N_22837,N_22382,N_22378);
and U22838 (N_22838,N_22312,N_22088);
nor U22839 (N_22839,N_22092,N_22392);
and U22840 (N_22840,N_22245,N_22312);
or U22841 (N_22841,N_22496,N_22112);
xnor U22842 (N_22842,N_22374,N_22249);
xnor U22843 (N_22843,N_22075,N_22280);
and U22844 (N_22844,N_22095,N_22013);
nand U22845 (N_22845,N_22316,N_22411);
and U22846 (N_22846,N_22057,N_22375);
nand U22847 (N_22847,N_22027,N_22200);
nand U22848 (N_22848,N_22171,N_22134);
nand U22849 (N_22849,N_22466,N_22287);
xor U22850 (N_22850,N_22284,N_22430);
nor U22851 (N_22851,N_22365,N_22440);
nor U22852 (N_22852,N_22048,N_22346);
or U22853 (N_22853,N_22006,N_22294);
nor U22854 (N_22854,N_22117,N_22287);
nand U22855 (N_22855,N_22014,N_22389);
nor U22856 (N_22856,N_22438,N_22412);
xnor U22857 (N_22857,N_22117,N_22273);
nor U22858 (N_22858,N_22072,N_22162);
xnor U22859 (N_22859,N_22289,N_22089);
or U22860 (N_22860,N_22437,N_22106);
nor U22861 (N_22861,N_22133,N_22278);
or U22862 (N_22862,N_22370,N_22225);
nor U22863 (N_22863,N_22019,N_22487);
and U22864 (N_22864,N_22358,N_22033);
xor U22865 (N_22865,N_22162,N_22358);
nor U22866 (N_22866,N_22448,N_22056);
nor U22867 (N_22867,N_22283,N_22047);
nand U22868 (N_22868,N_22313,N_22283);
nor U22869 (N_22869,N_22430,N_22311);
nand U22870 (N_22870,N_22489,N_22132);
xnor U22871 (N_22871,N_22472,N_22045);
xor U22872 (N_22872,N_22218,N_22249);
xor U22873 (N_22873,N_22001,N_22039);
xnor U22874 (N_22874,N_22180,N_22494);
or U22875 (N_22875,N_22433,N_22450);
or U22876 (N_22876,N_22064,N_22356);
nor U22877 (N_22877,N_22075,N_22003);
and U22878 (N_22878,N_22067,N_22304);
nor U22879 (N_22879,N_22054,N_22247);
nor U22880 (N_22880,N_22118,N_22499);
nor U22881 (N_22881,N_22494,N_22155);
xor U22882 (N_22882,N_22377,N_22426);
or U22883 (N_22883,N_22442,N_22496);
nand U22884 (N_22884,N_22427,N_22221);
or U22885 (N_22885,N_22244,N_22360);
xor U22886 (N_22886,N_22235,N_22116);
nand U22887 (N_22887,N_22265,N_22386);
xor U22888 (N_22888,N_22113,N_22151);
or U22889 (N_22889,N_22434,N_22145);
or U22890 (N_22890,N_22054,N_22006);
nand U22891 (N_22891,N_22136,N_22082);
xor U22892 (N_22892,N_22200,N_22489);
or U22893 (N_22893,N_22179,N_22340);
or U22894 (N_22894,N_22459,N_22277);
and U22895 (N_22895,N_22099,N_22348);
or U22896 (N_22896,N_22078,N_22456);
or U22897 (N_22897,N_22017,N_22415);
nand U22898 (N_22898,N_22298,N_22160);
xor U22899 (N_22899,N_22151,N_22015);
or U22900 (N_22900,N_22218,N_22358);
and U22901 (N_22901,N_22368,N_22372);
xnor U22902 (N_22902,N_22229,N_22452);
nor U22903 (N_22903,N_22090,N_22282);
nand U22904 (N_22904,N_22453,N_22186);
or U22905 (N_22905,N_22289,N_22305);
nor U22906 (N_22906,N_22079,N_22017);
and U22907 (N_22907,N_22443,N_22188);
xor U22908 (N_22908,N_22267,N_22350);
nor U22909 (N_22909,N_22095,N_22089);
and U22910 (N_22910,N_22275,N_22399);
and U22911 (N_22911,N_22359,N_22184);
or U22912 (N_22912,N_22166,N_22408);
or U22913 (N_22913,N_22311,N_22061);
or U22914 (N_22914,N_22103,N_22094);
nor U22915 (N_22915,N_22023,N_22242);
and U22916 (N_22916,N_22372,N_22323);
nor U22917 (N_22917,N_22332,N_22279);
nand U22918 (N_22918,N_22472,N_22239);
nor U22919 (N_22919,N_22289,N_22144);
or U22920 (N_22920,N_22414,N_22379);
or U22921 (N_22921,N_22257,N_22423);
and U22922 (N_22922,N_22309,N_22376);
or U22923 (N_22923,N_22104,N_22234);
nand U22924 (N_22924,N_22272,N_22454);
or U22925 (N_22925,N_22276,N_22249);
xor U22926 (N_22926,N_22250,N_22184);
xnor U22927 (N_22927,N_22007,N_22281);
nand U22928 (N_22928,N_22272,N_22283);
or U22929 (N_22929,N_22446,N_22138);
xor U22930 (N_22930,N_22124,N_22143);
xor U22931 (N_22931,N_22451,N_22019);
or U22932 (N_22932,N_22311,N_22283);
nor U22933 (N_22933,N_22210,N_22299);
and U22934 (N_22934,N_22437,N_22390);
nor U22935 (N_22935,N_22204,N_22456);
nand U22936 (N_22936,N_22036,N_22273);
and U22937 (N_22937,N_22324,N_22424);
xnor U22938 (N_22938,N_22247,N_22232);
xor U22939 (N_22939,N_22108,N_22277);
or U22940 (N_22940,N_22340,N_22276);
xnor U22941 (N_22941,N_22226,N_22444);
and U22942 (N_22942,N_22004,N_22331);
nor U22943 (N_22943,N_22489,N_22378);
and U22944 (N_22944,N_22331,N_22060);
nand U22945 (N_22945,N_22388,N_22391);
nor U22946 (N_22946,N_22065,N_22132);
nor U22947 (N_22947,N_22228,N_22183);
or U22948 (N_22948,N_22478,N_22037);
nor U22949 (N_22949,N_22366,N_22053);
xor U22950 (N_22950,N_22030,N_22372);
nor U22951 (N_22951,N_22062,N_22081);
xor U22952 (N_22952,N_22063,N_22277);
nand U22953 (N_22953,N_22180,N_22176);
xor U22954 (N_22954,N_22200,N_22055);
nor U22955 (N_22955,N_22231,N_22031);
and U22956 (N_22956,N_22050,N_22001);
and U22957 (N_22957,N_22458,N_22492);
xnor U22958 (N_22958,N_22173,N_22401);
xor U22959 (N_22959,N_22095,N_22203);
nor U22960 (N_22960,N_22044,N_22111);
and U22961 (N_22961,N_22117,N_22257);
nand U22962 (N_22962,N_22115,N_22227);
xnor U22963 (N_22963,N_22460,N_22209);
nand U22964 (N_22964,N_22044,N_22010);
nor U22965 (N_22965,N_22472,N_22081);
xor U22966 (N_22966,N_22051,N_22483);
or U22967 (N_22967,N_22246,N_22124);
xor U22968 (N_22968,N_22304,N_22063);
nand U22969 (N_22969,N_22280,N_22492);
and U22970 (N_22970,N_22096,N_22236);
xnor U22971 (N_22971,N_22123,N_22206);
and U22972 (N_22972,N_22446,N_22250);
or U22973 (N_22973,N_22278,N_22051);
nand U22974 (N_22974,N_22346,N_22176);
or U22975 (N_22975,N_22411,N_22422);
nor U22976 (N_22976,N_22495,N_22182);
and U22977 (N_22977,N_22180,N_22348);
and U22978 (N_22978,N_22078,N_22297);
and U22979 (N_22979,N_22330,N_22343);
and U22980 (N_22980,N_22320,N_22355);
nand U22981 (N_22981,N_22466,N_22102);
nand U22982 (N_22982,N_22215,N_22309);
or U22983 (N_22983,N_22470,N_22319);
xor U22984 (N_22984,N_22343,N_22489);
nor U22985 (N_22985,N_22148,N_22100);
nand U22986 (N_22986,N_22246,N_22449);
xnor U22987 (N_22987,N_22016,N_22179);
and U22988 (N_22988,N_22280,N_22179);
or U22989 (N_22989,N_22142,N_22374);
nand U22990 (N_22990,N_22220,N_22315);
or U22991 (N_22991,N_22256,N_22402);
or U22992 (N_22992,N_22002,N_22391);
xor U22993 (N_22993,N_22041,N_22231);
nand U22994 (N_22994,N_22319,N_22215);
nor U22995 (N_22995,N_22248,N_22413);
nand U22996 (N_22996,N_22487,N_22050);
nand U22997 (N_22997,N_22230,N_22041);
xor U22998 (N_22998,N_22153,N_22027);
xnor U22999 (N_22999,N_22295,N_22064);
or U23000 (N_23000,N_22564,N_22825);
nand U23001 (N_23001,N_22765,N_22929);
and U23002 (N_23002,N_22840,N_22889);
nor U23003 (N_23003,N_22969,N_22565);
and U23004 (N_23004,N_22618,N_22714);
nand U23005 (N_23005,N_22536,N_22721);
nor U23006 (N_23006,N_22879,N_22936);
or U23007 (N_23007,N_22801,N_22973);
and U23008 (N_23008,N_22788,N_22830);
and U23009 (N_23009,N_22539,N_22573);
nand U23010 (N_23010,N_22997,N_22548);
xor U23011 (N_23011,N_22995,N_22815);
nand U23012 (N_23012,N_22975,N_22747);
xor U23013 (N_23013,N_22550,N_22594);
nor U23014 (N_23014,N_22692,N_22726);
xor U23015 (N_23015,N_22895,N_22526);
or U23016 (N_23016,N_22650,N_22639);
or U23017 (N_23017,N_22532,N_22857);
and U23018 (N_23018,N_22768,N_22655);
nor U23019 (N_23019,N_22921,N_22587);
nand U23020 (N_23020,N_22715,N_22898);
nor U23021 (N_23021,N_22876,N_22673);
and U23022 (N_23022,N_22933,N_22525);
nor U23023 (N_23023,N_22654,N_22880);
xor U23024 (N_23024,N_22704,N_22868);
or U23025 (N_23025,N_22771,N_22516);
nor U23026 (N_23026,N_22817,N_22527);
nand U23027 (N_23027,N_22711,N_22870);
xor U23028 (N_23028,N_22700,N_22632);
nand U23029 (N_23029,N_22619,N_22845);
nor U23030 (N_23030,N_22635,N_22897);
or U23031 (N_23031,N_22620,N_22719);
and U23032 (N_23032,N_22993,N_22987);
xor U23033 (N_23033,N_22598,N_22760);
and U23034 (N_23034,N_22580,N_22528);
or U23035 (N_23035,N_22784,N_22800);
or U23036 (N_23036,N_22685,N_22510);
nand U23037 (N_23037,N_22930,N_22579);
nor U23038 (N_23038,N_22605,N_22622);
xor U23039 (N_23039,N_22843,N_22855);
xor U23040 (N_23040,N_22574,N_22637);
nor U23041 (N_23041,N_22856,N_22699);
nand U23042 (N_23042,N_22575,N_22567);
xnor U23043 (N_23043,N_22546,N_22831);
and U23044 (N_23044,N_22976,N_22529);
xnor U23045 (N_23045,N_22810,N_22723);
xor U23046 (N_23046,N_22675,N_22996);
xnor U23047 (N_23047,N_22724,N_22982);
and U23048 (N_23048,N_22813,N_22649);
nand U23049 (N_23049,N_22871,N_22560);
nand U23050 (N_23050,N_22551,N_22906);
and U23051 (N_23051,N_22854,N_22980);
xor U23052 (N_23052,N_22506,N_22659);
nor U23053 (N_23053,N_22500,N_22571);
nand U23054 (N_23054,N_22803,N_22954);
nand U23055 (N_23055,N_22535,N_22645);
xor U23056 (N_23056,N_22629,N_22623);
or U23057 (N_23057,N_22584,N_22609);
xnor U23058 (N_23058,N_22802,N_22811);
xnor U23059 (N_23059,N_22823,N_22896);
nand U23060 (N_23060,N_22706,N_22901);
nor U23061 (N_23061,N_22660,N_22716);
or U23062 (N_23062,N_22948,N_22819);
nand U23063 (N_23063,N_22783,N_22967);
and U23064 (N_23064,N_22873,N_22977);
nand U23065 (N_23065,N_22824,N_22520);
and U23066 (N_23066,N_22956,N_22826);
or U23067 (N_23067,N_22713,N_22557);
nor U23068 (N_23068,N_22607,N_22989);
nor U23069 (N_23069,N_22661,N_22746);
xor U23070 (N_23070,N_22991,N_22778);
nand U23071 (N_23071,N_22985,N_22517);
and U23072 (N_23072,N_22644,N_22938);
nor U23073 (N_23073,N_22702,N_22545);
and U23074 (N_23074,N_22931,N_22749);
or U23075 (N_23075,N_22904,N_22730);
nor U23076 (N_23076,N_22616,N_22836);
nand U23077 (N_23077,N_22858,N_22828);
and U23078 (N_23078,N_22887,N_22566);
and U23079 (N_23079,N_22615,N_22795);
nand U23080 (N_23080,N_22552,N_22884);
nor U23081 (N_23081,N_22925,N_22841);
nand U23082 (N_23082,N_22842,N_22767);
nor U23083 (N_23083,N_22988,N_22847);
nor U23084 (N_23084,N_22701,N_22742);
xnor U23085 (N_23085,N_22777,N_22761);
nor U23086 (N_23086,N_22739,N_22533);
xnor U23087 (N_23087,N_22709,N_22790);
and U23088 (N_23088,N_22829,N_22658);
xor U23089 (N_23089,N_22869,N_22596);
xnor U23090 (N_23090,N_22792,N_22923);
nand U23091 (N_23091,N_22983,N_22643);
or U23092 (N_23092,N_22950,N_22791);
xnor U23093 (N_23093,N_22908,N_22787);
nand U23094 (N_23094,N_22591,N_22668);
nor U23095 (N_23095,N_22769,N_22772);
or U23096 (N_23096,N_22662,N_22505);
nor U23097 (N_23097,N_22537,N_22577);
or U23098 (N_23098,N_22612,N_22893);
or U23099 (N_23099,N_22611,N_22634);
or U23100 (N_23100,N_22762,N_22676);
nand U23101 (N_23101,N_22955,N_22720);
or U23102 (N_23102,N_22695,N_22859);
and U23103 (N_23103,N_22741,N_22670);
and U23104 (N_23104,N_22927,N_22883);
xor U23105 (N_23105,N_22912,N_22846);
nor U23106 (N_23106,N_22853,N_22542);
nor U23107 (N_23107,N_22899,N_22595);
nor U23108 (N_23108,N_22578,N_22894);
xor U23109 (N_23109,N_22852,N_22850);
nand U23110 (N_23110,N_22682,N_22652);
and U23111 (N_23111,N_22805,N_22888);
nand U23112 (N_23112,N_22759,N_22944);
and U23113 (N_23113,N_22610,N_22986);
and U23114 (N_23114,N_22885,N_22809);
or U23115 (N_23115,N_22971,N_22748);
xnor U23116 (N_23116,N_22530,N_22621);
nand U23117 (N_23117,N_22909,N_22672);
nor U23118 (N_23118,N_22903,N_22628);
nor U23119 (N_23119,N_22754,N_22559);
and U23120 (N_23120,N_22835,N_22625);
or U23121 (N_23121,N_22592,N_22642);
xor U23122 (N_23122,N_22934,N_22838);
xnor U23123 (N_23123,N_22796,N_22808);
nor U23124 (N_23124,N_22666,N_22816);
xnor U23125 (N_23125,N_22943,N_22866);
xnor U23126 (N_23126,N_22663,N_22501);
nor U23127 (N_23127,N_22907,N_22569);
nand U23128 (N_23128,N_22799,N_22555);
and U23129 (N_23129,N_22727,N_22910);
or U23130 (N_23130,N_22671,N_22820);
nand U23131 (N_23131,N_22599,N_22547);
xor U23132 (N_23132,N_22593,N_22696);
or U23133 (N_23133,N_22710,N_22738);
nand U23134 (N_23134,N_22538,N_22686);
xor U23135 (N_23135,N_22945,N_22729);
xor U23136 (N_23136,N_22960,N_22563);
nor U23137 (N_23137,N_22582,N_22914);
and U23138 (N_23138,N_22583,N_22750);
and U23139 (N_23139,N_22794,N_22689);
nand U23140 (N_23140,N_22863,N_22683);
nor U23141 (N_23141,N_22981,N_22603);
nor U23142 (N_23142,N_22917,N_22946);
or U23143 (N_23143,N_22608,N_22782);
nand U23144 (N_23144,N_22740,N_22998);
nand U23145 (N_23145,N_22614,N_22789);
or U23146 (N_23146,N_22941,N_22890);
nor U23147 (N_23147,N_22877,N_22556);
or U23148 (N_23148,N_22703,N_22600);
and U23149 (N_23149,N_22631,N_22867);
and U23150 (N_23150,N_22648,N_22543);
nand U23151 (N_23151,N_22734,N_22679);
xor U23152 (N_23152,N_22667,N_22776);
and U23153 (N_23153,N_22570,N_22743);
and U23154 (N_23154,N_22990,N_22961);
and U23155 (N_23155,N_22900,N_22509);
or U23156 (N_23156,N_22585,N_22959);
and U23157 (N_23157,N_22544,N_22725);
xor U23158 (N_23158,N_22681,N_22504);
nand U23159 (N_23159,N_22974,N_22606);
nand U23160 (N_23160,N_22572,N_22953);
nor U23161 (N_23161,N_22744,N_22657);
nor U23162 (N_23162,N_22522,N_22979);
nor U23163 (N_23163,N_22718,N_22844);
nand U23164 (N_23164,N_22892,N_22833);
nand U23165 (N_23165,N_22602,N_22732);
xnor U23166 (N_23166,N_22865,N_22878);
nor U23167 (N_23167,N_22839,N_22753);
and U23168 (N_23168,N_22804,N_22807);
and U23169 (N_23169,N_22766,N_22786);
nor U23170 (N_23170,N_22519,N_22669);
xor U23171 (N_23171,N_22736,N_22947);
and U23172 (N_23172,N_22624,N_22687);
nand U23173 (N_23173,N_22864,N_22656);
or U23174 (N_23174,N_22638,N_22968);
and U23175 (N_23175,N_22940,N_22832);
and U23176 (N_23176,N_22994,N_22918);
and U23177 (N_23177,N_22674,N_22779);
nor U23178 (N_23178,N_22881,N_22717);
and U23179 (N_23179,N_22919,N_22935);
nor U23180 (N_23180,N_22920,N_22797);
nand U23181 (N_23181,N_22874,N_22922);
and U23182 (N_23182,N_22680,N_22722);
nor U23183 (N_23183,N_22688,N_22756);
nor U23184 (N_23184,N_22951,N_22735);
and U23185 (N_23185,N_22641,N_22834);
xnor U23186 (N_23186,N_22949,N_22640);
and U23187 (N_23187,N_22693,N_22586);
nor U23188 (N_23188,N_22952,N_22626);
and U23189 (N_23189,N_22678,N_22916);
nor U23190 (N_23190,N_22915,N_22924);
nor U23191 (N_23191,N_22745,N_22524);
xnor U23192 (N_23192,N_22939,N_22707);
nand U23193 (N_23193,N_22531,N_22646);
xnor U23194 (N_23194,N_22515,N_22962);
xor U23195 (N_23195,N_22568,N_22964);
xnor U23196 (N_23196,N_22601,N_22875);
and U23197 (N_23197,N_22554,N_22627);
or U23198 (N_23198,N_22633,N_22502);
and U23199 (N_23199,N_22540,N_22647);
nand U23200 (N_23200,N_22913,N_22905);
or U23201 (N_23201,N_22957,N_22507);
or U23202 (N_23202,N_22882,N_22958);
nand U23203 (N_23203,N_22733,N_22926);
nand U23204 (N_23204,N_22798,N_22508);
and U23205 (N_23205,N_22780,N_22827);
or U23206 (N_23206,N_22891,N_22549);
nand U23207 (N_23207,N_22764,N_22757);
xnor U23208 (N_23208,N_22512,N_22597);
nor U23209 (N_23209,N_22773,N_22763);
nor U23210 (N_23210,N_22511,N_22561);
nor U23211 (N_23211,N_22590,N_22698);
and U23212 (N_23212,N_22851,N_22806);
nor U23213 (N_23213,N_22992,N_22849);
xnor U23214 (N_23214,N_22966,N_22665);
nor U23215 (N_23215,N_22902,N_22755);
xnor U23216 (N_23216,N_22861,N_22770);
and U23217 (N_23217,N_22581,N_22651);
nand U23218 (N_23218,N_22814,N_22588);
or U23219 (N_23219,N_22937,N_22705);
nor U23220 (N_23220,N_22793,N_22630);
nand U23221 (N_23221,N_22697,N_22664);
nand U23222 (N_23222,N_22728,N_22822);
nor U23223 (N_23223,N_22928,N_22576);
and U23224 (N_23224,N_22751,N_22514);
nand U23225 (N_23225,N_22694,N_22541);
xnor U23226 (N_23226,N_22589,N_22818);
nor U23227 (N_23227,N_22691,N_22558);
or U23228 (N_23228,N_22523,N_22684);
or U23229 (N_23229,N_22562,N_22617);
nor U23230 (N_23230,N_22848,N_22821);
nor U23231 (N_23231,N_22503,N_22984);
or U23232 (N_23232,N_22812,N_22911);
nand U23233 (N_23233,N_22653,N_22636);
nand U23234 (N_23234,N_22752,N_22978);
xor U23235 (N_23235,N_22872,N_22712);
xnor U23236 (N_23236,N_22999,N_22862);
xor U23237 (N_23237,N_22521,N_22860);
xor U23238 (N_23238,N_22534,N_22518);
nand U23239 (N_23239,N_22690,N_22972);
or U23240 (N_23240,N_22731,N_22708);
and U23241 (N_23241,N_22963,N_22942);
and U23242 (N_23242,N_22775,N_22785);
xnor U23243 (N_23243,N_22837,N_22513);
nor U23244 (N_23244,N_22932,N_22965);
nor U23245 (N_23245,N_22774,N_22758);
or U23246 (N_23246,N_22613,N_22553);
or U23247 (N_23247,N_22604,N_22970);
xor U23248 (N_23248,N_22737,N_22886);
xnor U23249 (N_23249,N_22781,N_22677);
nor U23250 (N_23250,N_22514,N_22646);
nor U23251 (N_23251,N_22563,N_22610);
xnor U23252 (N_23252,N_22736,N_22943);
or U23253 (N_23253,N_22924,N_22591);
nor U23254 (N_23254,N_22696,N_22574);
xnor U23255 (N_23255,N_22949,N_22876);
nand U23256 (N_23256,N_22896,N_22718);
and U23257 (N_23257,N_22785,N_22759);
or U23258 (N_23258,N_22677,N_22618);
nor U23259 (N_23259,N_22971,N_22747);
or U23260 (N_23260,N_22948,N_22544);
xnor U23261 (N_23261,N_22509,N_22672);
and U23262 (N_23262,N_22619,N_22927);
or U23263 (N_23263,N_22634,N_22768);
nand U23264 (N_23264,N_22988,N_22718);
xor U23265 (N_23265,N_22704,N_22922);
nand U23266 (N_23266,N_22542,N_22790);
nand U23267 (N_23267,N_22864,N_22989);
and U23268 (N_23268,N_22948,N_22921);
or U23269 (N_23269,N_22569,N_22969);
and U23270 (N_23270,N_22686,N_22556);
or U23271 (N_23271,N_22651,N_22860);
or U23272 (N_23272,N_22967,N_22898);
nor U23273 (N_23273,N_22813,N_22801);
xor U23274 (N_23274,N_22509,N_22502);
or U23275 (N_23275,N_22738,N_22744);
nand U23276 (N_23276,N_22913,N_22572);
and U23277 (N_23277,N_22649,N_22583);
or U23278 (N_23278,N_22784,N_22778);
nor U23279 (N_23279,N_22637,N_22821);
nor U23280 (N_23280,N_22778,N_22677);
and U23281 (N_23281,N_22855,N_22798);
nand U23282 (N_23282,N_22865,N_22750);
nor U23283 (N_23283,N_22681,N_22651);
nand U23284 (N_23284,N_22853,N_22962);
nand U23285 (N_23285,N_22524,N_22711);
nand U23286 (N_23286,N_22976,N_22908);
or U23287 (N_23287,N_22631,N_22747);
nor U23288 (N_23288,N_22875,N_22703);
nor U23289 (N_23289,N_22840,N_22559);
or U23290 (N_23290,N_22840,N_22685);
xnor U23291 (N_23291,N_22901,N_22755);
nor U23292 (N_23292,N_22605,N_22681);
nor U23293 (N_23293,N_22554,N_22980);
nand U23294 (N_23294,N_22785,N_22680);
and U23295 (N_23295,N_22983,N_22712);
and U23296 (N_23296,N_22500,N_22890);
nand U23297 (N_23297,N_22951,N_22979);
nor U23298 (N_23298,N_22781,N_22510);
or U23299 (N_23299,N_22837,N_22670);
and U23300 (N_23300,N_22555,N_22557);
and U23301 (N_23301,N_22772,N_22691);
xor U23302 (N_23302,N_22894,N_22655);
and U23303 (N_23303,N_22608,N_22991);
and U23304 (N_23304,N_22868,N_22884);
xnor U23305 (N_23305,N_22610,N_22689);
nor U23306 (N_23306,N_22591,N_22595);
xor U23307 (N_23307,N_22683,N_22600);
and U23308 (N_23308,N_22891,N_22821);
nand U23309 (N_23309,N_22718,N_22559);
nor U23310 (N_23310,N_22623,N_22884);
or U23311 (N_23311,N_22581,N_22621);
xor U23312 (N_23312,N_22846,N_22551);
or U23313 (N_23313,N_22619,N_22892);
nor U23314 (N_23314,N_22759,N_22624);
nand U23315 (N_23315,N_22816,N_22689);
nand U23316 (N_23316,N_22966,N_22894);
nor U23317 (N_23317,N_22755,N_22834);
or U23318 (N_23318,N_22615,N_22582);
or U23319 (N_23319,N_22583,N_22691);
or U23320 (N_23320,N_22821,N_22546);
nor U23321 (N_23321,N_22704,N_22808);
xnor U23322 (N_23322,N_22768,N_22833);
xnor U23323 (N_23323,N_22605,N_22507);
nand U23324 (N_23324,N_22791,N_22508);
and U23325 (N_23325,N_22916,N_22806);
nand U23326 (N_23326,N_22948,N_22803);
and U23327 (N_23327,N_22732,N_22918);
xnor U23328 (N_23328,N_22967,N_22789);
xnor U23329 (N_23329,N_22919,N_22874);
or U23330 (N_23330,N_22859,N_22733);
or U23331 (N_23331,N_22940,N_22977);
or U23332 (N_23332,N_22971,N_22655);
and U23333 (N_23333,N_22610,N_22898);
nand U23334 (N_23334,N_22776,N_22857);
nor U23335 (N_23335,N_22826,N_22976);
nand U23336 (N_23336,N_22556,N_22748);
nand U23337 (N_23337,N_22584,N_22665);
nor U23338 (N_23338,N_22838,N_22517);
or U23339 (N_23339,N_22622,N_22792);
nand U23340 (N_23340,N_22965,N_22865);
nor U23341 (N_23341,N_22980,N_22728);
nor U23342 (N_23342,N_22561,N_22856);
nand U23343 (N_23343,N_22946,N_22902);
xor U23344 (N_23344,N_22895,N_22509);
xnor U23345 (N_23345,N_22705,N_22863);
or U23346 (N_23346,N_22917,N_22803);
nand U23347 (N_23347,N_22806,N_22736);
or U23348 (N_23348,N_22828,N_22632);
nand U23349 (N_23349,N_22650,N_22583);
nor U23350 (N_23350,N_22826,N_22555);
xor U23351 (N_23351,N_22911,N_22853);
nor U23352 (N_23352,N_22772,N_22583);
nor U23353 (N_23353,N_22578,N_22612);
nor U23354 (N_23354,N_22572,N_22801);
and U23355 (N_23355,N_22663,N_22930);
nor U23356 (N_23356,N_22894,N_22757);
xor U23357 (N_23357,N_22930,N_22871);
or U23358 (N_23358,N_22753,N_22676);
and U23359 (N_23359,N_22768,N_22958);
nand U23360 (N_23360,N_22986,N_22740);
nor U23361 (N_23361,N_22797,N_22521);
or U23362 (N_23362,N_22801,N_22918);
xor U23363 (N_23363,N_22896,N_22846);
nand U23364 (N_23364,N_22627,N_22987);
xor U23365 (N_23365,N_22732,N_22667);
or U23366 (N_23366,N_22507,N_22561);
and U23367 (N_23367,N_22555,N_22525);
nor U23368 (N_23368,N_22628,N_22910);
xor U23369 (N_23369,N_22920,N_22809);
and U23370 (N_23370,N_22506,N_22743);
nor U23371 (N_23371,N_22638,N_22646);
nand U23372 (N_23372,N_22777,N_22709);
and U23373 (N_23373,N_22786,N_22558);
nand U23374 (N_23374,N_22870,N_22733);
and U23375 (N_23375,N_22895,N_22898);
or U23376 (N_23376,N_22548,N_22825);
nand U23377 (N_23377,N_22899,N_22538);
and U23378 (N_23378,N_22720,N_22518);
xnor U23379 (N_23379,N_22561,N_22873);
nand U23380 (N_23380,N_22882,N_22976);
nor U23381 (N_23381,N_22967,N_22843);
or U23382 (N_23382,N_22939,N_22740);
nand U23383 (N_23383,N_22564,N_22936);
or U23384 (N_23384,N_22524,N_22797);
and U23385 (N_23385,N_22951,N_22739);
or U23386 (N_23386,N_22730,N_22731);
or U23387 (N_23387,N_22549,N_22511);
nand U23388 (N_23388,N_22648,N_22688);
nand U23389 (N_23389,N_22611,N_22755);
nand U23390 (N_23390,N_22896,N_22951);
nand U23391 (N_23391,N_22507,N_22813);
or U23392 (N_23392,N_22751,N_22667);
xor U23393 (N_23393,N_22854,N_22761);
and U23394 (N_23394,N_22526,N_22574);
and U23395 (N_23395,N_22725,N_22966);
or U23396 (N_23396,N_22809,N_22944);
or U23397 (N_23397,N_22669,N_22585);
nand U23398 (N_23398,N_22682,N_22522);
and U23399 (N_23399,N_22739,N_22592);
nor U23400 (N_23400,N_22908,N_22659);
nor U23401 (N_23401,N_22699,N_22590);
nor U23402 (N_23402,N_22827,N_22566);
and U23403 (N_23403,N_22547,N_22647);
or U23404 (N_23404,N_22571,N_22867);
and U23405 (N_23405,N_22940,N_22679);
xor U23406 (N_23406,N_22613,N_22659);
or U23407 (N_23407,N_22813,N_22667);
nand U23408 (N_23408,N_22632,N_22640);
xor U23409 (N_23409,N_22786,N_22956);
and U23410 (N_23410,N_22705,N_22639);
nor U23411 (N_23411,N_22550,N_22845);
nor U23412 (N_23412,N_22658,N_22503);
nor U23413 (N_23413,N_22592,N_22839);
or U23414 (N_23414,N_22829,N_22786);
xor U23415 (N_23415,N_22857,N_22897);
xnor U23416 (N_23416,N_22569,N_22739);
nor U23417 (N_23417,N_22640,N_22760);
nand U23418 (N_23418,N_22650,N_22969);
nand U23419 (N_23419,N_22616,N_22624);
nor U23420 (N_23420,N_22910,N_22725);
nor U23421 (N_23421,N_22706,N_22686);
xnor U23422 (N_23422,N_22819,N_22665);
nand U23423 (N_23423,N_22702,N_22598);
xor U23424 (N_23424,N_22998,N_22671);
nor U23425 (N_23425,N_22613,N_22743);
nor U23426 (N_23426,N_22731,N_22654);
nor U23427 (N_23427,N_22888,N_22943);
and U23428 (N_23428,N_22526,N_22855);
or U23429 (N_23429,N_22561,N_22521);
and U23430 (N_23430,N_22597,N_22727);
xor U23431 (N_23431,N_22924,N_22541);
xnor U23432 (N_23432,N_22701,N_22800);
xnor U23433 (N_23433,N_22738,N_22798);
xnor U23434 (N_23434,N_22819,N_22532);
and U23435 (N_23435,N_22892,N_22814);
and U23436 (N_23436,N_22574,N_22661);
nor U23437 (N_23437,N_22541,N_22848);
nor U23438 (N_23438,N_22899,N_22738);
or U23439 (N_23439,N_22810,N_22756);
nand U23440 (N_23440,N_22932,N_22668);
nor U23441 (N_23441,N_22576,N_22804);
nor U23442 (N_23442,N_22623,N_22967);
and U23443 (N_23443,N_22742,N_22915);
xnor U23444 (N_23444,N_22539,N_22662);
nand U23445 (N_23445,N_22807,N_22968);
nand U23446 (N_23446,N_22900,N_22647);
or U23447 (N_23447,N_22576,N_22577);
nand U23448 (N_23448,N_22537,N_22642);
xor U23449 (N_23449,N_22690,N_22930);
nand U23450 (N_23450,N_22821,N_22631);
or U23451 (N_23451,N_22926,N_22805);
nand U23452 (N_23452,N_22718,N_22585);
nand U23453 (N_23453,N_22892,N_22562);
and U23454 (N_23454,N_22511,N_22582);
nor U23455 (N_23455,N_22911,N_22819);
nor U23456 (N_23456,N_22612,N_22860);
xor U23457 (N_23457,N_22582,N_22882);
nor U23458 (N_23458,N_22712,N_22789);
nor U23459 (N_23459,N_22974,N_22800);
and U23460 (N_23460,N_22871,N_22892);
nor U23461 (N_23461,N_22907,N_22909);
xnor U23462 (N_23462,N_22529,N_22807);
and U23463 (N_23463,N_22905,N_22672);
or U23464 (N_23464,N_22765,N_22762);
and U23465 (N_23465,N_22561,N_22692);
nand U23466 (N_23466,N_22500,N_22522);
or U23467 (N_23467,N_22836,N_22719);
xor U23468 (N_23468,N_22788,N_22995);
xor U23469 (N_23469,N_22512,N_22800);
and U23470 (N_23470,N_22570,N_22738);
or U23471 (N_23471,N_22986,N_22527);
nand U23472 (N_23472,N_22944,N_22956);
nand U23473 (N_23473,N_22595,N_22588);
and U23474 (N_23474,N_22567,N_22876);
nand U23475 (N_23475,N_22660,N_22971);
nand U23476 (N_23476,N_22520,N_22731);
or U23477 (N_23477,N_22741,N_22727);
nand U23478 (N_23478,N_22728,N_22521);
and U23479 (N_23479,N_22782,N_22563);
and U23480 (N_23480,N_22679,N_22521);
or U23481 (N_23481,N_22982,N_22865);
nor U23482 (N_23482,N_22767,N_22641);
and U23483 (N_23483,N_22847,N_22741);
nand U23484 (N_23484,N_22933,N_22864);
nand U23485 (N_23485,N_22715,N_22645);
xnor U23486 (N_23486,N_22648,N_22826);
nand U23487 (N_23487,N_22623,N_22707);
and U23488 (N_23488,N_22838,N_22920);
and U23489 (N_23489,N_22643,N_22657);
xnor U23490 (N_23490,N_22692,N_22873);
or U23491 (N_23491,N_22956,N_22782);
or U23492 (N_23492,N_22880,N_22529);
xnor U23493 (N_23493,N_22852,N_22806);
or U23494 (N_23494,N_22606,N_22839);
xnor U23495 (N_23495,N_22684,N_22708);
or U23496 (N_23496,N_22976,N_22659);
nor U23497 (N_23497,N_22955,N_22607);
nand U23498 (N_23498,N_22591,N_22610);
and U23499 (N_23499,N_22705,N_22743);
nor U23500 (N_23500,N_23385,N_23118);
xnor U23501 (N_23501,N_23192,N_23453);
xnor U23502 (N_23502,N_23282,N_23085);
nand U23503 (N_23503,N_23316,N_23045);
xor U23504 (N_23504,N_23186,N_23163);
nor U23505 (N_23505,N_23059,N_23173);
nor U23506 (N_23506,N_23187,N_23129);
nor U23507 (N_23507,N_23137,N_23180);
nor U23508 (N_23508,N_23367,N_23031);
nand U23509 (N_23509,N_23162,N_23196);
or U23510 (N_23510,N_23165,N_23462);
nor U23511 (N_23511,N_23489,N_23077);
and U23512 (N_23512,N_23238,N_23281);
and U23513 (N_23513,N_23213,N_23407);
nand U23514 (N_23514,N_23363,N_23134);
nor U23515 (N_23515,N_23465,N_23270);
and U23516 (N_23516,N_23368,N_23028);
and U23517 (N_23517,N_23430,N_23008);
xor U23518 (N_23518,N_23132,N_23350);
nor U23519 (N_23519,N_23191,N_23420);
nor U23520 (N_23520,N_23037,N_23354);
and U23521 (N_23521,N_23380,N_23067);
nor U23522 (N_23522,N_23408,N_23386);
and U23523 (N_23523,N_23004,N_23322);
and U23524 (N_23524,N_23349,N_23185);
nand U23525 (N_23525,N_23271,N_23497);
xor U23526 (N_23526,N_23361,N_23161);
or U23527 (N_23527,N_23095,N_23178);
nor U23528 (N_23528,N_23327,N_23246);
and U23529 (N_23529,N_23082,N_23069);
xor U23530 (N_23530,N_23038,N_23343);
nand U23531 (N_23531,N_23306,N_23344);
nand U23532 (N_23532,N_23023,N_23133);
nor U23533 (N_23533,N_23036,N_23445);
nor U23534 (N_23534,N_23240,N_23156);
and U23535 (N_23535,N_23131,N_23402);
xnor U23536 (N_23536,N_23109,N_23202);
or U23537 (N_23537,N_23464,N_23245);
xnor U23538 (N_23538,N_23216,N_23395);
and U23539 (N_23539,N_23140,N_23377);
xnor U23540 (N_23540,N_23406,N_23431);
or U23541 (N_23541,N_23034,N_23040);
nor U23542 (N_23542,N_23397,N_23401);
nor U23543 (N_23543,N_23112,N_23138);
xor U23544 (N_23544,N_23189,N_23257);
nand U23545 (N_23545,N_23084,N_23236);
xnor U23546 (N_23546,N_23154,N_23292);
or U23547 (N_23547,N_23151,N_23164);
nor U23548 (N_23548,N_23381,N_23475);
nor U23549 (N_23549,N_23247,N_23106);
or U23550 (N_23550,N_23107,N_23054);
xor U23551 (N_23551,N_23105,N_23244);
or U23552 (N_23552,N_23002,N_23280);
or U23553 (N_23553,N_23101,N_23288);
xnor U23554 (N_23554,N_23025,N_23451);
and U23555 (N_23555,N_23211,N_23201);
and U23556 (N_23556,N_23048,N_23374);
or U23557 (N_23557,N_23099,N_23452);
and U23558 (N_23558,N_23291,N_23404);
or U23559 (N_23559,N_23320,N_23449);
or U23560 (N_23560,N_23274,N_23114);
xor U23561 (N_23561,N_23339,N_23179);
nor U23562 (N_23562,N_23149,N_23237);
or U23563 (N_23563,N_23362,N_23424);
nand U23564 (N_23564,N_23071,N_23078);
xor U23565 (N_23565,N_23057,N_23460);
xnor U23566 (N_23566,N_23287,N_23195);
xor U23567 (N_23567,N_23220,N_23044);
and U23568 (N_23568,N_23126,N_23455);
xor U23569 (N_23569,N_23313,N_23013);
nor U23570 (N_23570,N_23072,N_23086);
nand U23571 (N_23571,N_23174,N_23064);
nor U23572 (N_23572,N_23074,N_23221);
nor U23573 (N_23573,N_23056,N_23215);
xor U23574 (N_23574,N_23318,N_23442);
xor U23575 (N_23575,N_23136,N_23041);
xnor U23576 (N_23576,N_23169,N_23359);
or U23577 (N_23577,N_23295,N_23243);
and U23578 (N_23578,N_23388,N_23393);
nor U23579 (N_23579,N_23003,N_23047);
xor U23580 (N_23580,N_23482,N_23428);
and U23581 (N_23581,N_23273,N_23448);
nor U23582 (N_23582,N_23263,N_23269);
nor U23583 (N_23583,N_23447,N_23441);
or U23584 (N_23584,N_23224,N_23414);
xor U23585 (N_23585,N_23396,N_23265);
xnor U23586 (N_23586,N_23294,N_23005);
and U23587 (N_23587,N_23300,N_23321);
nand U23588 (N_23588,N_23190,N_23150);
or U23589 (N_23589,N_23128,N_23471);
nand U23590 (N_23590,N_23100,N_23091);
xnor U23591 (N_23591,N_23345,N_23139);
xnor U23592 (N_23592,N_23432,N_23090);
nor U23593 (N_23593,N_23000,N_23039);
nor U23594 (N_23594,N_23060,N_23168);
nand U23595 (N_23595,N_23143,N_23260);
xnor U23596 (N_23596,N_23250,N_23459);
nor U23597 (N_23597,N_23093,N_23252);
xor U23598 (N_23598,N_23022,N_23365);
nand U23599 (N_23599,N_23469,N_23423);
nor U23600 (N_23600,N_23094,N_23089);
and U23601 (N_23601,N_23261,N_23007);
and U23602 (N_23602,N_23239,N_23166);
nor U23603 (N_23603,N_23398,N_23334);
nor U23604 (N_23604,N_23499,N_23487);
nand U23605 (N_23605,N_23417,N_23443);
xnor U23606 (N_23606,N_23116,N_23015);
xnor U23607 (N_23607,N_23314,N_23207);
and U23608 (N_23608,N_23326,N_23217);
nor U23609 (N_23609,N_23457,N_23286);
xor U23610 (N_23610,N_23283,N_23266);
or U23611 (N_23611,N_23026,N_23358);
nor U23612 (N_23612,N_23421,N_23251);
and U23613 (N_23613,N_23272,N_23102);
nor U23614 (N_23614,N_23478,N_23248);
nand U23615 (N_23615,N_23030,N_23389);
nor U23616 (N_23616,N_23279,N_23035);
nand U23617 (N_23617,N_23193,N_23098);
nor U23618 (N_23618,N_23092,N_23223);
xor U23619 (N_23619,N_23172,N_23384);
xor U23620 (N_23620,N_23391,N_23068);
and U23621 (N_23621,N_23419,N_23338);
nand U23622 (N_23622,N_23336,N_23332);
xor U23623 (N_23623,N_23081,N_23214);
nor U23624 (N_23624,N_23016,N_23076);
and U23625 (N_23625,N_23467,N_23160);
or U23626 (N_23626,N_23461,N_23144);
and U23627 (N_23627,N_23230,N_23142);
or U23628 (N_23628,N_23019,N_23141);
xor U23629 (N_23629,N_23222,N_23175);
nand U23630 (N_23630,N_23167,N_23400);
or U23631 (N_23631,N_23063,N_23231);
or U23632 (N_23632,N_23413,N_23337);
nor U23633 (N_23633,N_23331,N_23159);
and U23634 (N_23634,N_23474,N_23333);
nor U23635 (N_23635,N_23120,N_23148);
or U23636 (N_23636,N_23188,N_23328);
nand U23637 (N_23637,N_23278,N_23050);
nand U23638 (N_23638,N_23297,N_23394);
or U23639 (N_23639,N_23470,N_23021);
xnor U23640 (N_23640,N_23229,N_23051);
xor U23641 (N_23641,N_23110,N_23479);
or U23642 (N_23642,N_23360,N_23152);
nor U23643 (N_23643,N_23147,N_23371);
nand U23644 (N_23644,N_23204,N_23418);
nand U23645 (N_23645,N_23476,N_23198);
nand U23646 (N_23646,N_23483,N_23249);
nand U23647 (N_23647,N_23104,N_23234);
nand U23648 (N_23648,N_23171,N_23427);
and U23649 (N_23649,N_23289,N_23258);
xnor U23650 (N_23650,N_23058,N_23182);
and U23651 (N_23651,N_23032,N_23267);
xnor U23652 (N_23652,N_23262,N_23477);
xor U23653 (N_23653,N_23315,N_23364);
nand U23654 (N_23654,N_23219,N_23450);
nor U23655 (N_23655,N_23387,N_23111);
or U23656 (N_23656,N_23061,N_23438);
nor U23657 (N_23657,N_23435,N_23307);
xnor U23658 (N_23658,N_23075,N_23153);
xor U23659 (N_23659,N_23181,N_23422);
nor U23660 (N_23660,N_23301,N_23115);
xor U23661 (N_23661,N_23199,N_23484);
or U23662 (N_23662,N_23323,N_23018);
xnor U23663 (N_23663,N_23200,N_23355);
nand U23664 (N_23664,N_23255,N_23225);
nor U23665 (N_23665,N_23342,N_23205);
and U23666 (N_23666,N_23042,N_23227);
nor U23667 (N_23667,N_23472,N_23403);
nand U23668 (N_23668,N_23065,N_23329);
and U23669 (N_23669,N_23382,N_23122);
and U23670 (N_23670,N_23308,N_23488);
nand U23671 (N_23671,N_23259,N_23378);
or U23672 (N_23672,N_23212,N_23351);
or U23673 (N_23673,N_23241,N_23296);
nand U23674 (N_23674,N_23001,N_23463);
and U23675 (N_23675,N_23194,N_23073);
xnor U23676 (N_23676,N_23029,N_23020);
nor U23677 (N_23677,N_23305,N_23302);
nor U23678 (N_23678,N_23303,N_23325);
xor U23679 (N_23679,N_23197,N_23330);
and U23680 (N_23680,N_23373,N_23498);
xnor U23681 (N_23681,N_23357,N_23304);
and U23682 (N_23682,N_23145,N_23097);
or U23683 (N_23683,N_23379,N_23285);
xnor U23684 (N_23684,N_23411,N_23226);
or U23685 (N_23685,N_23083,N_23006);
xnor U23686 (N_23686,N_23087,N_23233);
nor U23687 (N_23687,N_23235,N_23473);
or U23688 (N_23688,N_23317,N_23412);
xor U23689 (N_23689,N_23079,N_23121);
and U23690 (N_23690,N_23046,N_23372);
xnor U23691 (N_23691,N_23218,N_23480);
and U23692 (N_23692,N_23176,N_23298);
and U23693 (N_23693,N_23203,N_23375);
and U23694 (N_23694,N_23492,N_23390);
xnor U23695 (N_23695,N_23158,N_23127);
nand U23696 (N_23696,N_23275,N_23184);
xor U23697 (N_23697,N_23446,N_23440);
nor U23698 (N_23698,N_23009,N_23495);
and U23699 (N_23699,N_23253,N_23494);
xnor U23700 (N_23700,N_23155,N_23399);
and U23701 (N_23701,N_23410,N_23309);
nor U23702 (N_23702,N_23299,N_23206);
nand U23703 (N_23703,N_23405,N_23392);
xor U23704 (N_23704,N_23012,N_23183);
and U23705 (N_23705,N_23366,N_23014);
nor U23706 (N_23706,N_23177,N_23070);
nor U23707 (N_23707,N_23466,N_23210);
nor U23708 (N_23708,N_23256,N_23346);
nor U23709 (N_23709,N_23103,N_23146);
and U23710 (N_23710,N_23080,N_23055);
nor U23711 (N_23711,N_23415,N_23268);
nand U23712 (N_23712,N_23348,N_23439);
xnor U23713 (N_23713,N_23437,N_23383);
or U23714 (N_23714,N_23311,N_23335);
xnor U23715 (N_23715,N_23456,N_23376);
nand U23716 (N_23716,N_23444,N_23228);
or U23717 (N_23717,N_23496,N_23356);
or U23718 (N_23718,N_23347,N_23324);
nor U23719 (N_23719,N_23033,N_23277);
nor U23720 (N_23720,N_23157,N_23353);
nand U23721 (N_23721,N_23108,N_23319);
or U23722 (N_23722,N_23486,N_23052);
or U23723 (N_23723,N_23066,N_23242);
nand U23724 (N_23724,N_23254,N_23468);
nor U23725 (N_23725,N_23130,N_23209);
nor U23726 (N_23726,N_23124,N_23370);
nand U23727 (N_23727,N_23049,N_23088);
and U23728 (N_23728,N_23096,N_23312);
and U23729 (N_23729,N_23436,N_23011);
and U23730 (N_23730,N_23341,N_23017);
nor U23731 (N_23731,N_23493,N_23416);
nand U23732 (N_23732,N_23433,N_23491);
and U23733 (N_23733,N_23135,N_23290);
xnor U23734 (N_23734,N_23352,N_23208);
xnor U23735 (N_23735,N_23232,N_23284);
xnor U23736 (N_23736,N_23276,N_23043);
nor U23737 (N_23737,N_23429,N_23113);
or U23738 (N_23738,N_23454,N_23010);
or U23739 (N_23739,N_23434,N_23125);
and U23740 (N_23740,N_23117,N_23485);
nor U23741 (N_23741,N_23053,N_23481);
or U23742 (N_23742,N_23024,N_23027);
and U23743 (N_23743,N_23264,N_23123);
xor U23744 (N_23744,N_23425,N_23340);
xnor U23745 (N_23745,N_23426,N_23119);
xor U23746 (N_23746,N_23293,N_23170);
nand U23747 (N_23747,N_23409,N_23310);
xnor U23748 (N_23748,N_23369,N_23062);
nor U23749 (N_23749,N_23490,N_23458);
xnor U23750 (N_23750,N_23008,N_23390);
or U23751 (N_23751,N_23155,N_23148);
xor U23752 (N_23752,N_23459,N_23298);
nor U23753 (N_23753,N_23324,N_23278);
nor U23754 (N_23754,N_23082,N_23007);
xnor U23755 (N_23755,N_23276,N_23434);
nand U23756 (N_23756,N_23195,N_23143);
nand U23757 (N_23757,N_23038,N_23033);
or U23758 (N_23758,N_23197,N_23084);
nand U23759 (N_23759,N_23485,N_23180);
xnor U23760 (N_23760,N_23085,N_23348);
xor U23761 (N_23761,N_23412,N_23063);
nand U23762 (N_23762,N_23136,N_23106);
nand U23763 (N_23763,N_23092,N_23125);
or U23764 (N_23764,N_23089,N_23116);
or U23765 (N_23765,N_23044,N_23270);
and U23766 (N_23766,N_23069,N_23185);
nand U23767 (N_23767,N_23028,N_23190);
and U23768 (N_23768,N_23399,N_23313);
or U23769 (N_23769,N_23102,N_23367);
nor U23770 (N_23770,N_23020,N_23108);
nand U23771 (N_23771,N_23435,N_23308);
or U23772 (N_23772,N_23019,N_23339);
nand U23773 (N_23773,N_23211,N_23457);
or U23774 (N_23774,N_23366,N_23353);
nor U23775 (N_23775,N_23139,N_23056);
xnor U23776 (N_23776,N_23241,N_23124);
and U23777 (N_23777,N_23278,N_23193);
and U23778 (N_23778,N_23280,N_23377);
xor U23779 (N_23779,N_23017,N_23095);
and U23780 (N_23780,N_23162,N_23157);
xor U23781 (N_23781,N_23404,N_23330);
nor U23782 (N_23782,N_23303,N_23096);
nand U23783 (N_23783,N_23356,N_23274);
nand U23784 (N_23784,N_23137,N_23272);
xor U23785 (N_23785,N_23442,N_23195);
xnor U23786 (N_23786,N_23198,N_23083);
xor U23787 (N_23787,N_23197,N_23209);
nand U23788 (N_23788,N_23450,N_23496);
or U23789 (N_23789,N_23038,N_23308);
or U23790 (N_23790,N_23411,N_23498);
or U23791 (N_23791,N_23060,N_23030);
and U23792 (N_23792,N_23239,N_23082);
nand U23793 (N_23793,N_23153,N_23113);
and U23794 (N_23794,N_23447,N_23393);
or U23795 (N_23795,N_23443,N_23397);
xor U23796 (N_23796,N_23234,N_23383);
nand U23797 (N_23797,N_23069,N_23413);
nand U23798 (N_23798,N_23016,N_23185);
nor U23799 (N_23799,N_23229,N_23405);
nor U23800 (N_23800,N_23230,N_23431);
or U23801 (N_23801,N_23112,N_23221);
or U23802 (N_23802,N_23198,N_23365);
or U23803 (N_23803,N_23045,N_23404);
xor U23804 (N_23804,N_23020,N_23145);
nand U23805 (N_23805,N_23439,N_23005);
and U23806 (N_23806,N_23196,N_23287);
or U23807 (N_23807,N_23335,N_23355);
xnor U23808 (N_23808,N_23096,N_23268);
and U23809 (N_23809,N_23469,N_23162);
or U23810 (N_23810,N_23205,N_23038);
and U23811 (N_23811,N_23493,N_23496);
nand U23812 (N_23812,N_23469,N_23167);
nand U23813 (N_23813,N_23457,N_23363);
or U23814 (N_23814,N_23305,N_23343);
xor U23815 (N_23815,N_23036,N_23025);
xnor U23816 (N_23816,N_23214,N_23390);
xnor U23817 (N_23817,N_23391,N_23334);
or U23818 (N_23818,N_23285,N_23295);
nor U23819 (N_23819,N_23208,N_23126);
nand U23820 (N_23820,N_23363,N_23246);
nand U23821 (N_23821,N_23119,N_23087);
nand U23822 (N_23822,N_23076,N_23209);
or U23823 (N_23823,N_23013,N_23010);
nor U23824 (N_23824,N_23085,N_23290);
or U23825 (N_23825,N_23488,N_23002);
or U23826 (N_23826,N_23046,N_23166);
nand U23827 (N_23827,N_23022,N_23158);
nand U23828 (N_23828,N_23254,N_23312);
nor U23829 (N_23829,N_23421,N_23460);
nand U23830 (N_23830,N_23255,N_23252);
nor U23831 (N_23831,N_23094,N_23113);
nand U23832 (N_23832,N_23284,N_23342);
nor U23833 (N_23833,N_23059,N_23240);
xnor U23834 (N_23834,N_23116,N_23190);
or U23835 (N_23835,N_23226,N_23147);
nor U23836 (N_23836,N_23133,N_23204);
nor U23837 (N_23837,N_23056,N_23455);
nand U23838 (N_23838,N_23196,N_23209);
xor U23839 (N_23839,N_23367,N_23157);
nor U23840 (N_23840,N_23370,N_23123);
and U23841 (N_23841,N_23227,N_23010);
nand U23842 (N_23842,N_23412,N_23329);
nand U23843 (N_23843,N_23167,N_23188);
nor U23844 (N_23844,N_23044,N_23370);
nand U23845 (N_23845,N_23008,N_23278);
nor U23846 (N_23846,N_23107,N_23376);
nor U23847 (N_23847,N_23017,N_23440);
and U23848 (N_23848,N_23397,N_23208);
and U23849 (N_23849,N_23327,N_23384);
nor U23850 (N_23850,N_23227,N_23162);
and U23851 (N_23851,N_23214,N_23305);
nor U23852 (N_23852,N_23313,N_23238);
and U23853 (N_23853,N_23273,N_23161);
xnor U23854 (N_23854,N_23242,N_23229);
xor U23855 (N_23855,N_23329,N_23472);
or U23856 (N_23856,N_23315,N_23060);
or U23857 (N_23857,N_23012,N_23077);
and U23858 (N_23858,N_23032,N_23455);
or U23859 (N_23859,N_23292,N_23419);
nand U23860 (N_23860,N_23482,N_23111);
xor U23861 (N_23861,N_23151,N_23133);
xnor U23862 (N_23862,N_23357,N_23241);
and U23863 (N_23863,N_23303,N_23354);
nand U23864 (N_23864,N_23163,N_23254);
nor U23865 (N_23865,N_23044,N_23254);
xnor U23866 (N_23866,N_23243,N_23083);
and U23867 (N_23867,N_23400,N_23334);
xnor U23868 (N_23868,N_23450,N_23029);
and U23869 (N_23869,N_23492,N_23142);
or U23870 (N_23870,N_23139,N_23318);
nor U23871 (N_23871,N_23478,N_23427);
and U23872 (N_23872,N_23269,N_23052);
xor U23873 (N_23873,N_23372,N_23248);
nor U23874 (N_23874,N_23054,N_23477);
nand U23875 (N_23875,N_23151,N_23055);
xnor U23876 (N_23876,N_23456,N_23125);
nand U23877 (N_23877,N_23214,N_23226);
or U23878 (N_23878,N_23220,N_23418);
nand U23879 (N_23879,N_23082,N_23210);
xor U23880 (N_23880,N_23335,N_23173);
xor U23881 (N_23881,N_23262,N_23446);
nor U23882 (N_23882,N_23273,N_23291);
and U23883 (N_23883,N_23360,N_23055);
nor U23884 (N_23884,N_23148,N_23444);
and U23885 (N_23885,N_23009,N_23319);
or U23886 (N_23886,N_23093,N_23048);
nand U23887 (N_23887,N_23127,N_23384);
xor U23888 (N_23888,N_23308,N_23372);
or U23889 (N_23889,N_23228,N_23299);
and U23890 (N_23890,N_23266,N_23216);
nor U23891 (N_23891,N_23455,N_23333);
or U23892 (N_23892,N_23137,N_23003);
nor U23893 (N_23893,N_23147,N_23413);
nor U23894 (N_23894,N_23040,N_23344);
or U23895 (N_23895,N_23021,N_23396);
nand U23896 (N_23896,N_23409,N_23053);
nand U23897 (N_23897,N_23040,N_23127);
nor U23898 (N_23898,N_23200,N_23287);
nor U23899 (N_23899,N_23244,N_23493);
xnor U23900 (N_23900,N_23323,N_23082);
nand U23901 (N_23901,N_23402,N_23042);
xor U23902 (N_23902,N_23225,N_23027);
nand U23903 (N_23903,N_23070,N_23223);
nor U23904 (N_23904,N_23265,N_23159);
xor U23905 (N_23905,N_23054,N_23403);
xnor U23906 (N_23906,N_23262,N_23097);
nand U23907 (N_23907,N_23191,N_23124);
and U23908 (N_23908,N_23332,N_23147);
nand U23909 (N_23909,N_23488,N_23380);
xor U23910 (N_23910,N_23221,N_23452);
xnor U23911 (N_23911,N_23124,N_23089);
nand U23912 (N_23912,N_23480,N_23295);
xnor U23913 (N_23913,N_23177,N_23366);
nand U23914 (N_23914,N_23184,N_23377);
nand U23915 (N_23915,N_23455,N_23148);
xor U23916 (N_23916,N_23470,N_23358);
or U23917 (N_23917,N_23065,N_23323);
and U23918 (N_23918,N_23304,N_23487);
nand U23919 (N_23919,N_23145,N_23340);
and U23920 (N_23920,N_23382,N_23295);
and U23921 (N_23921,N_23314,N_23029);
or U23922 (N_23922,N_23143,N_23436);
and U23923 (N_23923,N_23277,N_23268);
nor U23924 (N_23924,N_23177,N_23099);
or U23925 (N_23925,N_23091,N_23027);
and U23926 (N_23926,N_23199,N_23083);
xnor U23927 (N_23927,N_23400,N_23289);
xor U23928 (N_23928,N_23346,N_23133);
nand U23929 (N_23929,N_23427,N_23351);
nand U23930 (N_23930,N_23194,N_23217);
xor U23931 (N_23931,N_23325,N_23300);
and U23932 (N_23932,N_23025,N_23082);
nor U23933 (N_23933,N_23075,N_23156);
xnor U23934 (N_23934,N_23169,N_23313);
nand U23935 (N_23935,N_23201,N_23370);
and U23936 (N_23936,N_23079,N_23090);
or U23937 (N_23937,N_23461,N_23229);
xnor U23938 (N_23938,N_23011,N_23218);
nor U23939 (N_23939,N_23020,N_23093);
or U23940 (N_23940,N_23352,N_23271);
nand U23941 (N_23941,N_23427,N_23275);
nand U23942 (N_23942,N_23146,N_23133);
nand U23943 (N_23943,N_23077,N_23470);
or U23944 (N_23944,N_23309,N_23384);
and U23945 (N_23945,N_23299,N_23499);
or U23946 (N_23946,N_23012,N_23133);
xnor U23947 (N_23947,N_23090,N_23450);
xnor U23948 (N_23948,N_23391,N_23344);
or U23949 (N_23949,N_23236,N_23009);
and U23950 (N_23950,N_23430,N_23255);
nor U23951 (N_23951,N_23121,N_23093);
and U23952 (N_23952,N_23444,N_23445);
or U23953 (N_23953,N_23430,N_23143);
or U23954 (N_23954,N_23363,N_23178);
and U23955 (N_23955,N_23296,N_23325);
nand U23956 (N_23956,N_23486,N_23369);
nor U23957 (N_23957,N_23352,N_23209);
nand U23958 (N_23958,N_23391,N_23325);
and U23959 (N_23959,N_23387,N_23219);
nor U23960 (N_23960,N_23158,N_23067);
nor U23961 (N_23961,N_23099,N_23208);
and U23962 (N_23962,N_23452,N_23079);
nand U23963 (N_23963,N_23134,N_23150);
nand U23964 (N_23964,N_23475,N_23387);
xor U23965 (N_23965,N_23356,N_23140);
nand U23966 (N_23966,N_23390,N_23382);
nand U23967 (N_23967,N_23347,N_23421);
and U23968 (N_23968,N_23004,N_23453);
and U23969 (N_23969,N_23263,N_23187);
xnor U23970 (N_23970,N_23202,N_23331);
nor U23971 (N_23971,N_23034,N_23005);
xor U23972 (N_23972,N_23050,N_23100);
nand U23973 (N_23973,N_23362,N_23110);
xor U23974 (N_23974,N_23255,N_23385);
and U23975 (N_23975,N_23253,N_23479);
and U23976 (N_23976,N_23422,N_23168);
nor U23977 (N_23977,N_23415,N_23222);
nand U23978 (N_23978,N_23230,N_23235);
nand U23979 (N_23979,N_23139,N_23337);
nand U23980 (N_23980,N_23091,N_23076);
or U23981 (N_23981,N_23054,N_23349);
or U23982 (N_23982,N_23142,N_23052);
and U23983 (N_23983,N_23458,N_23287);
and U23984 (N_23984,N_23272,N_23114);
nor U23985 (N_23985,N_23357,N_23153);
nor U23986 (N_23986,N_23255,N_23017);
or U23987 (N_23987,N_23480,N_23238);
nor U23988 (N_23988,N_23032,N_23288);
xor U23989 (N_23989,N_23420,N_23395);
xnor U23990 (N_23990,N_23322,N_23016);
xor U23991 (N_23991,N_23199,N_23320);
nor U23992 (N_23992,N_23176,N_23393);
and U23993 (N_23993,N_23294,N_23388);
nor U23994 (N_23994,N_23006,N_23488);
nor U23995 (N_23995,N_23212,N_23110);
and U23996 (N_23996,N_23194,N_23413);
nor U23997 (N_23997,N_23017,N_23231);
nand U23998 (N_23998,N_23224,N_23076);
or U23999 (N_23999,N_23083,N_23355);
nand U24000 (N_24000,N_23969,N_23535);
or U24001 (N_24001,N_23665,N_23864);
nand U24002 (N_24002,N_23915,N_23580);
nor U24003 (N_24003,N_23690,N_23532);
xnor U24004 (N_24004,N_23845,N_23642);
nor U24005 (N_24005,N_23918,N_23954);
and U24006 (N_24006,N_23601,N_23741);
and U24007 (N_24007,N_23659,N_23545);
or U24008 (N_24008,N_23970,N_23671);
or U24009 (N_24009,N_23655,N_23895);
or U24010 (N_24010,N_23920,N_23966);
nor U24011 (N_24011,N_23861,N_23809);
and U24012 (N_24012,N_23544,N_23981);
xnor U24013 (N_24013,N_23960,N_23764);
nand U24014 (N_24014,N_23579,N_23967);
xor U24015 (N_24015,N_23590,N_23843);
nor U24016 (N_24016,N_23592,N_23801);
xnor U24017 (N_24017,N_23924,N_23982);
nor U24018 (N_24018,N_23605,N_23974);
or U24019 (N_24019,N_23501,N_23702);
xnor U24020 (N_24020,N_23778,N_23834);
or U24021 (N_24021,N_23567,N_23968);
or U24022 (N_24022,N_23693,N_23546);
nor U24023 (N_24023,N_23957,N_23562);
or U24024 (N_24024,N_23746,N_23927);
or U24025 (N_24025,N_23743,N_23850);
and U24026 (N_24026,N_23514,N_23761);
nor U24027 (N_24027,N_23903,N_23612);
xor U24028 (N_24028,N_23561,N_23696);
nor U24029 (N_24029,N_23963,N_23638);
and U24030 (N_24030,N_23507,N_23557);
xnor U24031 (N_24031,N_23653,N_23713);
nor U24032 (N_24032,N_23932,N_23961);
or U24033 (N_24033,N_23921,N_23904);
nor U24034 (N_24034,N_23737,N_23839);
xor U24035 (N_24035,N_23600,N_23805);
xnor U24036 (N_24036,N_23931,N_23807);
nand U24037 (N_24037,N_23623,N_23523);
or U24038 (N_24038,N_23979,N_23525);
nand U24039 (N_24039,N_23799,N_23657);
or U24040 (N_24040,N_23571,N_23621);
xnor U24041 (N_24041,N_23858,N_23747);
nand U24042 (N_24042,N_23710,N_23650);
xor U24043 (N_24043,N_23964,N_23875);
nor U24044 (N_24044,N_23832,N_23877);
nor U24045 (N_24045,N_23842,N_23991);
nand U24046 (N_24046,N_23824,N_23660);
nand U24047 (N_24047,N_23643,N_23733);
and U24048 (N_24048,N_23700,N_23548);
nand U24049 (N_24049,N_23999,N_23817);
nand U24050 (N_24050,N_23632,N_23563);
nand U24051 (N_24051,N_23663,N_23553);
nor U24052 (N_24052,N_23588,N_23706);
xnor U24053 (N_24053,N_23698,N_23854);
or U24054 (N_24054,N_23517,N_23773);
or U24055 (N_24055,N_23995,N_23729);
nor U24056 (N_24056,N_23512,N_23962);
nor U24057 (N_24057,N_23528,N_23855);
nand U24058 (N_24058,N_23917,N_23822);
nand U24059 (N_24059,N_23504,N_23891);
nand U24060 (N_24060,N_23593,N_23651);
and U24061 (N_24061,N_23851,N_23724);
nor U24062 (N_24062,N_23583,N_23753);
nor U24063 (N_24063,N_23763,N_23505);
or U24064 (N_24064,N_23806,N_23811);
nor U24065 (N_24065,N_23831,N_23661);
or U24066 (N_24066,N_23998,N_23866);
nand U24067 (N_24067,N_23797,N_23620);
nand U24068 (N_24068,N_23727,N_23862);
and U24069 (N_24069,N_23871,N_23765);
and U24070 (N_24070,N_23630,N_23758);
or U24071 (N_24071,N_23644,N_23551);
nor U24072 (N_24072,N_23719,N_23547);
nand U24073 (N_24073,N_23827,N_23609);
nor U24074 (N_24074,N_23518,N_23914);
or U24075 (N_24075,N_23886,N_23752);
and U24076 (N_24076,N_23716,N_23956);
nor U24077 (N_24077,N_23565,N_23513);
nand U24078 (N_24078,N_23876,N_23925);
nor U24079 (N_24079,N_23977,N_23935);
nor U24080 (N_24080,N_23691,N_23989);
and U24081 (N_24081,N_23826,N_23516);
xor U24082 (N_24082,N_23508,N_23581);
nor U24083 (N_24083,N_23755,N_23971);
and U24084 (N_24084,N_23736,N_23742);
or U24085 (N_24085,N_23537,N_23684);
nand U24086 (N_24086,N_23669,N_23933);
nand U24087 (N_24087,N_23534,N_23550);
nor U24088 (N_24088,N_23522,N_23772);
xnor U24089 (N_24089,N_23686,N_23930);
nor U24090 (N_24090,N_23515,N_23756);
xnor U24091 (N_24091,N_23636,N_23846);
nor U24092 (N_24092,N_23622,N_23538);
xor U24093 (N_24093,N_23893,N_23506);
nor U24094 (N_24094,N_23952,N_23734);
nor U24095 (N_24095,N_23800,N_23986);
nor U24096 (N_24096,N_23649,N_23709);
or U24097 (N_24097,N_23785,N_23882);
or U24098 (N_24098,N_23591,N_23944);
and U24099 (N_24099,N_23595,N_23788);
nand U24100 (N_24100,N_23558,N_23692);
and U24101 (N_24101,N_23992,N_23808);
nand U24102 (N_24102,N_23770,N_23828);
xor U24103 (N_24103,N_23802,N_23783);
nand U24104 (N_24104,N_23880,N_23840);
and U24105 (N_24105,N_23934,N_23972);
nand U24106 (N_24106,N_23889,N_23714);
or U24107 (N_24107,N_23735,N_23870);
or U24108 (N_24108,N_23697,N_23767);
nor U24109 (N_24109,N_23844,N_23946);
xor U24110 (N_24110,N_23695,N_23884);
xor U24111 (N_24111,N_23949,N_23509);
and U24112 (N_24112,N_23611,N_23524);
xnor U24113 (N_24113,N_23645,N_23586);
or U24114 (N_24114,N_23725,N_23577);
and U24115 (N_24115,N_23652,N_23941);
and U24116 (N_24116,N_23674,N_23835);
or U24117 (N_24117,N_23955,N_23582);
or U24118 (N_24118,N_23721,N_23994);
xor U24119 (N_24119,N_23887,N_23527);
xnor U24120 (N_24120,N_23744,N_23899);
xor U24121 (N_24121,N_23879,N_23973);
nor U24122 (N_24122,N_23614,N_23984);
or U24123 (N_24123,N_23782,N_23570);
nand U24124 (N_24124,N_23720,N_23503);
or U24125 (N_24125,N_23739,N_23993);
nor U24126 (N_24126,N_23618,N_23656);
or U24127 (N_24127,N_23607,N_23678);
and U24128 (N_24128,N_23852,N_23740);
xnor U24129 (N_24129,N_23819,N_23745);
nor U24130 (N_24130,N_23694,N_23860);
nor U24131 (N_24131,N_23911,N_23908);
and U24132 (N_24132,N_23947,N_23901);
nand U24133 (N_24133,N_23667,N_23816);
and U24134 (N_24134,N_23682,N_23726);
and U24135 (N_24135,N_23502,N_23705);
nand U24136 (N_24136,N_23602,N_23732);
or U24137 (N_24137,N_23731,N_23784);
nand U24138 (N_24138,N_23634,N_23648);
nor U24139 (N_24139,N_23637,N_23707);
nand U24140 (N_24140,N_23730,N_23794);
nor U24141 (N_24141,N_23874,N_23987);
and U24142 (N_24142,N_23578,N_23939);
nand U24143 (N_24143,N_23781,N_23780);
nand U24144 (N_24144,N_23728,N_23938);
nor U24145 (N_24145,N_23883,N_23530);
nor U24146 (N_24146,N_23500,N_23658);
nand U24147 (N_24147,N_23815,N_23814);
nor U24148 (N_24148,N_23774,N_23959);
nand U24149 (N_24149,N_23672,N_23608);
or U24150 (N_24150,N_23937,N_23873);
xnor U24151 (N_24151,N_23790,N_23519);
nor U24152 (N_24152,N_23775,N_23897);
nor U24153 (N_24153,N_23813,N_23627);
xnor U24154 (N_24154,N_23894,N_23666);
or U24155 (N_24155,N_23615,N_23520);
nand U24156 (N_24156,N_23791,N_23679);
nor U24157 (N_24157,N_23521,N_23923);
nor U24158 (N_24158,N_23596,N_23597);
nor U24159 (N_24159,N_23685,N_23942);
or U24160 (N_24160,N_23631,N_23531);
or U24161 (N_24161,N_23549,N_23857);
and U24162 (N_24162,N_23635,N_23760);
nand U24163 (N_24163,N_23625,N_23610);
nand U24164 (N_24164,N_23922,N_23829);
or U24165 (N_24165,N_23867,N_23865);
or U24166 (N_24166,N_23640,N_23511);
and U24167 (N_24167,N_23759,N_23795);
xnor U24168 (N_24168,N_23560,N_23681);
or U24169 (N_24169,N_23606,N_23830);
or U24170 (N_24170,N_23976,N_23950);
nand U24171 (N_24171,N_23769,N_23670);
and U24172 (N_24172,N_23892,N_23568);
xnor U24173 (N_24173,N_23738,N_23985);
xor U24174 (N_24174,N_23863,N_23668);
nor U24175 (N_24175,N_23569,N_23540);
or U24176 (N_24176,N_23587,N_23572);
nor U24177 (N_24177,N_23566,N_23542);
xnor U24178 (N_24178,N_23945,N_23613);
and U24179 (N_24179,N_23617,N_23552);
or U24180 (N_24180,N_23654,N_23902);
or U24181 (N_24181,N_23900,N_23878);
xnor U24182 (N_24182,N_23750,N_23754);
or U24183 (N_24183,N_23885,N_23526);
nor U24184 (N_24184,N_23820,N_23712);
xnor U24185 (N_24185,N_23633,N_23536);
nand U24186 (N_24186,N_23766,N_23912);
and U24187 (N_24187,N_23529,N_23890);
and U24188 (N_24188,N_23818,N_23916);
xnor U24189 (N_24189,N_23787,N_23929);
nand U24190 (N_24190,N_23810,N_23677);
xor U24191 (N_24191,N_23599,N_23803);
nand U24192 (N_24192,N_23905,N_23604);
xnor U24193 (N_24193,N_23965,N_23943);
nand U24194 (N_24194,N_23837,N_23913);
nor U24195 (N_24195,N_23958,N_23928);
or U24196 (N_24196,N_23848,N_23624);
nand U24197 (N_24197,N_23589,N_23626);
and U24198 (N_24198,N_23988,N_23825);
nand U24199 (N_24199,N_23792,N_23539);
nand U24200 (N_24200,N_23639,N_23510);
and U24201 (N_24201,N_23821,N_23748);
and U24202 (N_24202,N_23833,N_23662);
nor U24203 (N_24203,N_23708,N_23849);
xnor U24204 (N_24204,N_23898,N_23704);
and U24205 (N_24205,N_23907,N_23575);
nor U24206 (N_24206,N_23715,N_23990);
nand U24207 (N_24207,N_23953,N_23836);
xor U24208 (N_24208,N_23762,N_23554);
nor U24209 (N_24209,N_23859,N_23838);
xor U24210 (N_24210,N_23688,N_23676);
and U24211 (N_24211,N_23948,N_23975);
nand U24212 (N_24212,N_23768,N_23680);
or U24213 (N_24213,N_23646,N_23598);
xor U24214 (N_24214,N_23779,N_23823);
or U24215 (N_24215,N_23798,N_23980);
nand U24216 (N_24216,N_23919,N_23703);
nor U24217 (N_24217,N_23564,N_23576);
nand U24218 (N_24218,N_23776,N_23717);
and U24219 (N_24219,N_23749,N_23628);
and U24220 (N_24220,N_23793,N_23556);
nand U24221 (N_24221,N_23603,N_23853);
xnor U24222 (N_24222,N_23629,N_23584);
xnor U24223 (N_24223,N_23574,N_23847);
nand U24224 (N_24224,N_23812,N_23841);
nor U24225 (N_24225,N_23868,N_23910);
nand U24226 (N_24226,N_23997,N_23573);
nor U24227 (N_24227,N_23906,N_23647);
nand U24228 (N_24228,N_23616,N_23664);
xor U24229 (N_24229,N_23701,N_23909);
nand U24230 (N_24230,N_23543,N_23896);
and U24231 (N_24231,N_23711,N_23751);
or U24232 (N_24232,N_23789,N_23699);
nand U24233 (N_24233,N_23983,N_23978);
xnor U24234 (N_24234,N_23722,N_23926);
and U24235 (N_24235,N_23619,N_23541);
xnor U24236 (N_24236,N_23951,N_23555);
or U24237 (N_24237,N_23796,N_23533);
xnor U24238 (N_24238,N_23771,N_23673);
nor U24239 (N_24239,N_23777,N_23675);
nor U24240 (N_24240,N_23888,N_23757);
nor U24241 (N_24241,N_23996,N_23687);
xnor U24242 (N_24242,N_23940,N_23804);
or U24243 (N_24243,N_23723,N_23936);
nand U24244 (N_24244,N_23594,N_23641);
xnor U24245 (N_24245,N_23786,N_23881);
nor U24246 (N_24246,N_23689,N_23559);
xnor U24247 (N_24247,N_23856,N_23585);
nor U24248 (N_24248,N_23718,N_23683);
or U24249 (N_24249,N_23869,N_23872);
or U24250 (N_24250,N_23546,N_23682);
nand U24251 (N_24251,N_23715,N_23982);
nand U24252 (N_24252,N_23558,N_23507);
and U24253 (N_24253,N_23587,N_23671);
xnor U24254 (N_24254,N_23550,N_23716);
and U24255 (N_24255,N_23546,N_23771);
nand U24256 (N_24256,N_23934,N_23541);
or U24257 (N_24257,N_23533,N_23504);
nand U24258 (N_24258,N_23964,N_23600);
and U24259 (N_24259,N_23683,N_23807);
nand U24260 (N_24260,N_23569,N_23526);
and U24261 (N_24261,N_23758,N_23822);
nand U24262 (N_24262,N_23886,N_23711);
nand U24263 (N_24263,N_23541,N_23545);
or U24264 (N_24264,N_23730,N_23550);
and U24265 (N_24265,N_23507,N_23941);
and U24266 (N_24266,N_23803,N_23557);
nand U24267 (N_24267,N_23657,N_23509);
and U24268 (N_24268,N_23505,N_23823);
or U24269 (N_24269,N_23579,N_23667);
nand U24270 (N_24270,N_23945,N_23777);
xnor U24271 (N_24271,N_23738,N_23577);
and U24272 (N_24272,N_23911,N_23783);
and U24273 (N_24273,N_23538,N_23951);
xor U24274 (N_24274,N_23685,N_23994);
and U24275 (N_24275,N_23549,N_23589);
or U24276 (N_24276,N_23714,N_23802);
or U24277 (N_24277,N_23919,N_23779);
nor U24278 (N_24278,N_23979,N_23688);
or U24279 (N_24279,N_23622,N_23928);
nor U24280 (N_24280,N_23898,N_23627);
and U24281 (N_24281,N_23932,N_23551);
xnor U24282 (N_24282,N_23865,N_23576);
or U24283 (N_24283,N_23783,N_23916);
nand U24284 (N_24284,N_23945,N_23708);
xor U24285 (N_24285,N_23917,N_23547);
xor U24286 (N_24286,N_23802,N_23624);
xnor U24287 (N_24287,N_23975,N_23704);
xor U24288 (N_24288,N_23682,N_23629);
or U24289 (N_24289,N_23536,N_23750);
xor U24290 (N_24290,N_23715,N_23994);
nand U24291 (N_24291,N_23565,N_23723);
and U24292 (N_24292,N_23789,N_23660);
or U24293 (N_24293,N_23805,N_23847);
nand U24294 (N_24294,N_23832,N_23954);
nand U24295 (N_24295,N_23864,N_23729);
nand U24296 (N_24296,N_23965,N_23557);
and U24297 (N_24297,N_23694,N_23639);
nor U24298 (N_24298,N_23960,N_23923);
nand U24299 (N_24299,N_23729,N_23983);
nor U24300 (N_24300,N_23726,N_23739);
nor U24301 (N_24301,N_23602,N_23638);
xor U24302 (N_24302,N_23882,N_23847);
nor U24303 (N_24303,N_23536,N_23651);
nor U24304 (N_24304,N_23681,N_23773);
and U24305 (N_24305,N_23975,N_23556);
nor U24306 (N_24306,N_23914,N_23564);
nor U24307 (N_24307,N_23705,N_23545);
xor U24308 (N_24308,N_23988,N_23880);
xnor U24309 (N_24309,N_23641,N_23782);
xor U24310 (N_24310,N_23639,N_23665);
nand U24311 (N_24311,N_23961,N_23951);
or U24312 (N_24312,N_23992,N_23605);
nand U24313 (N_24313,N_23945,N_23721);
nor U24314 (N_24314,N_23833,N_23888);
and U24315 (N_24315,N_23800,N_23565);
nand U24316 (N_24316,N_23596,N_23627);
or U24317 (N_24317,N_23882,N_23925);
and U24318 (N_24318,N_23955,N_23782);
nor U24319 (N_24319,N_23897,N_23734);
xnor U24320 (N_24320,N_23837,N_23500);
nor U24321 (N_24321,N_23685,N_23758);
xnor U24322 (N_24322,N_23908,N_23518);
or U24323 (N_24323,N_23986,N_23733);
nor U24324 (N_24324,N_23878,N_23991);
xnor U24325 (N_24325,N_23900,N_23929);
or U24326 (N_24326,N_23647,N_23892);
nand U24327 (N_24327,N_23943,N_23622);
nor U24328 (N_24328,N_23920,N_23758);
and U24329 (N_24329,N_23931,N_23761);
and U24330 (N_24330,N_23600,N_23875);
xor U24331 (N_24331,N_23680,N_23666);
or U24332 (N_24332,N_23990,N_23924);
nand U24333 (N_24333,N_23644,N_23640);
nor U24334 (N_24334,N_23847,N_23842);
xor U24335 (N_24335,N_23715,N_23898);
nor U24336 (N_24336,N_23575,N_23624);
or U24337 (N_24337,N_23954,N_23583);
and U24338 (N_24338,N_23520,N_23712);
nor U24339 (N_24339,N_23899,N_23564);
nand U24340 (N_24340,N_23611,N_23942);
or U24341 (N_24341,N_23515,N_23684);
xnor U24342 (N_24342,N_23624,N_23989);
or U24343 (N_24343,N_23957,N_23816);
nor U24344 (N_24344,N_23670,N_23761);
or U24345 (N_24345,N_23822,N_23770);
and U24346 (N_24346,N_23765,N_23713);
nor U24347 (N_24347,N_23881,N_23594);
xnor U24348 (N_24348,N_23682,N_23690);
or U24349 (N_24349,N_23871,N_23675);
nand U24350 (N_24350,N_23559,N_23726);
xor U24351 (N_24351,N_23696,N_23911);
nand U24352 (N_24352,N_23623,N_23617);
xor U24353 (N_24353,N_23767,N_23577);
nor U24354 (N_24354,N_23870,N_23695);
nand U24355 (N_24355,N_23908,N_23809);
nor U24356 (N_24356,N_23645,N_23864);
nor U24357 (N_24357,N_23812,N_23942);
nor U24358 (N_24358,N_23702,N_23941);
nor U24359 (N_24359,N_23581,N_23960);
and U24360 (N_24360,N_23816,N_23862);
and U24361 (N_24361,N_23986,N_23967);
nand U24362 (N_24362,N_23877,N_23500);
or U24363 (N_24363,N_23606,N_23659);
xor U24364 (N_24364,N_23773,N_23576);
nand U24365 (N_24365,N_23983,N_23847);
xor U24366 (N_24366,N_23655,N_23669);
or U24367 (N_24367,N_23820,N_23686);
and U24368 (N_24368,N_23838,N_23967);
nand U24369 (N_24369,N_23956,N_23597);
and U24370 (N_24370,N_23951,N_23969);
or U24371 (N_24371,N_23716,N_23898);
xor U24372 (N_24372,N_23568,N_23825);
and U24373 (N_24373,N_23716,N_23884);
xor U24374 (N_24374,N_23936,N_23638);
nand U24375 (N_24375,N_23747,N_23583);
or U24376 (N_24376,N_23883,N_23659);
and U24377 (N_24377,N_23912,N_23609);
nand U24378 (N_24378,N_23696,N_23630);
xor U24379 (N_24379,N_23897,N_23999);
nor U24380 (N_24380,N_23786,N_23593);
or U24381 (N_24381,N_23515,N_23634);
and U24382 (N_24382,N_23886,N_23787);
xor U24383 (N_24383,N_23812,N_23639);
nor U24384 (N_24384,N_23935,N_23563);
nor U24385 (N_24385,N_23973,N_23784);
or U24386 (N_24386,N_23889,N_23685);
or U24387 (N_24387,N_23928,N_23588);
nor U24388 (N_24388,N_23877,N_23713);
nor U24389 (N_24389,N_23767,N_23559);
and U24390 (N_24390,N_23849,N_23765);
nand U24391 (N_24391,N_23776,N_23760);
and U24392 (N_24392,N_23837,N_23797);
nand U24393 (N_24393,N_23965,N_23642);
nor U24394 (N_24394,N_23943,N_23939);
and U24395 (N_24395,N_23539,N_23746);
or U24396 (N_24396,N_23701,N_23666);
nor U24397 (N_24397,N_23701,N_23600);
or U24398 (N_24398,N_23846,N_23739);
and U24399 (N_24399,N_23539,N_23560);
nand U24400 (N_24400,N_23687,N_23726);
or U24401 (N_24401,N_23529,N_23685);
or U24402 (N_24402,N_23821,N_23989);
xor U24403 (N_24403,N_23997,N_23584);
nand U24404 (N_24404,N_23540,N_23937);
and U24405 (N_24405,N_23925,N_23602);
and U24406 (N_24406,N_23969,N_23758);
nand U24407 (N_24407,N_23779,N_23603);
nor U24408 (N_24408,N_23962,N_23921);
and U24409 (N_24409,N_23815,N_23961);
xnor U24410 (N_24410,N_23619,N_23550);
or U24411 (N_24411,N_23733,N_23937);
and U24412 (N_24412,N_23622,N_23643);
xnor U24413 (N_24413,N_23563,N_23868);
or U24414 (N_24414,N_23931,N_23939);
xor U24415 (N_24415,N_23669,N_23639);
xnor U24416 (N_24416,N_23673,N_23570);
nand U24417 (N_24417,N_23891,N_23721);
xnor U24418 (N_24418,N_23626,N_23973);
or U24419 (N_24419,N_23810,N_23979);
xor U24420 (N_24420,N_23535,N_23678);
or U24421 (N_24421,N_23647,N_23925);
nand U24422 (N_24422,N_23567,N_23849);
nor U24423 (N_24423,N_23684,N_23920);
nand U24424 (N_24424,N_23767,N_23663);
nor U24425 (N_24425,N_23619,N_23521);
nand U24426 (N_24426,N_23562,N_23673);
nand U24427 (N_24427,N_23776,N_23657);
and U24428 (N_24428,N_23570,N_23708);
or U24429 (N_24429,N_23676,N_23897);
or U24430 (N_24430,N_23838,N_23873);
nand U24431 (N_24431,N_23883,N_23813);
nand U24432 (N_24432,N_23989,N_23692);
or U24433 (N_24433,N_23584,N_23620);
and U24434 (N_24434,N_23791,N_23805);
and U24435 (N_24435,N_23721,N_23962);
nand U24436 (N_24436,N_23729,N_23844);
xor U24437 (N_24437,N_23726,N_23573);
xnor U24438 (N_24438,N_23744,N_23800);
nand U24439 (N_24439,N_23729,N_23666);
and U24440 (N_24440,N_23855,N_23599);
nand U24441 (N_24441,N_23896,N_23952);
nor U24442 (N_24442,N_23797,N_23996);
and U24443 (N_24443,N_23936,N_23800);
nor U24444 (N_24444,N_23598,N_23717);
nor U24445 (N_24445,N_23596,N_23632);
xnor U24446 (N_24446,N_23760,N_23813);
nor U24447 (N_24447,N_23579,N_23997);
xor U24448 (N_24448,N_23552,N_23842);
nor U24449 (N_24449,N_23767,N_23816);
xnor U24450 (N_24450,N_23737,N_23607);
nor U24451 (N_24451,N_23998,N_23500);
xnor U24452 (N_24452,N_23683,N_23797);
xor U24453 (N_24453,N_23602,N_23822);
or U24454 (N_24454,N_23942,N_23718);
nor U24455 (N_24455,N_23500,N_23961);
nand U24456 (N_24456,N_23679,N_23936);
nand U24457 (N_24457,N_23919,N_23504);
xnor U24458 (N_24458,N_23641,N_23958);
nand U24459 (N_24459,N_23628,N_23535);
nand U24460 (N_24460,N_23898,N_23516);
nor U24461 (N_24461,N_23676,N_23620);
nor U24462 (N_24462,N_23916,N_23812);
xor U24463 (N_24463,N_23558,N_23850);
and U24464 (N_24464,N_23855,N_23843);
nor U24465 (N_24465,N_23835,N_23518);
and U24466 (N_24466,N_23810,N_23945);
and U24467 (N_24467,N_23609,N_23508);
nor U24468 (N_24468,N_23682,N_23532);
or U24469 (N_24469,N_23918,N_23703);
nor U24470 (N_24470,N_23945,N_23702);
nor U24471 (N_24471,N_23546,N_23792);
nand U24472 (N_24472,N_23809,N_23943);
nor U24473 (N_24473,N_23994,N_23686);
xnor U24474 (N_24474,N_23765,N_23933);
xnor U24475 (N_24475,N_23682,N_23971);
and U24476 (N_24476,N_23863,N_23531);
xor U24477 (N_24477,N_23770,N_23682);
nor U24478 (N_24478,N_23696,N_23804);
and U24479 (N_24479,N_23986,N_23935);
xor U24480 (N_24480,N_23543,N_23609);
and U24481 (N_24481,N_23958,N_23662);
nand U24482 (N_24482,N_23764,N_23542);
or U24483 (N_24483,N_23839,N_23933);
xnor U24484 (N_24484,N_23830,N_23610);
nand U24485 (N_24485,N_23590,N_23694);
and U24486 (N_24486,N_23511,N_23710);
or U24487 (N_24487,N_23527,N_23733);
nand U24488 (N_24488,N_23992,N_23937);
nor U24489 (N_24489,N_23939,N_23707);
and U24490 (N_24490,N_23724,N_23903);
and U24491 (N_24491,N_23674,N_23925);
xor U24492 (N_24492,N_23646,N_23617);
or U24493 (N_24493,N_23691,N_23848);
nor U24494 (N_24494,N_23830,N_23732);
and U24495 (N_24495,N_23996,N_23823);
nor U24496 (N_24496,N_23501,N_23520);
nand U24497 (N_24497,N_23690,N_23704);
nand U24498 (N_24498,N_23991,N_23531);
and U24499 (N_24499,N_23756,N_23874);
xor U24500 (N_24500,N_24366,N_24210);
xor U24501 (N_24501,N_24135,N_24243);
nand U24502 (N_24502,N_24102,N_24132);
xor U24503 (N_24503,N_24426,N_24400);
and U24504 (N_24504,N_24436,N_24496);
nand U24505 (N_24505,N_24052,N_24125);
and U24506 (N_24506,N_24450,N_24414);
and U24507 (N_24507,N_24489,N_24474);
or U24508 (N_24508,N_24226,N_24267);
and U24509 (N_24509,N_24310,N_24439);
and U24510 (N_24510,N_24148,N_24271);
nor U24511 (N_24511,N_24260,N_24358);
nand U24512 (N_24512,N_24315,N_24121);
or U24513 (N_24513,N_24368,N_24070);
nor U24514 (N_24514,N_24238,N_24168);
nand U24515 (N_24515,N_24107,N_24209);
and U24516 (N_24516,N_24208,N_24246);
nand U24517 (N_24517,N_24009,N_24118);
nor U24518 (N_24518,N_24266,N_24265);
nand U24519 (N_24519,N_24312,N_24307);
and U24520 (N_24520,N_24375,N_24175);
and U24521 (N_24521,N_24328,N_24424);
nor U24522 (N_24522,N_24099,N_24372);
nand U24523 (N_24523,N_24022,N_24254);
nand U24524 (N_24524,N_24441,N_24104);
or U24525 (N_24525,N_24454,N_24395);
xor U24526 (N_24526,N_24134,N_24300);
nor U24527 (N_24527,N_24288,N_24402);
and U24528 (N_24528,N_24113,N_24393);
nor U24529 (N_24529,N_24153,N_24061);
xor U24530 (N_24530,N_24183,N_24201);
nand U24531 (N_24531,N_24230,N_24001);
xnor U24532 (N_24532,N_24244,N_24075);
and U24533 (N_24533,N_24290,N_24354);
nand U24534 (N_24534,N_24074,N_24455);
xnor U24535 (N_24535,N_24045,N_24004);
nor U24536 (N_24536,N_24369,N_24190);
xor U24537 (N_24537,N_24396,N_24007);
xnor U24538 (N_24538,N_24055,N_24343);
xor U24539 (N_24539,N_24071,N_24464);
or U24540 (N_24540,N_24186,N_24410);
xnor U24541 (N_24541,N_24305,N_24083);
nand U24542 (N_24542,N_24345,N_24385);
xnor U24543 (N_24543,N_24258,N_24398);
nor U24544 (N_24544,N_24108,N_24239);
xor U24545 (N_24545,N_24479,N_24337);
xor U24546 (N_24546,N_24249,N_24157);
or U24547 (N_24547,N_24191,N_24438);
nand U24548 (N_24548,N_24332,N_24042);
nand U24549 (N_24549,N_24361,N_24162);
nor U24550 (N_24550,N_24169,N_24333);
or U24551 (N_24551,N_24459,N_24432);
nand U24552 (N_24552,N_24259,N_24469);
xnor U24553 (N_24553,N_24392,N_24016);
and U24554 (N_24554,N_24470,N_24090);
xor U24555 (N_24555,N_24484,N_24377);
or U24556 (N_24556,N_24199,N_24040);
nand U24557 (N_24557,N_24261,N_24308);
or U24558 (N_24558,N_24468,N_24032);
or U24559 (N_24559,N_24026,N_24081);
xor U24560 (N_24560,N_24110,N_24068);
nor U24561 (N_24561,N_24476,N_24498);
nand U24562 (N_24562,N_24364,N_24471);
and U24563 (N_24563,N_24024,N_24417);
nand U24564 (N_24564,N_24423,N_24281);
nand U24565 (N_24565,N_24050,N_24064);
or U24566 (N_24566,N_24286,N_24115);
xor U24567 (N_24567,N_24403,N_24296);
or U24568 (N_24568,N_24171,N_24399);
nand U24569 (N_24569,N_24039,N_24228);
nor U24570 (N_24570,N_24091,N_24120);
or U24571 (N_24571,N_24105,N_24270);
xnor U24572 (N_24572,N_24057,N_24204);
nor U24573 (N_24573,N_24356,N_24043);
or U24574 (N_24574,N_24287,N_24317);
or U24575 (N_24575,N_24303,N_24086);
nand U24576 (N_24576,N_24234,N_24044);
nand U24577 (N_24577,N_24323,N_24320);
nand U24578 (N_24578,N_24252,N_24179);
or U24579 (N_24579,N_24198,N_24140);
and U24580 (N_24580,N_24486,N_24145);
nor U24581 (N_24581,N_24236,N_24311);
or U24582 (N_24582,N_24406,N_24445);
or U24583 (N_24583,N_24477,N_24394);
nor U24584 (N_24584,N_24442,N_24389);
or U24585 (N_24585,N_24006,N_24018);
or U24586 (N_24586,N_24340,N_24370);
nor U24587 (N_24587,N_24079,N_24376);
or U24588 (N_24588,N_24452,N_24487);
xnor U24589 (N_24589,N_24176,N_24314);
nor U24590 (N_24590,N_24313,N_24278);
nor U24591 (N_24591,N_24355,N_24129);
or U24592 (N_24592,N_24078,N_24206);
nand U24593 (N_24593,N_24002,N_24294);
or U24594 (N_24594,N_24401,N_24297);
nor U24595 (N_24595,N_24242,N_24391);
or U24596 (N_24596,N_24147,N_24447);
nor U24597 (N_24597,N_24155,N_24382);
and U24598 (N_24598,N_24380,N_24212);
xor U24599 (N_24599,N_24381,N_24025);
nand U24600 (N_24600,N_24084,N_24149);
and U24601 (N_24601,N_24128,N_24041);
or U24602 (N_24602,N_24109,N_24008);
nor U24603 (N_24603,N_24282,N_24137);
and U24604 (N_24604,N_24304,N_24427);
nor U24605 (N_24605,N_24180,N_24360);
nand U24606 (N_24606,N_24458,N_24248);
nor U24607 (N_24607,N_24233,N_24220);
nand U24608 (N_24608,N_24425,N_24164);
xnor U24609 (N_24609,N_24273,N_24136);
xor U24610 (N_24610,N_24388,N_24184);
and U24611 (N_24611,N_24031,N_24037);
or U24612 (N_24612,N_24231,N_24250);
nand U24613 (N_24613,N_24344,N_24059);
xor U24614 (N_24614,N_24222,N_24257);
xor U24615 (N_24615,N_24036,N_24277);
nand U24616 (N_24616,N_24205,N_24094);
nor U24617 (N_24617,N_24373,N_24213);
nand U24618 (N_24618,N_24139,N_24269);
xor U24619 (N_24619,N_24080,N_24336);
xnor U24620 (N_24620,N_24338,N_24207);
nor U24621 (N_24621,N_24299,N_24418);
nor U24622 (N_24622,N_24416,N_24272);
and U24623 (N_24623,N_24325,N_24367);
xor U24624 (N_24624,N_24131,N_24027);
nor U24625 (N_24625,N_24289,N_24499);
and U24626 (N_24626,N_24219,N_24327);
or U24627 (N_24627,N_24122,N_24405);
nand U24628 (N_24628,N_24189,N_24283);
or U24629 (N_24629,N_24173,N_24331);
and U24630 (N_24630,N_24152,N_24457);
and U24631 (N_24631,N_24359,N_24443);
or U24632 (N_24632,N_24019,N_24194);
or U24633 (N_24633,N_24185,N_24293);
and U24634 (N_24634,N_24188,N_24444);
nand U24635 (N_24635,N_24143,N_24263);
nor U24636 (N_24636,N_24088,N_24456);
or U24637 (N_24637,N_24352,N_24211);
nor U24638 (N_24638,N_24103,N_24437);
or U24639 (N_24639,N_24229,N_24285);
or U24640 (N_24640,N_24158,N_24430);
and U24641 (N_24641,N_24005,N_24011);
nor U24642 (N_24642,N_24021,N_24256);
or U24643 (N_24643,N_24390,N_24077);
and U24644 (N_24644,N_24087,N_24478);
nor U24645 (N_24645,N_24141,N_24166);
or U24646 (N_24646,N_24003,N_24174);
xnor U24647 (N_24647,N_24497,N_24161);
and U24648 (N_24648,N_24200,N_24112);
or U24649 (N_24649,N_24227,N_24034);
or U24650 (N_24650,N_24301,N_24495);
xnor U24651 (N_24651,N_24097,N_24329);
nor U24652 (N_24652,N_24067,N_24448);
or U24653 (N_24653,N_24472,N_24347);
nor U24654 (N_24654,N_24156,N_24216);
nor U24655 (N_24655,N_24494,N_24069);
or U24656 (N_24656,N_24054,N_24089);
and U24657 (N_24657,N_24339,N_24415);
and U24658 (N_24658,N_24365,N_24202);
and U24659 (N_24659,N_24126,N_24383);
nand U24660 (N_24660,N_24335,N_24453);
or U24661 (N_24661,N_24306,N_24093);
or U24662 (N_24662,N_24363,N_24051);
nand U24663 (N_24663,N_24225,N_24351);
or U24664 (N_24664,N_24013,N_24170);
or U24665 (N_24665,N_24408,N_24435);
or U24666 (N_24666,N_24076,N_24151);
xor U24667 (N_24667,N_24130,N_24350);
or U24668 (N_24668,N_24318,N_24062);
xor U24669 (N_24669,N_24197,N_24488);
xnor U24670 (N_24670,N_24085,N_24462);
or U24671 (N_24671,N_24275,N_24224);
and U24672 (N_24672,N_24292,N_24138);
xnor U24673 (N_24673,N_24480,N_24466);
nor U24674 (N_24674,N_24193,N_24411);
or U24675 (N_24675,N_24124,N_24241);
nand U24676 (N_24676,N_24465,N_24284);
xor U24677 (N_24677,N_24374,N_24413);
nor U24678 (N_24678,N_24251,N_24295);
and U24679 (N_24679,N_24235,N_24181);
and U24680 (N_24680,N_24167,N_24106);
xor U24681 (N_24681,N_24150,N_24023);
nand U24682 (N_24682,N_24268,N_24123);
nor U24683 (N_24683,N_24060,N_24142);
nand U24684 (N_24684,N_24274,N_24279);
or U24685 (N_24685,N_24178,N_24154);
or U24686 (N_24686,N_24264,N_24073);
nor U24687 (N_24687,N_24195,N_24397);
nand U24688 (N_24688,N_24485,N_24255);
or U24689 (N_24689,N_24431,N_24082);
xor U24690 (N_24690,N_24028,N_24460);
or U24691 (N_24691,N_24223,N_24237);
xor U24692 (N_24692,N_24096,N_24117);
nand U24693 (N_24693,N_24187,N_24298);
xor U24694 (N_24694,N_24111,N_24280);
or U24695 (N_24695,N_24326,N_24232);
xnor U24696 (N_24696,N_24262,N_24101);
nand U24697 (N_24697,N_24419,N_24420);
or U24698 (N_24698,N_24066,N_24428);
and U24699 (N_24699,N_24353,N_24046);
nand U24700 (N_24700,N_24362,N_24000);
nor U24701 (N_24701,N_24379,N_24033);
nor U24702 (N_24702,N_24349,N_24483);
and U24703 (N_24703,N_24245,N_24172);
or U24704 (N_24704,N_24330,N_24014);
nand U24705 (N_24705,N_24119,N_24482);
or U24706 (N_24706,N_24160,N_24481);
xor U24707 (N_24707,N_24334,N_24475);
and U24708 (N_24708,N_24063,N_24072);
or U24709 (N_24709,N_24133,N_24467);
xnor U24710 (N_24710,N_24384,N_24029);
xnor U24711 (N_24711,N_24203,N_24053);
and U24712 (N_24712,N_24342,N_24017);
nor U24713 (N_24713,N_24493,N_24449);
nand U24714 (N_24714,N_24341,N_24092);
nand U24715 (N_24715,N_24422,N_24182);
and U24716 (N_24716,N_24433,N_24217);
nand U24717 (N_24717,N_24127,N_24035);
xor U24718 (N_24718,N_24302,N_24463);
xnor U24719 (N_24719,N_24404,N_24065);
nand U24720 (N_24720,N_24215,N_24461);
xnor U24721 (N_24721,N_24163,N_24192);
or U24722 (N_24722,N_24144,N_24049);
and U24723 (N_24723,N_24409,N_24309);
nand U24724 (N_24724,N_24490,N_24316);
nand U24725 (N_24725,N_24319,N_24221);
nand U24726 (N_24726,N_24095,N_24177);
nor U24727 (N_24727,N_24165,N_24159);
xnor U24728 (N_24728,N_24012,N_24214);
xnor U24729 (N_24729,N_24348,N_24386);
nand U24730 (N_24730,N_24446,N_24015);
or U24731 (N_24731,N_24324,N_24357);
xor U24732 (N_24732,N_24412,N_24440);
or U24733 (N_24733,N_24473,N_24491);
nor U24734 (N_24734,N_24346,N_24321);
nor U24735 (N_24735,N_24100,N_24451);
nor U24736 (N_24736,N_24378,N_24291);
and U24737 (N_24737,N_24056,N_24010);
and U24738 (N_24738,N_24020,N_24146);
and U24739 (N_24739,N_24098,N_24048);
and U24740 (N_24740,N_24371,N_24116);
xor U24741 (N_24741,N_24030,N_24429);
and U24742 (N_24742,N_24038,N_24387);
and U24743 (N_24743,N_24434,N_24276);
nand U24744 (N_24744,N_24114,N_24247);
nor U24745 (N_24745,N_24421,N_24322);
or U24746 (N_24746,N_24240,N_24218);
nor U24747 (N_24747,N_24492,N_24047);
and U24748 (N_24748,N_24407,N_24196);
nand U24749 (N_24749,N_24253,N_24058);
and U24750 (N_24750,N_24470,N_24186);
or U24751 (N_24751,N_24438,N_24095);
or U24752 (N_24752,N_24225,N_24045);
nand U24753 (N_24753,N_24282,N_24361);
and U24754 (N_24754,N_24130,N_24116);
nor U24755 (N_24755,N_24228,N_24079);
and U24756 (N_24756,N_24288,N_24474);
nor U24757 (N_24757,N_24296,N_24050);
or U24758 (N_24758,N_24168,N_24180);
or U24759 (N_24759,N_24287,N_24202);
nand U24760 (N_24760,N_24164,N_24145);
and U24761 (N_24761,N_24073,N_24015);
and U24762 (N_24762,N_24286,N_24082);
and U24763 (N_24763,N_24086,N_24296);
and U24764 (N_24764,N_24424,N_24156);
and U24765 (N_24765,N_24283,N_24471);
and U24766 (N_24766,N_24007,N_24275);
or U24767 (N_24767,N_24008,N_24105);
or U24768 (N_24768,N_24393,N_24345);
and U24769 (N_24769,N_24327,N_24024);
xor U24770 (N_24770,N_24034,N_24306);
nand U24771 (N_24771,N_24273,N_24270);
nand U24772 (N_24772,N_24279,N_24373);
xnor U24773 (N_24773,N_24461,N_24126);
nand U24774 (N_24774,N_24488,N_24108);
nand U24775 (N_24775,N_24218,N_24319);
xor U24776 (N_24776,N_24009,N_24086);
or U24777 (N_24777,N_24255,N_24367);
or U24778 (N_24778,N_24027,N_24426);
nand U24779 (N_24779,N_24021,N_24471);
nor U24780 (N_24780,N_24006,N_24126);
and U24781 (N_24781,N_24342,N_24232);
or U24782 (N_24782,N_24166,N_24117);
and U24783 (N_24783,N_24024,N_24357);
nand U24784 (N_24784,N_24188,N_24006);
or U24785 (N_24785,N_24365,N_24207);
or U24786 (N_24786,N_24072,N_24161);
nor U24787 (N_24787,N_24164,N_24473);
xnor U24788 (N_24788,N_24399,N_24247);
xnor U24789 (N_24789,N_24398,N_24130);
or U24790 (N_24790,N_24093,N_24444);
nor U24791 (N_24791,N_24467,N_24200);
xor U24792 (N_24792,N_24411,N_24172);
and U24793 (N_24793,N_24396,N_24314);
xor U24794 (N_24794,N_24346,N_24159);
nor U24795 (N_24795,N_24446,N_24429);
and U24796 (N_24796,N_24175,N_24386);
xor U24797 (N_24797,N_24249,N_24301);
nand U24798 (N_24798,N_24353,N_24148);
or U24799 (N_24799,N_24185,N_24158);
nor U24800 (N_24800,N_24074,N_24111);
nand U24801 (N_24801,N_24195,N_24386);
and U24802 (N_24802,N_24150,N_24055);
nand U24803 (N_24803,N_24209,N_24188);
and U24804 (N_24804,N_24099,N_24373);
and U24805 (N_24805,N_24095,N_24339);
nand U24806 (N_24806,N_24453,N_24009);
nor U24807 (N_24807,N_24188,N_24149);
and U24808 (N_24808,N_24265,N_24175);
nand U24809 (N_24809,N_24338,N_24276);
nand U24810 (N_24810,N_24213,N_24226);
nand U24811 (N_24811,N_24146,N_24353);
xor U24812 (N_24812,N_24251,N_24358);
xor U24813 (N_24813,N_24055,N_24076);
nand U24814 (N_24814,N_24000,N_24170);
xnor U24815 (N_24815,N_24321,N_24317);
or U24816 (N_24816,N_24005,N_24285);
nor U24817 (N_24817,N_24228,N_24277);
or U24818 (N_24818,N_24010,N_24041);
nor U24819 (N_24819,N_24352,N_24480);
nand U24820 (N_24820,N_24449,N_24434);
xnor U24821 (N_24821,N_24116,N_24294);
and U24822 (N_24822,N_24348,N_24288);
xnor U24823 (N_24823,N_24290,N_24178);
and U24824 (N_24824,N_24269,N_24423);
nand U24825 (N_24825,N_24344,N_24171);
or U24826 (N_24826,N_24012,N_24089);
and U24827 (N_24827,N_24168,N_24005);
or U24828 (N_24828,N_24336,N_24240);
nor U24829 (N_24829,N_24367,N_24298);
or U24830 (N_24830,N_24477,N_24412);
and U24831 (N_24831,N_24497,N_24065);
or U24832 (N_24832,N_24233,N_24459);
nand U24833 (N_24833,N_24152,N_24211);
and U24834 (N_24834,N_24446,N_24426);
nand U24835 (N_24835,N_24142,N_24337);
nor U24836 (N_24836,N_24169,N_24353);
xor U24837 (N_24837,N_24028,N_24330);
xnor U24838 (N_24838,N_24338,N_24489);
nand U24839 (N_24839,N_24353,N_24189);
or U24840 (N_24840,N_24032,N_24470);
and U24841 (N_24841,N_24343,N_24114);
or U24842 (N_24842,N_24369,N_24069);
nor U24843 (N_24843,N_24415,N_24067);
and U24844 (N_24844,N_24334,N_24258);
nand U24845 (N_24845,N_24259,N_24445);
and U24846 (N_24846,N_24142,N_24057);
and U24847 (N_24847,N_24244,N_24495);
nor U24848 (N_24848,N_24474,N_24249);
nor U24849 (N_24849,N_24101,N_24298);
or U24850 (N_24850,N_24231,N_24271);
nor U24851 (N_24851,N_24212,N_24364);
or U24852 (N_24852,N_24053,N_24027);
nand U24853 (N_24853,N_24259,N_24406);
or U24854 (N_24854,N_24397,N_24436);
or U24855 (N_24855,N_24222,N_24480);
xor U24856 (N_24856,N_24185,N_24318);
xnor U24857 (N_24857,N_24148,N_24053);
nand U24858 (N_24858,N_24254,N_24019);
xor U24859 (N_24859,N_24002,N_24199);
nor U24860 (N_24860,N_24058,N_24227);
and U24861 (N_24861,N_24290,N_24469);
and U24862 (N_24862,N_24395,N_24166);
nand U24863 (N_24863,N_24499,N_24072);
nor U24864 (N_24864,N_24129,N_24000);
nor U24865 (N_24865,N_24327,N_24496);
xnor U24866 (N_24866,N_24169,N_24250);
nand U24867 (N_24867,N_24344,N_24354);
xnor U24868 (N_24868,N_24052,N_24020);
or U24869 (N_24869,N_24475,N_24461);
and U24870 (N_24870,N_24233,N_24054);
nand U24871 (N_24871,N_24379,N_24278);
and U24872 (N_24872,N_24164,N_24357);
nand U24873 (N_24873,N_24313,N_24245);
nand U24874 (N_24874,N_24081,N_24400);
or U24875 (N_24875,N_24000,N_24162);
or U24876 (N_24876,N_24216,N_24478);
nand U24877 (N_24877,N_24123,N_24265);
or U24878 (N_24878,N_24449,N_24077);
xnor U24879 (N_24879,N_24426,N_24305);
and U24880 (N_24880,N_24265,N_24386);
nand U24881 (N_24881,N_24187,N_24495);
and U24882 (N_24882,N_24082,N_24217);
and U24883 (N_24883,N_24046,N_24172);
and U24884 (N_24884,N_24493,N_24166);
or U24885 (N_24885,N_24058,N_24497);
or U24886 (N_24886,N_24118,N_24495);
or U24887 (N_24887,N_24462,N_24070);
or U24888 (N_24888,N_24192,N_24259);
and U24889 (N_24889,N_24303,N_24457);
xnor U24890 (N_24890,N_24206,N_24291);
xor U24891 (N_24891,N_24268,N_24055);
or U24892 (N_24892,N_24402,N_24416);
nor U24893 (N_24893,N_24499,N_24194);
nor U24894 (N_24894,N_24278,N_24358);
nand U24895 (N_24895,N_24087,N_24264);
nor U24896 (N_24896,N_24209,N_24252);
nand U24897 (N_24897,N_24066,N_24025);
xnor U24898 (N_24898,N_24458,N_24356);
nor U24899 (N_24899,N_24230,N_24428);
xnor U24900 (N_24900,N_24324,N_24289);
nand U24901 (N_24901,N_24072,N_24012);
and U24902 (N_24902,N_24283,N_24413);
xor U24903 (N_24903,N_24155,N_24079);
or U24904 (N_24904,N_24358,N_24456);
and U24905 (N_24905,N_24139,N_24129);
and U24906 (N_24906,N_24132,N_24014);
xnor U24907 (N_24907,N_24466,N_24489);
and U24908 (N_24908,N_24272,N_24257);
and U24909 (N_24909,N_24480,N_24357);
and U24910 (N_24910,N_24286,N_24297);
nand U24911 (N_24911,N_24187,N_24218);
and U24912 (N_24912,N_24199,N_24284);
nand U24913 (N_24913,N_24108,N_24216);
xor U24914 (N_24914,N_24309,N_24174);
xor U24915 (N_24915,N_24087,N_24053);
nor U24916 (N_24916,N_24481,N_24112);
nand U24917 (N_24917,N_24156,N_24361);
nor U24918 (N_24918,N_24187,N_24031);
xor U24919 (N_24919,N_24001,N_24247);
xnor U24920 (N_24920,N_24115,N_24435);
or U24921 (N_24921,N_24483,N_24161);
nor U24922 (N_24922,N_24186,N_24029);
xnor U24923 (N_24923,N_24289,N_24109);
nor U24924 (N_24924,N_24352,N_24066);
xnor U24925 (N_24925,N_24074,N_24424);
nor U24926 (N_24926,N_24098,N_24119);
nand U24927 (N_24927,N_24338,N_24359);
nor U24928 (N_24928,N_24454,N_24099);
nor U24929 (N_24929,N_24036,N_24271);
xor U24930 (N_24930,N_24071,N_24467);
xor U24931 (N_24931,N_24300,N_24167);
nand U24932 (N_24932,N_24315,N_24282);
and U24933 (N_24933,N_24147,N_24123);
and U24934 (N_24934,N_24382,N_24117);
nand U24935 (N_24935,N_24132,N_24443);
and U24936 (N_24936,N_24060,N_24417);
nor U24937 (N_24937,N_24071,N_24325);
nand U24938 (N_24938,N_24238,N_24227);
xnor U24939 (N_24939,N_24085,N_24308);
and U24940 (N_24940,N_24357,N_24316);
xor U24941 (N_24941,N_24073,N_24295);
nor U24942 (N_24942,N_24325,N_24108);
and U24943 (N_24943,N_24129,N_24496);
and U24944 (N_24944,N_24457,N_24426);
or U24945 (N_24945,N_24238,N_24117);
nand U24946 (N_24946,N_24157,N_24026);
and U24947 (N_24947,N_24216,N_24314);
and U24948 (N_24948,N_24352,N_24196);
xnor U24949 (N_24949,N_24433,N_24099);
and U24950 (N_24950,N_24266,N_24268);
nor U24951 (N_24951,N_24121,N_24340);
or U24952 (N_24952,N_24126,N_24313);
nor U24953 (N_24953,N_24170,N_24038);
or U24954 (N_24954,N_24337,N_24480);
and U24955 (N_24955,N_24349,N_24079);
and U24956 (N_24956,N_24422,N_24073);
and U24957 (N_24957,N_24107,N_24009);
xor U24958 (N_24958,N_24185,N_24219);
or U24959 (N_24959,N_24344,N_24302);
nand U24960 (N_24960,N_24014,N_24418);
and U24961 (N_24961,N_24259,N_24011);
and U24962 (N_24962,N_24446,N_24471);
xor U24963 (N_24963,N_24285,N_24034);
nor U24964 (N_24964,N_24272,N_24291);
xnor U24965 (N_24965,N_24294,N_24242);
or U24966 (N_24966,N_24103,N_24465);
or U24967 (N_24967,N_24226,N_24234);
nor U24968 (N_24968,N_24014,N_24271);
nor U24969 (N_24969,N_24155,N_24356);
and U24970 (N_24970,N_24015,N_24376);
nor U24971 (N_24971,N_24477,N_24009);
or U24972 (N_24972,N_24191,N_24365);
xor U24973 (N_24973,N_24011,N_24324);
and U24974 (N_24974,N_24010,N_24318);
or U24975 (N_24975,N_24392,N_24107);
xor U24976 (N_24976,N_24034,N_24038);
nor U24977 (N_24977,N_24293,N_24267);
nand U24978 (N_24978,N_24197,N_24086);
or U24979 (N_24979,N_24448,N_24321);
xor U24980 (N_24980,N_24069,N_24176);
xnor U24981 (N_24981,N_24111,N_24393);
nand U24982 (N_24982,N_24288,N_24295);
xnor U24983 (N_24983,N_24365,N_24326);
nand U24984 (N_24984,N_24392,N_24196);
or U24985 (N_24985,N_24359,N_24168);
nand U24986 (N_24986,N_24118,N_24117);
and U24987 (N_24987,N_24241,N_24261);
nand U24988 (N_24988,N_24202,N_24175);
nand U24989 (N_24989,N_24220,N_24490);
nor U24990 (N_24990,N_24302,N_24113);
nor U24991 (N_24991,N_24073,N_24315);
nor U24992 (N_24992,N_24115,N_24402);
xor U24993 (N_24993,N_24499,N_24053);
nor U24994 (N_24994,N_24299,N_24013);
nor U24995 (N_24995,N_24401,N_24337);
nor U24996 (N_24996,N_24225,N_24322);
or U24997 (N_24997,N_24371,N_24008);
xnor U24998 (N_24998,N_24368,N_24416);
nor U24999 (N_24999,N_24368,N_24499);
or UO_0 (O_0,N_24500,N_24891);
xnor UO_1 (O_1,N_24897,N_24748);
nand UO_2 (O_2,N_24653,N_24989);
nor UO_3 (O_3,N_24684,N_24872);
and UO_4 (O_4,N_24736,N_24835);
xnor UO_5 (O_5,N_24717,N_24976);
or UO_6 (O_6,N_24559,N_24606);
nand UO_7 (O_7,N_24534,N_24594);
nor UO_8 (O_8,N_24861,N_24763);
or UO_9 (O_9,N_24902,N_24612);
nor UO_10 (O_10,N_24522,N_24659);
nor UO_11 (O_11,N_24850,N_24884);
nand UO_12 (O_12,N_24503,N_24889);
and UO_13 (O_13,N_24587,N_24845);
nand UO_14 (O_14,N_24535,N_24859);
nor UO_15 (O_15,N_24724,N_24993);
and UO_16 (O_16,N_24521,N_24570);
nand UO_17 (O_17,N_24805,N_24870);
or UO_18 (O_18,N_24580,N_24563);
and UO_19 (O_19,N_24704,N_24793);
or UO_20 (O_20,N_24557,N_24985);
xor UO_21 (O_21,N_24782,N_24525);
and UO_22 (O_22,N_24928,N_24914);
xnor UO_23 (O_23,N_24945,N_24990);
xor UO_24 (O_24,N_24556,N_24555);
nand UO_25 (O_25,N_24591,N_24548);
and UO_26 (O_26,N_24940,N_24955);
or UO_27 (O_27,N_24740,N_24616);
and UO_28 (O_28,N_24537,N_24597);
nand UO_29 (O_29,N_24953,N_24677);
and UO_30 (O_30,N_24607,N_24841);
nor UO_31 (O_31,N_24987,N_24689);
and UO_32 (O_32,N_24982,N_24577);
or UO_33 (O_33,N_24942,N_24600);
nor UO_34 (O_34,N_24718,N_24610);
and UO_35 (O_35,N_24957,N_24807);
nor UO_36 (O_36,N_24762,N_24691);
xnor UO_37 (O_37,N_24708,N_24731);
or UO_38 (O_38,N_24735,N_24648);
nand UO_39 (O_39,N_24703,N_24721);
or UO_40 (O_40,N_24560,N_24753);
nor UO_41 (O_41,N_24797,N_24780);
nand UO_42 (O_42,N_24714,N_24880);
or UO_43 (O_43,N_24871,N_24681);
nand UO_44 (O_44,N_24685,N_24988);
nor UO_45 (O_45,N_24937,N_24775);
or UO_46 (O_46,N_24778,N_24671);
nand UO_47 (O_47,N_24707,N_24628);
or UO_48 (O_48,N_24770,N_24886);
or UO_49 (O_49,N_24911,N_24565);
xor UO_50 (O_50,N_24929,N_24826);
nor UO_51 (O_51,N_24571,N_24562);
or UO_52 (O_52,N_24879,N_24792);
or UO_53 (O_53,N_24665,N_24692);
nand UO_54 (O_54,N_24833,N_24634);
nor UO_55 (O_55,N_24526,N_24668);
xnor UO_56 (O_56,N_24589,N_24925);
nand UO_57 (O_57,N_24547,N_24745);
nand UO_58 (O_58,N_24983,N_24979);
or UO_59 (O_59,N_24935,N_24933);
and UO_60 (O_60,N_24842,N_24764);
or UO_61 (O_61,N_24725,N_24854);
and UO_62 (O_62,N_24849,N_24794);
nand UO_63 (O_63,N_24661,N_24908);
and UO_64 (O_64,N_24912,N_24552);
or UO_65 (O_65,N_24791,N_24630);
nand UO_66 (O_66,N_24624,N_24734);
or UO_67 (O_67,N_24887,N_24952);
xnor UO_68 (O_68,N_24881,N_24575);
nand UO_69 (O_69,N_24650,N_24528);
xnor UO_70 (O_70,N_24705,N_24706);
or UO_71 (O_71,N_24649,N_24924);
and UO_72 (O_72,N_24781,N_24803);
xor UO_73 (O_73,N_24864,N_24601);
or UO_74 (O_74,N_24852,N_24651);
and UO_75 (O_75,N_24964,N_24515);
and UO_76 (O_76,N_24750,N_24939);
nand UO_77 (O_77,N_24627,N_24837);
nand UO_78 (O_78,N_24590,N_24638);
and UO_79 (O_79,N_24749,N_24669);
nor UO_80 (O_80,N_24509,N_24644);
and UO_81 (O_81,N_24569,N_24761);
and UO_82 (O_82,N_24822,N_24629);
xor UO_83 (O_83,N_24810,N_24848);
nand UO_84 (O_84,N_24965,N_24532);
nor UO_85 (O_85,N_24863,N_24844);
and UO_86 (O_86,N_24647,N_24585);
or UO_87 (O_87,N_24977,N_24802);
nor UO_88 (O_88,N_24742,N_24943);
and UO_89 (O_89,N_24814,N_24968);
nand UO_90 (O_90,N_24727,N_24954);
or UO_91 (O_91,N_24998,N_24790);
nand UO_92 (O_92,N_24632,N_24655);
nand UO_93 (O_93,N_24815,N_24769);
and UO_94 (O_94,N_24710,N_24550);
or UO_95 (O_95,N_24866,N_24816);
xnor UO_96 (O_96,N_24817,N_24739);
or UO_97 (O_97,N_24930,N_24843);
nand UO_98 (O_98,N_24916,N_24660);
nand UO_99 (O_99,N_24573,N_24679);
nor UO_100 (O_100,N_24905,N_24621);
and UO_101 (O_101,N_24549,N_24969);
nand UO_102 (O_102,N_24583,N_24698);
or UO_103 (O_103,N_24611,N_24546);
or UO_104 (O_104,N_24729,N_24959);
nand UO_105 (O_105,N_24862,N_24533);
and UO_106 (O_106,N_24609,N_24572);
xor UO_107 (O_107,N_24754,N_24923);
xor UO_108 (O_108,N_24658,N_24869);
nor UO_109 (O_109,N_24633,N_24512);
nand UO_110 (O_110,N_24819,N_24752);
or UO_111 (O_111,N_24619,N_24696);
xor UO_112 (O_112,N_24962,N_24919);
or UO_113 (O_113,N_24697,N_24637);
or UO_114 (O_114,N_24834,N_24922);
or UO_115 (O_115,N_24542,N_24950);
or UO_116 (O_116,N_24894,N_24558);
xnor UO_117 (O_117,N_24598,N_24530);
or UO_118 (O_118,N_24787,N_24757);
nor UO_119 (O_119,N_24733,N_24510);
nand UO_120 (O_120,N_24693,N_24830);
xnor UO_121 (O_121,N_24578,N_24504);
or UO_122 (O_122,N_24529,N_24910);
xor UO_123 (O_123,N_24980,N_24520);
xnor UO_124 (O_124,N_24788,N_24926);
nor UO_125 (O_125,N_24858,N_24978);
nand UO_126 (O_126,N_24992,N_24620);
nor UO_127 (O_127,N_24878,N_24865);
and UO_128 (O_128,N_24947,N_24813);
nand UO_129 (O_129,N_24799,N_24516);
or UO_130 (O_130,N_24544,N_24915);
nor UO_131 (O_131,N_24768,N_24643);
nand UO_132 (O_132,N_24818,N_24895);
or UO_133 (O_133,N_24801,N_24545);
nand UO_134 (O_134,N_24554,N_24673);
nor UO_135 (O_135,N_24743,N_24507);
or UO_136 (O_136,N_24672,N_24779);
xnor UO_137 (O_137,N_24682,N_24700);
nand UO_138 (O_138,N_24994,N_24795);
and UO_139 (O_139,N_24666,N_24613);
xnor UO_140 (O_140,N_24513,N_24851);
or UO_141 (O_141,N_24719,N_24900);
nand UO_142 (O_142,N_24896,N_24519);
nor UO_143 (O_143,N_24680,N_24756);
or UO_144 (O_144,N_24592,N_24899);
nor UO_145 (O_145,N_24586,N_24951);
or UO_146 (O_146,N_24765,N_24553);
or UO_147 (O_147,N_24995,N_24972);
nand UO_148 (O_148,N_24588,N_24543);
nand UO_149 (O_149,N_24662,N_24938);
nor UO_150 (O_150,N_24712,N_24695);
nand UO_151 (O_151,N_24747,N_24956);
or UO_152 (O_152,N_24986,N_24664);
nand UO_153 (O_153,N_24892,N_24738);
and UO_154 (O_154,N_24683,N_24511);
or UO_155 (O_155,N_24709,N_24767);
nor UO_156 (O_156,N_24966,N_24971);
and UO_157 (O_157,N_24776,N_24716);
or UO_158 (O_158,N_24564,N_24847);
nand UO_159 (O_159,N_24991,N_24856);
nand UO_160 (O_160,N_24614,N_24970);
and UO_161 (O_161,N_24702,N_24777);
xor UO_162 (O_162,N_24903,N_24825);
nand UO_163 (O_163,N_24618,N_24875);
xor UO_164 (O_164,N_24783,N_24800);
nand UO_165 (O_165,N_24631,N_24867);
and UO_166 (O_166,N_24687,N_24711);
or UO_167 (O_167,N_24723,N_24868);
and UO_168 (O_168,N_24674,N_24773);
or UO_169 (O_169,N_24882,N_24518);
nand UO_170 (O_170,N_24904,N_24806);
xnor UO_171 (O_171,N_24574,N_24934);
nor UO_172 (O_172,N_24646,N_24579);
nor UO_173 (O_173,N_24502,N_24804);
or UO_174 (O_174,N_24909,N_24656);
xnor UO_175 (O_175,N_24626,N_24999);
and UO_176 (O_176,N_24784,N_24888);
and UO_177 (O_177,N_24615,N_24785);
and UO_178 (O_178,N_24876,N_24744);
or UO_179 (O_179,N_24846,N_24786);
nor UO_180 (O_180,N_24766,N_24602);
xnor UO_181 (O_181,N_24809,N_24523);
nand UO_182 (O_182,N_24996,N_24675);
nand UO_183 (O_183,N_24531,N_24874);
and UO_184 (O_184,N_24949,N_24760);
xnor UO_185 (O_185,N_24857,N_24652);
nand UO_186 (O_186,N_24853,N_24737);
and UO_187 (O_187,N_24694,N_24877);
xor UO_188 (O_188,N_24936,N_24517);
xnor UO_189 (O_189,N_24829,N_24941);
or UO_190 (O_190,N_24824,N_24827);
nor UO_191 (O_191,N_24595,N_24932);
or UO_192 (O_192,N_24641,N_24603);
nor UO_193 (O_193,N_24541,N_24771);
or UO_194 (O_194,N_24622,N_24883);
nor UO_195 (O_195,N_24582,N_24623);
nor UO_196 (O_196,N_24981,N_24811);
nor UO_197 (O_197,N_24715,N_24840);
and UO_198 (O_198,N_24755,N_24561);
or UO_199 (O_199,N_24625,N_24774);
or UO_200 (O_200,N_24640,N_24593);
or UO_201 (O_201,N_24838,N_24820);
xor UO_202 (O_202,N_24596,N_24828);
nor UO_203 (O_203,N_24568,N_24720);
and UO_204 (O_204,N_24948,N_24686);
and UO_205 (O_205,N_24636,N_24821);
xor UO_206 (O_206,N_24690,N_24581);
nor UO_207 (O_207,N_24961,N_24997);
or UO_208 (O_208,N_24732,N_24812);
nand UO_209 (O_209,N_24927,N_24920);
nor UO_210 (O_210,N_24508,N_24974);
nand UO_211 (O_211,N_24642,N_24772);
nand UO_212 (O_212,N_24505,N_24676);
nor UO_213 (O_213,N_24890,N_24832);
or UO_214 (O_214,N_24701,N_24605);
xor UO_215 (O_215,N_24960,N_24808);
or UO_216 (O_216,N_24654,N_24670);
and UO_217 (O_217,N_24635,N_24963);
or UO_218 (O_218,N_24751,N_24688);
and UO_219 (O_219,N_24663,N_24873);
or UO_220 (O_220,N_24514,N_24893);
and UO_221 (O_221,N_24726,N_24678);
nand UO_222 (O_222,N_24713,N_24823);
nor UO_223 (O_223,N_24599,N_24758);
and UO_224 (O_224,N_24639,N_24608);
or UO_225 (O_225,N_24860,N_24931);
xnor UO_226 (O_226,N_24913,N_24501);
or UO_227 (O_227,N_24921,N_24898);
or UO_228 (O_228,N_24567,N_24789);
xor UO_229 (O_229,N_24831,N_24839);
or UO_230 (O_230,N_24527,N_24551);
or UO_231 (O_231,N_24566,N_24728);
or UO_232 (O_232,N_24657,N_24901);
xor UO_233 (O_233,N_24539,N_24958);
xor UO_234 (O_234,N_24918,N_24906);
nand UO_235 (O_235,N_24730,N_24538);
or UO_236 (O_236,N_24741,N_24984);
and UO_237 (O_237,N_24946,N_24645);
or UO_238 (O_238,N_24885,N_24944);
and UO_239 (O_239,N_24699,N_24576);
or UO_240 (O_240,N_24796,N_24975);
nand UO_241 (O_241,N_24973,N_24855);
nor UO_242 (O_242,N_24836,N_24524);
nor UO_243 (O_243,N_24536,N_24746);
or UO_244 (O_244,N_24967,N_24759);
nand UO_245 (O_245,N_24722,N_24667);
nand UO_246 (O_246,N_24506,N_24917);
or UO_247 (O_247,N_24617,N_24584);
xnor UO_248 (O_248,N_24604,N_24907);
nand UO_249 (O_249,N_24798,N_24540);
xor UO_250 (O_250,N_24866,N_24658);
or UO_251 (O_251,N_24803,N_24962);
xnor UO_252 (O_252,N_24866,N_24590);
nand UO_253 (O_253,N_24564,N_24846);
or UO_254 (O_254,N_24818,N_24936);
or UO_255 (O_255,N_24829,N_24567);
nand UO_256 (O_256,N_24519,N_24675);
or UO_257 (O_257,N_24508,N_24692);
and UO_258 (O_258,N_24551,N_24972);
or UO_259 (O_259,N_24899,N_24965);
and UO_260 (O_260,N_24655,N_24841);
nor UO_261 (O_261,N_24682,N_24703);
or UO_262 (O_262,N_24669,N_24958);
or UO_263 (O_263,N_24810,N_24720);
nand UO_264 (O_264,N_24893,N_24678);
nor UO_265 (O_265,N_24923,N_24893);
xnor UO_266 (O_266,N_24742,N_24846);
xor UO_267 (O_267,N_24934,N_24943);
nor UO_268 (O_268,N_24527,N_24803);
or UO_269 (O_269,N_24627,N_24985);
or UO_270 (O_270,N_24923,N_24591);
or UO_271 (O_271,N_24912,N_24521);
xor UO_272 (O_272,N_24525,N_24529);
or UO_273 (O_273,N_24978,N_24907);
or UO_274 (O_274,N_24817,N_24694);
or UO_275 (O_275,N_24942,N_24534);
and UO_276 (O_276,N_24549,N_24605);
xnor UO_277 (O_277,N_24677,N_24560);
xnor UO_278 (O_278,N_24537,N_24624);
nand UO_279 (O_279,N_24838,N_24580);
nor UO_280 (O_280,N_24981,N_24610);
xnor UO_281 (O_281,N_24732,N_24855);
and UO_282 (O_282,N_24621,N_24526);
nor UO_283 (O_283,N_24739,N_24529);
or UO_284 (O_284,N_24655,N_24978);
or UO_285 (O_285,N_24599,N_24866);
nand UO_286 (O_286,N_24946,N_24682);
nand UO_287 (O_287,N_24971,N_24917);
xnor UO_288 (O_288,N_24806,N_24649);
nand UO_289 (O_289,N_24711,N_24583);
xnor UO_290 (O_290,N_24932,N_24616);
nand UO_291 (O_291,N_24927,N_24864);
nor UO_292 (O_292,N_24719,N_24850);
or UO_293 (O_293,N_24898,N_24542);
nand UO_294 (O_294,N_24953,N_24617);
or UO_295 (O_295,N_24736,N_24926);
or UO_296 (O_296,N_24878,N_24614);
xor UO_297 (O_297,N_24799,N_24724);
or UO_298 (O_298,N_24644,N_24820);
or UO_299 (O_299,N_24898,N_24647);
and UO_300 (O_300,N_24921,N_24578);
or UO_301 (O_301,N_24513,N_24671);
or UO_302 (O_302,N_24970,N_24794);
and UO_303 (O_303,N_24688,N_24612);
xor UO_304 (O_304,N_24903,N_24645);
and UO_305 (O_305,N_24759,N_24952);
nand UO_306 (O_306,N_24577,N_24688);
nand UO_307 (O_307,N_24790,N_24604);
nor UO_308 (O_308,N_24677,N_24936);
xor UO_309 (O_309,N_24813,N_24591);
and UO_310 (O_310,N_24632,N_24894);
xor UO_311 (O_311,N_24505,N_24509);
nand UO_312 (O_312,N_24696,N_24944);
xor UO_313 (O_313,N_24963,N_24628);
nor UO_314 (O_314,N_24792,N_24767);
or UO_315 (O_315,N_24972,N_24630);
or UO_316 (O_316,N_24861,N_24723);
or UO_317 (O_317,N_24733,N_24505);
xor UO_318 (O_318,N_24584,N_24625);
and UO_319 (O_319,N_24936,N_24667);
nor UO_320 (O_320,N_24935,N_24510);
nor UO_321 (O_321,N_24917,N_24908);
nor UO_322 (O_322,N_24973,N_24874);
xnor UO_323 (O_323,N_24852,N_24918);
or UO_324 (O_324,N_24633,N_24782);
or UO_325 (O_325,N_24614,N_24518);
xor UO_326 (O_326,N_24842,N_24828);
xor UO_327 (O_327,N_24771,N_24593);
nor UO_328 (O_328,N_24819,N_24985);
xor UO_329 (O_329,N_24834,N_24876);
or UO_330 (O_330,N_24821,N_24544);
or UO_331 (O_331,N_24890,N_24796);
or UO_332 (O_332,N_24870,N_24751);
nand UO_333 (O_333,N_24509,N_24824);
and UO_334 (O_334,N_24627,N_24925);
nor UO_335 (O_335,N_24951,N_24853);
nand UO_336 (O_336,N_24765,N_24811);
nand UO_337 (O_337,N_24590,N_24707);
xor UO_338 (O_338,N_24837,N_24952);
and UO_339 (O_339,N_24674,N_24856);
nor UO_340 (O_340,N_24877,N_24925);
xor UO_341 (O_341,N_24895,N_24619);
nor UO_342 (O_342,N_24637,N_24828);
or UO_343 (O_343,N_24990,N_24859);
xnor UO_344 (O_344,N_24870,N_24844);
and UO_345 (O_345,N_24558,N_24706);
nand UO_346 (O_346,N_24761,N_24758);
nand UO_347 (O_347,N_24573,N_24893);
or UO_348 (O_348,N_24999,N_24609);
nand UO_349 (O_349,N_24566,N_24812);
nor UO_350 (O_350,N_24507,N_24582);
or UO_351 (O_351,N_24809,N_24801);
nand UO_352 (O_352,N_24614,N_24643);
xor UO_353 (O_353,N_24949,N_24506);
xor UO_354 (O_354,N_24924,N_24945);
xnor UO_355 (O_355,N_24665,N_24923);
nand UO_356 (O_356,N_24916,N_24854);
nor UO_357 (O_357,N_24951,N_24771);
and UO_358 (O_358,N_24704,N_24611);
nand UO_359 (O_359,N_24685,N_24712);
nor UO_360 (O_360,N_24555,N_24892);
and UO_361 (O_361,N_24530,N_24811);
or UO_362 (O_362,N_24922,N_24739);
and UO_363 (O_363,N_24553,N_24651);
nor UO_364 (O_364,N_24532,N_24606);
or UO_365 (O_365,N_24775,N_24993);
and UO_366 (O_366,N_24751,N_24848);
nand UO_367 (O_367,N_24535,N_24968);
nor UO_368 (O_368,N_24797,N_24777);
nor UO_369 (O_369,N_24927,N_24627);
and UO_370 (O_370,N_24677,N_24757);
or UO_371 (O_371,N_24522,N_24705);
nor UO_372 (O_372,N_24797,N_24727);
or UO_373 (O_373,N_24802,N_24706);
or UO_374 (O_374,N_24978,N_24722);
nand UO_375 (O_375,N_24729,N_24631);
nor UO_376 (O_376,N_24744,N_24544);
or UO_377 (O_377,N_24738,N_24817);
nor UO_378 (O_378,N_24723,N_24804);
nor UO_379 (O_379,N_24780,N_24596);
xnor UO_380 (O_380,N_24818,N_24637);
and UO_381 (O_381,N_24851,N_24990);
nor UO_382 (O_382,N_24907,N_24658);
xor UO_383 (O_383,N_24723,N_24765);
and UO_384 (O_384,N_24915,N_24769);
and UO_385 (O_385,N_24507,N_24737);
nor UO_386 (O_386,N_24622,N_24581);
and UO_387 (O_387,N_24728,N_24597);
and UO_388 (O_388,N_24656,N_24672);
nand UO_389 (O_389,N_24654,N_24788);
or UO_390 (O_390,N_24686,N_24939);
and UO_391 (O_391,N_24632,N_24889);
nor UO_392 (O_392,N_24671,N_24816);
nor UO_393 (O_393,N_24581,N_24579);
xor UO_394 (O_394,N_24681,N_24638);
nor UO_395 (O_395,N_24866,N_24871);
nor UO_396 (O_396,N_24808,N_24826);
nand UO_397 (O_397,N_24572,N_24714);
and UO_398 (O_398,N_24662,N_24715);
xnor UO_399 (O_399,N_24692,N_24774);
or UO_400 (O_400,N_24556,N_24581);
and UO_401 (O_401,N_24769,N_24622);
nor UO_402 (O_402,N_24741,N_24703);
and UO_403 (O_403,N_24526,N_24944);
xnor UO_404 (O_404,N_24884,N_24950);
or UO_405 (O_405,N_24999,N_24940);
and UO_406 (O_406,N_24943,N_24996);
nor UO_407 (O_407,N_24599,N_24563);
nand UO_408 (O_408,N_24545,N_24921);
or UO_409 (O_409,N_24982,N_24882);
nand UO_410 (O_410,N_24975,N_24690);
nand UO_411 (O_411,N_24765,N_24654);
or UO_412 (O_412,N_24617,N_24520);
nor UO_413 (O_413,N_24912,N_24939);
and UO_414 (O_414,N_24544,N_24623);
and UO_415 (O_415,N_24613,N_24614);
and UO_416 (O_416,N_24716,N_24789);
nor UO_417 (O_417,N_24841,N_24832);
xor UO_418 (O_418,N_24665,N_24689);
nand UO_419 (O_419,N_24954,N_24761);
nand UO_420 (O_420,N_24517,N_24860);
xnor UO_421 (O_421,N_24623,N_24919);
nor UO_422 (O_422,N_24575,N_24548);
nor UO_423 (O_423,N_24504,N_24510);
nor UO_424 (O_424,N_24537,N_24580);
and UO_425 (O_425,N_24658,N_24785);
and UO_426 (O_426,N_24819,N_24899);
and UO_427 (O_427,N_24740,N_24948);
nand UO_428 (O_428,N_24782,N_24582);
nor UO_429 (O_429,N_24806,N_24877);
nand UO_430 (O_430,N_24893,N_24666);
nor UO_431 (O_431,N_24686,N_24542);
and UO_432 (O_432,N_24536,N_24552);
and UO_433 (O_433,N_24508,N_24991);
xnor UO_434 (O_434,N_24954,N_24628);
xor UO_435 (O_435,N_24690,N_24880);
nor UO_436 (O_436,N_24821,N_24908);
nand UO_437 (O_437,N_24702,N_24811);
nor UO_438 (O_438,N_24590,N_24549);
nor UO_439 (O_439,N_24600,N_24643);
nor UO_440 (O_440,N_24628,N_24744);
nand UO_441 (O_441,N_24914,N_24835);
or UO_442 (O_442,N_24717,N_24548);
and UO_443 (O_443,N_24920,N_24605);
xnor UO_444 (O_444,N_24999,N_24731);
nor UO_445 (O_445,N_24887,N_24684);
nand UO_446 (O_446,N_24970,N_24883);
xnor UO_447 (O_447,N_24979,N_24809);
nor UO_448 (O_448,N_24537,N_24981);
xor UO_449 (O_449,N_24516,N_24853);
or UO_450 (O_450,N_24779,N_24629);
and UO_451 (O_451,N_24950,N_24833);
and UO_452 (O_452,N_24678,N_24849);
xnor UO_453 (O_453,N_24781,N_24895);
or UO_454 (O_454,N_24796,N_24816);
and UO_455 (O_455,N_24941,N_24652);
or UO_456 (O_456,N_24545,N_24530);
and UO_457 (O_457,N_24556,N_24585);
xor UO_458 (O_458,N_24791,N_24537);
or UO_459 (O_459,N_24782,N_24538);
xor UO_460 (O_460,N_24747,N_24772);
xnor UO_461 (O_461,N_24828,N_24638);
xnor UO_462 (O_462,N_24716,N_24528);
nand UO_463 (O_463,N_24940,N_24897);
or UO_464 (O_464,N_24686,N_24924);
or UO_465 (O_465,N_24527,N_24814);
nand UO_466 (O_466,N_24800,N_24805);
or UO_467 (O_467,N_24653,N_24830);
nor UO_468 (O_468,N_24524,N_24730);
nor UO_469 (O_469,N_24757,N_24513);
nand UO_470 (O_470,N_24653,N_24640);
or UO_471 (O_471,N_24533,N_24739);
nor UO_472 (O_472,N_24666,N_24791);
or UO_473 (O_473,N_24932,N_24594);
or UO_474 (O_474,N_24768,N_24682);
or UO_475 (O_475,N_24940,N_24828);
nor UO_476 (O_476,N_24519,N_24650);
xor UO_477 (O_477,N_24961,N_24881);
xnor UO_478 (O_478,N_24557,N_24643);
nand UO_479 (O_479,N_24802,N_24973);
and UO_480 (O_480,N_24783,N_24830);
nor UO_481 (O_481,N_24640,N_24610);
or UO_482 (O_482,N_24764,N_24925);
and UO_483 (O_483,N_24974,N_24640);
and UO_484 (O_484,N_24612,N_24954);
nor UO_485 (O_485,N_24561,N_24724);
nand UO_486 (O_486,N_24853,N_24747);
nor UO_487 (O_487,N_24686,N_24625);
and UO_488 (O_488,N_24574,N_24529);
xnor UO_489 (O_489,N_24589,N_24705);
or UO_490 (O_490,N_24655,N_24901);
nand UO_491 (O_491,N_24657,N_24886);
and UO_492 (O_492,N_24758,N_24968);
and UO_493 (O_493,N_24512,N_24994);
and UO_494 (O_494,N_24833,N_24545);
nand UO_495 (O_495,N_24700,N_24537);
nor UO_496 (O_496,N_24911,N_24949);
nor UO_497 (O_497,N_24912,N_24537);
xnor UO_498 (O_498,N_24940,N_24996);
nor UO_499 (O_499,N_24569,N_24813);
nor UO_500 (O_500,N_24656,N_24641);
nor UO_501 (O_501,N_24816,N_24874);
xnor UO_502 (O_502,N_24501,N_24997);
nand UO_503 (O_503,N_24614,N_24727);
nand UO_504 (O_504,N_24906,N_24551);
or UO_505 (O_505,N_24930,N_24519);
or UO_506 (O_506,N_24584,N_24895);
or UO_507 (O_507,N_24937,N_24770);
or UO_508 (O_508,N_24736,N_24878);
nor UO_509 (O_509,N_24848,N_24842);
or UO_510 (O_510,N_24872,N_24653);
xnor UO_511 (O_511,N_24581,N_24578);
and UO_512 (O_512,N_24592,N_24728);
or UO_513 (O_513,N_24805,N_24944);
or UO_514 (O_514,N_24535,N_24654);
xnor UO_515 (O_515,N_24605,N_24607);
nand UO_516 (O_516,N_24741,N_24889);
or UO_517 (O_517,N_24884,N_24956);
xnor UO_518 (O_518,N_24582,N_24629);
nor UO_519 (O_519,N_24525,N_24524);
and UO_520 (O_520,N_24577,N_24976);
and UO_521 (O_521,N_24815,N_24705);
xnor UO_522 (O_522,N_24832,N_24746);
and UO_523 (O_523,N_24700,N_24590);
xnor UO_524 (O_524,N_24872,N_24590);
nor UO_525 (O_525,N_24980,N_24699);
nand UO_526 (O_526,N_24680,N_24550);
or UO_527 (O_527,N_24513,N_24742);
nor UO_528 (O_528,N_24809,N_24791);
xnor UO_529 (O_529,N_24804,N_24564);
or UO_530 (O_530,N_24677,N_24963);
and UO_531 (O_531,N_24593,N_24878);
nor UO_532 (O_532,N_24947,N_24570);
and UO_533 (O_533,N_24582,N_24675);
xor UO_534 (O_534,N_24712,N_24999);
nand UO_535 (O_535,N_24578,N_24549);
or UO_536 (O_536,N_24534,N_24569);
nor UO_537 (O_537,N_24587,N_24801);
xor UO_538 (O_538,N_24727,N_24965);
nand UO_539 (O_539,N_24808,N_24845);
nor UO_540 (O_540,N_24924,N_24660);
nand UO_541 (O_541,N_24771,N_24740);
nor UO_542 (O_542,N_24901,N_24915);
xnor UO_543 (O_543,N_24931,N_24921);
nor UO_544 (O_544,N_24542,N_24629);
or UO_545 (O_545,N_24786,N_24878);
or UO_546 (O_546,N_24741,N_24632);
or UO_547 (O_547,N_24860,N_24774);
xnor UO_548 (O_548,N_24757,N_24616);
xnor UO_549 (O_549,N_24844,N_24693);
nand UO_550 (O_550,N_24867,N_24686);
and UO_551 (O_551,N_24663,N_24932);
and UO_552 (O_552,N_24701,N_24540);
nand UO_553 (O_553,N_24945,N_24514);
nor UO_554 (O_554,N_24657,N_24816);
nand UO_555 (O_555,N_24893,N_24715);
nand UO_556 (O_556,N_24943,N_24900);
xnor UO_557 (O_557,N_24660,N_24663);
nor UO_558 (O_558,N_24934,N_24571);
xnor UO_559 (O_559,N_24627,N_24770);
xnor UO_560 (O_560,N_24593,N_24875);
or UO_561 (O_561,N_24605,N_24674);
nor UO_562 (O_562,N_24874,N_24755);
nor UO_563 (O_563,N_24501,N_24712);
and UO_564 (O_564,N_24695,N_24551);
or UO_565 (O_565,N_24814,N_24735);
or UO_566 (O_566,N_24580,N_24540);
xnor UO_567 (O_567,N_24728,N_24695);
or UO_568 (O_568,N_24943,N_24510);
nand UO_569 (O_569,N_24977,N_24675);
xnor UO_570 (O_570,N_24966,N_24627);
xor UO_571 (O_571,N_24635,N_24849);
or UO_572 (O_572,N_24725,N_24840);
nand UO_573 (O_573,N_24836,N_24924);
xnor UO_574 (O_574,N_24559,N_24967);
or UO_575 (O_575,N_24527,N_24843);
xnor UO_576 (O_576,N_24830,N_24944);
nand UO_577 (O_577,N_24879,N_24531);
nand UO_578 (O_578,N_24791,N_24886);
xnor UO_579 (O_579,N_24613,N_24541);
nor UO_580 (O_580,N_24821,N_24846);
nor UO_581 (O_581,N_24616,N_24918);
nor UO_582 (O_582,N_24793,N_24551);
and UO_583 (O_583,N_24900,N_24753);
nand UO_584 (O_584,N_24989,N_24678);
and UO_585 (O_585,N_24588,N_24990);
nor UO_586 (O_586,N_24849,N_24961);
or UO_587 (O_587,N_24918,N_24706);
nor UO_588 (O_588,N_24796,N_24954);
xor UO_589 (O_589,N_24830,N_24768);
xnor UO_590 (O_590,N_24623,N_24878);
nor UO_591 (O_591,N_24796,N_24689);
nand UO_592 (O_592,N_24754,N_24572);
and UO_593 (O_593,N_24710,N_24554);
and UO_594 (O_594,N_24779,N_24815);
or UO_595 (O_595,N_24778,N_24787);
xnor UO_596 (O_596,N_24631,N_24721);
or UO_597 (O_597,N_24975,N_24587);
and UO_598 (O_598,N_24963,N_24701);
and UO_599 (O_599,N_24860,N_24547);
or UO_600 (O_600,N_24687,N_24732);
xnor UO_601 (O_601,N_24945,N_24731);
xor UO_602 (O_602,N_24950,N_24783);
xnor UO_603 (O_603,N_24929,N_24919);
nor UO_604 (O_604,N_24637,N_24503);
or UO_605 (O_605,N_24908,N_24533);
or UO_606 (O_606,N_24617,N_24773);
or UO_607 (O_607,N_24901,N_24721);
xor UO_608 (O_608,N_24818,N_24557);
xor UO_609 (O_609,N_24523,N_24667);
nor UO_610 (O_610,N_24517,N_24745);
nor UO_611 (O_611,N_24791,N_24701);
nor UO_612 (O_612,N_24605,N_24856);
nand UO_613 (O_613,N_24871,N_24913);
and UO_614 (O_614,N_24913,N_24852);
nor UO_615 (O_615,N_24934,N_24731);
or UO_616 (O_616,N_24794,N_24843);
and UO_617 (O_617,N_24701,N_24883);
or UO_618 (O_618,N_24547,N_24564);
and UO_619 (O_619,N_24507,N_24531);
nand UO_620 (O_620,N_24520,N_24957);
xor UO_621 (O_621,N_24726,N_24567);
or UO_622 (O_622,N_24551,N_24860);
or UO_623 (O_623,N_24691,N_24839);
nand UO_624 (O_624,N_24748,N_24760);
xnor UO_625 (O_625,N_24877,N_24858);
and UO_626 (O_626,N_24605,N_24968);
xnor UO_627 (O_627,N_24824,N_24676);
nor UO_628 (O_628,N_24787,N_24912);
xnor UO_629 (O_629,N_24715,N_24996);
nand UO_630 (O_630,N_24913,N_24862);
nor UO_631 (O_631,N_24777,N_24703);
or UO_632 (O_632,N_24616,N_24761);
and UO_633 (O_633,N_24567,N_24634);
nor UO_634 (O_634,N_24671,N_24918);
or UO_635 (O_635,N_24744,N_24840);
nand UO_636 (O_636,N_24628,N_24677);
nand UO_637 (O_637,N_24599,N_24627);
and UO_638 (O_638,N_24938,N_24685);
or UO_639 (O_639,N_24624,N_24916);
and UO_640 (O_640,N_24648,N_24984);
or UO_641 (O_641,N_24773,N_24574);
and UO_642 (O_642,N_24719,N_24696);
and UO_643 (O_643,N_24707,N_24901);
or UO_644 (O_644,N_24912,N_24868);
nand UO_645 (O_645,N_24518,N_24724);
nor UO_646 (O_646,N_24818,N_24837);
xnor UO_647 (O_647,N_24663,N_24502);
and UO_648 (O_648,N_24592,N_24626);
nand UO_649 (O_649,N_24686,N_24769);
nand UO_650 (O_650,N_24549,N_24709);
and UO_651 (O_651,N_24775,N_24923);
and UO_652 (O_652,N_24992,N_24874);
or UO_653 (O_653,N_24552,N_24628);
nand UO_654 (O_654,N_24683,N_24909);
nor UO_655 (O_655,N_24952,N_24602);
nor UO_656 (O_656,N_24890,N_24658);
xnor UO_657 (O_657,N_24966,N_24606);
xnor UO_658 (O_658,N_24504,N_24883);
xnor UO_659 (O_659,N_24781,N_24590);
nor UO_660 (O_660,N_24943,N_24532);
or UO_661 (O_661,N_24680,N_24903);
xor UO_662 (O_662,N_24838,N_24643);
and UO_663 (O_663,N_24583,N_24520);
or UO_664 (O_664,N_24796,N_24839);
or UO_665 (O_665,N_24886,N_24767);
nand UO_666 (O_666,N_24894,N_24975);
and UO_667 (O_667,N_24501,N_24548);
or UO_668 (O_668,N_24865,N_24949);
xnor UO_669 (O_669,N_24776,N_24874);
xor UO_670 (O_670,N_24531,N_24828);
nor UO_671 (O_671,N_24508,N_24680);
and UO_672 (O_672,N_24558,N_24919);
nor UO_673 (O_673,N_24602,N_24979);
or UO_674 (O_674,N_24516,N_24636);
or UO_675 (O_675,N_24907,N_24785);
nor UO_676 (O_676,N_24562,N_24993);
nor UO_677 (O_677,N_24924,N_24701);
or UO_678 (O_678,N_24535,N_24521);
and UO_679 (O_679,N_24708,N_24752);
nand UO_680 (O_680,N_24567,N_24880);
nor UO_681 (O_681,N_24568,N_24560);
nor UO_682 (O_682,N_24672,N_24897);
or UO_683 (O_683,N_24713,N_24557);
or UO_684 (O_684,N_24840,N_24852);
or UO_685 (O_685,N_24629,N_24739);
nand UO_686 (O_686,N_24816,N_24879);
nand UO_687 (O_687,N_24555,N_24646);
and UO_688 (O_688,N_24842,N_24906);
xor UO_689 (O_689,N_24849,N_24823);
and UO_690 (O_690,N_24826,N_24857);
or UO_691 (O_691,N_24518,N_24954);
nand UO_692 (O_692,N_24558,N_24855);
nor UO_693 (O_693,N_24976,N_24506);
nand UO_694 (O_694,N_24804,N_24921);
and UO_695 (O_695,N_24843,N_24659);
nor UO_696 (O_696,N_24887,N_24821);
nand UO_697 (O_697,N_24561,N_24729);
and UO_698 (O_698,N_24750,N_24902);
or UO_699 (O_699,N_24750,N_24566);
or UO_700 (O_700,N_24775,N_24795);
or UO_701 (O_701,N_24770,N_24715);
nor UO_702 (O_702,N_24912,N_24794);
xor UO_703 (O_703,N_24779,N_24541);
nor UO_704 (O_704,N_24525,N_24993);
nand UO_705 (O_705,N_24637,N_24812);
and UO_706 (O_706,N_24862,N_24772);
nand UO_707 (O_707,N_24647,N_24891);
or UO_708 (O_708,N_24715,N_24667);
or UO_709 (O_709,N_24783,N_24728);
nand UO_710 (O_710,N_24684,N_24919);
and UO_711 (O_711,N_24856,N_24990);
xor UO_712 (O_712,N_24830,N_24799);
or UO_713 (O_713,N_24855,N_24778);
nand UO_714 (O_714,N_24819,N_24787);
xor UO_715 (O_715,N_24998,N_24629);
nand UO_716 (O_716,N_24733,N_24867);
or UO_717 (O_717,N_24923,N_24840);
or UO_718 (O_718,N_24917,N_24888);
nand UO_719 (O_719,N_24558,N_24772);
xor UO_720 (O_720,N_24597,N_24824);
and UO_721 (O_721,N_24810,N_24521);
and UO_722 (O_722,N_24518,N_24690);
and UO_723 (O_723,N_24747,N_24977);
xnor UO_724 (O_724,N_24660,N_24532);
nand UO_725 (O_725,N_24538,N_24860);
xor UO_726 (O_726,N_24926,N_24843);
or UO_727 (O_727,N_24515,N_24942);
and UO_728 (O_728,N_24794,N_24745);
xor UO_729 (O_729,N_24665,N_24716);
xor UO_730 (O_730,N_24852,N_24527);
and UO_731 (O_731,N_24768,N_24529);
nor UO_732 (O_732,N_24984,N_24885);
or UO_733 (O_733,N_24874,N_24782);
xor UO_734 (O_734,N_24959,N_24972);
or UO_735 (O_735,N_24666,N_24672);
nand UO_736 (O_736,N_24557,N_24906);
xor UO_737 (O_737,N_24905,N_24661);
or UO_738 (O_738,N_24703,N_24951);
or UO_739 (O_739,N_24518,N_24616);
nand UO_740 (O_740,N_24704,N_24878);
or UO_741 (O_741,N_24618,N_24924);
or UO_742 (O_742,N_24701,N_24703);
nand UO_743 (O_743,N_24971,N_24653);
xnor UO_744 (O_744,N_24849,N_24586);
nor UO_745 (O_745,N_24531,N_24897);
or UO_746 (O_746,N_24555,N_24580);
or UO_747 (O_747,N_24845,N_24694);
xnor UO_748 (O_748,N_24824,N_24756);
xnor UO_749 (O_749,N_24970,N_24688);
nand UO_750 (O_750,N_24614,N_24829);
nor UO_751 (O_751,N_24662,N_24547);
nand UO_752 (O_752,N_24933,N_24666);
nor UO_753 (O_753,N_24774,N_24540);
or UO_754 (O_754,N_24920,N_24601);
xor UO_755 (O_755,N_24691,N_24510);
and UO_756 (O_756,N_24902,N_24787);
or UO_757 (O_757,N_24936,N_24993);
and UO_758 (O_758,N_24686,N_24610);
nor UO_759 (O_759,N_24757,N_24530);
or UO_760 (O_760,N_24877,N_24539);
and UO_761 (O_761,N_24574,N_24812);
nand UO_762 (O_762,N_24713,N_24638);
nand UO_763 (O_763,N_24620,N_24886);
or UO_764 (O_764,N_24629,N_24948);
or UO_765 (O_765,N_24897,N_24920);
nand UO_766 (O_766,N_24848,N_24799);
nor UO_767 (O_767,N_24723,N_24604);
or UO_768 (O_768,N_24580,N_24571);
or UO_769 (O_769,N_24962,N_24826);
nor UO_770 (O_770,N_24523,N_24966);
xor UO_771 (O_771,N_24976,N_24903);
nand UO_772 (O_772,N_24819,N_24884);
nor UO_773 (O_773,N_24970,N_24894);
and UO_774 (O_774,N_24506,N_24601);
xor UO_775 (O_775,N_24654,N_24716);
nor UO_776 (O_776,N_24626,N_24979);
and UO_777 (O_777,N_24649,N_24521);
or UO_778 (O_778,N_24734,N_24840);
nand UO_779 (O_779,N_24951,N_24881);
nor UO_780 (O_780,N_24652,N_24584);
or UO_781 (O_781,N_24779,N_24952);
nand UO_782 (O_782,N_24756,N_24936);
and UO_783 (O_783,N_24796,N_24789);
or UO_784 (O_784,N_24842,N_24954);
or UO_785 (O_785,N_24588,N_24822);
and UO_786 (O_786,N_24820,N_24797);
and UO_787 (O_787,N_24737,N_24843);
or UO_788 (O_788,N_24731,N_24831);
and UO_789 (O_789,N_24822,N_24556);
and UO_790 (O_790,N_24891,N_24666);
xnor UO_791 (O_791,N_24976,N_24993);
xnor UO_792 (O_792,N_24982,N_24719);
xor UO_793 (O_793,N_24639,N_24609);
nand UO_794 (O_794,N_24911,N_24753);
xnor UO_795 (O_795,N_24900,N_24628);
nor UO_796 (O_796,N_24977,N_24637);
and UO_797 (O_797,N_24687,N_24931);
nor UO_798 (O_798,N_24641,N_24565);
nor UO_799 (O_799,N_24722,N_24734);
nor UO_800 (O_800,N_24709,N_24894);
and UO_801 (O_801,N_24512,N_24906);
xnor UO_802 (O_802,N_24852,N_24648);
or UO_803 (O_803,N_24595,N_24541);
or UO_804 (O_804,N_24705,N_24675);
and UO_805 (O_805,N_24793,N_24941);
nand UO_806 (O_806,N_24736,N_24921);
or UO_807 (O_807,N_24532,N_24788);
or UO_808 (O_808,N_24817,N_24578);
or UO_809 (O_809,N_24618,N_24557);
nand UO_810 (O_810,N_24656,N_24785);
xnor UO_811 (O_811,N_24945,N_24590);
xnor UO_812 (O_812,N_24988,N_24720);
xor UO_813 (O_813,N_24971,N_24619);
and UO_814 (O_814,N_24997,N_24612);
or UO_815 (O_815,N_24911,N_24873);
nand UO_816 (O_816,N_24705,N_24613);
xor UO_817 (O_817,N_24592,N_24554);
nor UO_818 (O_818,N_24949,N_24666);
nor UO_819 (O_819,N_24939,N_24704);
xnor UO_820 (O_820,N_24802,N_24623);
or UO_821 (O_821,N_24982,N_24930);
and UO_822 (O_822,N_24510,N_24976);
nor UO_823 (O_823,N_24590,N_24975);
or UO_824 (O_824,N_24614,N_24562);
xor UO_825 (O_825,N_24714,N_24847);
xnor UO_826 (O_826,N_24925,N_24669);
xnor UO_827 (O_827,N_24997,N_24668);
nor UO_828 (O_828,N_24879,N_24568);
xnor UO_829 (O_829,N_24803,N_24575);
and UO_830 (O_830,N_24517,N_24850);
and UO_831 (O_831,N_24729,N_24765);
nor UO_832 (O_832,N_24561,N_24959);
xor UO_833 (O_833,N_24805,N_24530);
nor UO_834 (O_834,N_24563,N_24808);
nor UO_835 (O_835,N_24527,N_24747);
or UO_836 (O_836,N_24529,N_24785);
nand UO_837 (O_837,N_24596,N_24578);
nand UO_838 (O_838,N_24983,N_24507);
and UO_839 (O_839,N_24820,N_24790);
nor UO_840 (O_840,N_24746,N_24684);
and UO_841 (O_841,N_24579,N_24613);
nor UO_842 (O_842,N_24751,N_24916);
or UO_843 (O_843,N_24525,N_24705);
or UO_844 (O_844,N_24718,N_24661);
nor UO_845 (O_845,N_24890,N_24990);
or UO_846 (O_846,N_24924,N_24596);
or UO_847 (O_847,N_24976,N_24753);
nand UO_848 (O_848,N_24723,N_24615);
or UO_849 (O_849,N_24634,N_24901);
nor UO_850 (O_850,N_24750,N_24697);
xnor UO_851 (O_851,N_24939,N_24572);
or UO_852 (O_852,N_24566,N_24780);
nor UO_853 (O_853,N_24579,N_24836);
or UO_854 (O_854,N_24762,N_24626);
xor UO_855 (O_855,N_24878,N_24726);
and UO_856 (O_856,N_24952,N_24623);
xor UO_857 (O_857,N_24918,N_24591);
xor UO_858 (O_858,N_24758,N_24515);
nor UO_859 (O_859,N_24667,N_24519);
and UO_860 (O_860,N_24810,N_24547);
nand UO_861 (O_861,N_24703,N_24879);
and UO_862 (O_862,N_24803,N_24511);
nand UO_863 (O_863,N_24941,N_24516);
and UO_864 (O_864,N_24769,N_24588);
or UO_865 (O_865,N_24571,N_24594);
nand UO_866 (O_866,N_24801,N_24682);
or UO_867 (O_867,N_24956,N_24999);
or UO_868 (O_868,N_24855,N_24683);
xnor UO_869 (O_869,N_24591,N_24891);
or UO_870 (O_870,N_24804,N_24760);
and UO_871 (O_871,N_24937,N_24716);
and UO_872 (O_872,N_24865,N_24699);
and UO_873 (O_873,N_24634,N_24795);
and UO_874 (O_874,N_24822,N_24745);
xor UO_875 (O_875,N_24933,N_24642);
and UO_876 (O_876,N_24838,N_24616);
nor UO_877 (O_877,N_24607,N_24623);
or UO_878 (O_878,N_24636,N_24875);
and UO_879 (O_879,N_24606,N_24727);
nor UO_880 (O_880,N_24851,N_24528);
nand UO_881 (O_881,N_24640,N_24558);
and UO_882 (O_882,N_24750,N_24995);
or UO_883 (O_883,N_24651,N_24989);
and UO_884 (O_884,N_24781,N_24904);
xnor UO_885 (O_885,N_24535,N_24798);
and UO_886 (O_886,N_24629,N_24992);
nand UO_887 (O_887,N_24566,N_24943);
or UO_888 (O_888,N_24608,N_24758);
xor UO_889 (O_889,N_24759,N_24521);
xnor UO_890 (O_890,N_24559,N_24610);
xnor UO_891 (O_891,N_24974,N_24889);
and UO_892 (O_892,N_24544,N_24548);
and UO_893 (O_893,N_24850,N_24663);
nand UO_894 (O_894,N_24836,N_24652);
or UO_895 (O_895,N_24863,N_24749);
nor UO_896 (O_896,N_24769,N_24537);
or UO_897 (O_897,N_24534,N_24768);
xor UO_898 (O_898,N_24881,N_24941);
xnor UO_899 (O_899,N_24942,N_24913);
or UO_900 (O_900,N_24750,N_24853);
nor UO_901 (O_901,N_24743,N_24878);
xnor UO_902 (O_902,N_24908,N_24612);
and UO_903 (O_903,N_24663,N_24654);
nor UO_904 (O_904,N_24967,N_24971);
and UO_905 (O_905,N_24554,N_24997);
and UO_906 (O_906,N_24853,N_24677);
nand UO_907 (O_907,N_24728,N_24588);
xor UO_908 (O_908,N_24746,N_24764);
nor UO_909 (O_909,N_24892,N_24878);
or UO_910 (O_910,N_24863,N_24791);
nand UO_911 (O_911,N_24797,N_24549);
nor UO_912 (O_912,N_24608,N_24511);
or UO_913 (O_913,N_24968,N_24659);
or UO_914 (O_914,N_24861,N_24521);
or UO_915 (O_915,N_24611,N_24950);
or UO_916 (O_916,N_24580,N_24916);
nand UO_917 (O_917,N_24507,N_24740);
xor UO_918 (O_918,N_24692,N_24945);
nor UO_919 (O_919,N_24654,N_24933);
xor UO_920 (O_920,N_24908,N_24554);
nand UO_921 (O_921,N_24825,N_24842);
xnor UO_922 (O_922,N_24852,N_24734);
xnor UO_923 (O_923,N_24610,N_24990);
xor UO_924 (O_924,N_24790,N_24635);
nor UO_925 (O_925,N_24880,N_24520);
and UO_926 (O_926,N_24699,N_24588);
nor UO_927 (O_927,N_24757,N_24653);
and UO_928 (O_928,N_24892,N_24685);
and UO_929 (O_929,N_24776,N_24579);
and UO_930 (O_930,N_24647,N_24867);
nand UO_931 (O_931,N_24661,N_24712);
nor UO_932 (O_932,N_24585,N_24904);
and UO_933 (O_933,N_24600,N_24944);
nor UO_934 (O_934,N_24860,N_24812);
nand UO_935 (O_935,N_24994,N_24986);
and UO_936 (O_936,N_24852,N_24778);
nand UO_937 (O_937,N_24856,N_24680);
and UO_938 (O_938,N_24525,N_24727);
or UO_939 (O_939,N_24961,N_24876);
xor UO_940 (O_940,N_24949,N_24566);
or UO_941 (O_941,N_24778,N_24747);
nor UO_942 (O_942,N_24855,N_24582);
or UO_943 (O_943,N_24833,N_24731);
xnor UO_944 (O_944,N_24841,N_24537);
and UO_945 (O_945,N_24961,N_24917);
and UO_946 (O_946,N_24583,N_24661);
nor UO_947 (O_947,N_24957,N_24904);
and UO_948 (O_948,N_24520,N_24685);
and UO_949 (O_949,N_24975,N_24578);
or UO_950 (O_950,N_24734,N_24588);
nor UO_951 (O_951,N_24995,N_24659);
nor UO_952 (O_952,N_24620,N_24560);
nand UO_953 (O_953,N_24779,N_24992);
xor UO_954 (O_954,N_24826,N_24837);
and UO_955 (O_955,N_24611,N_24598);
and UO_956 (O_956,N_24759,N_24566);
and UO_957 (O_957,N_24734,N_24837);
and UO_958 (O_958,N_24538,N_24948);
nand UO_959 (O_959,N_24657,N_24740);
and UO_960 (O_960,N_24918,N_24746);
nor UO_961 (O_961,N_24719,N_24714);
and UO_962 (O_962,N_24564,N_24700);
nand UO_963 (O_963,N_24770,N_24841);
nor UO_964 (O_964,N_24909,N_24511);
xnor UO_965 (O_965,N_24802,N_24998);
or UO_966 (O_966,N_24856,N_24553);
nor UO_967 (O_967,N_24767,N_24870);
nand UO_968 (O_968,N_24777,N_24871);
xnor UO_969 (O_969,N_24967,N_24877);
or UO_970 (O_970,N_24871,N_24773);
xnor UO_971 (O_971,N_24659,N_24607);
or UO_972 (O_972,N_24802,N_24543);
xor UO_973 (O_973,N_24521,N_24824);
xnor UO_974 (O_974,N_24506,N_24938);
nand UO_975 (O_975,N_24724,N_24615);
xor UO_976 (O_976,N_24552,N_24688);
nand UO_977 (O_977,N_24847,N_24757);
and UO_978 (O_978,N_24552,N_24569);
xor UO_979 (O_979,N_24951,N_24682);
nand UO_980 (O_980,N_24654,N_24982);
xor UO_981 (O_981,N_24955,N_24759);
xor UO_982 (O_982,N_24951,N_24800);
and UO_983 (O_983,N_24863,N_24864);
or UO_984 (O_984,N_24850,N_24891);
and UO_985 (O_985,N_24994,N_24697);
nand UO_986 (O_986,N_24693,N_24984);
and UO_987 (O_987,N_24868,N_24926);
nor UO_988 (O_988,N_24677,N_24509);
nand UO_989 (O_989,N_24588,N_24913);
or UO_990 (O_990,N_24724,N_24956);
nand UO_991 (O_991,N_24984,N_24858);
and UO_992 (O_992,N_24660,N_24806);
xnor UO_993 (O_993,N_24559,N_24848);
nand UO_994 (O_994,N_24948,N_24632);
xor UO_995 (O_995,N_24988,N_24582);
or UO_996 (O_996,N_24532,N_24685);
nor UO_997 (O_997,N_24727,N_24623);
or UO_998 (O_998,N_24985,N_24778);
xnor UO_999 (O_999,N_24948,N_24993);
or UO_1000 (O_1000,N_24700,N_24912);
or UO_1001 (O_1001,N_24948,N_24685);
and UO_1002 (O_1002,N_24778,N_24615);
and UO_1003 (O_1003,N_24856,N_24844);
or UO_1004 (O_1004,N_24833,N_24508);
or UO_1005 (O_1005,N_24533,N_24826);
nand UO_1006 (O_1006,N_24804,N_24687);
and UO_1007 (O_1007,N_24536,N_24639);
and UO_1008 (O_1008,N_24935,N_24998);
or UO_1009 (O_1009,N_24641,N_24894);
nor UO_1010 (O_1010,N_24669,N_24629);
xor UO_1011 (O_1011,N_24998,N_24890);
and UO_1012 (O_1012,N_24937,N_24872);
and UO_1013 (O_1013,N_24902,N_24969);
xnor UO_1014 (O_1014,N_24812,N_24547);
or UO_1015 (O_1015,N_24619,N_24524);
and UO_1016 (O_1016,N_24752,N_24780);
nand UO_1017 (O_1017,N_24632,N_24757);
or UO_1018 (O_1018,N_24673,N_24937);
and UO_1019 (O_1019,N_24920,N_24848);
nor UO_1020 (O_1020,N_24897,N_24728);
nand UO_1021 (O_1021,N_24836,N_24814);
and UO_1022 (O_1022,N_24886,N_24903);
xor UO_1023 (O_1023,N_24965,N_24527);
nor UO_1024 (O_1024,N_24728,N_24762);
nand UO_1025 (O_1025,N_24861,N_24587);
nand UO_1026 (O_1026,N_24961,N_24552);
or UO_1027 (O_1027,N_24856,N_24803);
nor UO_1028 (O_1028,N_24671,N_24626);
xor UO_1029 (O_1029,N_24855,N_24964);
and UO_1030 (O_1030,N_24831,N_24799);
nor UO_1031 (O_1031,N_24588,N_24645);
or UO_1032 (O_1032,N_24618,N_24825);
nand UO_1033 (O_1033,N_24748,N_24782);
xnor UO_1034 (O_1034,N_24829,N_24676);
xnor UO_1035 (O_1035,N_24693,N_24542);
nand UO_1036 (O_1036,N_24563,N_24957);
nand UO_1037 (O_1037,N_24661,N_24628);
xnor UO_1038 (O_1038,N_24905,N_24696);
nand UO_1039 (O_1039,N_24813,N_24858);
nor UO_1040 (O_1040,N_24533,N_24603);
or UO_1041 (O_1041,N_24647,N_24611);
nor UO_1042 (O_1042,N_24923,N_24683);
or UO_1043 (O_1043,N_24911,N_24850);
xnor UO_1044 (O_1044,N_24637,N_24885);
and UO_1045 (O_1045,N_24643,N_24967);
and UO_1046 (O_1046,N_24533,N_24592);
or UO_1047 (O_1047,N_24990,N_24621);
and UO_1048 (O_1048,N_24587,N_24601);
nand UO_1049 (O_1049,N_24689,N_24534);
and UO_1050 (O_1050,N_24835,N_24722);
or UO_1051 (O_1051,N_24731,N_24906);
nor UO_1052 (O_1052,N_24571,N_24836);
or UO_1053 (O_1053,N_24628,N_24984);
xnor UO_1054 (O_1054,N_24945,N_24928);
or UO_1055 (O_1055,N_24808,N_24657);
xnor UO_1056 (O_1056,N_24897,N_24680);
xnor UO_1057 (O_1057,N_24915,N_24676);
or UO_1058 (O_1058,N_24844,N_24883);
and UO_1059 (O_1059,N_24768,N_24698);
xor UO_1060 (O_1060,N_24541,N_24946);
and UO_1061 (O_1061,N_24813,N_24786);
or UO_1062 (O_1062,N_24596,N_24519);
nor UO_1063 (O_1063,N_24593,N_24898);
and UO_1064 (O_1064,N_24909,N_24882);
nor UO_1065 (O_1065,N_24741,N_24672);
xor UO_1066 (O_1066,N_24568,N_24754);
xnor UO_1067 (O_1067,N_24602,N_24917);
nand UO_1068 (O_1068,N_24704,N_24506);
nor UO_1069 (O_1069,N_24719,N_24770);
xor UO_1070 (O_1070,N_24987,N_24540);
nand UO_1071 (O_1071,N_24527,N_24738);
xor UO_1072 (O_1072,N_24880,N_24563);
or UO_1073 (O_1073,N_24884,N_24852);
and UO_1074 (O_1074,N_24530,N_24744);
and UO_1075 (O_1075,N_24556,N_24508);
and UO_1076 (O_1076,N_24887,N_24552);
and UO_1077 (O_1077,N_24527,N_24716);
xnor UO_1078 (O_1078,N_24559,N_24979);
xnor UO_1079 (O_1079,N_24517,N_24792);
nor UO_1080 (O_1080,N_24998,N_24667);
nor UO_1081 (O_1081,N_24832,N_24938);
nor UO_1082 (O_1082,N_24672,N_24977);
xnor UO_1083 (O_1083,N_24821,N_24540);
xnor UO_1084 (O_1084,N_24725,N_24897);
xnor UO_1085 (O_1085,N_24767,N_24593);
nor UO_1086 (O_1086,N_24524,N_24838);
or UO_1087 (O_1087,N_24799,N_24956);
nor UO_1088 (O_1088,N_24587,N_24675);
nor UO_1089 (O_1089,N_24952,N_24678);
xnor UO_1090 (O_1090,N_24519,N_24938);
nor UO_1091 (O_1091,N_24905,N_24689);
nor UO_1092 (O_1092,N_24541,N_24782);
nor UO_1093 (O_1093,N_24824,N_24669);
and UO_1094 (O_1094,N_24754,N_24538);
nand UO_1095 (O_1095,N_24581,N_24785);
xnor UO_1096 (O_1096,N_24500,N_24965);
xor UO_1097 (O_1097,N_24550,N_24580);
and UO_1098 (O_1098,N_24931,N_24877);
nor UO_1099 (O_1099,N_24512,N_24831);
xnor UO_1100 (O_1100,N_24546,N_24648);
nor UO_1101 (O_1101,N_24555,N_24990);
nor UO_1102 (O_1102,N_24872,N_24864);
or UO_1103 (O_1103,N_24699,N_24780);
nor UO_1104 (O_1104,N_24624,N_24701);
nand UO_1105 (O_1105,N_24628,N_24690);
nand UO_1106 (O_1106,N_24814,N_24597);
xor UO_1107 (O_1107,N_24820,N_24683);
nand UO_1108 (O_1108,N_24691,N_24605);
and UO_1109 (O_1109,N_24971,N_24589);
nand UO_1110 (O_1110,N_24885,N_24925);
nor UO_1111 (O_1111,N_24784,N_24772);
nor UO_1112 (O_1112,N_24867,N_24952);
and UO_1113 (O_1113,N_24711,N_24671);
and UO_1114 (O_1114,N_24642,N_24583);
or UO_1115 (O_1115,N_24930,N_24972);
and UO_1116 (O_1116,N_24663,N_24922);
xnor UO_1117 (O_1117,N_24510,N_24596);
xnor UO_1118 (O_1118,N_24709,N_24501);
and UO_1119 (O_1119,N_24536,N_24738);
xor UO_1120 (O_1120,N_24720,N_24745);
or UO_1121 (O_1121,N_24553,N_24812);
xnor UO_1122 (O_1122,N_24783,N_24868);
and UO_1123 (O_1123,N_24784,N_24694);
and UO_1124 (O_1124,N_24864,N_24540);
xnor UO_1125 (O_1125,N_24716,N_24919);
and UO_1126 (O_1126,N_24747,N_24821);
nand UO_1127 (O_1127,N_24946,N_24973);
or UO_1128 (O_1128,N_24754,N_24527);
nor UO_1129 (O_1129,N_24863,N_24979);
xor UO_1130 (O_1130,N_24765,N_24599);
nor UO_1131 (O_1131,N_24978,N_24732);
nand UO_1132 (O_1132,N_24624,N_24967);
and UO_1133 (O_1133,N_24758,N_24598);
nand UO_1134 (O_1134,N_24545,N_24983);
nor UO_1135 (O_1135,N_24778,N_24722);
nand UO_1136 (O_1136,N_24999,N_24938);
or UO_1137 (O_1137,N_24510,N_24889);
and UO_1138 (O_1138,N_24800,N_24962);
nand UO_1139 (O_1139,N_24656,N_24547);
and UO_1140 (O_1140,N_24862,N_24861);
nor UO_1141 (O_1141,N_24608,N_24816);
xnor UO_1142 (O_1142,N_24904,N_24937);
xor UO_1143 (O_1143,N_24712,N_24899);
nor UO_1144 (O_1144,N_24911,N_24764);
nor UO_1145 (O_1145,N_24793,N_24900);
xnor UO_1146 (O_1146,N_24896,N_24508);
nand UO_1147 (O_1147,N_24878,N_24915);
xnor UO_1148 (O_1148,N_24999,N_24616);
nand UO_1149 (O_1149,N_24523,N_24525);
or UO_1150 (O_1150,N_24749,N_24664);
nand UO_1151 (O_1151,N_24921,N_24676);
nor UO_1152 (O_1152,N_24782,N_24613);
or UO_1153 (O_1153,N_24760,N_24635);
nand UO_1154 (O_1154,N_24605,N_24565);
nand UO_1155 (O_1155,N_24982,N_24517);
and UO_1156 (O_1156,N_24726,N_24584);
or UO_1157 (O_1157,N_24833,N_24887);
nand UO_1158 (O_1158,N_24925,N_24508);
xor UO_1159 (O_1159,N_24723,N_24740);
and UO_1160 (O_1160,N_24983,N_24844);
nand UO_1161 (O_1161,N_24712,N_24727);
or UO_1162 (O_1162,N_24595,N_24659);
or UO_1163 (O_1163,N_24824,N_24909);
or UO_1164 (O_1164,N_24929,N_24962);
xnor UO_1165 (O_1165,N_24875,N_24625);
nand UO_1166 (O_1166,N_24832,N_24752);
and UO_1167 (O_1167,N_24833,N_24982);
or UO_1168 (O_1168,N_24917,N_24779);
or UO_1169 (O_1169,N_24938,N_24800);
xnor UO_1170 (O_1170,N_24938,N_24571);
nand UO_1171 (O_1171,N_24950,N_24547);
nand UO_1172 (O_1172,N_24762,N_24612);
or UO_1173 (O_1173,N_24807,N_24794);
or UO_1174 (O_1174,N_24833,N_24922);
nand UO_1175 (O_1175,N_24530,N_24914);
and UO_1176 (O_1176,N_24810,N_24878);
and UO_1177 (O_1177,N_24809,N_24567);
xnor UO_1178 (O_1178,N_24906,N_24956);
nand UO_1179 (O_1179,N_24639,N_24673);
or UO_1180 (O_1180,N_24692,N_24906);
nor UO_1181 (O_1181,N_24779,N_24738);
and UO_1182 (O_1182,N_24949,N_24732);
nand UO_1183 (O_1183,N_24743,N_24907);
or UO_1184 (O_1184,N_24869,N_24500);
nand UO_1185 (O_1185,N_24886,N_24830);
nor UO_1186 (O_1186,N_24665,N_24905);
and UO_1187 (O_1187,N_24508,N_24958);
nor UO_1188 (O_1188,N_24583,N_24900);
nor UO_1189 (O_1189,N_24884,N_24541);
or UO_1190 (O_1190,N_24676,N_24736);
xor UO_1191 (O_1191,N_24808,N_24810);
or UO_1192 (O_1192,N_24544,N_24604);
xor UO_1193 (O_1193,N_24903,N_24504);
nand UO_1194 (O_1194,N_24739,N_24656);
and UO_1195 (O_1195,N_24845,N_24513);
nand UO_1196 (O_1196,N_24760,N_24939);
nor UO_1197 (O_1197,N_24801,N_24603);
nor UO_1198 (O_1198,N_24704,N_24898);
xnor UO_1199 (O_1199,N_24735,N_24583);
xnor UO_1200 (O_1200,N_24622,N_24846);
and UO_1201 (O_1201,N_24861,N_24832);
nand UO_1202 (O_1202,N_24964,N_24895);
nand UO_1203 (O_1203,N_24630,N_24831);
xor UO_1204 (O_1204,N_24876,N_24610);
and UO_1205 (O_1205,N_24741,N_24634);
nor UO_1206 (O_1206,N_24904,N_24923);
nor UO_1207 (O_1207,N_24730,N_24894);
xor UO_1208 (O_1208,N_24908,N_24852);
nand UO_1209 (O_1209,N_24816,N_24536);
nor UO_1210 (O_1210,N_24728,N_24894);
nand UO_1211 (O_1211,N_24554,N_24629);
xnor UO_1212 (O_1212,N_24643,N_24914);
nor UO_1213 (O_1213,N_24949,N_24609);
xnor UO_1214 (O_1214,N_24562,N_24694);
and UO_1215 (O_1215,N_24698,N_24662);
or UO_1216 (O_1216,N_24709,N_24755);
or UO_1217 (O_1217,N_24617,N_24873);
xnor UO_1218 (O_1218,N_24645,N_24912);
and UO_1219 (O_1219,N_24651,N_24806);
and UO_1220 (O_1220,N_24563,N_24920);
and UO_1221 (O_1221,N_24514,N_24671);
and UO_1222 (O_1222,N_24790,N_24904);
nand UO_1223 (O_1223,N_24744,N_24974);
nand UO_1224 (O_1224,N_24902,N_24517);
or UO_1225 (O_1225,N_24962,N_24814);
or UO_1226 (O_1226,N_24594,N_24500);
or UO_1227 (O_1227,N_24529,N_24864);
or UO_1228 (O_1228,N_24634,N_24891);
or UO_1229 (O_1229,N_24690,N_24635);
or UO_1230 (O_1230,N_24828,N_24772);
nand UO_1231 (O_1231,N_24655,N_24532);
and UO_1232 (O_1232,N_24553,N_24762);
nor UO_1233 (O_1233,N_24768,N_24634);
and UO_1234 (O_1234,N_24899,N_24653);
xor UO_1235 (O_1235,N_24504,N_24979);
nand UO_1236 (O_1236,N_24650,N_24695);
nand UO_1237 (O_1237,N_24573,N_24825);
nor UO_1238 (O_1238,N_24907,N_24527);
xor UO_1239 (O_1239,N_24749,N_24929);
nand UO_1240 (O_1240,N_24774,N_24934);
or UO_1241 (O_1241,N_24812,N_24810);
xnor UO_1242 (O_1242,N_24563,N_24749);
nand UO_1243 (O_1243,N_24500,N_24899);
nand UO_1244 (O_1244,N_24815,N_24774);
and UO_1245 (O_1245,N_24886,N_24900);
xnor UO_1246 (O_1246,N_24638,N_24997);
or UO_1247 (O_1247,N_24884,N_24708);
nand UO_1248 (O_1248,N_24956,N_24778);
nand UO_1249 (O_1249,N_24970,N_24861);
and UO_1250 (O_1250,N_24569,N_24862);
xnor UO_1251 (O_1251,N_24758,N_24509);
and UO_1252 (O_1252,N_24500,N_24885);
or UO_1253 (O_1253,N_24906,N_24671);
or UO_1254 (O_1254,N_24729,N_24544);
or UO_1255 (O_1255,N_24672,N_24604);
or UO_1256 (O_1256,N_24773,N_24996);
nor UO_1257 (O_1257,N_24571,N_24920);
nor UO_1258 (O_1258,N_24749,N_24913);
and UO_1259 (O_1259,N_24520,N_24920);
nor UO_1260 (O_1260,N_24662,N_24536);
and UO_1261 (O_1261,N_24796,N_24930);
or UO_1262 (O_1262,N_24917,N_24720);
nand UO_1263 (O_1263,N_24955,N_24653);
xnor UO_1264 (O_1264,N_24629,N_24561);
and UO_1265 (O_1265,N_24549,N_24935);
xnor UO_1266 (O_1266,N_24730,N_24974);
or UO_1267 (O_1267,N_24704,N_24724);
nand UO_1268 (O_1268,N_24887,N_24914);
nand UO_1269 (O_1269,N_24569,N_24783);
nand UO_1270 (O_1270,N_24700,N_24502);
xor UO_1271 (O_1271,N_24541,N_24516);
or UO_1272 (O_1272,N_24656,N_24604);
and UO_1273 (O_1273,N_24727,N_24811);
or UO_1274 (O_1274,N_24606,N_24703);
nand UO_1275 (O_1275,N_24947,N_24754);
nand UO_1276 (O_1276,N_24611,N_24959);
xor UO_1277 (O_1277,N_24693,N_24758);
nor UO_1278 (O_1278,N_24947,N_24972);
xnor UO_1279 (O_1279,N_24730,N_24760);
and UO_1280 (O_1280,N_24752,N_24531);
nor UO_1281 (O_1281,N_24843,N_24968);
or UO_1282 (O_1282,N_24962,N_24865);
or UO_1283 (O_1283,N_24953,N_24738);
xor UO_1284 (O_1284,N_24694,N_24739);
and UO_1285 (O_1285,N_24940,N_24725);
nor UO_1286 (O_1286,N_24699,N_24561);
xnor UO_1287 (O_1287,N_24661,N_24596);
nand UO_1288 (O_1288,N_24540,N_24550);
nor UO_1289 (O_1289,N_24764,N_24856);
xnor UO_1290 (O_1290,N_24783,N_24882);
or UO_1291 (O_1291,N_24778,N_24861);
nand UO_1292 (O_1292,N_24528,N_24891);
and UO_1293 (O_1293,N_24510,N_24776);
and UO_1294 (O_1294,N_24685,N_24537);
nand UO_1295 (O_1295,N_24656,N_24899);
and UO_1296 (O_1296,N_24915,N_24617);
nand UO_1297 (O_1297,N_24910,N_24659);
and UO_1298 (O_1298,N_24796,N_24877);
and UO_1299 (O_1299,N_24716,N_24724);
xnor UO_1300 (O_1300,N_24519,N_24567);
nand UO_1301 (O_1301,N_24760,N_24948);
xnor UO_1302 (O_1302,N_24538,N_24755);
xnor UO_1303 (O_1303,N_24795,N_24714);
nor UO_1304 (O_1304,N_24907,N_24523);
xor UO_1305 (O_1305,N_24771,N_24922);
nand UO_1306 (O_1306,N_24646,N_24761);
xor UO_1307 (O_1307,N_24908,N_24866);
and UO_1308 (O_1308,N_24945,N_24844);
or UO_1309 (O_1309,N_24851,N_24536);
and UO_1310 (O_1310,N_24596,N_24814);
and UO_1311 (O_1311,N_24963,N_24692);
nand UO_1312 (O_1312,N_24727,N_24600);
and UO_1313 (O_1313,N_24517,N_24804);
or UO_1314 (O_1314,N_24890,N_24605);
nor UO_1315 (O_1315,N_24753,N_24886);
or UO_1316 (O_1316,N_24957,N_24767);
or UO_1317 (O_1317,N_24930,N_24710);
xor UO_1318 (O_1318,N_24503,N_24645);
nor UO_1319 (O_1319,N_24884,N_24860);
xor UO_1320 (O_1320,N_24691,N_24997);
or UO_1321 (O_1321,N_24503,N_24977);
nor UO_1322 (O_1322,N_24544,N_24608);
nand UO_1323 (O_1323,N_24719,N_24678);
nor UO_1324 (O_1324,N_24539,N_24700);
nor UO_1325 (O_1325,N_24738,N_24790);
nand UO_1326 (O_1326,N_24529,N_24893);
nor UO_1327 (O_1327,N_24798,N_24570);
nand UO_1328 (O_1328,N_24766,N_24951);
or UO_1329 (O_1329,N_24576,N_24894);
or UO_1330 (O_1330,N_24916,N_24896);
and UO_1331 (O_1331,N_24970,N_24717);
nand UO_1332 (O_1332,N_24627,N_24573);
nor UO_1333 (O_1333,N_24530,N_24973);
and UO_1334 (O_1334,N_24601,N_24894);
or UO_1335 (O_1335,N_24676,N_24892);
xor UO_1336 (O_1336,N_24734,N_24661);
xor UO_1337 (O_1337,N_24827,N_24778);
nand UO_1338 (O_1338,N_24877,N_24969);
nand UO_1339 (O_1339,N_24561,N_24691);
nand UO_1340 (O_1340,N_24857,N_24625);
or UO_1341 (O_1341,N_24594,N_24922);
or UO_1342 (O_1342,N_24945,N_24603);
nand UO_1343 (O_1343,N_24985,N_24502);
nand UO_1344 (O_1344,N_24562,N_24669);
xor UO_1345 (O_1345,N_24571,N_24673);
and UO_1346 (O_1346,N_24511,N_24790);
nor UO_1347 (O_1347,N_24859,N_24959);
or UO_1348 (O_1348,N_24811,N_24620);
or UO_1349 (O_1349,N_24592,N_24974);
xor UO_1350 (O_1350,N_24655,N_24684);
or UO_1351 (O_1351,N_24733,N_24506);
or UO_1352 (O_1352,N_24671,N_24910);
xor UO_1353 (O_1353,N_24818,N_24906);
and UO_1354 (O_1354,N_24825,N_24509);
and UO_1355 (O_1355,N_24924,N_24590);
nor UO_1356 (O_1356,N_24992,N_24838);
xnor UO_1357 (O_1357,N_24668,N_24566);
nand UO_1358 (O_1358,N_24880,N_24929);
nand UO_1359 (O_1359,N_24903,N_24954);
xnor UO_1360 (O_1360,N_24733,N_24772);
xor UO_1361 (O_1361,N_24518,N_24844);
nand UO_1362 (O_1362,N_24908,N_24647);
nor UO_1363 (O_1363,N_24742,N_24695);
xor UO_1364 (O_1364,N_24632,N_24844);
and UO_1365 (O_1365,N_24747,N_24516);
nor UO_1366 (O_1366,N_24628,N_24760);
nand UO_1367 (O_1367,N_24930,N_24590);
or UO_1368 (O_1368,N_24760,N_24571);
nand UO_1369 (O_1369,N_24985,N_24877);
xor UO_1370 (O_1370,N_24704,N_24782);
nor UO_1371 (O_1371,N_24775,N_24895);
xnor UO_1372 (O_1372,N_24896,N_24812);
and UO_1373 (O_1373,N_24956,N_24687);
xnor UO_1374 (O_1374,N_24594,N_24557);
or UO_1375 (O_1375,N_24909,N_24700);
or UO_1376 (O_1376,N_24857,N_24809);
nor UO_1377 (O_1377,N_24885,N_24808);
nor UO_1378 (O_1378,N_24909,N_24669);
nor UO_1379 (O_1379,N_24797,N_24847);
nor UO_1380 (O_1380,N_24822,N_24826);
xnor UO_1381 (O_1381,N_24795,N_24666);
nand UO_1382 (O_1382,N_24876,N_24886);
nand UO_1383 (O_1383,N_24617,N_24616);
xor UO_1384 (O_1384,N_24555,N_24997);
nand UO_1385 (O_1385,N_24757,N_24810);
nor UO_1386 (O_1386,N_24602,N_24671);
nor UO_1387 (O_1387,N_24891,N_24809);
or UO_1388 (O_1388,N_24563,N_24814);
or UO_1389 (O_1389,N_24532,N_24908);
nand UO_1390 (O_1390,N_24962,N_24879);
nand UO_1391 (O_1391,N_24912,N_24749);
xnor UO_1392 (O_1392,N_24903,N_24862);
xor UO_1393 (O_1393,N_24561,N_24847);
nor UO_1394 (O_1394,N_24860,N_24663);
nand UO_1395 (O_1395,N_24614,N_24644);
and UO_1396 (O_1396,N_24777,N_24664);
and UO_1397 (O_1397,N_24500,N_24986);
or UO_1398 (O_1398,N_24558,N_24593);
nor UO_1399 (O_1399,N_24645,N_24701);
nor UO_1400 (O_1400,N_24877,N_24548);
xor UO_1401 (O_1401,N_24662,N_24844);
xnor UO_1402 (O_1402,N_24652,N_24776);
nor UO_1403 (O_1403,N_24877,N_24544);
and UO_1404 (O_1404,N_24638,N_24986);
or UO_1405 (O_1405,N_24676,N_24802);
or UO_1406 (O_1406,N_24981,N_24903);
and UO_1407 (O_1407,N_24803,N_24653);
nor UO_1408 (O_1408,N_24694,N_24613);
nor UO_1409 (O_1409,N_24558,N_24762);
or UO_1410 (O_1410,N_24504,N_24778);
xor UO_1411 (O_1411,N_24620,N_24646);
xnor UO_1412 (O_1412,N_24929,N_24731);
xnor UO_1413 (O_1413,N_24619,N_24538);
xnor UO_1414 (O_1414,N_24621,N_24773);
nand UO_1415 (O_1415,N_24855,N_24828);
or UO_1416 (O_1416,N_24507,N_24898);
nand UO_1417 (O_1417,N_24689,N_24612);
nor UO_1418 (O_1418,N_24926,N_24808);
or UO_1419 (O_1419,N_24803,N_24630);
xor UO_1420 (O_1420,N_24943,N_24817);
nand UO_1421 (O_1421,N_24948,N_24991);
or UO_1422 (O_1422,N_24709,N_24795);
nand UO_1423 (O_1423,N_24662,N_24533);
and UO_1424 (O_1424,N_24667,N_24685);
and UO_1425 (O_1425,N_24718,N_24905);
xor UO_1426 (O_1426,N_24534,N_24716);
and UO_1427 (O_1427,N_24615,N_24743);
or UO_1428 (O_1428,N_24991,N_24766);
and UO_1429 (O_1429,N_24523,N_24891);
nor UO_1430 (O_1430,N_24557,N_24900);
or UO_1431 (O_1431,N_24531,N_24622);
and UO_1432 (O_1432,N_24532,N_24851);
nor UO_1433 (O_1433,N_24632,N_24831);
and UO_1434 (O_1434,N_24829,N_24873);
nor UO_1435 (O_1435,N_24509,N_24944);
and UO_1436 (O_1436,N_24620,N_24870);
and UO_1437 (O_1437,N_24636,N_24924);
or UO_1438 (O_1438,N_24827,N_24989);
and UO_1439 (O_1439,N_24810,N_24949);
xor UO_1440 (O_1440,N_24788,N_24753);
nand UO_1441 (O_1441,N_24834,N_24908);
nor UO_1442 (O_1442,N_24628,N_24733);
nand UO_1443 (O_1443,N_24576,N_24812);
and UO_1444 (O_1444,N_24745,N_24923);
nor UO_1445 (O_1445,N_24936,N_24748);
xnor UO_1446 (O_1446,N_24997,N_24558);
nand UO_1447 (O_1447,N_24723,N_24808);
and UO_1448 (O_1448,N_24999,N_24714);
nand UO_1449 (O_1449,N_24590,N_24921);
and UO_1450 (O_1450,N_24742,N_24705);
xor UO_1451 (O_1451,N_24871,N_24547);
and UO_1452 (O_1452,N_24910,N_24739);
xnor UO_1453 (O_1453,N_24659,N_24889);
or UO_1454 (O_1454,N_24610,N_24825);
nand UO_1455 (O_1455,N_24990,N_24968);
nor UO_1456 (O_1456,N_24788,N_24666);
nor UO_1457 (O_1457,N_24527,N_24693);
and UO_1458 (O_1458,N_24663,N_24534);
or UO_1459 (O_1459,N_24905,N_24556);
and UO_1460 (O_1460,N_24647,N_24793);
nor UO_1461 (O_1461,N_24644,N_24593);
and UO_1462 (O_1462,N_24573,N_24554);
or UO_1463 (O_1463,N_24660,N_24867);
xnor UO_1464 (O_1464,N_24930,N_24806);
xnor UO_1465 (O_1465,N_24694,N_24624);
and UO_1466 (O_1466,N_24531,N_24916);
xor UO_1467 (O_1467,N_24909,N_24777);
nand UO_1468 (O_1468,N_24967,N_24632);
xnor UO_1469 (O_1469,N_24830,N_24745);
and UO_1470 (O_1470,N_24940,N_24717);
nand UO_1471 (O_1471,N_24585,N_24640);
nor UO_1472 (O_1472,N_24633,N_24928);
and UO_1473 (O_1473,N_24639,N_24625);
and UO_1474 (O_1474,N_24736,N_24859);
xor UO_1475 (O_1475,N_24624,N_24505);
and UO_1476 (O_1476,N_24924,N_24541);
nor UO_1477 (O_1477,N_24963,N_24784);
and UO_1478 (O_1478,N_24632,N_24788);
and UO_1479 (O_1479,N_24855,N_24568);
and UO_1480 (O_1480,N_24690,N_24776);
xnor UO_1481 (O_1481,N_24783,N_24749);
xor UO_1482 (O_1482,N_24903,N_24527);
or UO_1483 (O_1483,N_24970,N_24799);
nor UO_1484 (O_1484,N_24583,N_24619);
nor UO_1485 (O_1485,N_24617,N_24726);
and UO_1486 (O_1486,N_24787,N_24617);
xor UO_1487 (O_1487,N_24896,N_24823);
xnor UO_1488 (O_1488,N_24628,N_24761);
nand UO_1489 (O_1489,N_24944,N_24704);
nand UO_1490 (O_1490,N_24849,N_24892);
nor UO_1491 (O_1491,N_24928,N_24732);
and UO_1492 (O_1492,N_24573,N_24505);
or UO_1493 (O_1493,N_24646,N_24823);
and UO_1494 (O_1494,N_24562,N_24812);
or UO_1495 (O_1495,N_24990,N_24812);
nor UO_1496 (O_1496,N_24532,N_24982);
xnor UO_1497 (O_1497,N_24827,N_24781);
and UO_1498 (O_1498,N_24696,N_24721);
nand UO_1499 (O_1499,N_24694,N_24941);
and UO_1500 (O_1500,N_24682,N_24878);
nand UO_1501 (O_1501,N_24558,N_24698);
xnor UO_1502 (O_1502,N_24579,N_24634);
nor UO_1503 (O_1503,N_24705,N_24832);
xnor UO_1504 (O_1504,N_24780,N_24501);
or UO_1505 (O_1505,N_24960,N_24654);
and UO_1506 (O_1506,N_24588,N_24901);
nand UO_1507 (O_1507,N_24693,N_24871);
and UO_1508 (O_1508,N_24652,N_24958);
nand UO_1509 (O_1509,N_24845,N_24818);
xor UO_1510 (O_1510,N_24956,N_24960);
nand UO_1511 (O_1511,N_24846,N_24593);
nand UO_1512 (O_1512,N_24532,N_24813);
or UO_1513 (O_1513,N_24867,N_24708);
xnor UO_1514 (O_1514,N_24944,N_24574);
or UO_1515 (O_1515,N_24648,N_24563);
xnor UO_1516 (O_1516,N_24702,N_24518);
nand UO_1517 (O_1517,N_24945,N_24688);
and UO_1518 (O_1518,N_24972,N_24638);
or UO_1519 (O_1519,N_24739,N_24762);
xnor UO_1520 (O_1520,N_24866,N_24844);
nand UO_1521 (O_1521,N_24806,N_24855);
or UO_1522 (O_1522,N_24740,N_24927);
or UO_1523 (O_1523,N_24893,N_24542);
nand UO_1524 (O_1524,N_24645,N_24735);
nand UO_1525 (O_1525,N_24881,N_24770);
nand UO_1526 (O_1526,N_24929,N_24994);
nand UO_1527 (O_1527,N_24509,N_24591);
or UO_1528 (O_1528,N_24963,N_24543);
and UO_1529 (O_1529,N_24827,N_24724);
or UO_1530 (O_1530,N_24940,N_24650);
and UO_1531 (O_1531,N_24673,N_24549);
nor UO_1532 (O_1532,N_24532,N_24578);
nand UO_1533 (O_1533,N_24993,N_24765);
or UO_1534 (O_1534,N_24704,N_24584);
nor UO_1535 (O_1535,N_24947,N_24547);
nor UO_1536 (O_1536,N_24568,N_24659);
or UO_1537 (O_1537,N_24541,N_24687);
nand UO_1538 (O_1538,N_24815,N_24658);
and UO_1539 (O_1539,N_24641,N_24797);
nand UO_1540 (O_1540,N_24722,N_24689);
or UO_1541 (O_1541,N_24837,N_24531);
nor UO_1542 (O_1542,N_24895,N_24816);
xnor UO_1543 (O_1543,N_24725,N_24659);
xnor UO_1544 (O_1544,N_24696,N_24647);
xor UO_1545 (O_1545,N_24827,N_24679);
and UO_1546 (O_1546,N_24826,N_24514);
or UO_1547 (O_1547,N_24820,N_24734);
and UO_1548 (O_1548,N_24910,N_24575);
and UO_1549 (O_1549,N_24809,N_24633);
and UO_1550 (O_1550,N_24681,N_24619);
xnor UO_1551 (O_1551,N_24842,N_24524);
or UO_1552 (O_1552,N_24915,N_24978);
nand UO_1553 (O_1553,N_24987,N_24791);
nand UO_1554 (O_1554,N_24941,N_24986);
xnor UO_1555 (O_1555,N_24631,N_24831);
nor UO_1556 (O_1556,N_24930,N_24515);
and UO_1557 (O_1557,N_24896,N_24541);
nand UO_1558 (O_1558,N_24887,N_24658);
or UO_1559 (O_1559,N_24960,N_24950);
nand UO_1560 (O_1560,N_24981,N_24759);
xnor UO_1561 (O_1561,N_24582,N_24912);
nand UO_1562 (O_1562,N_24840,N_24531);
or UO_1563 (O_1563,N_24805,N_24568);
xor UO_1564 (O_1564,N_24638,N_24868);
xnor UO_1565 (O_1565,N_24562,N_24738);
xor UO_1566 (O_1566,N_24751,N_24738);
xor UO_1567 (O_1567,N_24582,N_24929);
nand UO_1568 (O_1568,N_24509,N_24830);
nand UO_1569 (O_1569,N_24866,N_24606);
nor UO_1570 (O_1570,N_24559,N_24672);
xnor UO_1571 (O_1571,N_24887,N_24675);
and UO_1572 (O_1572,N_24919,N_24517);
xor UO_1573 (O_1573,N_24575,N_24639);
nand UO_1574 (O_1574,N_24908,N_24673);
or UO_1575 (O_1575,N_24875,N_24869);
nor UO_1576 (O_1576,N_24734,N_24860);
nand UO_1577 (O_1577,N_24929,N_24541);
and UO_1578 (O_1578,N_24705,N_24945);
xor UO_1579 (O_1579,N_24973,N_24803);
nor UO_1580 (O_1580,N_24583,N_24971);
or UO_1581 (O_1581,N_24921,N_24555);
and UO_1582 (O_1582,N_24956,N_24920);
xor UO_1583 (O_1583,N_24611,N_24739);
nand UO_1584 (O_1584,N_24565,N_24803);
xor UO_1585 (O_1585,N_24839,N_24867);
nor UO_1586 (O_1586,N_24946,N_24625);
and UO_1587 (O_1587,N_24994,N_24545);
nor UO_1588 (O_1588,N_24866,N_24781);
nor UO_1589 (O_1589,N_24889,N_24699);
and UO_1590 (O_1590,N_24941,N_24826);
xnor UO_1591 (O_1591,N_24676,N_24951);
nor UO_1592 (O_1592,N_24814,N_24652);
or UO_1593 (O_1593,N_24961,N_24828);
or UO_1594 (O_1594,N_24751,N_24699);
or UO_1595 (O_1595,N_24913,N_24769);
nor UO_1596 (O_1596,N_24901,N_24687);
xnor UO_1597 (O_1597,N_24620,N_24515);
nand UO_1598 (O_1598,N_24975,N_24505);
or UO_1599 (O_1599,N_24706,N_24628);
and UO_1600 (O_1600,N_24575,N_24509);
xor UO_1601 (O_1601,N_24828,N_24969);
nand UO_1602 (O_1602,N_24896,N_24581);
xnor UO_1603 (O_1603,N_24542,N_24682);
or UO_1604 (O_1604,N_24979,N_24753);
xnor UO_1605 (O_1605,N_24966,N_24765);
nand UO_1606 (O_1606,N_24768,N_24570);
and UO_1607 (O_1607,N_24587,N_24727);
and UO_1608 (O_1608,N_24929,N_24827);
or UO_1609 (O_1609,N_24706,N_24971);
nor UO_1610 (O_1610,N_24726,N_24951);
xnor UO_1611 (O_1611,N_24592,N_24620);
or UO_1612 (O_1612,N_24553,N_24563);
and UO_1613 (O_1613,N_24877,N_24567);
nand UO_1614 (O_1614,N_24621,N_24671);
and UO_1615 (O_1615,N_24648,N_24696);
and UO_1616 (O_1616,N_24963,N_24910);
and UO_1617 (O_1617,N_24538,N_24609);
and UO_1618 (O_1618,N_24642,N_24854);
and UO_1619 (O_1619,N_24718,N_24889);
xor UO_1620 (O_1620,N_24501,N_24782);
nand UO_1621 (O_1621,N_24853,N_24550);
and UO_1622 (O_1622,N_24719,N_24524);
nor UO_1623 (O_1623,N_24888,N_24987);
nor UO_1624 (O_1624,N_24841,N_24996);
nor UO_1625 (O_1625,N_24731,N_24707);
nor UO_1626 (O_1626,N_24508,N_24689);
and UO_1627 (O_1627,N_24962,N_24997);
nor UO_1628 (O_1628,N_24865,N_24562);
xnor UO_1629 (O_1629,N_24614,N_24711);
nor UO_1630 (O_1630,N_24632,N_24760);
nand UO_1631 (O_1631,N_24504,N_24927);
and UO_1632 (O_1632,N_24929,N_24975);
xor UO_1633 (O_1633,N_24624,N_24888);
nand UO_1634 (O_1634,N_24984,N_24518);
xor UO_1635 (O_1635,N_24631,N_24855);
xor UO_1636 (O_1636,N_24956,N_24891);
xnor UO_1637 (O_1637,N_24586,N_24543);
or UO_1638 (O_1638,N_24856,N_24611);
nand UO_1639 (O_1639,N_24854,N_24702);
nor UO_1640 (O_1640,N_24595,N_24507);
xnor UO_1641 (O_1641,N_24578,N_24607);
xnor UO_1642 (O_1642,N_24551,N_24664);
and UO_1643 (O_1643,N_24679,N_24634);
nor UO_1644 (O_1644,N_24500,N_24509);
or UO_1645 (O_1645,N_24890,N_24840);
xnor UO_1646 (O_1646,N_24988,N_24947);
nor UO_1647 (O_1647,N_24542,N_24817);
or UO_1648 (O_1648,N_24598,N_24834);
nor UO_1649 (O_1649,N_24583,N_24718);
xnor UO_1650 (O_1650,N_24995,N_24840);
nor UO_1651 (O_1651,N_24509,N_24652);
xor UO_1652 (O_1652,N_24614,N_24986);
xnor UO_1653 (O_1653,N_24707,N_24589);
xnor UO_1654 (O_1654,N_24677,N_24842);
nand UO_1655 (O_1655,N_24828,N_24714);
or UO_1656 (O_1656,N_24737,N_24979);
xor UO_1657 (O_1657,N_24832,N_24935);
or UO_1658 (O_1658,N_24934,N_24854);
nand UO_1659 (O_1659,N_24698,N_24552);
or UO_1660 (O_1660,N_24583,N_24965);
nor UO_1661 (O_1661,N_24658,N_24848);
or UO_1662 (O_1662,N_24874,N_24859);
or UO_1663 (O_1663,N_24728,N_24867);
xnor UO_1664 (O_1664,N_24944,N_24633);
and UO_1665 (O_1665,N_24637,N_24866);
nor UO_1666 (O_1666,N_24688,N_24921);
xnor UO_1667 (O_1667,N_24798,N_24914);
and UO_1668 (O_1668,N_24607,N_24791);
xor UO_1669 (O_1669,N_24692,N_24754);
and UO_1670 (O_1670,N_24554,N_24746);
or UO_1671 (O_1671,N_24923,N_24829);
nor UO_1672 (O_1672,N_24922,N_24658);
xor UO_1673 (O_1673,N_24654,N_24952);
and UO_1674 (O_1674,N_24959,N_24911);
xor UO_1675 (O_1675,N_24598,N_24868);
xnor UO_1676 (O_1676,N_24828,N_24884);
xor UO_1677 (O_1677,N_24624,N_24745);
and UO_1678 (O_1678,N_24723,N_24872);
xor UO_1679 (O_1679,N_24521,N_24585);
and UO_1680 (O_1680,N_24565,N_24601);
nor UO_1681 (O_1681,N_24648,N_24736);
or UO_1682 (O_1682,N_24842,N_24753);
xnor UO_1683 (O_1683,N_24718,N_24552);
nand UO_1684 (O_1684,N_24947,N_24860);
nand UO_1685 (O_1685,N_24776,N_24535);
nand UO_1686 (O_1686,N_24738,N_24952);
and UO_1687 (O_1687,N_24916,N_24732);
nor UO_1688 (O_1688,N_24606,N_24812);
and UO_1689 (O_1689,N_24829,N_24716);
nor UO_1690 (O_1690,N_24691,N_24728);
nor UO_1691 (O_1691,N_24828,N_24730);
and UO_1692 (O_1692,N_24884,N_24773);
nand UO_1693 (O_1693,N_24850,N_24761);
and UO_1694 (O_1694,N_24718,N_24743);
xor UO_1695 (O_1695,N_24723,N_24606);
and UO_1696 (O_1696,N_24774,N_24960);
nor UO_1697 (O_1697,N_24903,N_24971);
and UO_1698 (O_1698,N_24928,N_24804);
and UO_1699 (O_1699,N_24506,N_24769);
nor UO_1700 (O_1700,N_24843,N_24809);
and UO_1701 (O_1701,N_24712,N_24608);
and UO_1702 (O_1702,N_24784,N_24576);
nand UO_1703 (O_1703,N_24708,N_24838);
nor UO_1704 (O_1704,N_24511,N_24747);
nand UO_1705 (O_1705,N_24650,N_24776);
nand UO_1706 (O_1706,N_24691,N_24782);
nand UO_1707 (O_1707,N_24647,N_24823);
xnor UO_1708 (O_1708,N_24871,N_24869);
nor UO_1709 (O_1709,N_24710,N_24636);
or UO_1710 (O_1710,N_24740,N_24891);
nand UO_1711 (O_1711,N_24753,N_24772);
nor UO_1712 (O_1712,N_24591,N_24815);
xor UO_1713 (O_1713,N_24763,N_24546);
and UO_1714 (O_1714,N_24512,N_24672);
nand UO_1715 (O_1715,N_24985,N_24633);
and UO_1716 (O_1716,N_24801,N_24680);
and UO_1717 (O_1717,N_24826,N_24800);
or UO_1718 (O_1718,N_24937,N_24747);
or UO_1719 (O_1719,N_24893,N_24864);
or UO_1720 (O_1720,N_24939,N_24904);
or UO_1721 (O_1721,N_24578,N_24604);
xnor UO_1722 (O_1722,N_24793,N_24815);
nor UO_1723 (O_1723,N_24534,N_24946);
nand UO_1724 (O_1724,N_24812,N_24853);
or UO_1725 (O_1725,N_24846,N_24713);
nor UO_1726 (O_1726,N_24946,N_24572);
nand UO_1727 (O_1727,N_24948,N_24865);
or UO_1728 (O_1728,N_24865,N_24967);
and UO_1729 (O_1729,N_24554,N_24786);
nor UO_1730 (O_1730,N_24836,N_24840);
or UO_1731 (O_1731,N_24895,N_24911);
or UO_1732 (O_1732,N_24574,N_24897);
and UO_1733 (O_1733,N_24796,N_24668);
and UO_1734 (O_1734,N_24962,N_24878);
xnor UO_1735 (O_1735,N_24809,N_24946);
or UO_1736 (O_1736,N_24722,N_24535);
or UO_1737 (O_1737,N_24998,N_24861);
and UO_1738 (O_1738,N_24961,N_24937);
and UO_1739 (O_1739,N_24582,N_24902);
nor UO_1740 (O_1740,N_24683,N_24736);
xor UO_1741 (O_1741,N_24676,N_24872);
and UO_1742 (O_1742,N_24908,N_24806);
nand UO_1743 (O_1743,N_24562,N_24595);
nand UO_1744 (O_1744,N_24932,N_24725);
nand UO_1745 (O_1745,N_24933,N_24722);
or UO_1746 (O_1746,N_24697,N_24720);
or UO_1747 (O_1747,N_24604,N_24756);
nand UO_1748 (O_1748,N_24817,N_24882);
nand UO_1749 (O_1749,N_24721,N_24598);
nor UO_1750 (O_1750,N_24995,N_24753);
and UO_1751 (O_1751,N_24907,N_24859);
and UO_1752 (O_1752,N_24538,N_24691);
or UO_1753 (O_1753,N_24713,N_24513);
or UO_1754 (O_1754,N_24976,N_24842);
nand UO_1755 (O_1755,N_24567,N_24835);
nor UO_1756 (O_1756,N_24795,N_24839);
xor UO_1757 (O_1757,N_24534,N_24530);
nor UO_1758 (O_1758,N_24882,N_24522);
or UO_1759 (O_1759,N_24788,N_24541);
nand UO_1760 (O_1760,N_24731,N_24613);
and UO_1761 (O_1761,N_24504,N_24842);
nor UO_1762 (O_1762,N_24755,N_24862);
or UO_1763 (O_1763,N_24919,N_24878);
or UO_1764 (O_1764,N_24807,N_24639);
or UO_1765 (O_1765,N_24652,N_24602);
nor UO_1766 (O_1766,N_24502,N_24587);
and UO_1767 (O_1767,N_24558,N_24908);
or UO_1768 (O_1768,N_24711,N_24592);
xor UO_1769 (O_1769,N_24685,N_24580);
nor UO_1770 (O_1770,N_24613,N_24791);
xor UO_1771 (O_1771,N_24902,N_24877);
or UO_1772 (O_1772,N_24631,N_24791);
and UO_1773 (O_1773,N_24719,N_24671);
xnor UO_1774 (O_1774,N_24993,N_24952);
and UO_1775 (O_1775,N_24649,N_24568);
nor UO_1776 (O_1776,N_24546,N_24590);
xor UO_1777 (O_1777,N_24646,N_24914);
nor UO_1778 (O_1778,N_24722,N_24591);
or UO_1779 (O_1779,N_24663,N_24655);
xnor UO_1780 (O_1780,N_24920,N_24560);
nor UO_1781 (O_1781,N_24635,N_24586);
xnor UO_1782 (O_1782,N_24740,N_24998);
nand UO_1783 (O_1783,N_24981,N_24993);
xnor UO_1784 (O_1784,N_24635,N_24546);
xor UO_1785 (O_1785,N_24974,N_24761);
xnor UO_1786 (O_1786,N_24967,N_24697);
nor UO_1787 (O_1787,N_24585,N_24777);
xor UO_1788 (O_1788,N_24977,N_24526);
xor UO_1789 (O_1789,N_24866,N_24515);
nor UO_1790 (O_1790,N_24805,N_24598);
or UO_1791 (O_1791,N_24805,N_24814);
nor UO_1792 (O_1792,N_24860,N_24829);
and UO_1793 (O_1793,N_24951,N_24687);
nand UO_1794 (O_1794,N_24684,N_24942);
and UO_1795 (O_1795,N_24970,N_24554);
nor UO_1796 (O_1796,N_24605,N_24849);
nand UO_1797 (O_1797,N_24989,N_24808);
nor UO_1798 (O_1798,N_24520,N_24749);
nor UO_1799 (O_1799,N_24641,N_24847);
nor UO_1800 (O_1800,N_24767,N_24885);
or UO_1801 (O_1801,N_24966,N_24703);
or UO_1802 (O_1802,N_24782,N_24570);
or UO_1803 (O_1803,N_24821,N_24999);
or UO_1804 (O_1804,N_24882,N_24811);
xnor UO_1805 (O_1805,N_24795,N_24837);
nand UO_1806 (O_1806,N_24878,N_24750);
nand UO_1807 (O_1807,N_24929,N_24898);
and UO_1808 (O_1808,N_24960,N_24579);
xor UO_1809 (O_1809,N_24542,N_24551);
xor UO_1810 (O_1810,N_24785,N_24666);
and UO_1811 (O_1811,N_24903,N_24946);
nor UO_1812 (O_1812,N_24835,N_24728);
nor UO_1813 (O_1813,N_24962,N_24649);
and UO_1814 (O_1814,N_24596,N_24679);
nand UO_1815 (O_1815,N_24967,N_24845);
xor UO_1816 (O_1816,N_24775,N_24559);
nand UO_1817 (O_1817,N_24685,N_24977);
nand UO_1818 (O_1818,N_24954,N_24556);
xor UO_1819 (O_1819,N_24575,N_24856);
xor UO_1820 (O_1820,N_24832,N_24972);
or UO_1821 (O_1821,N_24621,N_24631);
and UO_1822 (O_1822,N_24562,N_24944);
nand UO_1823 (O_1823,N_24658,N_24993);
nor UO_1824 (O_1824,N_24812,N_24848);
nor UO_1825 (O_1825,N_24998,N_24794);
nand UO_1826 (O_1826,N_24551,N_24507);
nor UO_1827 (O_1827,N_24891,N_24683);
and UO_1828 (O_1828,N_24531,N_24530);
and UO_1829 (O_1829,N_24953,N_24697);
or UO_1830 (O_1830,N_24986,N_24603);
nand UO_1831 (O_1831,N_24843,N_24994);
and UO_1832 (O_1832,N_24966,N_24956);
nand UO_1833 (O_1833,N_24862,N_24682);
and UO_1834 (O_1834,N_24963,N_24667);
nor UO_1835 (O_1835,N_24717,N_24682);
xor UO_1836 (O_1836,N_24882,N_24822);
xnor UO_1837 (O_1837,N_24801,N_24750);
xor UO_1838 (O_1838,N_24609,N_24681);
and UO_1839 (O_1839,N_24757,N_24596);
or UO_1840 (O_1840,N_24817,N_24806);
xnor UO_1841 (O_1841,N_24713,N_24796);
nand UO_1842 (O_1842,N_24683,N_24772);
nor UO_1843 (O_1843,N_24754,N_24780);
nand UO_1844 (O_1844,N_24884,N_24922);
nand UO_1845 (O_1845,N_24895,N_24760);
or UO_1846 (O_1846,N_24848,N_24864);
or UO_1847 (O_1847,N_24665,N_24881);
nor UO_1848 (O_1848,N_24969,N_24533);
or UO_1849 (O_1849,N_24529,N_24871);
nand UO_1850 (O_1850,N_24968,N_24527);
nand UO_1851 (O_1851,N_24823,N_24573);
nand UO_1852 (O_1852,N_24751,N_24737);
nor UO_1853 (O_1853,N_24702,N_24558);
nand UO_1854 (O_1854,N_24967,N_24965);
and UO_1855 (O_1855,N_24893,N_24846);
nand UO_1856 (O_1856,N_24861,N_24827);
nor UO_1857 (O_1857,N_24908,N_24570);
and UO_1858 (O_1858,N_24586,N_24829);
or UO_1859 (O_1859,N_24662,N_24531);
or UO_1860 (O_1860,N_24801,N_24687);
and UO_1861 (O_1861,N_24573,N_24670);
xnor UO_1862 (O_1862,N_24845,N_24836);
or UO_1863 (O_1863,N_24823,N_24782);
and UO_1864 (O_1864,N_24770,N_24577);
or UO_1865 (O_1865,N_24615,N_24848);
nand UO_1866 (O_1866,N_24978,N_24678);
nand UO_1867 (O_1867,N_24601,N_24796);
or UO_1868 (O_1868,N_24927,N_24694);
nand UO_1869 (O_1869,N_24924,N_24978);
nor UO_1870 (O_1870,N_24943,N_24987);
or UO_1871 (O_1871,N_24915,N_24546);
nand UO_1872 (O_1872,N_24890,N_24996);
or UO_1873 (O_1873,N_24664,N_24617);
nand UO_1874 (O_1874,N_24943,N_24860);
xor UO_1875 (O_1875,N_24664,N_24707);
xnor UO_1876 (O_1876,N_24509,N_24998);
nand UO_1877 (O_1877,N_24826,N_24933);
or UO_1878 (O_1878,N_24903,N_24673);
nand UO_1879 (O_1879,N_24894,N_24510);
nor UO_1880 (O_1880,N_24867,N_24876);
and UO_1881 (O_1881,N_24796,N_24574);
and UO_1882 (O_1882,N_24708,N_24689);
or UO_1883 (O_1883,N_24697,N_24629);
xor UO_1884 (O_1884,N_24645,N_24637);
nand UO_1885 (O_1885,N_24620,N_24682);
xnor UO_1886 (O_1886,N_24526,N_24610);
and UO_1887 (O_1887,N_24640,N_24936);
nor UO_1888 (O_1888,N_24926,N_24925);
xnor UO_1889 (O_1889,N_24842,N_24832);
xor UO_1890 (O_1890,N_24623,N_24869);
nor UO_1891 (O_1891,N_24824,N_24887);
and UO_1892 (O_1892,N_24991,N_24530);
or UO_1893 (O_1893,N_24669,N_24525);
and UO_1894 (O_1894,N_24547,N_24843);
nand UO_1895 (O_1895,N_24779,N_24752);
nand UO_1896 (O_1896,N_24875,N_24872);
nand UO_1897 (O_1897,N_24645,N_24811);
nand UO_1898 (O_1898,N_24572,N_24702);
xor UO_1899 (O_1899,N_24692,N_24607);
and UO_1900 (O_1900,N_24613,N_24539);
and UO_1901 (O_1901,N_24974,N_24503);
nand UO_1902 (O_1902,N_24854,N_24929);
nor UO_1903 (O_1903,N_24894,N_24776);
and UO_1904 (O_1904,N_24683,N_24650);
and UO_1905 (O_1905,N_24603,N_24626);
xnor UO_1906 (O_1906,N_24736,N_24605);
xnor UO_1907 (O_1907,N_24517,N_24928);
nor UO_1908 (O_1908,N_24559,N_24712);
xor UO_1909 (O_1909,N_24562,N_24520);
and UO_1910 (O_1910,N_24997,N_24821);
nor UO_1911 (O_1911,N_24786,N_24628);
nand UO_1912 (O_1912,N_24642,N_24754);
xor UO_1913 (O_1913,N_24815,N_24877);
nand UO_1914 (O_1914,N_24962,N_24905);
nor UO_1915 (O_1915,N_24626,N_24790);
nand UO_1916 (O_1916,N_24655,N_24850);
or UO_1917 (O_1917,N_24751,N_24744);
xnor UO_1918 (O_1918,N_24622,N_24560);
xnor UO_1919 (O_1919,N_24981,N_24758);
nand UO_1920 (O_1920,N_24757,N_24914);
and UO_1921 (O_1921,N_24603,N_24816);
and UO_1922 (O_1922,N_24814,N_24808);
and UO_1923 (O_1923,N_24569,N_24584);
or UO_1924 (O_1924,N_24811,N_24940);
nand UO_1925 (O_1925,N_24832,N_24787);
nor UO_1926 (O_1926,N_24635,N_24625);
nor UO_1927 (O_1927,N_24988,N_24537);
nand UO_1928 (O_1928,N_24558,N_24978);
nand UO_1929 (O_1929,N_24569,N_24537);
or UO_1930 (O_1930,N_24559,N_24862);
nor UO_1931 (O_1931,N_24575,N_24690);
nor UO_1932 (O_1932,N_24612,N_24502);
and UO_1933 (O_1933,N_24760,N_24793);
and UO_1934 (O_1934,N_24899,N_24764);
and UO_1935 (O_1935,N_24781,N_24692);
xnor UO_1936 (O_1936,N_24739,N_24783);
or UO_1937 (O_1937,N_24670,N_24866);
and UO_1938 (O_1938,N_24636,N_24592);
or UO_1939 (O_1939,N_24687,N_24756);
and UO_1940 (O_1940,N_24545,N_24831);
nor UO_1941 (O_1941,N_24654,N_24755);
and UO_1942 (O_1942,N_24903,N_24624);
nand UO_1943 (O_1943,N_24784,N_24974);
and UO_1944 (O_1944,N_24791,N_24708);
xnor UO_1945 (O_1945,N_24732,N_24957);
nor UO_1946 (O_1946,N_24943,N_24759);
nand UO_1947 (O_1947,N_24909,N_24790);
xnor UO_1948 (O_1948,N_24786,N_24818);
or UO_1949 (O_1949,N_24968,N_24799);
or UO_1950 (O_1950,N_24972,N_24559);
and UO_1951 (O_1951,N_24729,N_24963);
or UO_1952 (O_1952,N_24732,N_24562);
nand UO_1953 (O_1953,N_24764,N_24627);
and UO_1954 (O_1954,N_24603,N_24823);
xnor UO_1955 (O_1955,N_24662,N_24508);
and UO_1956 (O_1956,N_24522,N_24561);
xnor UO_1957 (O_1957,N_24622,N_24553);
nor UO_1958 (O_1958,N_24534,N_24583);
xnor UO_1959 (O_1959,N_24655,N_24781);
and UO_1960 (O_1960,N_24717,N_24789);
and UO_1961 (O_1961,N_24585,N_24629);
or UO_1962 (O_1962,N_24711,N_24725);
and UO_1963 (O_1963,N_24868,N_24554);
xnor UO_1964 (O_1964,N_24835,N_24596);
or UO_1965 (O_1965,N_24545,N_24901);
nor UO_1966 (O_1966,N_24979,N_24688);
nor UO_1967 (O_1967,N_24749,N_24739);
nand UO_1968 (O_1968,N_24783,N_24517);
nand UO_1969 (O_1969,N_24985,N_24954);
nor UO_1970 (O_1970,N_24877,N_24947);
nor UO_1971 (O_1971,N_24573,N_24977);
nand UO_1972 (O_1972,N_24683,N_24748);
nand UO_1973 (O_1973,N_24857,N_24630);
nor UO_1974 (O_1974,N_24887,N_24817);
and UO_1975 (O_1975,N_24508,N_24851);
nand UO_1976 (O_1976,N_24980,N_24528);
nor UO_1977 (O_1977,N_24897,N_24612);
or UO_1978 (O_1978,N_24951,N_24793);
xnor UO_1979 (O_1979,N_24958,N_24916);
or UO_1980 (O_1980,N_24880,N_24584);
nand UO_1981 (O_1981,N_24676,N_24993);
or UO_1982 (O_1982,N_24862,N_24920);
nand UO_1983 (O_1983,N_24656,N_24559);
nand UO_1984 (O_1984,N_24608,N_24622);
xnor UO_1985 (O_1985,N_24902,N_24924);
nand UO_1986 (O_1986,N_24872,N_24898);
nand UO_1987 (O_1987,N_24976,N_24970);
nand UO_1988 (O_1988,N_24994,N_24629);
and UO_1989 (O_1989,N_24784,N_24511);
xor UO_1990 (O_1990,N_24928,N_24996);
nor UO_1991 (O_1991,N_24996,N_24525);
nand UO_1992 (O_1992,N_24911,N_24748);
xor UO_1993 (O_1993,N_24537,N_24545);
nor UO_1994 (O_1994,N_24968,N_24937);
or UO_1995 (O_1995,N_24843,N_24868);
nor UO_1996 (O_1996,N_24630,N_24946);
or UO_1997 (O_1997,N_24964,N_24731);
and UO_1998 (O_1998,N_24831,N_24778);
nor UO_1999 (O_1999,N_24994,N_24644);
nand UO_2000 (O_2000,N_24603,N_24853);
nor UO_2001 (O_2001,N_24707,N_24882);
xnor UO_2002 (O_2002,N_24930,N_24695);
xor UO_2003 (O_2003,N_24802,N_24839);
nor UO_2004 (O_2004,N_24932,N_24794);
nor UO_2005 (O_2005,N_24862,N_24768);
or UO_2006 (O_2006,N_24685,N_24725);
and UO_2007 (O_2007,N_24929,N_24925);
and UO_2008 (O_2008,N_24877,N_24913);
and UO_2009 (O_2009,N_24843,N_24674);
or UO_2010 (O_2010,N_24875,N_24710);
nor UO_2011 (O_2011,N_24907,N_24740);
nor UO_2012 (O_2012,N_24802,N_24781);
and UO_2013 (O_2013,N_24677,N_24752);
nand UO_2014 (O_2014,N_24740,N_24837);
and UO_2015 (O_2015,N_24536,N_24593);
and UO_2016 (O_2016,N_24573,N_24921);
or UO_2017 (O_2017,N_24907,N_24945);
xor UO_2018 (O_2018,N_24661,N_24923);
and UO_2019 (O_2019,N_24746,N_24670);
or UO_2020 (O_2020,N_24575,N_24842);
or UO_2021 (O_2021,N_24658,N_24648);
and UO_2022 (O_2022,N_24819,N_24753);
nor UO_2023 (O_2023,N_24509,N_24531);
nand UO_2024 (O_2024,N_24767,N_24623);
or UO_2025 (O_2025,N_24956,N_24952);
and UO_2026 (O_2026,N_24732,N_24631);
or UO_2027 (O_2027,N_24637,N_24978);
or UO_2028 (O_2028,N_24611,N_24566);
nor UO_2029 (O_2029,N_24527,N_24604);
nand UO_2030 (O_2030,N_24974,N_24971);
or UO_2031 (O_2031,N_24879,N_24667);
nand UO_2032 (O_2032,N_24792,N_24690);
xor UO_2033 (O_2033,N_24627,N_24625);
and UO_2034 (O_2034,N_24908,N_24549);
or UO_2035 (O_2035,N_24753,N_24659);
xnor UO_2036 (O_2036,N_24804,N_24596);
or UO_2037 (O_2037,N_24738,N_24960);
nor UO_2038 (O_2038,N_24998,N_24986);
and UO_2039 (O_2039,N_24620,N_24506);
xor UO_2040 (O_2040,N_24637,N_24921);
and UO_2041 (O_2041,N_24611,N_24571);
or UO_2042 (O_2042,N_24627,N_24522);
nand UO_2043 (O_2043,N_24673,N_24710);
nand UO_2044 (O_2044,N_24874,N_24876);
or UO_2045 (O_2045,N_24793,N_24944);
nand UO_2046 (O_2046,N_24843,N_24718);
and UO_2047 (O_2047,N_24871,N_24921);
nor UO_2048 (O_2048,N_24732,N_24911);
and UO_2049 (O_2049,N_24576,N_24518);
nor UO_2050 (O_2050,N_24645,N_24886);
xnor UO_2051 (O_2051,N_24881,N_24676);
and UO_2052 (O_2052,N_24918,N_24944);
or UO_2053 (O_2053,N_24806,N_24940);
nand UO_2054 (O_2054,N_24904,N_24960);
nand UO_2055 (O_2055,N_24853,N_24583);
xor UO_2056 (O_2056,N_24847,N_24906);
and UO_2057 (O_2057,N_24514,N_24525);
and UO_2058 (O_2058,N_24600,N_24846);
or UO_2059 (O_2059,N_24825,N_24855);
or UO_2060 (O_2060,N_24935,N_24843);
nand UO_2061 (O_2061,N_24930,N_24611);
or UO_2062 (O_2062,N_24590,N_24607);
nor UO_2063 (O_2063,N_24772,N_24535);
xor UO_2064 (O_2064,N_24658,N_24690);
xnor UO_2065 (O_2065,N_24668,N_24878);
nand UO_2066 (O_2066,N_24917,N_24855);
xor UO_2067 (O_2067,N_24726,N_24548);
nand UO_2068 (O_2068,N_24617,N_24693);
or UO_2069 (O_2069,N_24675,N_24759);
nor UO_2070 (O_2070,N_24941,N_24955);
nand UO_2071 (O_2071,N_24715,N_24942);
nand UO_2072 (O_2072,N_24517,N_24811);
nor UO_2073 (O_2073,N_24729,N_24993);
and UO_2074 (O_2074,N_24527,N_24666);
and UO_2075 (O_2075,N_24531,N_24721);
xnor UO_2076 (O_2076,N_24715,N_24564);
nor UO_2077 (O_2077,N_24835,N_24790);
nor UO_2078 (O_2078,N_24943,N_24920);
nor UO_2079 (O_2079,N_24562,N_24634);
xor UO_2080 (O_2080,N_24683,N_24758);
nor UO_2081 (O_2081,N_24840,N_24822);
nor UO_2082 (O_2082,N_24657,N_24700);
xnor UO_2083 (O_2083,N_24582,N_24934);
xor UO_2084 (O_2084,N_24748,N_24975);
and UO_2085 (O_2085,N_24586,N_24592);
or UO_2086 (O_2086,N_24659,N_24780);
nand UO_2087 (O_2087,N_24706,N_24605);
nor UO_2088 (O_2088,N_24827,N_24630);
xnor UO_2089 (O_2089,N_24949,N_24808);
nand UO_2090 (O_2090,N_24920,N_24834);
or UO_2091 (O_2091,N_24650,N_24813);
nand UO_2092 (O_2092,N_24904,N_24842);
nand UO_2093 (O_2093,N_24970,N_24918);
nand UO_2094 (O_2094,N_24582,N_24601);
nor UO_2095 (O_2095,N_24632,N_24763);
and UO_2096 (O_2096,N_24911,N_24852);
nand UO_2097 (O_2097,N_24785,N_24745);
xnor UO_2098 (O_2098,N_24812,N_24542);
and UO_2099 (O_2099,N_24663,N_24812);
or UO_2100 (O_2100,N_24984,N_24892);
xnor UO_2101 (O_2101,N_24588,N_24536);
and UO_2102 (O_2102,N_24898,N_24772);
xor UO_2103 (O_2103,N_24709,N_24518);
nand UO_2104 (O_2104,N_24752,N_24981);
or UO_2105 (O_2105,N_24994,N_24934);
or UO_2106 (O_2106,N_24727,N_24946);
or UO_2107 (O_2107,N_24751,N_24518);
nand UO_2108 (O_2108,N_24938,N_24995);
nor UO_2109 (O_2109,N_24508,N_24919);
nor UO_2110 (O_2110,N_24664,N_24583);
or UO_2111 (O_2111,N_24770,N_24842);
and UO_2112 (O_2112,N_24998,N_24595);
and UO_2113 (O_2113,N_24821,N_24610);
xor UO_2114 (O_2114,N_24684,N_24960);
and UO_2115 (O_2115,N_24849,N_24548);
nand UO_2116 (O_2116,N_24684,N_24778);
xnor UO_2117 (O_2117,N_24779,N_24734);
xnor UO_2118 (O_2118,N_24698,N_24677);
nor UO_2119 (O_2119,N_24837,N_24982);
or UO_2120 (O_2120,N_24520,N_24541);
nand UO_2121 (O_2121,N_24872,N_24555);
and UO_2122 (O_2122,N_24894,N_24826);
and UO_2123 (O_2123,N_24844,N_24733);
nor UO_2124 (O_2124,N_24828,N_24930);
or UO_2125 (O_2125,N_24985,N_24989);
nor UO_2126 (O_2126,N_24811,N_24816);
xnor UO_2127 (O_2127,N_24676,N_24678);
nand UO_2128 (O_2128,N_24775,N_24530);
and UO_2129 (O_2129,N_24796,N_24762);
xor UO_2130 (O_2130,N_24680,N_24544);
nor UO_2131 (O_2131,N_24568,N_24690);
and UO_2132 (O_2132,N_24513,N_24582);
or UO_2133 (O_2133,N_24546,N_24910);
xnor UO_2134 (O_2134,N_24989,N_24527);
and UO_2135 (O_2135,N_24511,N_24689);
and UO_2136 (O_2136,N_24763,N_24578);
and UO_2137 (O_2137,N_24808,N_24769);
or UO_2138 (O_2138,N_24684,N_24907);
xor UO_2139 (O_2139,N_24642,N_24546);
nor UO_2140 (O_2140,N_24907,N_24665);
xor UO_2141 (O_2141,N_24863,N_24805);
or UO_2142 (O_2142,N_24627,N_24730);
xnor UO_2143 (O_2143,N_24661,N_24630);
nand UO_2144 (O_2144,N_24976,N_24849);
nor UO_2145 (O_2145,N_24528,N_24947);
and UO_2146 (O_2146,N_24508,N_24815);
and UO_2147 (O_2147,N_24662,N_24771);
xor UO_2148 (O_2148,N_24776,N_24987);
xor UO_2149 (O_2149,N_24822,N_24885);
nor UO_2150 (O_2150,N_24916,N_24733);
xor UO_2151 (O_2151,N_24814,N_24794);
nor UO_2152 (O_2152,N_24701,N_24852);
or UO_2153 (O_2153,N_24763,N_24841);
or UO_2154 (O_2154,N_24929,N_24890);
xnor UO_2155 (O_2155,N_24944,N_24920);
nor UO_2156 (O_2156,N_24844,N_24755);
nor UO_2157 (O_2157,N_24952,N_24616);
or UO_2158 (O_2158,N_24805,N_24605);
and UO_2159 (O_2159,N_24626,N_24646);
xor UO_2160 (O_2160,N_24860,N_24873);
nor UO_2161 (O_2161,N_24959,N_24672);
nand UO_2162 (O_2162,N_24982,N_24943);
nand UO_2163 (O_2163,N_24979,N_24669);
nand UO_2164 (O_2164,N_24519,N_24887);
xor UO_2165 (O_2165,N_24911,N_24514);
xor UO_2166 (O_2166,N_24901,N_24857);
xor UO_2167 (O_2167,N_24647,N_24783);
nand UO_2168 (O_2168,N_24509,N_24629);
and UO_2169 (O_2169,N_24633,N_24854);
xnor UO_2170 (O_2170,N_24526,N_24728);
nand UO_2171 (O_2171,N_24769,N_24751);
or UO_2172 (O_2172,N_24553,N_24550);
xor UO_2173 (O_2173,N_24972,N_24882);
nor UO_2174 (O_2174,N_24956,N_24694);
nand UO_2175 (O_2175,N_24742,N_24831);
or UO_2176 (O_2176,N_24504,N_24797);
xnor UO_2177 (O_2177,N_24993,N_24513);
nand UO_2178 (O_2178,N_24963,N_24819);
or UO_2179 (O_2179,N_24827,N_24595);
and UO_2180 (O_2180,N_24985,N_24814);
or UO_2181 (O_2181,N_24908,N_24877);
nand UO_2182 (O_2182,N_24968,N_24920);
nand UO_2183 (O_2183,N_24632,N_24819);
and UO_2184 (O_2184,N_24631,N_24591);
or UO_2185 (O_2185,N_24773,N_24635);
xor UO_2186 (O_2186,N_24808,N_24531);
and UO_2187 (O_2187,N_24948,N_24794);
nand UO_2188 (O_2188,N_24952,N_24998);
xor UO_2189 (O_2189,N_24534,N_24661);
xnor UO_2190 (O_2190,N_24776,N_24745);
xnor UO_2191 (O_2191,N_24756,N_24886);
nand UO_2192 (O_2192,N_24613,N_24706);
xor UO_2193 (O_2193,N_24541,N_24627);
nor UO_2194 (O_2194,N_24796,N_24535);
nor UO_2195 (O_2195,N_24997,N_24656);
or UO_2196 (O_2196,N_24529,N_24773);
and UO_2197 (O_2197,N_24578,N_24592);
nor UO_2198 (O_2198,N_24829,N_24838);
and UO_2199 (O_2199,N_24510,N_24774);
nand UO_2200 (O_2200,N_24866,N_24769);
or UO_2201 (O_2201,N_24828,N_24689);
xnor UO_2202 (O_2202,N_24962,N_24734);
nand UO_2203 (O_2203,N_24605,N_24767);
and UO_2204 (O_2204,N_24955,N_24812);
and UO_2205 (O_2205,N_24510,N_24892);
and UO_2206 (O_2206,N_24533,N_24923);
nand UO_2207 (O_2207,N_24578,N_24779);
nand UO_2208 (O_2208,N_24563,N_24996);
and UO_2209 (O_2209,N_24932,N_24939);
nand UO_2210 (O_2210,N_24999,N_24503);
xnor UO_2211 (O_2211,N_24834,N_24694);
nor UO_2212 (O_2212,N_24600,N_24841);
nor UO_2213 (O_2213,N_24549,N_24700);
xnor UO_2214 (O_2214,N_24629,N_24962);
or UO_2215 (O_2215,N_24892,N_24917);
nor UO_2216 (O_2216,N_24668,N_24613);
xnor UO_2217 (O_2217,N_24913,N_24882);
or UO_2218 (O_2218,N_24746,N_24714);
or UO_2219 (O_2219,N_24890,N_24898);
nor UO_2220 (O_2220,N_24794,N_24740);
xnor UO_2221 (O_2221,N_24817,N_24597);
or UO_2222 (O_2222,N_24690,N_24659);
xor UO_2223 (O_2223,N_24913,N_24946);
or UO_2224 (O_2224,N_24860,N_24650);
xor UO_2225 (O_2225,N_24691,N_24729);
nand UO_2226 (O_2226,N_24541,N_24662);
xor UO_2227 (O_2227,N_24516,N_24930);
and UO_2228 (O_2228,N_24938,N_24965);
and UO_2229 (O_2229,N_24665,N_24791);
and UO_2230 (O_2230,N_24605,N_24815);
or UO_2231 (O_2231,N_24640,N_24718);
xor UO_2232 (O_2232,N_24775,N_24682);
and UO_2233 (O_2233,N_24998,N_24910);
and UO_2234 (O_2234,N_24702,N_24556);
nand UO_2235 (O_2235,N_24916,N_24933);
nand UO_2236 (O_2236,N_24792,N_24770);
nor UO_2237 (O_2237,N_24584,N_24610);
xnor UO_2238 (O_2238,N_24679,N_24586);
xor UO_2239 (O_2239,N_24788,N_24642);
xor UO_2240 (O_2240,N_24721,N_24890);
or UO_2241 (O_2241,N_24768,N_24819);
xnor UO_2242 (O_2242,N_24931,N_24922);
nor UO_2243 (O_2243,N_24634,N_24825);
nand UO_2244 (O_2244,N_24732,N_24807);
nand UO_2245 (O_2245,N_24637,N_24971);
or UO_2246 (O_2246,N_24945,N_24712);
nor UO_2247 (O_2247,N_24505,N_24535);
or UO_2248 (O_2248,N_24799,N_24596);
xor UO_2249 (O_2249,N_24514,N_24792);
and UO_2250 (O_2250,N_24711,N_24975);
nand UO_2251 (O_2251,N_24600,N_24602);
or UO_2252 (O_2252,N_24581,N_24840);
xnor UO_2253 (O_2253,N_24541,N_24749);
nand UO_2254 (O_2254,N_24706,N_24674);
nand UO_2255 (O_2255,N_24857,N_24972);
and UO_2256 (O_2256,N_24530,N_24960);
or UO_2257 (O_2257,N_24923,N_24871);
nand UO_2258 (O_2258,N_24948,N_24578);
xnor UO_2259 (O_2259,N_24593,N_24695);
and UO_2260 (O_2260,N_24518,N_24936);
nor UO_2261 (O_2261,N_24919,N_24515);
nor UO_2262 (O_2262,N_24780,N_24772);
nand UO_2263 (O_2263,N_24868,N_24802);
nand UO_2264 (O_2264,N_24563,N_24540);
or UO_2265 (O_2265,N_24600,N_24833);
or UO_2266 (O_2266,N_24548,N_24835);
or UO_2267 (O_2267,N_24565,N_24500);
nor UO_2268 (O_2268,N_24866,N_24536);
and UO_2269 (O_2269,N_24878,N_24817);
or UO_2270 (O_2270,N_24776,N_24575);
nand UO_2271 (O_2271,N_24920,N_24730);
xor UO_2272 (O_2272,N_24960,N_24689);
or UO_2273 (O_2273,N_24606,N_24942);
or UO_2274 (O_2274,N_24909,N_24678);
nor UO_2275 (O_2275,N_24919,N_24570);
nor UO_2276 (O_2276,N_24770,N_24963);
xor UO_2277 (O_2277,N_24978,N_24753);
nand UO_2278 (O_2278,N_24914,N_24801);
and UO_2279 (O_2279,N_24909,N_24978);
or UO_2280 (O_2280,N_24800,N_24629);
nor UO_2281 (O_2281,N_24992,N_24607);
nor UO_2282 (O_2282,N_24547,N_24928);
nor UO_2283 (O_2283,N_24926,N_24764);
xnor UO_2284 (O_2284,N_24953,N_24706);
xor UO_2285 (O_2285,N_24529,N_24509);
nor UO_2286 (O_2286,N_24833,N_24558);
and UO_2287 (O_2287,N_24632,N_24731);
nor UO_2288 (O_2288,N_24501,N_24620);
or UO_2289 (O_2289,N_24783,N_24741);
nand UO_2290 (O_2290,N_24547,N_24633);
nor UO_2291 (O_2291,N_24750,N_24506);
or UO_2292 (O_2292,N_24833,N_24840);
or UO_2293 (O_2293,N_24896,N_24662);
and UO_2294 (O_2294,N_24641,N_24696);
nand UO_2295 (O_2295,N_24869,N_24752);
nand UO_2296 (O_2296,N_24920,N_24504);
nand UO_2297 (O_2297,N_24802,N_24835);
nor UO_2298 (O_2298,N_24901,N_24769);
or UO_2299 (O_2299,N_24945,N_24998);
and UO_2300 (O_2300,N_24885,N_24681);
or UO_2301 (O_2301,N_24506,N_24780);
or UO_2302 (O_2302,N_24989,N_24895);
and UO_2303 (O_2303,N_24534,N_24933);
xnor UO_2304 (O_2304,N_24524,N_24935);
or UO_2305 (O_2305,N_24623,N_24995);
xor UO_2306 (O_2306,N_24920,N_24506);
xor UO_2307 (O_2307,N_24539,N_24681);
xnor UO_2308 (O_2308,N_24939,N_24613);
and UO_2309 (O_2309,N_24723,N_24570);
nor UO_2310 (O_2310,N_24774,N_24803);
xnor UO_2311 (O_2311,N_24952,N_24628);
nor UO_2312 (O_2312,N_24734,N_24915);
and UO_2313 (O_2313,N_24584,N_24922);
xnor UO_2314 (O_2314,N_24704,N_24875);
xnor UO_2315 (O_2315,N_24898,N_24864);
nor UO_2316 (O_2316,N_24606,N_24768);
xor UO_2317 (O_2317,N_24685,N_24830);
nand UO_2318 (O_2318,N_24734,N_24684);
nor UO_2319 (O_2319,N_24831,N_24828);
xnor UO_2320 (O_2320,N_24710,N_24544);
nand UO_2321 (O_2321,N_24687,N_24649);
or UO_2322 (O_2322,N_24891,N_24601);
nor UO_2323 (O_2323,N_24718,N_24655);
and UO_2324 (O_2324,N_24696,N_24938);
or UO_2325 (O_2325,N_24808,N_24713);
xor UO_2326 (O_2326,N_24681,N_24984);
nor UO_2327 (O_2327,N_24568,N_24500);
nor UO_2328 (O_2328,N_24853,N_24528);
or UO_2329 (O_2329,N_24558,N_24840);
nor UO_2330 (O_2330,N_24681,N_24850);
or UO_2331 (O_2331,N_24978,N_24712);
nand UO_2332 (O_2332,N_24809,N_24657);
nand UO_2333 (O_2333,N_24854,N_24869);
or UO_2334 (O_2334,N_24590,N_24593);
nor UO_2335 (O_2335,N_24974,N_24560);
xnor UO_2336 (O_2336,N_24540,N_24714);
nand UO_2337 (O_2337,N_24812,N_24581);
or UO_2338 (O_2338,N_24740,N_24576);
nand UO_2339 (O_2339,N_24731,N_24944);
xnor UO_2340 (O_2340,N_24746,N_24567);
nand UO_2341 (O_2341,N_24899,N_24971);
nor UO_2342 (O_2342,N_24723,N_24743);
xnor UO_2343 (O_2343,N_24970,N_24558);
xor UO_2344 (O_2344,N_24860,N_24716);
or UO_2345 (O_2345,N_24651,N_24963);
nor UO_2346 (O_2346,N_24609,N_24741);
nor UO_2347 (O_2347,N_24631,N_24873);
nor UO_2348 (O_2348,N_24568,N_24630);
or UO_2349 (O_2349,N_24649,N_24750);
nand UO_2350 (O_2350,N_24708,N_24537);
nor UO_2351 (O_2351,N_24708,N_24930);
nand UO_2352 (O_2352,N_24825,N_24780);
and UO_2353 (O_2353,N_24769,N_24599);
or UO_2354 (O_2354,N_24821,N_24996);
nor UO_2355 (O_2355,N_24844,N_24667);
nand UO_2356 (O_2356,N_24845,N_24685);
and UO_2357 (O_2357,N_24555,N_24505);
or UO_2358 (O_2358,N_24705,N_24937);
xnor UO_2359 (O_2359,N_24708,N_24830);
and UO_2360 (O_2360,N_24561,N_24927);
or UO_2361 (O_2361,N_24744,N_24960);
or UO_2362 (O_2362,N_24577,N_24894);
or UO_2363 (O_2363,N_24591,N_24944);
nand UO_2364 (O_2364,N_24602,N_24685);
and UO_2365 (O_2365,N_24917,N_24745);
or UO_2366 (O_2366,N_24653,N_24939);
nor UO_2367 (O_2367,N_24858,N_24910);
xor UO_2368 (O_2368,N_24678,N_24698);
and UO_2369 (O_2369,N_24520,N_24550);
or UO_2370 (O_2370,N_24812,N_24661);
or UO_2371 (O_2371,N_24596,N_24611);
or UO_2372 (O_2372,N_24902,N_24825);
nand UO_2373 (O_2373,N_24508,N_24511);
or UO_2374 (O_2374,N_24735,N_24737);
and UO_2375 (O_2375,N_24746,N_24956);
or UO_2376 (O_2376,N_24551,N_24915);
and UO_2377 (O_2377,N_24939,N_24515);
xor UO_2378 (O_2378,N_24659,N_24916);
nor UO_2379 (O_2379,N_24656,N_24952);
or UO_2380 (O_2380,N_24654,N_24870);
nor UO_2381 (O_2381,N_24550,N_24557);
and UO_2382 (O_2382,N_24856,N_24704);
or UO_2383 (O_2383,N_24968,N_24870);
nand UO_2384 (O_2384,N_24834,N_24604);
nand UO_2385 (O_2385,N_24913,N_24731);
xor UO_2386 (O_2386,N_24718,N_24537);
nand UO_2387 (O_2387,N_24619,N_24674);
and UO_2388 (O_2388,N_24520,N_24514);
and UO_2389 (O_2389,N_24742,N_24982);
xnor UO_2390 (O_2390,N_24608,N_24568);
and UO_2391 (O_2391,N_24570,N_24534);
nand UO_2392 (O_2392,N_24532,N_24528);
xor UO_2393 (O_2393,N_24562,N_24512);
nand UO_2394 (O_2394,N_24847,N_24587);
and UO_2395 (O_2395,N_24824,N_24567);
nand UO_2396 (O_2396,N_24983,N_24665);
and UO_2397 (O_2397,N_24790,N_24991);
nor UO_2398 (O_2398,N_24874,N_24965);
xnor UO_2399 (O_2399,N_24573,N_24900);
and UO_2400 (O_2400,N_24523,N_24773);
nor UO_2401 (O_2401,N_24834,N_24955);
nand UO_2402 (O_2402,N_24756,N_24892);
nor UO_2403 (O_2403,N_24794,N_24962);
xor UO_2404 (O_2404,N_24601,N_24846);
nor UO_2405 (O_2405,N_24732,N_24695);
nor UO_2406 (O_2406,N_24907,N_24834);
xnor UO_2407 (O_2407,N_24839,N_24926);
nand UO_2408 (O_2408,N_24969,N_24675);
nand UO_2409 (O_2409,N_24735,N_24881);
nor UO_2410 (O_2410,N_24682,N_24632);
or UO_2411 (O_2411,N_24712,N_24792);
and UO_2412 (O_2412,N_24632,N_24768);
xor UO_2413 (O_2413,N_24717,N_24810);
nand UO_2414 (O_2414,N_24898,N_24715);
xnor UO_2415 (O_2415,N_24573,N_24816);
or UO_2416 (O_2416,N_24630,N_24629);
nand UO_2417 (O_2417,N_24989,N_24671);
xnor UO_2418 (O_2418,N_24619,N_24967);
nand UO_2419 (O_2419,N_24899,N_24867);
nand UO_2420 (O_2420,N_24711,N_24704);
nand UO_2421 (O_2421,N_24546,N_24835);
nor UO_2422 (O_2422,N_24823,N_24585);
or UO_2423 (O_2423,N_24594,N_24971);
nor UO_2424 (O_2424,N_24527,N_24741);
nor UO_2425 (O_2425,N_24547,N_24923);
and UO_2426 (O_2426,N_24808,N_24576);
nor UO_2427 (O_2427,N_24898,N_24989);
nand UO_2428 (O_2428,N_24695,N_24882);
xnor UO_2429 (O_2429,N_24660,N_24747);
and UO_2430 (O_2430,N_24938,N_24827);
xnor UO_2431 (O_2431,N_24783,N_24655);
xor UO_2432 (O_2432,N_24648,N_24767);
xor UO_2433 (O_2433,N_24769,N_24950);
xor UO_2434 (O_2434,N_24503,N_24884);
and UO_2435 (O_2435,N_24834,N_24997);
nand UO_2436 (O_2436,N_24752,N_24763);
nand UO_2437 (O_2437,N_24579,N_24663);
and UO_2438 (O_2438,N_24882,N_24751);
xnor UO_2439 (O_2439,N_24775,N_24909);
xnor UO_2440 (O_2440,N_24559,N_24724);
nor UO_2441 (O_2441,N_24742,N_24997);
or UO_2442 (O_2442,N_24658,N_24872);
nor UO_2443 (O_2443,N_24623,N_24630);
or UO_2444 (O_2444,N_24780,N_24925);
and UO_2445 (O_2445,N_24703,N_24756);
nand UO_2446 (O_2446,N_24959,N_24971);
and UO_2447 (O_2447,N_24682,N_24651);
and UO_2448 (O_2448,N_24785,N_24750);
and UO_2449 (O_2449,N_24784,N_24725);
nand UO_2450 (O_2450,N_24913,N_24784);
xnor UO_2451 (O_2451,N_24627,N_24595);
nand UO_2452 (O_2452,N_24862,N_24586);
or UO_2453 (O_2453,N_24595,N_24626);
nor UO_2454 (O_2454,N_24990,N_24712);
nor UO_2455 (O_2455,N_24711,N_24625);
nor UO_2456 (O_2456,N_24740,N_24997);
xor UO_2457 (O_2457,N_24508,N_24887);
nand UO_2458 (O_2458,N_24550,N_24518);
nor UO_2459 (O_2459,N_24524,N_24620);
nand UO_2460 (O_2460,N_24675,N_24647);
nand UO_2461 (O_2461,N_24564,N_24515);
nand UO_2462 (O_2462,N_24515,N_24596);
nor UO_2463 (O_2463,N_24994,N_24619);
xor UO_2464 (O_2464,N_24509,N_24899);
xnor UO_2465 (O_2465,N_24519,N_24625);
or UO_2466 (O_2466,N_24992,N_24939);
nand UO_2467 (O_2467,N_24748,N_24525);
nor UO_2468 (O_2468,N_24703,N_24986);
xor UO_2469 (O_2469,N_24605,N_24905);
and UO_2470 (O_2470,N_24970,N_24620);
nand UO_2471 (O_2471,N_24506,N_24670);
xnor UO_2472 (O_2472,N_24724,N_24950);
or UO_2473 (O_2473,N_24757,N_24586);
nor UO_2474 (O_2474,N_24723,N_24880);
and UO_2475 (O_2475,N_24627,N_24829);
and UO_2476 (O_2476,N_24518,N_24893);
or UO_2477 (O_2477,N_24991,N_24760);
and UO_2478 (O_2478,N_24799,N_24702);
nand UO_2479 (O_2479,N_24527,N_24565);
xnor UO_2480 (O_2480,N_24567,N_24801);
xnor UO_2481 (O_2481,N_24714,N_24625);
and UO_2482 (O_2482,N_24601,N_24826);
nand UO_2483 (O_2483,N_24870,N_24920);
nand UO_2484 (O_2484,N_24843,N_24807);
nor UO_2485 (O_2485,N_24827,N_24881);
xnor UO_2486 (O_2486,N_24982,N_24974);
nor UO_2487 (O_2487,N_24597,N_24675);
and UO_2488 (O_2488,N_24865,N_24903);
xnor UO_2489 (O_2489,N_24551,N_24652);
or UO_2490 (O_2490,N_24633,N_24817);
and UO_2491 (O_2491,N_24781,N_24622);
nor UO_2492 (O_2492,N_24674,N_24668);
and UO_2493 (O_2493,N_24613,N_24828);
xor UO_2494 (O_2494,N_24734,N_24686);
nor UO_2495 (O_2495,N_24650,N_24671);
nor UO_2496 (O_2496,N_24575,N_24950);
or UO_2497 (O_2497,N_24621,N_24663);
nand UO_2498 (O_2498,N_24834,N_24755);
nand UO_2499 (O_2499,N_24937,N_24592);
nor UO_2500 (O_2500,N_24816,N_24817);
nor UO_2501 (O_2501,N_24937,N_24972);
nor UO_2502 (O_2502,N_24561,N_24948);
nor UO_2503 (O_2503,N_24690,N_24600);
nand UO_2504 (O_2504,N_24941,N_24749);
nor UO_2505 (O_2505,N_24578,N_24599);
nand UO_2506 (O_2506,N_24960,N_24898);
xnor UO_2507 (O_2507,N_24908,N_24680);
xor UO_2508 (O_2508,N_24797,N_24855);
and UO_2509 (O_2509,N_24898,N_24906);
and UO_2510 (O_2510,N_24664,N_24685);
or UO_2511 (O_2511,N_24658,N_24918);
and UO_2512 (O_2512,N_24659,N_24615);
and UO_2513 (O_2513,N_24837,N_24521);
or UO_2514 (O_2514,N_24837,N_24768);
xnor UO_2515 (O_2515,N_24869,N_24562);
xor UO_2516 (O_2516,N_24741,N_24830);
and UO_2517 (O_2517,N_24834,N_24697);
or UO_2518 (O_2518,N_24811,N_24676);
nor UO_2519 (O_2519,N_24672,N_24827);
nor UO_2520 (O_2520,N_24843,N_24947);
and UO_2521 (O_2521,N_24970,N_24560);
xnor UO_2522 (O_2522,N_24940,N_24880);
nand UO_2523 (O_2523,N_24521,N_24984);
nor UO_2524 (O_2524,N_24933,N_24829);
nor UO_2525 (O_2525,N_24687,N_24758);
nand UO_2526 (O_2526,N_24911,N_24941);
nand UO_2527 (O_2527,N_24764,N_24799);
or UO_2528 (O_2528,N_24763,N_24892);
and UO_2529 (O_2529,N_24669,N_24997);
nor UO_2530 (O_2530,N_24764,N_24585);
nand UO_2531 (O_2531,N_24740,N_24502);
nor UO_2532 (O_2532,N_24829,N_24789);
and UO_2533 (O_2533,N_24767,N_24762);
and UO_2534 (O_2534,N_24872,N_24620);
nand UO_2535 (O_2535,N_24602,N_24541);
xor UO_2536 (O_2536,N_24756,N_24778);
nor UO_2537 (O_2537,N_24507,N_24613);
xnor UO_2538 (O_2538,N_24987,N_24840);
and UO_2539 (O_2539,N_24905,N_24682);
or UO_2540 (O_2540,N_24597,N_24883);
nor UO_2541 (O_2541,N_24791,N_24840);
nand UO_2542 (O_2542,N_24734,N_24976);
nand UO_2543 (O_2543,N_24541,N_24639);
xor UO_2544 (O_2544,N_24808,N_24661);
nor UO_2545 (O_2545,N_24951,N_24672);
and UO_2546 (O_2546,N_24622,N_24513);
nor UO_2547 (O_2547,N_24696,N_24688);
nand UO_2548 (O_2548,N_24989,N_24611);
nand UO_2549 (O_2549,N_24675,N_24936);
nand UO_2550 (O_2550,N_24537,N_24929);
nor UO_2551 (O_2551,N_24734,N_24754);
and UO_2552 (O_2552,N_24536,N_24981);
or UO_2553 (O_2553,N_24728,N_24990);
or UO_2554 (O_2554,N_24854,N_24714);
nor UO_2555 (O_2555,N_24981,N_24833);
nand UO_2556 (O_2556,N_24696,N_24535);
nand UO_2557 (O_2557,N_24779,N_24623);
and UO_2558 (O_2558,N_24519,N_24624);
and UO_2559 (O_2559,N_24701,N_24634);
nand UO_2560 (O_2560,N_24689,N_24706);
nor UO_2561 (O_2561,N_24571,N_24781);
nand UO_2562 (O_2562,N_24575,N_24753);
nand UO_2563 (O_2563,N_24734,N_24824);
nand UO_2564 (O_2564,N_24866,N_24927);
nand UO_2565 (O_2565,N_24968,N_24684);
xnor UO_2566 (O_2566,N_24753,N_24643);
and UO_2567 (O_2567,N_24823,N_24622);
nor UO_2568 (O_2568,N_24577,N_24736);
or UO_2569 (O_2569,N_24922,N_24871);
nand UO_2570 (O_2570,N_24881,N_24595);
nor UO_2571 (O_2571,N_24610,N_24727);
nand UO_2572 (O_2572,N_24990,N_24803);
xnor UO_2573 (O_2573,N_24601,N_24777);
nand UO_2574 (O_2574,N_24888,N_24814);
nor UO_2575 (O_2575,N_24722,N_24594);
and UO_2576 (O_2576,N_24503,N_24771);
or UO_2577 (O_2577,N_24872,N_24647);
nand UO_2578 (O_2578,N_24883,N_24574);
nor UO_2579 (O_2579,N_24606,N_24721);
and UO_2580 (O_2580,N_24917,N_24906);
nor UO_2581 (O_2581,N_24986,N_24752);
and UO_2582 (O_2582,N_24571,N_24765);
nor UO_2583 (O_2583,N_24730,N_24548);
nand UO_2584 (O_2584,N_24704,N_24690);
or UO_2585 (O_2585,N_24959,N_24609);
nand UO_2586 (O_2586,N_24717,N_24736);
or UO_2587 (O_2587,N_24833,N_24891);
and UO_2588 (O_2588,N_24587,N_24852);
xnor UO_2589 (O_2589,N_24732,N_24884);
xnor UO_2590 (O_2590,N_24559,N_24818);
nor UO_2591 (O_2591,N_24668,N_24617);
xnor UO_2592 (O_2592,N_24529,N_24528);
or UO_2593 (O_2593,N_24912,N_24535);
xor UO_2594 (O_2594,N_24698,N_24810);
xnor UO_2595 (O_2595,N_24693,N_24981);
nor UO_2596 (O_2596,N_24786,N_24556);
xnor UO_2597 (O_2597,N_24940,N_24849);
xor UO_2598 (O_2598,N_24685,N_24581);
xnor UO_2599 (O_2599,N_24947,N_24808);
or UO_2600 (O_2600,N_24857,N_24956);
nand UO_2601 (O_2601,N_24526,N_24854);
xor UO_2602 (O_2602,N_24998,N_24987);
nor UO_2603 (O_2603,N_24713,N_24625);
or UO_2604 (O_2604,N_24518,N_24802);
nand UO_2605 (O_2605,N_24526,N_24754);
or UO_2606 (O_2606,N_24519,N_24665);
xnor UO_2607 (O_2607,N_24502,N_24940);
and UO_2608 (O_2608,N_24725,N_24756);
nor UO_2609 (O_2609,N_24816,N_24639);
nor UO_2610 (O_2610,N_24745,N_24621);
nor UO_2611 (O_2611,N_24506,N_24795);
xnor UO_2612 (O_2612,N_24976,N_24531);
or UO_2613 (O_2613,N_24653,N_24926);
nor UO_2614 (O_2614,N_24784,N_24510);
and UO_2615 (O_2615,N_24652,N_24568);
nand UO_2616 (O_2616,N_24717,N_24861);
xor UO_2617 (O_2617,N_24668,N_24522);
and UO_2618 (O_2618,N_24632,N_24696);
or UO_2619 (O_2619,N_24830,N_24669);
nor UO_2620 (O_2620,N_24754,N_24609);
and UO_2621 (O_2621,N_24608,N_24650);
and UO_2622 (O_2622,N_24858,N_24611);
nor UO_2623 (O_2623,N_24966,N_24764);
or UO_2624 (O_2624,N_24645,N_24612);
and UO_2625 (O_2625,N_24580,N_24598);
and UO_2626 (O_2626,N_24582,N_24992);
nor UO_2627 (O_2627,N_24937,N_24831);
and UO_2628 (O_2628,N_24756,N_24931);
xnor UO_2629 (O_2629,N_24869,N_24505);
or UO_2630 (O_2630,N_24842,N_24691);
nor UO_2631 (O_2631,N_24675,N_24638);
and UO_2632 (O_2632,N_24558,N_24864);
or UO_2633 (O_2633,N_24945,N_24634);
or UO_2634 (O_2634,N_24820,N_24872);
and UO_2635 (O_2635,N_24936,N_24776);
or UO_2636 (O_2636,N_24716,N_24988);
or UO_2637 (O_2637,N_24717,N_24871);
xnor UO_2638 (O_2638,N_24843,N_24618);
nand UO_2639 (O_2639,N_24995,N_24993);
nor UO_2640 (O_2640,N_24953,N_24978);
nand UO_2641 (O_2641,N_24590,N_24746);
nor UO_2642 (O_2642,N_24937,N_24934);
nand UO_2643 (O_2643,N_24894,N_24586);
nor UO_2644 (O_2644,N_24688,N_24992);
nand UO_2645 (O_2645,N_24820,N_24772);
and UO_2646 (O_2646,N_24691,N_24733);
nor UO_2647 (O_2647,N_24916,N_24653);
and UO_2648 (O_2648,N_24622,N_24549);
and UO_2649 (O_2649,N_24751,N_24850);
and UO_2650 (O_2650,N_24967,N_24615);
or UO_2651 (O_2651,N_24918,N_24888);
nand UO_2652 (O_2652,N_24991,N_24679);
nand UO_2653 (O_2653,N_24802,N_24933);
and UO_2654 (O_2654,N_24891,N_24690);
and UO_2655 (O_2655,N_24925,N_24525);
xnor UO_2656 (O_2656,N_24919,N_24873);
nor UO_2657 (O_2657,N_24698,N_24920);
xnor UO_2658 (O_2658,N_24967,N_24893);
xnor UO_2659 (O_2659,N_24580,N_24527);
and UO_2660 (O_2660,N_24535,N_24963);
or UO_2661 (O_2661,N_24585,N_24607);
or UO_2662 (O_2662,N_24544,N_24928);
nand UO_2663 (O_2663,N_24671,N_24505);
nand UO_2664 (O_2664,N_24672,N_24620);
or UO_2665 (O_2665,N_24770,N_24938);
and UO_2666 (O_2666,N_24698,N_24910);
or UO_2667 (O_2667,N_24785,N_24933);
or UO_2668 (O_2668,N_24880,N_24736);
nand UO_2669 (O_2669,N_24773,N_24706);
nor UO_2670 (O_2670,N_24620,N_24530);
or UO_2671 (O_2671,N_24818,N_24544);
nand UO_2672 (O_2672,N_24643,N_24821);
nand UO_2673 (O_2673,N_24923,N_24818);
nor UO_2674 (O_2674,N_24884,N_24749);
nand UO_2675 (O_2675,N_24877,N_24951);
nand UO_2676 (O_2676,N_24680,N_24945);
and UO_2677 (O_2677,N_24780,N_24960);
nand UO_2678 (O_2678,N_24503,N_24801);
and UO_2679 (O_2679,N_24651,N_24797);
xor UO_2680 (O_2680,N_24866,N_24904);
nand UO_2681 (O_2681,N_24876,N_24771);
xor UO_2682 (O_2682,N_24770,N_24979);
xor UO_2683 (O_2683,N_24758,N_24614);
nor UO_2684 (O_2684,N_24985,N_24808);
xnor UO_2685 (O_2685,N_24591,N_24804);
xnor UO_2686 (O_2686,N_24618,N_24686);
xor UO_2687 (O_2687,N_24564,N_24650);
or UO_2688 (O_2688,N_24530,N_24626);
or UO_2689 (O_2689,N_24512,N_24754);
xnor UO_2690 (O_2690,N_24593,N_24576);
nor UO_2691 (O_2691,N_24677,N_24585);
or UO_2692 (O_2692,N_24974,N_24981);
nand UO_2693 (O_2693,N_24620,N_24894);
xor UO_2694 (O_2694,N_24799,N_24819);
or UO_2695 (O_2695,N_24820,N_24852);
xnor UO_2696 (O_2696,N_24801,N_24729);
xnor UO_2697 (O_2697,N_24584,N_24656);
nand UO_2698 (O_2698,N_24861,N_24918);
and UO_2699 (O_2699,N_24762,N_24732);
and UO_2700 (O_2700,N_24921,N_24592);
or UO_2701 (O_2701,N_24569,N_24851);
nand UO_2702 (O_2702,N_24695,N_24558);
or UO_2703 (O_2703,N_24588,N_24520);
xnor UO_2704 (O_2704,N_24728,N_24875);
nand UO_2705 (O_2705,N_24659,N_24894);
and UO_2706 (O_2706,N_24728,N_24937);
xor UO_2707 (O_2707,N_24697,N_24564);
nor UO_2708 (O_2708,N_24724,N_24748);
and UO_2709 (O_2709,N_24733,N_24571);
or UO_2710 (O_2710,N_24647,N_24861);
or UO_2711 (O_2711,N_24987,N_24961);
and UO_2712 (O_2712,N_24749,N_24853);
nand UO_2713 (O_2713,N_24549,N_24922);
and UO_2714 (O_2714,N_24847,N_24702);
nand UO_2715 (O_2715,N_24905,N_24538);
or UO_2716 (O_2716,N_24763,N_24557);
or UO_2717 (O_2717,N_24845,N_24514);
xnor UO_2718 (O_2718,N_24897,N_24885);
and UO_2719 (O_2719,N_24878,N_24963);
nor UO_2720 (O_2720,N_24649,N_24656);
or UO_2721 (O_2721,N_24576,N_24804);
or UO_2722 (O_2722,N_24787,N_24873);
nand UO_2723 (O_2723,N_24772,N_24802);
xor UO_2724 (O_2724,N_24744,N_24791);
xor UO_2725 (O_2725,N_24572,N_24777);
xnor UO_2726 (O_2726,N_24990,N_24617);
and UO_2727 (O_2727,N_24574,N_24585);
nand UO_2728 (O_2728,N_24624,N_24951);
nand UO_2729 (O_2729,N_24546,N_24676);
or UO_2730 (O_2730,N_24809,N_24798);
nand UO_2731 (O_2731,N_24854,N_24682);
and UO_2732 (O_2732,N_24752,N_24797);
or UO_2733 (O_2733,N_24936,N_24898);
or UO_2734 (O_2734,N_24841,N_24649);
xor UO_2735 (O_2735,N_24705,N_24841);
or UO_2736 (O_2736,N_24855,N_24739);
nor UO_2737 (O_2737,N_24826,N_24597);
or UO_2738 (O_2738,N_24826,N_24621);
xor UO_2739 (O_2739,N_24571,N_24741);
nor UO_2740 (O_2740,N_24562,N_24605);
xor UO_2741 (O_2741,N_24629,N_24684);
xor UO_2742 (O_2742,N_24726,N_24675);
xnor UO_2743 (O_2743,N_24775,N_24573);
nor UO_2744 (O_2744,N_24611,N_24516);
and UO_2745 (O_2745,N_24928,N_24799);
nor UO_2746 (O_2746,N_24516,N_24735);
and UO_2747 (O_2747,N_24778,N_24516);
and UO_2748 (O_2748,N_24843,N_24980);
xnor UO_2749 (O_2749,N_24606,N_24751);
nor UO_2750 (O_2750,N_24938,N_24562);
or UO_2751 (O_2751,N_24545,N_24813);
or UO_2752 (O_2752,N_24852,N_24882);
nor UO_2753 (O_2753,N_24602,N_24655);
or UO_2754 (O_2754,N_24559,N_24843);
nor UO_2755 (O_2755,N_24592,N_24640);
or UO_2756 (O_2756,N_24970,N_24770);
xnor UO_2757 (O_2757,N_24950,N_24879);
xnor UO_2758 (O_2758,N_24670,N_24713);
and UO_2759 (O_2759,N_24707,N_24619);
nor UO_2760 (O_2760,N_24934,N_24573);
xnor UO_2761 (O_2761,N_24753,N_24676);
nand UO_2762 (O_2762,N_24994,N_24902);
or UO_2763 (O_2763,N_24578,N_24608);
and UO_2764 (O_2764,N_24929,N_24809);
nand UO_2765 (O_2765,N_24790,N_24776);
nand UO_2766 (O_2766,N_24630,N_24538);
nor UO_2767 (O_2767,N_24783,N_24632);
nand UO_2768 (O_2768,N_24667,N_24971);
xor UO_2769 (O_2769,N_24843,N_24881);
xor UO_2770 (O_2770,N_24964,N_24509);
nor UO_2771 (O_2771,N_24600,N_24796);
nand UO_2772 (O_2772,N_24729,N_24752);
or UO_2773 (O_2773,N_24725,N_24524);
nand UO_2774 (O_2774,N_24587,N_24962);
nor UO_2775 (O_2775,N_24868,N_24680);
nand UO_2776 (O_2776,N_24691,N_24955);
and UO_2777 (O_2777,N_24655,N_24542);
or UO_2778 (O_2778,N_24558,N_24516);
and UO_2779 (O_2779,N_24990,N_24706);
and UO_2780 (O_2780,N_24968,N_24983);
nand UO_2781 (O_2781,N_24666,N_24915);
and UO_2782 (O_2782,N_24743,N_24922);
or UO_2783 (O_2783,N_24723,N_24936);
nand UO_2784 (O_2784,N_24609,N_24518);
xor UO_2785 (O_2785,N_24805,N_24802);
nor UO_2786 (O_2786,N_24779,N_24560);
or UO_2787 (O_2787,N_24749,N_24882);
or UO_2788 (O_2788,N_24589,N_24734);
nand UO_2789 (O_2789,N_24632,N_24794);
xnor UO_2790 (O_2790,N_24524,N_24736);
nand UO_2791 (O_2791,N_24641,N_24904);
nand UO_2792 (O_2792,N_24747,N_24540);
and UO_2793 (O_2793,N_24810,N_24866);
xnor UO_2794 (O_2794,N_24509,N_24534);
nand UO_2795 (O_2795,N_24973,N_24933);
and UO_2796 (O_2796,N_24860,N_24768);
xnor UO_2797 (O_2797,N_24596,N_24958);
and UO_2798 (O_2798,N_24638,N_24823);
xnor UO_2799 (O_2799,N_24607,N_24810);
xor UO_2800 (O_2800,N_24813,N_24578);
nor UO_2801 (O_2801,N_24569,N_24574);
and UO_2802 (O_2802,N_24600,N_24818);
xor UO_2803 (O_2803,N_24649,N_24818);
or UO_2804 (O_2804,N_24593,N_24703);
and UO_2805 (O_2805,N_24584,N_24945);
nor UO_2806 (O_2806,N_24545,N_24773);
or UO_2807 (O_2807,N_24996,N_24755);
nand UO_2808 (O_2808,N_24507,N_24623);
nand UO_2809 (O_2809,N_24980,N_24955);
or UO_2810 (O_2810,N_24735,N_24519);
nand UO_2811 (O_2811,N_24541,N_24778);
nand UO_2812 (O_2812,N_24629,N_24996);
nor UO_2813 (O_2813,N_24989,N_24821);
nor UO_2814 (O_2814,N_24647,N_24881);
xor UO_2815 (O_2815,N_24615,N_24890);
nand UO_2816 (O_2816,N_24645,N_24539);
or UO_2817 (O_2817,N_24735,N_24842);
nand UO_2818 (O_2818,N_24820,N_24529);
and UO_2819 (O_2819,N_24570,N_24969);
xnor UO_2820 (O_2820,N_24685,N_24641);
xor UO_2821 (O_2821,N_24710,N_24873);
xor UO_2822 (O_2822,N_24527,N_24632);
nand UO_2823 (O_2823,N_24508,N_24559);
xor UO_2824 (O_2824,N_24785,N_24769);
and UO_2825 (O_2825,N_24618,N_24975);
or UO_2826 (O_2826,N_24976,N_24547);
nand UO_2827 (O_2827,N_24693,N_24553);
and UO_2828 (O_2828,N_24583,N_24667);
nor UO_2829 (O_2829,N_24918,N_24950);
nand UO_2830 (O_2830,N_24804,N_24639);
and UO_2831 (O_2831,N_24814,N_24946);
or UO_2832 (O_2832,N_24529,N_24920);
and UO_2833 (O_2833,N_24883,N_24784);
or UO_2834 (O_2834,N_24792,N_24861);
xnor UO_2835 (O_2835,N_24546,N_24787);
nand UO_2836 (O_2836,N_24710,N_24693);
nand UO_2837 (O_2837,N_24936,N_24538);
nand UO_2838 (O_2838,N_24620,N_24602);
nor UO_2839 (O_2839,N_24771,N_24761);
xor UO_2840 (O_2840,N_24646,N_24645);
and UO_2841 (O_2841,N_24541,N_24523);
or UO_2842 (O_2842,N_24765,N_24732);
and UO_2843 (O_2843,N_24511,N_24994);
xnor UO_2844 (O_2844,N_24523,N_24920);
and UO_2845 (O_2845,N_24925,N_24639);
nand UO_2846 (O_2846,N_24528,N_24710);
or UO_2847 (O_2847,N_24582,N_24634);
or UO_2848 (O_2848,N_24788,N_24925);
or UO_2849 (O_2849,N_24587,N_24856);
xnor UO_2850 (O_2850,N_24600,N_24605);
nor UO_2851 (O_2851,N_24685,N_24960);
or UO_2852 (O_2852,N_24508,N_24920);
nand UO_2853 (O_2853,N_24606,N_24765);
nor UO_2854 (O_2854,N_24913,N_24867);
nor UO_2855 (O_2855,N_24677,N_24793);
xnor UO_2856 (O_2856,N_24909,N_24617);
and UO_2857 (O_2857,N_24969,N_24906);
xnor UO_2858 (O_2858,N_24957,N_24648);
or UO_2859 (O_2859,N_24576,N_24653);
and UO_2860 (O_2860,N_24794,N_24761);
xor UO_2861 (O_2861,N_24626,N_24765);
nor UO_2862 (O_2862,N_24766,N_24597);
and UO_2863 (O_2863,N_24693,N_24966);
nor UO_2864 (O_2864,N_24892,N_24762);
or UO_2865 (O_2865,N_24862,N_24527);
and UO_2866 (O_2866,N_24857,N_24838);
xor UO_2867 (O_2867,N_24505,N_24701);
xnor UO_2868 (O_2868,N_24963,N_24780);
or UO_2869 (O_2869,N_24766,N_24961);
and UO_2870 (O_2870,N_24867,N_24912);
nand UO_2871 (O_2871,N_24624,N_24617);
or UO_2872 (O_2872,N_24780,N_24531);
and UO_2873 (O_2873,N_24881,N_24667);
and UO_2874 (O_2874,N_24798,N_24625);
and UO_2875 (O_2875,N_24671,N_24775);
xor UO_2876 (O_2876,N_24984,N_24771);
xnor UO_2877 (O_2877,N_24617,N_24632);
or UO_2878 (O_2878,N_24922,N_24607);
xnor UO_2879 (O_2879,N_24904,N_24814);
nand UO_2880 (O_2880,N_24722,N_24786);
or UO_2881 (O_2881,N_24630,N_24654);
nand UO_2882 (O_2882,N_24782,N_24540);
or UO_2883 (O_2883,N_24838,N_24718);
nor UO_2884 (O_2884,N_24941,N_24552);
xor UO_2885 (O_2885,N_24906,N_24967);
nor UO_2886 (O_2886,N_24905,N_24868);
or UO_2887 (O_2887,N_24848,N_24681);
nand UO_2888 (O_2888,N_24889,N_24915);
and UO_2889 (O_2889,N_24810,N_24517);
nor UO_2890 (O_2890,N_24758,N_24610);
or UO_2891 (O_2891,N_24605,N_24768);
xor UO_2892 (O_2892,N_24656,N_24702);
nand UO_2893 (O_2893,N_24891,N_24510);
xor UO_2894 (O_2894,N_24653,N_24942);
or UO_2895 (O_2895,N_24634,N_24681);
and UO_2896 (O_2896,N_24746,N_24884);
xnor UO_2897 (O_2897,N_24551,N_24529);
nor UO_2898 (O_2898,N_24887,N_24831);
nand UO_2899 (O_2899,N_24672,N_24578);
nand UO_2900 (O_2900,N_24953,N_24755);
or UO_2901 (O_2901,N_24788,N_24913);
nor UO_2902 (O_2902,N_24729,N_24935);
xnor UO_2903 (O_2903,N_24609,N_24818);
or UO_2904 (O_2904,N_24536,N_24712);
or UO_2905 (O_2905,N_24634,N_24740);
xnor UO_2906 (O_2906,N_24728,N_24624);
xor UO_2907 (O_2907,N_24688,N_24769);
nor UO_2908 (O_2908,N_24961,N_24603);
and UO_2909 (O_2909,N_24870,N_24957);
or UO_2910 (O_2910,N_24894,N_24768);
or UO_2911 (O_2911,N_24520,N_24605);
nor UO_2912 (O_2912,N_24968,N_24594);
nand UO_2913 (O_2913,N_24772,N_24618);
nor UO_2914 (O_2914,N_24927,N_24792);
nand UO_2915 (O_2915,N_24549,N_24794);
and UO_2916 (O_2916,N_24908,N_24679);
nand UO_2917 (O_2917,N_24766,N_24968);
and UO_2918 (O_2918,N_24999,N_24950);
and UO_2919 (O_2919,N_24965,N_24826);
nand UO_2920 (O_2920,N_24510,N_24692);
and UO_2921 (O_2921,N_24924,N_24789);
or UO_2922 (O_2922,N_24571,N_24631);
nand UO_2923 (O_2923,N_24988,N_24567);
xor UO_2924 (O_2924,N_24650,N_24660);
nand UO_2925 (O_2925,N_24844,N_24676);
xor UO_2926 (O_2926,N_24934,N_24875);
or UO_2927 (O_2927,N_24836,N_24830);
or UO_2928 (O_2928,N_24892,N_24870);
nor UO_2929 (O_2929,N_24648,N_24887);
xnor UO_2930 (O_2930,N_24724,N_24844);
and UO_2931 (O_2931,N_24625,N_24912);
xnor UO_2932 (O_2932,N_24540,N_24904);
xor UO_2933 (O_2933,N_24655,N_24779);
xnor UO_2934 (O_2934,N_24950,N_24899);
nor UO_2935 (O_2935,N_24851,N_24684);
xnor UO_2936 (O_2936,N_24940,N_24805);
xnor UO_2937 (O_2937,N_24748,N_24501);
xnor UO_2938 (O_2938,N_24590,N_24845);
or UO_2939 (O_2939,N_24545,N_24938);
and UO_2940 (O_2940,N_24848,N_24995);
xor UO_2941 (O_2941,N_24945,N_24917);
and UO_2942 (O_2942,N_24651,N_24709);
nand UO_2943 (O_2943,N_24649,N_24601);
nor UO_2944 (O_2944,N_24796,N_24970);
xor UO_2945 (O_2945,N_24641,N_24951);
xor UO_2946 (O_2946,N_24738,N_24761);
nand UO_2947 (O_2947,N_24557,N_24842);
nor UO_2948 (O_2948,N_24976,N_24733);
xnor UO_2949 (O_2949,N_24657,N_24767);
nor UO_2950 (O_2950,N_24769,N_24746);
or UO_2951 (O_2951,N_24912,N_24549);
nand UO_2952 (O_2952,N_24891,N_24817);
nand UO_2953 (O_2953,N_24700,N_24976);
xnor UO_2954 (O_2954,N_24915,N_24729);
nor UO_2955 (O_2955,N_24503,N_24928);
or UO_2956 (O_2956,N_24605,N_24724);
or UO_2957 (O_2957,N_24999,N_24780);
nand UO_2958 (O_2958,N_24570,N_24852);
and UO_2959 (O_2959,N_24858,N_24988);
xnor UO_2960 (O_2960,N_24521,N_24533);
nand UO_2961 (O_2961,N_24534,N_24896);
nand UO_2962 (O_2962,N_24518,N_24659);
or UO_2963 (O_2963,N_24522,N_24665);
nand UO_2964 (O_2964,N_24932,N_24503);
xnor UO_2965 (O_2965,N_24974,N_24510);
xnor UO_2966 (O_2966,N_24650,N_24990);
nand UO_2967 (O_2967,N_24850,N_24714);
and UO_2968 (O_2968,N_24969,N_24561);
nand UO_2969 (O_2969,N_24977,N_24842);
nand UO_2970 (O_2970,N_24805,N_24571);
or UO_2971 (O_2971,N_24974,N_24916);
xor UO_2972 (O_2972,N_24645,N_24998);
and UO_2973 (O_2973,N_24964,N_24923);
nor UO_2974 (O_2974,N_24563,N_24678);
xor UO_2975 (O_2975,N_24608,N_24961);
nor UO_2976 (O_2976,N_24738,N_24802);
or UO_2977 (O_2977,N_24948,N_24565);
nand UO_2978 (O_2978,N_24587,N_24891);
nor UO_2979 (O_2979,N_24614,N_24718);
and UO_2980 (O_2980,N_24552,N_24733);
nand UO_2981 (O_2981,N_24589,N_24569);
and UO_2982 (O_2982,N_24940,N_24993);
or UO_2983 (O_2983,N_24787,N_24926);
or UO_2984 (O_2984,N_24613,N_24885);
nor UO_2985 (O_2985,N_24936,N_24669);
and UO_2986 (O_2986,N_24892,N_24548);
nor UO_2987 (O_2987,N_24872,N_24797);
nand UO_2988 (O_2988,N_24823,N_24615);
or UO_2989 (O_2989,N_24774,N_24776);
and UO_2990 (O_2990,N_24591,N_24755);
and UO_2991 (O_2991,N_24843,N_24884);
or UO_2992 (O_2992,N_24779,N_24504);
nand UO_2993 (O_2993,N_24779,N_24853);
nand UO_2994 (O_2994,N_24947,N_24839);
nor UO_2995 (O_2995,N_24986,N_24993);
xor UO_2996 (O_2996,N_24740,N_24735);
nor UO_2997 (O_2997,N_24945,N_24709);
nand UO_2998 (O_2998,N_24864,N_24815);
nor UO_2999 (O_2999,N_24987,N_24551);
endmodule