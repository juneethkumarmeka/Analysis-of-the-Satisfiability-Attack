module basic_1500_15000_2000_5_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_1205,In_1475);
and U1 (N_1,In_834,In_326);
nand U2 (N_2,In_1221,In_229);
or U3 (N_3,In_235,In_1290);
or U4 (N_4,In_1279,In_664);
nor U5 (N_5,In_1206,In_1336);
nand U6 (N_6,In_1485,In_468);
nor U7 (N_7,In_1078,In_946);
or U8 (N_8,In_634,In_106);
and U9 (N_9,In_1249,In_1276);
and U10 (N_10,In_923,In_1006);
nor U11 (N_11,In_67,In_453);
nand U12 (N_12,In_1032,In_310);
or U13 (N_13,In_1478,In_733);
nand U14 (N_14,In_1218,In_254);
nor U15 (N_15,In_147,In_1196);
nand U16 (N_16,In_1202,In_550);
and U17 (N_17,In_433,In_915);
and U18 (N_18,In_971,In_1297);
or U19 (N_19,In_793,In_1161);
nor U20 (N_20,In_162,In_367);
or U21 (N_21,In_1317,In_1013);
and U22 (N_22,In_920,In_69);
or U23 (N_23,In_997,In_1396);
nand U24 (N_24,In_1285,In_1399);
or U25 (N_25,In_1381,In_341);
and U26 (N_26,In_14,In_752);
nand U27 (N_27,In_861,In_301);
or U28 (N_28,In_1146,In_1234);
and U29 (N_29,In_218,In_1088);
nor U30 (N_30,In_1471,In_762);
and U31 (N_31,In_1470,In_142);
or U32 (N_32,In_1347,In_182);
and U33 (N_33,In_383,In_1484);
or U34 (N_34,In_709,In_245);
nor U35 (N_35,In_394,In_812);
nor U36 (N_36,In_425,In_1282);
and U37 (N_37,In_1229,In_533);
nand U38 (N_38,In_968,In_1151);
or U39 (N_39,In_1014,In_952);
or U40 (N_40,In_52,In_74);
nor U41 (N_41,In_735,In_561);
and U42 (N_42,In_1355,In_1492);
nand U43 (N_43,In_272,In_62);
nor U44 (N_44,In_1265,In_872);
nand U45 (N_45,In_1203,In_189);
nand U46 (N_46,In_1188,In_58);
and U47 (N_47,In_841,In_919);
and U48 (N_48,In_642,In_204);
nand U49 (N_49,In_1000,In_798);
nand U50 (N_50,In_1315,In_80);
nand U51 (N_51,In_1043,In_721);
or U52 (N_52,In_930,In_379);
nor U53 (N_53,In_472,In_977);
nor U54 (N_54,In_519,In_1476);
and U55 (N_55,In_1159,In_710);
or U56 (N_56,In_1487,In_656);
and U57 (N_57,In_1149,In_888);
nor U58 (N_58,In_854,In_222);
nand U59 (N_59,In_848,In_403);
nand U60 (N_60,In_575,In_1152);
or U61 (N_61,In_465,In_178);
nor U62 (N_62,In_342,In_452);
and U63 (N_63,In_1209,In_393);
nand U64 (N_64,In_785,In_494);
nand U65 (N_65,In_1216,In_1294);
nand U66 (N_66,In_92,In_156);
or U67 (N_67,In_1403,In_270);
nor U68 (N_68,In_1250,In_37);
nor U69 (N_69,In_1037,In_138);
nand U70 (N_70,In_258,In_764);
and U71 (N_71,In_715,In_934);
nor U72 (N_72,In_381,In_784);
or U73 (N_73,In_51,In_1359);
and U74 (N_74,In_911,In_741);
and U75 (N_75,In_696,In_417);
nand U76 (N_76,In_716,In_605);
nor U77 (N_77,In_761,In_1240);
nor U78 (N_78,In_257,In_1246);
nor U79 (N_79,In_1133,In_464);
nor U80 (N_80,In_719,In_545);
or U81 (N_81,In_1155,In_451);
and U82 (N_82,In_1314,In_1486);
nand U83 (N_83,In_25,In_455);
nand U84 (N_84,In_1305,In_1357);
nor U85 (N_85,In_317,In_253);
and U86 (N_86,In_294,In_1447);
and U87 (N_87,In_1177,In_240);
or U88 (N_88,In_826,In_1056);
nand U89 (N_89,In_1431,In_763);
nor U90 (N_90,In_1456,In_401);
and U91 (N_91,In_1130,In_4);
xor U92 (N_92,In_905,In_1496);
or U93 (N_93,In_811,In_431);
nor U94 (N_94,In_284,In_543);
xnor U95 (N_95,In_1346,In_970);
and U96 (N_96,In_770,In_694);
or U97 (N_97,In_511,In_1147);
or U98 (N_98,In_1313,In_623);
and U99 (N_99,In_316,In_781);
and U100 (N_100,In_374,In_1068);
or U101 (N_101,In_833,In_410);
nor U102 (N_102,In_1343,In_951);
nand U103 (N_103,In_866,In_1049);
and U104 (N_104,In_1330,In_1375);
nand U105 (N_105,In_172,In_287);
and U106 (N_106,In_969,In_89);
nor U107 (N_107,In_46,In_73);
nand U108 (N_108,In_1195,In_980);
nand U109 (N_109,In_1121,In_1075);
and U110 (N_110,In_690,In_1325);
nand U111 (N_111,In_1423,In_1009);
and U112 (N_112,In_632,In_279);
or U113 (N_113,In_356,In_1488);
nor U114 (N_114,In_699,In_1170);
and U115 (N_115,In_1036,In_517);
or U116 (N_116,In_1318,In_382);
or U117 (N_117,In_1277,In_746);
xor U118 (N_118,In_1004,In_330);
and U119 (N_119,In_1235,In_129);
nand U120 (N_120,In_527,In_1142);
nor U121 (N_121,In_672,In_155);
and U122 (N_122,In_927,In_70);
or U123 (N_123,In_1232,In_547);
nand U124 (N_124,In_1081,In_1425);
or U125 (N_125,In_714,In_559);
and U126 (N_126,In_113,In_742);
nor U127 (N_127,In_313,In_684);
or U128 (N_128,In_975,In_909);
and U129 (N_129,In_31,In_1050);
or U130 (N_130,In_1062,In_288);
nor U131 (N_131,In_568,In_148);
nand U132 (N_132,In_1067,In_108);
or U133 (N_133,In_194,In_344);
nand U134 (N_134,In_759,In_502);
nor U135 (N_135,In_1319,In_844);
and U136 (N_136,In_1460,In_282);
or U137 (N_137,In_1380,In_136);
nor U138 (N_138,In_1176,In_1289);
and U139 (N_139,In_577,In_1472);
and U140 (N_140,In_482,In_1128);
and U141 (N_141,In_555,In_1204);
nand U142 (N_142,In_829,In_835);
or U143 (N_143,In_889,In_1045);
and U144 (N_144,In_1286,In_467);
nand U145 (N_145,In_593,In_99);
and U146 (N_146,In_260,In_495);
and U147 (N_147,In_179,In_1126);
nor U148 (N_148,In_1157,In_730);
and U149 (N_149,In_389,In_591);
nor U150 (N_150,In_1089,In_693);
or U151 (N_151,In_335,In_169);
and U152 (N_152,In_269,In_738);
nand U153 (N_153,In_558,In_857);
nand U154 (N_154,In_1163,In_756);
or U155 (N_155,In_560,In_987);
nor U156 (N_156,In_1057,In_203);
nor U157 (N_157,In_1140,In_1348);
nand U158 (N_158,In_1407,In_687);
nor U159 (N_159,In_497,In_685);
and U160 (N_160,In_666,In_243);
and U161 (N_161,In_1405,In_1100);
or U162 (N_162,In_375,In_63);
or U163 (N_163,In_510,In_1451);
and U164 (N_164,In_447,In_1054);
or U165 (N_165,In_94,In_1442);
xnor U166 (N_166,In_1253,In_101);
or U167 (N_167,In_925,In_123);
or U168 (N_168,In_406,In_163);
nor U169 (N_169,In_366,In_562);
or U170 (N_170,In_928,In_1386);
or U171 (N_171,In_816,In_1382);
or U172 (N_172,In_1239,In_348);
nor U173 (N_173,In_1263,In_552);
or U174 (N_174,In_1086,In_191);
and U175 (N_175,In_574,In_496);
nand U176 (N_176,In_1046,In_883);
and U177 (N_177,In_77,In_336);
nor U178 (N_178,In_1410,In_1421);
or U179 (N_179,In_1371,In_137);
or U180 (N_180,In_818,In_322);
and U181 (N_181,In_1010,In_1022);
nor U182 (N_182,In_328,In_198);
nand U183 (N_183,In_630,In_902);
nand U184 (N_184,In_1292,In_777);
or U185 (N_185,In_1303,In_786);
and U186 (N_186,In_1287,In_318);
or U187 (N_187,In_734,In_1061);
nor U188 (N_188,In_520,In_722);
nor U189 (N_189,In_851,In_1441);
or U190 (N_190,In_1102,In_1463);
nand U191 (N_191,In_910,In_731);
nand U192 (N_192,In_414,In_1224);
or U193 (N_193,In_19,In_567);
or U194 (N_194,In_1225,In_250);
nor U195 (N_195,In_964,In_512);
nor U196 (N_196,In_195,In_643);
and U197 (N_197,In_343,In_661);
nand U198 (N_198,In_15,In_723);
nand U199 (N_199,In_1400,In_388);
or U200 (N_200,In_659,In_1233);
and U201 (N_201,In_1422,In_184);
nand U202 (N_202,In_416,In_1115);
and U203 (N_203,In_481,In_614);
nand U204 (N_204,In_1254,In_1272);
or U205 (N_205,In_1110,In_200);
nand U206 (N_206,In_1454,In_1450);
nor U207 (N_207,In_1160,In_864);
nor U208 (N_208,In_1490,In_627);
nand U209 (N_209,In_1,In_529);
and U210 (N_210,In_350,In_1383);
and U211 (N_211,In_1109,In_845);
or U212 (N_212,In_650,In_128);
xor U213 (N_213,In_81,In_580);
nor U214 (N_214,In_1077,In_912);
nor U215 (N_215,In_1241,In_219);
or U216 (N_216,In_807,In_1270);
nand U217 (N_217,In_1212,In_90);
nor U218 (N_218,In_1499,In_779);
xor U219 (N_219,In_1015,In_1034);
nand U220 (N_220,In_1338,In_1440);
or U221 (N_221,In_105,In_958);
nand U222 (N_222,In_1200,In_1419);
nor U223 (N_223,In_1256,In_732);
and U224 (N_224,In_3,In_991);
nor U225 (N_225,In_594,In_206);
or U226 (N_226,In_739,In_936);
or U227 (N_227,In_1173,In_535);
nand U228 (N_228,In_399,In_1238);
nor U229 (N_229,In_941,In_385);
nor U230 (N_230,In_61,In_525);
and U231 (N_231,In_293,In_1041);
nor U232 (N_232,In_747,In_667);
or U233 (N_233,In_718,In_648);
or U234 (N_234,In_285,In_1458);
nor U235 (N_235,In_146,In_397);
nor U236 (N_236,In_996,In_620);
and U237 (N_237,In_469,In_1047);
or U238 (N_238,In_47,In_507);
nor U239 (N_239,In_1184,In_1274);
nand U240 (N_240,In_470,In_261);
and U241 (N_241,In_390,In_295);
or U242 (N_242,In_349,In_745);
and U243 (N_243,In_879,In_929);
nor U244 (N_244,In_772,In_68);
nor U245 (N_245,In_153,In_1326);
nand U246 (N_246,In_1342,In_300);
nor U247 (N_247,In_1174,In_333);
nor U248 (N_248,In_20,In_1153);
nor U249 (N_249,In_441,In_609);
nor U250 (N_250,In_140,In_1372);
and U251 (N_251,In_1025,In_100);
or U252 (N_252,In_1117,In_1031);
and U253 (N_253,In_949,In_1101);
nor U254 (N_254,In_59,In_773);
nand U255 (N_255,In_956,In_1213);
nand U256 (N_256,In_9,In_1210);
and U257 (N_257,In_542,In_10);
or U258 (N_258,In_1302,In_1363);
or U259 (N_259,In_411,In_449);
xor U260 (N_260,In_1390,In_116);
nand U261 (N_261,In_1103,In_654);
nand U262 (N_262,In_681,In_1427);
and U263 (N_263,In_112,In_249);
xor U264 (N_264,In_271,In_751);
nand U265 (N_265,In_66,In_1122);
or U266 (N_266,In_386,In_1226);
and U267 (N_267,In_278,In_1281);
nand U268 (N_268,In_556,In_1311);
nor U269 (N_269,In_1245,In_1280);
nand U270 (N_270,In_810,In_602);
nand U271 (N_271,In_1262,In_1242);
nand U272 (N_272,In_1299,In_358);
nor U273 (N_273,In_233,In_1323);
or U274 (N_274,In_624,In_637);
or U275 (N_275,In_1464,In_982);
nand U276 (N_276,In_57,In_782);
nor U277 (N_277,In_150,In_276);
nor U278 (N_278,In_1446,In_508);
nand U279 (N_279,In_315,In_228);
or U280 (N_280,In_1392,In_308);
nand U281 (N_281,In_445,In_1247);
nor U282 (N_282,In_776,In_774);
and U283 (N_283,In_1208,In_428);
xnor U284 (N_284,In_862,In_639);
or U285 (N_285,In_769,In_1179);
nand U286 (N_286,In_478,In_488);
or U287 (N_287,In_215,In_1308);
and U288 (N_288,In_387,In_1469);
and U289 (N_289,In_139,In_359);
xnor U290 (N_290,In_850,In_1296);
nand U291 (N_291,In_1401,In_154);
or U292 (N_292,In_1011,In_1304);
nor U293 (N_293,In_815,In_16);
or U294 (N_294,In_590,In_573);
or U295 (N_295,In_521,In_332);
and U296 (N_296,In_799,In_345);
or U297 (N_297,In_1430,In_585);
nand U298 (N_298,In_280,In_1020);
or U299 (N_299,In_413,In_462);
and U300 (N_300,In_407,In_1364);
and U301 (N_301,In_571,In_208);
nand U302 (N_302,In_1001,In_24);
nor U303 (N_303,In_838,In_1243);
nor U304 (N_304,In_1432,In_499);
or U305 (N_305,In_456,In_1275);
nor U306 (N_306,In_917,In_1428);
and U307 (N_307,In_853,In_901);
nand U308 (N_308,In_794,In_1096);
or U309 (N_309,In_130,In_423);
and U310 (N_310,In_466,In_539);
nand U311 (N_311,In_171,In_931);
nor U312 (N_312,In_662,In_117);
and U313 (N_313,In_658,In_576);
or U314 (N_314,In_115,In_1017);
or U315 (N_315,In_1331,In_1104);
nand U316 (N_316,In_126,In_242);
and U317 (N_317,In_489,In_87);
xnor U318 (N_318,In_1337,In_1350);
nor U319 (N_319,In_691,In_230);
nor U320 (N_320,In_298,In_788);
and U321 (N_321,In_223,In_541);
nand U322 (N_322,In_205,In_633);
nand U323 (N_323,In_484,In_444);
nand U324 (N_324,In_1076,In_876);
or U325 (N_325,In_60,In_1433);
and U326 (N_326,In_706,In_708);
or U327 (N_327,In_974,In_1353);
nand U328 (N_328,In_678,In_405);
or U329 (N_329,In_806,In_972);
nor U330 (N_330,In_1026,In_524);
and U331 (N_331,In_1093,In_789);
or U332 (N_332,In_363,In_1426);
or U333 (N_333,In_791,In_1066);
and U334 (N_334,In_1307,In_64);
or U335 (N_335,In_177,In_1029);
or U336 (N_336,In_28,In_1402);
nand U337 (N_337,In_954,In_553);
nand U338 (N_338,In_907,In_419);
nand U339 (N_339,In_1316,In_424);
xnor U340 (N_340,In_1333,In_754);
nand U341 (N_341,In_569,In_1288);
or U342 (N_342,In_1394,In_1420);
and U343 (N_343,In_647,In_1493);
nand U344 (N_344,In_868,In_852);
nor U345 (N_345,In_299,In_1108);
and U346 (N_346,In_1236,In_1082);
or U347 (N_347,In_645,In_107);
or U348 (N_348,In_141,In_697);
or U349 (N_349,In_688,In_1283);
nor U350 (N_350,In_582,In_961);
nor U351 (N_351,In_805,In_1462);
and U352 (N_352,In_225,In_291);
nand U353 (N_353,In_477,In_175);
nand U354 (N_354,In_832,In_668);
or U355 (N_355,In_583,In_304);
or U356 (N_356,In_32,In_947);
or U357 (N_357,In_1231,In_604);
nor U358 (N_358,In_1064,In_669);
and U359 (N_359,In_420,In_534);
nand U360 (N_360,In_161,In_408);
nor U361 (N_361,In_190,In_686);
or U362 (N_362,In_78,In_263);
and U363 (N_363,In_705,In_933);
and U364 (N_364,In_29,In_8);
nor U365 (N_365,In_1003,In_893);
and U366 (N_366,In_683,In_1291);
nor U367 (N_367,In_1434,In_1328);
nor U368 (N_368,In_995,In_1495);
or U369 (N_369,In_167,In_768);
nor U370 (N_370,In_531,In_1158);
nor U371 (N_371,In_1145,In_102);
and U372 (N_372,In_1370,In_783);
and U373 (N_373,In_563,In_606);
nor U374 (N_374,In_505,In_702);
nand U375 (N_375,In_196,In_720);
nor U376 (N_376,In_7,In_860);
and U377 (N_377,In_960,In_646);
or U378 (N_378,In_890,In_611);
nor U379 (N_379,In_1335,In_174);
nand U380 (N_380,In_682,In_274);
nor U381 (N_381,In_1220,In_625);
nand U382 (N_382,In_474,In_290);
and U383 (N_383,In_579,In_698);
nand U384 (N_384,In_922,In_820);
nand U385 (N_385,In_373,In_1028);
or U386 (N_386,In_22,In_460);
and U387 (N_387,In_679,In_1069);
nor U388 (N_388,In_825,In_370);
or U389 (N_389,In_1139,In_760);
and U390 (N_390,In_873,In_790);
nand U391 (N_391,In_652,In_617);
and U392 (N_392,In_765,In_18);
or U393 (N_393,In_940,In_264);
nand U394 (N_394,In_1124,In_1373);
xor U395 (N_395,In_50,In_409);
and U396 (N_396,In_1268,In_849);
or U397 (N_397,In_1119,In_908);
or U398 (N_398,In_950,In_821);
nor U399 (N_399,In_1189,In_942);
nor U400 (N_400,In_612,In_214);
and U401 (N_401,In_1019,In_338);
and U402 (N_402,In_622,In_948);
and U403 (N_403,In_1237,In_1138);
nand U404 (N_404,In_1118,In_1106);
nor U405 (N_405,In_135,In_839);
nor U406 (N_406,In_368,In_145);
nand U407 (N_407,In_267,In_36);
nand U408 (N_408,In_1483,In_30);
and U409 (N_409,In_504,In_376);
and U410 (N_410,In_578,In_689);
nand U411 (N_411,In_1360,In_717);
nand U412 (N_412,In_479,In_1070);
nor U413 (N_413,In_490,In_186);
nor U414 (N_414,In_40,In_748);
nor U415 (N_415,In_628,In_327);
and U416 (N_416,In_439,In_778);
and U417 (N_417,In_1023,In_1468);
or U418 (N_418,In_766,In_395);
and U419 (N_419,In_1387,In_629);
and U420 (N_420,In_79,In_216);
nand U421 (N_421,In_323,In_1084);
nor U422 (N_422,In_1367,In_187);
nand U423 (N_423,In_538,In_896);
or U424 (N_424,In_899,In_989);
nor U425 (N_425,In_1098,In_1024);
nor U426 (N_426,In_98,In_448);
or U427 (N_427,In_1466,In_1259);
nor U428 (N_428,In_631,In_544);
nand U429 (N_429,In_518,In_657);
and U430 (N_430,In_962,In_823);
nand U431 (N_431,In_1339,In_663);
and U432 (N_432,In_985,In_953);
and U433 (N_433,In_1379,In_796);
nand U434 (N_434,In_516,In_158);
and U435 (N_435,In_422,In_1060);
or U436 (N_436,In_75,In_1168);
and U437 (N_437,In_471,In_227);
or U438 (N_438,In_1085,In_2);
and U439 (N_439,In_289,In_34);
and U440 (N_440,In_586,In_320);
or U441 (N_441,In_1191,In_1480);
or U442 (N_442,In_601,In_724);
nand U443 (N_443,In_744,In_476);
or U444 (N_444,In_592,In_1199);
nor U445 (N_445,In_45,In_1306);
xnor U446 (N_446,In_443,In_251);
and U447 (N_447,In_755,In_1412);
nor U448 (N_448,In_843,In_607);
and U449 (N_449,In_900,In_640);
xnor U450 (N_450,In_1175,In_725);
and U451 (N_451,In_1351,In_378);
nand U452 (N_452,In_252,In_675);
and U453 (N_453,In_1154,In_1007);
and U454 (N_454,In_1278,In_392);
or U455 (N_455,In_1356,In_226);
nor U456 (N_456,In_132,In_38);
nand U457 (N_457,In_380,In_729);
and U458 (N_458,In_677,In_878);
nor U459 (N_459,In_938,In_1376);
nand U460 (N_460,In_1352,In_1123);
nor U461 (N_461,In_509,In_551);
and U462 (N_462,In_1477,In_450);
nand U463 (N_463,In_871,In_118);
or U464 (N_464,In_181,In_528);
and U465 (N_465,In_1435,In_339);
or U466 (N_466,In_916,In_1457);
or U467 (N_467,In_673,In_597);
or U468 (N_468,In_49,In_1120);
or U469 (N_469,In_711,In_319);
and U470 (N_470,In_88,In_43);
nand U471 (N_471,In_1181,In_207);
or U472 (N_472,In_565,In_603);
nor U473 (N_473,In_877,In_372);
nor U474 (N_474,In_1071,In_454);
and U475 (N_475,In_302,In_211);
or U476 (N_476,In_334,In_231);
nand U477 (N_477,In_1354,In_1398);
or U478 (N_478,In_831,In_114);
nand U479 (N_479,In_149,In_491);
or U480 (N_480,In_822,In_159);
or U481 (N_481,In_72,In_166);
or U482 (N_482,In_740,In_939);
xnor U483 (N_483,In_522,In_351);
and U484 (N_484,In_473,In_6);
and U485 (N_485,In_268,In_1332);
or U486 (N_486,In_17,In_1300);
or U487 (N_487,In_1345,In_1193);
and U488 (N_488,In_42,In_638);
nand U489 (N_489,In_296,In_506);
nor U490 (N_490,In_1094,In_286);
and U491 (N_491,In_458,In_712);
nor U492 (N_492,In_858,In_1374);
and U493 (N_493,In_170,In_1039);
or U494 (N_494,In_546,In_1125);
nand U495 (N_495,In_93,In_1295);
or U496 (N_496,In_0,In_800);
or U497 (N_497,In_1207,In_1385);
and U498 (N_498,In_665,In_993);
and U499 (N_499,In_157,In_750);
and U500 (N_500,In_1406,In_589);
or U501 (N_501,In_122,In_1150);
and U502 (N_502,In_737,In_1180);
and U503 (N_503,In_1388,In_446);
or U504 (N_504,In_91,In_236);
or U505 (N_505,In_1107,In_1111);
nand U506 (N_506,In_875,In_259);
nor U507 (N_507,In_1309,In_1413);
or U508 (N_508,In_1248,In_202);
nor U509 (N_509,In_986,In_151);
or U510 (N_510,In_224,In_311);
nand U511 (N_511,In_641,In_1453);
nor U512 (N_512,In_340,In_213);
and U513 (N_513,In_897,In_1257);
nor U514 (N_514,In_808,In_780);
nor U515 (N_515,In_1048,In_427);
or U516 (N_516,In_1051,In_1197);
nor U517 (N_517,In_830,In_1198);
or U518 (N_518,In_1143,In_435);
and U519 (N_519,In_1172,In_514);
nor U520 (N_520,In_121,In_353);
or U521 (N_521,In_983,In_160);
and U522 (N_522,In_35,In_217);
nand U523 (N_523,In_1448,In_847);
and U524 (N_524,In_1134,In_165);
and U525 (N_525,In_1087,In_885);
or U526 (N_526,In_842,In_1378);
nor U527 (N_527,In_840,In_1312);
nand U528 (N_528,In_434,In_1228);
and U529 (N_529,In_1095,In_1252);
and U530 (N_530,In_440,In_266);
nor U531 (N_531,In_999,In_674);
and U532 (N_532,In_131,In_212);
nand U533 (N_533,In_247,In_354);
nor U534 (N_534,In_1194,In_1341);
or U535 (N_535,In_421,In_1227);
or U536 (N_536,In_957,In_127);
or U537 (N_537,In_1391,In_273);
or U538 (N_538,In_1171,In_1053);
and U539 (N_539,In_307,In_1298);
or U540 (N_540,In_391,In_1473);
nand U541 (N_541,In_526,In_881);
or U542 (N_542,In_437,In_736);
nor U543 (N_543,In_44,In_981);
or U544 (N_544,In_1042,In_39);
and U545 (N_545,In_41,In_703);
or U546 (N_546,In_973,In_314);
xor U547 (N_547,In_581,In_1395);
or U548 (N_548,In_1349,In_192);
nor U549 (N_549,In_1044,In_97);
or U550 (N_550,In_500,In_1255);
or U551 (N_551,In_880,In_670);
nor U552 (N_552,In_1183,In_1135);
and U553 (N_553,In_1362,In_554);
nand U554 (N_554,In_649,In_5);
or U555 (N_555,In_362,In_1097);
and U556 (N_556,In_1244,In_1452);
or U557 (N_557,In_461,In_1321);
or U558 (N_558,In_83,In_183);
and U559 (N_559,In_707,In_1033);
and U560 (N_560,In_1012,In_635);
and U561 (N_561,In_891,In_1489);
nand U562 (N_562,In_86,In_570);
and U563 (N_563,In_26,In_1058);
nand U564 (N_564,In_1429,In_859);
nor U565 (N_565,In_1008,In_185);
or U566 (N_566,In_817,In_713);
nand U567 (N_567,In_935,In_771);
nor U568 (N_568,In_775,In_1408);
nor U569 (N_569,In_201,In_1494);
nand U570 (N_570,In_809,In_221);
or U571 (N_571,In_232,In_1293);
or U572 (N_572,In_56,In_1165);
nand U573 (N_573,In_1411,In_608);
or U574 (N_574,In_1273,In_95);
nand U575 (N_575,In_855,In_1491);
nand U576 (N_576,In_265,In_487);
or U577 (N_577,In_1127,In_802);
or U578 (N_578,In_325,In_1092);
nand U579 (N_579,In_671,In_867);
or U580 (N_580,In_653,In_119);
or U581 (N_581,In_1059,In_598);
nor U582 (N_582,In_1148,In_1162);
and U583 (N_583,In_990,In_613);
or U584 (N_584,In_870,In_1324);
and U585 (N_585,In_1099,In_1424);
or U586 (N_586,In_588,In_111);
and U587 (N_587,In_152,In_210);
nor U588 (N_588,In_1465,In_1340);
and U589 (N_589,In_1261,In_882);
nand U590 (N_590,In_12,In_1327);
or U591 (N_591,In_238,In_587);
nand U592 (N_592,In_176,In_1393);
or U593 (N_593,In_874,In_1271);
or U594 (N_594,In_1409,In_1404);
and U595 (N_595,In_1040,In_887);
and U596 (N_596,In_1481,In_188);
nand U597 (N_597,In_1397,In_994);
nand U598 (N_598,In_965,In_365);
nand U599 (N_599,In_13,In_1474);
or U600 (N_600,In_863,In_1479);
and U601 (N_601,In_944,In_143);
nor U602 (N_602,In_1005,In_400);
and U603 (N_603,In_54,In_655);
or U604 (N_604,In_926,In_1443);
nand U605 (N_605,In_676,In_1377);
and U606 (N_606,In_1083,In_1251);
and U607 (N_607,In_109,In_932);
and U608 (N_608,In_1439,In_914);
nand U609 (N_609,In_1063,In_1222);
or U610 (N_610,In_549,In_480);
or U611 (N_611,In_1021,In_27);
nor U612 (N_612,In_636,In_1116);
nor U613 (N_613,In_438,In_564);
nand U614 (N_614,In_797,In_96);
nor U615 (N_615,In_836,In_804);
nor U616 (N_616,In_988,In_1201);
or U617 (N_617,In_197,In_803);
and U618 (N_618,In_398,In_801);
and U619 (N_619,In_321,In_1185);
nand U620 (N_620,In_819,In_610);
or U621 (N_621,In_1437,In_728);
and U622 (N_622,In_483,In_513);
nor U623 (N_623,In_1438,In_331);
and U624 (N_624,In_1073,In_1467);
and U625 (N_625,In_199,In_626);
and U626 (N_626,In_415,In_234);
nand U627 (N_627,In_244,In_303);
nand U628 (N_628,In_644,In_246);
and U629 (N_629,In_1112,In_692);
nand U630 (N_630,In_1344,In_937);
and U631 (N_631,In_753,In_795);
xor U632 (N_632,In_1052,In_727);
nand U633 (N_633,In_700,In_680);
and U634 (N_634,In_281,In_898);
and U635 (N_635,In_1266,In_1445);
or U636 (N_636,In_1186,In_21);
nand U637 (N_637,In_1264,In_701);
nor U638 (N_638,In_1090,In_125);
nor U639 (N_639,In_704,In_1365);
or U640 (N_640,In_943,In_1214);
and U641 (N_641,In_306,In_329);
or U642 (N_642,In_1219,In_537);
and U643 (N_643,In_486,In_856);
or U644 (N_644,In_361,In_758);
nand U645 (N_645,In_1091,In_892);
nand U646 (N_646,In_384,In_364);
nor U647 (N_647,In_530,In_103);
nand U648 (N_648,In_1418,In_283);
and U649 (N_649,In_1368,In_337);
nand U650 (N_650,In_110,In_1461);
and U651 (N_651,In_621,In_787);
nand U652 (N_652,In_1436,In_85);
and U653 (N_653,In_48,In_1190);
xor U654 (N_654,In_404,In_1030);
nor U655 (N_655,In_492,In_743);
and U656 (N_656,In_924,In_1074);
nor U657 (N_657,In_992,In_33);
nand U658 (N_658,In_292,In_485);
or U659 (N_659,In_168,In_180);
or U660 (N_660,In_846,In_357);
or U661 (N_661,In_572,In_955);
or U662 (N_662,In_305,In_501);
nand U663 (N_663,In_1384,In_436);
or U664 (N_664,In_1369,In_599);
or U665 (N_665,In_979,In_1215);
or U666 (N_666,In_355,In_824);
nor U667 (N_667,In_475,In_1027);
or U668 (N_668,In_792,In_426);
and U669 (N_669,In_1414,In_498);
xnor U670 (N_670,In_1132,In_523);
and U671 (N_671,In_1284,In_402);
xor U672 (N_672,In_1449,In_651);
or U673 (N_673,In_324,In_55);
nor U674 (N_674,In_757,In_726);
and U675 (N_675,In_828,In_1415);
or U676 (N_676,In_503,In_412);
and U677 (N_677,In_813,In_463);
or U678 (N_678,In_963,In_959);
or U679 (N_679,In_277,In_241);
and U680 (N_680,In_104,In_566);
or U681 (N_681,In_1334,In_600);
or U682 (N_682,In_894,In_584);
or U683 (N_683,In_1156,In_369);
and U684 (N_684,In_945,In_1217);
nand U685 (N_685,In_536,In_618);
nand U686 (N_686,In_84,In_1322);
nor U687 (N_687,In_256,In_442);
and U688 (N_688,In_869,In_1105);
nand U689 (N_689,In_430,In_1182);
nand U690 (N_690,In_1055,In_1310);
nor U691 (N_691,In_71,In_124);
and U692 (N_692,In_23,In_1080);
nand U693 (N_693,In_173,In_429);
nor U694 (N_694,In_275,In_886);
nand U695 (N_695,In_297,In_1301);
and U696 (N_696,In_220,In_1329);
nor U697 (N_697,In_1079,In_616);
nand U698 (N_698,In_193,In_1459);
or U699 (N_699,In_615,In_248);
or U700 (N_700,In_1166,In_1187);
nand U701 (N_701,In_1223,In_1167);
or U702 (N_702,In_540,In_53);
nand U703 (N_703,In_1417,In_1455);
nand U704 (N_704,In_1038,In_1389);
nand U705 (N_705,In_493,In_1269);
or U706 (N_706,In_209,In_903);
nand U707 (N_707,In_11,In_906);
or U708 (N_708,In_749,In_1129);
nor U709 (N_709,In_120,In_978);
nor U710 (N_710,In_884,In_1497);
and U711 (N_711,In_695,In_457);
or U712 (N_712,In_360,In_1416);
nor U713 (N_713,In_837,In_913);
and U714 (N_714,In_827,In_619);
nand U715 (N_715,In_237,In_1230);
nor U716 (N_716,In_1358,In_895);
and U717 (N_717,In_967,In_1211);
nand U718 (N_718,In_1141,In_76);
nand U719 (N_719,In_865,In_921);
or U720 (N_720,In_377,In_1192);
nor U721 (N_721,In_595,In_532);
nor U722 (N_722,In_239,In_1267);
and U723 (N_723,In_1361,In_984);
nand U724 (N_724,In_1260,In_814);
nand U725 (N_725,In_1137,In_1444);
or U726 (N_726,In_1320,In_1114);
nand U727 (N_727,In_1164,In_1144);
nand U728 (N_728,In_396,In_557);
and U729 (N_729,In_347,In_144);
nand U730 (N_730,In_1136,In_1482);
or U731 (N_731,In_515,In_82);
nand U732 (N_732,In_1178,In_432);
or U733 (N_733,In_352,In_1366);
xor U734 (N_734,In_1131,In_1065);
and U735 (N_735,In_976,In_371);
and U736 (N_736,In_596,In_1002);
or U737 (N_737,In_1035,In_1016);
or U738 (N_738,In_1169,In_1258);
nor U739 (N_739,In_164,In_312);
and U740 (N_740,In_660,In_918);
xnor U741 (N_741,In_134,In_133);
and U742 (N_742,In_1018,In_548);
or U743 (N_743,In_418,In_262);
or U744 (N_744,In_255,In_459);
or U745 (N_745,In_65,In_1072);
and U746 (N_746,In_998,In_767);
and U747 (N_747,In_904,In_346);
nand U748 (N_748,In_1113,In_1498);
nor U749 (N_749,In_309,In_966);
and U750 (N_750,In_248,In_229);
and U751 (N_751,In_1393,In_119);
and U752 (N_752,In_1498,In_1479);
or U753 (N_753,In_451,In_453);
nor U754 (N_754,In_1024,In_404);
and U755 (N_755,In_1039,In_507);
nor U756 (N_756,In_371,In_210);
nand U757 (N_757,In_329,In_81);
or U758 (N_758,In_1067,In_134);
and U759 (N_759,In_491,In_1054);
nor U760 (N_760,In_689,In_718);
and U761 (N_761,In_1406,In_708);
or U762 (N_762,In_1457,In_1436);
or U763 (N_763,In_1474,In_539);
nor U764 (N_764,In_897,In_371);
nor U765 (N_765,In_1004,In_1144);
and U766 (N_766,In_1016,In_1024);
nand U767 (N_767,In_438,In_580);
nor U768 (N_768,In_293,In_989);
and U769 (N_769,In_176,In_375);
and U770 (N_770,In_614,In_134);
and U771 (N_771,In_189,In_624);
nor U772 (N_772,In_788,In_123);
nand U773 (N_773,In_655,In_188);
or U774 (N_774,In_456,In_1117);
nand U775 (N_775,In_819,In_1199);
or U776 (N_776,In_1128,In_1131);
and U777 (N_777,In_1133,In_946);
and U778 (N_778,In_217,In_572);
or U779 (N_779,In_1163,In_1478);
or U780 (N_780,In_675,In_834);
and U781 (N_781,In_181,In_1274);
nand U782 (N_782,In_886,In_1438);
nor U783 (N_783,In_1460,In_548);
nand U784 (N_784,In_1271,In_1120);
nor U785 (N_785,In_260,In_1451);
nor U786 (N_786,In_1107,In_1461);
nand U787 (N_787,In_1325,In_651);
nand U788 (N_788,In_38,In_296);
and U789 (N_789,In_1310,In_623);
or U790 (N_790,In_654,In_893);
or U791 (N_791,In_1198,In_533);
and U792 (N_792,In_644,In_678);
nand U793 (N_793,In_1445,In_163);
nor U794 (N_794,In_1349,In_468);
nand U795 (N_795,In_489,In_783);
nand U796 (N_796,In_1123,In_334);
and U797 (N_797,In_1400,In_898);
nand U798 (N_798,In_981,In_912);
or U799 (N_799,In_45,In_932);
or U800 (N_800,In_1085,In_120);
nor U801 (N_801,In_871,In_579);
or U802 (N_802,In_726,In_650);
or U803 (N_803,In_693,In_1267);
and U804 (N_804,In_562,In_849);
nor U805 (N_805,In_355,In_789);
or U806 (N_806,In_261,In_266);
nand U807 (N_807,In_79,In_492);
nand U808 (N_808,In_183,In_857);
or U809 (N_809,In_471,In_1125);
nor U810 (N_810,In_848,In_934);
nand U811 (N_811,In_344,In_765);
nand U812 (N_812,In_717,In_1054);
xnor U813 (N_813,In_376,In_668);
and U814 (N_814,In_276,In_121);
xor U815 (N_815,In_249,In_115);
and U816 (N_816,In_1257,In_295);
nand U817 (N_817,In_1231,In_326);
and U818 (N_818,In_1229,In_1215);
or U819 (N_819,In_345,In_109);
and U820 (N_820,In_1208,In_214);
nor U821 (N_821,In_911,In_238);
or U822 (N_822,In_14,In_462);
nor U823 (N_823,In_1229,In_392);
nor U824 (N_824,In_775,In_404);
nor U825 (N_825,In_616,In_317);
and U826 (N_826,In_427,In_1355);
nand U827 (N_827,In_1318,In_914);
nand U828 (N_828,In_1033,In_396);
nand U829 (N_829,In_583,In_853);
and U830 (N_830,In_804,In_894);
or U831 (N_831,In_885,In_125);
and U832 (N_832,In_1310,In_345);
and U833 (N_833,In_1002,In_916);
or U834 (N_834,In_577,In_167);
nor U835 (N_835,In_419,In_794);
or U836 (N_836,In_234,In_1398);
or U837 (N_837,In_89,In_75);
or U838 (N_838,In_277,In_701);
or U839 (N_839,In_444,In_1276);
nand U840 (N_840,In_34,In_447);
nor U841 (N_841,In_726,In_588);
nor U842 (N_842,In_46,In_1236);
or U843 (N_843,In_1152,In_547);
or U844 (N_844,In_536,In_1106);
or U845 (N_845,In_362,In_126);
nor U846 (N_846,In_684,In_165);
nor U847 (N_847,In_884,In_203);
or U848 (N_848,In_1472,In_286);
and U849 (N_849,In_999,In_460);
xnor U850 (N_850,In_43,In_1234);
and U851 (N_851,In_370,In_366);
and U852 (N_852,In_408,In_385);
and U853 (N_853,In_1067,In_964);
and U854 (N_854,In_682,In_1291);
or U855 (N_855,In_862,In_690);
nor U856 (N_856,In_459,In_972);
or U857 (N_857,In_966,In_357);
and U858 (N_858,In_514,In_483);
and U859 (N_859,In_345,In_965);
and U860 (N_860,In_305,In_1069);
and U861 (N_861,In_1108,In_346);
nand U862 (N_862,In_221,In_461);
xnor U863 (N_863,In_1378,In_871);
or U864 (N_864,In_1419,In_255);
and U865 (N_865,In_526,In_430);
or U866 (N_866,In_512,In_956);
nor U867 (N_867,In_1334,In_327);
nand U868 (N_868,In_1350,In_1298);
nor U869 (N_869,In_137,In_200);
nor U870 (N_870,In_1003,In_1159);
and U871 (N_871,In_287,In_262);
or U872 (N_872,In_1181,In_290);
nand U873 (N_873,In_574,In_1196);
nor U874 (N_874,In_142,In_151);
nand U875 (N_875,In_382,In_201);
nand U876 (N_876,In_846,In_457);
or U877 (N_877,In_1345,In_19);
nor U878 (N_878,In_1209,In_1207);
nand U879 (N_879,In_624,In_336);
and U880 (N_880,In_1297,In_1442);
or U881 (N_881,In_270,In_1027);
and U882 (N_882,In_303,In_352);
or U883 (N_883,In_624,In_948);
nand U884 (N_884,In_370,In_884);
nand U885 (N_885,In_1447,In_38);
or U886 (N_886,In_634,In_1106);
nor U887 (N_887,In_427,In_199);
nor U888 (N_888,In_1399,In_1100);
nor U889 (N_889,In_403,In_1189);
nor U890 (N_890,In_24,In_1398);
and U891 (N_891,In_1321,In_381);
and U892 (N_892,In_843,In_1429);
and U893 (N_893,In_1368,In_1278);
nor U894 (N_894,In_1125,In_11);
nor U895 (N_895,In_968,In_784);
nor U896 (N_896,In_923,In_1238);
nand U897 (N_897,In_1425,In_1328);
nor U898 (N_898,In_461,In_1468);
or U899 (N_899,In_1468,In_1121);
nor U900 (N_900,In_794,In_337);
and U901 (N_901,In_1083,In_251);
nor U902 (N_902,In_1041,In_213);
nor U903 (N_903,In_1278,In_189);
nor U904 (N_904,In_1124,In_815);
nor U905 (N_905,In_1436,In_906);
and U906 (N_906,In_620,In_329);
or U907 (N_907,In_671,In_855);
or U908 (N_908,In_1225,In_1094);
and U909 (N_909,In_440,In_963);
and U910 (N_910,In_631,In_1038);
or U911 (N_911,In_958,In_1312);
and U912 (N_912,In_1185,In_495);
xor U913 (N_913,In_1422,In_946);
and U914 (N_914,In_1088,In_1393);
nand U915 (N_915,In_667,In_157);
nand U916 (N_916,In_832,In_897);
and U917 (N_917,In_988,In_83);
nor U918 (N_918,In_891,In_781);
or U919 (N_919,In_34,In_82);
nand U920 (N_920,In_885,In_1178);
nor U921 (N_921,In_1322,In_268);
or U922 (N_922,In_1356,In_229);
nor U923 (N_923,In_733,In_90);
nand U924 (N_924,In_1269,In_209);
nand U925 (N_925,In_990,In_44);
nand U926 (N_926,In_296,In_144);
nand U927 (N_927,In_1378,In_924);
and U928 (N_928,In_1057,In_488);
and U929 (N_929,In_633,In_997);
and U930 (N_930,In_199,In_1221);
and U931 (N_931,In_440,In_1025);
or U932 (N_932,In_1011,In_1284);
nand U933 (N_933,In_809,In_695);
and U934 (N_934,In_1144,In_132);
or U935 (N_935,In_760,In_1248);
or U936 (N_936,In_1415,In_1479);
or U937 (N_937,In_35,In_1014);
nor U938 (N_938,In_836,In_641);
nand U939 (N_939,In_273,In_1189);
and U940 (N_940,In_1394,In_1342);
and U941 (N_941,In_800,In_1097);
and U942 (N_942,In_1317,In_647);
or U943 (N_943,In_1154,In_1374);
nand U944 (N_944,In_1478,In_233);
nand U945 (N_945,In_951,In_228);
nand U946 (N_946,In_1355,In_26);
nor U947 (N_947,In_261,In_433);
xnor U948 (N_948,In_157,In_576);
or U949 (N_949,In_1002,In_89);
nand U950 (N_950,In_999,In_182);
or U951 (N_951,In_1097,In_611);
and U952 (N_952,In_307,In_811);
nand U953 (N_953,In_844,In_885);
nand U954 (N_954,In_564,In_644);
nand U955 (N_955,In_417,In_226);
nor U956 (N_956,In_473,In_509);
nor U957 (N_957,In_854,In_392);
and U958 (N_958,In_46,In_665);
and U959 (N_959,In_120,In_663);
nor U960 (N_960,In_1159,In_420);
or U961 (N_961,In_1097,In_213);
xor U962 (N_962,In_1465,In_1258);
xor U963 (N_963,In_872,In_568);
or U964 (N_964,In_1202,In_1298);
and U965 (N_965,In_1077,In_1142);
nor U966 (N_966,In_1158,In_986);
nor U967 (N_967,In_972,In_138);
or U968 (N_968,In_330,In_277);
or U969 (N_969,In_276,In_892);
xor U970 (N_970,In_1065,In_904);
nor U971 (N_971,In_672,In_477);
nor U972 (N_972,In_335,In_515);
or U973 (N_973,In_1319,In_432);
or U974 (N_974,In_1295,In_75);
or U975 (N_975,In_718,In_986);
or U976 (N_976,In_487,In_993);
nand U977 (N_977,In_628,In_389);
and U978 (N_978,In_638,In_873);
and U979 (N_979,In_289,In_357);
or U980 (N_980,In_932,In_446);
nor U981 (N_981,In_343,In_540);
nand U982 (N_982,In_1135,In_474);
nor U983 (N_983,In_1235,In_958);
nor U984 (N_984,In_785,In_1351);
or U985 (N_985,In_1355,In_288);
nand U986 (N_986,In_1101,In_718);
and U987 (N_987,In_1130,In_1250);
nor U988 (N_988,In_215,In_25);
and U989 (N_989,In_1415,In_57);
or U990 (N_990,In_1101,In_32);
or U991 (N_991,In_678,In_626);
and U992 (N_992,In_1349,In_1261);
and U993 (N_993,In_372,In_1007);
nand U994 (N_994,In_500,In_84);
and U995 (N_995,In_1109,In_493);
nor U996 (N_996,In_716,In_614);
or U997 (N_997,In_388,In_621);
nand U998 (N_998,In_404,In_174);
and U999 (N_999,In_590,In_50);
or U1000 (N_1000,In_1153,In_867);
and U1001 (N_1001,In_173,In_306);
nor U1002 (N_1002,In_1426,In_1469);
nor U1003 (N_1003,In_68,In_271);
nand U1004 (N_1004,In_796,In_1228);
and U1005 (N_1005,In_101,In_531);
nor U1006 (N_1006,In_632,In_400);
nor U1007 (N_1007,In_1117,In_293);
nand U1008 (N_1008,In_311,In_955);
and U1009 (N_1009,In_1355,In_1057);
nor U1010 (N_1010,In_601,In_203);
nand U1011 (N_1011,In_312,In_377);
nand U1012 (N_1012,In_711,In_877);
or U1013 (N_1013,In_166,In_740);
nand U1014 (N_1014,In_402,In_554);
xnor U1015 (N_1015,In_604,In_1221);
or U1016 (N_1016,In_486,In_496);
nand U1017 (N_1017,In_499,In_477);
nand U1018 (N_1018,In_1187,In_716);
or U1019 (N_1019,In_506,In_310);
or U1020 (N_1020,In_525,In_1016);
nand U1021 (N_1021,In_1259,In_268);
nand U1022 (N_1022,In_1276,In_1385);
nor U1023 (N_1023,In_631,In_316);
nand U1024 (N_1024,In_264,In_1301);
or U1025 (N_1025,In_1233,In_714);
nand U1026 (N_1026,In_356,In_718);
and U1027 (N_1027,In_990,In_1339);
and U1028 (N_1028,In_306,In_879);
and U1029 (N_1029,In_1327,In_1037);
nor U1030 (N_1030,In_1020,In_1044);
or U1031 (N_1031,In_299,In_89);
nor U1032 (N_1032,In_1234,In_1389);
or U1033 (N_1033,In_1063,In_1298);
and U1034 (N_1034,In_287,In_1416);
xnor U1035 (N_1035,In_1244,In_48);
or U1036 (N_1036,In_1441,In_886);
nand U1037 (N_1037,In_104,In_159);
and U1038 (N_1038,In_898,In_1491);
or U1039 (N_1039,In_694,In_1072);
or U1040 (N_1040,In_1108,In_1282);
nand U1041 (N_1041,In_449,In_499);
or U1042 (N_1042,In_270,In_1326);
or U1043 (N_1043,In_1202,In_961);
or U1044 (N_1044,In_744,In_706);
and U1045 (N_1045,In_1282,In_603);
or U1046 (N_1046,In_807,In_1325);
nor U1047 (N_1047,In_1297,In_295);
or U1048 (N_1048,In_1468,In_1105);
nor U1049 (N_1049,In_1201,In_659);
xor U1050 (N_1050,In_871,In_630);
or U1051 (N_1051,In_538,In_766);
nor U1052 (N_1052,In_1469,In_367);
nor U1053 (N_1053,In_125,In_1409);
nor U1054 (N_1054,In_779,In_257);
nand U1055 (N_1055,In_31,In_909);
nand U1056 (N_1056,In_106,In_1357);
nand U1057 (N_1057,In_941,In_160);
or U1058 (N_1058,In_564,In_1267);
and U1059 (N_1059,In_755,In_1402);
nand U1060 (N_1060,In_990,In_1227);
nand U1061 (N_1061,In_1373,In_907);
nand U1062 (N_1062,In_1175,In_248);
nand U1063 (N_1063,In_710,In_1266);
or U1064 (N_1064,In_1445,In_915);
or U1065 (N_1065,In_638,In_185);
nor U1066 (N_1066,In_480,In_1405);
nor U1067 (N_1067,In_395,In_893);
or U1068 (N_1068,In_468,In_1453);
nand U1069 (N_1069,In_476,In_264);
and U1070 (N_1070,In_583,In_1332);
or U1071 (N_1071,In_304,In_1219);
nor U1072 (N_1072,In_338,In_529);
or U1073 (N_1073,In_1253,In_1302);
nor U1074 (N_1074,In_930,In_668);
nor U1075 (N_1075,In_1263,In_970);
or U1076 (N_1076,In_670,In_521);
nand U1077 (N_1077,In_1074,In_888);
nand U1078 (N_1078,In_668,In_906);
nand U1079 (N_1079,In_91,In_1276);
nor U1080 (N_1080,In_866,In_1054);
and U1081 (N_1081,In_795,In_0);
nand U1082 (N_1082,In_1405,In_1162);
xnor U1083 (N_1083,In_241,In_1298);
nor U1084 (N_1084,In_383,In_510);
and U1085 (N_1085,In_626,In_1088);
nor U1086 (N_1086,In_611,In_1362);
and U1087 (N_1087,In_571,In_847);
xor U1088 (N_1088,In_403,In_341);
nand U1089 (N_1089,In_848,In_874);
and U1090 (N_1090,In_1372,In_1127);
and U1091 (N_1091,In_440,In_268);
and U1092 (N_1092,In_343,In_1014);
or U1093 (N_1093,In_661,In_777);
xor U1094 (N_1094,In_720,In_321);
xor U1095 (N_1095,In_879,In_904);
and U1096 (N_1096,In_1227,In_1463);
nand U1097 (N_1097,In_523,In_693);
or U1098 (N_1098,In_14,In_721);
nand U1099 (N_1099,In_1422,In_772);
nand U1100 (N_1100,In_693,In_486);
and U1101 (N_1101,In_428,In_1233);
or U1102 (N_1102,In_944,In_1466);
nor U1103 (N_1103,In_224,In_397);
or U1104 (N_1104,In_297,In_284);
and U1105 (N_1105,In_475,In_1128);
or U1106 (N_1106,In_952,In_596);
nand U1107 (N_1107,In_986,In_1343);
or U1108 (N_1108,In_151,In_12);
or U1109 (N_1109,In_472,In_456);
or U1110 (N_1110,In_1470,In_98);
nor U1111 (N_1111,In_927,In_1006);
or U1112 (N_1112,In_1228,In_500);
or U1113 (N_1113,In_120,In_1057);
xor U1114 (N_1114,In_12,In_1137);
and U1115 (N_1115,In_543,In_1295);
nor U1116 (N_1116,In_573,In_206);
nand U1117 (N_1117,In_257,In_772);
nor U1118 (N_1118,In_251,In_944);
and U1119 (N_1119,In_168,In_918);
nand U1120 (N_1120,In_1259,In_1359);
nor U1121 (N_1121,In_120,In_446);
xnor U1122 (N_1122,In_598,In_112);
and U1123 (N_1123,In_1237,In_404);
and U1124 (N_1124,In_284,In_301);
nand U1125 (N_1125,In_94,In_615);
or U1126 (N_1126,In_830,In_1363);
nand U1127 (N_1127,In_518,In_497);
xnor U1128 (N_1128,In_138,In_692);
xor U1129 (N_1129,In_353,In_61);
nand U1130 (N_1130,In_262,In_1166);
nor U1131 (N_1131,In_253,In_1459);
nand U1132 (N_1132,In_1325,In_1242);
or U1133 (N_1133,In_1179,In_350);
nor U1134 (N_1134,In_1004,In_941);
and U1135 (N_1135,In_447,In_1196);
or U1136 (N_1136,In_1445,In_321);
and U1137 (N_1137,In_1468,In_1424);
xnor U1138 (N_1138,In_91,In_1209);
or U1139 (N_1139,In_404,In_1275);
or U1140 (N_1140,In_169,In_559);
or U1141 (N_1141,In_362,In_107);
nor U1142 (N_1142,In_652,In_262);
and U1143 (N_1143,In_191,In_143);
and U1144 (N_1144,In_1027,In_301);
or U1145 (N_1145,In_914,In_1484);
nor U1146 (N_1146,In_802,In_874);
nand U1147 (N_1147,In_1285,In_701);
nand U1148 (N_1148,In_129,In_1373);
nand U1149 (N_1149,In_1453,In_76);
or U1150 (N_1150,In_13,In_1086);
nor U1151 (N_1151,In_338,In_353);
or U1152 (N_1152,In_1232,In_464);
or U1153 (N_1153,In_1441,In_371);
or U1154 (N_1154,In_830,In_101);
or U1155 (N_1155,In_952,In_236);
nor U1156 (N_1156,In_218,In_132);
or U1157 (N_1157,In_228,In_1192);
and U1158 (N_1158,In_1344,In_1483);
xnor U1159 (N_1159,In_482,In_605);
xor U1160 (N_1160,In_164,In_126);
nand U1161 (N_1161,In_1112,In_333);
and U1162 (N_1162,In_1222,In_821);
nand U1163 (N_1163,In_1131,In_5);
nor U1164 (N_1164,In_1231,In_318);
nand U1165 (N_1165,In_597,In_875);
and U1166 (N_1166,In_537,In_402);
and U1167 (N_1167,In_1039,In_1366);
nand U1168 (N_1168,In_1175,In_1351);
or U1169 (N_1169,In_523,In_195);
and U1170 (N_1170,In_1164,In_483);
nor U1171 (N_1171,In_559,In_1051);
nand U1172 (N_1172,In_181,In_1021);
nor U1173 (N_1173,In_60,In_758);
or U1174 (N_1174,In_618,In_429);
and U1175 (N_1175,In_211,In_71);
and U1176 (N_1176,In_859,In_538);
and U1177 (N_1177,In_1252,In_147);
and U1178 (N_1178,In_1309,In_1184);
nor U1179 (N_1179,In_818,In_869);
and U1180 (N_1180,In_818,In_1333);
nor U1181 (N_1181,In_893,In_634);
and U1182 (N_1182,In_672,In_856);
or U1183 (N_1183,In_1292,In_101);
nor U1184 (N_1184,In_224,In_1000);
nor U1185 (N_1185,In_1136,In_1078);
xnor U1186 (N_1186,In_855,In_1391);
and U1187 (N_1187,In_1066,In_164);
nand U1188 (N_1188,In_286,In_451);
and U1189 (N_1189,In_942,In_950);
nand U1190 (N_1190,In_262,In_520);
nand U1191 (N_1191,In_906,In_1291);
nor U1192 (N_1192,In_900,In_620);
or U1193 (N_1193,In_89,In_143);
nand U1194 (N_1194,In_1349,In_1163);
and U1195 (N_1195,In_941,In_1188);
nand U1196 (N_1196,In_1435,In_853);
nor U1197 (N_1197,In_1263,In_987);
or U1198 (N_1198,In_394,In_1083);
nor U1199 (N_1199,In_703,In_112);
and U1200 (N_1200,In_1170,In_581);
nor U1201 (N_1201,In_827,In_155);
and U1202 (N_1202,In_1486,In_864);
nor U1203 (N_1203,In_556,In_1413);
nor U1204 (N_1204,In_1487,In_550);
or U1205 (N_1205,In_1434,In_1059);
and U1206 (N_1206,In_888,In_1441);
nor U1207 (N_1207,In_1351,In_1314);
or U1208 (N_1208,In_1464,In_861);
nand U1209 (N_1209,In_96,In_56);
nand U1210 (N_1210,In_94,In_435);
and U1211 (N_1211,In_867,In_124);
or U1212 (N_1212,In_871,In_343);
or U1213 (N_1213,In_858,In_64);
nor U1214 (N_1214,In_476,In_98);
nand U1215 (N_1215,In_951,In_528);
nand U1216 (N_1216,In_879,In_0);
nor U1217 (N_1217,In_571,In_832);
nor U1218 (N_1218,In_768,In_330);
and U1219 (N_1219,In_320,In_763);
or U1220 (N_1220,In_314,In_1171);
nand U1221 (N_1221,In_937,In_460);
and U1222 (N_1222,In_199,In_72);
nand U1223 (N_1223,In_122,In_181);
and U1224 (N_1224,In_1060,In_11);
nand U1225 (N_1225,In_110,In_903);
nand U1226 (N_1226,In_995,In_979);
and U1227 (N_1227,In_1123,In_282);
or U1228 (N_1228,In_27,In_1402);
nand U1229 (N_1229,In_1102,In_344);
nor U1230 (N_1230,In_781,In_1255);
nor U1231 (N_1231,In_596,In_1141);
and U1232 (N_1232,In_915,In_107);
or U1233 (N_1233,In_66,In_1139);
or U1234 (N_1234,In_1440,In_747);
or U1235 (N_1235,In_1461,In_1192);
nor U1236 (N_1236,In_1218,In_451);
and U1237 (N_1237,In_520,In_856);
nand U1238 (N_1238,In_1274,In_85);
or U1239 (N_1239,In_1080,In_565);
nor U1240 (N_1240,In_1135,In_74);
or U1241 (N_1241,In_4,In_1337);
xnor U1242 (N_1242,In_896,In_315);
nand U1243 (N_1243,In_960,In_1132);
and U1244 (N_1244,In_1420,In_1449);
nand U1245 (N_1245,In_1042,In_365);
and U1246 (N_1246,In_268,In_1199);
nand U1247 (N_1247,In_521,In_1256);
nor U1248 (N_1248,In_247,In_953);
nand U1249 (N_1249,In_660,In_782);
and U1250 (N_1250,In_542,In_587);
or U1251 (N_1251,In_699,In_626);
nand U1252 (N_1252,In_704,In_299);
or U1253 (N_1253,In_627,In_105);
and U1254 (N_1254,In_1430,In_1406);
nand U1255 (N_1255,In_861,In_1388);
or U1256 (N_1256,In_1357,In_1428);
nand U1257 (N_1257,In_935,In_1041);
nand U1258 (N_1258,In_1388,In_1390);
nand U1259 (N_1259,In_103,In_546);
or U1260 (N_1260,In_743,In_411);
and U1261 (N_1261,In_1345,In_557);
and U1262 (N_1262,In_317,In_132);
and U1263 (N_1263,In_1333,In_232);
and U1264 (N_1264,In_1131,In_1178);
nor U1265 (N_1265,In_1157,In_1387);
or U1266 (N_1266,In_933,In_869);
nand U1267 (N_1267,In_238,In_949);
or U1268 (N_1268,In_1314,In_1167);
nor U1269 (N_1269,In_92,In_184);
or U1270 (N_1270,In_462,In_263);
nand U1271 (N_1271,In_1249,In_1291);
nor U1272 (N_1272,In_1465,In_1281);
and U1273 (N_1273,In_825,In_1352);
nand U1274 (N_1274,In_1014,In_885);
and U1275 (N_1275,In_1332,In_504);
or U1276 (N_1276,In_424,In_719);
nor U1277 (N_1277,In_536,In_380);
nor U1278 (N_1278,In_1080,In_908);
or U1279 (N_1279,In_1015,In_1445);
nor U1280 (N_1280,In_801,In_569);
or U1281 (N_1281,In_629,In_398);
and U1282 (N_1282,In_271,In_1307);
or U1283 (N_1283,In_656,In_707);
nand U1284 (N_1284,In_281,In_313);
and U1285 (N_1285,In_1327,In_1086);
or U1286 (N_1286,In_1310,In_9);
nor U1287 (N_1287,In_1026,In_190);
nand U1288 (N_1288,In_1485,In_1250);
nand U1289 (N_1289,In_1102,In_182);
or U1290 (N_1290,In_1310,In_35);
nand U1291 (N_1291,In_1231,In_174);
and U1292 (N_1292,In_885,In_1209);
or U1293 (N_1293,In_1066,In_354);
or U1294 (N_1294,In_157,In_609);
nor U1295 (N_1295,In_980,In_432);
nor U1296 (N_1296,In_282,In_206);
nor U1297 (N_1297,In_896,In_679);
nor U1298 (N_1298,In_371,In_32);
nor U1299 (N_1299,In_908,In_1254);
or U1300 (N_1300,In_200,In_339);
nor U1301 (N_1301,In_1310,In_131);
nor U1302 (N_1302,In_801,In_1007);
and U1303 (N_1303,In_194,In_677);
nor U1304 (N_1304,In_450,In_666);
nor U1305 (N_1305,In_603,In_183);
nand U1306 (N_1306,In_887,In_828);
or U1307 (N_1307,In_1485,In_945);
nor U1308 (N_1308,In_12,In_999);
nor U1309 (N_1309,In_653,In_244);
nor U1310 (N_1310,In_534,In_352);
nor U1311 (N_1311,In_524,In_698);
nand U1312 (N_1312,In_876,In_509);
nor U1313 (N_1313,In_1119,In_734);
and U1314 (N_1314,In_727,In_1277);
or U1315 (N_1315,In_415,In_618);
nor U1316 (N_1316,In_353,In_380);
nand U1317 (N_1317,In_1003,In_78);
xor U1318 (N_1318,In_797,In_277);
or U1319 (N_1319,In_544,In_1101);
or U1320 (N_1320,In_506,In_1218);
nand U1321 (N_1321,In_639,In_297);
nand U1322 (N_1322,In_469,In_400);
or U1323 (N_1323,In_691,In_770);
or U1324 (N_1324,In_107,In_597);
and U1325 (N_1325,In_1101,In_198);
nor U1326 (N_1326,In_934,In_530);
nand U1327 (N_1327,In_269,In_554);
or U1328 (N_1328,In_1325,In_641);
and U1329 (N_1329,In_747,In_1041);
nor U1330 (N_1330,In_911,In_1138);
and U1331 (N_1331,In_1157,In_942);
and U1332 (N_1332,In_711,In_182);
or U1333 (N_1333,In_87,In_235);
nand U1334 (N_1334,In_335,In_972);
and U1335 (N_1335,In_985,In_1201);
and U1336 (N_1336,In_363,In_95);
or U1337 (N_1337,In_379,In_948);
or U1338 (N_1338,In_902,In_765);
or U1339 (N_1339,In_784,In_641);
or U1340 (N_1340,In_1111,In_226);
xor U1341 (N_1341,In_743,In_129);
or U1342 (N_1342,In_1213,In_361);
xor U1343 (N_1343,In_321,In_948);
nor U1344 (N_1344,In_811,In_932);
or U1345 (N_1345,In_958,In_1098);
or U1346 (N_1346,In_608,In_1238);
or U1347 (N_1347,In_764,In_590);
nand U1348 (N_1348,In_909,In_1132);
nand U1349 (N_1349,In_1395,In_670);
xor U1350 (N_1350,In_532,In_1002);
or U1351 (N_1351,In_1321,In_1290);
nor U1352 (N_1352,In_216,In_1009);
nor U1353 (N_1353,In_1321,In_114);
nor U1354 (N_1354,In_944,In_635);
nand U1355 (N_1355,In_1416,In_1043);
or U1356 (N_1356,In_1011,In_153);
or U1357 (N_1357,In_57,In_967);
nor U1358 (N_1358,In_1255,In_213);
and U1359 (N_1359,In_1450,In_520);
nand U1360 (N_1360,In_912,In_1265);
and U1361 (N_1361,In_1119,In_751);
nor U1362 (N_1362,In_868,In_444);
or U1363 (N_1363,In_143,In_39);
nand U1364 (N_1364,In_1379,In_1331);
or U1365 (N_1365,In_700,In_817);
nand U1366 (N_1366,In_357,In_780);
and U1367 (N_1367,In_295,In_946);
nand U1368 (N_1368,In_401,In_930);
nor U1369 (N_1369,In_23,In_1385);
nor U1370 (N_1370,In_1493,In_1453);
nand U1371 (N_1371,In_1427,In_241);
nor U1372 (N_1372,In_1321,In_1377);
nand U1373 (N_1373,In_581,In_172);
or U1374 (N_1374,In_1448,In_746);
xnor U1375 (N_1375,In_626,In_801);
nor U1376 (N_1376,In_728,In_176);
nor U1377 (N_1377,In_422,In_620);
nor U1378 (N_1378,In_346,In_68);
or U1379 (N_1379,In_743,In_1388);
and U1380 (N_1380,In_406,In_162);
nand U1381 (N_1381,In_1365,In_1046);
nor U1382 (N_1382,In_1033,In_168);
nor U1383 (N_1383,In_85,In_1314);
nand U1384 (N_1384,In_265,In_889);
nand U1385 (N_1385,In_1074,In_811);
and U1386 (N_1386,In_912,In_10);
nor U1387 (N_1387,In_1451,In_1287);
nor U1388 (N_1388,In_897,In_538);
and U1389 (N_1389,In_671,In_233);
nor U1390 (N_1390,In_1008,In_388);
nor U1391 (N_1391,In_456,In_298);
or U1392 (N_1392,In_1310,In_752);
nor U1393 (N_1393,In_1378,In_333);
or U1394 (N_1394,In_1114,In_1105);
nor U1395 (N_1395,In_207,In_1174);
nand U1396 (N_1396,In_1018,In_1347);
xnor U1397 (N_1397,In_1045,In_34);
and U1398 (N_1398,In_785,In_625);
and U1399 (N_1399,In_451,In_292);
and U1400 (N_1400,In_382,In_889);
or U1401 (N_1401,In_1486,In_660);
xor U1402 (N_1402,In_1404,In_1474);
nand U1403 (N_1403,In_434,In_308);
or U1404 (N_1404,In_1421,In_139);
nor U1405 (N_1405,In_1285,In_319);
nor U1406 (N_1406,In_782,In_996);
nor U1407 (N_1407,In_890,In_1451);
or U1408 (N_1408,In_276,In_1004);
nand U1409 (N_1409,In_559,In_1053);
nor U1410 (N_1410,In_837,In_942);
nand U1411 (N_1411,In_1015,In_1220);
xnor U1412 (N_1412,In_1343,In_130);
and U1413 (N_1413,In_1136,In_218);
nor U1414 (N_1414,In_1376,In_269);
or U1415 (N_1415,In_1480,In_1095);
and U1416 (N_1416,In_396,In_1434);
and U1417 (N_1417,In_794,In_1426);
or U1418 (N_1418,In_1268,In_1220);
nor U1419 (N_1419,In_604,In_436);
or U1420 (N_1420,In_91,In_637);
nor U1421 (N_1421,In_181,In_613);
or U1422 (N_1422,In_1089,In_471);
and U1423 (N_1423,In_55,In_837);
xor U1424 (N_1424,In_111,In_457);
nand U1425 (N_1425,In_1411,In_118);
nand U1426 (N_1426,In_1323,In_972);
xnor U1427 (N_1427,In_65,In_1418);
or U1428 (N_1428,In_1301,In_1478);
or U1429 (N_1429,In_873,In_559);
or U1430 (N_1430,In_1246,In_1021);
and U1431 (N_1431,In_1233,In_57);
nand U1432 (N_1432,In_294,In_305);
xor U1433 (N_1433,In_900,In_956);
nor U1434 (N_1434,In_969,In_188);
or U1435 (N_1435,In_528,In_1072);
nand U1436 (N_1436,In_1042,In_895);
and U1437 (N_1437,In_1366,In_912);
nor U1438 (N_1438,In_26,In_84);
nor U1439 (N_1439,In_117,In_155);
nand U1440 (N_1440,In_641,In_939);
nor U1441 (N_1441,In_726,In_652);
nand U1442 (N_1442,In_193,In_689);
nand U1443 (N_1443,In_874,In_675);
or U1444 (N_1444,In_149,In_752);
nand U1445 (N_1445,In_1168,In_859);
nor U1446 (N_1446,In_166,In_720);
nor U1447 (N_1447,In_35,In_1295);
nor U1448 (N_1448,In_723,In_1110);
nor U1449 (N_1449,In_1102,In_1166);
and U1450 (N_1450,In_596,In_1409);
nor U1451 (N_1451,In_382,In_1112);
and U1452 (N_1452,In_226,In_971);
or U1453 (N_1453,In_346,In_1288);
nand U1454 (N_1454,In_1332,In_566);
or U1455 (N_1455,In_60,In_157);
nor U1456 (N_1456,In_524,In_518);
nand U1457 (N_1457,In_695,In_955);
or U1458 (N_1458,In_566,In_345);
and U1459 (N_1459,In_1032,In_330);
nand U1460 (N_1460,In_185,In_1053);
and U1461 (N_1461,In_816,In_206);
and U1462 (N_1462,In_76,In_550);
and U1463 (N_1463,In_1494,In_987);
or U1464 (N_1464,In_1272,In_1230);
and U1465 (N_1465,In_283,In_310);
nor U1466 (N_1466,In_1312,In_1290);
nand U1467 (N_1467,In_527,In_70);
or U1468 (N_1468,In_21,In_559);
nand U1469 (N_1469,In_509,In_1093);
nand U1470 (N_1470,In_498,In_798);
nor U1471 (N_1471,In_931,In_749);
nor U1472 (N_1472,In_989,In_358);
nor U1473 (N_1473,In_1395,In_80);
nor U1474 (N_1474,In_616,In_164);
nand U1475 (N_1475,In_1055,In_1070);
nor U1476 (N_1476,In_317,In_1356);
nor U1477 (N_1477,In_1182,In_182);
nor U1478 (N_1478,In_507,In_1498);
nor U1479 (N_1479,In_1308,In_330);
nor U1480 (N_1480,In_292,In_76);
and U1481 (N_1481,In_1319,In_422);
nor U1482 (N_1482,In_642,In_36);
and U1483 (N_1483,In_1441,In_115);
nor U1484 (N_1484,In_1240,In_1060);
or U1485 (N_1485,In_304,In_1063);
nor U1486 (N_1486,In_847,In_545);
nand U1487 (N_1487,In_281,In_438);
or U1488 (N_1488,In_881,In_822);
nand U1489 (N_1489,In_692,In_7);
nor U1490 (N_1490,In_779,In_394);
nor U1491 (N_1491,In_1281,In_579);
nor U1492 (N_1492,In_1423,In_822);
or U1493 (N_1493,In_61,In_73);
nand U1494 (N_1494,In_144,In_1211);
and U1495 (N_1495,In_1169,In_369);
and U1496 (N_1496,In_1104,In_245);
and U1497 (N_1497,In_1098,In_468);
or U1498 (N_1498,In_168,In_513);
nand U1499 (N_1499,In_1021,In_1277);
or U1500 (N_1500,In_662,In_1038);
and U1501 (N_1501,In_632,In_864);
and U1502 (N_1502,In_220,In_1083);
nor U1503 (N_1503,In_323,In_82);
or U1504 (N_1504,In_756,In_1184);
and U1505 (N_1505,In_1223,In_804);
or U1506 (N_1506,In_244,In_245);
nand U1507 (N_1507,In_161,In_1275);
nand U1508 (N_1508,In_1438,In_31);
nor U1509 (N_1509,In_980,In_397);
and U1510 (N_1510,In_1287,In_915);
nand U1511 (N_1511,In_1427,In_1011);
or U1512 (N_1512,In_878,In_1359);
and U1513 (N_1513,In_1182,In_106);
nor U1514 (N_1514,In_725,In_213);
nand U1515 (N_1515,In_893,In_932);
nand U1516 (N_1516,In_1115,In_1248);
nand U1517 (N_1517,In_1246,In_156);
and U1518 (N_1518,In_1192,In_583);
or U1519 (N_1519,In_1165,In_199);
nand U1520 (N_1520,In_157,In_1214);
or U1521 (N_1521,In_1364,In_1310);
nand U1522 (N_1522,In_1247,In_1256);
nand U1523 (N_1523,In_102,In_1283);
nor U1524 (N_1524,In_1471,In_1423);
nand U1525 (N_1525,In_645,In_812);
or U1526 (N_1526,In_861,In_722);
nand U1527 (N_1527,In_32,In_156);
and U1528 (N_1528,In_1049,In_1111);
nor U1529 (N_1529,In_285,In_314);
nor U1530 (N_1530,In_847,In_231);
nor U1531 (N_1531,In_1266,In_231);
nor U1532 (N_1532,In_410,In_605);
or U1533 (N_1533,In_1063,In_1311);
nor U1534 (N_1534,In_838,In_50);
or U1535 (N_1535,In_943,In_1409);
xnor U1536 (N_1536,In_168,In_1099);
or U1537 (N_1537,In_1335,In_301);
nand U1538 (N_1538,In_631,In_1332);
nor U1539 (N_1539,In_1332,In_1045);
nor U1540 (N_1540,In_1354,In_1305);
nor U1541 (N_1541,In_1269,In_436);
and U1542 (N_1542,In_318,In_663);
or U1543 (N_1543,In_19,In_315);
and U1544 (N_1544,In_361,In_914);
nand U1545 (N_1545,In_711,In_332);
or U1546 (N_1546,In_1283,In_951);
or U1547 (N_1547,In_693,In_1184);
nand U1548 (N_1548,In_1239,In_427);
nor U1549 (N_1549,In_352,In_867);
nand U1550 (N_1550,In_540,In_803);
nand U1551 (N_1551,In_688,In_1167);
and U1552 (N_1552,In_379,In_259);
nor U1553 (N_1553,In_1297,In_648);
and U1554 (N_1554,In_1078,In_651);
and U1555 (N_1555,In_67,In_73);
nor U1556 (N_1556,In_1179,In_1408);
nand U1557 (N_1557,In_438,In_579);
or U1558 (N_1558,In_125,In_466);
or U1559 (N_1559,In_810,In_70);
nand U1560 (N_1560,In_1254,In_626);
nand U1561 (N_1561,In_488,In_1035);
or U1562 (N_1562,In_223,In_605);
and U1563 (N_1563,In_21,In_343);
and U1564 (N_1564,In_784,In_1035);
or U1565 (N_1565,In_716,In_415);
nand U1566 (N_1566,In_700,In_1357);
xor U1567 (N_1567,In_909,In_126);
or U1568 (N_1568,In_923,In_1221);
and U1569 (N_1569,In_527,In_396);
nand U1570 (N_1570,In_217,In_1388);
nor U1571 (N_1571,In_385,In_933);
or U1572 (N_1572,In_865,In_251);
nand U1573 (N_1573,In_1096,In_571);
and U1574 (N_1574,In_714,In_257);
or U1575 (N_1575,In_831,In_1218);
or U1576 (N_1576,In_363,In_1417);
nor U1577 (N_1577,In_727,In_610);
and U1578 (N_1578,In_1464,In_437);
or U1579 (N_1579,In_902,In_1203);
nor U1580 (N_1580,In_1273,In_644);
nand U1581 (N_1581,In_1468,In_1337);
and U1582 (N_1582,In_1453,In_312);
xor U1583 (N_1583,In_60,In_1445);
or U1584 (N_1584,In_1262,In_493);
or U1585 (N_1585,In_713,In_168);
nor U1586 (N_1586,In_1204,In_1364);
or U1587 (N_1587,In_323,In_1495);
or U1588 (N_1588,In_1408,In_1198);
and U1589 (N_1589,In_1303,In_334);
nand U1590 (N_1590,In_1347,In_264);
or U1591 (N_1591,In_295,In_146);
nor U1592 (N_1592,In_742,In_713);
and U1593 (N_1593,In_451,In_1420);
or U1594 (N_1594,In_1433,In_408);
and U1595 (N_1595,In_454,In_1297);
nor U1596 (N_1596,In_857,In_1397);
nor U1597 (N_1597,In_1442,In_393);
or U1598 (N_1598,In_1420,In_161);
or U1599 (N_1599,In_783,In_883);
and U1600 (N_1600,In_170,In_218);
nor U1601 (N_1601,In_1148,In_853);
nand U1602 (N_1602,In_657,In_501);
and U1603 (N_1603,In_101,In_1315);
nor U1604 (N_1604,In_171,In_204);
nor U1605 (N_1605,In_1444,In_191);
nor U1606 (N_1606,In_1135,In_1456);
nor U1607 (N_1607,In_102,In_193);
or U1608 (N_1608,In_802,In_1203);
nand U1609 (N_1609,In_1046,In_1008);
and U1610 (N_1610,In_1303,In_1085);
nand U1611 (N_1611,In_414,In_1263);
or U1612 (N_1612,In_1262,In_1232);
nand U1613 (N_1613,In_31,In_199);
or U1614 (N_1614,In_1429,In_1124);
nand U1615 (N_1615,In_398,In_344);
nand U1616 (N_1616,In_31,In_35);
and U1617 (N_1617,In_505,In_448);
and U1618 (N_1618,In_1485,In_938);
nor U1619 (N_1619,In_1441,In_777);
nor U1620 (N_1620,In_184,In_543);
and U1621 (N_1621,In_1242,In_844);
nor U1622 (N_1622,In_1431,In_1250);
nand U1623 (N_1623,In_723,In_912);
nor U1624 (N_1624,In_1149,In_975);
and U1625 (N_1625,In_104,In_1189);
nand U1626 (N_1626,In_36,In_429);
nand U1627 (N_1627,In_259,In_784);
nor U1628 (N_1628,In_1083,In_94);
nor U1629 (N_1629,In_767,In_335);
or U1630 (N_1630,In_1260,In_870);
and U1631 (N_1631,In_692,In_1018);
nor U1632 (N_1632,In_1098,In_113);
or U1633 (N_1633,In_10,In_457);
and U1634 (N_1634,In_171,In_609);
nor U1635 (N_1635,In_1446,In_659);
and U1636 (N_1636,In_1467,In_1310);
nor U1637 (N_1637,In_788,In_646);
or U1638 (N_1638,In_1106,In_1296);
nor U1639 (N_1639,In_1163,In_794);
nor U1640 (N_1640,In_856,In_37);
and U1641 (N_1641,In_1022,In_275);
nor U1642 (N_1642,In_1352,In_1470);
or U1643 (N_1643,In_367,In_111);
or U1644 (N_1644,In_1388,In_344);
nor U1645 (N_1645,In_394,In_616);
nand U1646 (N_1646,In_973,In_851);
or U1647 (N_1647,In_856,In_935);
or U1648 (N_1648,In_171,In_1406);
or U1649 (N_1649,In_1278,In_833);
nand U1650 (N_1650,In_1205,In_1396);
and U1651 (N_1651,In_1318,In_1113);
or U1652 (N_1652,In_524,In_180);
nor U1653 (N_1653,In_991,In_556);
xor U1654 (N_1654,In_161,In_949);
and U1655 (N_1655,In_645,In_1157);
xnor U1656 (N_1656,In_687,In_29);
nor U1657 (N_1657,In_388,In_1419);
or U1658 (N_1658,In_794,In_18);
nand U1659 (N_1659,In_1410,In_770);
nor U1660 (N_1660,In_1242,In_601);
nand U1661 (N_1661,In_1281,In_621);
and U1662 (N_1662,In_1331,In_446);
or U1663 (N_1663,In_822,In_73);
xor U1664 (N_1664,In_681,In_126);
or U1665 (N_1665,In_359,In_0);
xor U1666 (N_1666,In_1486,In_1344);
nor U1667 (N_1667,In_1153,In_1415);
and U1668 (N_1668,In_294,In_1038);
or U1669 (N_1669,In_288,In_348);
nand U1670 (N_1670,In_752,In_948);
nand U1671 (N_1671,In_757,In_71);
and U1672 (N_1672,In_876,In_1454);
nor U1673 (N_1673,In_1419,In_878);
nand U1674 (N_1674,In_967,In_871);
and U1675 (N_1675,In_908,In_838);
or U1676 (N_1676,In_936,In_555);
and U1677 (N_1677,In_873,In_54);
and U1678 (N_1678,In_101,In_988);
nand U1679 (N_1679,In_34,In_874);
and U1680 (N_1680,In_435,In_502);
nor U1681 (N_1681,In_1293,In_1350);
and U1682 (N_1682,In_580,In_1344);
nor U1683 (N_1683,In_410,In_258);
nor U1684 (N_1684,In_731,In_1382);
nor U1685 (N_1685,In_125,In_1345);
nor U1686 (N_1686,In_76,In_890);
or U1687 (N_1687,In_987,In_387);
nand U1688 (N_1688,In_494,In_860);
nor U1689 (N_1689,In_1207,In_770);
or U1690 (N_1690,In_180,In_60);
and U1691 (N_1691,In_931,In_668);
xor U1692 (N_1692,In_1323,In_1107);
nor U1693 (N_1693,In_1299,In_1089);
and U1694 (N_1694,In_835,In_684);
nor U1695 (N_1695,In_519,In_356);
nor U1696 (N_1696,In_185,In_1465);
nand U1697 (N_1697,In_1333,In_273);
nand U1698 (N_1698,In_264,In_541);
or U1699 (N_1699,In_502,In_986);
nand U1700 (N_1700,In_1137,In_737);
xor U1701 (N_1701,In_253,In_797);
and U1702 (N_1702,In_816,In_539);
or U1703 (N_1703,In_1071,In_320);
or U1704 (N_1704,In_974,In_1287);
nor U1705 (N_1705,In_948,In_99);
and U1706 (N_1706,In_149,In_1026);
nor U1707 (N_1707,In_1197,In_245);
nand U1708 (N_1708,In_1003,In_86);
and U1709 (N_1709,In_15,In_36);
nor U1710 (N_1710,In_901,In_1287);
or U1711 (N_1711,In_1088,In_388);
and U1712 (N_1712,In_554,In_488);
nor U1713 (N_1713,In_297,In_340);
and U1714 (N_1714,In_753,In_161);
nand U1715 (N_1715,In_1256,In_342);
nor U1716 (N_1716,In_137,In_257);
nor U1717 (N_1717,In_607,In_733);
or U1718 (N_1718,In_1190,In_1329);
nor U1719 (N_1719,In_808,In_545);
and U1720 (N_1720,In_1111,In_909);
nand U1721 (N_1721,In_527,In_99);
or U1722 (N_1722,In_1344,In_688);
nor U1723 (N_1723,In_568,In_1149);
and U1724 (N_1724,In_808,In_519);
and U1725 (N_1725,In_1366,In_498);
or U1726 (N_1726,In_424,In_1193);
and U1727 (N_1727,In_185,In_393);
and U1728 (N_1728,In_1340,In_739);
or U1729 (N_1729,In_1431,In_719);
or U1730 (N_1730,In_1066,In_1058);
nor U1731 (N_1731,In_511,In_616);
nand U1732 (N_1732,In_1363,In_591);
and U1733 (N_1733,In_578,In_383);
nand U1734 (N_1734,In_1266,In_167);
or U1735 (N_1735,In_974,In_1142);
and U1736 (N_1736,In_1388,In_1201);
nor U1737 (N_1737,In_798,In_841);
or U1738 (N_1738,In_462,In_1018);
nand U1739 (N_1739,In_119,In_1142);
and U1740 (N_1740,In_541,In_325);
and U1741 (N_1741,In_79,In_1204);
nor U1742 (N_1742,In_42,In_1378);
or U1743 (N_1743,In_261,In_1492);
nor U1744 (N_1744,In_111,In_1275);
and U1745 (N_1745,In_846,In_1052);
nand U1746 (N_1746,In_1383,In_903);
and U1747 (N_1747,In_464,In_345);
nand U1748 (N_1748,In_133,In_42);
and U1749 (N_1749,In_669,In_1209);
nand U1750 (N_1750,In_833,In_1301);
nor U1751 (N_1751,In_183,In_804);
nor U1752 (N_1752,In_1400,In_451);
nor U1753 (N_1753,In_1325,In_78);
xor U1754 (N_1754,In_330,In_82);
and U1755 (N_1755,In_123,In_1350);
nand U1756 (N_1756,In_919,In_1141);
and U1757 (N_1757,In_446,In_1360);
and U1758 (N_1758,In_43,In_798);
and U1759 (N_1759,In_659,In_356);
or U1760 (N_1760,In_283,In_1081);
and U1761 (N_1761,In_684,In_251);
nor U1762 (N_1762,In_813,In_1247);
nand U1763 (N_1763,In_396,In_217);
or U1764 (N_1764,In_1377,In_554);
nand U1765 (N_1765,In_1159,In_544);
nor U1766 (N_1766,In_980,In_822);
and U1767 (N_1767,In_1182,In_660);
nor U1768 (N_1768,In_1384,In_1400);
xnor U1769 (N_1769,In_1333,In_938);
and U1770 (N_1770,In_585,In_717);
and U1771 (N_1771,In_124,In_696);
or U1772 (N_1772,In_399,In_756);
or U1773 (N_1773,In_874,In_868);
nor U1774 (N_1774,In_279,In_236);
nand U1775 (N_1775,In_1463,In_1299);
nand U1776 (N_1776,In_1008,In_160);
nand U1777 (N_1777,In_1090,In_1459);
and U1778 (N_1778,In_769,In_1480);
nor U1779 (N_1779,In_527,In_811);
and U1780 (N_1780,In_1282,In_844);
or U1781 (N_1781,In_648,In_263);
and U1782 (N_1782,In_1368,In_131);
or U1783 (N_1783,In_576,In_587);
or U1784 (N_1784,In_374,In_1363);
nand U1785 (N_1785,In_1227,In_116);
and U1786 (N_1786,In_7,In_1325);
nand U1787 (N_1787,In_226,In_521);
xor U1788 (N_1788,In_214,In_913);
or U1789 (N_1789,In_246,In_1056);
and U1790 (N_1790,In_640,In_1495);
or U1791 (N_1791,In_1117,In_671);
nor U1792 (N_1792,In_1398,In_852);
nand U1793 (N_1793,In_949,In_346);
nand U1794 (N_1794,In_1332,In_905);
or U1795 (N_1795,In_476,In_823);
and U1796 (N_1796,In_1386,In_1462);
nor U1797 (N_1797,In_1070,In_1087);
nor U1798 (N_1798,In_1399,In_500);
nand U1799 (N_1799,In_1435,In_90);
nand U1800 (N_1800,In_1283,In_806);
nand U1801 (N_1801,In_1244,In_781);
and U1802 (N_1802,In_453,In_967);
nand U1803 (N_1803,In_470,In_709);
or U1804 (N_1804,In_4,In_333);
or U1805 (N_1805,In_874,In_31);
or U1806 (N_1806,In_270,In_809);
and U1807 (N_1807,In_1467,In_1275);
nand U1808 (N_1808,In_978,In_661);
nor U1809 (N_1809,In_642,In_717);
or U1810 (N_1810,In_938,In_1036);
nand U1811 (N_1811,In_1223,In_876);
or U1812 (N_1812,In_48,In_1385);
nor U1813 (N_1813,In_1200,In_935);
or U1814 (N_1814,In_780,In_1466);
nor U1815 (N_1815,In_384,In_74);
xor U1816 (N_1816,In_938,In_1161);
nand U1817 (N_1817,In_441,In_630);
nor U1818 (N_1818,In_872,In_1425);
nand U1819 (N_1819,In_1133,In_567);
nor U1820 (N_1820,In_795,In_785);
nand U1821 (N_1821,In_223,In_13);
xor U1822 (N_1822,In_129,In_682);
nor U1823 (N_1823,In_322,In_1116);
nor U1824 (N_1824,In_1041,In_143);
or U1825 (N_1825,In_267,In_1319);
or U1826 (N_1826,In_141,In_601);
or U1827 (N_1827,In_35,In_852);
or U1828 (N_1828,In_565,In_194);
nor U1829 (N_1829,In_712,In_744);
nor U1830 (N_1830,In_1284,In_79);
nand U1831 (N_1831,In_716,In_1403);
or U1832 (N_1832,In_1430,In_656);
nand U1833 (N_1833,In_599,In_1207);
nand U1834 (N_1834,In_153,In_1100);
or U1835 (N_1835,In_185,In_998);
nand U1836 (N_1836,In_674,In_186);
and U1837 (N_1837,In_1456,In_403);
or U1838 (N_1838,In_918,In_214);
xor U1839 (N_1839,In_861,In_431);
or U1840 (N_1840,In_1464,In_235);
nand U1841 (N_1841,In_104,In_1161);
nand U1842 (N_1842,In_228,In_745);
or U1843 (N_1843,In_700,In_268);
nor U1844 (N_1844,In_972,In_104);
nand U1845 (N_1845,In_1050,In_293);
nand U1846 (N_1846,In_955,In_120);
nor U1847 (N_1847,In_1314,In_1287);
xnor U1848 (N_1848,In_1214,In_375);
and U1849 (N_1849,In_1395,In_1463);
and U1850 (N_1850,In_326,In_584);
or U1851 (N_1851,In_1266,In_34);
nand U1852 (N_1852,In_610,In_1162);
or U1853 (N_1853,In_1184,In_938);
nor U1854 (N_1854,In_169,In_713);
nor U1855 (N_1855,In_401,In_894);
nor U1856 (N_1856,In_1207,In_1323);
nand U1857 (N_1857,In_1176,In_61);
or U1858 (N_1858,In_1356,In_1196);
and U1859 (N_1859,In_213,In_148);
and U1860 (N_1860,In_662,In_176);
and U1861 (N_1861,In_1258,In_646);
nand U1862 (N_1862,In_332,In_111);
and U1863 (N_1863,In_114,In_1240);
nand U1864 (N_1864,In_321,In_917);
nor U1865 (N_1865,In_1254,In_1348);
and U1866 (N_1866,In_370,In_1281);
nor U1867 (N_1867,In_1235,In_940);
or U1868 (N_1868,In_152,In_673);
nor U1869 (N_1869,In_1134,In_739);
or U1870 (N_1870,In_1239,In_1241);
or U1871 (N_1871,In_1276,In_505);
and U1872 (N_1872,In_606,In_329);
nand U1873 (N_1873,In_63,In_1177);
and U1874 (N_1874,In_707,In_100);
xnor U1875 (N_1875,In_24,In_2);
nor U1876 (N_1876,In_783,In_1383);
nand U1877 (N_1877,In_1493,In_378);
nand U1878 (N_1878,In_1486,In_296);
or U1879 (N_1879,In_860,In_987);
nor U1880 (N_1880,In_816,In_1326);
nor U1881 (N_1881,In_893,In_49);
and U1882 (N_1882,In_958,In_1439);
nor U1883 (N_1883,In_854,In_76);
or U1884 (N_1884,In_791,In_153);
nand U1885 (N_1885,In_1311,In_300);
or U1886 (N_1886,In_1435,In_670);
and U1887 (N_1887,In_562,In_1125);
nor U1888 (N_1888,In_769,In_205);
nor U1889 (N_1889,In_43,In_538);
nor U1890 (N_1890,In_1181,In_1099);
or U1891 (N_1891,In_1284,In_447);
or U1892 (N_1892,In_152,In_1237);
and U1893 (N_1893,In_1486,In_417);
or U1894 (N_1894,In_825,In_183);
nor U1895 (N_1895,In_1451,In_1077);
and U1896 (N_1896,In_723,In_108);
or U1897 (N_1897,In_1241,In_1336);
nor U1898 (N_1898,In_120,In_16);
and U1899 (N_1899,In_1262,In_701);
nor U1900 (N_1900,In_734,In_1207);
nand U1901 (N_1901,In_598,In_791);
nand U1902 (N_1902,In_25,In_799);
or U1903 (N_1903,In_968,In_1317);
or U1904 (N_1904,In_1431,In_1376);
nor U1905 (N_1905,In_145,In_1051);
or U1906 (N_1906,In_1252,In_260);
nor U1907 (N_1907,In_1107,In_1125);
nor U1908 (N_1908,In_959,In_698);
nand U1909 (N_1909,In_1073,In_287);
nor U1910 (N_1910,In_1090,In_628);
nand U1911 (N_1911,In_1481,In_1074);
nand U1912 (N_1912,In_540,In_272);
nor U1913 (N_1913,In_206,In_539);
nand U1914 (N_1914,In_52,In_612);
nand U1915 (N_1915,In_1408,In_1037);
or U1916 (N_1916,In_947,In_464);
xnor U1917 (N_1917,In_315,In_630);
and U1918 (N_1918,In_741,In_482);
nor U1919 (N_1919,In_971,In_1467);
or U1920 (N_1920,In_312,In_840);
nor U1921 (N_1921,In_523,In_909);
nor U1922 (N_1922,In_87,In_164);
and U1923 (N_1923,In_1201,In_824);
and U1924 (N_1924,In_63,In_536);
or U1925 (N_1925,In_92,In_940);
nor U1926 (N_1926,In_493,In_1140);
nand U1927 (N_1927,In_1466,In_333);
or U1928 (N_1928,In_431,In_695);
or U1929 (N_1929,In_540,In_556);
nor U1930 (N_1930,In_1029,In_985);
nor U1931 (N_1931,In_158,In_1134);
nand U1932 (N_1932,In_912,In_1037);
nand U1933 (N_1933,In_316,In_1004);
and U1934 (N_1934,In_1250,In_1017);
xor U1935 (N_1935,In_677,In_459);
or U1936 (N_1936,In_203,In_50);
and U1937 (N_1937,In_505,In_626);
nor U1938 (N_1938,In_1491,In_1075);
and U1939 (N_1939,In_199,In_846);
nor U1940 (N_1940,In_382,In_840);
and U1941 (N_1941,In_68,In_1436);
and U1942 (N_1942,In_424,In_1367);
nand U1943 (N_1943,In_1329,In_1114);
or U1944 (N_1944,In_746,In_278);
nand U1945 (N_1945,In_152,In_558);
nor U1946 (N_1946,In_1014,In_672);
nor U1947 (N_1947,In_126,In_1306);
and U1948 (N_1948,In_712,In_424);
nand U1949 (N_1949,In_189,In_1214);
nor U1950 (N_1950,In_429,In_996);
xor U1951 (N_1951,In_538,In_635);
xor U1952 (N_1952,In_624,In_38);
or U1953 (N_1953,In_1167,In_111);
nand U1954 (N_1954,In_1036,In_334);
or U1955 (N_1955,In_1020,In_705);
xnor U1956 (N_1956,In_318,In_203);
nand U1957 (N_1957,In_988,In_1066);
or U1958 (N_1958,In_1482,In_1486);
nand U1959 (N_1959,In_505,In_816);
or U1960 (N_1960,In_1047,In_128);
nand U1961 (N_1961,In_802,In_817);
or U1962 (N_1962,In_803,In_610);
or U1963 (N_1963,In_62,In_1400);
nor U1964 (N_1964,In_589,In_920);
or U1965 (N_1965,In_128,In_1363);
and U1966 (N_1966,In_1165,In_223);
or U1967 (N_1967,In_144,In_392);
or U1968 (N_1968,In_529,In_276);
and U1969 (N_1969,In_435,In_774);
or U1970 (N_1970,In_606,In_1046);
and U1971 (N_1971,In_768,In_698);
and U1972 (N_1972,In_1179,In_390);
and U1973 (N_1973,In_528,In_1096);
nand U1974 (N_1974,In_696,In_1012);
nor U1975 (N_1975,In_922,In_330);
nand U1976 (N_1976,In_1062,In_304);
nor U1977 (N_1977,In_764,In_722);
or U1978 (N_1978,In_915,In_237);
nor U1979 (N_1979,In_1436,In_1181);
nand U1980 (N_1980,In_830,In_935);
nor U1981 (N_1981,In_728,In_754);
nand U1982 (N_1982,In_635,In_340);
nand U1983 (N_1983,In_1112,In_691);
nor U1984 (N_1984,In_1385,In_974);
nand U1985 (N_1985,In_489,In_1232);
nand U1986 (N_1986,In_643,In_1191);
nand U1987 (N_1987,In_1228,In_1117);
nand U1988 (N_1988,In_64,In_1263);
and U1989 (N_1989,In_938,In_263);
nand U1990 (N_1990,In_1486,In_1086);
or U1991 (N_1991,In_1222,In_5);
nor U1992 (N_1992,In_1105,In_47);
nor U1993 (N_1993,In_822,In_901);
and U1994 (N_1994,In_640,In_824);
nor U1995 (N_1995,In_147,In_894);
nand U1996 (N_1996,In_1334,In_388);
nand U1997 (N_1997,In_840,In_856);
xnor U1998 (N_1998,In_1316,In_124);
xor U1999 (N_1999,In_916,In_974);
nand U2000 (N_2000,In_1268,In_1100);
and U2001 (N_2001,In_1125,In_1247);
nand U2002 (N_2002,In_827,In_467);
nand U2003 (N_2003,In_1483,In_589);
nand U2004 (N_2004,In_1393,In_723);
nand U2005 (N_2005,In_989,In_159);
nand U2006 (N_2006,In_793,In_753);
nor U2007 (N_2007,In_1401,In_1069);
or U2008 (N_2008,In_1186,In_482);
nand U2009 (N_2009,In_80,In_779);
or U2010 (N_2010,In_1284,In_740);
or U2011 (N_2011,In_1454,In_592);
nand U2012 (N_2012,In_783,In_937);
and U2013 (N_2013,In_71,In_1459);
and U2014 (N_2014,In_804,In_950);
nand U2015 (N_2015,In_569,In_1031);
or U2016 (N_2016,In_543,In_588);
nand U2017 (N_2017,In_190,In_1001);
or U2018 (N_2018,In_971,In_100);
nor U2019 (N_2019,In_43,In_1197);
or U2020 (N_2020,In_656,In_244);
and U2021 (N_2021,In_422,In_848);
nor U2022 (N_2022,In_241,In_1215);
or U2023 (N_2023,In_749,In_1177);
or U2024 (N_2024,In_1146,In_759);
nor U2025 (N_2025,In_395,In_1102);
or U2026 (N_2026,In_55,In_1351);
nor U2027 (N_2027,In_1213,In_172);
nand U2028 (N_2028,In_72,In_746);
nor U2029 (N_2029,In_681,In_982);
nand U2030 (N_2030,In_265,In_1411);
nor U2031 (N_2031,In_284,In_577);
nor U2032 (N_2032,In_1428,In_1007);
nand U2033 (N_2033,In_138,In_1452);
and U2034 (N_2034,In_915,In_1376);
nand U2035 (N_2035,In_456,In_1194);
nor U2036 (N_2036,In_298,In_803);
nor U2037 (N_2037,In_887,In_1362);
or U2038 (N_2038,In_1139,In_863);
and U2039 (N_2039,In_1301,In_815);
and U2040 (N_2040,In_1410,In_864);
nand U2041 (N_2041,In_275,In_67);
or U2042 (N_2042,In_1497,In_1224);
and U2043 (N_2043,In_1419,In_42);
or U2044 (N_2044,In_567,In_860);
nor U2045 (N_2045,In_901,In_1372);
nor U2046 (N_2046,In_254,In_66);
or U2047 (N_2047,In_1324,In_1315);
nor U2048 (N_2048,In_942,In_341);
nand U2049 (N_2049,In_100,In_1343);
and U2050 (N_2050,In_490,In_789);
or U2051 (N_2051,In_1459,In_1267);
or U2052 (N_2052,In_397,In_169);
nor U2053 (N_2053,In_1091,In_492);
nor U2054 (N_2054,In_1288,In_733);
or U2055 (N_2055,In_603,In_616);
and U2056 (N_2056,In_1066,In_1437);
nand U2057 (N_2057,In_434,In_45);
and U2058 (N_2058,In_1030,In_1243);
and U2059 (N_2059,In_1434,In_129);
nor U2060 (N_2060,In_1300,In_1369);
and U2061 (N_2061,In_997,In_1086);
nand U2062 (N_2062,In_518,In_76);
nor U2063 (N_2063,In_606,In_849);
or U2064 (N_2064,In_1172,In_443);
or U2065 (N_2065,In_1,In_379);
and U2066 (N_2066,In_568,In_416);
xnor U2067 (N_2067,In_343,In_697);
nor U2068 (N_2068,In_562,In_1006);
nand U2069 (N_2069,In_106,In_1344);
nand U2070 (N_2070,In_431,In_1467);
or U2071 (N_2071,In_431,In_888);
or U2072 (N_2072,In_86,In_365);
or U2073 (N_2073,In_130,In_1061);
and U2074 (N_2074,In_1386,In_508);
or U2075 (N_2075,In_1007,In_638);
and U2076 (N_2076,In_496,In_1100);
nor U2077 (N_2077,In_482,In_278);
or U2078 (N_2078,In_555,In_1160);
nor U2079 (N_2079,In_363,In_121);
nand U2080 (N_2080,In_1118,In_53);
or U2081 (N_2081,In_909,In_1426);
xor U2082 (N_2082,In_650,In_1392);
or U2083 (N_2083,In_623,In_458);
or U2084 (N_2084,In_456,In_182);
nand U2085 (N_2085,In_880,In_585);
nand U2086 (N_2086,In_1364,In_1253);
or U2087 (N_2087,In_178,In_740);
nand U2088 (N_2088,In_1258,In_608);
nor U2089 (N_2089,In_856,In_1147);
nand U2090 (N_2090,In_807,In_1031);
or U2091 (N_2091,In_1414,In_645);
nand U2092 (N_2092,In_699,In_695);
nor U2093 (N_2093,In_1170,In_986);
nand U2094 (N_2094,In_800,In_663);
nand U2095 (N_2095,In_312,In_279);
nand U2096 (N_2096,In_784,In_148);
nand U2097 (N_2097,In_1332,In_863);
or U2098 (N_2098,In_560,In_30);
nand U2099 (N_2099,In_1339,In_682);
or U2100 (N_2100,In_1285,In_293);
or U2101 (N_2101,In_537,In_1163);
nor U2102 (N_2102,In_1456,In_71);
nor U2103 (N_2103,In_1220,In_958);
nor U2104 (N_2104,In_1139,In_647);
nand U2105 (N_2105,In_688,In_129);
nand U2106 (N_2106,In_1077,In_716);
or U2107 (N_2107,In_363,In_1345);
and U2108 (N_2108,In_1251,In_1358);
nor U2109 (N_2109,In_676,In_1167);
or U2110 (N_2110,In_460,In_161);
and U2111 (N_2111,In_1244,In_113);
nand U2112 (N_2112,In_1458,In_195);
nor U2113 (N_2113,In_912,In_434);
and U2114 (N_2114,In_1296,In_79);
xor U2115 (N_2115,In_1025,In_320);
nand U2116 (N_2116,In_175,In_785);
nor U2117 (N_2117,In_787,In_627);
nor U2118 (N_2118,In_1372,In_1214);
nand U2119 (N_2119,In_1325,In_890);
and U2120 (N_2120,In_1320,In_1021);
or U2121 (N_2121,In_683,In_1473);
or U2122 (N_2122,In_971,In_903);
nor U2123 (N_2123,In_1387,In_1492);
nor U2124 (N_2124,In_1230,In_740);
and U2125 (N_2125,In_868,In_603);
xor U2126 (N_2126,In_49,In_816);
nor U2127 (N_2127,In_1268,In_1001);
and U2128 (N_2128,In_798,In_835);
and U2129 (N_2129,In_1442,In_239);
nor U2130 (N_2130,In_965,In_351);
or U2131 (N_2131,In_814,In_1210);
and U2132 (N_2132,In_590,In_115);
nand U2133 (N_2133,In_232,In_1161);
nand U2134 (N_2134,In_267,In_785);
nand U2135 (N_2135,In_1042,In_908);
or U2136 (N_2136,In_1032,In_1131);
nand U2137 (N_2137,In_180,In_295);
nor U2138 (N_2138,In_361,In_1406);
nand U2139 (N_2139,In_83,In_1393);
xnor U2140 (N_2140,In_947,In_137);
and U2141 (N_2141,In_922,In_1446);
and U2142 (N_2142,In_696,In_1070);
nor U2143 (N_2143,In_479,In_805);
and U2144 (N_2144,In_816,In_1042);
or U2145 (N_2145,In_541,In_1363);
nor U2146 (N_2146,In_816,In_330);
and U2147 (N_2147,In_498,In_879);
nor U2148 (N_2148,In_164,In_899);
or U2149 (N_2149,In_188,In_117);
nor U2150 (N_2150,In_858,In_1488);
nor U2151 (N_2151,In_869,In_1418);
or U2152 (N_2152,In_1221,In_532);
nand U2153 (N_2153,In_1063,In_1356);
nor U2154 (N_2154,In_420,In_857);
or U2155 (N_2155,In_731,In_1126);
nor U2156 (N_2156,In_1376,In_712);
or U2157 (N_2157,In_765,In_250);
and U2158 (N_2158,In_1247,In_1305);
nand U2159 (N_2159,In_543,In_1046);
nor U2160 (N_2160,In_651,In_1209);
or U2161 (N_2161,In_28,In_652);
nand U2162 (N_2162,In_699,In_257);
nand U2163 (N_2163,In_217,In_693);
nand U2164 (N_2164,In_1073,In_730);
nand U2165 (N_2165,In_406,In_559);
nand U2166 (N_2166,In_550,In_112);
or U2167 (N_2167,In_750,In_377);
or U2168 (N_2168,In_1121,In_471);
nand U2169 (N_2169,In_1269,In_1149);
nand U2170 (N_2170,In_978,In_585);
or U2171 (N_2171,In_1225,In_961);
nor U2172 (N_2172,In_13,In_917);
and U2173 (N_2173,In_825,In_1228);
nand U2174 (N_2174,In_952,In_1189);
nor U2175 (N_2175,In_1333,In_849);
or U2176 (N_2176,In_762,In_390);
or U2177 (N_2177,In_522,In_1069);
nand U2178 (N_2178,In_1142,In_1370);
nand U2179 (N_2179,In_876,In_1171);
and U2180 (N_2180,In_1020,In_1483);
nor U2181 (N_2181,In_1248,In_27);
nand U2182 (N_2182,In_248,In_75);
or U2183 (N_2183,In_978,In_1350);
and U2184 (N_2184,In_591,In_106);
or U2185 (N_2185,In_7,In_1135);
xnor U2186 (N_2186,In_410,In_404);
nor U2187 (N_2187,In_762,In_804);
nand U2188 (N_2188,In_37,In_1320);
or U2189 (N_2189,In_1110,In_377);
and U2190 (N_2190,In_852,In_936);
nand U2191 (N_2191,In_273,In_451);
nor U2192 (N_2192,In_1184,In_1402);
or U2193 (N_2193,In_122,In_1272);
nor U2194 (N_2194,In_764,In_1423);
and U2195 (N_2195,In_26,In_1246);
and U2196 (N_2196,In_277,In_1492);
nor U2197 (N_2197,In_469,In_120);
nor U2198 (N_2198,In_77,In_402);
and U2199 (N_2199,In_36,In_871);
and U2200 (N_2200,In_1355,In_428);
nor U2201 (N_2201,In_529,In_728);
and U2202 (N_2202,In_745,In_32);
nand U2203 (N_2203,In_482,In_468);
nand U2204 (N_2204,In_1475,In_885);
or U2205 (N_2205,In_483,In_194);
and U2206 (N_2206,In_330,In_788);
nand U2207 (N_2207,In_656,In_617);
nand U2208 (N_2208,In_566,In_418);
xor U2209 (N_2209,In_119,In_756);
or U2210 (N_2210,In_880,In_6);
and U2211 (N_2211,In_1101,In_342);
nand U2212 (N_2212,In_713,In_1144);
nand U2213 (N_2213,In_324,In_525);
nand U2214 (N_2214,In_821,In_218);
nand U2215 (N_2215,In_193,In_79);
or U2216 (N_2216,In_434,In_583);
nand U2217 (N_2217,In_1042,In_1165);
nand U2218 (N_2218,In_1222,In_324);
nand U2219 (N_2219,In_808,In_593);
and U2220 (N_2220,In_553,In_182);
or U2221 (N_2221,In_761,In_32);
nand U2222 (N_2222,In_661,In_800);
or U2223 (N_2223,In_1087,In_1439);
or U2224 (N_2224,In_1393,In_1268);
and U2225 (N_2225,In_257,In_980);
nor U2226 (N_2226,In_576,In_1264);
and U2227 (N_2227,In_121,In_812);
and U2228 (N_2228,In_281,In_148);
and U2229 (N_2229,In_1123,In_46);
and U2230 (N_2230,In_140,In_210);
nor U2231 (N_2231,In_299,In_1173);
and U2232 (N_2232,In_797,In_370);
or U2233 (N_2233,In_1244,In_697);
nand U2234 (N_2234,In_973,In_1227);
and U2235 (N_2235,In_259,In_859);
or U2236 (N_2236,In_511,In_222);
and U2237 (N_2237,In_175,In_1491);
nor U2238 (N_2238,In_58,In_751);
nand U2239 (N_2239,In_222,In_1410);
or U2240 (N_2240,In_1282,In_91);
xor U2241 (N_2241,In_52,In_1048);
nor U2242 (N_2242,In_657,In_611);
nor U2243 (N_2243,In_509,In_369);
and U2244 (N_2244,In_745,In_679);
nor U2245 (N_2245,In_301,In_312);
nor U2246 (N_2246,In_77,In_913);
nor U2247 (N_2247,In_1017,In_159);
nor U2248 (N_2248,In_1415,In_1172);
nand U2249 (N_2249,In_44,In_246);
or U2250 (N_2250,In_1240,In_802);
nand U2251 (N_2251,In_873,In_665);
or U2252 (N_2252,In_91,In_299);
and U2253 (N_2253,In_186,In_814);
nand U2254 (N_2254,In_578,In_612);
nor U2255 (N_2255,In_1413,In_134);
and U2256 (N_2256,In_530,In_783);
nand U2257 (N_2257,In_216,In_183);
nand U2258 (N_2258,In_408,In_288);
nand U2259 (N_2259,In_604,In_670);
nor U2260 (N_2260,In_44,In_1154);
and U2261 (N_2261,In_468,In_509);
nand U2262 (N_2262,In_821,In_561);
nor U2263 (N_2263,In_638,In_1306);
nor U2264 (N_2264,In_912,In_306);
nor U2265 (N_2265,In_733,In_1376);
nand U2266 (N_2266,In_1229,In_442);
or U2267 (N_2267,In_1166,In_214);
and U2268 (N_2268,In_473,In_971);
nand U2269 (N_2269,In_1145,In_1255);
or U2270 (N_2270,In_1223,In_1344);
nor U2271 (N_2271,In_211,In_286);
and U2272 (N_2272,In_1340,In_186);
nor U2273 (N_2273,In_877,In_973);
nor U2274 (N_2274,In_1483,In_718);
and U2275 (N_2275,In_316,In_103);
nor U2276 (N_2276,In_634,In_752);
nand U2277 (N_2277,In_192,In_807);
or U2278 (N_2278,In_551,In_1498);
and U2279 (N_2279,In_914,In_776);
xor U2280 (N_2280,In_1009,In_394);
nor U2281 (N_2281,In_1268,In_248);
or U2282 (N_2282,In_1178,In_262);
nor U2283 (N_2283,In_266,In_1396);
and U2284 (N_2284,In_257,In_1462);
and U2285 (N_2285,In_1020,In_221);
nor U2286 (N_2286,In_734,In_1339);
nor U2287 (N_2287,In_158,In_119);
nand U2288 (N_2288,In_1209,In_24);
xor U2289 (N_2289,In_1274,In_1298);
and U2290 (N_2290,In_255,In_1280);
or U2291 (N_2291,In_241,In_1410);
nor U2292 (N_2292,In_29,In_1288);
and U2293 (N_2293,In_162,In_493);
nor U2294 (N_2294,In_1108,In_1378);
or U2295 (N_2295,In_1421,In_532);
nor U2296 (N_2296,In_868,In_239);
and U2297 (N_2297,In_1412,In_217);
nand U2298 (N_2298,In_422,In_19);
nor U2299 (N_2299,In_729,In_937);
and U2300 (N_2300,In_1497,In_891);
or U2301 (N_2301,In_614,In_341);
nand U2302 (N_2302,In_1318,In_505);
nor U2303 (N_2303,In_256,In_759);
nand U2304 (N_2304,In_1266,In_1124);
or U2305 (N_2305,In_31,In_60);
nand U2306 (N_2306,In_931,In_318);
or U2307 (N_2307,In_472,In_605);
or U2308 (N_2308,In_349,In_141);
or U2309 (N_2309,In_557,In_682);
or U2310 (N_2310,In_1078,In_1391);
nor U2311 (N_2311,In_1300,In_843);
nor U2312 (N_2312,In_509,In_752);
and U2313 (N_2313,In_526,In_621);
or U2314 (N_2314,In_424,In_851);
or U2315 (N_2315,In_817,In_777);
xnor U2316 (N_2316,In_332,In_1478);
nor U2317 (N_2317,In_448,In_1213);
or U2318 (N_2318,In_955,In_1415);
nor U2319 (N_2319,In_854,In_91);
nor U2320 (N_2320,In_1338,In_1104);
and U2321 (N_2321,In_510,In_228);
nor U2322 (N_2322,In_945,In_76);
or U2323 (N_2323,In_1087,In_1260);
nand U2324 (N_2324,In_125,In_572);
nand U2325 (N_2325,In_632,In_479);
xor U2326 (N_2326,In_588,In_512);
or U2327 (N_2327,In_547,In_278);
and U2328 (N_2328,In_985,In_215);
nand U2329 (N_2329,In_361,In_1179);
nand U2330 (N_2330,In_633,In_317);
and U2331 (N_2331,In_462,In_238);
nor U2332 (N_2332,In_1428,In_239);
nand U2333 (N_2333,In_1237,In_499);
and U2334 (N_2334,In_1213,In_1480);
or U2335 (N_2335,In_1478,In_525);
or U2336 (N_2336,In_551,In_943);
nand U2337 (N_2337,In_114,In_389);
and U2338 (N_2338,In_1217,In_907);
or U2339 (N_2339,In_943,In_252);
and U2340 (N_2340,In_699,In_1461);
nand U2341 (N_2341,In_55,In_667);
or U2342 (N_2342,In_1019,In_1241);
or U2343 (N_2343,In_347,In_494);
and U2344 (N_2344,In_1197,In_367);
and U2345 (N_2345,In_1216,In_1328);
nor U2346 (N_2346,In_565,In_463);
nor U2347 (N_2347,In_1340,In_15);
nor U2348 (N_2348,In_1365,In_1134);
nand U2349 (N_2349,In_337,In_887);
nor U2350 (N_2350,In_1306,In_574);
or U2351 (N_2351,In_1087,In_1014);
nor U2352 (N_2352,In_578,In_230);
or U2353 (N_2353,In_571,In_800);
and U2354 (N_2354,In_1029,In_73);
nor U2355 (N_2355,In_371,In_943);
or U2356 (N_2356,In_493,In_1208);
nor U2357 (N_2357,In_77,In_872);
nor U2358 (N_2358,In_1227,In_1162);
nand U2359 (N_2359,In_1046,In_425);
or U2360 (N_2360,In_545,In_190);
or U2361 (N_2361,In_272,In_86);
or U2362 (N_2362,In_202,In_1279);
nor U2363 (N_2363,In_1194,In_1332);
and U2364 (N_2364,In_708,In_1369);
nor U2365 (N_2365,In_1279,In_604);
or U2366 (N_2366,In_144,In_1352);
or U2367 (N_2367,In_441,In_1482);
nor U2368 (N_2368,In_398,In_907);
xor U2369 (N_2369,In_768,In_489);
or U2370 (N_2370,In_834,In_1050);
nand U2371 (N_2371,In_583,In_772);
nor U2372 (N_2372,In_559,In_1489);
or U2373 (N_2373,In_931,In_340);
and U2374 (N_2374,In_703,In_1470);
or U2375 (N_2375,In_829,In_416);
and U2376 (N_2376,In_256,In_866);
xor U2377 (N_2377,In_921,In_793);
or U2378 (N_2378,In_918,In_903);
and U2379 (N_2379,In_257,In_966);
nand U2380 (N_2380,In_215,In_68);
nand U2381 (N_2381,In_452,In_247);
and U2382 (N_2382,In_641,In_1334);
nand U2383 (N_2383,In_1324,In_332);
or U2384 (N_2384,In_673,In_670);
and U2385 (N_2385,In_711,In_284);
nand U2386 (N_2386,In_897,In_743);
nor U2387 (N_2387,In_254,In_515);
and U2388 (N_2388,In_81,In_998);
nand U2389 (N_2389,In_19,In_847);
or U2390 (N_2390,In_1475,In_116);
and U2391 (N_2391,In_268,In_828);
nand U2392 (N_2392,In_50,In_661);
nor U2393 (N_2393,In_879,In_290);
or U2394 (N_2394,In_1299,In_877);
and U2395 (N_2395,In_1156,In_858);
and U2396 (N_2396,In_1000,In_1010);
nor U2397 (N_2397,In_520,In_806);
and U2398 (N_2398,In_620,In_1021);
and U2399 (N_2399,In_1078,In_105);
xnor U2400 (N_2400,In_786,In_553);
nand U2401 (N_2401,In_1173,In_950);
and U2402 (N_2402,In_314,In_450);
and U2403 (N_2403,In_550,In_480);
and U2404 (N_2404,In_721,In_280);
and U2405 (N_2405,In_571,In_1006);
or U2406 (N_2406,In_1462,In_424);
or U2407 (N_2407,In_156,In_1069);
and U2408 (N_2408,In_917,In_706);
nor U2409 (N_2409,In_1349,In_963);
nor U2410 (N_2410,In_977,In_894);
and U2411 (N_2411,In_567,In_1271);
nand U2412 (N_2412,In_565,In_313);
nor U2413 (N_2413,In_772,In_1005);
nand U2414 (N_2414,In_266,In_501);
nor U2415 (N_2415,In_804,In_352);
or U2416 (N_2416,In_1067,In_643);
or U2417 (N_2417,In_644,In_1373);
nor U2418 (N_2418,In_866,In_209);
nor U2419 (N_2419,In_1491,In_35);
or U2420 (N_2420,In_1352,In_409);
nand U2421 (N_2421,In_825,In_257);
and U2422 (N_2422,In_302,In_878);
nor U2423 (N_2423,In_332,In_952);
nor U2424 (N_2424,In_541,In_265);
and U2425 (N_2425,In_270,In_509);
nand U2426 (N_2426,In_305,In_513);
nand U2427 (N_2427,In_192,In_14);
nor U2428 (N_2428,In_1354,In_837);
or U2429 (N_2429,In_1184,In_1471);
nor U2430 (N_2430,In_693,In_578);
or U2431 (N_2431,In_1296,In_727);
or U2432 (N_2432,In_52,In_539);
nor U2433 (N_2433,In_597,In_1088);
nor U2434 (N_2434,In_1472,In_658);
nor U2435 (N_2435,In_943,In_8);
nand U2436 (N_2436,In_545,In_841);
or U2437 (N_2437,In_653,In_986);
nor U2438 (N_2438,In_816,In_850);
nor U2439 (N_2439,In_861,In_745);
nand U2440 (N_2440,In_850,In_1446);
and U2441 (N_2441,In_593,In_935);
nand U2442 (N_2442,In_21,In_716);
or U2443 (N_2443,In_619,In_895);
nand U2444 (N_2444,In_1226,In_504);
nor U2445 (N_2445,In_1062,In_1338);
or U2446 (N_2446,In_1386,In_800);
or U2447 (N_2447,In_979,In_1318);
nor U2448 (N_2448,In_456,In_277);
nand U2449 (N_2449,In_922,In_1166);
nor U2450 (N_2450,In_115,In_162);
xnor U2451 (N_2451,In_1253,In_516);
nor U2452 (N_2452,In_1344,In_1493);
or U2453 (N_2453,In_888,In_1062);
nand U2454 (N_2454,In_1241,In_1268);
and U2455 (N_2455,In_1076,In_341);
nand U2456 (N_2456,In_613,In_689);
nor U2457 (N_2457,In_757,In_1010);
and U2458 (N_2458,In_887,In_514);
or U2459 (N_2459,In_619,In_921);
or U2460 (N_2460,In_153,In_1347);
and U2461 (N_2461,In_726,In_294);
nor U2462 (N_2462,In_281,In_741);
or U2463 (N_2463,In_1311,In_590);
nor U2464 (N_2464,In_44,In_346);
nor U2465 (N_2465,In_646,In_313);
and U2466 (N_2466,In_1241,In_374);
nand U2467 (N_2467,In_12,In_1320);
or U2468 (N_2468,In_717,In_131);
or U2469 (N_2469,In_1229,In_1355);
or U2470 (N_2470,In_1235,In_407);
nand U2471 (N_2471,In_681,In_303);
xnor U2472 (N_2472,In_669,In_485);
and U2473 (N_2473,In_1489,In_329);
or U2474 (N_2474,In_299,In_513);
and U2475 (N_2475,In_1088,In_1456);
nor U2476 (N_2476,In_369,In_407);
nor U2477 (N_2477,In_294,In_85);
nor U2478 (N_2478,In_1000,In_1060);
nor U2479 (N_2479,In_297,In_408);
nor U2480 (N_2480,In_851,In_1159);
or U2481 (N_2481,In_58,In_565);
nor U2482 (N_2482,In_789,In_383);
nor U2483 (N_2483,In_1346,In_1340);
and U2484 (N_2484,In_1138,In_807);
nor U2485 (N_2485,In_952,In_924);
nor U2486 (N_2486,In_906,In_146);
or U2487 (N_2487,In_1067,In_1395);
or U2488 (N_2488,In_141,In_1248);
and U2489 (N_2489,In_893,In_1241);
and U2490 (N_2490,In_828,In_473);
nor U2491 (N_2491,In_448,In_1478);
nand U2492 (N_2492,In_463,In_1387);
nand U2493 (N_2493,In_1014,In_1490);
xnor U2494 (N_2494,In_286,In_480);
or U2495 (N_2495,In_763,In_1405);
or U2496 (N_2496,In_1092,In_385);
and U2497 (N_2497,In_1417,In_1060);
xnor U2498 (N_2498,In_256,In_1467);
nor U2499 (N_2499,In_554,In_810);
and U2500 (N_2500,In_1285,In_1121);
and U2501 (N_2501,In_277,In_712);
nand U2502 (N_2502,In_1099,In_394);
and U2503 (N_2503,In_364,In_841);
and U2504 (N_2504,In_801,In_467);
nor U2505 (N_2505,In_849,In_54);
nor U2506 (N_2506,In_711,In_667);
and U2507 (N_2507,In_1211,In_526);
nand U2508 (N_2508,In_1227,In_43);
and U2509 (N_2509,In_1033,In_509);
nand U2510 (N_2510,In_330,In_924);
and U2511 (N_2511,In_837,In_24);
nor U2512 (N_2512,In_473,In_508);
or U2513 (N_2513,In_25,In_694);
and U2514 (N_2514,In_300,In_620);
nor U2515 (N_2515,In_828,In_53);
or U2516 (N_2516,In_817,In_1105);
and U2517 (N_2517,In_817,In_513);
and U2518 (N_2518,In_806,In_385);
nor U2519 (N_2519,In_1108,In_366);
and U2520 (N_2520,In_1347,In_917);
or U2521 (N_2521,In_92,In_441);
xnor U2522 (N_2522,In_78,In_674);
nor U2523 (N_2523,In_945,In_670);
nand U2524 (N_2524,In_1047,In_362);
and U2525 (N_2525,In_104,In_1243);
and U2526 (N_2526,In_790,In_392);
and U2527 (N_2527,In_1015,In_738);
and U2528 (N_2528,In_724,In_1012);
nor U2529 (N_2529,In_236,In_500);
or U2530 (N_2530,In_1200,In_1334);
nand U2531 (N_2531,In_312,In_222);
or U2532 (N_2532,In_1192,In_1173);
nand U2533 (N_2533,In_784,In_175);
nor U2534 (N_2534,In_1003,In_228);
or U2535 (N_2535,In_939,In_1229);
and U2536 (N_2536,In_921,In_1424);
nor U2537 (N_2537,In_1088,In_1399);
xnor U2538 (N_2538,In_660,In_1298);
nand U2539 (N_2539,In_626,In_974);
nand U2540 (N_2540,In_370,In_123);
or U2541 (N_2541,In_1443,In_261);
nand U2542 (N_2542,In_1172,In_1025);
and U2543 (N_2543,In_1471,In_599);
nand U2544 (N_2544,In_783,In_1117);
nand U2545 (N_2545,In_47,In_551);
and U2546 (N_2546,In_386,In_34);
nor U2547 (N_2547,In_1028,In_53);
and U2548 (N_2548,In_8,In_623);
nand U2549 (N_2549,In_1386,In_30);
nor U2550 (N_2550,In_731,In_649);
or U2551 (N_2551,In_669,In_781);
nand U2552 (N_2552,In_392,In_1162);
or U2553 (N_2553,In_574,In_326);
nand U2554 (N_2554,In_7,In_1006);
nand U2555 (N_2555,In_1336,In_431);
or U2556 (N_2556,In_211,In_182);
nor U2557 (N_2557,In_1381,In_1026);
nand U2558 (N_2558,In_249,In_37);
or U2559 (N_2559,In_1303,In_518);
nor U2560 (N_2560,In_1384,In_439);
and U2561 (N_2561,In_1176,In_780);
and U2562 (N_2562,In_1024,In_717);
nand U2563 (N_2563,In_818,In_917);
or U2564 (N_2564,In_239,In_520);
or U2565 (N_2565,In_1383,In_1323);
nand U2566 (N_2566,In_412,In_695);
and U2567 (N_2567,In_142,In_562);
or U2568 (N_2568,In_118,In_485);
or U2569 (N_2569,In_969,In_1251);
nor U2570 (N_2570,In_505,In_19);
and U2571 (N_2571,In_205,In_1198);
nor U2572 (N_2572,In_138,In_703);
or U2573 (N_2573,In_1051,In_937);
or U2574 (N_2574,In_1486,In_1313);
and U2575 (N_2575,In_1367,In_1133);
nand U2576 (N_2576,In_1068,In_501);
or U2577 (N_2577,In_236,In_1098);
nor U2578 (N_2578,In_1280,In_1099);
or U2579 (N_2579,In_210,In_45);
nand U2580 (N_2580,In_731,In_821);
or U2581 (N_2581,In_583,In_421);
and U2582 (N_2582,In_267,In_1056);
nor U2583 (N_2583,In_1346,In_74);
and U2584 (N_2584,In_957,In_1208);
nand U2585 (N_2585,In_167,In_773);
nand U2586 (N_2586,In_542,In_810);
nand U2587 (N_2587,In_729,In_851);
nand U2588 (N_2588,In_143,In_1211);
and U2589 (N_2589,In_1067,In_1081);
nor U2590 (N_2590,In_1282,In_1372);
or U2591 (N_2591,In_290,In_349);
nand U2592 (N_2592,In_427,In_921);
nor U2593 (N_2593,In_1238,In_886);
or U2594 (N_2594,In_1098,In_987);
nor U2595 (N_2595,In_611,In_1152);
nand U2596 (N_2596,In_580,In_283);
or U2597 (N_2597,In_67,In_869);
nand U2598 (N_2598,In_139,In_2);
or U2599 (N_2599,In_48,In_559);
nand U2600 (N_2600,In_1418,In_1121);
nand U2601 (N_2601,In_205,In_1289);
xor U2602 (N_2602,In_1206,In_1045);
nor U2603 (N_2603,In_39,In_730);
nand U2604 (N_2604,In_1438,In_987);
and U2605 (N_2605,In_464,In_257);
nor U2606 (N_2606,In_764,In_667);
and U2607 (N_2607,In_1499,In_215);
and U2608 (N_2608,In_608,In_714);
nand U2609 (N_2609,In_849,In_1370);
and U2610 (N_2610,In_1429,In_403);
and U2611 (N_2611,In_1262,In_397);
nor U2612 (N_2612,In_247,In_893);
nand U2613 (N_2613,In_230,In_284);
nand U2614 (N_2614,In_692,In_740);
nand U2615 (N_2615,In_276,In_261);
or U2616 (N_2616,In_99,In_692);
or U2617 (N_2617,In_1258,In_1076);
or U2618 (N_2618,In_279,In_1096);
or U2619 (N_2619,In_1131,In_1278);
and U2620 (N_2620,In_1456,In_405);
nor U2621 (N_2621,In_0,In_1168);
xnor U2622 (N_2622,In_14,In_835);
nor U2623 (N_2623,In_1344,In_354);
nand U2624 (N_2624,In_778,In_1211);
nor U2625 (N_2625,In_8,In_1430);
nand U2626 (N_2626,In_618,In_495);
nand U2627 (N_2627,In_252,In_443);
nor U2628 (N_2628,In_975,In_1306);
and U2629 (N_2629,In_1355,In_927);
and U2630 (N_2630,In_1464,In_923);
nand U2631 (N_2631,In_825,In_665);
nor U2632 (N_2632,In_1185,In_929);
or U2633 (N_2633,In_782,In_957);
or U2634 (N_2634,In_602,In_724);
or U2635 (N_2635,In_626,In_328);
and U2636 (N_2636,In_1488,In_419);
or U2637 (N_2637,In_647,In_280);
xnor U2638 (N_2638,In_1411,In_151);
nor U2639 (N_2639,In_19,In_555);
xnor U2640 (N_2640,In_392,In_265);
nor U2641 (N_2641,In_648,In_1425);
nand U2642 (N_2642,In_904,In_570);
or U2643 (N_2643,In_247,In_1216);
and U2644 (N_2644,In_392,In_654);
or U2645 (N_2645,In_1188,In_659);
nand U2646 (N_2646,In_1,In_272);
nor U2647 (N_2647,In_820,In_235);
nor U2648 (N_2648,In_1302,In_758);
or U2649 (N_2649,In_580,In_748);
nor U2650 (N_2650,In_666,In_285);
nand U2651 (N_2651,In_760,In_1208);
nand U2652 (N_2652,In_398,In_917);
and U2653 (N_2653,In_1476,In_736);
and U2654 (N_2654,In_430,In_912);
nand U2655 (N_2655,In_1261,In_1110);
nand U2656 (N_2656,In_713,In_423);
and U2657 (N_2657,In_341,In_117);
nand U2658 (N_2658,In_1183,In_98);
and U2659 (N_2659,In_202,In_696);
xor U2660 (N_2660,In_398,In_345);
and U2661 (N_2661,In_40,In_438);
nand U2662 (N_2662,In_284,In_1039);
and U2663 (N_2663,In_772,In_974);
and U2664 (N_2664,In_691,In_1263);
nor U2665 (N_2665,In_95,In_644);
or U2666 (N_2666,In_1018,In_1239);
xnor U2667 (N_2667,In_17,In_1259);
and U2668 (N_2668,In_323,In_1458);
nand U2669 (N_2669,In_1484,In_1175);
or U2670 (N_2670,In_1403,In_423);
and U2671 (N_2671,In_1051,In_991);
nor U2672 (N_2672,In_557,In_1322);
nor U2673 (N_2673,In_794,In_1330);
nor U2674 (N_2674,In_1313,In_1495);
or U2675 (N_2675,In_913,In_672);
or U2676 (N_2676,In_13,In_52);
and U2677 (N_2677,In_682,In_462);
nor U2678 (N_2678,In_23,In_389);
nand U2679 (N_2679,In_1030,In_974);
nor U2680 (N_2680,In_421,In_447);
nand U2681 (N_2681,In_1399,In_614);
and U2682 (N_2682,In_1012,In_354);
nor U2683 (N_2683,In_399,In_1325);
nand U2684 (N_2684,In_1185,In_1073);
nor U2685 (N_2685,In_1493,In_933);
nand U2686 (N_2686,In_1381,In_1375);
or U2687 (N_2687,In_584,In_1371);
nand U2688 (N_2688,In_1343,In_551);
or U2689 (N_2689,In_818,In_511);
and U2690 (N_2690,In_1095,In_345);
nand U2691 (N_2691,In_1257,In_920);
nor U2692 (N_2692,In_1094,In_1177);
nand U2693 (N_2693,In_567,In_647);
nor U2694 (N_2694,In_1483,In_1355);
nand U2695 (N_2695,In_911,In_572);
nor U2696 (N_2696,In_1489,In_1432);
nor U2697 (N_2697,In_402,In_1122);
and U2698 (N_2698,In_428,In_116);
nand U2699 (N_2699,In_31,In_1392);
or U2700 (N_2700,In_669,In_92);
nand U2701 (N_2701,In_508,In_788);
or U2702 (N_2702,In_1232,In_1478);
or U2703 (N_2703,In_1364,In_146);
or U2704 (N_2704,In_901,In_13);
xor U2705 (N_2705,In_16,In_1270);
nand U2706 (N_2706,In_1150,In_214);
nand U2707 (N_2707,In_1003,In_1436);
nand U2708 (N_2708,In_985,In_1499);
nand U2709 (N_2709,In_854,In_422);
nor U2710 (N_2710,In_923,In_987);
and U2711 (N_2711,In_1116,In_815);
nand U2712 (N_2712,In_998,In_1079);
and U2713 (N_2713,In_141,In_711);
nand U2714 (N_2714,In_3,In_1042);
nand U2715 (N_2715,In_112,In_227);
or U2716 (N_2716,In_1034,In_1347);
nand U2717 (N_2717,In_1143,In_1138);
nand U2718 (N_2718,In_1160,In_140);
and U2719 (N_2719,In_1261,In_1401);
nor U2720 (N_2720,In_36,In_955);
nand U2721 (N_2721,In_1033,In_331);
and U2722 (N_2722,In_676,In_1045);
or U2723 (N_2723,In_1471,In_178);
or U2724 (N_2724,In_1456,In_1207);
and U2725 (N_2725,In_974,In_605);
nor U2726 (N_2726,In_633,In_874);
nor U2727 (N_2727,In_791,In_960);
or U2728 (N_2728,In_193,In_667);
and U2729 (N_2729,In_1291,In_513);
nor U2730 (N_2730,In_140,In_942);
or U2731 (N_2731,In_335,In_3);
and U2732 (N_2732,In_663,In_875);
nor U2733 (N_2733,In_571,In_867);
nand U2734 (N_2734,In_836,In_330);
or U2735 (N_2735,In_760,In_446);
and U2736 (N_2736,In_813,In_1492);
or U2737 (N_2737,In_985,In_280);
and U2738 (N_2738,In_1168,In_1244);
and U2739 (N_2739,In_297,In_118);
nor U2740 (N_2740,In_796,In_1213);
nand U2741 (N_2741,In_141,In_309);
nor U2742 (N_2742,In_1182,In_60);
or U2743 (N_2743,In_83,In_1398);
or U2744 (N_2744,In_834,In_1017);
or U2745 (N_2745,In_1156,In_418);
or U2746 (N_2746,In_1089,In_1406);
or U2747 (N_2747,In_922,In_1461);
nor U2748 (N_2748,In_1280,In_194);
nor U2749 (N_2749,In_1489,In_207);
or U2750 (N_2750,In_990,In_941);
nand U2751 (N_2751,In_100,In_1291);
or U2752 (N_2752,In_82,In_95);
or U2753 (N_2753,In_729,In_418);
nor U2754 (N_2754,In_373,In_220);
and U2755 (N_2755,In_759,In_946);
and U2756 (N_2756,In_1358,In_918);
nor U2757 (N_2757,In_719,In_1183);
or U2758 (N_2758,In_1004,In_1497);
nor U2759 (N_2759,In_1049,In_551);
and U2760 (N_2760,In_149,In_1029);
or U2761 (N_2761,In_297,In_286);
nor U2762 (N_2762,In_715,In_976);
and U2763 (N_2763,In_1340,In_1008);
or U2764 (N_2764,In_1432,In_361);
nand U2765 (N_2765,In_919,In_610);
xnor U2766 (N_2766,In_307,In_1166);
nand U2767 (N_2767,In_83,In_771);
or U2768 (N_2768,In_412,In_941);
or U2769 (N_2769,In_1428,In_1080);
and U2770 (N_2770,In_967,In_1358);
and U2771 (N_2771,In_346,In_6);
and U2772 (N_2772,In_1137,In_1254);
and U2773 (N_2773,In_1388,In_1406);
and U2774 (N_2774,In_794,In_1381);
and U2775 (N_2775,In_763,In_1426);
or U2776 (N_2776,In_87,In_211);
nor U2777 (N_2777,In_286,In_1346);
nor U2778 (N_2778,In_1360,In_119);
xnor U2779 (N_2779,In_1157,In_555);
or U2780 (N_2780,In_848,In_1427);
or U2781 (N_2781,In_1003,In_1356);
and U2782 (N_2782,In_1097,In_1195);
nand U2783 (N_2783,In_1424,In_1068);
nand U2784 (N_2784,In_88,In_1450);
and U2785 (N_2785,In_1110,In_146);
or U2786 (N_2786,In_36,In_1183);
nor U2787 (N_2787,In_1241,In_1498);
or U2788 (N_2788,In_23,In_523);
and U2789 (N_2789,In_990,In_421);
and U2790 (N_2790,In_557,In_16);
nand U2791 (N_2791,In_333,In_682);
nor U2792 (N_2792,In_1248,In_89);
nor U2793 (N_2793,In_730,In_1097);
nand U2794 (N_2794,In_138,In_966);
and U2795 (N_2795,In_588,In_60);
nor U2796 (N_2796,In_1388,In_1034);
nor U2797 (N_2797,In_329,In_1143);
nor U2798 (N_2798,In_718,In_344);
or U2799 (N_2799,In_693,In_301);
xor U2800 (N_2800,In_1356,In_1396);
nand U2801 (N_2801,In_1119,In_214);
or U2802 (N_2802,In_481,In_916);
xor U2803 (N_2803,In_46,In_137);
nand U2804 (N_2804,In_1193,In_330);
and U2805 (N_2805,In_565,In_281);
nor U2806 (N_2806,In_1194,In_1306);
and U2807 (N_2807,In_675,In_944);
and U2808 (N_2808,In_1006,In_1411);
or U2809 (N_2809,In_240,In_7);
nor U2810 (N_2810,In_454,In_164);
or U2811 (N_2811,In_275,In_143);
xor U2812 (N_2812,In_1435,In_572);
nor U2813 (N_2813,In_1481,In_321);
and U2814 (N_2814,In_1184,In_1302);
or U2815 (N_2815,In_844,In_352);
nor U2816 (N_2816,In_543,In_223);
nand U2817 (N_2817,In_27,In_275);
or U2818 (N_2818,In_391,In_122);
nor U2819 (N_2819,In_113,In_1093);
and U2820 (N_2820,In_631,In_780);
nor U2821 (N_2821,In_557,In_463);
nor U2822 (N_2822,In_88,In_1234);
or U2823 (N_2823,In_827,In_313);
nand U2824 (N_2824,In_323,In_1440);
or U2825 (N_2825,In_227,In_295);
xnor U2826 (N_2826,In_790,In_974);
nor U2827 (N_2827,In_1359,In_1495);
or U2828 (N_2828,In_913,In_1011);
or U2829 (N_2829,In_640,In_1104);
or U2830 (N_2830,In_1079,In_87);
nand U2831 (N_2831,In_989,In_888);
xnor U2832 (N_2832,In_110,In_1315);
or U2833 (N_2833,In_137,In_1107);
nor U2834 (N_2834,In_919,In_1344);
nor U2835 (N_2835,In_908,In_86);
and U2836 (N_2836,In_1212,In_1019);
or U2837 (N_2837,In_273,In_242);
nand U2838 (N_2838,In_422,In_1492);
nor U2839 (N_2839,In_175,In_1293);
or U2840 (N_2840,In_1277,In_1434);
or U2841 (N_2841,In_862,In_697);
and U2842 (N_2842,In_431,In_37);
or U2843 (N_2843,In_1297,In_121);
nand U2844 (N_2844,In_625,In_1363);
and U2845 (N_2845,In_150,In_610);
and U2846 (N_2846,In_69,In_4);
and U2847 (N_2847,In_1120,In_1075);
or U2848 (N_2848,In_147,In_537);
or U2849 (N_2849,In_1162,In_244);
nor U2850 (N_2850,In_569,In_1413);
or U2851 (N_2851,In_515,In_1234);
and U2852 (N_2852,In_848,In_1072);
nand U2853 (N_2853,In_597,In_1344);
nor U2854 (N_2854,In_554,In_715);
nor U2855 (N_2855,In_113,In_952);
and U2856 (N_2856,In_1467,In_771);
and U2857 (N_2857,In_945,In_270);
nor U2858 (N_2858,In_806,In_355);
nor U2859 (N_2859,In_819,In_455);
or U2860 (N_2860,In_358,In_797);
or U2861 (N_2861,In_25,In_864);
and U2862 (N_2862,In_510,In_608);
nand U2863 (N_2863,In_1155,In_369);
xor U2864 (N_2864,In_380,In_76);
nor U2865 (N_2865,In_100,In_1165);
nand U2866 (N_2866,In_577,In_52);
or U2867 (N_2867,In_161,In_525);
or U2868 (N_2868,In_52,In_1448);
xor U2869 (N_2869,In_668,In_1234);
nand U2870 (N_2870,In_1350,In_225);
nand U2871 (N_2871,In_803,In_375);
xor U2872 (N_2872,In_791,In_115);
nand U2873 (N_2873,In_759,In_1063);
xnor U2874 (N_2874,In_488,In_794);
xnor U2875 (N_2875,In_859,In_1194);
nand U2876 (N_2876,In_375,In_1008);
and U2877 (N_2877,In_1210,In_924);
nor U2878 (N_2878,In_1084,In_862);
nor U2879 (N_2879,In_845,In_644);
or U2880 (N_2880,In_569,In_283);
or U2881 (N_2881,In_91,In_49);
nand U2882 (N_2882,In_1314,In_1384);
nand U2883 (N_2883,In_272,In_1248);
nor U2884 (N_2884,In_100,In_1316);
or U2885 (N_2885,In_29,In_1332);
and U2886 (N_2886,In_1296,In_587);
nand U2887 (N_2887,In_363,In_571);
nand U2888 (N_2888,In_1078,In_240);
or U2889 (N_2889,In_539,In_146);
nor U2890 (N_2890,In_910,In_758);
nand U2891 (N_2891,In_1392,In_826);
nor U2892 (N_2892,In_316,In_655);
nor U2893 (N_2893,In_292,In_1148);
nor U2894 (N_2894,In_1217,In_1021);
or U2895 (N_2895,In_1175,In_1012);
or U2896 (N_2896,In_657,In_1157);
or U2897 (N_2897,In_611,In_282);
nand U2898 (N_2898,In_1406,In_216);
or U2899 (N_2899,In_950,In_564);
or U2900 (N_2900,In_323,In_1444);
or U2901 (N_2901,In_716,In_622);
nand U2902 (N_2902,In_1293,In_318);
or U2903 (N_2903,In_1204,In_1390);
and U2904 (N_2904,In_532,In_296);
or U2905 (N_2905,In_406,In_533);
or U2906 (N_2906,In_398,In_321);
or U2907 (N_2907,In_687,In_111);
and U2908 (N_2908,In_258,In_1091);
nor U2909 (N_2909,In_895,In_286);
nand U2910 (N_2910,In_483,In_721);
xor U2911 (N_2911,In_1033,In_1052);
nand U2912 (N_2912,In_241,In_1217);
nand U2913 (N_2913,In_1288,In_544);
and U2914 (N_2914,In_181,In_132);
xor U2915 (N_2915,In_314,In_202);
and U2916 (N_2916,In_599,In_777);
nor U2917 (N_2917,In_1131,In_568);
xor U2918 (N_2918,In_624,In_997);
nor U2919 (N_2919,In_281,In_1375);
or U2920 (N_2920,In_1133,In_210);
nand U2921 (N_2921,In_1071,In_388);
and U2922 (N_2922,In_594,In_600);
and U2923 (N_2923,In_1183,In_92);
or U2924 (N_2924,In_1143,In_1089);
xnor U2925 (N_2925,In_591,In_1477);
or U2926 (N_2926,In_669,In_95);
and U2927 (N_2927,In_109,In_513);
and U2928 (N_2928,In_1026,In_223);
and U2929 (N_2929,In_52,In_435);
and U2930 (N_2930,In_1166,In_784);
or U2931 (N_2931,In_1309,In_715);
or U2932 (N_2932,In_1340,In_1368);
nor U2933 (N_2933,In_166,In_480);
nor U2934 (N_2934,In_735,In_465);
and U2935 (N_2935,In_818,In_1450);
and U2936 (N_2936,In_870,In_18);
nor U2937 (N_2937,In_510,In_926);
and U2938 (N_2938,In_1373,In_1437);
or U2939 (N_2939,In_297,In_1479);
nor U2940 (N_2940,In_642,In_1223);
and U2941 (N_2941,In_144,In_1364);
nor U2942 (N_2942,In_14,In_1397);
nor U2943 (N_2943,In_1400,In_667);
nand U2944 (N_2944,In_805,In_1425);
nand U2945 (N_2945,In_617,In_100);
xor U2946 (N_2946,In_760,In_243);
nor U2947 (N_2947,In_761,In_1260);
nand U2948 (N_2948,In_1283,In_1235);
and U2949 (N_2949,In_921,In_1184);
and U2950 (N_2950,In_82,In_20);
and U2951 (N_2951,In_571,In_1132);
or U2952 (N_2952,In_1144,In_473);
nor U2953 (N_2953,In_1063,In_400);
nor U2954 (N_2954,In_690,In_932);
or U2955 (N_2955,In_1419,In_1394);
nor U2956 (N_2956,In_289,In_375);
or U2957 (N_2957,In_1294,In_1386);
and U2958 (N_2958,In_984,In_741);
nand U2959 (N_2959,In_349,In_332);
nor U2960 (N_2960,In_158,In_1016);
or U2961 (N_2961,In_1199,In_1246);
or U2962 (N_2962,In_791,In_26);
nor U2963 (N_2963,In_783,In_1365);
or U2964 (N_2964,In_982,In_210);
nor U2965 (N_2965,In_511,In_747);
or U2966 (N_2966,In_1333,In_614);
nor U2967 (N_2967,In_1028,In_727);
and U2968 (N_2968,In_1250,In_712);
or U2969 (N_2969,In_972,In_102);
or U2970 (N_2970,In_258,In_1064);
and U2971 (N_2971,In_226,In_632);
nand U2972 (N_2972,In_1000,In_593);
nand U2973 (N_2973,In_333,In_978);
nand U2974 (N_2974,In_991,In_400);
nand U2975 (N_2975,In_1420,In_503);
nand U2976 (N_2976,In_282,In_1091);
nand U2977 (N_2977,In_890,In_1305);
and U2978 (N_2978,In_177,In_296);
nor U2979 (N_2979,In_152,In_1034);
nand U2980 (N_2980,In_1087,In_266);
or U2981 (N_2981,In_378,In_1027);
nand U2982 (N_2982,In_883,In_342);
and U2983 (N_2983,In_1202,In_1479);
and U2984 (N_2984,In_894,In_830);
nor U2985 (N_2985,In_685,In_408);
and U2986 (N_2986,In_17,In_469);
or U2987 (N_2987,In_1168,In_537);
and U2988 (N_2988,In_511,In_1058);
nor U2989 (N_2989,In_1169,In_496);
and U2990 (N_2990,In_141,In_1022);
nand U2991 (N_2991,In_1062,In_696);
nand U2992 (N_2992,In_958,In_332);
or U2993 (N_2993,In_32,In_1378);
nand U2994 (N_2994,In_42,In_632);
and U2995 (N_2995,In_1206,In_804);
nand U2996 (N_2996,In_110,In_596);
and U2997 (N_2997,In_623,In_1112);
or U2998 (N_2998,In_790,In_1249);
or U2999 (N_2999,In_97,In_794);
or U3000 (N_3000,N_782,N_2263);
xnor U3001 (N_3001,N_2891,N_2833);
nor U3002 (N_3002,N_2397,N_972);
nor U3003 (N_3003,N_476,N_2754);
nand U3004 (N_3004,N_284,N_1341);
or U3005 (N_3005,N_1586,N_1089);
nor U3006 (N_3006,N_2528,N_64);
nor U3007 (N_3007,N_421,N_1969);
nand U3008 (N_3008,N_467,N_2423);
nand U3009 (N_3009,N_1285,N_470);
or U3010 (N_3010,N_672,N_334);
and U3011 (N_3011,N_2285,N_1434);
nand U3012 (N_3012,N_1303,N_127);
and U3013 (N_3013,N_1782,N_986);
nor U3014 (N_3014,N_1919,N_1231);
nand U3015 (N_3015,N_2934,N_712);
nand U3016 (N_3016,N_387,N_179);
and U3017 (N_3017,N_1554,N_425);
and U3018 (N_3018,N_2885,N_2452);
nand U3019 (N_3019,N_2957,N_1471);
nor U3020 (N_3020,N_1843,N_975);
or U3021 (N_3021,N_803,N_552);
and U3022 (N_3022,N_397,N_1062);
nand U3023 (N_3023,N_2499,N_1272);
nand U3024 (N_3024,N_978,N_227);
nand U3025 (N_3025,N_2883,N_579);
or U3026 (N_3026,N_1465,N_435);
and U3027 (N_3027,N_1882,N_120);
or U3028 (N_3028,N_2098,N_2215);
nand U3029 (N_3029,N_1731,N_2630);
nor U3030 (N_3030,N_1711,N_1803);
or U3031 (N_3031,N_2081,N_2448);
xnor U3032 (N_3032,N_1028,N_2677);
and U3033 (N_3033,N_598,N_2194);
xor U3034 (N_3034,N_2907,N_573);
or U3035 (N_3035,N_1794,N_2763);
nand U3036 (N_3036,N_2653,N_1440);
and U3037 (N_3037,N_1175,N_2616);
nor U3038 (N_3038,N_523,N_1823);
nand U3039 (N_3039,N_2935,N_1141);
nand U3040 (N_3040,N_1489,N_2968);
nor U3041 (N_3041,N_87,N_423);
or U3042 (N_3042,N_2994,N_2889);
xor U3043 (N_3043,N_502,N_2880);
and U3044 (N_3044,N_2472,N_2925);
or U3045 (N_3045,N_100,N_1431);
nand U3046 (N_3046,N_492,N_2627);
nand U3047 (N_3047,N_1599,N_1212);
nand U3048 (N_3048,N_2158,N_939);
nor U3049 (N_3049,N_2972,N_900);
nand U3050 (N_3050,N_1043,N_1490);
or U3051 (N_3051,N_335,N_2240);
or U3052 (N_3052,N_2720,N_1933);
nor U3053 (N_3053,N_165,N_633);
nor U3054 (N_3054,N_796,N_834);
nor U3055 (N_3055,N_1537,N_2013);
nor U3056 (N_3056,N_711,N_1940);
nor U3057 (N_3057,N_2118,N_1432);
nand U3058 (N_3058,N_2529,N_2679);
or U3059 (N_3059,N_657,N_327);
xnor U3060 (N_3060,N_2702,N_136);
or U3061 (N_3061,N_2817,N_866);
nor U3062 (N_3062,N_2888,N_2712);
nand U3063 (N_3063,N_2606,N_2212);
nand U3064 (N_3064,N_2143,N_1023);
and U3065 (N_3065,N_38,N_1099);
nor U3066 (N_3066,N_790,N_2183);
nor U3067 (N_3067,N_65,N_613);
and U3068 (N_3068,N_2553,N_1515);
nand U3069 (N_3069,N_482,N_1118);
nand U3070 (N_3070,N_2100,N_2947);
or U3071 (N_3071,N_715,N_2083);
or U3072 (N_3072,N_2485,N_1397);
and U3073 (N_3073,N_609,N_2929);
xnor U3074 (N_3074,N_1092,N_1138);
nand U3075 (N_3075,N_670,N_125);
and U3076 (N_3076,N_1759,N_2357);
nand U3077 (N_3077,N_1616,N_1946);
and U3078 (N_3078,N_1750,N_1693);
and U3079 (N_3079,N_2231,N_181);
nor U3080 (N_3080,N_36,N_1084);
or U3081 (N_3081,N_1646,N_649);
nand U3082 (N_3082,N_2569,N_692);
nand U3083 (N_3083,N_2159,N_2096);
nand U3084 (N_3084,N_1144,N_2905);
nand U3085 (N_3085,N_2807,N_704);
nor U3086 (N_3086,N_753,N_519);
or U3087 (N_3087,N_389,N_211);
nor U3088 (N_3088,N_708,N_437);
nor U3089 (N_3089,N_70,N_529);
and U3090 (N_3090,N_2172,N_539);
and U3091 (N_3091,N_743,N_1522);
nor U3092 (N_3092,N_2871,N_1863);
and U3093 (N_3093,N_1159,N_1547);
nor U3094 (N_3094,N_2146,N_2078);
and U3095 (N_3095,N_2654,N_2042);
and U3096 (N_3096,N_1565,N_2694);
and U3097 (N_3097,N_62,N_841);
nand U3098 (N_3098,N_1211,N_1247);
or U3099 (N_3099,N_1149,N_213);
and U3100 (N_3100,N_2649,N_1480);
and U3101 (N_3101,N_1900,N_2419);
nor U3102 (N_3102,N_113,N_1825);
nor U3103 (N_3103,N_2239,N_1716);
and U3104 (N_3104,N_989,N_1418);
or U3105 (N_3105,N_1333,N_2467);
nand U3106 (N_3106,N_1178,N_2281);
nor U3107 (N_3107,N_1326,N_373);
and U3108 (N_3108,N_1987,N_757);
nand U3109 (N_3109,N_2121,N_2208);
nand U3110 (N_3110,N_407,N_2801);
and U3111 (N_3111,N_655,N_2560);
or U3112 (N_3112,N_1475,N_2830);
nor U3113 (N_3113,N_1888,N_688);
nor U3114 (N_3114,N_808,N_2797);
or U3115 (N_3115,N_1009,N_945);
nor U3116 (N_3116,N_2303,N_675);
nor U3117 (N_3117,N_2005,N_1730);
and U3118 (N_3118,N_325,N_1602);
and U3119 (N_3119,N_1678,N_2837);
or U3120 (N_3120,N_1464,N_72);
nand U3121 (N_3121,N_2267,N_1820);
nor U3122 (N_3122,N_1064,N_542);
or U3123 (N_3123,N_2374,N_1875);
and U3124 (N_3124,N_2603,N_261);
or U3125 (N_3125,N_2794,N_488);
nor U3126 (N_3126,N_318,N_651);
nor U3127 (N_3127,N_172,N_2761);
nor U3128 (N_3128,N_1074,N_2021);
nand U3129 (N_3129,N_415,N_22);
nor U3130 (N_3130,N_668,N_2946);
and U3131 (N_3131,N_178,N_196);
and U3132 (N_3132,N_1133,N_1265);
nor U3133 (N_3133,N_1577,N_281);
and U3134 (N_3134,N_1007,N_2373);
nand U3135 (N_3135,N_910,N_99);
and U3136 (N_3136,N_2219,N_1421);
nand U3137 (N_3137,N_53,N_164);
and U3138 (N_3138,N_2381,N_357);
nand U3139 (N_3139,N_2813,N_2524);
nand U3140 (N_3140,N_2298,N_2044);
nand U3141 (N_3141,N_1327,N_1637);
nand U3142 (N_3142,N_1839,N_2046);
nor U3143 (N_3143,N_1787,N_2953);
and U3144 (N_3144,N_684,N_1708);
nand U3145 (N_3145,N_1792,N_2256);
nand U3146 (N_3146,N_2597,N_1562);
or U3147 (N_3147,N_1136,N_471);
or U3148 (N_3148,N_1992,N_2144);
and U3149 (N_3149,N_1758,N_755);
nand U3150 (N_3150,N_746,N_1891);
nand U3151 (N_3151,N_1512,N_880);
or U3152 (N_3152,N_163,N_2908);
nand U3153 (N_3153,N_1015,N_2362);
and U3154 (N_3154,N_1184,N_951);
and U3155 (N_3155,N_1558,N_162);
nor U3156 (N_3156,N_703,N_1228);
and U3157 (N_3157,N_2402,N_1776);
nand U3158 (N_3158,N_2189,N_1568);
nor U3159 (N_3159,N_1544,N_671);
or U3160 (N_3160,N_665,N_915);
and U3161 (N_3161,N_408,N_2293);
nand U3162 (N_3162,N_266,N_760);
nor U3163 (N_3163,N_2490,N_1328);
nor U3164 (N_3164,N_1923,N_2228);
and U3165 (N_3165,N_1504,N_13);
nor U3166 (N_3166,N_2344,N_438);
xnor U3167 (N_3167,N_52,N_1438);
nor U3168 (N_3168,N_1106,N_117);
and U3169 (N_3169,N_355,N_999);
or U3170 (N_3170,N_931,N_93);
and U3171 (N_3171,N_2138,N_2136);
and U3172 (N_3172,N_1514,N_1619);
and U3173 (N_3173,N_2253,N_454);
nor U3174 (N_3174,N_1350,N_2310);
nand U3175 (N_3175,N_67,N_1194);
nor U3176 (N_3176,N_991,N_933);
or U3177 (N_3177,N_565,N_1035);
and U3178 (N_3178,N_2699,N_37);
nand U3179 (N_3179,N_2409,N_1456);
or U3180 (N_3180,N_1393,N_1296);
xnor U3181 (N_3181,N_2437,N_2148);
nor U3182 (N_3182,N_1847,N_1835);
and U3183 (N_3183,N_98,N_2909);
and U3184 (N_3184,N_43,N_2950);
nand U3185 (N_3185,N_2930,N_2024);
and U3186 (N_3186,N_733,N_1713);
or U3187 (N_3187,N_2967,N_1202);
nand U3188 (N_3188,N_1830,N_1760);
nand U3189 (N_3189,N_1698,N_1983);
and U3190 (N_3190,N_1498,N_1058);
nor U3191 (N_3191,N_2716,N_2886);
and U3192 (N_3192,N_922,N_1310);
nor U3193 (N_3193,N_2713,N_546);
or U3194 (N_3194,N_1376,N_1061);
or U3195 (N_3195,N_2488,N_16);
nand U3196 (N_3196,N_2345,N_617);
or U3197 (N_3197,N_2459,N_371);
nor U3198 (N_3198,N_914,N_1429);
nor U3199 (N_3199,N_63,N_2273);
nand U3200 (N_3200,N_2951,N_1487);
nor U3201 (N_3201,N_647,N_2846);
nor U3202 (N_3202,N_1679,N_1234);
nand U3203 (N_3203,N_1103,N_2390);
nor U3204 (N_3204,N_1628,N_584);
nand U3205 (N_3205,N_2366,N_1420);
or U3206 (N_3206,N_304,N_2764);
and U3207 (N_3207,N_1896,N_1805);
nor U3208 (N_3208,N_2386,N_2068);
or U3209 (N_3209,N_2657,N_1137);
and U3210 (N_3210,N_1907,N_2135);
and U3211 (N_3211,N_1351,N_484);
and U3212 (N_3212,N_2161,N_1812);
or U3213 (N_3213,N_126,N_2855);
nor U3214 (N_3214,N_2703,N_2401);
nand U3215 (N_3215,N_771,N_2475);
or U3216 (N_3216,N_1460,N_1986);
nand U3217 (N_3217,N_2970,N_909);
nand U3218 (N_3218,N_2006,N_1689);
nand U3219 (N_3219,N_2035,N_2000);
or U3220 (N_3220,N_83,N_2014);
nor U3221 (N_3221,N_728,N_851);
nand U3222 (N_3222,N_223,N_1171);
and U3223 (N_3223,N_2230,N_890);
nor U3224 (N_3224,N_1183,N_1337);
and U3225 (N_3225,N_2268,N_1871);
and U3226 (N_3226,N_868,N_2457);
and U3227 (N_3227,N_1786,N_509);
nand U3228 (N_3228,N_2988,N_2640);
or U3229 (N_3229,N_1281,N_1564);
nor U3230 (N_3230,N_1959,N_124);
nand U3231 (N_3231,N_1380,N_554);
nor U3232 (N_3232,N_2085,N_2261);
xor U3233 (N_3233,N_938,N_2382);
nand U3234 (N_3234,N_450,N_2019);
or U3235 (N_3235,N_2308,N_2283);
nor U3236 (N_3236,N_1665,N_255);
nor U3237 (N_3237,N_1469,N_1849);
nand U3238 (N_3238,N_2567,N_1260);
nand U3239 (N_3239,N_2999,N_436);
nand U3240 (N_3240,N_953,N_754);
or U3241 (N_3241,N_2140,N_800);
and U3242 (N_3242,N_528,N_904);
nand U3243 (N_3243,N_2965,N_2609);
and U3244 (N_3244,N_1790,N_1248);
nor U3245 (N_3245,N_2119,N_1755);
and U3246 (N_3246,N_2915,N_602);
nor U3247 (N_3247,N_2549,N_2070);
and U3248 (N_3248,N_1629,N_342);
nand U3249 (N_3249,N_987,N_12);
or U3250 (N_3250,N_1675,N_252);
nand U3251 (N_3251,N_535,N_1415);
or U3252 (N_3252,N_2949,N_2058);
and U3253 (N_3253,N_2760,N_858);
and U3254 (N_3254,N_2464,N_1978);
nor U3255 (N_3255,N_2975,N_385);
or U3256 (N_3256,N_1065,N_420);
or U3257 (N_3257,N_2828,N_2132);
nor U3258 (N_3258,N_2103,N_1917);
and U3259 (N_3259,N_2963,N_1170);
xor U3260 (N_3260,N_2288,N_2184);
nand U3261 (N_3261,N_1697,N_1266);
nor U3262 (N_3262,N_630,N_1941);
or U3263 (N_3263,N_935,N_226);
xor U3264 (N_3264,N_1439,N_1404);
nor U3265 (N_3265,N_849,N_1717);
nor U3266 (N_3266,N_1683,N_644);
or U3267 (N_3267,N_620,N_2432);
nand U3268 (N_3268,N_2449,N_925);
and U3269 (N_3269,N_2856,N_738);
nand U3270 (N_3270,N_2751,N_1390);
nor U3271 (N_3271,N_1254,N_225);
nor U3272 (N_3272,N_2595,N_1667);
or U3273 (N_3273,N_1041,N_1507);
xor U3274 (N_3274,N_1867,N_2433);
and U3275 (N_3275,N_1233,N_1278);
nor U3276 (N_3276,N_2789,N_1014);
nand U3277 (N_3277,N_375,N_2061);
nand U3278 (N_3278,N_1344,N_430);
nor U3279 (N_3279,N_2196,N_2167);
or U3280 (N_3280,N_1597,N_2107);
nand U3281 (N_3281,N_974,N_958);
and U3282 (N_3282,N_446,N_71);
or U3283 (N_3283,N_2723,N_802);
or U3284 (N_3284,N_1673,N_1771);
and U3285 (N_3285,N_1524,N_2139);
or U3286 (N_3286,N_869,N_201);
or U3287 (N_3287,N_2580,N_795);
and U3288 (N_3288,N_68,N_706);
and U3289 (N_3289,N_2768,N_2708);
or U3290 (N_3290,N_1088,N_1077);
nand U3291 (N_3291,N_2496,N_57);
or U3292 (N_3292,N_537,N_1966);
or U3293 (N_3293,N_2665,N_727);
nor U3294 (N_3294,N_2666,N_1476);
or U3295 (N_3295,N_831,N_2939);
and U3296 (N_3296,N_253,N_2769);
and U3297 (N_3297,N_964,N_534);
and U3298 (N_3298,N_2474,N_929);
or U3299 (N_3299,N_612,N_2674);
nor U3300 (N_3300,N_320,N_97);
or U3301 (N_3301,N_1880,N_76);
nand U3302 (N_3302,N_2351,N_2274);
and U3303 (N_3303,N_2910,N_2495);
and U3304 (N_3304,N_1611,N_639);
nand U3305 (N_3305,N_1095,N_2927);
nand U3306 (N_3306,N_2105,N_1243);
nor U3307 (N_3307,N_1938,N_2180);
xnor U3308 (N_3308,N_597,N_2384);
or U3309 (N_3309,N_2914,N_607);
nand U3310 (N_3310,N_2672,N_2901);
and U3311 (N_3311,N_2557,N_2340);
nand U3312 (N_3312,N_513,N_1063);
nand U3313 (N_3313,N_1899,N_17);
nor U3314 (N_3314,N_992,N_589);
nor U3315 (N_3315,N_1040,N_2541);
and U3316 (N_3316,N_517,N_2259);
nor U3317 (N_3317,N_1798,N_547);
or U3318 (N_3318,N_353,N_702);
and U3319 (N_3319,N_1180,N_739);
nor U3320 (N_3320,N_1027,N_2408);
or U3321 (N_3321,N_1943,N_1579);
and U3322 (N_3322,N_369,N_1773);
or U3323 (N_3323,N_2932,N_182);
and U3324 (N_3324,N_242,N_2727);
or U3325 (N_3325,N_2550,N_326);
or U3326 (N_3326,N_824,N_440);
nand U3327 (N_3327,N_2337,N_1594);
xor U3328 (N_3328,N_2015,N_26);
nand U3329 (N_3329,N_2395,N_1079);
nor U3330 (N_3330,N_891,N_409);
nor U3331 (N_3331,N_2733,N_1988);
or U3332 (N_3332,N_1696,N_1687);
nand U3333 (N_3333,N_1046,N_235);
or U3334 (N_3334,N_525,N_1898);
nand U3335 (N_3335,N_215,N_1459);
and U3336 (N_3336,N_526,N_1056);
and U3337 (N_3337,N_2063,N_2181);
nand U3338 (N_3338,N_1383,N_2434);
and U3339 (N_3339,N_246,N_1080);
and U3340 (N_3340,N_2282,N_751);
nand U3341 (N_3341,N_2348,N_2387);
nand U3342 (N_3342,N_2556,N_2793);
or U3343 (N_3343,N_2808,N_1906);
nand U3344 (N_3344,N_2882,N_347);
or U3345 (N_3345,N_2077,N_1268);
nand U3346 (N_3346,N_1370,N_1030);
nand U3347 (N_3347,N_2466,N_2695);
nor U3348 (N_3348,N_2091,N_2523);
nand U3349 (N_3349,N_2349,N_1883);
nor U3350 (N_3350,N_2329,N_112);
nor U3351 (N_3351,N_1740,N_2564);
nand U3352 (N_3352,N_2027,N_1197);
and U3353 (N_3353,N_1378,N_1783);
nor U3354 (N_3354,N_146,N_604);
nand U3355 (N_3355,N_1997,N_1779);
nor U3356 (N_3356,N_1831,N_530);
and U3357 (N_3357,N_394,N_2581);
nand U3358 (N_3358,N_645,N_399);
and U3359 (N_3359,N_2859,N_2185);
and U3360 (N_3360,N_2637,N_2418);
nor U3361 (N_3361,N_2048,N_1976);
nand U3362 (N_3362,N_2037,N_2735);
and U3363 (N_3363,N_1734,N_1904);
nand U3364 (N_3364,N_937,N_966);
nand U3365 (N_3365,N_853,N_475);
and U3366 (N_3366,N_2451,N_2060);
nand U3367 (N_3367,N_2179,N_901);
and U3368 (N_3368,N_2050,N_9);
xor U3369 (N_3369,N_204,N_581);
nand U3370 (N_3370,N_1190,N_562);
nand U3371 (N_3371,N_264,N_1625);
nand U3372 (N_3372,N_228,N_2290);
and U3373 (N_3373,N_2617,N_2810);
or U3374 (N_3374,N_973,N_2300);
or U3375 (N_3375,N_289,N_638);
or U3376 (N_3376,N_1336,N_2217);
nor U3377 (N_3377,N_902,N_2029);
nand U3378 (N_3378,N_1642,N_449);
nand U3379 (N_3379,N_810,N_2403);
nand U3380 (N_3380,N_1405,N_1176);
nand U3381 (N_3381,N_263,N_2691);
or U3382 (N_3382,N_156,N_1712);
and U3383 (N_3383,N_1008,N_1146);
nand U3384 (N_3384,N_969,N_683);
or U3385 (N_3385,N_2704,N_1198);
and U3386 (N_3386,N_536,N_2728);
nand U3387 (N_3387,N_2811,N_1715);
and U3388 (N_3388,N_2527,N_1105);
and U3389 (N_3389,N_2088,N_1321);
or U3390 (N_3390,N_2056,N_781);
nor U3391 (N_3391,N_1879,N_48);
nor U3392 (N_3392,N_701,N_2547);
and U3393 (N_3393,N_2854,N_1935);
or U3394 (N_3394,N_2770,N_1513);
and U3395 (N_3395,N_1042,N_1339);
nor U3396 (N_3396,N_777,N_2791);
nor U3397 (N_3397,N_7,N_1723);
and U3398 (N_3398,N_2201,N_1873);
and U3399 (N_3399,N_2780,N_1525);
nand U3400 (N_3400,N_871,N_2752);
and U3401 (N_3401,N_600,N_451);
nand U3402 (N_3402,N_734,N_1800);
and U3403 (N_3403,N_1727,N_20);
nor U3404 (N_3404,N_2235,N_1261);
or U3405 (N_3405,N_2198,N_2645);
xor U3406 (N_3406,N_2683,N_431);
or U3407 (N_3407,N_981,N_985);
and U3408 (N_3408,N_1177,N_2876);
or U3409 (N_3409,N_2945,N_1038);
nand U3410 (N_3410,N_898,N_1414);
and U3411 (N_3411,N_2004,N_2725);
and U3412 (N_3412,N_2842,N_761);
nor U3413 (N_3413,N_1214,N_2410);
or U3414 (N_3414,N_485,N_1477);
nand U3415 (N_3415,N_2636,N_216);
and U3416 (N_3416,N_2250,N_1705);
or U3417 (N_3417,N_150,N_1618);
or U3418 (N_3418,N_1312,N_2921);
and U3419 (N_3419,N_2090,N_310);
nand U3420 (N_3420,N_1129,N_1559);
nor U3421 (N_3421,N_1290,N_2203);
nor U3422 (N_3422,N_128,N_1340);
and U3423 (N_3423,N_846,N_1529);
and U3424 (N_3424,N_386,N_2629);
or U3425 (N_3425,N_2193,N_908);
nor U3426 (N_3426,N_2772,N_884);
nor U3427 (N_3427,N_1990,N_283);
or U3428 (N_3428,N_131,N_1965);
and U3429 (N_3429,N_1520,N_141);
nor U3430 (N_3430,N_280,N_2598);
nand U3431 (N_3431,N_2835,N_2894);
or U3432 (N_3432,N_1454,N_586);
nor U3433 (N_3433,N_1767,N_578);
and U3434 (N_3434,N_2851,N_2788);
nand U3435 (N_3435,N_2822,N_1864);
or U3436 (N_3436,N_927,N_2758);
or U3437 (N_3437,N_2840,N_726);
or U3438 (N_3438,N_1195,N_1004);
nand U3439 (N_3439,N_877,N_2530);
and U3440 (N_3440,N_2361,N_873);
nor U3441 (N_3441,N_393,N_434);
nor U3442 (N_3442,N_1098,N_1242);
nor U3443 (N_3443,N_2831,N_1603);
nor U3444 (N_3444,N_2229,N_1109);
or U3445 (N_3445,N_153,N_1848);
nand U3446 (N_3446,N_833,N_561);
nand U3447 (N_3447,N_1349,N_158);
and U3448 (N_3448,N_835,N_2919);
nor U3449 (N_3449,N_1001,N_1430);
nor U3450 (N_3450,N_319,N_1196);
or U3451 (N_3451,N_2347,N_2848);
and U3452 (N_3452,N_2570,N_2426);
or U3453 (N_3453,N_247,N_527);
xnor U3454 (N_3454,N_2336,N_1838);
or U3455 (N_3455,N_1968,N_2912);
and U3456 (N_3456,N_524,N_1914);
or U3457 (N_3457,N_2425,N_35);
nor U3458 (N_3458,N_2514,N_2613);
or U3459 (N_3459,N_1122,N_2540);
and U3460 (N_3460,N_286,N_2631);
or U3461 (N_3461,N_1235,N_2860);
or U3462 (N_3462,N_2818,N_2322);
nand U3463 (N_3463,N_2978,N_961);
and U3464 (N_3464,N_205,N_1829);
or U3465 (N_3465,N_1925,N_2572);
nor U3466 (N_3466,N_2486,N_149);
nor U3467 (N_3467,N_1467,N_2221);
or U3468 (N_3468,N_2320,N_220);
and U3469 (N_3469,N_2753,N_2684);
or U3470 (N_3470,N_2985,N_190);
or U3471 (N_3471,N_241,N_2987);
nand U3472 (N_3472,N_2034,N_2507);
nand U3473 (N_3473,N_291,N_2031);
and U3474 (N_3474,N_1449,N_1424);
nor U3475 (N_3475,N_934,N_1240);
nor U3476 (N_3476,N_2623,N_1018);
and U3477 (N_3477,N_2815,N_404);
or U3478 (N_3478,N_742,N_2385);
or U3479 (N_3479,N_1182,N_370);
nand U3480 (N_3480,N_2800,N_1039);
nand U3481 (N_3481,N_2602,N_1259);
or U3482 (N_3482,N_2120,N_2324);
and U3483 (N_3483,N_277,N_2421);
and U3484 (N_3484,N_222,N_236);
or U3485 (N_3485,N_1550,N_2380);
nor U3486 (N_3486,N_693,N_480);
and U3487 (N_3487,N_1412,N_1486);
and U3488 (N_3488,N_2454,N_1590);
nor U3489 (N_3489,N_1518,N_1125);
nor U3490 (N_3490,N_1895,N_997);
or U3491 (N_3491,N_576,N_1656);
nor U3492 (N_3492,N_154,N_270);
and U3493 (N_3493,N_1435,N_1016);
and U3494 (N_3494,N_1273,N_2620);
xnor U3495 (N_3495,N_151,N_2295);
nor U3496 (N_3496,N_231,N_2600);
nor U3497 (N_3497,N_2424,N_2717);
or U3498 (N_3498,N_1037,N_1457);
and U3499 (N_3499,N_1905,N_29);
or U3500 (N_3500,N_234,N_40);
and U3501 (N_3501,N_2829,N_957);
or U3502 (N_3502,N_1720,N_1609);
or U3503 (N_3503,N_823,N_1617);
and U3504 (N_3504,N_721,N_2497);
nor U3505 (N_3505,N_1366,N_1192);
or U3506 (N_3506,N_427,N_621);
and U3507 (N_3507,N_2786,N_1506);
nand U3508 (N_3508,N_1497,N_2825);
and U3509 (N_3509,N_2151,N_1021);
and U3510 (N_3510,N_1725,N_248);
nand U3511 (N_3511,N_1657,N_1494);
nand U3512 (N_3512,N_696,N_2095);
nor U3513 (N_3513,N_1174,N_1870);
nand U3514 (N_3514,N_41,N_1142);
nor U3515 (N_3515,N_122,N_1269);
xor U3516 (N_3516,N_1299,N_794);
and U3517 (N_3517,N_1499,N_2160);
or U3518 (N_3518,N_949,N_744);
nor U3519 (N_3519,N_1592,N_198);
and U3520 (N_3520,N_2644,N_2589);
nand U3521 (N_3521,N_2494,N_1294);
nor U3522 (N_3522,N_510,N_2745);
nor U3523 (N_3523,N_2413,N_1956);
or U3524 (N_3524,N_2591,N_89);
or U3525 (N_3525,N_1680,N_1822);
or U3526 (N_3526,N_2548,N_2099);
or U3527 (N_3527,N_1502,N_109);
or U3528 (N_3528,N_1574,N_1277);
and U3529 (N_3529,N_1119,N_1381);
or U3530 (N_3530,N_2918,N_243);
or U3531 (N_3531,N_1655,N_555);
and U3532 (N_3532,N_1833,N_2022);
and U3533 (N_3533,N_88,N_1630);
or U3534 (N_3534,N_2202,N_1691);
nand U3535 (N_3535,N_1958,N_1924);
nand U3536 (N_3536,N_2671,N_2785);
nand U3537 (N_3537,N_160,N_1495);
nor U3538 (N_3538,N_82,N_115);
nor U3539 (N_3539,N_741,N_923);
nor U3540 (N_3540,N_2370,N_2513);
nor U3541 (N_3541,N_2043,N_1156);
and U3542 (N_3542,N_1379,N_1582);
and U3543 (N_3543,N_1926,N_2872);
or U3544 (N_3544,N_2371,N_1868);
or U3545 (N_3545,N_2109,N_2162);
or U3546 (N_3546,N_2359,N_1066);
nand U3547 (N_3547,N_1053,N_2481);
xnor U3548 (N_3548,N_219,N_1663);
and U3549 (N_3549,N_1560,N_134);
or U3550 (N_3550,N_1633,N_2510);
nor U3551 (N_3551,N_1401,N_2590);
nor U3552 (N_3552,N_918,N_2059);
nand U3553 (N_3553,N_1036,N_1073);
nand U3554 (N_3554,N_2866,N_1410);
or U3555 (N_3555,N_2269,N_570);
or U3556 (N_3556,N_2920,N_368);
and U3557 (N_3557,N_59,N_79);
or U3558 (N_3558,N_1396,N_2933);
nand U3559 (N_3559,N_1521,N_424);
and U3560 (N_3560,N_155,N_148);
nand U3561 (N_3561,N_518,N_316);
or U3562 (N_3562,N_874,N_784);
and U3563 (N_3563,N_1892,N_1912);
xor U3564 (N_3564,N_1911,N_1082);
nor U3565 (N_3565,N_2445,N_1112);
nor U3566 (N_3566,N_322,N_1793);
nor U3567 (N_3567,N_770,N_2803);
or U3568 (N_3568,N_658,N_2688);
nand U3569 (N_3569,N_1121,N_1885);
or U3570 (N_3570,N_2304,N_129);
or U3571 (N_3571,N_1527,N_60);
nand U3572 (N_3572,N_2440,N_2960);
xor U3573 (N_3573,N_1050,N_1147);
or U3574 (N_3574,N_372,N_2465);
nand U3575 (N_3575,N_2664,N_2869);
nand U3576 (N_3576,N_2177,N_1332);
nand U3577 (N_3577,N_383,N_2565);
xor U3578 (N_3578,N_865,N_1484);
nor U3579 (N_3579,N_2102,N_952);
or U3580 (N_3580,N_1881,N_1069);
and U3581 (N_3581,N_1749,N_723);
nand U3582 (N_3582,N_585,N_1827);
or U3583 (N_3583,N_2777,N_2321);
or U3584 (N_3584,N_2016,N_1186);
nor U3585 (N_3585,N_2325,N_1011);
and U3586 (N_3586,N_1950,N_2149);
or U3587 (N_3587,N_186,N_2864);
nand U3588 (N_3588,N_1491,N_736);
or U3589 (N_3589,N_844,N_1160);
and U3590 (N_3590,N_2867,N_787);
and U3591 (N_3591,N_351,N_615);
nor U3592 (N_3592,N_1335,N_1428);
xor U3593 (N_3593,N_2928,N_998);
nor U3594 (N_3594,N_478,N_1552);
and U3595 (N_3595,N_1834,N_27);
nor U3596 (N_3596,N_698,N_2075);
or U3597 (N_3597,N_2447,N_558);
nor U3598 (N_3598,N_2868,N_883);
nand U3599 (N_3599,N_116,N_606);
nand U3600 (N_3600,N_1419,N_707);
or U3601 (N_3601,N_2922,N_1230);
and U3602 (N_3602,N_897,N_946);
xnor U3603 (N_3603,N_2204,N_474);
or U3604 (N_3604,N_161,N_1246);
or U3605 (N_3605,N_419,N_1047);
nand U3606 (N_3606,N_309,N_2233);
nor U3607 (N_3607,N_2076,N_1115);
or U3608 (N_3608,N_531,N_6);
nand U3609 (N_3609,N_2053,N_2906);
or U3610 (N_3610,N_24,N_80);
nor U3611 (N_3611,N_1446,N_1761);
nand U3612 (N_3612,N_2125,N_183);
or U3613 (N_3613,N_2936,N_2741);
and U3614 (N_3614,N_1086,N_1669);
or U3615 (N_3615,N_2213,N_1973);
nand U3616 (N_3616,N_2651,N_1263);
and U3617 (N_3617,N_324,N_2458);
and U3618 (N_3618,N_2008,N_1096);
nor U3619 (N_3619,N_457,N_544);
nor U3620 (N_3620,N_2895,N_455);
and U3621 (N_3621,N_2503,N_81);
or U3622 (N_3622,N_577,N_1903);
or U3623 (N_3623,N_95,N_2036);
or U3624 (N_3624,N_2116,N_58);
and U3625 (N_3625,N_2110,N_2147);
nand U3626 (N_3626,N_830,N_1785);
or U3627 (N_3627,N_1048,N_1291);
or U3628 (N_3628,N_354,N_2774);
or U3629 (N_3629,N_1635,N_993);
nand U3630 (N_3630,N_2072,N_1662);
and U3631 (N_3631,N_2893,N_402);
nor U3632 (N_3632,N_384,N_167);
and U3633 (N_3633,N_2017,N_477);
nor U3634 (N_3634,N_896,N_2973);
or U3635 (N_3635,N_395,N_1596);
or U3636 (N_3636,N_955,N_507);
nor U3637 (N_3637,N_2218,N_2087);
nand U3638 (N_3638,N_2615,N_2117);
or U3639 (N_3639,N_2301,N_1688);
and U3640 (N_3640,N_230,N_1598);
xor U3641 (N_3641,N_572,N_718);
or U3642 (N_3642,N_976,N_1051);
nand U3643 (N_3643,N_119,N_2314);
nor U3644 (N_3644,N_2245,N_2991);
nor U3645 (N_3645,N_2171,N_1846);
and U3646 (N_3646,N_240,N_1681);
or U3647 (N_3647,N_2379,N_616);
nor U3648 (N_3648,N_2209,N_1166);
nand U3649 (N_3649,N_2237,N_2621);
or U3650 (N_3650,N_406,N_2812);
nand U3651 (N_3651,N_1044,N_1006);
nand U3652 (N_3652,N_2254,N_2378);
nand U3653 (N_3653,N_2980,N_462);
and U3654 (N_3654,N_1049,N_1163);
nand U3655 (N_3655,N_2427,N_2498);
nor U3656 (N_3656,N_1478,N_105);
and U3657 (N_3657,N_1463,N_1954);
nor U3658 (N_3658,N_379,N_1207);
nor U3659 (N_3659,N_889,N_412);
or U3660 (N_3660,N_2724,N_988);
or U3661 (N_3661,N_893,N_256);
nor U3662 (N_3662,N_2632,N_2066);
and U3663 (N_3663,N_1570,N_1288);
nand U3664 (N_3664,N_2765,N_608);
and U3665 (N_3665,N_1641,N_380);
or U3666 (N_3666,N_990,N_486);
or U3667 (N_3667,N_2141,N_629);
and U3668 (N_3668,N_1540,N_2009);
and U3669 (N_3669,N_1394,N_2816);
or U3670 (N_3670,N_500,N_595);
nor U3671 (N_3671,N_1399,N_1241);
or U3672 (N_3672,N_297,N_1753);
and U3673 (N_3673,N_1022,N_392);
nand U3674 (N_3674,N_2265,N_2896);
nor U3675 (N_3675,N_674,N_1710);
nand U3676 (N_3676,N_1531,N_2291);
and U3677 (N_3677,N_522,N_599);
nand U3678 (N_3678,N_175,N_31);
or U3679 (N_3679,N_276,N_268);
nand U3680 (N_3680,N_2289,N_333);
and U3681 (N_3681,N_2676,N_2940);
or U3682 (N_3682,N_188,N_2108);
nand U3683 (N_3683,N_1541,N_410);
nor U3684 (N_3684,N_2272,N_2618);
and U3685 (N_3685,N_2571,N_1777);
and U3686 (N_3686,N_2853,N_690);
and U3687 (N_3687,N_1581,N_1724);
and U3688 (N_3688,N_2511,N_2252);
or U3689 (N_3689,N_2354,N_2614);
or U3690 (N_3690,N_730,N_2264);
nand U3691 (N_3691,N_1901,N_1811);
xor U3692 (N_3692,N_85,N_941);
and U3693 (N_3693,N_936,N_1075);
or U3694 (N_3694,N_1632,N_709);
and U3695 (N_3695,N_2535,N_1855);
and U3696 (N_3696,N_2128,N_1928);
nand U3697 (N_3697,N_2335,N_921);
and U3698 (N_3698,N_1757,N_511);
nand U3699 (N_3699,N_1301,N_716);
nand U3700 (N_3700,N_1320,N_468);
nand U3701 (N_3701,N_1150,N_18);
nor U3702 (N_3702,N_2546,N_2332);
nand U3703 (N_3703,N_2686,N_1032);
nor U3704 (N_3704,N_315,N_114);
xor U3705 (N_3705,N_185,N_152);
and U3706 (N_3706,N_1701,N_1778);
nor U3707 (N_3707,N_258,N_766);
or U3708 (N_3708,N_1548,N_2478);
nand U3709 (N_3709,N_2446,N_453);
nand U3710 (N_3710,N_1887,N_2628);
or U3711 (N_3711,N_1964,N_177);
nor U3712 (N_3712,N_94,N_2520);
nand U3713 (N_3713,N_2093,N_2966);
or U3714 (N_3714,N_2943,N_1154);
nor U3715 (N_3715,N_2767,N_1173);
or U3716 (N_3716,N_2435,N_202);
nand U3717 (N_3717,N_646,N_2079);
nand U3718 (N_3718,N_1819,N_1221);
or U3719 (N_3719,N_1738,N_1076);
nand U3720 (N_3720,N_1865,N_50);
nor U3721 (N_3721,N_2500,N_2275);
or U3722 (N_3722,N_737,N_1752);
nand U3723 (N_3723,N_2026,N_1091);
and U3724 (N_3724,N_2607,N_1474);
or U3725 (N_3725,N_11,N_2879);
nor U3726 (N_3726,N_2493,N_2396);
or U3727 (N_3727,N_2205,N_1422);
xnor U3728 (N_3728,N_875,N_1253);
nand U3729 (N_3729,N_1929,N_2574);
nand U3730 (N_3730,N_1226,N_2663);
nand U3731 (N_3731,N_278,N_2838);
or U3732 (N_3732,N_2175,N_296);
or U3733 (N_3733,N_2658,N_816);
or U3734 (N_3734,N_827,N_1227);
nor U3735 (N_3735,N_2545,N_1203);
nand U3736 (N_3736,N_257,N_2227);
and U3737 (N_3737,N_2047,N_2187);
and U3738 (N_3738,N_2106,N_1356);
nor U3739 (N_3739,N_1692,N_1453);
or U3740 (N_3740,N_1921,N_2092);
or U3741 (N_3741,N_2392,N_2526);
or U3742 (N_3742,N_195,N_1600);
nand U3743 (N_3743,N_2718,N_56);
xor U3744 (N_3744,N_2206,N_2566);
and U3745 (N_3745,N_1916,N_350);
and U3746 (N_3746,N_717,N_2152);
nor U3747 (N_3747,N_944,N_2726);
nand U3748 (N_3748,N_2067,N_2874);
xor U3749 (N_3749,N_2689,N_2255);
xnor U3750 (N_3750,N_239,N_560);
nor U3751 (N_3751,N_1280,N_2962);
nor U3752 (N_3752,N_812,N_2841);
or U3753 (N_3753,N_159,N_1726);
or U3754 (N_3754,N_403,N_1818);
or U3755 (N_3755,N_2461,N_170);
nor U3756 (N_3756,N_1648,N_1741);
nand U3757 (N_3757,N_1010,N_2033);
nor U3758 (N_3758,N_460,N_635);
or U3759 (N_3759,N_1215,N_1398);
and U3760 (N_3760,N_1844,N_1443);
and U3761 (N_3761,N_1877,N_791);
nor U3762 (N_3762,N_458,N_1325);
and U3763 (N_3763,N_1338,N_982);
and U3764 (N_3764,N_625,N_2534);
and U3765 (N_3765,N_2537,N_2338);
or U3766 (N_3766,N_2519,N_850);
nor U3767 (N_3767,N_2756,N_2584);
nand U3768 (N_3768,N_779,N_2536);
and U3769 (N_3769,N_983,N_867);
or U3770 (N_3770,N_1482,N_1181);
nand U3771 (N_3771,N_1893,N_1127);
or U3772 (N_3772,N_2641,N_441);
and U3773 (N_3773,N_610,N_336);
and U3774 (N_3774,N_1158,N_414);
and U3775 (N_3775,N_339,N_1113);
and U3776 (N_3776,N_731,N_1774);
nand U3777 (N_3777,N_1539,N_2248);
xnor U3778 (N_3778,N_2330,N_2197);
and U3779 (N_3779,N_132,N_302);
nor U3780 (N_3780,N_493,N_272);
xnor U3781 (N_3781,N_2169,N_1345);
nor U3782 (N_3782,N_2417,N_497);
or U3783 (N_3783,N_2827,N_2052);
nor U3784 (N_3784,N_2681,N_2462);
nor U3785 (N_3785,N_47,N_2583);
nor U3786 (N_3786,N_1557,N_2163);
nand U3787 (N_3787,N_1837,N_1139);
nor U3788 (N_3788,N_46,N_1229);
nor U3789 (N_3789,N_358,N_2407);
and U3790 (N_3790,N_174,N_967);
nand U3791 (N_3791,N_1974,N_947);
nand U3792 (N_3792,N_2739,N_2802);
and U3793 (N_3793,N_2834,N_1816);
nand U3794 (N_3794,N_550,N_2049);
or U3795 (N_3795,N_1806,N_864);
nand U3796 (N_3796,N_2771,N_251);
nor U3797 (N_3797,N_439,N_1772);
nand U3798 (N_3798,N_2783,N_917);
nor U3799 (N_3799,N_2276,N_1193);
or U3800 (N_3800,N_1377,N_1742);
xnor U3801 (N_3801,N_735,N_1623);
nor U3802 (N_3802,N_700,N_4);
nor U3803 (N_3803,N_2367,N_2823);
nand U3804 (N_3804,N_61,N_634);
nor U3805 (N_3805,N_825,N_1309);
or U3806 (N_3806,N_287,N_515);
or U3807 (N_3807,N_1388,N_2740);
nor U3808 (N_3808,N_2341,N_2164);
nand U3809 (N_3809,N_465,N_2782);
or U3810 (N_3810,N_959,N_2271);
nand U3811 (N_3811,N_2469,N_2242);
nand U3812 (N_3812,N_1850,N_664);
and U3813 (N_3813,N_490,N_448);
nand U3814 (N_3814,N_1153,N_282);
nor U3815 (N_3815,N_1369,N_814);
nor U3816 (N_3816,N_2383,N_1536);
nor U3817 (N_3817,N_1485,N_214);
or U3818 (N_3818,N_2531,N_1052);
and U3819 (N_3819,N_1854,N_1155);
and U3820 (N_3820,N_2174,N_1733);
nand U3821 (N_3821,N_1238,N_2544);
and U3822 (N_3822,N_2191,N_1610);
and U3823 (N_3823,N_341,N_489);
nand U3824 (N_3824,N_1300,N_1068);
nand U3825 (N_3825,N_2492,N_1622);
nand U3826 (N_3826,N_400,N_2257);
and U3827 (N_3827,N_483,N_1416);
and U3828 (N_3828,N_356,N_2319);
nor U3829 (N_3829,N_1913,N_1187);
and U3830 (N_3830,N_2002,N_1389);
and U3831 (N_3831,N_432,N_1306);
and U3832 (N_3832,N_2824,N_426);
or U3833 (N_3833,N_1365,N_138);
nor U3834 (N_3834,N_2155,N_1167);
or U3835 (N_3835,N_631,N_2007);
and U3836 (N_3836,N_2892,N_2306);
and U3837 (N_3837,N_75,N_1589);
and U3838 (N_3838,N_648,N_345);
or U3839 (N_3839,N_789,N_2706);
nor U3840 (N_3840,N_2995,N_2165);
nand U3841 (N_3841,N_1358,N_1872);
nand U3842 (N_3842,N_363,N_1308);
nand U3843 (N_3843,N_1595,N_396);
or U3844 (N_3844,N_2236,N_1417);
or U3845 (N_3845,N_118,N_2964);
or U3846 (N_3846,N_882,N_2931);
nand U3847 (N_3847,N_956,N_847);
or U3848 (N_3848,N_1859,N_2561);
and U3849 (N_3849,N_780,N_2956);
nand U3850 (N_3850,N_413,N_2312);
and U3851 (N_3851,N_8,N_1251);
nand U3852 (N_3852,N_2277,N_1575);
xor U3853 (N_3853,N_2039,N_1658);
or U3854 (N_3854,N_1029,N_838);
nand U3855 (N_3855,N_224,N_2626);
nand U3856 (N_3856,N_2862,N_2398);
nand U3857 (N_3857,N_1523,N_1764);
nor U3858 (N_3858,N_666,N_2593);
nor U3859 (N_3859,N_714,N_557);
and U3860 (N_3860,N_2012,N_2114);
or U3861 (N_3861,N_137,N_401);
nand U3862 (N_3862,N_1072,N_1511);
or U3863 (N_3863,N_365,N_2678);
nor U3864 (N_3864,N_540,N_2515);
and U3865 (N_3865,N_1804,N_447);
and U3866 (N_3866,N_142,N_2670);
or U3867 (N_3867,N_1128,N_1450);
and U3868 (N_3868,N_2608,N_90);
nand U3869 (N_3869,N_2489,N_622);
nor U3870 (N_3870,N_21,N_2460);
and U3871 (N_3871,N_1939,N_1447);
or U3872 (N_3872,N_855,N_2484);
and U3873 (N_3873,N_2873,N_769);
nor U3874 (N_3874,N_1647,N_2154);
nor U3875 (N_3875,N_2,N_2316);
and U3876 (N_3876,N_1963,N_1437);
or U3877 (N_3877,N_1702,N_2405);
nand U3878 (N_3878,N_2364,N_2585);
and U3879 (N_3879,N_1955,N_2744);
nor U3880 (N_3880,N_1836,N_1411);
nor U3881 (N_3881,N_108,N_2877);
xor U3882 (N_3882,N_2884,N_1670);
nor U3883 (N_3883,N_1555,N_954);
and U3884 (N_3884,N_2731,N_2416);
nand U3885 (N_3885,N_1140,N_1384);
nor U3886 (N_3886,N_783,N_292);
and U3887 (N_3887,N_1860,N_828);
and U3888 (N_3888,N_1363,N_2453);
nand U3889 (N_3889,N_2284,N_1481);
nor U3890 (N_3890,N_1775,N_1179);
or U3891 (N_3891,N_2113,N_676);
nand U3892 (N_3892,N_1034,N_1472);
or U3893 (N_3893,N_805,N_839);
or U3894 (N_3894,N_2302,N_344);
and U3895 (N_3895,N_906,N_1651);
nor U3896 (N_3896,N_1902,N_1081);
or U3897 (N_3897,N_1313,N_1110);
nor U3898 (N_3898,N_2675,N_2455);
and U3899 (N_3899,N_2852,N_461);
nor U3900 (N_3900,N_2622,N_1631);
nand U3901 (N_3901,N_752,N_775);
or U3902 (N_3902,N_1751,N_429);
nand U3903 (N_3903,N_1024,N_563);
and U3904 (N_3904,N_763,N_2826);
nor U3905 (N_3905,N_2270,N_364);
and U3906 (N_3906,N_2555,N_1245);
or U3907 (N_3907,N_308,N_1162);
or U3908 (N_3908,N_2244,N_1461);
or U3909 (N_3909,N_685,N_1948);
nand U3910 (N_3910,N_1012,N_262);
or U3911 (N_3911,N_809,N_237);
nand U3912 (N_3912,N_2071,N_3);
and U3913 (N_3913,N_2887,N_905);
or U3914 (N_3914,N_288,N_2097);
or U3915 (N_3915,N_2126,N_1682);
nor U3916 (N_3916,N_2479,N_1452);
nor U3917 (N_3917,N_1795,N_699);
nor U3918 (N_3918,N_303,N_1218);
nand U3919 (N_3919,N_1984,N_788);
or U3920 (N_3920,N_686,N_2647);
or U3921 (N_3921,N_2755,N_2168);
and U3922 (N_3922,N_806,N_1817);
nand U3923 (N_3923,N_2334,N_653);
and U3924 (N_3924,N_556,N_2742);
and U3925 (N_3925,N_863,N_1359);
nand U3926 (N_3926,N_1252,N_995);
or U3927 (N_3927,N_2073,N_192);
nand U3928 (N_3928,N_2210,N_797);
or U3929 (N_3929,N_1519,N_1462);
or U3930 (N_3930,N_1427,N_2692);
nor U3931 (N_3931,N_340,N_1747);
nand U3932 (N_3932,N_2241,N_1094);
or U3933 (N_3933,N_2062,N_2997);
and U3934 (N_3934,N_15,N_2057);
nand U3935 (N_3935,N_91,N_1375);
or U3936 (N_3936,N_1114,N_1334);
nor U3937 (N_3937,N_1676,N_1908);
nand U3938 (N_3938,N_691,N_740);
nor U3939 (N_3939,N_2902,N_673);
or U3940 (N_3940,N_314,N_2480);
nand U3941 (N_3941,N_2133,N_2926);
nor U3942 (N_3942,N_618,N_2130);
nor U3943 (N_3943,N_209,N_2342);
nor U3944 (N_3944,N_2504,N_101);
nor U3945 (N_3945,N_588,N_25);
nor U3946 (N_3946,N_854,N_1814);
nor U3947 (N_3947,N_1739,N_376);
and U3948 (N_3948,N_2969,N_433);
or U3949 (N_3949,N_2350,N_1445);
or U3950 (N_3950,N_221,N_199);
and U3951 (N_3951,N_2558,N_2596);
or U3952 (N_3952,N_374,N_2903);
nand U3953 (N_3953,N_2353,N_1591);
or U3954 (N_3954,N_2020,N_382);
nand U3955 (N_3955,N_2682,N_217);
xnor U3956 (N_3956,N_2532,N_2979);
nand U3957 (N_3957,N_2094,N_2778);
or U3958 (N_3958,N_1323,N_1572);
and U3959 (N_3959,N_2784,N_1942);
or U3960 (N_3960,N_2732,N_1426);
or U3961 (N_3961,N_1927,N_169);
and U3962 (N_3962,N_232,N_212);
nor U3963 (N_3963,N_1055,N_1442);
and U3964 (N_3964,N_1853,N_494);
xor U3965 (N_3965,N_1840,N_135);
or U3966 (N_3966,N_1003,N_2156);
nor U3967 (N_3967,N_84,N_1993);
and U3968 (N_3968,N_2089,N_2192);
nor U3969 (N_3969,N_2115,N_388);
nand U3970 (N_3970,N_662,N_456);
and U3971 (N_3971,N_1528,N_1406);
nand U3972 (N_3972,N_2065,N_2011);
and U3973 (N_3973,N_2792,N_843);
nor U3974 (N_3974,N_1297,N_2318);
or U3975 (N_3975,N_1551,N_2512);
nand U3976 (N_3976,N_293,N_2238);
and U3977 (N_3977,N_2278,N_1674);
nor U3978 (N_3978,N_2573,N_1473);
and U3979 (N_3979,N_1980,N_271);
nor U3980 (N_3980,N_2746,N_1403);
or U3981 (N_3981,N_2438,N_1026);
and U3982 (N_3982,N_965,N_2028);
xnor U3983 (N_3983,N_1799,N_472);
or U3984 (N_3984,N_1479,N_1078);
or U3985 (N_3985,N_1302,N_1743);
nor U3986 (N_3986,N_2509,N_2938);
or U3987 (N_3987,N_857,N_343);
or U3988 (N_3988,N_2333,N_1706);
nand U3989 (N_3989,N_2311,N_1151);
or U3990 (N_3990,N_1244,N_980);
nand U3991 (N_3991,N_2955,N_2635);
or U3992 (N_3992,N_2705,N_811);
nor U3993 (N_3993,N_2157,N_469);
nor U3994 (N_3994,N_590,N_2127);
or U3995 (N_3995,N_2176,N_1318);
and U3996 (N_3996,N_749,N_2222);
and U3997 (N_3997,N_2660,N_104);
and U3998 (N_3998,N_1945,N_623);
xor U3999 (N_3999,N_1508,N_1566);
nand U4000 (N_4000,N_860,N_2648);
nor U4001 (N_4001,N_1549,N_2223);
nor U4002 (N_4002,N_930,N_1961);
and U4003 (N_4003,N_491,N_2989);
and U4004 (N_4004,N_294,N_147);
nor U4005 (N_4005,N_1236,N_2611);
nor U4006 (N_4006,N_2436,N_51);
or U4007 (N_4007,N_2559,N_145);
nand U4008 (N_4008,N_669,N_166);
nor U4009 (N_4009,N_328,N_69);
nand U4010 (N_4010,N_1947,N_1107);
and U4011 (N_4011,N_1824,N_77);
and U4012 (N_4012,N_1148,N_1451);
and U4013 (N_4013,N_1613,N_1526);
xor U4014 (N_4014,N_1059,N_2260);
nor U4015 (N_4015,N_2279,N_2086);
nor U4016 (N_4016,N_2897,N_1343);
and U4017 (N_4017,N_2959,N_245);
nor U4018 (N_4018,N_1407,N_2917);
and U4019 (N_4019,N_848,N_650);
nand U4020 (N_4020,N_2656,N_1856);
nor U4021 (N_4021,N_1262,N_2506);
nor U4022 (N_4022,N_2604,N_878);
and U4023 (N_4023,N_2594,N_1975);
and U4024 (N_4024,N_244,N_2796);
nor U4025 (N_4025,N_143,N_2363);
and U4026 (N_4026,N_1382,N_1994);
nand U4027 (N_4027,N_1168,N_1821);
nand U4028 (N_4028,N_1304,N_1569);
nor U4029 (N_4029,N_200,N_210);
nand U4030 (N_4030,N_892,N_422);
nand U4031 (N_4031,N_2483,N_1886);
or U4032 (N_4032,N_1556,N_2280);
nor U4033 (N_4033,N_2400,N_1671);
nand U4034 (N_4034,N_667,N_2038);
nand U4035 (N_4035,N_592,N_1311);
nor U4036 (N_4036,N_2582,N_501);
nand U4037 (N_4037,N_2655,N_2870);
nand U4038 (N_4038,N_1769,N_1191);
nor U4039 (N_4039,N_1561,N_2456);
and U4040 (N_4040,N_745,N_1949);
nand U4041 (N_4041,N_2069,N_1534);
xor U4042 (N_4042,N_1093,N_1161);
nand U4043 (N_4043,N_2476,N_1275);
and U4044 (N_4044,N_107,N_2781);
nor U4045 (N_4045,N_1111,N_1815);
or U4046 (N_4046,N_267,N_2251);
nor U4047 (N_4047,N_2294,N_596);
or U4048 (N_4048,N_762,N_411);
nand U4049 (N_4049,N_948,N_2941);
or U4050 (N_4050,N_42,N_2414);
nor U4051 (N_4051,N_1957,N_1123);
or U4052 (N_4052,N_2173,N_2505);
or U4053 (N_4053,N_1257,N_2482);
nand U4054 (N_4054,N_2913,N_1813);
nor U4055 (N_4055,N_1315,N_2748);
and U4056 (N_4056,N_842,N_2323);
or U4057 (N_4057,N_894,N_2576);
xnor U4058 (N_4058,N_2736,N_928);
and U4059 (N_4059,N_1626,N_2698);
and U4060 (N_4060,N_594,N_2200);
nor U4061 (N_4061,N_417,N_1402);
nor U4062 (N_4062,N_924,N_1530);
nor U4063 (N_4063,N_2673,N_1845);
and U4064 (N_4064,N_1553,N_663);
or U4065 (N_4065,N_121,N_2612);
and U4066 (N_4066,N_312,N_2552);
nor U4067 (N_4067,N_2214,N_2865);
nor U4068 (N_4068,N_654,N_1862);
or U4069 (N_4069,N_887,N_1287);
nor U4070 (N_4070,N_2220,N_1493);
and U4071 (N_4071,N_2977,N_2766);
or U4072 (N_4072,N_2667,N_2990);
nor U4073 (N_4073,N_2211,N_1387);
or U4074 (N_4074,N_54,N_583);
nand U4075 (N_4075,N_817,N_1981);
nand U4076 (N_4076,N_2188,N_1316);
nor U4077 (N_4077,N_2715,N_1516);
nor U4078 (N_4078,N_1385,N_2661);
and U4079 (N_4079,N_1097,N_2738);
and U4080 (N_4080,N_1020,N_39);
nand U4081 (N_4081,N_1319,N_2471);
or U4082 (N_4082,N_2262,N_2470);
nand U4083 (N_4083,N_601,N_2624);
xor U4084 (N_4084,N_1780,N_2983);
and U4085 (N_4085,N_1322,N_2450);
and U4086 (N_4086,N_1996,N_2875);
nor U4087 (N_4087,N_1567,N_1361);
nand U4088 (N_4088,N_1143,N_2685);
and U4089 (N_4089,N_2577,N_656);
nand U4090 (N_4090,N_960,N_1222);
and U4091 (N_4091,N_360,N_1728);
or U4092 (N_4092,N_1002,N_346);
nand U4093 (N_4093,N_2296,N_994);
nor U4094 (N_4094,N_566,N_140);
nor U4095 (N_4095,N_1436,N_888);
nor U4096 (N_4096,N_2832,N_1910);
and U4097 (N_4097,N_2568,N_301);
or U4098 (N_4098,N_2775,N_1533);
nor U4099 (N_4099,N_1878,N_2331);
and U4100 (N_4100,N_626,N_2579);
nand U4101 (N_4101,N_2734,N_2080);
nor U4102 (N_4102,N_300,N_2477);
and U4103 (N_4103,N_719,N_2372);
nor U4104 (N_4104,N_1124,N_1444);
and U4105 (N_4105,N_1930,N_919);
or U4106 (N_4106,N_1237,N_78);
nand U4107 (N_4107,N_1909,N_2134);
or U4108 (N_4108,N_2592,N_1330);
nor U4109 (N_4109,N_503,N_390);
or U4110 (N_4110,N_1861,N_2543);
nand U4111 (N_4111,N_2729,N_2587);
xor U4112 (N_4112,N_254,N_1283);
nand U4113 (N_4113,N_2605,N_968);
or U4114 (N_4114,N_2368,N_756);
and U4115 (N_4115,N_1694,N_2904);
or U4116 (N_4116,N_2701,N_1117);
and U4117 (N_4117,N_1578,N_1789);
nand U4118 (N_4118,N_1543,N_778);
xnor U4119 (N_4119,N_1920,N_1639);
or U4120 (N_4120,N_1685,N_807);
nand U4121 (N_4121,N_1025,N_574);
nand U4122 (N_4122,N_2224,N_2074);
nand U4123 (N_4123,N_2411,N_2420);
nand U4124 (N_4124,N_2101,N_2010);
nand U4125 (N_4125,N_1636,N_1213);
or U4126 (N_4126,N_2634,N_2586);
and U4127 (N_4127,N_970,N_1517);
or U4128 (N_4128,N_1276,N_1971);
or U4129 (N_4129,N_1587,N_516);
nor U4130 (N_4130,N_950,N_1897);
and U4131 (N_4131,N_2412,N_2431);
nor U4132 (N_4132,N_2787,N_2064);
and U4133 (N_4133,N_1985,N_464);
nor U4134 (N_4134,N_2804,N_2150);
nand U4135 (N_4135,N_1347,N_466);
or U4136 (N_4136,N_836,N_1982);
or U4137 (N_4137,N_496,N_1746);
or U4138 (N_4138,N_2737,N_2820);
or U4139 (N_4139,N_1500,N_45);
nand U4140 (N_4140,N_767,N_1748);
nor U4141 (N_4141,N_391,N_1209);
or U4142 (N_4142,N_1067,N_2170);
and U4143 (N_4143,N_2525,N_1256);
nand U4144 (N_4144,N_538,N_49);
nand U4145 (N_4145,N_377,N_1643);
nand U4146 (N_4146,N_2601,N_1217);
or U4147 (N_4147,N_852,N_695);
or U4148 (N_4148,N_445,N_416);
or U4149 (N_4149,N_86,N_1801);
nand U4150 (N_4150,N_661,N_1085);
nor U4151 (N_4151,N_1386,N_361);
nor U4152 (N_4152,N_1225,N_2388);
or U4153 (N_4153,N_321,N_1791);
or U4154 (N_4154,N_2502,N_2001);
nand U4155 (N_4155,N_2773,N_1654);
and U4156 (N_4156,N_1284,N_1360);
or U4157 (N_4157,N_1346,N_1585);
nor U4158 (N_4158,N_2195,N_2190);
and U4159 (N_4159,N_418,N_2861);
and U4160 (N_4160,N_776,N_171);
or U4161 (N_4161,N_1307,N_1342);
nand U4162 (N_4162,N_568,N_1807);
nand U4163 (N_4163,N_1423,N_920);
or U4164 (N_4164,N_916,N_1722);
nand U4165 (N_4165,N_680,N_1483);
nand U4166 (N_4166,N_2809,N_1546);
nor U4167 (N_4167,N_911,N_2944);
nand U4168 (N_4168,N_764,N_2025);
or U4169 (N_4169,N_5,N_1200);
nor U4170 (N_4170,N_2538,N_505);
and U4171 (N_4171,N_1392,N_1766);
or U4172 (N_4172,N_1677,N_520);
or U4173 (N_4173,N_1802,N_305);
or U4174 (N_4174,N_1017,N_829);
nor U4175 (N_4175,N_139,N_359);
nor U4176 (N_4176,N_349,N_2145);
nand U4177 (N_4177,N_2954,N_2610);
and U4178 (N_4178,N_2937,N_498);
nand U4179 (N_4179,N_543,N_2984);
nand U4180 (N_4180,N_512,N_2993);
and U4181 (N_4181,N_2317,N_1620);
or U4182 (N_4182,N_499,N_2721);
and U4183 (N_4183,N_1664,N_1448);
nand U4184 (N_4184,N_1298,N_459);
and U4185 (N_4185,N_2315,N_1937);
nor U4186 (N_4186,N_1653,N_2040);
and U4187 (N_4187,N_913,N_2023);
nand U4188 (N_4188,N_1841,N_1991);
and U4189 (N_4189,N_678,N_1874);
or U4190 (N_4190,N_567,N_2806);
and U4191 (N_4191,N_1255,N_1721);
or U4192 (N_4192,N_1425,N_1271);
and U4193 (N_4193,N_473,N_832);
and U4194 (N_4194,N_1729,N_44);
nand U4195 (N_4195,N_1132,N_748);
nand U4196 (N_4196,N_191,N_785);
nor U4197 (N_4197,N_912,N_2652);
or U4198 (N_4198,N_637,N_2844);
nor U4199 (N_4199,N_2377,N_2857);
nor U4200 (N_4200,N_331,N_1509);
nand U4201 (N_4201,N_750,N_1952);
nor U4202 (N_4202,N_1934,N_92);
nor U4203 (N_4203,N_1102,N_311);
and U4204 (N_4204,N_1989,N_660);
and U4205 (N_4205,N_2297,N_2693);
or U4206 (N_4206,N_2924,N_208);
xnor U4207 (N_4207,N_1735,N_10);
nand U4208 (N_4208,N_1756,N_541);
xor U4209 (N_4209,N_2563,N_1126);
nor U4210 (N_4210,N_290,N_2182);
and U4211 (N_4211,N_337,N_1189);
nor U4212 (N_4212,N_1100,N_732);
or U4213 (N_4213,N_1953,N_2722);
or U4214 (N_4214,N_1019,N_2863);
and U4215 (N_4215,N_1488,N_495);
or U4216 (N_4216,N_587,N_1922);
nor U4217 (N_4217,N_1305,N_2487);
or U4218 (N_4218,N_768,N_2948);
nor U4219 (N_4219,N_2749,N_1054);
or U4220 (N_4220,N_1593,N_2790);
nor U4221 (N_4221,N_481,N_1605);
or U4222 (N_4222,N_689,N_804);
and U4223 (N_4223,N_2328,N_603);
and U4224 (N_4224,N_249,N_1134);
nand U4225 (N_4225,N_1071,N_2441);
nor U4226 (N_4226,N_932,N_1372);
or U4227 (N_4227,N_1573,N_1468);
and U4228 (N_4228,N_840,N_551);
and U4229 (N_4229,N_2207,N_553);
nand U4230 (N_4230,N_1650,N_2389);
nor U4231 (N_4231,N_1295,N_2762);
nand U4232 (N_4232,N_2112,N_168);
and U4233 (N_4233,N_870,N_2533);
nor U4234 (N_4234,N_758,N_881);
or U4235 (N_4235,N_2982,N_1232);
and U4236 (N_4236,N_786,N_677);
and U4237 (N_4237,N_2952,N_2178);
and U4238 (N_4238,N_571,N_1206);
nor U4239 (N_4239,N_1889,N_1510);
and U4240 (N_4240,N_879,N_2030);
nand U4241 (N_4241,N_2669,N_1135);
nor U4242 (N_4242,N_1890,N_1866);
and U4243 (N_4243,N_2961,N_2798);
or U4244 (N_4244,N_963,N_1354);
nor U4245 (N_4245,N_298,N_2082);
nor U4246 (N_4246,N_19,N_1210);
or U4247 (N_4247,N_2971,N_2142);
nand U4248 (N_4248,N_1033,N_628);
or U4249 (N_4249,N_463,N_2539);
and U4250 (N_4250,N_2343,N_549);
nor U4251 (N_4251,N_876,N_2339);
nand U4252 (N_4252,N_1057,N_2650);
nor U4253 (N_4253,N_1704,N_1542);
or U4254 (N_4254,N_176,N_2898);
or U4255 (N_4255,N_2643,N_564);
nor U4256 (N_4256,N_2365,N_642);
and U4257 (N_4257,N_559,N_1199);
nand U4258 (N_4258,N_2299,N_1267);
or U4259 (N_4259,N_238,N_1409);
nor U4260 (N_4260,N_1972,N_1580);
nor U4261 (N_4261,N_1223,N_2444);
and U4262 (N_4262,N_33,N_317);
nor U4263 (N_4263,N_1788,N_2258);
or U4264 (N_4264,N_259,N_330);
and U4265 (N_4265,N_1699,N_362);
and U4266 (N_4266,N_1317,N_103);
or U4267 (N_4267,N_1031,N_279);
or U4268 (N_4268,N_682,N_2923);
nand U4269 (N_4269,N_679,N_1331);
and U4270 (N_4270,N_2084,N_845);
nand U4271 (N_4271,N_1828,N_1503);
nand U4272 (N_4272,N_1441,N_452);
and U4273 (N_4273,N_1796,N_2391);
or U4274 (N_4274,N_1087,N_1634);
or U4275 (N_4275,N_1250,N_1977);
and U4276 (N_4276,N_2394,N_1612);
and U4277 (N_4277,N_2588,N_1944);
or U4278 (N_4278,N_724,N_1492);
nor U4279 (N_4279,N_2958,N_2286);
and U4280 (N_4280,N_1070,N_521);
and U4281 (N_4281,N_123,N_2730);
or U4282 (N_4282,N_575,N_2858);
and U4283 (N_4283,N_2266,N_886);
nor U4284 (N_4284,N_1090,N_2697);
nor U4285 (N_4285,N_971,N_640);
and U4286 (N_4286,N_2599,N_32);
nand U4287 (N_4287,N_133,N_1608);
and U4288 (N_4288,N_1652,N_504);
or U4289 (N_4289,N_1374,N_299);
nor U4290 (N_4290,N_295,N_2821);
nand U4291 (N_4291,N_1810,N_2633);
and U4292 (N_4292,N_765,N_1604);
nor U4293 (N_4293,N_265,N_1045);
nand U4294 (N_4294,N_636,N_1104);
and U4295 (N_4295,N_110,N_96);
and U4296 (N_4296,N_569,N_2166);
nand U4297 (N_4297,N_1709,N_962);
nand U4298 (N_4298,N_818,N_2750);
nand U4299 (N_4299,N_348,N_792);
nand U4300 (N_4300,N_2562,N_826);
and U4301 (N_4301,N_1152,N_2779);
nor U4302 (N_4302,N_23,N_687);
nor U4303 (N_4303,N_907,N_2439);
nor U4304 (N_4304,N_1584,N_1876);
and U4305 (N_4305,N_1274,N_2759);
nand U4306 (N_4306,N_1352,N_1101);
nand U4307 (N_4307,N_2799,N_1413);
nor U4308 (N_4308,N_2358,N_2415);
nand U4309 (N_4309,N_2795,N_1695);
or U4310 (N_4310,N_306,N_2890);
nor U4311 (N_4311,N_1852,N_1960);
nor U4312 (N_4312,N_2473,N_729);
and U4313 (N_4313,N_1538,N_307);
nand U4314 (N_4314,N_1400,N_1686);
nand U4315 (N_4315,N_1220,N_1784);
or U4316 (N_4316,N_157,N_1754);
or U4317 (N_4317,N_2517,N_2996);
or U4318 (N_4318,N_2747,N_378);
or U4319 (N_4319,N_2899,N_1967);
nand U4320 (N_4320,N_2508,N_0);
nor U4321 (N_4321,N_2805,N_1645);
or U4322 (N_4322,N_1208,N_979);
nor U4323 (N_4323,N_1286,N_2878);
nand U4324 (N_4324,N_206,N_1979);
or U4325 (N_4325,N_2836,N_203);
and U4326 (N_4326,N_1264,N_1505);
nand U4327 (N_4327,N_1736,N_705);
and U4328 (N_4328,N_1116,N_1145);
nor U4329 (N_4329,N_1638,N_332);
nand U4330 (N_4330,N_533,N_2104);
xor U4331 (N_4331,N_1367,N_184);
or U4332 (N_4332,N_1204,N_173);
or U4333 (N_4333,N_2054,N_1355);
nor U4334 (N_4334,N_30,N_1808);
or U4335 (N_4335,N_2369,N_313);
and U4336 (N_4336,N_444,N_273);
and U4337 (N_4337,N_2137,N_1999);
nand U4338 (N_4338,N_1884,N_1744);
and U4339 (N_4339,N_2662,N_2032);
nor U4340 (N_4340,N_1649,N_1700);
or U4341 (N_4341,N_428,N_2714);
nor U4342 (N_4342,N_74,N_2309);
nand U4343 (N_4343,N_1869,N_2422);
or U4344 (N_4344,N_1293,N_532);
nor U4345 (N_4345,N_1970,N_381);
or U4346 (N_4346,N_1762,N_2234);
and U4347 (N_4347,N_1576,N_1962);
and U4348 (N_4348,N_1289,N_895);
nand U4349 (N_4349,N_1395,N_111);
or U4350 (N_4350,N_2843,N_861);
or U4351 (N_4351,N_2463,N_899);
nand U4352 (N_4352,N_813,N_1998);
or U4353 (N_4353,N_2129,N_269);
nand U4354 (N_4354,N_2404,N_605);
nor U4355 (N_4355,N_659,N_2376);
or U4356 (N_4356,N_1684,N_1185);
nor U4357 (N_4357,N_697,N_903);
or U4358 (N_4358,N_1083,N_798);
xnor U4359 (N_4359,N_1770,N_275);
nand U4360 (N_4360,N_2491,N_1362);
or U4361 (N_4361,N_2186,N_641);
nand U4362 (N_4362,N_2719,N_2711);
or U4363 (N_4363,N_193,N_2687);
nand U4364 (N_4364,N_2041,N_1932);
nand U4365 (N_4365,N_2355,N_1292);
nor U4366 (N_4366,N_1931,N_722);
or U4367 (N_4367,N_1172,N_1249);
and U4368 (N_4368,N_2668,N_2313);
and U4369 (N_4369,N_2055,N_338);
or U4370 (N_4370,N_2226,N_66);
nand U4371 (N_4371,N_367,N_2900);
nor U4372 (N_4372,N_774,N_487);
or U4373 (N_4373,N_260,N_1588);
nand U4374 (N_4374,N_442,N_725);
xor U4375 (N_4375,N_2199,N_2327);
nor U4376 (N_4376,N_2521,N_2839);
nand U4377 (N_4377,N_366,N_2124);
or U4378 (N_4378,N_2111,N_274);
and U4379 (N_4379,N_1640,N_2292);
nand U4380 (N_4380,N_207,N_2428);
nand U4381 (N_4381,N_1672,N_1353);
nor U4382 (N_4382,N_1601,N_548);
xnor U4383 (N_4383,N_1765,N_2625);
nor U4384 (N_4384,N_793,N_2247);
and U4385 (N_4385,N_1005,N_1660);
and U4386 (N_4386,N_1936,N_1373);
nand U4387 (N_4387,N_2619,N_144);
nor U4388 (N_4388,N_1,N_2551);
nor U4389 (N_4389,N_1624,N_614);
and U4390 (N_4390,N_926,N_1621);
and U4391 (N_4391,N_14,N_822);
nand U4392 (N_4392,N_1060,N_2542);
nand U4393 (N_4393,N_1470,N_1563);
nor U4394 (N_4394,N_233,N_713);
nor U4395 (N_4395,N_1666,N_2911);
or U4396 (N_4396,N_2287,N_106);
or U4397 (N_4397,N_2406,N_2743);
or U4398 (N_4398,N_2243,N_189);
and U4399 (N_4399,N_821,N_984);
or U4400 (N_4400,N_996,N_1157);
nor U4401 (N_4401,N_1615,N_1583);
nand U4402 (N_4402,N_197,N_1661);
nor U4403 (N_4403,N_2710,N_443);
nor U4404 (N_4404,N_1614,N_194);
or U4405 (N_4405,N_352,N_1108);
and U4406 (N_4406,N_1357,N_1164);
nor U4407 (N_4407,N_1763,N_624);
and U4408 (N_4408,N_2429,N_2916);
nor U4409 (N_4409,N_2776,N_2981);
or U4410 (N_4410,N_1408,N_102);
nand U4411 (N_4411,N_2249,N_2018);
or U4412 (N_4412,N_2516,N_2578);
and U4413 (N_4413,N_2122,N_681);
and U4414 (N_4414,N_1851,N_1714);
and U4415 (N_4415,N_773,N_2976);
xor U4416 (N_4416,N_2443,N_2153);
nand U4417 (N_4417,N_1894,N_2123);
or U4418 (N_4418,N_1607,N_508);
or U4419 (N_4419,N_772,N_2045);
nor U4420 (N_4420,N_1364,N_1718);
and U4421 (N_4421,N_593,N_1832);
or U4422 (N_4422,N_710,N_2707);
nand U4423 (N_4423,N_1314,N_187);
nand U4424 (N_4424,N_1781,N_2942);
nor U4425 (N_4425,N_506,N_2468);
and U4426 (N_4426,N_819,N_2659);
nor U4427 (N_4427,N_323,N_2700);
nand U4428 (N_4428,N_856,N_1668);
xor U4429 (N_4429,N_859,N_2307);
and U4430 (N_4430,N_2216,N_2881);
nand U4431 (N_4431,N_1239,N_2642);
nand U4432 (N_4432,N_1201,N_2305);
and U4433 (N_4433,N_2709,N_942);
nand U4434 (N_4434,N_2003,N_34);
and U4435 (N_4435,N_1130,N_1768);
or U4436 (N_4436,N_1707,N_1329);
and U4437 (N_4437,N_1644,N_2849);
or U4438 (N_4438,N_1732,N_940);
nand U4439 (N_4439,N_872,N_1809);
nand U4440 (N_4440,N_250,N_1391);
nand U4441 (N_4441,N_2845,N_1368);
nand U4442 (N_4442,N_1205,N_815);
nor U4443 (N_4443,N_2819,N_1258);
nor U4444 (N_4444,N_2518,N_1737);
or U4445 (N_4445,N_1188,N_2814);
nor U4446 (N_4446,N_694,N_229);
and U4447 (N_4447,N_2554,N_720);
or U4448 (N_4448,N_837,N_1013);
nand U4449 (N_4449,N_55,N_2757);
or U4450 (N_4450,N_2051,N_2360);
nand U4451 (N_4451,N_747,N_1797);
and U4452 (N_4452,N_1545,N_218);
and U4453 (N_4453,N_1000,N_1995);
and U4454 (N_4454,N_582,N_1571);
and U4455 (N_4455,N_1324,N_1279);
nand U4456 (N_4456,N_2847,N_943);
and U4457 (N_4457,N_885,N_2232);
or U4458 (N_4458,N_627,N_2690);
nand U4459 (N_4459,N_405,N_329);
nand U4460 (N_4460,N_2430,N_2246);
and U4461 (N_4461,N_977,N_1224);
nand U4462 (N_4462,N_759,N_2346);
nand U4463 (N_4463,N_1433,N_285);
or U4464 (N_4464,N_1703,N_2131);
nand U4465 (N_4465,N_2399,N_1690);
nand U4466 (N_4466,N_1455,N_2998);
or U4467 (N_4467,N_619,N_2393);
nand U4468 (N_4468,N_1532,N_2986);
nand U4469 (N_4469,N_2680,N_1719);
nand U4470 (N_4470,N_2522,N_820);
and U4471 (N_4471,N_862,N_2225);
nor U4472 (N_4472,N_580,N_1131);
and U4473 (N_4473,N_1826,N_1659);
nor U4474 (N_4474,N_1842,N_2992);
and U4475 (N_4475,N_1918,N_1627);
and U4476 (N_4476,N_2352,N_180);
nand U4477 (N_4477,N_28,N_2375);
nand U4478 (N_4478,N_801,N_591);
and U4479 (N_4479,N_2974,N_1371);
nor U4480 (N_4480,N_1270,N_1219);
nand U4481 (N_4481,N_2638,N_1282);
nor U4482 (N_4482,N_2696,N_632);
and U4483 (N_4483,N_1458,N_398);
or U4484 (N_4484,N_1466,N_2850);
xnor U4485 (N_4485,N_1858,N_1606);
and U4486 (N_4486,N_799,N_1857);
nor U4487 (N_4487,N_130,N_1348);
nor U4488 (N_4488,N_1915,N_73);
or U4489 (N_4489,N_1496,N_2501);
nor U4490 (N_4490,N_1120,N_652);
and U4491 (N_4491,N_1165,N_1535);
and U4492 (N_4492,N_479,N_545);
or U4493 (N_4493,N_1745,N_514);
nor U4494 (N_4494,N_2442,N_2575);
nand U4495 (N_4495,N_611,N_2326);
and U4496 (N_4496,N_643,N_2356);
or U4497 (N_4497,N_1169,N_2639);
and U4498 (N_4498,N_1501,N_2646);
and U4499 (N_4499,N_1951,N_1216);
nand U4500 (N_4500,N_1161,N_1440);
nand U4501 (N_4501,N_2786,N_699);
and U4502 (N_4502,N_2166,N_2069);
nor U4503 (N_4503,N_1269,N_1645);
or U4504 (N_4504,N_1753,N_850);
nand U4505 (N_4505,N_853,N_293);
or U4506 (N_4506,N_2868,N_1633);
xnor U4507 (N_4507,N_1117,N_25);
and U4508 (N_4508,N_2156,N_1935);
or U4509 (N_4509,N_2359,N_2226);
xor U4510 (N_4510,N_2127,N_948);
or U4511 (N_4511,N_1242,N_1894);
nand U4512 (N_4512,N_2223,N_429);
nor U4513 (N_4513,N_1548,N_2572);
or U4514 (N_4514,N_1577,N_2277);
or U4515 (N_4515,N_836,N_1537);
nor U4516 (N_4516,N_430,N_100);
nor U4517 (N_4517,N_1177,N_251);
nand U4518 (N_4518,N_2438,N_1489);
or U4519 (N_4519,N_5,N_358);
or U4520 (N_4520,N_2493,N_966);
nand U4521 (N_4521,N_784,N_304);
xor U4522 (N_4522,N_2227,N_2630);
or U4523 (N_4523,N_1328,N_481);
nand U4524 (N_4524,N_2202,N_2727);
or U4525 (N_4525,N_2216,N_1871);
nor U4526 (N_4526,N_861,N_2842);
or U4527 (N_4527,N_2008,N_1733);
and U4528 (N_4528,N_268,N_140);
and U4529 (N_4529,N_1895,N_2484);
nand U4530 (N_4530,N_1829,N_1846);
and U4531 (N_4531,N_1814,N_1383);
or U4532 (N_4532,N_1515,N_2659);
nor U4533 (N_4533,N_2819,N_189);
nand U4534 (N_4534,N_2186,N_169);
nand U4535 (N_4535,N_2389,N_455);
and U4536 (N_4536,N_2257,N_1431);
nand U4537 (N_4537,N_1007,N_1468);
nor U4538 (N_4538,N_2495,N_1765);
or U4539 (N_4539,N_1926,N_2727);
or U4540 (N_4540,N_2734,N_2018);
nand U4541 (N_4541,N_747,N_728);
or U4542 (N_4542,N_1640,N_2433);
and U4543 (N_4543,N_1819,N_444);
nand U4544 (N_4544,N_1424,N_1651);
nor U4545 (N_4545,N_1626,N_1417);
and U4546 (N_4546,N_1530,N_1335);
or U4547 (N_4547,N_2725,N_2120);
nor U4548 (N_4548,N_2522,N_669);
and U4549 (N_4549,N_636,N_1423);
nor U4550 (N_4550,N_2599,N_421);
nor U4551 (N_4551,N_357,N_169);
nand U4552 (N_4552,N_881,N_2338);
or U4553 (N_4553,N_2701,N_1307);
or U4554 (N_4554,N_1668,N_178);
nand U4555 (N_4555,N_1016,N_373);
and U4556 (N_4556,N_2027,N_1957);
nor U4557 (N_4557,N_480,N_1635);
nor U4558 (N_4558,N_1299,N_2119);
nand U4559 (N_4559,N_1267,N_2278);
or U4560 (N_4560,N_2360,N_1216);
nor U4561 (N_4561,N_57,N_2271);
and U4562 (N_4562,N_627,N_934);
nand U4563 (N_4563,N_1663,N_362);
nand U4564 (N_4564,N_1950,N_621);
nor U4565 (N_4565,N_1231,N_1005);
nand U4566 (N_4566,N_1532,N_195);
and U4567 (N_4567,N_2423,N_2373);
nor U4568 (N_4568,N_1364,N_916);
or U4569 (N_4569,N_2387,N_624);
and U4570 (N_4570,N_1611,N_2439);
or U4571 (N_4571,N_1993,N_1708);
nor U4572 (N_4572,N_1412,N_410);
nor U4573 (N_4573,N_525,N_1326);
nand U4574 (N_4574,N_2858,N_2882);
nor U4575 (N_4575,N_2830,N_2124);
xor U4576 (N_4576,N_2719,N_2402);
nand U4577 (N_4577,N_71,N_1909);
nand U4578 (N_4578,N_2903,N_2323);
or U4579 (N_4579,N_591,N_162);
nand U4580 (N_4580,N_1578,N_858);
and U4581 (N_4581,N_1313,N_296);
nor U4582 (N_4582,N_1704,N_1249);
and U4583 (N_4583,N_2491,N_1159);
or U4584 (N_4584,N_1595,N_1183);
nor U4585 (N_4585,N_1767,N_637);
and U4586 (N_4586,N_1456,N_1484);
or U4587 (N_4587,N_2529,N_2400);
or U4588 (N_4588,N_880,N_85);
nor U4589 (N_4589,N_1944,N_2898);
nand U4590 (N_4590,N_513,N_2930);
or U4591 (N_4591,N_1249,N_1385);
xnor U4592 (N_4592,N_1701,N_2151);
and U4593 (N_4593,N_1907,N_1494);
or U4594 (N_4594,N_584,N_1417);
nor U4595 (N_4595,N_2460,N_1002);
and U4596 (N_4596,N_2382,N_1860);
or U4597 (N_4597,N_2728,N_350);
or U4598 (N_4598,N_812,N_2530);
nand U4599 (N_4599,N_1285,N_565);
and U4600 (N_4600,N_2315,N_918);
nand U4601 (N_4601,N_279,N_1918);
and U4602 (N_4602,N_1558,N_2093);
nor U4603 (N_4603,N_306,N_2838);
nand U4604 (N_4604,N_2580,N_195);
and U4605 (N_4605,N_1825,N_763);
nor U4606 (N_4606,N_2685,N_279);
and U4607 (N_4607,N_2282,N_2143);
or U4608 (N_4608,N_1570,N_756);
nand U4609 (N_4609,N_2214,N_842);
and U4610 (N_4610,N_1557,N_659);
and U4611 (N_4611,N_105,N_867);
and U4612 (N_4612,N_1611,N_2465);
and U4613 (N_4613,N_692,N_376);
nor U4614 (N_4614,N_331,N_2431);
nand U4615 (N_4615,N_258,N_653);
nand U4616 (N_4616,N_1465,N_1332);
nor U4617 (N_4617,N_1647,N_2537);
nor U4618 (N_4618,N_2867,N_2404);
nor U4619 (N_4619,N_277,N_1358);
nor U4620 (N_4620,N_1737,N_743);
or U4621 (N_4621,N_619,N_1504);
and U4622 (N_4622,N_264,N_1046);
or U4623 (N_4623,N_1947,N_313);
or U4624 (N_4624,N_1063,N_1512);
and U4625 (N_4625,N_1365,N_946);
nor U4626 (N_4626,N_1832,N_785);
or U4627 (N_4627,N_2247,N_2248);
nor U4628 (N_4628,N_2770,N_1971);
and U4629 (N_4629,N_2436,N_798);
nor U4630 (N_4630,N_29,N_1470);
nand U4631 (N_4631,N_2406,N_1164);
or U4632 (N_4632,N_944,N_631);
nand U4633 (N_4633,N_1970,N_2379);
and U4634 (N_4634,N_1354,N_672);
or U4635 (N_4635,N_2201,N_1515);
and U4636 (N_4636,N_2720,N_425);
nor U4637 (N_4637,N_2579,N_1600);
nand U4638 (N_4638,N_362,N_2831);
nor U4639 (N_4639,N_755,N_2466);
nor U4640 (N_4640,N_2956,N_1056);
or U4641 (N_4641,N_351,N_2082);
nand U4642 (N_4642,N_1176,N_2385);
or U4643 (N_4643,N_2271,N_496);
and U4644 (N_4644,N_491,N_2666);
nand U4645 (N_4645,N_727,N_591);
nand U4646 (N_4646,N_449,N_1021);
nor U4647 (N_4647,N_579,N_2683);
nor U4648 (N_4648,N_2090,N_1355);
and U4649 (N_4649,N_1050,N_951);
and U4650 (N_4650,N_2903,N_2202);
nand U4651 (N_4651,N_1653,N_822);
nand U4652 (N_4652,N_753,N_2443);
nor U4653 (N_4653,N_2742,N_1404);
and U4654 (N_4654,N_2071,N_646);
nor U4655 (N_4655,N_84,N_1553);
and U4656 (N_4656,N_2883,N_1656);
nor U4657 (N_4657,N_830,N_1292);
xnor U4658 (N_4658,N_1820,N_2695);
nor U4659 (N_4659,N_2209,N_1505);
and U4660 (N_4660,N_1043,N_2761);
nand U4661 (N_4661,N_1926,N_2842);
or U4662 (N_4662,N_1657,N_386);
or U4663 (N_4663,N_2239,N_2299);
nand U4664 (N_4664,N_1472,N_790);
and U4665 (N_4665,N_1010,N_2654);
nand U4666 (N_4666,N_567,N_1298);
nand U4667 (N_4667,N_2864,N_2119);
and U4668 (N_4668,N_2856,N_1298);
nand U4669 (N_4669,N_1929,N_286);
xnor U4670 (N_4670,N_2481,N_1527);
and U4671 (N_4671,N_2457,N_1402);
and U4672 (N_4672,N_2207,N_1227);
nand U4673 (N_4673,N_4,N_1599);
or U4674 (N_4674,N_2329,N_191);
and U4675 (N_4675,N_221,N_493);
nor U4676 (N_4676,N_1176,N_1974);
nand U4677 (N_4677,N_512,N_1493);
and U4678 (N_4678,N_339,N_1825);
nand U4679 (N_4679,N_906,N_2493);
and U4680 (N_4680,N_2465,N_2911);
nand U4681 (N_4681,N_2841,N_2875);
or U4682 (N_4682,N_92,N_2185);
or U4683 (N_4683,N_209,N_1985);
or U4684 (N_4684,N_1851,N_1975);
nor U4685 (N_4685,N_556,N_311);
nand U4686 (N_4686,N_907,N_2087);
xor U4687 (N_4687,N_2893,N_2428);
nor U4688 (N_4688,N_1366,N_2450);
nor U4689 (N_4689,N_2914,N_1716);
and U4690 (N_4690,N_2877,N_1294);
nand U4691 (N_4691,N_1901,N_652);
nand U4692 (N_4692,N_831,N_600);
nor U4693 (N_4693,N_1876,N_1103);
or U4694 (N_4694,N_2557,N_2394);
nand U4695 (N_4695,N_202,N_364);
nand U4696 (N_4696,N_1373,N_2347);
nor U4697 (N_4697,N_1802,N_2786);
nor U4698 (N_4698,N_807,N_125);
nor U4699 (N_4699,N_1472,N_1319);
nor U4700 (N_4700,N_707,N_1346);
or U4701 (N_4701,N_2093,N_632);
nor U4702 (N_4702,N_2012,N_1458);
or U4703 (N_4703,N_2909,N_2608);
nor U4704 (N_4704,N_1474,N_2612);
nor U4705 (N_4705,N_214,N_219);
nor U4706 (N_4706,N_149,N_1255);
and U4707 (N_4707,N_2807,N_689);
nor U4708 (N_4708,N_933,N_2753);
nor U4709 (N_4709,N_2836,N_2782);
nor U4710 (N_4710,N_361,N_529);
or U4711 (N_4711,N_1236,N_1043);
nor U4712 (N_4712,N_1482,N_1260);
nand U4713 (N_4713,N_1793,N_2655);
nor U4714 (N_4714,N_2588,N_1440);
or U4715 (N_4715,N_1720,N_2303);
and U4716 (N_4716,N_2637,N_2107);
nor U4717 (N_4717,N_213,N_1740);
or U4718 (N_4718,N_2212,N_550);
nand U4719 (N_4719,N_723,N_1123);
or U4720 (N_4720,N_431,N_2635);
and U4721 (N_4721,N_2915,N_1078);
and U4722 (N_4722,N_1209,N_364);
nor U4723 (N_4723,N_2243,N_2100);
nor U4724 (N_4724,N_1047,N_2840);
and U4725 (N_4725,N_2036,N_2629);
xor U4726 (N_4726,N_1967,N_993);
or U4727 (N_4727,N_1605,N_754);
and U4728 (N_4728,N_689,N_2186);
and U4729 (N_4729,N_256,N_279);
nor U4730 (N_4730,N_673,N_494);
and U4731 (N_4731,N_282,N_2365);
nor U4732 (N_4732,N_1053,N_1366);
nand U4733 (N_4733,N_1037,N_2874);
nor U4734 (N_4734,N_2105,N_2617);
or U4735 (N_4735,N_917,N_1930);
nand U4736 (N_4736,N_2170,N_2773);
and U4737 (N_4737,N_1807,N_540);
nand U4738 (N_4738,N_2499,N_1629);
nor U4739 (N_4739,N_2347,N_480);
or U4740 (N_4740,N_649,N_736);
nor U4741 (N_4741,N_211,N_1379);
nand U4742 (N_4742,N_2841,N_1084);
or U4743 (N_4743,N_375,N_2094);
nand U4744 (N_4744,N_189,N_412);
or U4745 (N_4745,N_1550,N_232);
or U4746 (N_4746,N_1090,N_2136);
xnor U4747 (N_4747,N_380,N_2615);
nor U4748 (N_4748,N_1342,N_1778);
nand U4749 (N_4749,N_2593,N_619);
xnor U4750 (N_4750,N_1889,N_2873);
and U4751 (N_4751,N_2852,N_2516);
and U4752 (N_4752,N_923,N_517);
nand U4753 (N_4753,N_2863,N_2644);
nor U4754 (N_4754,N_516,N_88);
and U4755 (N_4755,N_834,N_2391);
nand U4756 (N_4756,N_189,N_2473);
or U4757 (N_4757,N_1198,N_2773);
and U4758 (N_4758,N_674,N_1880);
nor U4759 (N_4759,N_1090,N_2587);
nand U4760 (N_4760,N_126,N_2841);
and U4761 (N_4761,N_1234,N_769);
xnor U4762 (N_4762,N_1106,N_271);
nor U4763 (N_4763,N_608,N_238);
and U4764 (N_4764,N_125,N_784);
nand U4765 (N_4765,N_868,N_828);
nor U4766 (N_4766,N_221,N_986);
and U4767 (N_4767,N_1532,N_2381);
or U4768 (N_4768,N_2194,N_2);
and U4769 (N_4769,N_568,N_137);
nor U4770 (N_4770,N_793,N_536);
nand U4771 (N_4771,N_15,N_2860);
or U4772 (N_4772,N_82,N_2966);
nor U4773 (N_4773,N_2411,N_1782);
nand U4774 (N_4774,N_415,N_2186);
or U4775 (N_4775,N_1337,N_642);
or U4776 (N_4776,N_1806,N_677);
nor U4777 (N_4777,N_2929,N_582);
nand U4778 (N_4778,N_74,N_2528);
or U4779 (N_4779,N_1600,N_2530);
nand U4780 (N_4780,N_1649,N_57);
or U4781 (N_4781,N_2192,N_1351);
nand U4782 (N_4782,N_780,N_2450);
nor U4783 (N_4783,N_389,N_289);
and U4784 (N_4784,N_1111,N_2649);
nor U4785 (N_4785,N_584,N_2224);
nor U4786 (N_4786,N_2804,N_1481);
and U4787 (N_4787,N_1611,N_1466);
nand U4788 (N_4788,N_2561,N_2188);
nor U4789 (N_4789,N_2396,N_1870);
and U4790 (N_4790,N_1338,N_349);
and U4791 (N_4791,N_698,N_1470);
nand U4792 (N_4792,N_1716,N_164);
and U4793 (N_4793,N_1888,N_2124);
nor U4794 (N_4794,N_1327,N_978);
and U4795 (N_4795,N_1026,N_2824);
or U4796 (N_4796,N_2598,N_2210);
nor U4797 (N_4797,N_943,N_2209);
and U4798 (N_4798,N_2982,N_1428);
and U4799 (N_4799,N_1492,N_2241);
nor U4800 (N_4800,N_726,N_2270);
and U4801 (N_4801,N_2975,N_1907);
nor U4802 (N_4802,N_213,N_2593);
nor U4803 (N_4803,N_2088,N_2478);
nor U4804 (N_4804,N_2452,N_246);
and U4805 (N_4805,N_2983,N_1349);
nor U4806 (N_4806,N_2830,N_702);
and U4807 (N_4807,N_1182,N_81);
nor U4808 (N_4808,N_2690,N_2840);
nor U4809 (N_4809,N_612,N_2729);
and U4810 (N_4810,N_2611,N_1188);
nand U4811 (N_4811,N_1084,N_808);
or U4812 (N_4812,N_2237,N_2892);
nor U4813 (N_4813,N_933,N_2855);
nor U4814 (N_4814,N_314,N_897);
or U4815 (N_4815,N_2745,N_959);
and U4816 (N_4816,N_1669,N_1954);
or U4817 (N_4817,N_2346,N_388);
nor U4818 (N_4818,N_1537,N_1538);
and U4819 (N_4819,N_367,N_2326);
and U4820 (N_4820,N_1139,N_148);
nor U4821 (N_4821,N_232,N_999);
nand U4822 (N_4822,N_1412,N_2717);
and U4823 (N_4823,N_1857,N_1172);
or U4824 (N_4824,N_1067,N_2678);
nor U4825 (N_4825,N_468,N_1088);
or U4826 (N_4826,N_2933,N_1191);
nor U4827 (N_4827,N_2997,N_2394);
nor U4828 (N_4828,N_904,N_2085);
and U4829 (N_4829,N_2722,N_2724);
or U4830 (N_4830,N_748,N_2431);
or U4831 (N_4831,N_1534,N_2872);
nor U4832 (N_4832,N_1376,N_2468);
and U4833 (N_4833,N_1416,N_29);
or U4834 (N_4834,N_1940,N_430);
nand U4835 (N_4835,N_1176,N_1334);
nand U4836 (N_4836,N_2099,N_899);
nand U4837 (N_4837,N_1193,N_1398);
nor U4838 (N_4838,N_2381,N_988);
nand U4839 (N_4839,N_603,N_737);
or U4840 (N_4840,N_177,N_154);
nor U4841 (N_4841,N_2471,N_2917);
and U4842 (N_4842,N_910,N_1803);
nand U4843 (N_4843,N_2125,N_427);
or U4844 (N_4844,N_1664,N_1202);
or U4845 (N_4845,N_1063,N_2675);
and U4846 (N_4846,N_33,N_2024);
nand U4847 (N_4847,N_1313,N_1941);
nor U4848 (N_4848,N_895,N_634);
nand U4849 (N_4849,N_2881,N_1416);
or U4850 (N_4850,N_2889,N_2910);
nand U4851 (N_4851,N_129,N_231);
and U4852 (N_4852,N_551,N_492);
and U4853 (N_4853,N_1996,N_1203);
or U4854 (N_4854,N_2302,N_1975);
or U4855 (N_4855,N_96,N_2765);
or U4856 (N_4856,N_1092,N_2667);
or U4857 (N_4857,N_209,N_2371);
nand U4858 (N_4858,N_1758,N_2423);
nor U4859 (N_4859,N_2246,N_22);
nand U4860 (N_4860,N_656,N_2788);
nand U4861 (N_4861,N_2050,N_2012);
nand U4862 (N_4862,N_2319,N_400);
nand U4863 (N_4863,N_465,N_1639);
or U4864 (N_4864,N_815,N_515);
or U4865 (N_4865,N_2796,N_1892);
nand U4866 (N_4866,N_1308,N_2516);
nor U4867 (N_4867,N_1730,N_2488);
nand U4868 (N_4868,N_2692,N_2797);
nor U4869 (N_4869,N_2995,N_1731);
nor U4870 (N_4870,N_1991,N_2394);
or U4871 (N_4871,N_1146,N_2636);
or U4872 (N_4872,N_1923,N_267);
nand U4873 (N_4873,N_90,N_661);
nand U4874 (N_4874,N_1827,N_969);
and U4875 (N_4875,N_161,N_2143);
nor U4876 (N_4876,N_1051,N_2419);
nor U4877 (N_4877,N_432,N_761);
xor U4878 (N_4878,N_2387,N_280);
nor U4879 (N_4879,N_757,N_2116);
nand U4880 (N_4880,N_1667,N_1741);
nand U4881 (N_4881,N_993,N_1584);
and U4882 (N_4882,N_1029,N_1965);
nor U4883 (N_4883,N_1178,N_561);
nor U4884 (N_4884,N_1033,N_1235);
nor U4885 (N_4885,N_612,N_701);
or U4886 (N_4886,N_1719,N_2166);
xor U4887 (N_4887,N_1569,N_2975);
nand U4888 (N_4888,N_483,N_718);
nand U4889 (N_4889,N_1545,N_627);
and U4890 (N_4890,N_1596,N_1168);
nor U4891 (N_4891,N_898,N_964);
and U4892 (N_4892,N_2851,N_207);
or U4893 (N_4893,N_418,N_480);
nand U4894 (N_4894,N_601,N_2436);
nand U4895 (N_4895,N_2011,N_2361);
nand U4896 (N_4896,N_1613,N_1650);
and U4897 (N_4897,N_2627,N_2348);
or U4898 (N_4898,N_1445,N_623);
or U4899 (N_4899,N_906,N_1535);
nor U4900 (N_4900,N_2633,N_2754);
or U4901 (N_4901,N_1881,N_2160);
or U4902 (N_4902,N_877,N_2659);
nor U4903 (N_4903,N_1733,N_1853);
or U4904 (N_4904,N_170,N_1458);
nor U4905 (N_4905,N_1753,N_1717);
nor U4906 (N_4906,N_1401,N_1774);
and U4907 (N_4907,N_192,N_1084);
nor U4908 (N_4908,N_1332,N_2155);
nand U4909 (N_4909,N_336,N_2692);
and U4910 (N_4910,N_2253,N_1930);
nor U4911 (N_4911,N_1312,N_941);
and U4912 (N_4912,N_2839,N_1717);
nand U4913 (N_4913,N_2861,N_2953);
nor U4914 (N_4914,N_2800,N_585);
nand U4915 (N_4915,N_88,N_243);
or U4916 (N_4916,N_1777,N_2970);
and U4917 (N_4917,N_82,N_210);
and U4918 (N_4918,N_88,N_2108);
or U4919 (N_4919,N_2943,N_1664);
or U4920 (N_4920,N_1310,N_2764);
nand U4921 (N_4921,N_548,N_702);
nand U4922 (N_4922,N_132,N_2817);
nor U4923 (N_4923,N_2988,N_2263);
nand U4924 (N_4924,N_417,N_1059);
nor U4925 (N_4925,N_245,N_662);
nand U4926 (N_4926,N_1484,N_1234);
nand U4927 (N_4927,N_2508,N_562);
and U4928 (N_4928,N_424,N_1233);
nor U4929 (N_4929,N_1914,N_2989);
nor U4930 (N_4930,N_276,N_2825);
nand U4931 (N_4931,N_2427,N_2623);
or U4932 (N_4932,N_928,N_2527);
nand U4933 (N_4933,N_2069,N_2293);
nor U4934 (N_4934,N_523,N_1737);
or U4935 (N_4935,N_754,N_1528);
or U4936 (N_4936,N_1926,N_8);
nor U4937 (N_4937,N_2737,N_1198);
nand U4938 (N_4938,N_1781,N_598);
and U4939 (N_4939,N_2135,N_1283);
and U4940 (N_4940,N_368,N_1248);
or U4941 (N_4941,N_2153,N_2689);
and U4942 (N_4942,N_471,N_455);
and U4943 (N_4943,N_2843,N_1005);
nand U4944 (N_4944,N_2607,N_393);
and U4945 (N_4945,N_2472,N_1062);
nor U4946 (N_4946,N_1907,N_270);
and U4947 (N_4947,N_1049,N_1480);
and U4948 (N_4948,N_1870,N_2480);
nand U4949 (N_4949,N_2937,N_1105);
and U4950 (N_4950,N_1792,N_922);
and U4951 (N_4951,N_408,N_360);
nand U4952 (N_4952,N_217,N_1885);
xor U4953 (N_4953,N_688,N_1620);
nor U4954 (N_4954,N_1107,N_1920);
nand U4955 (N_4955,N_2858,N_976);
nand U4956 (N_4956,N_394,N_2018);
and U4957 (N_4957,N_2541,N_522);
and U4958 (N_4958,N_855,N_1624);
nor U4959 (N_4959,N_863,N_2153);
xnor U4960 (N_4960,N_1966,N_1063);
nor U4961 (N_4961,N_602,N_1758);
nand U4962 (N_4962,N_1048,N_1901);
and U4963 (N_4963,N_1847,N_2534);
and U4964 (N_4964,N_111,N_2247);
or U4965 (N_4965,N_1647,N_2139);
nor U4966 (N_4966,N_1936,N_453);
and U4967 (N_4967,N_546,N_684);
nand U4968 (N_4968,N_454,N_2382);
and U4969 (N_4969,N_888,N_169);
or U4970 (N_4970,N_2113,N_1903);
and U4971 (N_4971,N_1827,N_2859);
and U4972 (N_4972,N_2130,N_1826);
or U4973 (N_4973,N_2097,N_527);
or U4974 (N_4974,N_2851,N_1751);
nand U4975 (N_4975,N_2230,N_1729);
and U4976 (N_4976,N_352,N_61);
nor U4977 (N_4977,N_932,N_2235);
nor U4978 (N_4978,N_451,N_2256);
xnor U4979 (N_4979,N_2973,N_2855);
or U4980 (N_4980,N_2272,N_1453);
and U4981 (N_4981,N_371,N_1974);
and U4982 (N_4982,N_718,N_1547);
nand U4983 (N_4983,N_1287,N_643);
nor U4984 (N_4984,N_1607,N_1853);
and U4985 (N_4985,N_2311,N_742);
or U4986 (N_4986,N_769,N_65);
nor U4987 (N_4987,N_281,N_1867);
and U4988 (N_4988,N_756,N_603);
nand U4989 (N_4989,N_1254,N_1758);
nor U4990 (N_4990,N_1109,N_984);
and U4991 (N_4991,N_1628,N_1813);
nor U4992 (N_4992,N_783,N_890);
nand U4993 (N_4993,N_1096,N_1472);
nor U4994 (N_4994,N_2790,N_1078);
xnor U4995 (N_4995,N_690,N_353);
and U4996 (N_4996,N_1827,N_318);
and U4997 (N_4997,N_2017,N_2236);
nand U4998 (N_4998,N_635,N_409);
nand U4999 (N_4999,N_2519,N_136);
and U5000 (N_5000,N_887,N_2014);
nand U5001 (N_5001,N_2212,N_1150);
nor U5002 (N_5002,N_2957,N_2772);
nor U5003 (N_5003,N_2230,N_2245);
nor U5004 (N_5004,N_1679,N_2200);
nor U5005 (N_5005,N_877,N_1311);
nor U5006 (N_5006,N_501,N_2486);
nor U5007 (N_5007,N_1177,N_1413);
nand U5008 (N_5008,N_792,N_2195);
nand U5009 (N_5009,N_1820,N_486);
nand U5010 (N_5010,N_1664,N_2262);
nand U5011 (N_5011,N_2230,N_2987);
nand U5012 (N_5012,N_2081,N_1837);
nand U5013 (N_5013,N_456,N_866);
nor U5014 (N_5014,N_1927,N_457);
xnor U5015 (N_5015,N_2645,N_2973);
nor U5016 (N_5016,N_2851,N_1123);
or U5017 (N_5017,N_312,N_2579);
or U5018 (N_5018,N_1262,N_2355);
and U5019 (N_5019,N_868,N_2161);
or U5020 (N_5020,N_151,N_2915);
or U5021 (N_5021,N_833,N_586);
or U5022 (N_5022,N_1404,N_120);
nand U5023 (N_5023,N_76,N_736);
nor U5024 (N_5024,N_2010,N_2029);
or U5025 (N_5025,N_2180,N_1309);
nand U5026 (N_5026,N_1664,N_2924);
and U5027 (N_5027,N_208,N_915);
or U5028 (N_5028,N_2188,N_1479);
nor U5029 (N_5029,N_996,N_2809);
nand U5030 (N_5030,N_2794,N_318);
and U5031 (N_5031,N_772,N_1970);
nand U5032 (N_5032,N_219,N_928);
or U5033 (N_5033,N_271,N_635);
nor U5034 (N_5034,N_675,N_600);
nand U5035 (N_5035,N_1882,N_2276);
nor U5036 (N_5036,N_1773,N_775);
and U5037 (N_5037,N_514,N_465);
nand U5038 (N_5038,N_2505,N_822);
and U5039 (N_5039,N_2026,N_1766);
and U5040 (N_5040,N_2243,N_1400);
nand U5041 (N_5041,N_2792,N_2452);
nand U5042 (N_5042,N_1780,N_2243);
nor U5043 (N_5043,N_2303,N_1285);
nor U5044 (N_5044,N_2629,N_893);
and U5045 (N_5045,N_2422,N_964);
nand U5046 (N_5046,N_2798,N_2864);
or U5047 (N_5047,N_1684,N_2521);
or U5048 (N_5048,N_2078,N_2024);
and U5049 (N_5049,N_603,N_431);
nand U5050 (N_5050,N_2816,N_1260);
or U5051 (N_5051,N_1893,N_1562);
nor U5052 (N_5052,N_2332,N_1727);
xor U5053 (N_5053,N_2077,N_2729);
and U5054 (N_5054,N_455,N_2735);
or U5055 (N_5055,N_2596,N_2734);
nand U5056 (N_5056,N_2664,N_2515);
or U5057 (N_5057,N_1234,N_1204);
or U5058 (N_5058,N_54,N_361);
and U5059 (N_5059,N_591,N_387);
or U5060 (N_5060,N_641,N_745);
nand U5061 (N_5061,N_1749,N_1349);
and U5062 (N_5062,N_2377,N_2949);
nand U5063 (N_5063,N_292,N_2872);
xnor U5064 (N_5064,N_1973,N_312);
nand U5065 (N_5065,N_2601,N_1821);
and U5066 (N_5066,N_2410,N_2294);
and U5067 (N_5067,N_2689,N_821);
nor U5068 (N_5068,N_341,N_1470);
nand U5069 (N_5069,N_1073,N_1133);
and U5070 (N_5070,N_1866,N_1588);
nand U5071 (N_5071,N_983,N_672);
nor U5072 (N_5072,N_2417,N_1060);
and U5073 (N_5073,N_76,N_474);
nor U5074 (N_5074,N_386,N_710);
nand U5075 (N_5075,N_1695,N_1313);
nor U5076 (N_5076,N_417,N_810);
and U5077 (N_5077,N_1661,N_2);
nand U5078 (N_5078,N_585,N_2836);
nor U5079 (N_5079,N_788,N_2158);
or U5080 (N_5080,N_1838,N_1912);
nor U5081 (N_5081,N_2258,N_1833);
nor U5082 (N_5082,N_1645,N_2087);
nand U5083 (N_5083,N_2246,N_201);
nor U5084 (N_5084,N_766,N_2012);
nor U5085 (N_5085,N_2291,N_188);
nor U5086 (N_5086,N_1944,N_1013);
or U5087 (N_5087,N_25,N_1571);
nor U5088 (N_5088,N_1016,N_2042);
and U5089 (N_5089,N_2070,N_1974);
nand U5090 (N_5090,N_1221,N_832);
and U5091 (N_5091,N_1898,N_2660);
or U5092 (N_5092,N_643,N_697);
nand U5093 (N_5093,N_874,N_1052);
and U5094 (N_5094,N_2479,N_772);
nor U5095 (N_5095,N_1138,N_1777);
and U5096 (N_5096,N_2245,N_2279);
nand U5097 (N_5097,N_1878,N_2084);
nand U5098 (N_5098,N_908,N_761);
and U5099 (N_5099,N_1558,N_31);
nor U5100 (N_5100,N_2214,N_1447);
nor U5101 (N_5101,N_87,N_2984);
or U5102 (N_5102,N_1911,N_2574);
nor U5103 (N_5103,N_2767,N_2119);
or U5104 (N_5104,N_2546,N_2114);
and U5105 (N_5105,N_2614,N_1244);
nor U5106 (N_5106,N_851,N_1696);
and U5107 (N_5107,N_952,N_244);
xor U5108 (N_5108,N_968,N_1865);
nor U5109 (N_5109,N_1355,N_1871);
nand U5110 (N_5110,N_460,N_2538);
nor U5111 (N_5111,N_1546,N_1795);
nand U5112 (N_5112,N_2867,N_2912);
or U5113 (N_5113,N_1924,N_1562);
and U5114 (N_5114,N_363,N_884);
and U5115 (N_5115,N_1623,N_241);
and U5116 (N_5116,N_2427,N_1724);
or U5117 (N_5117,N_477,N_2417);
and U5118 (N_5118,N_1989,N_458);
or U5119 (N_5119,N_1693,N_1821);
nor U5120 (N_5120,N_2019,N_2412);
nand U5121 (N_5121,N_1715,N_423);
or U5122 (N_5122,N_87,N_2513);
and U5123 (N_5123,N_2955,N_1914);
and U5124 (N_5124,N_846,N_835);
nand U5125 (N_5125,N_1507,N_2471);
xor U5126 (N_5126,N_174,N_1063);
nand U5127 (N_5127,N_2059,N_1422);
nand U5128 (N_5128,N_1622,N_2969);
and U5129 (N_5129,N_415,N_1362);
nand U5130 (N_5130,N_562,N_2241);
and U5131 (N_5131,N_1339,N_1040);
or U5132 (N_5132,N_2787,N_2045);
and U5133 (N_5133,N_742,N_2910);
and U5134 (N_5134,N_1556,N_1886);
nand U5135 (N_5135,N_1643,N_579);
nand U5136 (N_5136,N_2041,N_1842);
nand U5137 (N_5137,N_75,N_1747);
or U5138 (N_5138,N_632,N_303);
or U5139 (N_5139,N_1799,N_2654);
and U5140 (N_5140,N_1784,N_2616);
or U5141 (N_5141,N_1828,N_1050);
or U5142 (N_5142,N_2889,N_260);
and U5143 (N_5143,N_2,N_2575);
and U5144 (N_5144,N_1558,N_406);
xor U5145 (N_5145,N_213,N_552);
nand U5146 (N_5146,N_741,N_1824);
nand U5147 (N_5147,N_464,N_255);
nand U5148 (N_5148,N_602,N_2849);
or U5149 (N_5149,N_77,N_427);
or U5150 (N_5150,N_1646,N_1557);
or U5151 (N_5151,N_2439,N_102);
and U5152 (N_5152,N_2889,N_1955);
and U5153 (N_5153,N_1845,N_151);
and U5154 (N_5154,N_2886,N_1460);
or U5155 (N_5155,N_822,N_1719);
or U5156 (N_5156,N_2353,N_2640);
nand U5157 (N_5157,N_567,N_286);
nor U5158 (N_5158,N_2581,N_592);
and U5159 (N_5159,N_1835,N_1274);
nor U5160 (N_5160,N_875,N_1324);
nor U5161 (N_5161,N_1882,N_573);
nor U5162 (N_5162,N_1168,N_1457);
xor U5163 (N_5163,N_2614,N_2958);
or U5164 (N_5164,N_823,N_1821);
or U5165 (N_5165,N_2401,N_1021);
or U5166 (N_5166,N_2215,N_79);
nand U5167 (N_5167,N_940,N_120);
or U5168 (N_5168,N_1110,N_2679);
nor U5169 (N_5169,N_2104,N_284);
or U5170 (N_5170,N_2880,N_1459);
and U5171 (N_5171,N_423,N_404);
and U5172 (N_5172,N_2816,N_1673);
nand U5173 (N_5173,N_1218,N_232);
nor U5174 (N_5174,N_2694,N_2236);
nor U5175 (N_5175,N_2322,N_2036);
or U5176 (N_5176,N_1432,N_774);
or U5177 (N_5177,N_2134,N_893);
or U5178 (N_5178,N_460,N_2722);
or U5179 (N_5179,N_281,N_1363);
and U5180 (N_5180,N_1970,N_1580);
or U5181 (N_5181,N_771,N_460);
and U5182 (N_5182,N_268,N_570);
xor U5183 (N_5183,N_2790,N_1733);
or U5184 (N_5184,N_1638,N_100);
nor U5185 (N_5185,N_1708,N_736);
or U5186 (N_5186,N_1209,N_2009);
xnor U5187 (N_5187,N_1839,N_1945);
nand U5188 (N_5188,N_1949,N_1964);
or U5189 (N_5189,N_1340,N_1048);
nor U5190 (N_5190,N_2800,N_859);
nor U5191 (N_5191,N_228,N_1005);
nor U5192 (N_5192,N_2371,N_2108);
or U5193 (N_5193,N_579,N_1815);
nor U5194 (N_5194,N_1058,N_2710);
nand U5195 (N_5195,N_1112,N_1683);
nand U5196 (N_5196,N_1552,N_153);
nor U5197 (N_5197,N_291,N_1356);
or U5198 (N_5198,N_150,N_2824);
or U5199 (N_5199,N_302,N_776);
and U5200 (N_5200,N_2939,N_2974);
and U5201 (N_5201,N_1477,N_1949);
or U5202 (N_5202,N_799,N_2183);
and U5203 (N_5203,N_2633,N_228);
nand U5204 (N_5204,N_732,N_1137);
nor U5205 (N_5205,N_1770,N_2567);
nand U5206 (N_5206,N_606,N_1427);
nor U5207 (N_5207,N_2347,N_812);
nand U5208 (N_5208,N_2594,N_729);
or U5209 (N_5209,N_131,N_2635);
or U5210 (N_5210,N_2852,N_1558);
xnor U5211 (N_5211,N_2130,N_1598);
nor U5212 (N_5212,N_949,N_86);
nor U5213 (N_5213,N_231,N_407);
and U5214 (N_5214,N_912,N_515);
nand U5215 (N_5215,N_2745,N_619);
or U5216 (N_5216,N_2652,N_2109);
or U5217 (N_5217,N_1332,N_1159);
or U5218 (N_5218,N_1202,N_672);
or U5219 (N_5219,N_931,N_2065);
xor U5220 (N_5220,N_607,N_507);
nand U5221 (N_5221,N_1551,N_2336);
or U5222 (N_5222,N_2697,N_2618);
and U5223 (N_5223,N_94,N_2239);
or U5224 (N_5224,N_137,N_2205);
and U5225 (N_5225,N_2967,N_1263);
nor U5226 (N_5226,N_796,N_1275);
nor U5227 (N_5227,N_1447,N_2767);
nand U5228 (N_5228,N_2835,N_1305);
and U5229 (N_5229,N_334,N_2376);
or U5230 (N_5230,N_1447,N_787);
nor U5231 (N_5231,N_1642,N_228);
nor U5232 (N_5232,N_57,N_1192);
and U5233 (N_5233,N_2309,N_1037);
or U5234 (N_5234,N_2653,N_2160);
nand U5235 (N_5235,N_1724,N_1648);
nor U5236 (N_5236,N_1990,N_2433);
nand U5237 (N_5237,N_834,N_64);
and U5238 (N_5238,N_71,N_1752);
nand U5239 (N_5239,N_1399,N_1616);
or U5240 (N_5240,N_1941,N_2000);
nor U5241 (N_5241,N_1251,N_1094);
nand U5242 (N_5242,N_2145,N_366);
nor U5243 (N_5243,N_1206,N_1129);
nand U5244 (N_5244,N_1894,N_2785);
and U5245 (N_5245,N_800,N_2886);
xor U5246 (N_5246,N_1022,N_860);
and U5247 (N_5247,N_1004,N_2139);
nor U5248 (N_5248,N_2155,N_144);
and U5249 (N_5249,N_775,N_1516);
or U5250 (N_5250,N_757,N_852);
and U5251 (N_5251,N_125,N_1797);
and U5252 (N_5252,N_2047,N_2940);
and U5253 (N_5253,N_1170,N_2703);
xor U5254 (N_5254,N_671,N_1863);
or U5255 (N_5255,N_2525,N_2438);
nor U5256 (N_5256,N_2670,N_1125);
xor U5257 (N_5257,N_2488,N_868);
nor U5258 (N_5258,N_1485,N_860);
nand U5259 (N_5259,N_84,N_2982);
nand U5260 (N_5260,N_1175,N_932);
and U5261 (N_5261,N_276,N_1875);
or U5262 (N_5262,N_2250,N_472);
nand U5263 (N_5263,N_2247,N_2774);
nand U5264 (N_5264,N_978,N_25);
and U5265 (N_5265,N_798,N_70);
or U5266 (N_5266,N_423,N_645);
nand U5267 (N_5267,N_2821,N_1638);
and U5268 (N_5268,N_2670,N_2969);
or U5269 (N_5269,N_1177,N_1789);
nand U5270 (N_5270,N_1587,N_2120);
nor U5271 (N_5271,N_98,N_2150);
nand U5272 (N_5272,N_271,N_1553);
and U5273 (N_5273,N_2888,N_2589);
and U5274 (N_5274,N_766,N_2671);
and U5275 (N_5275,N_2336,N_2004);
or U5276 (N_5276,N_2799,N_598);
nor U5277 (N_5277,N_1612,N_2635);
or U5278 (N_5278,N_966,N_926);
nor U5279 (N_5279,N_945,N_362);
or U5280 (N_5280,N_264,N_2789);
or U5281 (N_5281,N_2002,N_2013);
or U5282 (N_5282,N_1544,N_2481);
nand U5283 (N_5283,N_2348,N_1379);
nor U5284 (N_5284,N_1963,N_2128);
and U5285 (N_5285,N_1917,N_1050);
or U5286 (N_5286,N_1401,N_1714);
or U5287 (N_5287,N_66,N_2242);
nor U5288 (N_5288,N_2481,N_2240);
or U5289 (N_5289,N_572,N_1588);
and U5290 (N_5290,N_2122,N_2253);
nor U5291 (N_5291,N_1797,N_2382);
and U5292 (N_5292,N_398,N_2453);
and U5293 (N_5293,N_192,N_1142);
nor U5294 (N_5294,N_2333,N_502);
and U5295 (N_5295,N_500,N_1370);
and U5296 (N_5296,N_2888,N_581);
and U5297 (N_5297,N_2006,N_2835);
nand U5298 (N_5298,N_2753,N_463);
nand U5299 (N_5299,N_211,N_1456);
nand U5300 (N_5300,N_2749,N_1991);
nand U5301 (N_5301,N_1559,N_772);
xnor U5302 (N_5302,N_2053,N_1975);
nand U5303 (N_5303,N_264,N_1438);
nor U5304 (N_5304,N_288,N_1558);
nand U5305 (N_5305,N_874,N_1183);
or U5306 (N_5306,N_2701,N_1464);
or U5307 (N_5307,N_2300,N_2501);
and U5308 (N_5308,N_698,N_1434);
nor U5309 (N_5309,N_1123,N_60);
xor U5310 (N_5310,N_2721,N_1703);
nand U5311 (N_5311,N_1698,N_300);
xor U5312 (N_5312,N_723,N_788);
or U5313 (N_5313,N_84,N_1658);
nor U5314 (N_5314,N_2695,N_2002);
and U5315 (N_5315,N_2463,N_1185);
nor U5316 (N_5316,N_1503,N_1829);
and U5317 (N_5317,N_2050,N_785);
nor U5318 (N_5318,N_793,N_2219);
nand U5319 (N_5319,N_224,N_2150);
nand U5320 (N_5320,N_531,N_936);
and U5321 (N_5321,N_1227,N_1322);
and U5322 (N_5322,N_1334,N_1726);
and U5323 (N_5323,N_1587,N_576);
or U5324 (N_5324,N_2684,N_738);
nor U5325 (N_5325,N_972,N_1433);
or U5326 (N_5326,N_2252,N_1735);
nand U5327 (N_5327,N_2096,N_2336);
nor U5328 (N_5328,N_1400,N_2131);
or U5329 (N_5329,N_1202,N_382);
or U5330 (N_5330,N_1409,N_743);
nor U5331 (N_5331,N_122,N_2691);
and U5332 (N_5332,N_615,N_1819);
nor U5333 (N_5333,N_1507,N_257);
and U5334 (N_5334,N_358,N_1387);
xnor U5335 (N_5335,N_1819,N_1712);
nor U5336 (N_5336,N_2141,N_1354);
xor U5337 (N_5337,N_223,N_925);
and U5338 (N_5338,N_1200,N_2101);
or U5339 (N_5339,N_1383,N_435);
or U5340 (N_5340,N_1901,N_125);
or U5341 (N_5341,N_1593,N_1143);
xor U5342 (N_5342,N_1390,N_2869);
or U5343 (N_5343,N_1227,N_1781);
or U5344 (N_5344,N_953,N_732);
and U5345 (N_5345,N_2926,N_2260);
nor U5346 (N_5346,N_371,N_2145);
and U5347 (N_5347,N_1706,N_315);
nor U5348 (N_5348,N_2231,N_733);
or U5349 (N_5349,N_18,N_1089);
or U5350 (N_5350,N_2184,N_2125);
and U5351 (N_5351,N_811,N_521);
nand U5352 (N_5352,N_1125,N_1001);
nor U5353 (N_5353,N_2472,N_2145);
nand U5354 (N_5354,N_491,N_2304);
and U5355 (N_5355,N_1229,N_1294);
or U5356 (N_5356,N_2307,N_1758);
nand U5357 (N_5357,N_203,N_459);
or U5358 (N_5358,N_3,N_1872);
nor U5359 (N_5359,N_2792,N_1295);
or U5360 (N_5360,N_542,N_1761);
nand U5361 (N_5361,N_2209,N_193);
and U5362 (N_5362,N_1237,N_2920);
nand U5363 (N_5363,N_190,N_2115);
and U5364 (N_5364,N_476,N_957);
nor U5365 (N_5365,N_1683,N_2464);
nor U5366 (N_5366,N_1726,N_621);
and U5367 (N_5367,N_858,N_1823);
and U5368 (N_5368,N_19,N_1105);
nor U5369 (N_5369,N_1259,N_50);
nand U5370 (N_5370,N_954,N_125);
or U5371 (N_5371,N_2378,N_2308);
nor U5372 (N_5372,N_2625,N_2822);
or U5373 (N_5373,N_225,N_2472);
xor U5374 (N_5374,N_1699,N_1877);
and U5375 (N_5375,N_1531,N_143);
and U5376 (N_5376,N_2450,N_2860);
xor U5377 (N_5377,N_1504,N_2192);
or U5378 (N_5378,N_1014,N_1433);
nor U5379 (N_5379,N_137,N_905);
nand U5380 (N_5380,N_1218,N_1155);
or U5381 (N_5381,N_2578,N_90);
nand U5382 (N_5382,N_630,N_802);
nand U5383 (N_5383,N_2387,N_71);
and U5384 (N_5384,N_53,N_910);
nand U5385 (N_5385,N_2785,N_2733);
nand U5386 (N_5386,N_812,N_996);
or U5387 (N_5387,N_1630,N_1408);
nor U5388 (N_5388,N_392,N_1776);
nor U5389 (N_5389,N_1159,N_1791);
nand U5390 (N_5390,N_1378,N_1210);
nand U5391 (N_5391,N_1364,N_1013);
nand U5392 (N_5392,N_1234,N_7);
and U5393 (N_5393,N_542,N_1640);
nor U5394 (N_5394,N_1146,N_261);
nand U5395 (N_5395,N_539,N_2581);
nand U5396 (N_5396,N_1758,N_1028);
nor U5397 (N_5397,N_2457,N_1793);
or U5398 (N_5398,N_1409,N_1094);
and U5399 (N_5399,N_476,N_1555);
nand U5400 (N_5400,N_2753,N_1835);
nand U5401 (N_5401,N_1499,N_335);
nor U5402 (N_5402,N_2815,N_2083);
or U5403 (N_5403,N_1283,N_873);
and U5404 (N_5404,N_2204,N_1482);
or U5405 (N_5405,N_2670,N_1906);
or U5406 (N_5406,N_587,N_2453);
nor U5407 (N_5407,N_402,N_133);
or U5408 (N_5408,N_966,N_2213);
xor U5409 (N_5409,N_2563,N_1462);
nand U5410 (N_5410,N_2846,N_1471);
nand U5411 (N_5411,N_150,N_887);
or U5412 (N_5412,N_926,N_164);
nor U5413 (N_5413,N_2890,N_1941);
or U5414 (N_5414,N_1687,N_2813);
nor U5415 (N_5415,N_757,N_161);
or U5416 (N_5416,N_591,N_639);
and U5417 (N_5417,N_675,N_2751);
or U5418 (N_5418,N_607,N_1996);
nor U5419 (N_5419,N_1194,N_1270);
xor U5420 (N_5420,N_2021,N_2255);
or U5421 (N_5421,N_402,N_2907);
or U5422 (N_5422,N_1661,N_1044);
nand U5423 (N_5423,N_468,N_2910);
nand U5424 (N_5424,N_2696,N_2673);
and U5425 (N_5425,N_2115,N_546);
and U5426 (N_5426,N_2493,N_2015);
and U5427 (N_5427,N_1472,N_559);
and U5428 (N_5428,N_2406,N_692);
and U5429 (N_5429,N_2590,N_45);
and U5430 (N_5430,N_1526,N_1931);
and U5431 (N_5431,N_2576,N_2476);
nand U5432 (N_5432,N_1976,N_568);
nand U5433 (N_5433,N_341,N_1727);
or U5434 (N_5434,N_2403,N_1610);
nor U5435 (N_5435,N_2399,N_2749);
nand U5436 (N_5436,N_205,N_774);
nor U5437 (N_5437,N_1870,N_943);
or U5438 (N_5438,N_1366,N_424);
nand U5439 (N_5439,N_2829,N_38);
nor U5440 (N_5440,N_2680,N_139);
nor U5441 (N_5441,N_785,N_2913);
and U5442 (N_5442,N_2415,N_2022);
nor U5443 (N_5443,N_399,N_423);
or U5444 (N_5444,N_2606,N_56);
nor U5445 (N_5445,N_2993,N_406);
or U5446 (N_5446,N_626,N_462);
nor U5447 (N_5447,N_369,N_522);
and U5448 (N_5448,N_2502,N_57);
or U5449 (N_5449,N_1274,N_1437);
and U5450 (N_5450,N_2506,N_965);
and U5451 (N_5451,N_979,N_1038);
and U5452 (N_5452,N_1157,N_2711);
nor U5453 (N_5453,N_2623,N_1211);
nand U5454 (N_5454,N_801,N_2061);
nor U5455 (N_5455,N_305,N_1590);
and U5456 (N_5456,N_1420,N_934);
nor U5457 (N_5457,N_1754,N_2916);
nand U5458 (N_5458,N_57,N_100);
nand U5459 (N_5459,N_1006,N_2284);
xnor U5460 (N_5460,N_2088,N_443);
or U5461 (N_5461,N_2126,N_1791);
and U5462 (N_5462,N_1362,N_2037);
nor U5463 (N_5463,N_1554,N_2916);
nor U5464 (N_5464,N_2787,N_414);
nor U5465 (N_5465,N_2854,N_514);
and U5466 (N_5466,N_756,N_1909);
and U5467 (N_5467,N_2612,N_900);
nor U5468 (N_5468,N_1851,N_2093);
nand U5469 (N_5469,N_2072,N_1012);
or U5470 (N_5470,N_2099,N_2250);
nand U5471 (N_5471,N_524,N_1086);
nor U5472 (N_5472,N_2532,N_1032);
nor U5473 (N_5473,N_2195,N_1398);
or U5474 (N_5474,N_904,N_1809);
nand U5475 (N_5475,N_2680,N_2524);
nand U5476 (N_5476,N_493,N_2383);
or U5477 (N_5477,N_138,N_1374);
or U5478 (N_5478,N_898,N_2017);
or U5479 (N_5479,N_2052,N_2044);
nor U5480 (N_5480,N_1492,N_1686);
nand U5481 (N_5481,N_2462,N_2591);
nand U5482 (N_5482,N_2343,N_1330);
and U5483 (N_5483,N_1641,N_2753);
nor U5484 (N_5484,N_2051,N_465);
nand U5485 (N_5485,N_2172,N_2342);
nor U5486 (N_5486,N_2185,N_2371);
nor U5487 (N_5487,N_5,N_1990);
and U5488 (N_5488,N_76,N_717);
and U5489 (N_5489,N_1028,N_1620);
nor U5490 (N_5490,N_2845,N_1085);
nor U5491 (N_5491,N_831,N_2132);
nand U5492 (N_5492,N_11,N_47);
or U5493 (N_5493,N_1994,N_1692);
nor U5494 (N_5494,N_598,N_1472);
nor U5495 (N_5495,N_2441,N_2490);
and U5496 (N_5496,N_833,N_826);
nand U5497 (N_5497,N_1280,N_2784);
nand U5498 (N_5498,N_1747,N_2336);
or U5499 (N_5499,N_1517,N_1672);
or U5500 (N_5500,N_2908,N_1094);
or U5501 (N_5501,N_1753,N_1367);
or U5502 (N_5502,N_1021,N_295);
and U5503 (N_5503,N_929,N_4);
and U5504 (N_5504,N_1889,N_2629);
xnor U5505 (N_5505,N_1338,N_103);
nor U5506 (N_5506,N_1736,N_2657);
or U5507 (N_5507,N_1375,N_2563);
and U5508 (N_5508,N_1154,N_2574);
nand U5509 (N_5509,N_2764,N_2295);
nor U5510 (N_5510,N_1454,N_657);
or U5511 (N_5511,N_2216,N_434);
or U5512 (N_5512,N_621,N_1877);
nor U5513 (N_5513,N_2318,N_1512);
and U5514 (N_5514,N_2661,N_1152);
nand U5515 (N_5515,N_2765,N_662);
and U5516 (N_5516,N_1902,N_162);
nand U5517 (N_5517,N_2964,N_2453);
nand U5518 (N_5518,N_2279,N_1779);
nand U5519 (N_5519,N_1139,N_1903);
and U5520 (N_5520,N_1611,N_2921);
and U5521 (N_5521,N_960,N_1520);
or U5522 (N_5522,N_2768,N_586);
and U5523 (N_5523,N_2264,N_1538);
nand U5524 (N_5524,N_596,N_1040);
or U5525 (N_5525,N_2587,N_372);
nor U5526 (N_5526,N_2693,N_2854);
nand U5527 (N_5527,N_2593,N_690);
and U5528 (N_5528,N_2120,N_1253);
nor U5529 (N_5529,N_927,N_1682);
or U5530 (N_5530,N_448,N_1516);
xor U5531 (N_5531,N_823,N_318);
or U5532 (N_5532,N_2757,N_1519);
nor U5533 (N_5533,N_1316,N_318);
or U5534 (N_5534,N_2912,N_694);
or U5535 (N_5535,N_824,N_1310);
or U5536 (N_5536,N_2063,N_373);
or U5537 (N_5537,N_2911,N_375);
nor U5538 (N_5538,N_1823,N_1222);
and U5539 (N_5539,N_2231,N_1010);
nand U5540 (N_5540,N_1069,N_1790);
nor U5541 (N_5541,N_537,N_917);
nand U5542 (N_5542,N_2362,N_1406);
nor U5543 (N_5543,N_700,N_2982);
and U5544 (N_5544,N_873,N_478);
or U5545 (N_5545,N_2770,N_2556);
nand U5546 (N_5546,N_89,N_1407);
nor U5547 (N_5547,N_409,N_1984);
and U5548 (N_5548,N_1572,N_2613);
and U5549 (N_5549,N_1018,N_605);
or U5550 (N_5550,N_752,N_993);
nand U5551 (N_5551,N_2282,N_2648);
and U5552 (N_5552,N_2988,N_1865);
or U5553 (N_5553,N_736,N_822);
xnor U5554 (N_5554,N_1028,N_380);
or U5555 (N_5555,N_852,N_59);
or U5556 (N_5556,N_1416,N_2734);
xor U5557 (N_5557,N_28,N_1115);
or U5558 (N_5558,N_543,N_656);
or U5559 (N_5559,N_880,N_1158);
nor U5560 (N_5560,N_1299,N_133);
or U5561 (N_5561,N_50,N_1540);
and U5562 (N_5562,N_554,N_61);
xor U5563 (N_5563,N_320,N_2691);
nand U5564 (N_5564,N_1058,N_1611);
nor U5565 (N_5565,N_498,N_1838);
or U5566 (N_5566,N_1310,N_2081);
and U5567 (N_5567,N_633,N_816);
nand U5568 (N_5568,N_1996,N_2196);
or U5569 (N_5569,N_1015,N_703);
nor U5570 (N_5570,N_1568,N_2126);
or U5571 (N_5571,N_1693,N_523);
nor U5572 (N_5572,N_2259,N_1622);
xor U5573 (N_5573,N_953,N_34);
or U5574 (N_5574,N_2091,N_2133);
and U5575 (N_5575,N_1034,N_2787);
nor U5576 (N_5576,N_2368,N_1401);
xor U5577 (N_5577,N_1443,N_1096);
nand U5578 (N_5578,N_645,N_261);
and U5579 (N_5579,N_419,N_230);
or U5580 (N_5580,N_1890,N_423);
nor U5581 (N_5581,N_162,N_1012);
nor U5582 (N_5582,N_1839,N_1327);
nand U5583 (N_5583,N_2485,N_123);
nor U5584 (N_5584,N_2423,N_2768);
nand U5585 (N_5585,N_28,N_2881);
and U5586 (N_5586,N_1764,N_327);
or U5587 (N_5587,N_1322,N_952);
nor U5588 (N_5588,N_41,N_908);
or U5589 (N_5589,N_1729,N_2459);
nand U5590 (N_5590,N_2299,N_2214);
xor U5591 (N_5591,N_162,N_27);
and U5592 (N_5592,N_2955,N_1315);
or U5593 (N_5593,N_649,N_506);
or U5594 (N_5594,N_1777,N_2793);
and U5595 (N_5595,N_496,N_2420);
nand U5596 (N_5596,N_2801,N_1442);
and U5597 (N_5597,N_205,N_447);
nand U5598 (N_5598,N_1848,N_1873);
nor U5599 (N_5599,N_2530,N_1049);
nand U5600 (N_5600,N_1566,N_2079);
nand U5601 (N_5601,N_2301,N_1439);
nor U5602 (N_5602,N_2707,N_2284);
and U5603 (N_5603,N_137,N_619);
nand U5604 (N_5604,N_323,N_324);
and U5605 (N_5605,N_624,N_401);
nand U5606 (N_5606,N_881,N_753);
or U5607 (N_5607,N_51,N_343);
nor U5608 (N_5608,N_528,N_2064);
nand U5609 (N_5609,N_983,N_1352);
nor U5610 (N_5610,N_2450,N_2836);
nor U5611 (N_5611,N_2205,N_2959);
nor U5612 (N_5612,N_2675,N_2937);
nor U5613 (N_5613,N_397,N_275);
nor U5614 (N_5614,N_1426,N_2247);
nand U5615 (N_5615,N_2250,N_2671);
nor U5616 (N_5616,N_220,N_1761);
nand U5617 (N_5617,N_996,N_1578);
nand U5618 (N_5618,N_2308,N_1386);
nor U5619 (N_5619,N_859,N_688);
or U5620 (N_5620,N_1588,N_2336);
and U5621 (N_5621,N_1245,N_1803);
or U5622 (N_5622,N_1475,N_1193);
or U5623 (N_5623,N_807,N_2290);
or U5624 (N_5624,N_1182,N_246);
nor U5625 (N_5625,N_991,N_1635);
and U5626 (N_5626,N_1579,N_74);
and U5627 (N_5627,N_1314,N_2051);
and U5628 (N_5628,N_2560,N_375);
and U5629 (N_5629,N_2708,N_577);
nand U5630 (N_5630,N_1991,N_500);
and U5631 (N_5631,N_2837,N_1870);
or U5632 (N_5632,N_1686,N_1056);
and U5633 (N_5633,N_300,N_539);
xnor U5634 (N_5634,N_530,N_2286);
and U5635 (N_5635,N_1802,N_1885);
nand U5636 (N_5636,N_1275,N_1154);
xnor U5637 (N_5637,N_2429,N_1784);
and U5638 (N_5638,N_2304,N_541);
or U5639 (N_5639,N_1869,N_92);
and U5640 (N_5640,N_2163,N_577);
nand U5641 (N_5641,N_1249,N_1419);
nand U5642 (N_5642,N_1639,N_1559);
xnor U5643 (N_5643,N_2841,N_1745);
nor U5644 (N_5644,N_2392,N_2907);
and U5645 (N_5645,N_387,N_1107);
or U5646 (N_5646,N_1830,N_1913);
or U5647 (N_5647,N_2058,N_2468);
or U5648 (N_5648,N_834,N_2699);
nor U5649 (N_5649,N_1555,N_2301);
and U5650 (N_5650,N_1389,N_2692);
nor U5651 (N_5651,N_1456,N_403);
nor U5652 (N_5652,N_2965,N_2330);
and U5653 (N_5653,N_86,N_2981);
nand U5654 (N_5654,N_487,N_90);
nor U5655 (N_5655,N_1334,N_894);
or U5656 (N_5656,N_1715,N_1641);
nand U5657 (N_5657,N_903,N_346);
nand U5658 (N_5658,N_2736,N_1973);
or U5659 (N_5659,N_1360,N_91);
or U5660 (N_5660,N_2885,N_1723);
nand U5661 (N_5661,N_2899,N_2623);
and U5662 (N_5662,N_358,N_2530);
nor U5663 (N_5663,N_1180,N_1895);
nand U5664 (N_5664,N_2304,N_1410);
xnor U5665 (N_5665,N_2059,N_1014);
and U5666 (N_5666,N_2190,N_1206);
nor U5667 (N_5667,N_1682,N_2908);
or U5668 (N_5668,N_407,N_741);
nor U5669 (N_5669,N_918,N_356);
nor U5670 (N_5670,N_265,N_488);
nor U5671 (N_5671,N_1513,N_2971);
or U5672 (N_5672,N_2158,N_162);
nor U5673 (N_5673,N_2,N_1329);
nand U5674 (N_5674,N_1944,N_2367);
nand U5675 (N_5675,N_293,N_878);
nand U5676 (N_5676,N_2820,N_1405);
nand U5677 (N_5677,N_1458,N_1135);
nor U5678 (N_5678,N_200,N_322);
and U5679 (N_5679,N_211,N_2728);
or U5680 (N_5680,N_744,N_736);
or U5681 (N_5681,N_815,N_2498);
or U5682 (N_5682,N_2602,N_948);
nand U5683 (N_5683,N_2640,N_2566);
and U5684 (N_5684,N_2240,N_639);
nor U5685 (N_5685,N_1132,N_727);
or U5686 (N_5686,N_2666,N_1362);
or U5687 (N_5687,N_17,N_2187);
and U5688 (N_5688,N_2347,N_2997);
nand U5689 (N_5689,N_468,N_2864);
nand U5690 (N_5690,N_1673,N_786);
or U5691 (N_5691,N_2601,N_2223);
or U5692 (N_5692,N_863,N_2081);
and U5693 (N_5693,N_1935,N_2016);
or U5694 (N_5694,N_2772,N_2921);
nor U5695 (N_5695,N_1588,N_634);
nand U5696 (N_5696,N_686,N_1288);
or U5697 (N_5697,N_2201,N_702);
or U5698 (N_5698,N_2566,N_1653);
or U5699 (N_5699,N_1326,N_1665);
nor U5700 (N_5700,N_214,N_2292);
or U5701 (N_5701,N_2390,N_1796);
nor U5702 (N_5702,N_2217,N_1012);
and U5703 (N_5703,N_73,N_1099);
or U5704 (N_5704,N_1599,N_2258);
nor U5705 (N_5705,N_1576,N_1844);
nand U5706 (N_5706,N_141,N_915);
nand U5707 (N_5707,N_1753,N_2314);
nand U5708 (N_5708,N_1096,N_1014);
or U5709 (N_5709,N_804,N_1021);
or U5710 (N_5710,N_2569,N_342);
or U5711 (N_5711,N_2216,N_2530);
and U5712 (N_5712,N_2638,N_923);
nor U5713 (N_5713,N_347,N_2947);
and U5714 (N_5714,N_2708,N_359);
or U5715 (N_5715,N_2705,N_958);
or U5716 (N_5716,N_1089,N_2792);
or U5717 (N_5717,N_2419,N_2498);
nor U5718 (N_5718,N_1194,N_2591);
or U5719 (N_5719,N_1187,N_659);
nor U5720 (N_5720,N_2136,N_1357);
nand U5721 (N_5721,N_2073,N_2513);
nand U5722 (N_5722,N_129,N_358);
nand U5723 (N_5723,N_2741,N_1565);
nor U5724 (N_5724,N_2783,N_575);
nand U5725 (N_5725,N_1728,N_346);
and U5726 (N_5726,N_601,N_2248);
nand U5727 (N_5727,N_1761,N_2292);
xnor U5728 (N_5728,N_1103,N_2507);
or U5729 (N_5729,N_2876,N_2878);
nand U5730 (N_5730,N_1226,N_2453);
or U5731 (N_5731,N_2251,N_288);
and U5732 (N_5732,N_966,N_1298);
and U5733 (N_5733,N_1036,N_2630);
nor U5734 (N_5734,N_550,N_2205);
or U5735 (N_5735,N_2812,N_749);
nor U5736 (N_5736,N_657,N_2122);
or U5737 (N_5737,N_278,N_2419);
and U5738 (N_5738,N_2616,N_2003);
or U5739 (N_5739,N_836,N_1529);
nand U5740 (N_5740,N_2068,N_1907);
and U5741 (N_5741,N_2959,N_2931);
nand U5742 (N_5742,N_1438,N_2682);
nor U5743 (N_5743,N_2669,N_772);
xor U5744 (N_5744,N_1335,N_229);
nand U5745 (N_5745,N_422,N_1764);
and U5746 (N_5746,N_227,N_1133);
and U5747 (N_5747,N_672,N_2764);
nor U5748 (N_5748,N_1331,N_2595);
or U5749 (N_5749,N_871,N_1252);
nor U5750 (N_5750,N_1813,N_608);
nand U5751 (N_5751,N_68,N_460);
and U5752 (N_5752,N_1745,N_421);
or U5753 (N_5753,N_222,N_2390);
nand U5754 (N_5754,N_1856,N_2458);
nor U5755 (N_5755,N_1898,N_1959);
nand U5756 (N_5756,N_126,N_73);
or U5757 (N_5757,N_449,N_428);
or U5758 (N_5758,N_2420,N_1565);
nand U5759 (N_5759,N_2089,N_1652);
nor U5760 (N_5760,N_93,N_2600);
or U5761 (N_5761,N_616,N_1077);
nor U5762 (N_5762,N_2399,N_2947);
nor U5763 (N_5763,N_1836,N_2884);
or U5764 (N_5764,N_1045,N_1418);
nand U5765 (N_5765,N_1746,N_1943);
nand U5766 (N_5766,N_1571,N_1720);
or U5767 (N_5767,N_1432,N_1916);
nor U5768 (N_5768,N_1302,N_2857);
or U5769 (N_5769,N_1203,N_1529);
nor U5770 (N_5770,N_372,N_2277);
and U5771 (N_5771,N_994,N_784);
or U5772 (N_5772,N_1605,N_2402);
nor U5773 (N_5773,N_1329,N_761);
nand U5774 (N_5774,N_1093,N_2690);
nor U5775 (N_5775,N_53,N_2858);
nor U5776 (N_5776,N_669,N_1029);
or U5777 (N_5777,N_1210,N_2643);
nor U5778 (N_5778,N_620,N_1252);
nand U5779 (N_5779,N_2407,N_216);
nor U5780 (N_5780,N_143,N_2514);
nand U5781 (N_5781,N_493,N_1563);
or U5782 (N_5782,N_1352,N_2170);
and U5783 (N_5783,N_2510,N_2711);
and U5784 (N_5784,N_1843,N_1525);
nand U5785 (N_5785,N_1693,N_2878);
nand U5786 (N_5786,N_1380,N_449);
nand U5787 (N_5787,N_220,N_2114);
or U5788 (N_5788,N_2003,N_634);
nand U5789 (N_5789,N_222,N_2954);
nand U5790 (N_5790,N_2652,N_612);
nand U5791 (N_5791,N_1332,N_2470);
or U5792 (N_5792,N_648,N_2076);
and U5793 (N_5793,N_1163,N_1951);
and U5794 (N_5794,N_90,N_2432);
nor U5795 (N_5795,N_2060,N_2906);
nor U5796 (N_5796,N_530,N_112);
nand U5797 (N_5797,N_2942,N_1836);
or U5798 (N_5798,N_696,N_2581);
or U5799 (N_5799,N_1591,N_301);
and U5800 (N_5800,N_236,N_2371);
and U5801 (N_5801,N_2690,N_1789);
and U5802 (N_5802,N_1979,N_828);
nand U5803 (N_5803,N_1800,N_1125);
nor U5804 (N_5804,N_2063,N_375);
or U5805 (N_5805,N_2467,N_2636);
and U5806 (N_5806,N_726,N_603);
nand U5807 (N_5807,N_466,N_1526);
nor U5808 (N_5808,N_626,N_2886);
or U5809 (N_5809,N_1022,N_2460);
nand U5810 (N_5810,N_521,N_2039);
and U5811 (N_5811,N_412,N_1803);
and U5812 (N_5812,N_2181,N_863);
nand U5813 (N_5813,N_199,N_1576);
and U5814 (N_5814,N_1957,N_1993);
nand U5815 (N_5815,N_2430,N_6);
nand U5816 (N_5816,N_2430,N_1710);
nand U5817 (N_5817,N_1685,N_719);
nand U5818 (N_5818,N_590,N_23);
or U5819 (N_5819,N_2210,N_1946);
and U5820 (N_5820,N_1464,N_133);
or U5821 (N_5821,N_1199,N_2057);
nor U5822 (N_5822,N_1149,N_1219);
and U5823 (N_5823,N_102,N_699);
nor U5824 (N_5824,N_683,N_2870);
nor U5825 (N_5825,N_1096,N_2372);
nand U5826 (N_5826,N_350,N_932);
nand U5827 (N_5827,N_2342,N_772);
nand U5828 (N_5828,N_118,N_106);
nand U5829 (N_5829,N_1072,N_2135);
or U5830 (N_5830,N_1746,N_2578);
or U5831 (N_5831,N_2128,N_885);
or U5832 (N_5832,N_1786,N_615);
nor U5833 (N_5833,N_1141,N_247);
nor U5834 (N_5834,N_2317,N_1845);
or U5835 (N_5835,N_982,N_118);
xor U5836 (N_5836,N_2916,N_1405);
nor U5837 (N_5837,N_2041,N_2975);
or U5838 (N_5838,N_1133,N_975);
nand U5839 (N_5839,N_483,N_444);
or U5840 (N_5840,N_1534,N_2835);
nor U5841 (N_5841,N_1570,N_1754);
nor U5842 (N_5842,N_2645,N_954);
nand U5843 (N_5843,N_419,N_2973);
nand U5844 (N_5844,N_2756,N_2634);
nor U5845 (N_5845,N_2255,N_2164);
nor U5846 (N_5846,N_1950,N_1703);
nand U5847 (N_5847,N_1135,N_2754);
and U5848 (N_5848,N_2423,N_1249);
and U5849 (N_5849,N_631,N_2014);
nor U5850 (N_5850,N_596,N_850);
or U5851 (N_5851,N_749,N_1690);
and U5852 (N_5852,N_2713,N_2845);
or U5853 (N_5853,N_2049,N_2658);
or U5854 (N_5854,N_1925,N_1923);
xor U5855 (N_5855,N_2511,N_2386);
nor U5856 (N_5856,N_2855,N_1481);
and U5857 (N_5857,N_2301,N_1749);
nor U5858 (N_5858,N_1109,N_2621);
xnor U5859 (N_5859,N_769,N_1325);
nor U5860 (N_5860,N_874,N_1032);
and U5861 (N_5861,N_1399,N_1689);
nand U5862 (N_5862,N_2199,N_2442);
or U5863 (N_5863,N_48,N_2225);
xor U5864 (N_5864,N_359,N_1672);
nand U5865 (N_5865,N_2803,N_2232);
or U5866 (N_5866,N_1520,N_1318);
xor U5867 (N_5867,N_2103,N_2990);
nor U5868 (N_5868,N_2329,N_1297);
or U5869 (N_5869,N_1819,N_1878);
or U5870 (N_5870,N_1191,N_2170);
or U5871 (N_5871,N_669,N_1809);
nor U5872 (N_5872,N_48,N_1803);
xnor U5873 (N_5873,N_927,N_1000);
nand U5874 (N_5874,N_781,N_2283);
or U5875 (N_5875,N_648,N_459);
and U5876 (N_5876,N_1004,N_1717);
or U5877 (N_5877,N_103,N_702);
or U5878 (N_5878,N_484,N_43);
and U5879 (N_5879,N_294,N_875);
or U5880 (N_5880,N_485,N_2544);
or U5881 (N_5881,N_2902,N_2844);
nand U5882 (N_5882,N_1954,N_2);
or U5883 (N_5883,N_2280,N_1443);
nor U5884 (N_5884,N_2237,N_2116);
nor U5885 (N_5885,N_1383,N_801);
and U5886 (N_5886,N_1602,N_1341);
or U5887 (N_5887,N_1860,N_476);
and U5888 (N_5888,N_1601,N_1228);
nor U5889 (N_5889,N_2808,N_524);
or U5890 (N_5890,N_2076,N_925);
or U5891 (N_5891,N_193,N_1045);
nor U5892 (N_5892,N_1397,N_752);
nor U5893 (N_5893,N_173,N_1832);
nor U5894 (N_5894,N_2218,N_1093);
nand U5895 (N_5895,N_2092,N_272);
or U5896 (N_5896,N_522,N_2547);
or U5897 (N_5897,N_291,N_2023);
or U5898 (N_5898,N_753,N_629);
nand U5899 (N_5899,N_927,N_2634);
nand U5900 (N_5900,N_295,N_1742);
and U5901 (N_5901,N_1204,N_2941);
nor U5902 (N_5902,N_358,N_1709);
nor U5903 (N_5903,N_2260,N_2089);
nor U5904 (N_5904,N_1165,N_2957);
nor U5905 (N_5905,N_2732,N_954);
nor U5906 (N_5906,N_554,N_930);
nand U5907 (N_5907,N_1293,N_1018);
nor U5908 (N_5908,N_2704,N_1473);
nor U5909 (N_5909,N_379,N_403);
nor U5910 (N_5910,N_2814,N_1792);
xnor U5911 (N_5911,N_1120,N_1081);
nand U5912 (N_5912,N_1739,N_2886);
nand U5913 (N_5913,N_1518,N_1895);
nor U5914 (N_5914,N_1268,N_1937);
or U5915 (N_5915,N_84,N_940);
and U5916 (N_5916,N_200,N_1018);
nor U5917 (N_5917,N_147,N_337);
nor U5918 (N_5918,N_1137,N_23);
nand U5919 (N_5919,N_34,N_1052);
and U5920 (N_5920,N_1843,N_829);
or U5921 (N_5921,N_607,N_1375);
and U5922 (N_5922,N_1086,N_1980);
and U5923 (N_5923,N_188,N_2777);
nor U5924 (N_5924,N_1620,N_1330);
nand U5925 (N_5925,N_2366,N_2130);
and U5926 (N_5926,N_109,N_1337);
xnor U5927 (N_5927,N_1219,N_211);
or U5928 (N_5928,N_605,N_158);
nor U5929 (N_5929,N_57,N_2155);
nor U5930 (N_5930,N_2932,N_655);
nor U5931 (N_5931,N_450,N_2039);
nor U5932 (N_5932,N_2385,N_181);
nand U5933 (N_5933,N_2943,N_2370);
nor U5934 (N_5934,N_2403,N_711);
and U5935 (N_5935,N_2732,N_366);
nor U5936 (N_5936,N_520,N_1682);
nand U5937 (N_5937,N_531,N_3);
nor U5938 (N_5938,N_1238,N_2600);
or U5939 (N_5939,N_208,N_1998);
and U5940 (N_5940,N_339,N_69);
nand U5941 (N_5941,N_23,N_1997);
or U5942 (N_5942,N_2231,N_772);
nor U5943 (N_5943,N_460,N_2212);
nand U5944 (N_5944,N_1952,N_454);
or U5945 (N_5945,N_148,N_1238);
or U5946 (N_5946,N_2312,N_902);
and U5947 (N_5947,N_1042,N_1651);
or U5948 (N_5948,N_2010,N_2349);
nand U5949 (N_5949,N_2946,N_734);
or U5950 (N_5950,N_607,N_2602);
xor U5951 (N_5951,N_2481,N_2937);
nor U5952 (N_5952,N_750,N_525);
nand U5953 (N_5953,N_831,N_2629);
or U5954 (N_5954,N_2888,N_894);
xor U5955 (N_5955,N_1260,N_1280);
and U5956 (N_5956,N_1316,N_163);
or U5957 (N_5957,N_2865,N_2536);
nand U5958 (N_5958,N_2456,N_2625);
nor U5959 (N_5959,N_2694,N_2714);
nor U5960 (N_5960,N_2615,N_960);
or U5961 (N_5961,N_1392,N_1701);
nand U5962 (N_5962,N_1621,N_2953);
nor U5963 (N_5963,N_1437,N_2143);
nand U5964 (N_5964,N_1658,N_561);
or U5965 (N_5965,N_1104,N_2198);
or U5966 (N_5966,N_2376,N_33);
nand U5967 (N_5967,N_2533,N_2959);
and U5968 (N_5968,N_2393,N_2707);
nand U5969 (N_5969,N_940,N_828);
nand U5970 (N_5970,N_2326,N_2888);
nor U5971 (N_5971,N_148,N_2330);
and U5972 (N_5972,N_115,N_1905);
nand U5973 (N_5973,N_2011,N_1565);
or U5974 (N_5974,N_1087,N_963);
or U5975 (N_5975,N_1411,N_284);
and U5976 (N_5976,N_105,N_481);
nor U5977 (N_5977,N_1760,N_1384);
nor U5978 (N_5978,N_2656,N_2286);
nor U5979 (N_5979,N_277,N_2822);
nand U5980 (N_5980,N_346,N_1765);
or U5981 (N_5981,N_535,N_636);
or U5982 (N_5982,N_542,N_1696);
nand U5983 (N_5983,N_1112,N_2103);
and U5984 (N_5984,N_2093,N_1470);
xnor U5985 (N_5985,N_2538,N_1490);
and U5986 (N_5986,N_1503,N_2068);
and U5987 (N_5987,N_748,N_2162);
nand U5988 (N_5988,N_1589,N_357);
nand U5989 (N_5989,N_271,N_737);
and U5990 (N_5990,N_1763,N_1056);
nor U5991 (N_5991,N_2746,N_144);
nor U5992 (N_5992,N_1391,N_286);
and U5993 (N_5993,N_2827,N_1534);
or U5994 (N_5994,N_1974,N_1844);
nor U5995 (N_5995,N_797,N_1167);
and U5996 (N_5996,N_2551,N_2014);
and U5997 (N_5997,N_2879,N_2818);
nand U5998 (N_5998,N_673,N_1878);
nor U5999 (N_5999,N_2731,N_2494);
and U6000 (N_6000,N_4880,N_5036);
nor U6001 (N_6001,N_3792,N_3890);
nand U6002 (N_6002,N_3615,N_5021);
nor U6003 (N_6003,N_5913,N_4676);
or U6004 (N_6004,N_3800,N_4619);
and U6005 (N_6005,N_4855,N_3225);
or U6006 (N_6006,N_5956,N_3494);
and U6007 (N_6007,N_3435,N_5899);
nand U6008 (N_6008,N_5345,N_5249);
or U6009 (N_6009,N_4284,N_4344);
nor U6010 (N_6010,N_3720,N_3399);
or U6011 (N_6011,N_3819,N_4446);
nor U6012 (N_6012,N_4348,N_4399);
nand U6013 (N_6013,N_4701,N_3981);
nor U6014 (N_6014,N_3026,N_5178);
nand U6015 (N_6015,N_5033,N_3319);
and U6016 (N_6016,N_4991,N_5675);
xor U6017 (N_6017,N_5644,N_5415);
and U6018 (N_6018,N_3680,N_4747);
xor U6019 (N_6019,N_5313,N_4064);
nand U6020 (N_6020,N_5383,N_4174);
nand U6021 (N_6021,N_5124,N_5615);
and U6022 (N_6022,N_4459,N_3577);
or U6023 (N_6023,N_5564,N_5301);
nand U6024 (N_6024,N_3022,N_4390);
nand U6025 (N_6025,N_3484,N_4552);
or U6026 (N_6026,N_3357,N_3204);
or U6027 (N_6027,N_4292,N_4997);
and U6028 (N_6028,N_5584,N_3360);
nand U6029 (N_6029,N_3491,N_5820);
or U6030 (N_6030,N_3813,N_4389);
nand U6031 (N_6031,N_5420,N_4048);
nor U6032 (N_6032,N_4050,N_3700);
nor U6033 (N_6033,N_3596,N_3305);
xor U6034 (N_6034,N_4498,N_5869);
nor U6035 (N_6035,N_5575,N_4103);
nand U6036 (N_6036,N_5507,N_5755);
nand U6037 (N_6037,N_4758,N_3730);
nor U6038 (N_6038,N_5333,N_5695);
nor U6039 (N_6039,N_5825,N_5491);
nor U6040 (N_6040,N_3231,N_5561);
and U6041 (N_6041,N_3387,N_5327);
and U6042 (N_6042,N_5375,N_5960);
or U6043 (N_6043,N_4753,N_4748);
nor U6044 (N_6044,N_4232,N_4071);
nor U6045 (N_6045,N_5851,N_3843);
and U6046 (N_6046,N_5012,N_4208);
and U6047 (N_6047,N_4806,N_3628);
xnor U6048 (N_6048,N_5321,N_3308);
nor U6049 (N_6049,N_4236,N_4728);
nand U6050 (N_6050,N_4388,N_3546);
and U6051 (N_6051,N_3595,N_3023);
nor U6052 (N_6052,N_4745,N_3649);
nand U6053 (N_6053,N_4912,N_5076);
and U6054 (N_6054,N_4260,N_4702);
or U6055 (N_6055,N_4072,N_4562);
or U6056 (N_6056,N_4206,N_5132);
nor U6057 (N_6057,N_5798,N_5019);
and U6058 (N_6058,N_4682,N_3573);
nand U6059 (N_6059,N_3108,N_3073);
or U6060 (N_6060,N_5216,N_3802);
nand U6061 (N_6061,N_5891,N_5051);
nor U6062 (N_6062,N_3423,N_4909);
nand U6063 (N_6063,N_5055,N_3531);
nand U6064 (N_6064,N_3449,N_5933);
nand U6065 (N_6065,N_5112,N_5119);
and U6066 (N_6066,N_5719,N_4804);
and U6067 (N_6067,N_4386,N_5058);
nor U6068 (N_6068,N_3529,N_5640);
or U6069 (N_6069,N_3816,N_4622);
nand U6070 (N_6070,N_5867,N_4955);
nand U6071 (N_6071,N_3236,N_5264);
or U6072 (N_6072,N_4125,N_3696);
or U6073 (N_6073,N_5560,N_3911);
nor U6074 (N_6074,N_4861,N_5011);
xor U6075 (N_6075,N_4707,N_4913);
and U6076 (N_6076,N_3099,N_3294);
xnor U6077 (N_6077,N_4863,N_4918);
nand U6078 (N_6078,N_4587,N_4944);
nand U6079 (N_6079,N_4611,N_5905);
or U6080 (N_6080,N_4014,N_3874);
or U6081 (N_6081,N_5666,N_5031);
nor U6082 (N_6082,N_5768,N_3162);
and U6083 (N_6083,N_3672,N_4340);
or U6084 (N_6084,N_5281,N_5393);
and U6085 (N_6085,N_3187,N_4146);
or U6086 (N_6086,N_3368,N_3454);
or U6087 (N_6087,N_4249,N_3543);
nand U6088 (N_6088,N_5062,N_5654);
or U6089 (N_6089,N_5118,N_3740);
or U6090 (N_6090,N_3509,N_4590);
or U6091 (N_6091,N_3223,N_5775);
nand U6092 (N_6092,N_3989,N_4524);
nor U6093 (N_6093,N_4418,N_5919);
and U6094 (N_6094,N_4414,N_5849);
and U6095 (N_6095,N_5512,N_4180);
and U6096 (N_6096,N_4519,N_4521);
and U6097 (N_6097,N_4083,N_4835);
and U6098 (N_6098,N_3355,N_4914);
nor U6099 (N_6099,N_4948,N_4550);
and U6100 (N_6100,N_5590,N_4999);
or U6101 (N_6101,N_5680,N_3642);
nor U6102 (N_6102,N_3971,N_3378);
nor U6103 (N_6103,N_5063,N_5910);
or U6104 (N_6104,N_4279,N_5045);
nor U6105 (N_6105,N_5066,N_3041);
or U6106 (N_6106,N_5211,N_4150);
nor U6107 (N_6107,N_5160,N_5609);
nand U6108 (N_6108,N_4520,N_4966);
nor U6109 (N_6109,N_3967,N_5370);
nor U6110 (N_6110,N_3520,N_5110);
or U6111 (N_6111,N_3882,N_5284);
and U6112 (N_6112,N_3806,N_4423);
and U6113 (N_6113,N_3128,N_5901);
nand U6114 (N_6114,N_3548,N_4842);
nor U6115 (N_6115,N_3519,N_5291);
and U6116 (N_6116,N_5462,N_4652);
and U6117 (N_6117,N_5734,N_5490);
and U6118 (N_6118,N_5607,N_4043);
nor U6119 (N_6119,N_3171,N_5368);
nor U6120 (N_6120,N_3182,N_4924);
or U6121 (N_6121,N_4987,N_4537);
and U6122 (N_6122,N_5835,N_4427);
or U6123 (N_6123,N_4343,N_4668);
xnor U6124 (N_6124,N_4685,N_4518);
and U6125 (N_6125,N_4073,N_5109);
nor U6126 (N_6126,N_5423,N_5679);
nor U6127 (N_6127,N_4410,N_3147);
nand U6128 (N_6128,N_4588,N_3918);
and U6129 (N_6129,N_4528,N_5971);
or U6130 (N_6130,N_3149,N_3785);
or U6131 (N_6131,N_5535,N_4505);
nand U6132 (N_6132,N_4516,N_4038);
and U6133 (N_6133,N_5625,N_5060);
nor U6134 (N_6134,N_3310,N_4396);
and U6135 (N_6135,N_3951,N_5986);
nand U6136 (N_6136,N_4679,N_3893);
and U6137 (N_6137,N_5214,N_4886);
nand U6138 (N_6138,N_5141,N_5907);
nand U6139 (N_6139,N_4998,N_3561);
nand U6140 (N_6140,N_3823,N_3324);
nand U6141 (N_6141,N_3719,N_3228);
or U6142 (N_6142,N_5107,N_4198);
and U6143 (N_6143,N_5510,N_4456);
nand U6144 (N_6144,N_3748,N_5702);
nand U6145 (N_6145,N_3196,N_3239);
or U6146 (N_6146,N_5198,N_4627);
nor U6147 (N_6147,N_3943,N_5145);
and U6148 (N_6148,N_3253,N_5186);
and U6149 (N_6149,N_4434,N_4349);
or U6150 (N_6150,N_5422,N_3880);
and U6151 (N_6151,N_3928,N_3051);
nand U6152 (N_6152,N_3970,N_3944);
or U6153 (N_6153,N_3653,N_5858);
nor U6154 (N_6154,N_5877,N_3537);
and U6155 (N_6155,N_4608,N_4440);
nor U6156 (N_6156,N_4219,N_4931);
nor U6157 (N_6157,N_4959,N_4297);
nor U6158 (N_6158,N_5041,N_4579);
and U6159 (N_6159,N_4828,N_5280);
or U6160 (N_6160,N_5022,N_4052);
and U6161 (N_6161,N_3973,N_3629);
or U6162 (N_6162,N_4098,N_5880);
nor U6163 (N_6163,N_4658,N_4022);
or U6164 (N_6164,N_4650,N_3156);
nor U6165 (N_6165,N_5992,N_3503);
or U6166 (N_6166,N_5928,N_3047);
nand U6167 (N_6167,N_3058,N_5606);
or U6168 (N_6168,N_5771,N_5085);
nor U6169 (N_6169,N_3431,N_5073);
nor U6170 (N_6170,N_4877,N_5233);
nor U6171 (N_6171,N_3042,N_3082);
nor U6172 (N_6172,N_5424,N_4294);
nor U6173 (N_6173,N_4323,N_4178);
or U6174 (N_6174,N_5830,N_5528);
nor U6175 (N_6175,N_5935,N_5317);
nand U6176 (N_6176,N_3814,N_3780);
nand U6177 (N_6177,N_5452,N_4218);
nand U6178 (N_6178,N_3832,N_3158);
nor U6179 (N_6179,N_4547,N_4827);
or U6180 (N_6180,N_3822,N_5075);
and U6181 (N_6181,N_3933,N_4181);
or U6182 (N_6182,N_3617,N_5430);
nand U6183 (N_6183,N_4559,N_4350);
or U6184 (N_6184,N_4517,N_4534);
and U6185 (N_6185,N_4599,N_5900);
or U6186 (N_6186,N_4648,N_4223);
nor U6187 (N_6187,N_4803,N_5427);
nand U6188 (N_6188,N_5797,N_5187);
and U6189 (N_6189,N_3066,N_4781);
nor U6190 (N_6190,N_4357,N_4193);
and U6191 (N_6191,N_3424,N_5217);
or U6192 (N_6192,N_3110,N_5572);
nand U6193 (N_6193,N_5256,N_3927);
and U6194 (N_6194,N_5213,N_5508);
or U6195 (N_6195,N_4846,N_4560);
or U6196 (N_6196,N_5436,N_4354);
or U6197 (N_6197,N_5026,N_3350);
nor U6198 (N_6198,N_4976,N_4871);
and U6199 (N_6199,N_3276,N_3601);
nand U6200 (N_6200,N_4603,N_5769);
nand U6201 (N_6201,N_5359,N_4908);
nand U6202 (N_6202,N_3952,N_4610);
xor U6203 (N_6203,N_4556,N_4761);
and U6204 (N_6204,N_4080,N_3351);
nor U6205 (N_6205,N_5738,N_4017);
or U6206 (N_6206,N_4653,N_3311);
nand U6207 (N_6207,N_4383,N_3554);
and U6208 (N_6208,N_5384,N_4175);
nor U6209 (N_6209,N_4958,N_4123);
or U6210 (N_6210,N_5509,N_4536);
nor U6211 (N_6211,N_5040,N_4407);
nand U6212 (N_6212,N_5319,N_4813);
nor U6213 (N_6213,N_5613,N_5114);
nor U6214 (N_6214,N_4647,N_5276);
and U6215 (N_6215,N_4420,N_4903);
or U6216 (N_6216,N_3032,N_5895);
and U6217 (N_6217,N_3133,N_3039);
nand U6218 (N_6218,N_5067,N_5565);
nor U6219 (N_6219,N_3797,N_3815);
nor U6220 (N_6220,N_3398,N_4093);
or U6221 (N_6221,N_4030,N_5599);
or U6222 (N_6222,N_5294,N_4309);
and U6223 (N_6223,N_4172,N_5721);
nand U6224 (N_6224,N_4584,N_4697);
or U6225 (N_6225,N_3328,N_3272);
and U6226 (N_6226,N_3244,N_3539);
xor U6227 (N_6227,N_4024,N_4283);
and U6228 (N_6228,N_4878,N_5586);
or U6229 (N_6229,N_4811,N_5405);
or U6230 (N_6230,N_4027,N_4122);
and U6231 (N_6231,N_3549,N_5378);
nor U6232 (N_6232,N_4896,N_5224);
nor U6233 (N_6233,N_5275,N_3791);
nand U6234 (N_6234,N_3768,N_5887);
and U6235 (N_6235,N_4392,N_5172);
or U6236 (N_6236,N_5543,N_5581);
or U6237 (N_6237,N_3869,N_5837);
nor U6238 (N_6238,N_4327,N_3480);
and U6239 (N_6239,N_4995,N_3285);
nor U6240 (N_6240,N_5697,N_5957);
or U6241 (N_6241,N_5096,N_5540);
xor U6242 (N_6242,N_5763,N_3887);
nand U6243 (N_6243,N_4034,N_3312);
and U6244 (N_6244,N_4960,N_3591);
and U6245 (N_6245,N_3116,N_5161);
nor U6246 (N_6246,N_3662,N_3979);
nand U6247 (N_6247,N_5857,N_4177);
nand U6248 (N_6248,N_3313,N_3137);
and U6249 (N_6249,N_3950,N_5008);
and U6250 (N_6250,N_4594,N_5013);
nor U6251 (N_6251,N_4969,N_3482);
nand U6252 (N_6252,N_5637,N_5757);
nand U6253 (N_6253,N_3930,N_5329);
or U6254 (N_6254,N_5652,N_3232);
nand U6255 (N_6255,N_4737,N_5821);
nor U6256 (N_6256,N_4214,N_5382);
nand U6257 (N_6257,N_3264,N_5533);
nand U6258 (N_6258,N_5875,N_4629);
nor U6259 (N_6259,N_4502,N_3870);
nor U6260 (N_6260,N_5188,N_3582);
or U6261 (N_6261,N_5944,N_4130);
and U6262 (N_6262,N_3361,N_3624);
or U6263 (N_6263,N_5443,N_5046);
and U6264 (N_6264,N_3417,N_3220);
nor U6265 (N_6265,N_5770,N_3931);
xor U6266 (N_6266,N_4710,N_4290);
nor U6267 (N_6267,N_3980,N_3863);
and U6268 (N_6268,N_3851,N_3160);
or U6269 (N_6269,N_5277,N_4503);
xor U6270 (N_6270,N_4540,N_4137);
and U6271 (N_6271,N_5983,N_4089);
nand U6272 (N_6272,N_4090,N_3540);
nor U6273 (N_6273,N_3117,N_3325);
nand U6274 (N_6274,N_3884,N_5774);
nor U6275 (N_6275,N_4962,N_5271);
nor U6276 (N_6276,N_4194,N_5180);
and U6277 (N_6277,N_4621,N_5628);
and U6278 (N_6278,N_4894,N_3080);
and U6279 (N_6279,N_5461,N_5673);
nor U6280 (N_6280,N_3407,N_5408);
nand U6281 (N_6281,N_5658,N_3044);
nor U6282 (N_6282,N_3912,N_4437);
nand U6283 (N_6283,N_4041,N_3640);
and U6284 (N_6284,N_4287,N_4779);
and U6285 (N_6285,N_3966,N_4527);
nand U6286 (N_6286,N_4453,N_3450);
and U6287 (N_6287,N_5671,N_5121);
or U6288 (N_6288,N_4809,N_3523);
xnor U6289 (N_6289,N_5446,N_5065);
and U6290 (N_6290,N_4170,N_4363);
nor U6291 (N_6291,N_3567,N_4149);
and U6292 (N_6292,N_5215,N_4495);
nand U6293 (N_6293,N_5845,N_5634);
nor U6294 (N_6294,N_4443,N_5521);
and U6295 (N_6295,N_4321,N_5197);
and U6296 (N_6296,N_5890,N_5125);
nor U6297 (N_6297,N_4585,N_5647);
or U6298 (N_6298,N_5164,N_3152);
and U6299 (N_6299,N_3704,N_4639);
nor U6300 (N_6300,N_5137,N_5764);
nor U6301 (N_6301,N_3476,N_5136);
nor U6302 (N_6302,N_5113,N_5292);
nand U6303 (N_6303,N_3899,N_5678);
or U6304 (N_6304,N_3607,N_4810);
nand U6305 (N_6305,N_4266,N_4649);
and U6306 (N_6306,N_5357,N_3692);
and U6307 (N_6307,N_5082,N_5266);
nand U6308 (N_6308,N_3521,N_4142);
and U6309 (N_6309,N_3306,N_4815);
nand U6310 (N_6310,N_3530,N_3825);
nand U6311 (N_6311,N_3203,N_5142);
nor U6312 (N_6312,N_5632,N_3467);
nand U6313 (N_6313,N_4651,N_5482);
xor U6314 (N_6314,N_4830,N_4672);
nor U6315 (N_6315,N_5143,N_4841);
and U6316 (N_6316,N_3637,N_3910);
nor U6317 (N_6317,N_4765,N_4139);
or U6318 (N_6318,N_5953,N_5873);
nand U6319 (N_6319,N_4738,N_5445);
nor U6320 (N_6320,N_5601,N_3742);
nor U6321 (N_6321,N_5318,N_5513);
nor U6322 (N_6322,N_3600,N_5230);
or U6323 (N_6323,N_4952,N_3217);
and U6324 (N_6324,N_3292,N_4016);
nand U6325 (N_6325,N_3769,N_5963);
xor U6326 (N_6326,N_5871,N_4107);
or U6327 (N_6327,N_4526,N_4417);
and U6328 (N_6328,N_3716,N_5544);
nor U6329 (N_6329,N_3677,N_4636);
nand U6330 (N_6330,N_3382,N_5348);
or U6331 (N_6331,N_4581,N_5103);
and U6332 (N_6332,N_5812,N_3273);
nand U6333 (N_6333,N_5573,N_4342);
and U6334 (N_6334,N_3248,N_5629);
and U6335 (N_6335,N_3396,N_3060);
and U6336 (N_6336,N_5816,N_3773);
and U6337 (N_6337,N_4691,N_4138);
and U6338 (N_6338,N_5403,N_5169);
or U6339 (N_6339,N_3991,N_5638);
and U6340 (N_6340,N_4833,N_3782);
nand U6341 (N_6341,N_5688,N_5016);
and U6342 (N_6342,N_5195,N_3500);
or U6343 (N_6343,N_5725,N_3404);
nand U6344 (N_6344,N_4447,N_4703);
nor U6345 (N_6345,N_5039,N_5718);
and U6346 (N_6346,N_5807,N_5773);
and U6347 (N_6347,N_3315,N_3603);
and U6348 (N_6348,N_4654,N_5475);
nor U6349 (N_6349,N_5438,N_4352);
nand U6350 (N_6350,N_4021,N_4766);
and U6351 (N_6351,N_4325,N_4129);
nor U6352 (N_6352,N_5135,N_4431);
nand U6353 (N_6353,N_3438,N_5296);
nand U6354 (N_6354,N_4868,N_4413);
or U6355 (N_6355,N_3380,N_4244);
nand U6356 (N_6356,N_5200,N_4949);
nand U6357 (N_6357,N_4727,N_3620);
nand U6358 (N_6358,N_4449,N_3316);
or U6359 (N_6359,N_5848,N_3317);
nor U6360 (N_6360,N_4280,N_5585);
or U6361 (N_6361,N_4274,N_5054);
or U6362 (N_6362,N_4213,N_4961);
or U6363 (N_6363,N_4749,N_5795);
or U6364 (N_6364,N_4905,N_3455);
and U6365 (N_6365,N_4533,N_4785);
nor U6366 (N_6366,N_5978,N_3916);
nor U6367 (N_6367,N_5399,N_3111);
nand U6368 (N_6368,N_5068,N_5226);
or U6369 (N_6369,N_5084,N_3124);
nand U6370 (N_6370,N_3635,N_4106);
and U6371 (N_6371,N_5713,N_4971);
and U6372 (N_6372,N_4049,N_5940);
nand U6373 (N_6373,N_5150,N_3760);
nand U6374 (N_6374,N_4576,N_5733);
and U6375 (N_6375,N_4817,N_5939);
or U6376 (N_6376,N_4255,N_3437);
nor U6377 (N_6377,N_5843,N_4736);
nor U6378 (N_6378,N_4299,N_4561);
nand U6379 (N_6379,N_3820,N_3250);
nor U6380 (N_6380,N_5083,N_3447);
nor U6381 (N_6381,N_3095,N_3372);
nor U6382 (N_6382,N_4442,N_4293);
nor U6383 (N_6383,N_3440,N_4018);
nand U6384 (N_6384,N_5251,N_5456);
nand U6385 (N_6385,N_3982,N_4631);
nor U6386 (N_6386,N_3441,N_4922);
and U6387 (N_6387,N_4486,N_3934);
nand U6388 (N_6388,N_5295,N_4563);
or U6389 (N_6389,N_4009,N_4628);
and U6390 (N_6390,N_4468,N_4834);
or U6391 (N_6391,N_3593,N_5254);
nor U6392 (N_6392,N_5754,N_3353);
or U6393 (N_6393,N_4450,N_5496);
nor U6394 (N_6394,N_5554,N_3733);
and U6395 (N_6395,N_4644,N_3788);
and U6396 (N_6396,N_4539,N_3063);
and U6397 (N_6397,N_3075,N_4037);
nor U6398 (N_6398,N_5583,N_3551);
nor U6399 (N_6399,N_4775,N_3706);
nand U6400 (N_6400,N_4469,N_5874);
or U6401 (N_6401,N_5307,N_5931);
nor U6402 (N_6402,N_5672,N_3255);
nand U6403 (N_6403,N_5222,N_5884);
or U6404 (N_6404,N_4439,N_3631);
nor U6405 (N_6405,N_4932,N_3889);
or U6406 (N_6406,N_5975,N_4496);
nor U6407 (N_6407,N_3609,N_3400);
nand U6408 (N_6408,N_3610,N_4531);
nand U6409 (N_6409,N_5498,N_5947);
or U6410 (N_6410,N_3469,N_3190);
or U6411 (N_6411,N_5273,N_4699);
or U6412 (N_6412,N_5166,N_4771);
or U6413 (N_6413,N_4548,N_3138);
and U6414 (N_6414,N_5151,N_4858);
nand U6415 (N_6415,N_4336,N_5993);
nor U6416 (N_6416,N_5650,N_4215);
and U6417 (N_6417,N_4480,N_4289);
and U6418 (N_6418,N_4023,N_4514);
or U6419 (N_6419,N_5023,N_3611);
and U6420 (N_6420,N_5095,N_4015);
or U6421 (N_6421,N_3290,N_5193);
and U6422 (N_6422,N_5229,N_5147);
nor U6423 (N_6423,N_3192,N_4711);
or U6424 (N_6424,N_3411,N_3188);
and U6425 (N_6425,N_3794,N_4378);
nand U6426 (N_6426,N_5704,N_4782);
nor U6427 (N_6427,N_3046,N_3233);
and U6428 (N_6428,N_5171,N_5645);
nor U6429 (N_6429,N_5537,N_4394);
and U6430 (N_6430,N_4572,N_4245);
or U6431 (N_6431,N_4821,N_3571);
and U6432 (N_6432,N_4147,N_4272);
xor U6433 (N_6433,N_3146,N_4867);
or U6434 (N_6434,N_3043,N_3120);
and U6435 (N_6435,N_4953,N_4360);
nand U6436 (N_6436,N_3029,N_5239);
nand U6437 (N_6437,N_5850,N_5826);
or U6438 (N_6438,N_4473,N_5322);
nand U6439 (N_6439,N_4400,N_4330);
or U6440 (N_6440,N_3459,N_3959);
nor U6441 (N_6441,N_4010,N_3925);
nor U6442 (N_6442,N_3122,N_5010);
nor U6443 (N_6443,N_3714,N_5942);
and U6444 (N_6444,N_5979,N_3402);
nor U6445 (N_6445,N_5969,N_4973);
nor U6446 (N_6446,N_3388,N_5842);
nand U6447 (N_6447,N_3256,N_5397);
nor U6448 (N_6448,N_4241,N_3365);
nor U6449 (N_6449,N_3155,N_4315);
nor U6450 (N_6450,N_5231,N_5111);
and U6451 (N_6451,N_3613,N_5819);
and U6452 (N_6452,N_3185,N_5964);
and U6453 (N_6453,N_4318,N_4543);
xnor U6454 (N_6454,N_5344,N_4509);
or U6455 (N_6455,N_3334,N_4915);
or U6456 (N_6456,N_4371,N_5449);
nand U6457 (N_6457,N_3215,N_4954);
nor U6458 (N_6458,N_3049,N_5080);
or U6459 (N_6459,N_5745,N_3344);
nand U6460 (N_6460,N_5790,N_3321);
nor U6461 (N_6461,N_3650,N_4109);
or U6462 (N_6462,N_4798,N_3105);
and U6463 (N_6463,N_3267,N_3581);
nor U6464 (N_6464,N_5471,N_3406);
or U6465 (N_6465,N_4783,N_3015);
nor U6466 (N_6466,N_4185,N_4838);
or U6467 (N_6467,N_5306,N_5911);
and U6468 (N_6468,N_5104,N_4688);
nor U6469 (N_6469,N_5473,N_4927);
and U6470 (N_6470,N_5053,N_5582);
nor U6471 (N_6471,N_4381,N_4689);
nor U6472 (N_6472,N_5888,N_5700);
or U6473 (N_6473,N_5300,N_3299);
or U6474 (N_6474,N_4092,N_4430);
or U6475 (N_6475,N_3926,N_4096);
nand U6476 (N_6476,N_5959,N_5002);
or U6477 (N_6477,N_3209,N_3987);
and U6478 (N_6478,N_4176,N_3641);
and U6479 (N_6479,N_5434,N_3142);
or U6480 (N_6480,N_3920,N_3002);
and U6481 (N_6481,N_5189,N_4425);
nor U6482 (N_6482,N_3131,N_5641);
and U6483 (N_6483,N_5199,N_4704);
nand U6484 (N_6484,N_3622,N_4899);
nand U6485 (N_6485,N_4577,N_3505);
and U6486 (N_6486,N_3818,N_4458);
nor U6487 (N_6487,N_4351,N_5432);
nand U6488 (N_6488,N_4698,N_5343);
nand U6489 (N_6489,N_5676,N_4529);
and U6490 (N_6490,N_5278,N_5201);
or U6491 (N_6491,N_5057,N_5183);
and U6492 (N_6492,N_5894,N_5932);
nor U6493 (N_6493,N_4079,N_4011);
and U6494 (N_6494,N_5868,N_4823);
nor U6495 (N_6495,N_3180,N_4724);
nand U6496 (N_6496,N_4718,N_4086);
nor U6497 (N_6497,N_4666,N_5860);
xnor U6498 (N_6498,N_4310,N_3550);
or U6499 (N_6499,N_3143,N_4714);
nor U6500 (N_6500,N_5555,N_3456);
or U6501 (N_6501,N_5780,N_5206);
and U6502 (N_6502,N_3405,N_4421);
and U6503 (N_6503,N_3102,N_3556);
nor U6504 (N_6504,N_4209,N_3140);
nand U6505 (N_6505,N_4075,N_5766);
and U6506 (N_6506,N_4586,N_4108);
nor U6507 (N_6507,N_5810,N_5389);
and U6508 (N_6508,N_4907,N_3309);
and U6509 (N_6509,N_3734,N_3830);
nor U6510 (N_6510,N_5624,N_5937);
or U6511 (N_6511,N_5973,N_4706);
nand U6512 (N_6512,N_5556,N_5392);
or U6513 (N_6513,N_4269,N_3498);
or U6514 (N_6514,N_4569,N_3961);
and U6515 (N_6515,N_3169,N_5364);
and U6516 (N_6516,N_4984,N_5316);
and U6517 (N_6517,N_4883,N_5889);
nor U6518 (N_6518,N_3647,N_4121);
nor U6519 (N_6519,N_5488,N_3897);
and U6520 (N_6520,N_4069,N_3359);
or U6521 (N_6521,N_4893,N_4445);
nand U6522 (N_6522,N_4365,N_3875);
and U6523 (N_6523,N_4754,N_4136);
nor U6524 (N_6524,N_4433,N_5786);
nor U6525 (N_6525,N_4002,N_3369);
or U6526 (N_6526,N_5362,N_3625);
or U6527 (N_6527,N_5639,N_4339);
xor U6528 (N_6528,N_5182,N_4712);
and U6529 (N_6529,N_4379,N_3762);
and U6530 (N_6530,N_4265,N_3205);
nor U6531 (N_6531,N_5015,N_5863);
or U6532 (N_6532,N_5627,N_5374);
and U6533 (N_6533,N_3495,N_3167);
nand U6534 (N_6534,N_5325,N_5502);
and U6535 (N_6535,N_5800,N_5758);
or U6536 (N_6536,N_4790,N_5562);
nor U6537 (N_6537,N_3332,N_4491);
or U6538 (N_6538,N_3514,N_4237);
or U6539 (N_6539,N_3024,N_4723);
nand U6540 (N_6540,N_3847,N_3903);
nor U6541 (N_6541,N_4901,N_4159);
or U6542 (N_6542,N_4278,N_4930);
or U6543 (N_6543,N_5043,N_3393);
and U6544 (N_6544,N_4945,N_3774);
nor U6545 (N_6545,N_4849,N_4497);
nor U6546 (N_6546,N_4767,N_3084);
nor U6547 (N_6547,N_3094,N_4338);
or U6548 (N_6548,N_4470,N_4741);
or U6549 (N_6549,N_3811,N_5717);
or U6550 (N_6550,N_5037,N_3793);
nand U6551 (N_6551,N_5551,N_4326);
and U6552 (N_6552,N_3426,N_4462);
and U6553 (N_6553,N_4163,N_5824);
nand U6554 (N_6554,N_4929,N_5386);
nor U6555 (N_6555,N_4201,N_3079);
nor U6556 (N_6556,N_5994,N_5148);
or U6557 (N_6557,N_5709,N_5252);
nor U6558 (N_6558,N_3003,N_3483);
or U6559 (N_6559,N_3604,N_4722);
or U6560 (N_6560,N_3086,N_3681);
and U6561 (N_6561,N_5155,N_4145);
and U6562 (N_6562,N_3468,N_5728);
nor U6563 (N_6563,N_5227,N_3472);
and U6564 (N_6564,N_3807,N_5173);
nand U6565 (N_6565,N_3686,N_4268);
or U6566 (N_6566,N_4637,N_3990);
and U6567 (N_6567,N_4787,N_4906);
or U6568 (N_6568,N_3163,N_3856);
nand U6569 (N_6569,N_4385,N_5175);
nor U6570 (N_6570,N_4441,N_5866);
nand U6571 (N_6571,N_5970,N_3858);
nand U6572 (N_6572,N_3835,N_3842);
nand U6573 (N_6573,N_3141,N_5219);
xor U6574 (N_6574,N_3565,N_4670);
and U6575 (N_6575,N_4799,N_5335);
nor U6576 (N_6576,N_5377,N_4935);
and U6577 (N_6577,N_4068,N_3756);
or U6578 (N_6578,N_4974,N_3374);
and U6579 (N_6579,N_5701,N_3866);
or U6580 (N_6580,N_3885,N_3779);
nand U6581 (N_6581,N_5366,N_5355);
and U6582 (N_6582,N_4361,N_3569);
nor U6583 (N_6583,N_4696,N_5588);
nor U6584 (N_6584,N_4493,N_5149);
nor U6585 (N_6585,N_4478,N_5245);
or U6586 (N_6586,N_3287,N_3261);
or U6587 (N_6587,N_3501,N_5662);
nand U6588 (N_6588,N_4300,N_3969);
or U6589 (N_6589,N_3366,N_4544);
nor U6590 (N_6590,N_3999,N_5834);
and U6591 (N_6591,N_3988,N_4964);
nor U6592 (N_6592,N_3583,N_4380);
and U6593 (N_6593,N_4674,N_3743);
xnor U6594 (N_6594,N_4408,N_5394);
or U6595 (N_6595,N_4892,N_4965);
nand U6596 (N_6596,N_5747,N_4919);
and U6597 (N_6597,N_4763,N_3302);
nand U6598 (N_6598,N_5504,N_3729);
nand U6599 (N_6599,N_5417,N_3207);
and U6600 (N_6600,N_3178,N_3279);
nand U6601 (N_6601,N_3853,N_3542);
and U6602 (N_6602,N_3331,N_4940);
nor U6603 (N_6603,N_4832,N_3865);
nand U6604 (N_6604,N_4968,N_3293);
nand U6605 (N_6605,N_3848,N_4364);
or U6606 (N_6606,N_4731,N_5493);
and U6607 (N_6607,N_4881,N_4313);
and U6608 (N_6608,N_4542,N_3083);
nand U6609 (N_6609,N_4298,N_3172);
or U6610 (N_6610,N_3957,N_5122);
nand U6611 (N_6611,N_3247,N_4217);
nand U6612 (N_6612,N_4609,N_3845);
nor U6613 (N_6613,N_4184,N_3208);
nor U6614 (N_6614,N_5987,N_4179);
and U6615 (N_6615,N_3367,N_5838);
xnor U6616 (N_6616,N_5035,N_4690);
xor U6617 (N_6617,N_3055,N_3707);
or U6618 (N_6618,N_4680,N_5988);
or U6619 (N_6619,N_5727,N_5981);
nor U6620 (N_6620,N_5744,N_5761);
nor U6621 (N_6621,N_4405,N_4571);
or U6622 (N_6622,N_5138,N_4156);
nor U6623 (N_6623,N_3682,N_4488);
and U6624 (N_6624,N_5623,N_3941);
and U6625 (N_6625,N_4625,N_5339);
and U6626 (N_6626,N_4398,N_4140);
or U6627 (N_6627,N_5547,N_3466);
and U6628 (N_6628,N_4725,N_5401);
and U6629 (N_6629,N_4205,N_5265);
and U6630 (N_6630,N_5946,N_5440);
or U6631 (N_6631,N_3258,N_5192);
xnor U6632 (N_6632,N_5480,N_5828);
or U6633 (N_6633,N_5591,N_5395);
and U6634 (N_6634,N_3106,N_4155);
nand U6635 (N_6635,N_5270,N_4525);
or U6636 (N_6636,N_3998,N_5854);
and U6637 (N_6637,N_3206,N_5353);
nor U6638 (N_6638,N_5003,N_5024);
and U6639 (N_6639,N_3096,N_3280);
and U6640 (N_6640,N_4370,N_4665);
nand U6641 (N_6641,N_3275,N_5501);
and U6642 (N_6642,N_5739,N_5391);
and U6643 (N_6643,N_5202,N_4596);
nand U6644 (N_6644,N_5998,N_5027);
and U6645 (N_6645,N_3968,N_3129);
nor U6646 (N_6646,N_5376,N_5603);
nor U6647 (N_6647,N_4535,N_3139);
nor U6648 (N_6648,N_3775,N_5017);
or U6649 (N_6649,N_3379,N_5594);
and U6650 (N_6650,N_4059,N_5833);
xor U6651 (N_6651,N_3906,N_4800);
or U6652 (N_6652,N_3538,N_5494);
nor U6653 (N_6653,N_4291,N_4302);
nand U6654 (N_6654,N_4742,N_4947);
and U6655 (N_6655,N_3329,N_5787);
or U6656 (N_6656,N_3909,N_3744);
nand U6657 (N_6657,N_4733,N_3829);
nor U6658 (N_6658,N_4951,N_3154);
or U6659 (N_6659,N_3020,N_3009);
nand U6660 (N_6660,N_5742,N_4384);
nor U6661 (N_6661,N_3460,N_4276);
nor U6662 (N_6662,N_3303,N_5269);
nor U6663 (N_6663,N_4359,N_4675);
nor U6664 (N_6664,N_4530,N_3341);
and U6665 (N_6665,N_3453,N_3214);
and U6666 (N_6666,N_3027,N_4808);
and U6667 (N_6667,N_4891,N_4247);
and U6668 (N_6668,N_4239,N_4721);
or U6669 (N_6669,N_4864,N_4911);
and U6670 (N_6670,N_5611,N_3471);
nor U6671 (N_6671,N_4161,N_5237);
nor U6672 (N_6672,N_4258,N_3854);
or U6673 (N_6673,N_5238,N_4660);
and U6674 (N_6674,N_4492,N_5620);
nand U6675 (N_6675,N_4415,N_3960);
nor U6676 (N_6676,N_5885,N_5441);
or U6677 (N_6677,N_3975,N_4546);
and U6678 (N_6678,N_5915,N_4613);
and U6679 (N_6679,N_3668,N_5365);
nor U6680 (N_6680,N_4739,N_3691);
or U6681 (N_6681,N_3318,N_5570);
or U6682 (N_6682,N_5892,N_3001);
nand U6683 (N_6683,N_3200,N_3913);
and U6684 (N_6684,N_4663,N_3948);
or U6685 (N_6685,N_4709,N_3757);
and U6686 (N_6686,N_5893,N_3497);
nor U6687 (N_6687,N_3655,N_4195);
or U6688 (N_6688,N_4840,N_5268);
nor U6689 (N_6689,N_3462,N_5293);
nand U6690 (N_6690,N_4921,N_3241);
nor U6691 (N_6691,N_3592,N_5737);
nand U6692 (N_6692,N_4317,N_5592);
nand U6693 (N_6693,N_3761,N_3251);
and U6694 (N_6694,N_3758,N_5663);
nand U6695 (N_6695,N_4780,N_3871);
nand U6696 (N_6696,N_4481,N_4677);
and U6697 (N_6697,N_4700,N_4046);
nand U6698 (N_6698,N_3608,N_5822);
nor U6699 (N_6699,N_4889,N_3929);
nand U6700 (N_6700,N_3867,N_5660);
or U6701 (N_6701,N_4490,N_5442);
nand U6702 (N_6702,N_4693,N_3410);
nor U6703 (N_6703,N_5352,N_5435);
and U6704 (N_6704,N_3419,N_5538);
or U6705 (N_6705,N_3010,N_4183);
or U6706 (N_6706,N_4282,N_4013);
nor U6707 (N_6707,N_5479,N_3589);
and U6708 (N_6708,N_4664,N_5267);
nand U6709 (N_6709,N_4851,N_4638);
nor U6710 (N_6710,N_3803,N_4204);
or U6711 (N_6711,N_3463,N_4522);
or U6712 (N_6712,N_5476,N_4487);
and U6713 (N_6713,N_3457,N_5954);
and U6714 (N_6714,N_5949,N_3715);
and U6715 (N_6715,N_5859,N_5205);
nor U6716 (N_6716,N_4601,N_3654);
nor U6717 (N_6717,N_5589,N_3183);
nor U6718 (N_6718,N_4252,N_4684);
nand U6719 (N_6719,N_5428,N_4243);
or U6720 (N_6720,N_3900,N_4512);
nand U6721 (N_6721,N_5466,N_5878);
nor U6722 (N_6722,N_4012,N_3738);
nand U6723 (N_6723,N_3487,N_5534);
and U6724 (N_6724,N_3614,N_3661);
or U6725 (N_6725,N_5996,N_5668);
and U6726 (N_6726,N_3211,N_5478);
nor U6727 (N_6727,N_5714,N_5861);
or U6728 (N_6728,N_4824,N_4845);
nor U6729 (N_6729,N_3186,N_4157);
nor U6730 (N_6730,N_4314,N_5552);
nand U6731 (N_6731,N_5130,N_5710);
nand U6732 (N_6732,N_5303,N_4331);
and U6733 (N_6733,N_4006,N_4740);
nor U6734 (N_6734,N_5741,N_5283);
xor U6735 (N_6735,N_5792,N_4101);
nand U6736 (N_6736,N_4566,N_5788);
and U6737 (N_6737,N_5363,N_3701);
xnor U6738 (N_6738,N_5324,N_5789);
nor U6739 (N_6739,N_5091,N_3174);
nand U6740 (N_6740,N_4567,N_5917);
nand U6741 (N_6741,N_3274,N_4412);
and U6742 (N_6742,N_5157,N_5681);
nor U6743 (N_6743,N_5736,N_3088);
nand U6744 (N_6744,N_5579,N_5451);
and U6745 (N_6745,N_3336,N_3346);
nand U6746 (N_6746,N_5261,N_4859);
or U6747 (N_6747,N_3291,N_3731);
or U6748 (N_6748,N_3089,N_4866);
nor U6749 (N_6749,N_3709,N_5000);
nand U6750 (N_6750,N_5659,N_3876);
and U6751 (N_6751,N_3844,N_3978);
nor U6752 (N_6752,N_4791,N_5914);
nand U6753 (N_6753,N_4882,N_4085);
or U6754 (N_6754,N_4328,N_3559);
and U6755 (N_6755,N_3741,N_3667);
and U6756 (N_6756,N_3846,N_4646);
and U6757 (N_6757,N_3132,N_3808);
and U6758 (N_6758,N_5315,N_3937);
nand U6759 (N_6759,N_3562,N_4257);
and U6760 (N_6760,N_4655,N_4132);
or U6761 (N_6761,N_5548,N_5686);
nand U6762 (N_6762,N_5367,N_3659);
nand U6763 (N_6763,N_5760,N_3511);
nor U6764 (N_6764,N_5328,N_3218);
nor U6765 (N_6765,N_5783,N_5087);
and U6766 (N_6766,N_5791,N_4117);
nor U6767 (N_6767,N_4678,N_5703);
and U6768 (N_6768,N_4554,N_5934);
nand U6769 (N_6769,N_3636,N_4029);
nor U6770 (N_6770,N_4077,N_4403);
and U6771 (N_6771,N_5077,N_4203);
nand U6772 (N_6772,N_4067,N_3330);
or U6773 (N_6773,N_5373,N_4938);
nand U6774 (N_6774,N_5730,N_4375);
or U6775 (N_6775,N_4411,N_5839);
nand U6776 (N_6776,N_5938,N_3427);
or U6777 (N_6777,N_4126,N_5152);
nand U6778 (N_6778,N_5715,N_3954);
and U6779 (N_6779,N_5568,N_3385);
xnor U6780 (N_6780,N_5649,N_3252);
nor U6781 (N_6781,N_4988,N_4578);
xor U6782 (N_6782,N_5484,N_4879);
nor U6783 (N_6783,N_3557,N_5289);
nor U6784 (N_6784,N_3091,N_5685);
or U6785 (N_6785,N_5413,N_4719);
nand U6786 (N_6786,N_5489,N_4296);
nand U6787 (N_6787,N_4135,N_5236);
or U6788 (N_6788,N_5724,N_4113);
or U6789 (N_6789,N_4826,N_4472);
and U6790 (N_6790,N_4460,N_3518);
nand U6791 (N_6791,N_3119,N_3340);
or U6792 (N_6792,N_3752,N_3109);
and U6793 (N_6793,N_4221,N_5351);
nand U6794 (N_6794,N_4382,N_5748);
nand U6795 (N_6795,N_3019,N_4111);
nand U6796 (N_6796,N_4933,N_5431);
and U6797 (N_6797,N_5809,N_4091);
nand U6798 (N_6798,N_4801,N_4970);
nor U6799 (N_6799,N_5576,N_4169);
nand U6800 (N_6800,N_5069,N_5259);
nor U6801 (N_6801,N_3087,N_5455);
nor U6802 (N_6802,N_4055,N_4105);
xnor U6803 (N_6803,N_3201,N_5951);
nor U6804 (N_6804,N_4395,N_4641);
nand U6805 (N_6805,N_3695,N_3688);
or U6806 (N_6806,N_5371,N_4900);
and U6807 (N_6807,N_5836,N_3515);
nand U6808 (N_6808,N_4116,N_3739);
or U6809 (N_6809,N_5872,N_5388);
xor U6810 (N_6810,N_4053,N_4617);
and U6811 (N_6811,N_3690,N_4056);
or U6812 (N_6812,N_5577,N_4788);
nand U6813 (N_6813,N_3278,N_4337);
nor U6814 (N_6814,N_3839,N_3684);
or U6815 (N_6815,N_4972,N_5185);
or U6816 (N_6816,N_3342,N_4471);
or U6817 (N_6817,N_4920,N_5042);
nand U6818 (N_6818,N_3216,N_3297);
and U6819 (N_6819,N_4028,N_5784);
nor U6820 (N_6820,N_5312,N_3796);
and U6821 (N_6821,N_5048,N_5904);
nand U6822 (N_6822,N_3648,N_4642);
nand U6823 (N_6823,N_3224,N_5018);
or U6824 (N_6824,N_4366,N_3219);
nand U6825 (N_6825,N_3597,N_4167);
nand U6826 (N_6826,N_5811,N_4078);
nand U6827 (N_6827,N_3489,N_3266);
and U6828 (N_6828,N_3114,N_5347);
xnor U6829 (N_6829,N_3126,N_4264);
nor U6830 (N_6830,N_3736,N_5897);
nand U6831 (N_6831,N_3052,N_3765);
or U6832 (N_6832,N_3588,N_3977);
xor U6833 (N_6833,N_5453,N_5726);
nor U6834 (N_6834,N_5458,N_4996);
nor U6835 (N_6835,N_3326,N_4890);
nor U6836 (N_6836,N_5470,N_3408);
nand U6837 (N_6837,N_5304,N_3135);
nor U6838 (N_6838,N_4612,N_3585);
nand U6839 (N_6839,N_3917,N_3717);
or U6840 (N_6840,N_3323,N_5580);
nor U6841 (N_6841,N_4957,N_4623);
and U6842 (N_6842,N_5670,N_3371);
nand U6843 (N_6843,N_5262,N_3151);
nor U6844 (N_6844,N_5350,N_4872);
nand U6845 (N_6845,N_3834,N_4393);
nand U6846 (N_6846,N_4853,N_5404);
nand U6847 (N_6847,N_5460,N_5474);
nand U6848 (N_6848,N_5823,N_3415);
or U6849 (N_6849,N_5439,N_5129);
nor U6850 (N_6850,N_4025,N_3873);
and U6851 (N_6851,N_3000,N_3528);
nand U6852 (N_6852,N_5078,N_5648);
nor U6853 (N_6853,N_4705,N_4367);
or U6854 (N_6854,N_4484,N_5168);
nand U6855 (N_6855,N_4047,N_3919);
nor U6856 (N_6856,N_3092,N_3809);
and U6857 (N_6857,N_4898,N_5194);
nand U6858 (N_6858,N_4735,N_5159);
nor U6859 (N_6859,N_3107,N_4451);
xor U6860 (N_6860,N_3996,N_4839);
nor U6861 (N_6861,N_4333,N_4483);
or U6862 (N_6862,N_3777,N_4216);
or U6863 (N_6863,N_5898,N_4253);
nand U6864 (N_6864,N_5167,N_4874);
and U6865 (N_6865,N_3045,N_3104);
and U6866 (N_6866,N_5674,N_4504);
nand U6867 (N_6867,N_3222,N_5631);
nand U6868 (N_6868,N_3907,N_4597);
xnor U6869 (N_6869,N_4202,N_4240);
and U6870 (N_6870,N_4171,N_4506);
nand U6871 (N_6871,N_3067,N_5081);
or U6872 (N_6872,N_4669,N_5163);
nand U6873 (N_6873,N_3485,N_3564);
or U6874 (N_6874,N_4477,N_5282);
nor U6875 (N_6875,N_3283,N_3598);
or U6876 (N_6876,N_5072,N_4285);
nand U6877 (N_6877,N_3381,N_4489);
and U6878 (N_6878,N_3513,N_4402);
nand U6879 (N_6879,N_5948,N_3646);
nand U6880 (N_6880,N_4683,N_4549);
and U6881 (N_6881,N_3237,N_3011);
nor U6882 (N_6882,N_5495,N_3112);
nand U6883 (N_6883,N_4592,N_3445);
nand U6884 (N_6884,N_4227,N_4589);
and U6885 (N_6885,N_3286,N_4757);
or U6886 (N_6886,N_3263,N_4829);
nand U6887 (N_6887,N_3008,N_4424);
nor U6888 (N_6888,N_5099,N_4173);
nor U6889 (N_6889,N_3210,N_4936);
or U6890 (N_6890,N_3533,N_5089);
nand U6891 (N_6891,N_4744,N_5146);
and U6892 (N_6892,N_3421,N_5153);
nor U6893 (N_6893,N_4095,N_5061);
or U6894 (N_6894,N_4807,N_3563);
or U6895 (N_6895,N_3226,N_4600);
and U6896 (N_6896,N_4985,N_3268);
nor U6897 (N_6897,N_3638,N_3735);
and U6898 (N_6898,N_3434,N_4870);
or U6899 (N_6899,N_3433,N_3193);
nand U6900 (N_6900,N_4368,N_4225);
nor U6901 (N_6901,N_4144,N_5170);
nor U6902 (N_6902,N_5001,N_5071);
or U6903 (N_6903,N_3439,N_5532);
nor U6904 (N_6904,N_4238,N_4081);
and U6905 (N_6905,N_5247,N_3879);
or U6906 (N_6906,N_5524,N_3924);
and U6907 (N_6907,N_3177,N_4802);
or U6908 (N_6908,N_3446,N_5767);
or U6909 (N_6909,N_3535,N_4604);
nand U6910 (N_6910,N_3077,N_4770);
nor U6911 (N_6911,N_5832,N_5086);
and U6912 (N_6912,N_5429,N_3390);
nor U6913 (N_6913,N_5108,N_5184);
nor U6914 (N_6914,N_5336,N_4633);
or U6915 (N_6915,N_5126,N_3040);
nor U6916 (N_6916,N_3175,N_3499);
nor U6917 (N_6917,N_3354,N_5014);
and U6918 (N_6918,N_3413,N_4304);
nor U6919 (N_6919,N_5633,N_3964);
nor U6920 (N_6920,N_5618,N_4467);
and U6921 (N_6921,N_3553,N_4598);
nand U6922 (N_6922,N_3663,N_3072);
and U6923 (N_6923,N_5827,N_4812);
nand U6924 (N_6924,N_5481,N_5829);
or U6925 (N_6925,N_5358,N_3831);
nor U6926 (N_6926,N_4570,N_3801);
nor U6927 (N_6927,N_3383,N_3878);
or U6928 (N_6928,N_5777,N_4345);
and U6929 (N_6929,N_3676,N_3810);
and U6930 (N_6930,N_3904,N_3963);
and U6931 (N_6931,N_5433,N_4661);
nor U6932 (N_6932,N_5665,N_5862);
nor U6933 (N_6933,N_4937,N_3493);
or U6934 (N_6934,N_3377,N_5550);
or U6935 (N_6935,N_5655,N_4941);
nand U6936 (N_6936,N_3855,N_4902);
nor U6937 (N_6937,N_3213,N_5047);
or U6938 (N_6938,N_5985,N_3994);
nor U6939 (N_6939,N_3868,N_4261);
and U6940 (N_6940,N_4242,N_4259);
xor U6941 (N_6941,N_3337,N_3665);
or U6942 (N_6942,N_5621,N_5514);
nand U6943 (N_6943,N_5608,N_5472);
xor U6944 (N_6944,N_3558,N_5448);
nor U6945 (N_6945,N_4541,N_3249);
nor U6946 (N_6946,N_4377,N_3356);
nor U6947 (N_6947,N_3452,N_4626);
and U6948 (N_6948,N_5567,N_3578);
nand U6949 (N_6949,N_5302,N_5360);
or U6950 (N_6950,N_4212,N_3877);
nor U6951 (N_6951,N_3048,N_3118);
nor U6952 (N_6952,N_4124,N_3304);
nor U6953 (N_6953,N_5499,N_3857);
or U6954 (N_6954,N_4319,N_3623);
nand U6955 (N_6955,N_3227,N_4778);
or U6956 (N_6956,N_4776,N_5684);
and U6957 (N_6957,N_3444,N_5258);
or U6958 (N_6958,N_3301,N_3824);
and U6959 (N_6959,N_5320,N_3643);
and U6960 (N_6960,N_5693,N_3902);
and U6961 (N_6961,N_3414,N_4500);
nor U6962 (N_6962,N_4564,N_4946);
or U6963 (N_6963,N_5468,N_4070);
nor U6964 (N_6964,N_3284,N_5396);
xor U6965 (N_6965,N_3246,N_4916);
nor U6966 (N_6966,N_3296,N_4404);
and U6967 (N_6967,N_5257,N_5605);
or U6968 (N_6968,N_4234,N_3522);
or U6969 (N_6969,N_4708,N_3144);
nor U6970 (N_6970,N_5309,N_3790);
nor U6971 (N_6971,N_3432,N_4406);
or U6972 (N_6972,N_4635,N_3693);
nand U6973 (N_6973,N_3921,N_3478);
nand U6974 (N_6974,N_3745,N_3007);
nand U6975 (N_6975,N_3683,N_4076);
and U6976 (N_6976,N_5906,N_4186);
nor U6977 (N_6977,N_4275,N_4713);
nand U6978 (N_6978,N_3384,N_5074);
or U6979 (N_6979,N_3605,N_3616);
or U6980 (N_6980,N_5955,N_4448);
and U6981 (N_6981,N_5483,N_3703);
and U6982 (N_6982,N_4583,N_5600);
nor U6983 (N_6983,N_5707,N_3905);
nor U6984 (N_6984,N_4231,N_4270);
or U6985 (N_6985,N_3516,N_4307);
or U6986 (N_6986,N_3723,N_5379);
or U6987 (N_6987,N_3078,N_3199);
xnor U6988 (N_6988,N_3348,N_5669);
nand U6989 (N_6989,N_5879,N_5691);
nand U6990 (N_6990,N_5916,N_5566);
xnor U6991 (N_6991,N_3392,N_3799);
or U6992 (N_6992,N_3547,N_5557);
or U6993 (N_6993,N_5912,N_3269);
and U6994 (N_6994,N_3136,N_3767);
and U6995 (N_6995,N_4751,N_4233);
nand U6996 (N_6996,N_3984,N_3674);
nor U6997 (N_6997,N_5342,N_4235);
nor U6998 (N_6998,N_3895,N_3660);
nor U6999 (N_6999,N_5846,N_3025);
and U7000 (N_7000,N_4031,N_3872);
or U7001 (N_7001,N_3005,N_4112);
and U7002 (N_7002,N_5426,N_5380);
or U7003 (N_7003,N_4288,N_4084);
nor U7004 (N_7004,N_3524,N_4455);
nor U7005 (N_7005,N_4277,N_4391);
nand U7006 (N_7006,N_3295,N_4869);
nand U7007 (N_7007,N_4825,N_4355);
and U7008 (N_7008,N_4362,N_4158);
or U7009 (N_7009,N_4045,N_5698);
or U7010 (N_7010,N_5517,N_5870);
nor U7011 (N_7011,N_4164,N_4062);
and U7012 (N_7012,N_3504,N_3755);
or U7013 (N_7013,N_3658,N_5500);
and U7014 (N_7014,N_3037,N_4463);
nor U7015 (N_7015,N_4281,N_5406);
and U7016 (N_7016,N_3013,N_4004);
or U7017 (N_7017,N_4591,N_3666);
nand U7018 (N_7018,N_4273,N_3028);
nand U7019 (N_7019,N_3429,N_5511);
nor U7020 (N_7020,N_5759,N_3566);
or U7021 (N_7021,N_5667,N_3036);
and U7022 (N_7022,N_3732,N_5694);
or U7023 (N_7023,N_4032,N_4695);
nor U7024 (N_7024,N_4939,N_3260);
nand U7025 (N_7025,N_5223,N_4454);
or U7026 (N_7026,N_4320,N_3234);
nand U7027 (N_7027,N_5242,N_3718);
and U7028 (N_7028,N_5154,N_4836);
or U7029 (N_7029,N_5962,N_4322);
and U7030 (N_7030,N_5997,N_3630);
nor U7031 (N_7031,N_4796,N_3481);
or U7032 (N_7032,N_5134,N_3474);
nor U7033 (N_7033,N_5852,N_4429);
nor U7034 (N_7034,N_3552,N_5664);
or U7035 (N_7035,N_5007,N_5162);
xor U7036 (N_7036,N_5299,N_5604);
nor U7037 (N_7037,N_5722,N_3289);
nand U7038 (N_7038,N_5746,N_4848);
nand U7039 (N_7039,N_5574,N_3070);
and U7040 (N_7040,N_4717,N_3841);
nor U7041 (N_7041,N_4620,N_5005);
or U7042 (N_7042,N_4850,N_4794);
and U7043 (N_7043,N_4982,N_3759);
nand U7044 (N_7044,N_3673,N_4444);
nand U7045 (N_7045,N_5990,N_5656);
or U7046 (N_7046,N_5756,N_3034);
or U7047 (N_7047,N_4419,N_5418);
or U7048 (N_7048,N_5210,N_3751);
nor U7049 (N_7049,N_3093,N_3430);
or U7050 (N_7050,N_3675,N_3014);
and U7051 (N_7051,N_5553,N_3403);
nand U7052 (N_7052,N_3270,N_5492);
nand U7053 (N_7053,N_4888,N_5092);
nor U7054 (N_7054,N_3479,N_4772);
and U7055 (N_7055,N_4466,N_4774);
and U7056 (N_7056,N_4797,N_3657);
nor U7057 (N_7057,N_5311,N_5106);
or U7058 (N_7058,N_4659,N_4983);
xnor U7059 (N_7059,N_4248,N_4228);
and U7060 (N_7060,N_3115,N_5597);
or U7061 (N_7061,N_4553,N_3076);
or U7062 (N_7062,N_5952,N_4119);
nand U7063 (N_7063,N_4980,N_4476);
or U7064 (N_7064,N_4795,N_3103);
nand U7065 (N_7065,N_4263,N_5179);
xor U7066 (N_7066,N_4857,N_5749);
and U7067 (N_7067,N_5234,N_3164);
nand U7068 (N_7068,N_5467,N_4197);
and U7069 (N_7069,N_3035,N_4934);
and U7070 (N_7070,N_3195,N_4532);
nand U7071 (N_7071,N_3194,N_4066);
nor U7072 (N_7072,N_5793,N_3883);
nor U7073 (N_7073,N_5006,N_3544);
nand U7074 (N_7074,N_3245,N_4324);
nand U7075 (N_7075,N_4793,N_3307);
nand U7076 (N_7076,N_3619,N_4494);
and U7077 (N_7077,N_5314,N_5982);
nand U7078 (N_7078,N_3123,N_5409);
or U7079 (N_7079,N_5781,N_3370);
xnor U7080 (N_7080,N_5980,N_5525);
xnor U7081 (N_7081,N_4474,N_3397);
nor U7082 (N_7082,N_5541,N_4042);
or U7083 (N_7083,N_4574,N_4992);
or U7084 (N_7084,N_4033,N_4686);
nand U7085 (N_7085,N_3587,N_3724);
and U7086 (N_7086,N_3862,N_5369);
and U7087 (N_7087,N_5794,N_3746);
and U7088 (N_7088,N_4329,N_5207);
nor U7089 (N_7089,N_4295,N_3985);
nor U7090 (N_7090,N_4308,N_3669);
and U7091 (N_7091,N_3898,N_3864);
and U7092 (N_7092,N_5337,N_3259);
or U7093 (N_7093,N_3492,N_3953);
nand U7094 (N_7094,N_5117,N_4256);
nand U7095 (N_7095,N_4306,N_5779);
nor U7096 (N_7096,N_5050,N_3510);
nor U7097 (N_7097,N_4820,N_5288);
nand U7098 (N_7098,N_4990,N_3699);
xnor U7099 (N_7099,N_4720,N_5923);
and U7100 (N_7100,N_4580,N_4087);
or U7101 (N_7101,N_4865,N_4656);
nor U7102 (N_7102,N_3345,N_4928);
nand U7103 (N_7103,N_3753,N_5805);
and U7104 (N_7104,N_3376,N_5232);
and U7105 (N_7105,N_3238,N_5297);
and U7106 (N_7106,N_5070,N_5596);
nor U7107 (N_7107,N_5630,N_3545);
or U7108 (N_7108,N_5097,N_3394);
xnor U7109 (N_7109,N_3097,N_5356);
nand U7110 (N_7110,N_4873,N_4165);
and U7111 (N_7111,N_4875,N_4977);
nor U7112 (N_7112,N_3314,N_5209);
and U7113 (N_7113,N_3242,N_3687);
or U7114 (N_7114,N_5139,N_4814);
and U7115 (N_7115,N_4088,N_3710);
xor U7116 (N_7116,N_4557,N_3363);
and U7117 (N_7117,N_4967,N_5610);
and U7118 (N_7118,N_5841,N_4852);
and U7119 (N_7119,N_5115,N_3789);
or U7120 (N_7120,N_4153,N_4538);
or U7121 (N_7121,N_5818,N_5753);
nand U7122 (N_7122,N_5272,N_3962);
and U7123 (N_7123,N_4334,N_4099);
nor U7124 (N_7124,N_4211,N_4485);
or U7125 (N_7125,N_3458,N_3054);
nand U7126 (N_7126,N_4729,N_3006);
or U7127 (N_7127,N_3837,N_4229);
nand U7128 (N_7128,N_4819,N_3257);
or U7129 (N_7129,N_5131,N_5571);
or U7130 (N_7130,N_5093,N_5465);
nand U7131 (N_7131,N_4436,N_5385);
and U7132 (N_7132,N_4254,N_4769);
and U7133 (N_7133,N_3184,N_5450);
xor U7134 (N_7134,N_4191,N_3708);
nand U7135 (N_7135,N_4614,N_5263);
nor U7136 (N_7136,N_4220,N_3161);
nor U7137 (N_7137,N_5814,N_4301);
and U7138 (N_7138,N_3085,N_4060);
nor U7139 (N_7139,N_5349,N_4856);
nand U7140 (N_7140,N_5619,N_5922);
or U7141 (N_7141,N_3678,N_5972);
nand U7142 (N_7142,N_5677,N_4844);
and U7143 (N_7143,N_5387,N_4565);
nand U7144 (N_7144,N_3702,N_5090);
or U7145 (N_7145,N_4764,N_3300);
or U7146 (N_7146,N_5260,N_5088);
nand U7147 (N_7147,N_5799,N_5354);
and U7148 (N_7148,N_4618,N_5929);
and U7149 (N_7149,N_3121,N_3101);
and U7150 (N_7150,N_5765,N_3946);
or U7151 (N_7151,N_4575,N_3861);
or U7152 (N_7152,N_4346,N_3541);
nand U7153 (N_7153,N_4632,N_5140);
or U7154 (N_7154,N_3389,N_5250);
nor U7155 (N_7155,N_4816,N_5855);
nor U7156 (N_7156,N_4251,N_4692);
nand U7157 (N_7157,N_5762,N_5966);
nand U7158 (N_7158,N_3150,N_3418);
nor U7159 (N_7159,N_3347,N_5326);
and U7160 (N_7160,N_3770,N_3992);
nor U7161 (N_7161,N_3612,N_5683);
nand U7162 (N_7162,N_5909,N_5323);
or U7163 (N_7163,N_3891,N_5622);
nor U7164 (N_7164,N_5536,N_5025);
nor U7165 (N_7165,N_3145,N_5563);
nor U7166 (N_7166,N_4615,N_5416);
nand U7167 (N_7167,N_5285,N_4210);
nand U7168 (N_7168,N_3574,N_5105);
and U7169 (N_7169,N_4616,N_3443);
or U7170 (N_7170,N_5228,N_5999);
nand U7171 (N_7171,N_5255,N_4923);
nor U7172 (N_7172,N_4501,N_4376);
xor U7173 (N_7173,N_3849,N_3580);
nor U7174 (N_7174,N_4943,N_4120);
or U7175 (N_7175,N_5203,N_4822);
or U7176 (N_7176,N_3711,N_3243);
nor U7177 (N_7177,N_5156,N_4162);
and U7178 (N_7178,N_3532,N_4097);
nand U7179 (N_7179,N_5750,N_4464);
and U7180 (N_7180,N_3974,N_3804);
or U7181 (N_7181,N_5004,N_5918);
or U7182 (N_7182,N_5246,N_3881);
xor U7183 (N_7183,N_3338,N_5518);
nand U7184 (N_7184,N_4457,N_5936);
nand U7185 (N_7185,N_5925,N_5643);
or U7186 (N_7186,N_5908,N_3781);
nor U7187 (N_7187,N_5976,N_3694);
and U7188 (N_7188,N_4141,N_5945);
nand U7189 (N_7189,N_4950,N_3229);
nor U7190 (N_7190,N_5731,N_3949);
or U7191 (N_7191,N_4199,N_3590);
nor U7192 (N_7192,N_5485,N_3064);
nor U7193 (N_7193,N_4303,N_4805);
or U7194 (N_7194,N_5815,N_5398);
nor U7195 (N_7195,N_4595,N_3050);
or U7196 (N_7196,N_3555,N_5332);
nor U7197 (N_7197,N_4353,N_5699);
nor U7198 (N_7198,N_4854,N_4726);
nand U7199 (N_7199,N_5864,N_3473);
nor U7200 (N_7200,N_3420,N_4000);
nand U7201 (N_7201,N_5290,N_4786);
and U7202 (N_7202,N_5034,N_3922);
or U7203 (N_7203,N_5776,N_5578);
or U7204 (N_7204,N_4311,N_3670);
nand U7205 (N_7205,N_3859,N_4657);
nor U7206 (N_7206,N_3749,N_3947);
nand U7207 (N_7207,N_4152,N_3254);
nand U7208 (N_7208,N_5882,N_3176);
nand U7209 (N_7209,N_3375,N_3940);
or U7210 (N_7210,N_3113,N_5752);
xor U7211 (N_7211,N_5687,N_4573);
nor U7212 (N_7212,N_4409,N_4168);
nor U7213 (N_7213,N_3507,N_4643);
nor U7214 (N_7214,N_3888,N_5235);
or U7215 (N_7215,N_3901,N_4286);
or U7216 (N_7216,N_5410,N_3852);
nor U7217 (N_7217,N_5785,N_3938);
and U7218 (N_7218,N_5218,N_3364);
nand U7219 (N_7219,N_3838,N_3327);
nand U7220 (N_7220,N_3168,N_3560);
nor U7221 (N_7221,N_3584,N_3057);
or U7222 (N_7222,N_4040,N_3995);
or U7223 (N_7223,N_4428,N_5732);
nor U7224 (N_7224,N_3778,N_4226);
and U7225 (N_7225,N_3689,N_3576);
nand U7226 (N_7226,N_4582,N_4671);
and U7227 (N_7227,N_3798,N_3221);
nor U7228 (N_7228,N_5330,N_4461);
nor U7229 (N_7229,N_5523,N_4508);
nand U7230 (N_7230,N_3191,N_3722);
nand U7231 (N_7231,N_5657,N_3599);
and U7232 (N_7232,N_3783,N_4511);
and U7233 (N_7233,N_5346,N_3763);
nor U7234 (N_7234,N_3697,N_5927);
or U7235 (N_7235,N_5361,N_3134);
nor U7236 (N_7236,N_3826,N_4019);
or U7237 (N_7237,N_5965,N_3896);
nor U7238 (N_7238,N_4897,N_5305);
nor U7239 (N_7239,N_3277,N_4768);
nor U7240 (N_7240,N_3639,N_5447);
and U7241 (N_7241,N_5464,N_3409);
nand U7242 (N_7242,N_5661,N_4143);
nand U7243 (N_7243,N_4732,N_3502);
and U7244 (N_7244,N_5617,N_4104);
and U7245 (N_7245,N_4640,N_3976);
nand U7246 (N_7246,N_4662,N_5522);
and U7247 (N_7247,N_3512,N_3165);
and U7248 (N_7248,N_5190,N_3181);
or U7249 (N_7249,N_5196,N_4192);
or U7250 (N_7250,N_4860,N_3100);
nand U7251 (N_7251,N_4981,N_5920);
nor U7252 (N_7252,N_4224,N_5032);
nor U7253 (N_7253,N_5853,N_3527);
nand U7254 (N_7254,N_3725,N_5690);
or U7255 (N_7255,N_3153,N_5390);
nor U7256 (N_7256,N_4267,N_3339);
or U7257 (N_7257,N_3618,N_4154);
nor U7258 (N_7258,N_4777,N_3021);
and U7259 (N_7259,N_5883,N_5402);
nand U7260 (N_7260,N_4756,N_5469);
nor U7261 (N_7261,N_3914,N_3477);
nor U7262 (N_7262,N_3068,N_3656);
and U7263 (N_7263,N_5902,N_5708);
nand U7264 (N_7264,N_3936,N_4358);
nand U7265 (N_7265,N_5696,N_5204);
and U7266 (N_7266,N_4734,N_5038);
or U7267 (N_7267,N_5740,N_5123);
or U7268 (N_7268,N_4545,N_5341);
and U7269 (N_7269,N_5559,N_5516);
nor U7270 (N_7270,N_4602,N_4063);
or U7271 (N_7271,N_3664,N_3570);
and U7272 (N_7272,N_4102,N_5856);
nor U7273 (N_7273,N_5030,N_4910);
or U7274 (N_7274,N_5692,N_5720);
or U7275 (N_7275,N_5444,N_3281);
and U7276 (N_7276,N_5116,N_4523);
nor U7277 (N_7277,N_3333,N_5240);
or U7278 (N_7278,N_4039,N_3945);
or U7279 (N_7279,N_3062,N_5653);
or U7280 (N_7280,N_4789,N_5995);
nor U7281 (N_7281,N_5526,N_3451);
nor U7282 (N_7282,N_3651,N_3362);
nand U7283 (N_7283,N_3335,N_3197);
or U7284 (N_7284,N_5158,N_3386);
nand U7285 (N_7285,N_5477,N_5454);
and U7286 (N_7286,N_5808,N_4160);
nor U7287 (N_7287,N_5595,N_4510);
and U7288 (N_7288,N_5381,N_5802);
nand U7289 (N_7289,N_3983,N_5165);
nand U7290 (N_7290,N_3705,N_5958);
nand U7291 (N_7291,N_4035,N_5459);
or U7292 (N_7292,N_3428,N_4188);
nor U7293 (N_7293,N_5102,N_3644);
nor U7294 (N_7294,N_5711,N_3074);
nand U7295 (N_7295,N_5689,N_3517);
nor U7296 (N_7296,N_3915,N_4312);
or U7297 (N_7297,N_3713,N_4989);
and U7298 (N_7298,N_5414,N_3827);
and U7299 (N_7299,N_4332,N_5635);
nor U7300 (N_7300,N_5991,N_4515);
nand U7301 (N_7301,N_5840,N_4387);
nor U7302 (N_7302,N_3017,N_4624);
nand U7303 (N_7303,N_3349,N_5796);
nor U7304 (N_7304,N_3805,N_3090);
nor U7305 (N_7305,N_5463,N_3506);
or U7306 (N_7306,N_4305,N_3602);
xor U7307 (N_7307,N_3795,N_5729);
or U7308 (N_7308,N_4005,N_3525);
nor U7309 (N_7309,N_4687,N_5372);
nor U7310 (N_7310,N_3470,N_3464);
nand U7311 (N_7311,N_4818,N_3776);
and U7312 (N_7312,N_3125,N_3727);
nand U7313 (N_7313,N_5208,N_4847);
nor U7314 (N_7314,N_4356,N_3772);
nor U7315 (N_7315,N_3298,N_5778);
nor U7316 (N_7316,N_5587,N_4673);
or U7317 (N_7317,N_3240,N_5804);
nand U7318 (N_7318,N_3166,N_3212);
nor U7319 (N_7319,N_5094,N_3993);
or U7320 (N_7320,N_5279,N_5191);
or U7321 (N_7321,N_4743,N_5334);
or U7322 (N_7322,N_5924,N_3997);
nor U7323 (N_7323,N_3053,N_4716);
or U7324 (N_7324,N_3579,N_5974);
and U7325 (N_7325,N_4895,N_5801);
and U7326 (N_7326,N_3679,N_3448);
nand U7327 (N_7327,N_3747,N_3436);
or U7328 (N_7328,N_5847,N_4246);
nand U7329 (N_7329,N_3894,N_3496);
or U7330 (N_7330,N_5120,N_5530);
and U7331 (N_7331,N_5128,N_5950);
nand U7332 (N_7332,N_4134,N_4773);
nor U7333 (N_7333,N_4058,N_3771);
and U7334 (N_7334,N_3422,N_4475);
nand U7335 (N_7335,N_5331,N_4606);
and U7336 (N_7336,N_3425,N_3908);
nand U7337 (N_7337,N_4681,N_4507);
nor U7338 (N_7338,N_3892,N_4792);
nand U7339 (N_7339,N_5419,N_4094);
nor U7340 (N_7340,N_4755,N_4001);
or U7341 (N_7341,N_3442,N_3170);
nor U7342 (N_7342,N_3098,N_4207);
nand U7343 (N_7343,N_3148,N_4003);
nor U7344 (N_7344,N_5682,N_3282);
or U7345 (N_7345,N_5079,N_5253);
or U7346 (N_7346,N_3626,N_4513);
and U7347 (N_7347,N_4222,N_3069);
nand U7348 (N_7348,N_5338,N_4730);
or U7349 (N_7349,N_3265,N_3271);
or U7350 (N_7350,N_4694,N_5782);
nand U7351 (N_7351,N_5248,N_4862);
nor U7352 (N_7352,N_4465,N_5967);
or U7353 (N_7353,N_4978,N_4925);
and U7354 (N_7354,N_4369,N_3685);
and U7355 (N_7355,N_4189,N_3071);
or U7356 (N_7356,N_4100,N_4127);
and U7357 (N_7357,N_3288,N_4422);
nor U7358 (N_7358,N_3712,N_4993);
and U7359 (N_7359,N_4114,N_3412);
nor U7360 (N_7360,N_4128,N_3401);
or U7361 (N_7361,N_4262,N_4843);
nor U7362 (N_7362,N_4316,N_4607);
nor U7363 (N_7363,N_5569,N_3766);
nand U7364 (N_7364,N_5977,N_4044);
xor U7365 (N_7365,N_4479,N_5503);
or U7366 (N_7366,N_4884,N_3056);
and U7367 (N_7367,N_3159,N_5984);
nand U7368 (N_7368,N_3632,N_3932);
and U7369 (N_7369,N_4020,N_3787);
or U7370 (N_7370,N_3230,N_3860);
xor U7371 (N_7371,N_5881,N_4196);
or U7372 (N_7372,N_5421,N_4416);
or U7373 (N_7373,N_3817,N_5941);
nor U7374 (N_7374,N_5723,N_4759);
or U7375 (N_7375,N_4131,N_4975);
nor U7376 (N_7376,N_5243,N_4438);
or U7377 (N_7377,N_4904,N_3202);
or U7378 (N_7378,N_5487,N_3958);
nor U7379 (N_7379,N_5225,N_4187);
nor U7380 (N_7380,N_3833,N_3018);
nor U7381 (N_7381,N_4036,N_3939);
or U7382 (N_7382,N_5220,N_4885);
and U7383 (N_7383,N_5903,N_5497);
and U7384 (N_7384,N_5174,N_3737);
nor U7385 (N_7385,N_5506,N_5286);
nor U7386 (N_7386,N_5340,N_3721);
nor U7387 (N_7387,N_5865,N_3965);
nor U7388 (N_7388,N_4917,N_4341);
and U7389 (N_7389,N_4082,N_3508);
nand U7390 (N_7390,N_3923,N_4667);
and U7391 (N_7391,N_5705,N_3955);
nand U7392 (N_7392,N_5049,N_3728);
nor U7393 (N_7393,N_4057,N_5052);
nand U7394 (N_7394,N_5886,N_4397);
nand U7395 (N_7395,N_5298,N_5921);
nand U7396 (N_7396,N_4760,N_5029);
or U7397 (N_7397,N_4118,N_3490);
nand U7398 (N_7398,N_4190,N_5539);
or U7399 (N_7399,N_3031,N_3575);
or U7400 (N_7400,N_4182,N_5926);
and U7401 (N_7401,N_5519,N_4645);
nor U7402 (N_7402,N_4762,N_4752);
or U7403 (N_7403,N_5310,N_3754);
and U7404 (N_7404,N_4166,N_5407);
nand U7405 (N_7405,N_4110,N_3812);
and U7406 (N_7406,N_5101,N_5241);
nand U7407 (N_7407,N_5176,N_4250);
nor U7408 (N_7408,N_4435,N_3726);
and U7409 (N_7409,N_3004,N_3850);
or U7410 (N_7410,N_3750,N_5221);
nand U7411 (N_7411,N_5425,N_5772);
or U7412 (N_7412,N_3645,N_3127);
nor U7413 (N_7413,N_4051,N_4374);
nand U7414 (N_7414,N_4499,N_4432);
or U7415 (N_7415,N_3606,N_5457);
nand U7416 (N_7416,N_3358,N_3784);
or U7417 (N_7417,N_3536,N_5542);
or U7418 (N_7418,N_5612,N_5831);
nand U7419 (N_7419,N_5646,N_4605);
nand U7420 (N_7420,N_5593,N_5616);
and U7421 (N_7421,N_5531,N_3594);
nand U7422 (N_7422,N_4482,N_5056);
nor U7423 (N_7423,N_5520,N_5144);
nand U7424 (N_7424,N_5876,N_4061);
nand U7425 (N_7425,N_4148,N_4630);
nand U7426 (N_7426,N_3828,N_5059);
or U7427 (N_7427,N_3322,N_3572);
or U7428 (N_7428,N_5817,N_5813);
and U7429 (N_7429,N_4994,N_3130);
nor U7430 (N_7430,N_3173,N_5411);
and U7431 (N_7431,N_4784,N_5009);
or U7432 (N_7432,N_4568,N_5803);
and U7433 (N_7433,N_3065,N_5651);
nor U7434 (N_7434,N_5546,N_4115);
nand U7435 (N_7435,N_3030,N_4750);
and U7436 (N_7436,N_3956,N_5100);
and U7437 (N_7437,N_4746,N_5735);
or U7438 (N_7438,N_5133,N_5943);
nand U7439 (N_7439,N_3016,N_4373);
or U7440 (N_7440,N_3179,N_5486);
nand U7441 (N_7441,N_5287,N_3343);
or U7442 (N_7442,N_3840,N_4133);
nor U7443 (N_7443,N_5712,N_3059);
and U7444 (N_7444,N_4074,N_3373);
or U7445 (N_7445,N_3486,N_4926);
nand U7446 (N_7446,N_5743,N_4008);
nor U7447 (N_7447,N_5558,N_5274);
nor U7448 (N_7448,N_3534,N_5127);
nand U7449 (N_7449,N_5515,N_3465);
or U7450 (N_7450,N_3461,N_4372);
nor U7451 (N_7451,N_3836,N_3081);
and U7452 (N_7452,N_5527,N_3568);
and U7453 (N_7453,N_5181,N_5529);
nor U7454 (N_7454,N_4335,N_4837);
or U7455 (N_7455,N_4887,N_3262);
or U7456 (N_7456,N_5626,N_5806);
nand U7457 (N_7457,N_4026,N_3526);
or U7458 (N_7458,N_4054,N_3488);
or U7459 (N_7459,N_3634,N_3621);
or U7460 (N_7460,N_5020,N_4831);
and U7461 (N_7461,N_3235,N_5989);
or U7462 (N_7462,N_3157,N_5602);
nand U7463 (N_7463,N_3935,N_5930);
nor U7464 (N_7464,N_3352,N_3189);
and U7465 (N_7465,N_3821,N_4555);
or U7466 (N_7466,N_5844,N_3633);
nor U7467 (N_7467,N_3986,N_5706);
and U7468 (N_7468,N_4551,N_5751);
xor U7469 (N_7469,N_3671,N_3586);
and U7470 (N_7470,N_4558,N_3786);
or U7471 (N_7471,N_3320,N_4634);
nand U7472 (N_7472,N_3886,N_4593);
or U7473 (N_7473,N_3012,N_5028);
nor U7474 (N_7474,N_4963,N_5716);
nor U7475 (N_7475,N_3038,N_5308);
or U7476 (N_7476,N_3698,N_3198);
nor U7477 (N_7477,N_5212,N_5064);
and U7478 (N_7478,N_4942,N_5598);
nor U7479 (N_7479,N_5642,N_5244);
or U7480 (N_7480,N_3416,N_5098);
or U7481 (N_7481,N_5400,N_5545);
and U7482 (N_7482,N_4715,N_4007);
nand U7483 (N_7483,N_5961,N_5549);
nand U7484 (N_7484,N_3942,N_5614);
nand U7485 (N_7485,N_5636,N_5177);
and U7486 (N_7486,N_5896,N_4401);
nand U7487 (N_7487,N_4347,N_4151);
nor U7488 (N_7488,N_4986,N_3391);
nor U7489 (N_7489,N_3627,N_4426);
nor U7490 (N_7490,N_3033,N_5968);
nor U7491 (N_7491,N_4200,N_3652);
and U7492 (N_7492,N_3395,N_3475);
or U7493 (N_7493,N_5412,N_4271);
nor U7494 (N_7494,N_4230,N_4876);
and U7495 (N_7495,N_3972,N_3764);
and U7496 (N_7496,N_4452,N_5044);
or U7497 (N_7497,N_4979,N_5505);
nor U7498 (N_7498,N_4956,N_4065);
nor U7499 (N_7499,N_5437,N_3061);
xnor U7500 (N_7500,N_5766,N_4707);
nand U7501 (N_7501,N_5037,N_4503);
and U7502 (N_7502,N_3344,N_4562);
nor U7503 (N_7503,N_3560,N_4652);
nor U7504 (N_7504,N_3647,N_3234);
and U7505 (N_7505,N_4146,N_3012);
and U7506 (N_7506,N_4484,N_4113);
or U7507 (N_7507,N_4102,N_4441);
and U7508 (N_7508,N_3461,N_5617);
or U7509 (N_7509,N_5529,N_4242);
nand U7510 (N_7510,N_4515,N_4413);
nand U7511 (N_7511,N_5861,N_5151);
nor U7512 (N_7512,N_3805,N_3018);
nand U7513 (N_7513,N_4378,N_5509);
or U7514 (N_7514,N_3339,N_4494);
nand U7515 (N_7515,N_4478,N_4262);
nand U7516 (N_7516,N_3756,N_4481);
nor U7517 (N_7517,N_4386,N_3398);
nor U7518 (N_7518,N_4683,N_4684);
nor U7519 (N_7519,N_5575,N_4395);
nor U7520 (N_7520,N_3148,N_5124);
or U7521 (N_7521,N_3127,N_4715);
nand U7522 (N_7522,N_4098,N_5177);
nand U7523 (N_7523,N_4818,N_4844);
nand U7524 (N_7524,N_4878,N_4747);
nand U7525 (N_7525,N_4974,N_4032);
xnor U7526 (N_7526,N_5685,N_5160);
and U7527 (N_7527,N_3193,N_3344);
nor U7528 (N_7528,N_3094,N_4496);
xor U7529 (N_7529,N_4533,N_5160);
or U7530 (N_7530,N_3854,N_5626);
nand U7531 (N_7531,N_3857,N_5997);
nand U7532 (N_7532,N_3636,N_5528);
nor U7533 (N_7533,N_4967,N_4706);
xor U7534 (N_7534,N_3498,N_4351);
nand U7535 (N_7535,N_4317,N_5292);
xor U7536 (N_7536,N_5813,N_5361);
and U7537 (N_7537,N_5356,N_5307);
nor U7538 (N_7538,N_3099,N_5222);
nand U7539 (N_7539,N_5448,N_4448);
and U7540 (N_7540,N_4389,N_3588);
nand U7541 (N_7541,N_3746,N_5338);
nor U7542 (N_7542,N_4331,N_5069);
nand U7543 (N_7543,N_5819,N_5090);
or U7544 (N_7544,N_5597,N_5537);
nand U7545 (N_7545,N_3137,N_3551);
or U7546 (N_7546,N_5009,N_4576);
nand U7547 (N_7547,N_3024,N_4383);
or U7548 (N_7548,N_3716,N_5049);
nor U7549 (N_7549,N_3606,N_3043);
nor U7550 (N_7550,N_5166,N_4633);
or U7551 (N_7551,N_5243,N_5292);
nor U7552 (N_7552,N_4157,N_5501);
nand U7553 (N_7553,N_4511,N_3084);
and U7554 (N_7554,N_4966,N_5019);
nand U7555 (N_7555,N_5233,N_3528);
nor U7556 (N_7556,N_3059,N_4445);
nor U7557 (N_7557,N_4975,N_3437);
and U7558 (N_7558,N_4927,N_5329);
and U7559 (N_7559,N_5939,N_5281);
and U7560 (N_7560,N_5672,N_4301);
xnor U7561 (N_7561,N_5420,N_4178);
nand U7562 (N_7562,N_4291,N_5889);
or U7563 (N_7563,N_3683,N_5388);
nor U7564 (N_7564,N_3765,N_4313);
xnor U7565 (N_7565,N_4138,N_5027);
nand U7566 (N_7566,N_4381,N_5453);
and U7567 (N_7567,N_3548,N_3496);
and U7568 (N_7568,N_3154,N_4384);
nor U7569 (N_7569,N_5066,N_5926);
nor U7570 (N_7570,N_3364,N_4225);
nor U7571 (N_7571,N_3184,N_4097);
or U7572 (N_7572,N_4400,N_3528);
nand U7573 (N_7573,N_5027,N_3470);
or U7574 (N_7574,N_3807,N_5742);
nor U7575 (N_7575,N_3423,N_4928);
xnor U7576 (N_7576,N_5037,N_5541);
xor U7577 (N_7577,N_3583,N_3958);
and U7578 (N_7578,N_3518,N_3763);
nor U7579 (N_7579,N_3660,N_4665);
nor U7580 (N_7580,N_5877,N_5415);
nand U7581 (N_7581,N_4516,N_5775);
or U7582 (N_7582,N_4567,N_4222);
nand U7583 (N_7583,N_5226,N_5653);
and U7584 (N_7584,N_4238,N_3064);
and U7585 (N_7585,N_5200,N_4272);
xnor U7586 (N_7586,N_4532,N_5295);
nand U7587 (N_7587,N_5214,N_4026);
nand U7588 (N_7588,N_5833,N_5473);
nand U7589 (N_7589,N_4643,N_4358);
nand U7590 (N_7590,N_5696,N_3314);
and U7591 (N_7591,N_3290,N_4465);
nor U7592 (N_7592,N_5609,N_3568);
nand U7593 (N_7593,N_3193,N_3435);
nor U7594 (N_7594,N_5871,N_5200);
nand U7595 (N_7595,N_3938,N_3753);
nand U7596 (N_7596,N_5878,N_5081);
nor U7597 (N_7597,N_5760,N_5513);
or U7598 (N_7598,N_5280,N_4744);
nor U7599 (N_7599,N_4743,N_3748);
or U7600 (N_7600,N_4108,N_3941);
nor U7601 (N_7601,N_5739,N_5496);
nand U7602 (N_7602,N_3040,N_3016);
nor U7603 (N_7603,N_4558,N_3943);
nand U7604 (N_7604,N_3616,N_5119);
and U7605 (N_7605,N_5807,N_5065);
or U7606 (N_7606,N_4299,N_5837);
nand U7607 (N_7607,N_3171,N_4260);
nand U7608 (N_7608,N_3282,N_3949);
or U7609 (N_7609,N_3010,N_3849);
and U7610 (N_7610,N_3739,N_3484);
xnor U7611 (N_7611,N_5446,N_3060);
or U7612 (N_7612,N_5979,N_4700);
or U7613 (N_7613,N_5273,N_5417);
nor U7614 (N_7614,N_5578,N_3589);
nor U7615 (N_7615,N_3556,N_4005);
or U7616 (N_7616,N_3839,N_3917);
and U7617 (N_7617,N_3378,N_3311);
and U7618 (N_7618,N_4725,N_3232);
nor U7619 (N_7619,N_5514,N_3864);
and U7620 (N_7620,N_4468,N_3181);
or U7621 (N_7621,N_3975,N_4956);
and U7622 (N_7622,N_5615,N_4806);
nand U7623 (N_7623,N_4781,N_5742);
nor U7624 (N_7624,N_4176,N_3518);
or U7625 (N_7625,N_5508,N_5993);
or U7626 (N_7626,N_5917,N_4074);
xnor U7627 (N_7627,N_4001,N_4277);
or U7628 (N_7628,N_4068,N_4897);
and U7629 (N_7629,N_3927,N_4831);
nor U7630 (N_7630,N_4873,N_4157);
or U7631 (N_7631,N_3896,N_3786);
nand U7632 (N_7632,N_5578,N_3112);
and U7633 (N_7633,N_3149,N_5625);
nor U7634 (N_7634,N_3509,N_5495);
and U7635 (N_7635,N_5557,N_5925);
nor U7636 (N_7636,N_5132,N_4501);
or U7637 (N_7637,N_3702,N_3042);
nor U7638 (N_7638,N_5897,N_3811);
and U7639 (N_7639,N_5505,N_5736);
nand U7640 (N_7640,N_3683,N_4809);
and U7641 (N_7641,N_5151,N_5299);
and U7642 (N_7642,N_4236,N_5907);
nor U7643 (N_7643,N_4961,N_4619);
or U7644 (N_7644,N_4887,N_5982);
or U7645 (N_7645,N_3078,N_5370);
or U7646 (N_7646,N_3683,N_5967);
and U7647 (N_7647,N_4404,N_3959);
nand U7648 (N_7648,N_5580,N_3341);
nand U7649 (N_7649,N_3095,N_5198);
nor U7650 (N_7650,N_3694,N_3503);
or U7651 (N_7651,N_5703,N_4580);
nor U7652 (N_7652,N_4473,N_3549);
and U7653 (N_7653,N_4141,N_4945);
and U7654 (N_7654,N_4232,N_3340);
and U7655 (N_7655,N_3065,N_4619);
nand U7656 (N_7656,N_3929,N_3934);
and U7657 (N_7657,N_4795,N_5195);
xnor U7658 (N_7658,N_3350,N_5192);
or U7659 (N_7659,N_4116,N_4966);
or U7660 (N_7660,N_3561,N_4964);
or U7661 (N_7661,N_5381,N_4334);
nor U7662 (N_7662,N_3630,N_3181);
and U7663 (N_7663,N_4446,N_4531);
nor U7664 (N_7664,N_3255,N_4454);
nand U7665 (N_7665,N_5154,N_3288);
and U7666 (N_7666,N_4948,N_5398);
xnor U7667 (N_7667,N_5585,N_4161);
nand U7668 (N_7668,N_5983,N_5729);
and U7669 (N_7669,N_4097,N_5928);
nand U7670 (N_7670,N_4015,N_5271);
nor U7671 (N_7671,N_4814,N_3820);
or U7672 (N_7672,N_5860,N_4026);
nand U7673 (N_7673,N_4058,N_4146);
and U7674 (N_7674,N_3943,N_5094);
nor U7675 (N_7675,N_3867,N_5485);
and U7676 (N_7676,N_4038,N_4735);
nor U7677 (N_7677,N_4368,N_5823);
and U7678 (N_7678,N_5515,N_3110);
xor U7679 (N_7679,N_3840,N_4384);
or U7680 (N_7680,N_3753,N_3514);
nand U7681 (N_7681,N_4947,N_5291);
and U7682 (N_7682,N_4327,N_5164);
or U7683 (N_7683,N_4381,N_4716);
and U7684 (N_7684,N_3504,N_3460);
and U7685 (N_7685,N_3067,N_3327);
or U7686 (N_7686,N_4289,N_4487);
nand U7687 (N_7687,N_5702,N_5532);
nor U7688 (N_7688,N_3335,N_3913);
nor U7689 (N_7689,N_3031,N_5582);
and U7690 (N_7690,N_4301,N_5763);
nand U7691 (N_7691,N_3074,N_5043);
and U7692 (N_7692,N_4024,N_3587);
or U7693 (N_7693,N_5248,N_5553);
and U7694 (N_7694,N_3328,N_4811);
nand U7695 (N_7695,N_3365,N_4052);
nor U7696 (N_7696,N_5746,N_4804);
or U7697 (N_7697,N_3478,N_3693);
and U7698 (N_7698,N_3055,N_5166);
nand U7699 (N_7699,N_5851,N_4050);
and U7700 (N_7700,N_4810,N_4637);
nor U7701 (N_7701,N_5507,N_3946);
or U7702 (N_7702,N_4846,N_4033);
nor U7703 (N_7703,N_4730,N_5129);
xor U7704 (N_7704,N_4916,N_4832);
nor U7705 (N_7705,N_5459,N_4004);
or U7706 (N_7706,N_5017,N_4505);
nand U7707 (N_7707,N_4896,N_4781);
and U7708 (N_7708,N_5791,N_3657);
nand U7709 (N_7709,N_3108,N_4149);
nor U7710 (N_7710,N_5274,N_3848);
or U7711 (N_7711,N_3600,N_5196);
nand U7712 (N_7712,N_4781,N_4585);
or U7713 (N_7713,N_5927,N_3563);
nor U7714 (N_7714,N_5663,N_5052);
or U7715 (N_7715,N_4788,N_4747);
nor U7716 (N_7716,N_5503,N_3213);
and U7717 (N_7717,N_3927,N_5838);
and U7718 (N_7718,N_3639,N_5694);
or U7719 (N_7719,N_3160,N_5486);
nand U7720 (N_7720,N_4439,N_4320);
nor U7721 (N_7721,N_3030,N_3773);
nor U7722 (N_7722,N_3703,N_4663);
or U7723 (N_7723,N_4537,N_5958);
and U7724 (N_7724,N_5615,N_3863);
nand U7725 (N_7725,N_3546,N_4118);
or U7726 (N_7726,N_5900,N_3131);
or U7727 (N_7727,N_4032,N_5446);
nor U7728 (N_7728,N_4129,N_5649);
nor U7729 (N_7729,N_5375,N_3243);
nand U7730 (N_7730,N_5369,N_4435);
nor U7731 (N_7731,N_5541,N_5834);
nor U7732 (N_7732,N_5455,N_5922);
and U7733 (N_7733,N_4766,N_5078);
nor U7734 (N_7734,N_4053,N_4137);
and U7735 (N_7735,N_3077,N_5738);
or U7736 (N_7736,N_5367,N_5255);
and U7737 (N_7737,N_3648,N_4656);
or U7738 (N_7738,N_4790,N_3736);
nand U7739 (N_7739,N_3625,N_3668);
nand U7740 (N_7740,N_5515,N_4628);
or U7741 (N_7741,N_3866,N_4342);
and U7742 (N_7742,N_5899,N_4037);
or U7743 (N_7743,N_3142,N_3945);
and U7744 (N_7744,N_5007,N_3993);
nor U7745 (N_7745,N_3800,N_4651);
nand U7746 (N_7746,N_4933,N_5183);
nand U7747 (N_7747,N_4999,N_4923);
nor U7748 (N_7748,N_3690,N_4996);
nor U7749 (N_7749,N_3909,N_5323);
nand U7750 (N_7750,N_3732,N_5051);
nand U7751 (N_7751,N_5289,N_4794);
nor U7752 (N_7752,N_3731,N_3922);
nand U7753 (N_7753,N_3369,N_4086);
nor U7754 (N_7754,N_3957,N_3599);
or U7755 (N_7755,N_5379,N_4652);
nor U7756 (N_7756,N_4804,N_5619);
and U7757 (N_7757,N_5602,N_3481);
and U7758 (N_7758,N_4339,N_5275);
and U7759 (N_7759,N_4456,N_5639);
nand U7760 (N_7760,N_3710,N_4971);
nor U7761 (N_7761,N_5759,N_3227);
nor U7762 (N_7762,N_5354,N_5378);
nor U7763 (N_7763,N_4557,N_4982);
and U7764 (N_7764,N_5215,N_5116);
nor U7765 (N_7765,N_4970,N_4624);
nor U7766 (N_7766,N_5934,N_5117);
and U7767 (N_7767,N_4098,N_5902);
and U7768 (N_7768,N_4837,N_3335);
and U7769 (N_7769,N_4873,N_5105);
or U7770 (N_7770,N_3287,N_4955);
and U7771 (N_7771,N_4111,N_3882);
nor U7772 (N_7772,N_3462,N_5805);
nor U7773 (N_7773,N_5994,N_4715);
nand U7774 (N_7774,N_4390,N_5262);
nand U7775 (N_7775,N_3130,N_5916);
or U7776 (N_7776,N_5268,N_5947);
nor U7777 (N_7777,N_5545,N_5339);
and U7778 (N_7778,N_3842,N_5636);
or U7779 (N_7779,N_5569,N_4780);
nand U7780 (N_7780,N_3880,N_3257);
and U7781 (N_7781,N_3217,N_3566);
nand U7782 (N_7782,N_3295,N_4300);
or U7783 (N_7783,N_5333,N_5859);
nand U7784 (N_7784,N_3224,N_5192);
nor U7785 (N_7785,N_3732,N_5047);
nand U7786 (N_7786,N_4869,N_3221);
and U7787 (N_7787,N_5957,N_5722);
and U7788 (N_7788,N_4200,N_3617);
xor U7789 (N_7789,N_5772,N_5203);
nand U7790 (N_7790,N_3928,N_3598);
nor U7791 (N_7791,N_5143,N_3515);
and U7792 (N_7792,N_4186,N_4370);
nand U7793 (N_7793,N_5166,N_3510);
nand U7794 (N_7794,N_4005,N_3819);
and U7795 (N_7795,N_4041,N_5786);
and U7796 (N_7796,N_4925,N_5124);
and U7797 (N_7797,N_3000,N_3584);
and U7798 (N_7798,N_3932,N_4097);
nor U7799 (N_7799,N_4841,N_3154);
nand U7800 (N_7800,N_4902,N_3551);
and U7801 (N_7801,N_5341,N_3041);
nor U7802 (N_7802,N_5329,N_5515);
or U7803 (N_7803,N_5938,N_5773);
or U7804 (N_7804,N_3131,N_3747);
nor U7805 (N_7805,N_3481,N_3217);
nand U7806 (N_7806,N_3967,N_3408);
and U7807 (N_7807,N_3498,N_3143);
nor U7808 (N_7808,N_3363,N_3137);
or U7809 (N_7809,N_4972,N_4059);
or U7810 (N_7810,N_5559,N_4766);
nand U7811 (N_7811,N_3442,N_3963);
or U7812 (N_7812,N_4544,N_3020);
and U7813 (N_7813,N_4874,N_4387);
and U7814 (N_7814,N_3301,N_3211);
and U7815 (N_7815,N_4891,N_3725);
and U7816 (N_7816,N_5066,N_4536);
nand U7817 (N_7817,N_4590,N_4035);
or U7818 (N_7818,N_4300,N_5047);
nor U7819 (N_7819,N_4810,N_5152);
or U7820 (N_7820,N_3939,N_3296);
nand U7821 (N_7821,N_4286,N_4552);
nor U7822 (N_7822,N_3523,N_5380);
nor U7823 (N_7823,N_3184,N_4696);
and U7824 (N_7824,N_5592,N_5902);
xor U7825 (N_7825,N_4262,N_4195);
or U7826 (N_7826,N_3317,N_5280);
or U7827 (N_7827,N_3223,N_3889);
and U7828 (N_7828,N_3512,N_5984);
or U7829 (N_7829,N_4689,N_5786);
or U7830 (N_7830,N_5931,N_5883);
nand U7831 (N_7831,N_5645,N_3741);
or U7832 (N_7832,N_5543,N_3454);
nor U7833 (N_7833,N_5591,N_4197);
nor U7834 (N_7834,N_3095,N_5106);
and U7835 (N_7835,N_5645,N_5703);
and U7836 (N_7836,N_4495,N_4889);
or U7837 (N_7837,N_5409,N_4126);
nand U7838 (N_7838,N_4248,N_4904);
or U7839 (N_7839,N_4676,N_5512);
or U7840 (N_7840,N_5118,N_3064);
nand U7841 (N_7841,N_4449,N_5596);
nor U7842 (N_7842,N_4324,N_4225);
nand U7843 (N_7843,N_3529,N_3879);
nand U7844 (N_7844,N_5868,N_3460);
nand U7845 (N_7845,N_4904,N_5836);
nand U7846 (N_7846,N_3747,N_3945);
and U7847 (N_7847,N_3982,N_5260);
nor U7848 (N_7848,N_4311,N_4809);
and U7849 (N_7849,N_5445,N_4569);
or U7850 (N_7850,N_4583,N_3509);
and U7851 (N_7851,N_3847,N_3189);
and U7852 (N_7852,N_4660,N_5512);
nand U7853 (N_7853,N_5041,N_5923);
and U7854 (N_7854,N_3458,N_3300);
nor U7855 (N_7855,N_3919,N_3152);
or U7856 (N_7856,N_5707,N_4444);
nand U7857 (N_7857,N_5429,N_5107);
or U7858 (N_7858,N_5717,N_5701);
or U7859 (N_7859,N_5432,N_5764);
nor U7860 (N_7860,N_4731,N_4331);
nand U7861 (N_7861,N_5683,N_4670);
or U7862 (N_7862,N_5041,N_5325);
xor U7863 (N_7863,N_3476,N_5996);
nor U7864 (N_7864,N_3470,N_4649);
xnor U7865 (N_7865,N_3242,N_3569);
nand U7866 (N_7866,N_3124,N_5274);
nand U7867 (N_7867,N_5141,N_5681);
nand U7868 (N_7868,N_5125,N_5609);
nor U7869 (N_7869,N_3491,N_4230);
or U7870 (N_7870,N_4123,N_5186);
and U7871 (N_7871,N_5332,N_4974);
or U7872 (N_7872,N_4128,N_4816);
or U7873 (N_7873,N_5324,N_3212);
or U7874 (N_7874,N_4190,N_3532);
or U7875 (N_7875,N_3459,N_4431);
or U7876 (N_7876,N_3606,N_4585);
nand U7877 (N_7877,N_3520,N_3670);
or U7878 (N_7878,N_5235,N_4312);
nand U7879 (N_7879,N_4566,N_5916);
nand U7880 (N_7880,N_3009,N_4250);
or U7881 (N_7881,N_3678,N_5072);
nor U7882 (N_7882,N_5576,N_4826);
nor U7883 (N_7883,N_4379,N_3720);
or U7884 (N_7884,N_3583,N_5404);
and U7885 (N_7885,N_5313,N_5806);
nor U7886 (N_7886,N_3237,N_3657);
nand U7887 (N_7887,N_4346,N_3223);
or U7888 (N_7888,N_3191,N_5395);
or U7889 (N_7889,N_4577,N_4765);
and U7890 (N_7890,N_4344,N_4607);
or U7891 (N_7891,N_3234,N_4123);
and U7892 (N_7892,N_4013,N_3140);
or U7893 (N_7893,N_4747,N_4604);
nor U7894 (N_7894,N_3574,N_4679);
nand U7895 (N_7895,N_5689,N_3195);
or U7896 (N_7896,N_4464,N_4865);
or U7897 (N_7897,N_5831,N_4015);
or U7898 (N_7898,N_5803,N_5209);
nand U7899 (N_7899,N_5687,N_5994);
nand U7900 (N_7900,N_3189,N_3386);
or U7901 (N_7901,N_3958,N_5987);
or U7902 (N_7902,N_4219,N_4385);
or U7903 (N_7903,N_5261,N_4246);
and U7904 (N_7904,N_5089,N_5927);
and U7905 (N_7905,N_3555,N_3703);
nand U7906 (N_7906,N_5796,N_5864);
nor U7907 (N_7907,N_3314,N_5780);
nand U7908 (N_7908,N_4836,N_4694);
and U7909 (N_7909,N_5500,N_4375);
nor U7910 (N_7910,N_5875,N_4880);
and U7911 (N_7911,N_4764,N_4800);
nor U7912 (N_7912,N_5821,N_5721);
or U7913 (N_7913,N_5643,N_4652);
nor U7914 (N_7914,N_4012,N_4009);
and U7915 (N_7915,N_4844,N_3121);
nand U7916 (N_7916,N_5678,N_3829);
nor U7917 (N_7917,N_3646,N_3958);
xnor U7918 (N_7918,N_4076,N_5397);
and U7919 (N_7919,N_3001,N_5106);
and U7920 (N_7920,N_5038,N_3418);
xor U7921 (N_7921,N_3098,N_4034);
nand U7922 (N_7922,N_3430,N_3687);
nor U7923 (N_7923,N_4546,N_3689);
nand U7924 (N_7924,N_4424,N_5301);
nand U7925 (N_7925,N_3430,N_3922);
or U7926 (N_7926,N_4864,N_5762);
and U7927 (N_7927,N_3426,N_4101);
nor U7928 (N_7928,N_3095,N_3692);
nor U7929 (N_7929,N_5909,N_5200);
nand U7930 (N_7930,N_5960,N_3840);
xor U7931 (N_7931,N_5374,N_5727);
or U7932 (N_7932,N_3284,N_4645);
nand U7933 (N_7933,N_3726,N_4621);
nand U7934 (N_7934,N_4291,N_4384);
and U7935 (N_7935,N_3563,N_5332);
or U7936 (N_7936,N_4846,N_3123);
nand U7937 (N_7937,N_4549,N_3615);
nand U7938 (N_7938,N_4192,N_4327);
and U7939 (N_7939,N_4653,N_3969);
and U7940 (N_7940,N_5895,N_5521);
and U7941 (N_7941,N_3215,N_5908);
nand U7942 (N_7942,N_3533,N_5773);
nand U7943 (N_7943,N_5468,N_3621);
nor U7944 (N_7944,N_4771,N_3050);
nor U7945 (N_7945,N_3625,N_3636);
and U7946 (N_7946,N_3552,N_5109);
nor U7947 (N_7947,N_4907,N_4433);
and U7948 (N_7948,N_5213,N_5761);
nor U7949 (N_7949,N_4799,N_5752);
or U7950 (N_7950,N_4622,N_4398);
and U7951 (N_7951,N_5108,N_4700);
nor U7952 (N_7952,N_4626,N_5714);
nand U7953 (N_7953,N_3029,N_5293);
nand U7954 (N_7954,N_4008,N_5003);
and U7955 (N_7955,N_4664,N_4196);
nor U7956 (N_7956,N_3734,N_4136);
nand U7957 (N_7957,N_5150,N_5363);
and U7958 (N_7958,N_4792,N_5769);
nor U7959 (N_7959,N_4513,N_3654);
or U7960 (N_7960,N_4068,N_3401);
and U7961 (N_7961,N_3116,N_3471);
nand U7962 (N_7962,N_5255,N_3710);
nand U7963 (N_7963,N_3069,N_3315);
or U7964 (N_7964,N_4926,N_4641);
nand U7965 (N_7965,N_5890,N_4698);
and U7966 (N_7966,N_3817,N_3557);
or U7967 (N_7967,N_3273,N_3857);
or U7968 (N_7968,N_4943,N_3894);
or U7969 (N_7969,N_5005,N_4361);
and U7970 (N_7970,N_5988,N_4355);
nor U7971 (N_7971,N_3438,N_3242);
or U7972 (N_7972,N_4785,N_3737);
nand U7973 (N_7973,N_5088,N_5200);
nor U7974 (N_7974,N_3110,N_4139);
nor U7975 (N_7975,N_3632,N_5254);
and U7976 (N_7976,N_4489,N_5391);
and U7977 (N_7977,N_3395,N_4332);
nor U7978 (N_7978,N_3756,N_3493);
or U7979 (N_7979,N_3036,N_4237);
or U7980 (N_7980,N_4279,N_3056);
nor U7981 (N_7981,N_3877,N_4247);
nand U7982 (N_7982,N_3139,N_4803);
or U7983 (N_7983,N_5844,N_4678);
nor U7984 (N_7984,N_3433,N_3229);
nor U7985 (N_7985,N_5994,N_4726);
nand U7986 (N_7986,N_4437,N_4933);
xnor U7987 (N_7987,N_3105,N_5347);
or U7988 (N_7988,N_5256,N_4881);
nor U7989 (N_7989,N_3811,N_3636);
or U7990 (N_7990,N_5125,N_4778);
and U7991 (N_7991,N_3421,N_4265);
nand U7992 (N_7992,N_5027,N_4358);
and U7993 (N_7993,N_5346,N_4589);
nand U7994 (N_7994,N_5979,N_5593);
nor U7995 (N_7995,N_5682,N_3925);
and U7996 (N_7996,N_3596,N_4118);
and U7997 (N_7997,N_5235,N_5574);
nand U7998 (N_7998,N_5588,N_5493);
or U7999 (N_7999,N_5390,N_3134);
nor U8000 (N_8000,N_4299,N_3485);
xnor U8001 (N_8001,N_3664,N_3207);
nand U8002 (N_8002,N_4019,N_4147);
nor U8003 (N_8003,N_3985,N_3587);
or U8004 (N_8004,N_4184,N_4666);
or U8005 (N_8005,N_3401,N_3035);
or U8006 (N_8006,N_4298,N_3419);
nor U8007 (N_8007,N_3182,N_3886);
nor U8008 (N_8008,N_3826,N_4823);
or U8009 (N_8009,N_5868,N_4118);
xnor U8010 (N_8010,N_5868,N_3660);
or U8011 (N_8011,N_4354,N_5240);
or U8012 (N_8012,N_4858,N_3400);
nor U8013 (N_8013,N_4370,N_4327);
or U8014 (N_8014,N_4185,N_3191);
and U8015 (N_8015,N_4780,N_4174);
nor U8016 (N_8016,N_4010,N_5490);
or U8017 (N_8017,N_4918,N_5993);
nor U8018 (N_8018,N_4521,N_3537);
nor U8019 (N_8019,N_4399,N_3155);
or U8020 (N_8020,N_5963,N_5620);
and U8021 (N_8021,N_4160,N_4373);
and U8022 (N_8022,N_3889,N_4757);
nor U8023 (N_8023,N_4406,N_5474);
or U8024 (N_8024,N_4516,N_3245);
or U8025 (N_8025,N_4219,N_5501);
and U8026 (N_8026,N_4550,N_5082);
or U8027 (N_8027,N_4582,N_4455);
nor U8028 (N_8028,N_5406,N_5524);
nor U8029 (N_8029,N_3006,N_3343);
nand U8030 (N_8030,N_3313,N_4931);
nand U8031 (N_8031,N_5377,N_3254);
nor U8032 (N_8032,N_4837,N_5574);
nor U8033 (N_8033,N_3660,N_5692);
or U8034 (N_8034,N_3855,N_3397);
xor U8035 (N_8035,N_5588,N_4180);
and U8036 (N_8036,N_3462,N_3445);
or U8037 (N_8037,N_4052,N_5686);
or U8038 (N_8038,N_5676,N_5386);
or U8039 (N_8039,N_5478,N_5200);
or U8040 (N_8040,N_4992,N_4824);
or U8041 (N_8041,N_4581,N_5833);
nand U8042 (N_8042,N_5348,N_5177);
nand U8043 (N_8043,N_5930,N_3830);
nand U8044 (N_8044,N_3425,N_3157);
nor U8045 (N_8045,N_5581,N_3767);
or U8046 (N_8046,N_3288,N_5763);
and U8047 (N_8047,N_3725,N_4578);
nor U8048 (N_8048,N_5173,N_4005);
nor U8049 (N_8049,N_5514,N_5679);
and U8050 (N_8050,N_4365,N_4820);
and U8051 (N_8051,N_4927,N_3462);
or U8052 (N_8052,N_3624,N_4376);
and U8053 (N_8053,N_4397,N_5631);
nor U8054 (N_8054,N_3178,N_3885);
and U8055 (N_8055,N_4181,N_4606);
nand U8056 (N_8056,N_3728,N_4212);
nor U8057 (N_8057,N_4419,N_3429);
or U8058 (N_8058,N_5955,N_4314);
nand U8059 (N_8059,N_4924,N_5195);
and U8060 (N_8060,N_5590,N_3060);
and U8061 (N_8061,N_4408,N_3061);
nor U8062 (N_8062,N_5222,N_4836);
or U8063 (N_8063,N_3388,N_5879);
nand U8064 (N_8064,N_3405,N_4904);
and U8065 (N_8065,N_4569,N_3700);
or U8066 (N_8066,N_3898,N_4674);
nor U8067 (N_8067,N_5426,N_3023);
and U8068 (N_8068,N_4768,N_5507);
and U8069 (N_8069,N_5244,N_3671);
nand U8070 (N_8070,N_5025,N_3110);
and U8071 (N_8071,N_5785,N_4823);
and U8072 (N_8072,N_4228,N_5761);
nand U8073 (N_8073,N_3575,N_5156);
or U8074 (N_8074,N_3367,N_3077);
nor U8075 (N_8075,N_4277,N_4984);
nor U8076 (N_8076,N_3190,N_4255);
and U8077 (N_8077,N_4515,N_4448);
nor U8078 (N_8078,N_4155,N_4455);
and U8079 (N_8079,N_4988,N_3635);
or U8080 (N_8080,N_5795,N_5546);
nor U8081 (N_8081,N_3974,N_4058);
nor U8082 (N_8082,N_4266,N_4836);
or U8083 (N_8083,N_4808,N_4285);
nand U8084 (N_8084,N_4277,N_5489);
nor U8085 (N_8085,N_5561,N_3506);
nor U8086 (N_8086,N_3272,N_5337);
nor U8087 (N_8087,N_5893,N_4572);
or U8088 (N_8088,N_3117,N_4903);
and U8089 (N_8089,N_3360,N_4915);
or U8090 (N_8090,N_4887,N_3055);
or U8091 (N_8091,N_4847,N_4550);
or U8092 (N_8092,N_4193,N_3038);
nor U8093 (N_8093,N_4037,N_5663);
nand U8094 (N_8094,N_4783,N_5691);
nor U8095 (N_8095,N_3134,N_3054);
nand U8096 (N_8096,N_3180,N_4369);
nand U8097 (N_8097,N_3682,N_4864);
or U8098 (N_8098,N_5602,N_4001);
nand U8099 (N_8099,N_5207,N_4059);
or U8100 (N_8100,N_3723,N_4503);
or U8101 (N_8101,N_4351,N_3139);
nor U8102 (N_8102,N_5972,N_5014);
and U8103 (N_8103,N_3939,N_5440);
nand U8104 (N_8104,N_3720,N_3431);
nand U8105 (N_8105,N_4389,N_5304);
nand U8106 (N_8106,N_5938,N_5004);
nand U8107 (N_8107,N_3490,N_4541);
and U8108 (N_8108,N_4480,N_5227);
nor U8109 (N_8109,N_4678,N_5285);
or U8110 (N_8110,N_5157,N_4217);
or U8111 (N_8111,N_4461,N_3521);
nor U8112 (N_8112,N_3100,N_4788);
nor U8113 (N_8113,N_5512,N_5461);
and U8114 (N_8114,N_5917,N_4271);
or U8115 (N_8115,N_5496,N_5429);
and U8116 (N_8116,N_5973,N_5243);
and U8117 (N_8117,N_3734,N_3632);
nor U8118 (N_8118,N_3834,N_5240);
nand U8119 (N_8119,N_3706,N_3785);
or U8120 (N_8120,N_4579,N_3247);
nand U8121 (N_8121,N_3043,N_5536);
and U8122 (N_8122,N_3609,N_4846);
or U8123 (N_8123,N_4392,N_4093);
nand U8124 (N_8124,N_4410,N_3977);
nor U8125 (N_8125,N_4173,N_5176);
and U8126 (N_8126,N_3417,N_3753);
nand U8127 (N_8127,N_3003,N_5337);
and U8128 (N_8128,N_4876,N_3431);
nand U8129 (N_8129,N_4859,N_4209);
nor U8130 (N_8130,N_3303,N_3821);
nor U8131 (N_8131,N_3397,N_4436);
and U8132 (N_8132,N_5041,N_3674);
or U8133 (N_8133,N_5147,N_4869);
nand U8134 (N_8134,N_4764,N_3621);
or U8135 (N_8135,N_4419,N_3683);
and U8136 (N_8136,N_3565,N_3385);
or U8137 (N_8137,N_5873,N_4335);
and U8138 (N_8138,N_4454,N_5251);
or U8139 (N_8139,N_4374,N_5398);
or U8140 (N_8140,N_4973,N_5209);
and U8141 (N_8141,N_3918,N_4439);
or U8142 (N_8142,N_5452,N_5152);
and U8143 (N_8143,N_4827,N_4939);
and U8144 (N_8144,N_5242,N_5306);
nor U8145 (N_8145,N_3698,N_4624);
nor U8146 (N_8146,N_4037,N_5801);
nor U8147 (N_8147,N_3483,N_3380);
nor U8148 (N_8148,N_3510,N_5917);
nand U8149 (N_8149,N_5655,N_3478);
nand U8150 (N_8150,N_3372,N_3412);
and U8151 (N_8151,N_3550,N_4776);
and U8152 (N_8152,N_5747,N_3762);
or U8153 (N_8153,N_4671,N_5068);
nor U8154 (N_8154,N_3619,N_3543);
nor U8155 (N_8155,N_3882,N_5152);
and U8156 (N_8156,N_3000,N_4392);
nand U8157 (N_8157,N_3825,N_3150);
nand U8158 (N_8158,N_3946,N_3351);
nand U8159 (N_8159,N_4282,N_4249);
and U8160 (N_8160,N_5210,N_3032);
and U8161 (N_8161,N_3858,N_3955);
nor U8162 (N_8162,N_4583,N_3283);
nand U8163 (N_8163,N_4108,N_5849);
or U8164 (N_8164,N_4357,N_3374);
and U8165 (N_8165,N_4726,N_3827);
or U8166 (N_8166,N_4790,N_5359);
and U8167 (N_8167,N_4279,N_5174);
or U8168 (N_8168,N_5928,N_4555);
nor U8169 (N_8169,N_5326,N_3789);
nor U8170 (N_8170,N_3993,N_4739);
and U8171 (N_8171,N_3022,N_5235);
or U8172 (N_8172,N_4538,N_3688);
and U8173 (N_8173,N_5929,N_3899);
or U8174 (N_8174,N_4191,N_3838);
nor U8175 (N_8175,N_5900,N_5475);
or U8176 (N_8176,N_4546,N_3847);
nor U8177 (N_8177,N_5698,N_5125);
nand U8178 (N_8178,N_3730,N_3968);
and U8179 (N_8179,N_5192,N_5437);
nand U8180 (N_8180,N_3090,N_3070);
nor U8181 (N_8181,N_3538,N_4565);
and U8182 (N_8182,N_5784,N_4375);
and U8183 (N_8183,N_5517,N_5891);
xor U8184 (N_8184,N_3860,N_5714);
nand U8185 (N_8185,N_5727,N_4619);
or U8186 (N_8186,N_5243,N_4467);
nor U8187 (N_8187,N_5688,N_4372);
and U8188 (N_8188,N_4993,N_5163);
or U8189 (N_8189,N_3282,N_4378);
and U8190 (N_8190,N_3855,N_4846);
nand U8191 (N_8191,N_3566,N_4761);
and U8192 (N_8192,N_4949,N_5739);
nor U8193 (N_8193,N_3308,N_4928);
and U8194 (N_8194,N_4023,N_3440);
or U8195 (N_8195,N_4258,N_4295);
or U8196 (N_8196,N_4428,N_4478);
nor U8197 (N_8197,N_5944,N_4011);
and U8198 (N_8198,N_5770,N_5805);
and U8199 (N_8199,N_4180,N_3880);
nor U8200 (N_8200,N_4491,N_3049);
nand U8201 (N_8201,N_4030,N_3050);
nand U8202 (N_8202,N_5318,N_3533);
and U8203 (N_8203,N_3281,N_4106);
and U8204 (N_8204,N_4672,N_3124);
nand U8205 (N_8205,N_4881,N_3087);
or U8206 (N_8206,N_5504,N_4855);
and U8207 (N_8207,N_5599,N_5520);
or U8208 (N_8208,N_4799,N_5716);
and U8209 (N_8209,N_3709,N_4660);
or U8210 (N_8210,N_5484,N_4527);
nand U8211 (N_8211,N_4880,N_3904);
nand U8212 (N_8212,N_4133,N_4764);
nand U8213 (N_8213,N_4262,N_3357);
nand U8214 (N_8214,N_4979,N_5884);
and U8215 (N_8215,N_5211,N_4455);
nand U8216 (N_8216,N_4711,N_5889);
nor U8217 (N_8217,N_3046,N_5379);
or U8218 (N_8218,N_5976,N_3419);
or U8219 (N_8219,N_4325,N_3151);
or U8220 (N_8220,N_4568,N_4148);
nand U8221 (N_8221,N_5970,N_5083);
nand U8222 (N_8222,N_4576,N_5099);
and U8223 (N_8223,N_5453,N_4367);
or U8224 (N_8224,N_5406,N_4896);
nor U8225 (N_8225,N_4313,N_5230);
and U8226 (N_8226,N_5781,N_5933);
or U8227 (N_8227,N_5795,N_3702);
nor U8228 (N_8228,N_3773,N_3080);
and U8229 (N_8229,N_3920,N_5534);
or U8230 (N_8230,N_4785,N_5053);
or U8231 (N_8231,N_5890,N_4532);
or U8232 (N_8232,N_4156,N_5825);
and U8233 (N_8233,N_5718,N_4669);
nand U8234 (N_8234,N_4721,N_3651);
or U8235 (N_8235,N_3699,N_3282);
or U8236 (N_8236,N_5646,N_4616);
and U8237 (N_8237,N_4005,N_4612);
or U8238 (N_8238,N_5850,N_5763);
nand U8239 (N_8239,N_5121,N_3161);
nor U8240 (N_8240,N_3911,N_5668);
nand U8241 (N_8241,N_3167,N_4592);
or U8242 (N_8242,N_4354,N_5378);
nand U8243 (N_8243,N_4005,N_4644);
nor U8244 (N_8244,N_4549,N_3461);
nand U8245 (N_8245,N_5132,N_5400);
and U8246 (N_8246,N_3428,N_5304);
nor U8247 (N_8247,N_3729,N_3569);
nand U8248 (N_8248,N_4151,N_4860);
xnor U8249 (N_8249,N_4315,N_3154);
and U8250 (N_8250,N_3095,N_4631);
and U8251 (N_8251,N_5036,N_5499);
nor U8252 (N_8252,N_5187,N_5199);
or U8253 (N_8253,N_5301,N_3046);
nand U8254 (N_8254,N_3840,N_5169);
and U8255 (N_8255,N_3421,N_3411);
xnor U8256 (N_8256,N_4315,N_4714);
nor U8257 (N_8257,N_3686,N_3871);
nor U8258 (N_8258,N_5619,N_3601);
nor U8259 (N_8259,N_3685,N_4022);
or U8260 (N_8260,N_4838,N_5961);
and U8261 (N_8261,N_3547,N_4903);
nor U8262 (N_8262,N_3903,N_3559);
nor U8263 (N_8263,N_4315,N_5433);
nor U8264 (N_8264,N_4237,N_3605);
and U8265 (N_8265,N_4288,N_3775);
and U8266 (N_8266,N_4123,N_3502);
nand U8267 (N_8267,N_3275,N_5576);
nand U8268 (N_8268,N_3106,N_5026);
nand U8269 (N_8269,N_4356,N_4390);
or U8270 (N_8270,N_4209,N_5592);
or U8271 (N_8271,N_3555,N_3578);
or U8272 (N_8272,N_4181,N_4952);
nand U8273 (N_8273,N_3797,N_3401);
nand U8274 (N_8274,N_5022,N_3731);
nand U8275 (N_8275,N_4918,N_4778);
or U8276 (N_8276,N_4451,N_5755);
nor U8277 (N_8277,N_5355,N_5490);
and U8278 (N_8278,N_5961,N_5814);
or U8279 (N_8279,N_5626,N_5263);
or U8280 (N_8280,N_4216,N_3880);
and U8281 (N_8281,N_3007,N_5483);
nor U8282 (N_8282,N_3658,N_4615);
nor U8283 (N_8283,N_3196,N_5047);
nor U8284 (N_8284,N_4327,N_4556);
and U8285 (N_8285,N_4161,N_4291);
and U8286 (N_8286,N_4135,N_5690);
and U8287 (N_8287,N_3258,N_3074);
nand U8288 (N_8288,N_4488,N_5111);
nand U8289 (N_8289,N_5067,N_4471);
and U8290 (N_8290,N_5582,N_4471);
nand U8291 (N_8291,N_5149,N_5240);
and U8292 (N_8292,N_5585,N_3171);
nor U8293 (N_8293,N_4063,N_5834);
xnor U8294 (N_8294,N_5466,N_3234);
or U8295 (N_8295,N_4464,N_5649);
nor U8296 (N_8296,N_4915,N_3658);
nor U8297 (N_8297,N_4315,N_5536);
and U8298 (N_8298,N_4725,N_4530);
and U8299 (N_8299,N_5570,N_5751);
or U8300 (N_8300,N_3645,N_4407);
nand U8301 (N_8301,N_5475,N_5644);
nand U8302 (N_8302,N_5583,N_4476);
nor U8303 (N_8303,N_4225,N_4741);
nand U8304 (N_8304,N_3915,N_3783);
or U8305 (N_8305,N_3819,N_4670);
nand U8306 (N_8306,N_3446,N_3439);
and U8307 (N_8307,N_4064,N_3567);
or U8308 (N_8308,N_5938,N_5647);
nor U8309 (N_8309,N_3916,N_3947);
or U8310 (N_8310,N_5655,N_3364);
and U8311 (N_8311,N_4151,N_4680);
nand U8312 (N_8312,N_3322,N_4607);
and U8313 (N_8313,N_4227,N_3487);
nand U8314 (N_8314,N_5947,N_4627);
or U8315 (N_8315,N_3241,N_4840);
nand U8316 (N_8316,N_5204,N_3080);
or U8317 (N_8317,N_5648,N_4248);
nand U8318 (N_8318,N_5144,N_5006);
nand U8319 (N_8319,N_5920,N_3758);
nand U8320 (N_8320,N_4635,N_5007);
nand U8321 (N_8321,N_4727,N_5883);
nor U8322 (N_8322,N_3571,N_4834);
nor U8323 (N_8323,N_3310,N_4836);
nor U8324 (N_8324,N_4633,N_3866);
and U8325 (N_8325,N_5520,N_4907);
nor U8326 (N_8326,N_5549,N_5053);
and U8327 (N_8327,N_5112,N_3132);
nand U8328 (N_8328,N_3126,N_5679);
nand U8329 (N_8329,N_5385,N_4254);
or U8330 (N_8330,N_4667,N_3917);
and U8331 (N_8331,N_5975,N_4127);
nor U8332 (N_8332,N_3368,N_4731);
and U8333 (N_8333,N_4383,N_4624);
nand U8334 (N_8334,N_5146,N_5479);
or U8335 (N_8335,N_3013,N_4835);
nand U8336 (N_8336,N_5629,N_5197);
or U8337 (N_8337,N_5178,N_3698);
nand U8338 (N_8338,N_4009,N_5283);
or U8339 (N_8339,N_4780,N_4720);
nand U8340 (N_8340,N_5173,N_3392);
and U8341 (N_8341,N_4784,N_4480);
and U8342 (N_8342,N_5692,N_4999);
and U8343 (N_8343,N_3060,N_5974);
nor U8344 (N_8344,N_3651,N_5955);
nor U8345 (N_8345,N_4754,N_4709);
nand U8346 (N_8346,N_5153,N_4437);
nor U8347 (N_8347,N_5946,N_5521);
nor U8348 (N_8348,N_5334,N_3046);
nor U8349 (N_8349,N_3732,N_4536);
nand U8350 (N_8350,N_3745,N_5762);
nand U8351 (N_8351,N_3432,N_3051);
nand U8352 (N_8352,N_5738,N_3220);
or U8353 (N_8353,N_3957,N_5642);
nand U8354 (N_8354,N_4580,N_4472);
nand U8355 (N_8355,N_4176,N_5755);
or U8356 (N_8356,N_3929,N_5453);
nor U8357 (N_8357,N_5909,N_5253);
nand U8358 (N_8358,N_3578,N_5492);
or U8359 (N_8359,N_5981,N_4610);
nor U8360 (N_8360,N_4222,N_5493);
nor U8361 (N_8361,N_5440,N_4967);
or U8362 (N_8362,N_5212,N_4625);
or U8363 (N_8363,N_4681,N_4663);
nor U8364 (N_8364,N_3965,N_5468);
and U8365 (N_8365,N_3717,N_4878);
nor U8366 (N_8366,N_5696,N_4435);
nor U8367 (N_8367,N_5684,N_5272);
nand U8368 (N_8368,N_5094,N_3677);
and U8369 (N_8369,N_3671,N_5080);
or U8370 (N_8370,N_3794,N_4017);
nand U8371 (N_8371,N_4934,N_4502);
or U8372 (N_8372,N_4853,N_3870);
nor U8373 (N_8373,N_5082,N_5013);
nand U8374 (N_8374,N_5940,N_5085);
and U8375 (N_8375,N_3170,N_3178);
nand U8376 (N_8376,N_3488,N_4237);
and U8377 (N_8377,N_5320,N_4084);
nor U8378 (N_8378,N_5212,N_5085);
and U8379 (N_8379,N_3539,N_3184);
nor U8380 (N_8380,N_3075,N_3761);
and U8381 (N_8381,N_3279,N_3725);
and U8382 (N_8382,N_3814,N_3343);
or U8383 (N_8383,N_3163,N_5697);
or U8384 (N_8384,N_5148,N_5130);
nand U8385 (N_8385,N_4420,N_3823);
nand U8386 (N_8386,N_5424,N_5724);
or U8387 (N_8387,N_4142,N_3217);
nor U8388 (N_8388,N_5843,N_5307);
nand U8389 (N_8389,N_3482,N_5956);
or U8390 (N_8390,N_4192,N_3009);
or U8391 (N_8391,N_4778,N_4740);
nand U8392 (N_8392,N_3802,N_4700);
nand U8393 (N_8393,N_4313,N_5296);
or U8394 (N_8394,N_5264,N_5801);
nand U8395 (N_8395,N_5351,N_3021);
and U8396 (N_8396,N_4965,N_3907);
or U8397 (N_8397,N_4843,N_5871);
or U8398 (N_8398,N_5262,N_5818);
or U8399 (N_8399,N_4321,N_3678);
nor U8400 (N_8400,N_4702,N_4820);
nor U8401 (N_8401,N_5525,N_4303);
or U8402 (N_8402,N_4970,N_5118);
nand U8403 (N_8403,N_4873,N_4845);
and U8404 (N_8404,N_5951,N_5424);
xor U8405 (N_8405,N_4603,N_5183);
and U8406 (N_8406,N_5880,N_5066);
nor U8407 (N_8407,N_4116,N_3041);
nand U8408 (N_8408,N_3665,N_3712);
and U8409 (N_8409,N_3422,N_5178);
and U8410 (N_8410,N_3282,N_3429);
nand U8411 (N_8411,N_4274,N_4150);
or U8412 (N_8412,N_5806,N_4819);
and U8413 (N_8413,N_3503,N_4949);
and U8414 (N_8414,N_3111,N_3924);
nor U8415 (N_8415,N_4082,N_4849);
and U8416 (N_8416,N_4203,N_4900);
nor U8417 (N_8417,N_5559,N_4006);
and U8418 (N_8418,N_4456,N_4935);
or U8419 (N_8419,N_5692,N_3795);
nand U8420 (N_8420,N_3123,N_4160);
and U8421 (N_8421,N_3289,N_4756);
nor U8422 (N_8422,N_4675,N_5249);
nor U8423 (N_8423,N_5264,N_4682);
or U8424 (N_8424,N_3892,N_4201);
nand U8425 (N_8425,N_3617,N_5139);
or U8426 (N_8426,N_5375,N_4717);
and U8427 (N_8427,N_4314,N_4338);
and U8428 (N_8428,N_5864,N_4288);
and U8429 (N_8429,N_5811,N_5286);
nor U8430 (N_8430,N_4007,N_5594);
nand U8431 (N_8431,N_3697,N_5558);
and U8432 (N_8432,N_5331,N_5775);
nand U8433 (N_8433,N_3440,N_5590);
nor U8434 (N_8434,N_5027,N_4076);
nor U8435 (N_8435,N_5745,N_3450);
and U8436 (N_8436,N_5168,N_4036);
nand U8437 (N_8437,N_3019,N_3719);
nand U8438 (N_8438,N_3980,N_4922);
and U8439 (N_8439,N_4247,N_3540);
nor U8440 (N_8440,N_3639,N_4676);
nor U8441 (N_8441,N_3650,N_3651);
nor U8442 (N_8442,N_5222,N_3606);
and U8443 (N_8443,N_4787,N_5022);
nor U8444 (N_8444,N_4716,N_5108);
or U8445 (N_8445,N_3846,N_3113);
nor U8446 (N_8446,N_5927,N_3470);
or U8447 (N_8447,N_3045,N_5325);
nor U8448 (N_8448,N_4125,N_4781);
nor U8449 (N_8449,N_3339,N_4886);
nand U8450 (N_8450,N_3210,N_5129);
xor U8451 (N_8451,N_4238,N_3523);
or U8452 (N_8452,N_5217,N_4569);
nor U8453 (N_8453,N_4319,N_5682);
and U8454 (N_8454,N_5282,N_4326);
nor U8455 (N_8455,N_3704,N_3412);
xor U8456 (N_8456,N_4580,N_5462);
nor U8457 (N_8457,N_3387,N_5536);
or U8458 (N_8458,N_3682,N_4346);
or U8459 (N_8459,N_3397,N_4956);
or U8460 (N_8460,N_5172,N_3454);
nand U8461 (N_8461,N_4557,N_4418);
nand U8462 (N_8462,N_4256,N_5238);
and U8463 (N_8463,N_5881,N_3787);
nor U8464 (N_8464,N_5305,N_4630);
nand U8465 (N_8465,N_3502,N_5832);
or U8466 (N_8466,N_3122,N_4091);
nor U8467 (N_8467,N_4185,N_3247);
nor U8468 (N_8468,N_4689,N_5301);
nor U8469 (N_8469,N_4739,N_5508);
nor U8470 (N_8470,N_3358,N_4740);
nand U8471 (N_8471,N_5793,N_4253);
nor U8472 (N_8472,N_4430,N_5882);
nor U8473 (N_8473,N_4992,N_5989);
nand U8474 (N_8474,N_4266,N_4383);
and U8475 (N_8475,N_5348,N_5655);
and U8476 (N_8476,N_3155,N_4100);
nor U8477 (N_8477,N_3163,N_4371);
nand U8478 (N_8478,N_4753,N_4972);
or U8479 (N_8479,N_5734,N_4944);
nor U8480 (N_8480,N_3333,N_5383);
nor U8481 (N_8481,N_3850,N_5529);
and U8482 (N_8482,N_3086,N_3931);
nor U8483 (N_8483,N_3528,N_5104);
nor U8484 (N_8484,N_3990,N_4091);
or U8485 (N_8485,N_3642,N_5577);
nor U8486 (N_8486,N_5022,N_4930);
or U8487 (N_8487,N_3913,N_5537);
or U8488 (N_8488,N_5844,N_5801);
nor U8489 (N_8489,N_5657,N_5047);
and U8490 (N_8490,N_4953,N_4248);
or U8491 (N_8491,N_5298,N_5292);
nor U8492 (N_8492,N_3297,N_5403);
and U8493 (N_8493,N_4533,N_3734);
and U8494 (N_8494,N_4909,N_4668);
nand U8495 (N_8495,N_5840,N_3025);
nand U8496 (N_8496,N_5563,N_5218);
nor U8497 (N_8497,N_3245,N_3445);
nor U8498 (N_8498,N_5365,N_5192);
or U8499 (N_8499,N_4351,N_3740);
nor U8500 (N_8500,N_5596,N_4979);
nor U8501 (N_8501,N_5979,N_5281);
or U8502 (N_8502,N_3491,N_4384);
nor U8503 (N_8503,N_4136,N_3369);
or U8504 (N_8504,N_4122,N_4579);
and U8505 (N_8505,N_3573,N_4659);
nand U8506 (N_8506,N_5903,N_3636);
or U8507 (N_8507,N_3401,N_5151);
and U8508 (N_8508,N_3418,N_4752);
and U8509 (N_8509,N_3980,N_4544);
or U8510 (N_8510,N_5858,N_3137);
or U8511 (N_8511,N_4537,N_5993);
nand U8512 (N_8512,N_5529,N_4666);
or U8513 (N_8513,N_5633,N_3968);
or U8514 (N_8514,N_4153,N_5231);
and U8515 (N_8515,N_3336,N_5474);
nor U8516 (N_8516,N_3619,N_4223);
or U8517 (N_8517,N_3244,N_4019);
and U8518 (N_8518,N_5205,N_5337);
or U8519 (N_8519,N_5111,N_5765);
nand U8520 (N_8520,N_4629,N_5621);
or U8521 (N_8521,N_5664,N_3447);
or U8522 (N_8522,N_5494,N_5189);
nor U8523 (N_8523,N_5770,N_5089);
nand U8524 (N_8524,N_4936,N_4565);
nor U8525 (N_8525,N_3391,N_5500);
and U8526 (N_8526,N_3116,N_5205);
or U8527 (N_8527,N_5370,N_5085);
nor U8528 (N_8528,N_3102,N_5781);
nand U8529 (N_8529,N_3437,N_3906);
nand U8530 (N_8530,N_3121,N_5490);
or U8531 (N_8531,N_5823,N_4794);
and U8532 (N_8532,N_4088,N_4167);
nand U8533 (N_8533,N_4520,N_4350);
nand U8534 (N_8534,N_3020,N_4674);
nand U8535 (N_8535,N_3084,N_5868);
nor U8536 (N_8536,N_4330,N_5780);
or U8537 (N_8537,N_4681,N_5608);
or U8538 (N_8538,N_3094,N_5735);
nand U8539 (N_8539,N_4311,N_3824);
or U8540 (N_8540,N_4890,N_5325);
and U8541 (N_8541,N_4202,N_3953);
or U8542 (N_8542,N_4738,N_5894);
xnor U8543 (N_8543,N_3762,N_5933);
or U8544 (N_8544,N_5372,N_3561);
or U8545 (N_8545,N_5502,N_3460);
nand U8546 (N_8546,N_3505,N_4164);
and U8547 (N_8547,N_5117,N_3615);
or U8548 (N_8548,N_5716,N_5568);
nor U8549 (N_8549,N_5154,N_5031);
nor U8550 (N_8550,N_4334,N_4635);
nor U8551 (N_8551,N_4258,N_5019);
or U8552 (N_8552,N_4465,N_4620);
nand U8553 (N_8553,N_3797,N_4842);
nor U8554 (N_8554,N_5676,N_3400);
nand U8555 (N_8555,N_4518,N_3887);
nand U8556 (N_8556,N_5952,N_5188);
nor U8557 (N_8557,N_4616,N_3548);
nor U8558 (N_8558,N_3690,N_5380);
and U8559 (N_8559,N_4192,N_3522);
xor U8560 (N_8560,N_4710,N_4097);
or U8561 (N_8561,N_4812,N_4216);
and U8562 (N_8562,N_4707,N_4068);
or U8563 (N_8563,N_3442,N_3234);
nor U8564 (N_8564,N_4932,N_3089);
and U8565 (N_8565,N_4923,N_5682);
or U8566 (N_8566,N_3586,N_3127);
nand U8567 (N_8567,N_4155,N_5335);
nor U8568 (N_8568,N_3820,N_3323);
or U8569 (N_8569,N_3920,N_4084);
or U8570 (N_8570,N_4088,N_5094);
or U8571 (N_8571,N_5691,N_4348);
or U8572 (N_8572,N_4786,N_5375);
or U8573 (N_8573,N_3019,N_3215);
nor U8574 (N_8574,N_3636,N_4360);
nand U8575 (N_8575,N_5425,N_3874);
nor U8576 (N_8576,N_5032,N_4136);
nor U8577 (N_8577,N_5346,N_5363);
nor U8578 (N_8578,N_5785,N_3561);
nand U8579 (N_8579,N_5885,N_3089);
nand U8580 (N_8580,N_3667,N_5392);
nor U8581 (N_8581,N_3477,N_3132);
or U8582 (N_8582,N_4169,N_3331);
nor U8583 (N_8583,N_5273,N_3214);
nand U8584 (N_8584,N_5482,N_3140);
nand U8585 (N_8585,N_5889,N_3250);
nand U8586 (N_8586,N_5626,N_5532);
and U8587 (N_8587,N_3720,N_4649);
nor U8588 (N_8588,N_5068,N_5436);
nor U8589 (N_8589,N_4685,N_4212);
or U8590 (N_8590,N_5769,N_5823);
nand U8591 (N_8591,N_4159,N_5324);
nand U8592 (N_8592,N_5494,N_5145);
nand U8593 (N_8593,N_4536,N_4001);
nand U8594 (N_8594,N_5676,N_4098);
nand U8595 (N_8595,N_5965,N_4215);
xnor U8596 (N_8596,N_5572,N_3353);
nand U8597 (N_8597,N_3400,N_5200);
or U8598 (N_8598,N_4508,N_4824);
nand U8599 (N_8599,N_5671,N_5034);
nand U8600 (N_8600,N_3358,N_3386);
and U8601 (N_8601,N_5327,N_4190);
and U8602 (N_8602,N_5534,N_3984);
or U8603 (N_8603,N_3855,N_3907);
or U8604 (N_8604,N_4447,N_3303);
nand U8605 (N_8605,N_5265,N_3356);
or U8606 (N_8606,N_3509,N_3857);
or U8607 (N_8607,N_3704,N_4810);
or U8608 (N_8608,N_3935,N_5222);
and U8609 (N_8609,N_3305,N_5499);
or U8610 (N_8610,N_3008,N_4473);
nor U8611 (N_8611,N_4711,N_4265);
nor U8612 (N_8612,N_3529,N_4189);
and U8613 (N_8613,N_5292,N_4719);
or U8614 (N_8614,N_4079,N_5542);
nand U8615 (N_8615,N_3272,N_5345);
or U8616 (N_8616,N_5560,N_4893);
or U8617 (N_8617,N_4818,N_5971);
nor U8618 (N_8618,N_5290,N_4229);
and U8619 (N_8619,N_3578,N_3403);
nand U8620 (N_8620,N_3404,N_5494);
nor U8621 (N_8621,N_4960,N_5027);
or U8622 (N_8622,N_4717,N_5413);
or U8623 (N_8623,N_4853,N_5548);
and U8624 (N_8624,N_3189,N_4358);
or U8625 (N_8625,N_4179,N_3095);
and U8626 (N_8626,N_4035,N_5095);
and U8627 (N_8627,N_5833,N_3729);
nand U8628 (N_8628,N_5057,N_5517);
nand U8629 (N_8629,N_3425,N_3184);
nor U8630 (N_8630,N_4585,N_4183);
and U8631 (N_8631,N_3399,N_3925);
nand U8632 (N_8632,N_3499,N_5980);
or U8633 (N_8633,N_3249,N_5030);
nor U8634 (N_8634,N_4166,N_3182);
and U8635 (N_8635,N_5108,N_3580);
or U8636 (N_8636,N_4195,N_4589);
or U8637 (N_8637,N_4574,N_4904);
or U8638 (N_8638,N_3319,N_4650);
nor U8639 (N_8639,N_5432,N_4302);
and U8640 (N_8640,N_4758,N_5970);
nand U8641 (N_8641,N_5053,N_4257);
or U8642 (N_8642,N_5780,N_4571);
and U8643 (N_8643,N_5288,N_4100);
nor U8644 (N_8644,N_3134,N_4878);
or U8645 (N_8645,N_5408,N_3935);
nand U8646 (N_8646,N_3430,N_4154);
and U8647 (N_8647,N_5108,N_3343);
or U8648 (N_8648,N_5537,N_4194);
and U8649 (N_8649,N_3184,N_5518);
nand U8650 (N_8650,N_3278,N_4863);
and U8651 (N_8651,N_3378,N_5652);
and U8652 (N_8652,N_3136,N_3703);
nor U8653 (N_8653,N_4261,N_3834);
nor U8654 (N_8654,N_5406,N_5137);
or U8655 (N_8655,N_4613,N_3409);
nand U8656 (N_8656,N_3589,N_5569);
and U8657 (N_8657,N_4459,N_5414);
or U8658 (N_8658,N_4193,N_5004);
xor U8659 (N_8659,N_5654,N_5621);
and U8660 (N_8660,N_3971,N_3401);
or U8661 (N_8661,N_5277,N_4027);
and U8662 (N_8662,N_4954,N_3937);
and U8663 (N_8663,N_5491,N_4132);
nand U8664 (N_8664,N_3150,N_4897);
nor U8665 (N_8665,N_5081,N_4103);
nand U8666 (N_8666,N_3260,N_4273);
or U8667 (N_8667,N_4434,N_3252);
xor U8668 (N_8668,N_5365,N_4351);
and U8669 (N_8669,N_3731,N_5346);
and U8670 (N_8670,N_3959,N_5865);
and U8671 (N_8671,N_5324,N_5993);
and U8672 (N_8672,N_4317,N_5751);
nand U8673 (N_8673,N_3886,N_4087);
nor U8674 (N_8674,N_3108,N_5377);
or U8675 (N_8675,N_3720,N_5702);
nor U8676 (N_8676,N_5847,N_3172);
nor U8677 (N_8677,N_3694,N_3510);
nand U8678 (N_8678,N_3285,N_5078);
nand U8679 (N_8679,N_3824,N_3434);
and U8680 (N_8680,N_4090,N_5524);
nand U8681 (N_8681,N_4753,N_5661);
nor U8682 (N_8682,N_5028,N_5409);
and U8683 (N_8683,N_5791,N_3164);
or U8684 (N_8684,N_3820,N_5582);
nor U8685 (N_8685,N_4472,N_5522);
nor U8686 (N_8686,N_3508,N_5050);
nand U8687 (N_8687,N_4615,N_4749);
nor U8688 (N_8688,N_4596,N_5054);
nand U8689 (N_8689,N_5188,N_3385);
or U8690 (N_8690,N_4226,N_4750);
or U8691 (N_8691,N_3589,N_5242);
or U8692 (N_8692,N_5912,N_3528);
nand U8693 (N_8693,N_5836,N_4945);
or U8694 (N_8694,N_5742,N_5631);
nand U8695 (N_8695,N_4474,N_4434);
and U8696 (N_8696,N_3841,N_5788);
and U8697 (N_8697,N_4590,N_3840);
or U8698 (N_8698,N_5541,N_5032);
and U8699 (N_8699,N_5963,N_5045);
or U8700 (N_8700,N_4266,N_5435);
nor U8701 (N_8701,N_3240,N_5306);
nand U8702 (N_8702,N_5513,N_5325);
nor U8703 (N_8703,N_3487,N_3274);
or U8704 (N_8704,N_5839,N_3117);
or U8705 (N_8705,N_3449,N_5361);
or U8706 (N_8706,N_5111,N_5210);
and U8707 (N_8707,N_5531,N_5990);
and U8708 (N_8708,N_5375,N_5753);
or U8709 (N_8709,N_3537,N_3407);
nand U8710 (N_8710,N_5960,N_4860);
xnor U8711 (N_8711,N_4221,N_5190);
nor U8712 (N_8712,N_5629,N_5996);
and U8713 (N_8713,N_3260,N_4107);
nand U8714 (N_8714,N_4711,N_3383);
nor U8715 (N_8715,N_5860,N_3737);
or U8716 (N_8716,N_4573,N_3471);
or U8717 (N_8717,N_3999,N_3621);
and U8718 (N_8718,N_3806,N_3205);
or U8719 (N_8719,N_4859,N_5231);
and U8720 (N_8720,N_5044,N_3377);
nand U8721 (N_8721,N_5838,N_4734);
or U8722 (N_8722,N_3047,N_3528);
nor U8723 (N_8723,N_4961,N_4571);
nand U8724 (N_8724,N_5299,N_4095);
and U8725 (N_8725,N_4516,N_4443);
nand U8726 (N_8726,N_5887,N_5029);
nor U8727 (N_8727,N_3025,N_4219);
nand U8728 (N_8728,N_4773,N_3420);
nand U8729 (N_8729,N_3086,N_3214);
nand U8730 (N_8730,N_4634,N_4922);
or U8731 (N_8731,N_3014,N_3105);
nor U8732 (N_8732,N_5531,N_3170);
and U8733 (N_8733,N_5414,N_3536);
nor U8734 (N_8734,N_4183,N_3595);
nor U8735 (N_8735,N_3003,N_3335);
nor U8736 (N_8736,N_4731,N_3023);
nor U8737 (N_8737,N_5507,N_4963);
nor U8738 (N_8738,N_4681,N_5388);
nor U8739 (N_8739,N_4469,N_5286);
and U8740 (N_8740,N_5349,N_4367);
or U8741 (N_8741,N_5798,N_5728);
nor U8742 (N_8742,N_4985,N_4728);
and U8743 (N_8743,N_5857,N_4641);
nor U8744 (N_8744,N_5551,N_5271);
nor U8745 (N_8745,N_4861,N_4458);
nand U8746 (N_8746,N_5755,N_4692);
or U8747 (N_8747,N_3178,N_4220);
and U8748 (N_8748,N_3042,N_4191);
nor U8749 (N_8749,N_4715,N_4860);
nand U8750 (N_8750,N_5279,N_5932);
nand U8751 (N_8751,N_4011,N_5954);
and U8752 (N_8752,N_4386,N_3378);
nor U8753 (N_8753,N_4893,N_4320);
or U8754 (N_8754,N_5865,N_5006);
nor U8755 (N_8755,N_3311,N_5070);
and U8756 (N_8756,N_4587,N_5795);
or U8757 (N_8757,N_5119,N_5559);
nand U8758 (N_8758,N_3943,N_4929);
nand U8759 (N_8759,N_5924,N_4281);
or U8760 (N_8760,N_3651,N_3222);
nand U8761 (N_8761,N_5479,N_4937);
nand U8762 (N_8762,N_4374,N_4390);
and U8763 (N_8763,N_3157,N_3926);
and U8764 (N_8764,N_3585,N_4953);
nand U8765 (N_8765,N_5721,N_4074);
nor U8766 (N_8766,N_5071,N_3888);
nor U8767 (N_8767,N_5364,N_4499);
nor U8768 (N_8768,N_4018,N_5535);
and U8769 (N_8769,N_3454,N_4698);
nand U8770 (N_8770,N_4474,N_3473);
and U8771 (N_8771,N_4539,N_5243);
and U8772 (N_8772,N_5335,N_4813);
nor U8773 (N_8773,N_4006,N_5148);
or U8774 (N_8774,N_5514,N_5083);
or U8775 (N_8775,N_5489,N_5570);
or U8776 (N_8776,N_4901,N_4988);
or U8777 (N_8777,N_5549,N_5212);
and U8778 (N_8778,N_4056,N_5228);
and U8779 (N_8779,N_5198,N_4066);
or U8780 (N_8780,N_5348,N_4504);
nor U8781 (N_8781,N_4770,N_3119);
or U8782 (N_8782,N_3218,N_3299);
nand U8783 (N_8783,N_4196,N_3424);
nand U8784 (N_8784,N_3692,N_4534);
and U8785 (N_8785,N_4387,N_5207);
nand U8786 (N_8786,N_5758,N_4451);
and U8787 (N_8787,N_4924,N_3268);
or U8788 (N_8788,N_5219,N_5715);
xnor U8789 (N_8789,N_3330,N_3209);
and U8790 (N_8790,N_5545,N_3989);
or U8791 (N_8791,N_3390,N_4721);
nand U8792 (N_8792,N_4030,N_5437);
nand U8793 (N_8793,N_4916,N_4858);
and U8794 (N_8794,N_4839,N_3383);
or U8795 (N_8795,N_3148,N_3360);
and U8796 (N_8796,N_4486,N_4086);
and U8797 (N_8797,N_5818,N_4952);
nand U8798 (N_8798,N_4200,N_3210);
nor U8799 (N_8799,N_5887,N_4029);
nand U8800 (N_8800,N_5555,N_5534);
nand U8801 (N_8801,N_4748,N_4623);
and U8802 (N_8802,N_3025,N_3828);
nor U8803 (N_8803,N_5720,N_3600);
nand U8804 (N_8804,N_3330,N_3076);
and U8805 (N_8805,N_5405,N_5958);
nand U8806 (N_8806,N_5085,N_3517);
or U8807 (N_8807,N_4667,N_5673);
nand U8808 (N_8808,N_4117,N_5259);
nor U8809 (N_8809,N_4715,N_3405);
nand U8810 (N_8810,N_5022,N_3408);
or U8811 (N_8811,N_3364,N_5429);
and U8812 (N_8812,N_4852,N_5804);
or U8813 (N_8813,N_5593,N_5992);
or U8814 (N_8814,N_5248,N_3030);
or U8815 (N_8815,N_3859,N_5994);
and U8816 (N_8816,N_5677,N_5072);
nand U8817 (N_8817,N_3211,N_4622);
and U8818 (N_8818,N_5812,N_5105);
nor U8819 (N_8819,N_3102,N_3830);
or U8820 (N_8820,N_4278,N_3357);
nand U8821 (N_8821,N_3729,N_4271);
or U8822 (N_8822,N_5019,N_5205);
or U8823 (N_8823,N_3804,N_4101);
nand U8824 (N_8824,N_4670,N_3957);
or U8825 (N_8825,N_3958,N_5083);
nand U8826 (N_8826,N_5442,N_4743);
nand U8827 (N_8827,N_4581,N_3799);
nor U8828 (N_8828,N_4176,N_3598);
and U8829 (N_8829,N_5938,N_4766);
nand U8830 (N_8830,N_3379,N_5516);
nand U8831 (N_8831,N_4120,N_3502);
and U8832 (N_8832,N_3850,N_4741);
and U8833 (N_8833,N_5814,N_3642);
nand U8834 (N_8834,N_3752,N_3664);
nor U8835 (N_8835,N_5125,N_3315);
or U8836 (N_8836,N_4000,N_3326);
and U8837 (N_8837,N_3454,N_4233);
nand U8838 (N_8838,N_3976,N_3411);
nand U8839 (N_8839,N_4284,N_4936);
or U8840 (N_8840,N_4938,N_4974);
or U8841 (N_8841,N_3799,N_4998);
or U8842 (N_8842,N_3469,N_4402);
nand U8843 (N_8843,N_5579,N_5127);
and U8844 (N_8844,N_5030,N_5886);
or U8845 (N_8845,N_5605,N_3155);
and U8846 (N_8846,N_5065,N_3086);
nor U8847 (N_8847,N_4841,N_3056);
nand U8848 (N_8848,N_5745,N_5760);
or U8849 (N_8849,N_3140,N_5040);
nor U8850 (N_8850,N_4699,N_5621);
nor U8851 (N_8851,N_5518,N_4468);
nor U8852 (N_8852,N_5894,N_5997);
or U8853 (N_8853,N_4815,N_3811);
nor U8854 (N_8854,N_5455,N_3716);
or U8855 (N_8855,N_3328,N_3354);
nand U8856 (N_8856,N_4636,N_5885);
nand U8857 (N_8857,N_3504,N_4298);
nand U8858 (N_8858,N_3262,N_4557);
or U8859 (N_8859,N_3940,N_4383);
and U8860 (N_8860,N_5896,N_4617);
or U8861 (N_8861,N_4760,N_3118);
nor U8862 (N_8862,N_4555,N_5671);
or U8863 (N_8863,N_4174,N_5889);
nand U8864 (N_8864,N_4481,N_4318);
nand U8865 (N_8865,N_5981,N_3104);
and U8866 (N_8866,N_3516,N_4989);
or U8867 (N_8867,N_4507,N_4491);
nor U8868 (N_8868,N_5376,N_3496);
and U8869 (N_8869,N_3951,N_5845);
nand U8870 (N_8870,N_4970,N_4031);
or U8871 (N_8871,N_4717,N_4239);
nor U8872 (N_8872,N_4119,N_5361);
and U8873 (N_8873,N_3889,N_5244);
nand U8874 (N_8874,N_4553,N_5914);
nand U8875 (N_8875,N_3383,N_5279);
nand U8876 (N_8876,N_4973,N_3236);
nor U8877 (N_8877,N_3654,N_3858);
nand U8878 (N_8878,N_5749,N_3303);
nor U8879 (N_8879,N_3397,N_4922);
nand U8880 (N_8880,N_5031,N_3484);
nor U8881 (N_8881,N_3410,N_5757);
nand U8882 (N_8882,N_4152,N_3251);
nand U8883 (N_8883,N_3379,N_4042);
or U8884 (N_8884,N_4947,N_5179);
nand U8885 (N_8885,N_3255,N_4416);
and U8886 (N_8886,N_4895,N_3416);
nand U8887 (N_8887,N_3769,N_3591);
and U8888 (N_8888,N_5179,N_3546);
and U8889 (N_8889,N_4660,N_3216);
nor U8890 (N_8890,N_4431,N_4230);
and U8891 (N_8891,N_3913,N_5342);
nor U8892 (N_8892,N_3166,N_3886);
nand U8893 (N_8893,N_5944,N_5745);
and U8894 (N_8894,N_5430,N_4894);
nand U8895 (N_8895,N_3464,N_3302);
nor U8896 (N_8896,N_4334,N_3404);
and U8897 (N_8897,N_4804,N_3964);
nor U8898 (N_8898,N_4528,N_5390);
or U8899 (N_8899,N_5441,N_3935);
nor U8900 (N_8900,N_5253,N_3016);
nor U8901 (N_8901,N_5229,N_4238);
nand U8902 (N_8902,N_5617,N_5671);
and U8903 (N_8903,N_4912,N_3303);
or U8904 (N_8904,N_5395,N_4924);
or U8905 (N_8905,N_5622,N_4483);
and U8906 (N_8906,N_4237,N_4056);
nor U8907 (N_8907,N_3704,N_3401);
or U8908 (N_8908,N_4372,N_4384);
or U8909 (N_8909,N_3593,N_5467);
nor U8910 (N_8910,N_5762,N_5965);
and U8911 (N_8911,N_5420,N_5499);
nor U8912 (N_8912,N_5151,N_3504);
xnor U8913 (N_8913,N_5438,N_4763);
nand U8914 (N_8914,N_3500,N_3213);
or U8915 (N_8915,N_3184,N_4024);
nand U8916 (N_8916,N_5927,N_4484);
xnor U8917 (N_8917,N_5416,N_4365);
or U8918 (N_8918,N_3680,N_3808);
nor U8919 (N_8919,N_4845,N_3501);
or U8920 (N_8920,N_4589,N_5859);
nand U8921 (N_8921,N_3674,N_5709);
or U8922 (N_8922,N_3739,N_3677);
and U8923 (N_8923,N_4143,N_3425);
nand U8924 (N_8924,N_4763,N_3051);
or U8925 (N_8925,N_3486,N_5795);
nor U8926 (N_8926,N_3447,N_5342);
or U8927 (N_8927,N_4286,N_5648);
nor U8928 (N_8928,N_4014,N_5813);
nand U8929 (N_8929,N_4019,N_4159);
nand U8930 (N_8930,N_3309,N_4526);
nor U8931 (N_8931,N_4084,N_5891);
and U8932 (N_8932,N_4949,N_5264);
nand U8933 (N_8933,N_5917,N_3437);
or U8934 (N_8934,N_3539,N_3552);
and U8935 (N_8935,N_4884,N_4679);
or U8936 (N_8936,N_5180,N_4462);
nor U8937 (N_8937,N_3924,N_3805);
nor U8938 (N_8938,N_3225,N_4440);
nand U8939 (N_8939,N_4564,N_4444);
nor U8940 (N_8940,N_3527,N_5560);
nor U8941 (N_8941,N_3726,N_4467);
and U8942 (N_8942,N_4330,N_4339);
nand U8943 (N_8943,N_3459,N_5164);
or U8944 (N_8944,N_4245,N_3204);
nand U8945 (N_8945,N_3847,N_4314);
nand U8946 (N_8946,N_5148,N_4100);
nand U8947 (N_8947,N_4257,N_5413);
and U8948 (N_8948,N_4688,N_5578);
nor U8949 (N_8949,N_5551,N_5370);
and U8950 (N_8950,N_4381,N_3705);
and U8951 (N_8951,N_4895,N_5169);
and U8952 (N_8952,N_4287,N_4403);
and U8953 (N_8953,N_3820,N_5407);
nand U8954 (N_8954,N_3988,N_4219);
and U8955 (N_8955,N_4646,N_4399);
or U8956 (N_8956,N_5445,N_4832);
and U8957 (N_8957,N_5758,N_3541);
or U8958 (N_8958,N_3061,N_3089);
nor U8959 (N_8959,N_5473,N_5910);
nand U8960 (N_8960,N_5949,N_4213);
and U8961 (N_8961,N_3524,N_4085);
and U8962 (N_8962,N_5759,N_3963);
nand U8963 (N_8963,N_3131,N_5241);
nor U8964 (N_8964,N_5289,N_3109);
nand U8965 (N_8965,N_5009,N_3778);
or U8966 (N_8966,N_3702,N_4869);
or U8967 (N_8967,N_3619,N_5956);
nor U8968 (N_8968,N_4068,N_4476);
and U8969 (N_8969,N_5821,N_5687);
or U8970 (N_8970,N_3178,N_3493);
nor U8971 (N_8971,N_5537,N_5692);
or U8972 (N_8972,N_4359,N_5550);
and U8973 (N_8973,N_4719,N_4021);
and U8974 (N_8974,N_4505,N_5765);
or U8975 (N_8975,N_4148,N_5666);
nor U8976 (N_8976,N_5392,N_4147);
or U8977 (N_8977,N_4568,N_3755);
nor U8978 (N_8978,N_5518,N_3280);
and U8979 (N_8979,N_5040,N_5064);
and U8980 (N_8980,N_5905,N_3561);
or U8981 (N_8981,N_3663,N_3313);
or U8982 (N_8982,N_5823,N_5106);
and U8983 (N_8983,N_5160,N_5659);
nand U8984 (N_8984,N_5522,N_3793);
or U8985 (N_8985,N_5848,N_5915);
or U8986 (N_8986,N_5505,N_4472);
nor U8987 (N_8987,N_4353,N_3091);
or U8988 (N_8988,N_4438,N_4495);
nand U8989 (N_8989,N_4286,N_5577);
nor U8990 (N_8990,N_4862,N_4574);
nand U8991 (N_8991,N_3668,N_3191);
or U8992 (N_8992,N_5200,N_5664);
or U8993 (N_8993,N_4733,N_5236);
nand U8994 (N_8994,N_5439,N_3737);
and U8995 (N_8995,N_5266,N_3499);
or U8996 (N_8996,N_3369,N_4268);
or U8997 (N_8997,N_3185,N_4243);
nand U8998 (N_8998,N_5386,N_4259);
xnor U8999 (N_8999,N_3015,N_5334);
nor U9000 (N_9000,N_7529,N_8473);
or U9001 (N_9001,N_7225,N_8435);
or U9002 (N_9002,N_7152,N_6656);
nand U9003 (N_9003,N_6214,N_7884);
nor U9004 (N_9004,N_6154,N_6477);
nand U9005 (N_9005,N_7218,N_6377);
or U9006 (N_9006,N_8373,N_7396);
and U9007 (N_9007,N_8086,N_7927);
nor U9008 (N_9008,N_8127,N_8080);
and U9009 (N_9009,N_6961,N_8837);
nand U9010 (N_9010,N_6193,N_6676);
or U9011 (N_9011,N_7999,N_7942);
and U9012 (N_9012,N_6055,N_8941);
nor U9013 (N_9013,N_7405,N_8747);
xnor U9014 (N_9014,N_6626,N_7374);
and U9015 (N_9015,N_8582,N_6038);
nor U9016 (N_9016,N_8072,N_6456);
nand U9017 (N_9017,N_6772,N_7462);
nand U9018 (N_9018,N_6727,N_6830);
or U9019 (N_9019,N_7475,N_7861);
or U9020 (N_9020,N_8372,N_8122);
and U9021 (N_9021,N_7757,N_8391);
or U9022 (N_9022,N_7793,N_8480);
and U9023 (N_9023,N_6853,N_7386);
nor U9024 (N_9024,N_8370,N_8802);
or U9025 (N_9025,N_7070,N_6339);
and U9026 (N_9026,N_6723,N_7361);
nand U9027 (N_9027,N_8056,N_6966);
nor U9028 (N_9028,N_8882,N_6500);
and U9029 (N_9029,N_6840,N_8828);
and U9030 (N_9030,N_7502,N_7780);
nor U9031 (N_9031,N_7878,N_8617);
nand U9032 (N_9032,N_7691,N_6642);
and U9033 (N_9033,N_7432,N_8458);
and U9034 (N_9034,N_7764,N_8919);
nand U9035 (N_9035,N_6632,N_7178);
or U9036 (N_9036,N_7843,N_6705);
nand U9037 (N_9037,N_6645,N_6893);
nand U9038 (N_9038,N_7029,N_7687);
xnor U9039 (N_9039,N_8599,N_8134);
xnor U9040 (N_9040,N_6802,N_6597);
nand U9041 (N_9041,N_6509,N_8417);
and U9042 (N_9042,N_6075,N_7379);
nor U9043 (N_9043,N_7819,N_6322);
and U9044 (N_9044,N_8764,N_6534);
or U9045 (N_9045,N_8931,N_6871);
nor U9046 (N_9046,N_6265,N_7748);
nand U9047 (N_9047,N_6163,N_8379);
and U9048 (N_9048,N_8783,N_8507);
nor U9049 (N_9049,N_8223,N_8785);
xnor U9050 (N_9050,N_8441,N_8903);
nor U9051 (N_9051,N_6362,N_6153);
nor U9052 (N_9052,N_7875,N_6269);
nand U9053 (N_9053,N_6810,N_7114);
and U9054 (N_9054,N_7438,N_8389);
nand U9055 (N_9055,N_8008,N_7362);
nand U9056 (N_9056,N_7447,N_8991);
or U9057 (N_9057,N_6122,N_8574);
or U9058 (N_9058,N_6764,N_8346);
nor U9059 (N_9059,N_7812,N_7328);
or U9060 (N_9060,N_6282,N_6601);
xnor U9061 (N_9061,N_7320,N_6683);
nand U9062 (N_9062,N_6140,N_6858);
and U9063 (N_9063,N_8815,N_8488);
nor U9064 (N_9064,N_8087,N_7209);
nand U9065 (N_9065,N_7799,N_8098);
nand U9066 (N_9066,N_8451,N_7571);
nor U9067 (N_9067,N_7236,N_6677);
and U9068 (N_9068,N_8757,N_8039);
nor U9069 (N_9069,N_7129,N_6901);
and U9070 (N_9070,N_7674,N_8581);
nand U9071 (N_9071,N_6717,N_7005);
or U9072 (N_9072,N_6742,N_8557);
xnor U9073 (N_9073,N_6932,N_8492);
nor U9074 (N_9074,N_6868,N_6841);
and U9075 (N_9075,N_7421,N_6510);
nor U9076 (N_9076,N_8609,N_6039);
and U9077 (N_9077,N_8795,N_6883);
and U9078 (N_9078,N_8212,N_8779);
and U9079 (N_9079,N_7511,N_6844);
and U9080 (N_9080,N_7338,N_6398);
nand U9081 (N_9081,N_8155,N_6958);
nand U9082 (N_9082,N_8014,N_7709);
and U9083 (N_9083,N_8528,N_7869);
nand U9084 (N_9084,N_7557,N_8425);
nor U9085 (N_9085,N_8844,N_6741);
nor U9086 (N_9086,N_7915,N_6201);
or U9087 (N_9087,N_6620,N_7616);
or U9088 (N_9088,N_6365,N_8199);
or U9089 (N_9089,N_7954,N_7656);
nand U9090 (N_9090,N_8894,N_6962);
nor U9091 (N_9091,N_7763,N_7901);
nand U9092 (N_9092,N_7606,N_7015);
and U9093 (N_9093,N_7309,N_6314);
nor U9094 (N_9094,N_7060,N_6704);
or U9095 (N_9095,N_6419,N_6141);
nor U9096 (N_9096,N_6526,N_7082);
and U9097 (N_9097,N_6939,N_7118);
and U9098 (N_9098,N_6591,N_6297);
nand U9099 (N_9099,N_8428,N_6785);
nand U9100 (N_9100,N_6286,N_8638);
nand U9101 (N_9101,N_8934,N_6607);
or U9102 (N_9102,N_7052,N_6112);
nor U9103 (N_9103,N_7248,N_7985);
and U9104 (N_9104,N_6831,N_8999);
nand U9105 (N_9105,N_7559,N_8801);
nor U9106 (N_9106,N_8926,N_7816);
or U9107 (N_9107,N_6832,N_7916);
or U9108 (N_9108,N_7684,N_6264);
and U9109 (N_9109,N_6346,N_8368);
or U9110 (N_9110,N_6430,N_7223);
nor U9111 (N_9111,N_6519,N_6133);
nor U9112 (N_9112,N_7403,N_6564);
nand U9113 (N_9113,N_8251,N_6424);
nor U9114 (N_9114,N_7750,N_8610);
and U9115 (N_9115,N_6266,N_6529);
nand U9116 (N_9116,N_8491,N_8294);
and U9117 (N_9117,N_8682,N_7470);
and U9118 (N_9118,N_6261,N_8347);
nor U9119 (N_9119,N_6064,N_7651);
nand U9120 (N_9120,N_6442,N_6945);
or U9121 (N_9121,N_8085,N_7220);
nand U9122 (N_9122,N_8915,N_7893);
or U9123 (N_9123,N_6439,N_8065);
xnor U9124 (N_9124,N_6572,N_6826);
and U9125 (N_9125,N_6040,N_7690);
or U9126 (N_9126,N_8258,N_8032);
nor U9127 (N_9127,N_8579,N_7887);
nor U9128 (N_9128,N_7425,N_7117);
nand U9129 (N_9129,N_6916,N_8414);
or U9130 (N_9130,N_7296,N_7215);
nand U9131 (N_9131,N_6944,N_6513);
nor U9132 (N_9132,N_7020,N_7105);
nand U9133 (N_9133,N_6602,N_7413);
nor U9134 (N_9134,N_6931,N_8268);
or U9135 (N_9135,N_7713,N_7370);
nor U9136 (N_9136,N_6582,N_6910);
nand U9137 (N_9137,N_8314,N_6919);
or U9138 (N_9138,N_6808,N_8699);
and U9139 (N_9139,N_8850,N_6964);
nand U9140 (N_9140,N_8386,N_7357);
xnor U9141 (N_9141,N_6045,N_6225);
or U9142 (N_9142,N_7930,N_6665);
nand U9143 (N_9143,N_6775,N_7935);
xnor U9144 (N_9144,N_8967,N_8929);
and U9145 (N_9145,N_7372,N_8271);
nor U9146 (N_9146,N_6761,N_8656);
nand U9147 (N_9147,N_7563,N_7364);
nor U9148 (N_9148,N_7092,N_8021);
nand U9149 (N_9149,N_7091,N_6807);
and U9150 (N_9150,N_6878,N_8880);
nand U9151 (N_9151,N_8918,N_7132);
nor U9152 (N_9152,N_6949,N_6943);
nor U9153 (N_9153,N_7094,N_8295);
nor U9154 (N_9154,N_7592,N_7756);
nor U9155 (N_9155,N_7172,N_7187);
nor U9156 (N_9156,N_8732,N_8781);
nand U9157 (N_9157,N_8627,N_8355);
nand U9158 (N_9158,N_6343,N_7961);
nor U9159 (N_9159,N_7801,N_6037);
nand U9160 (N_9160,N_6071,N_6034);
and U9161 (N_9161,N_8010,N_6559);
nand U9162 (N_9162,N_7791,N_6104);
and U9163 (N_9163,N_8674,N_8826);
nand U9164 (N_9164,N_7399,N_7337);
or U9165 (N_9165,N_8614,N_8561);
nand U9166 (N_9166,N_6938,N_7246);
or U9167 (N_9167,N_7648,N_7978);
nand U9168 (N_9168,N_6863,N_8711);
or U9169 (N_9169,N_7727,N_8529);
nor U9170 (N_9170,N_8165,N_6847);
and U9171 (N_9171,N_7979,N_6445);
nor U9172 (N_9172,N_7813,N_7620);
or U9173 (N_9173,N_7834,N_6864);
nor U9174 (N_9174,N_6058,N_7739);
or U9175 (N_9175,N_8825,N_6546);
or U9176 (N_9176,N_7782,N_7702);
and U9177 (N_9177,N_8168,N_7213);
and U9178 (N_9178,N_6794,N_6881);
and U9179 (N_9179,N_8615,N_8835);
nand U9180 (N_9180,N_7027,N_7058);
and U9181 (N_9181,N_8910,N_7423);
nor U9182 (N_9182,N_8486,N_7235);
xnor U9183 (N_9183,N_6896,N_7474);
or U9184 (N_9184,N_8806,N_6630);
nor U9185 (N_9185,N_6765,N_7800);
xnor U9186 (N_9186,N_8863,N_7877);
nor U9187 (N_9187,N_6169,N_6205);
nor U9188 (N_9188,N_7641,N_7351);
and U9189 (N_9189,N_8658,N_8317);
nand U9190 (N_9190,N_8696,N_6256);
or U9191 (N_9191,N_6004,N_6053);
nor U9192 (N_9192,N_6084,N_6707);
nor U9193 (N_9193,N_6484,N_6953);
and U9194 (N_9194,N_8680,N_6797);
or U9195 (N_9195,N_7039,N_8104);
nor U9196 (N_9196,N_6756,N_6976);
nor U9197 (N_9197,N_7322,N_6616);
nand U9198 (N_9198,N_7963,N_7941);
nand U9199 (N_9199,N_6784,N_8157);
or U9200 (N_9200,N_6651,N_8832);
nand U9201 (N_9201,N_8675,N_7504);
nand U9202 (N_9202,N_6793,N_8431);
nand U9203 (N_9203,N_7818,N_6215);
nand U9204 (N_9204,N_7456,N_6493);
xnor U9205 (N_9205,N_8963,N_6006);
and U9206 (N_9206,N_7131,N_8467);
and U9207 (N_9207,N_7140,N_6253);
nor U9208 (N_9208,N_7440,N_8814);
nand U9209 (N_9209,N_6934,N_7057);
nor U9210 (N_9210,N_7341,N_7852);
or U9211 (N_9211,N_8131,N_8113);
nor U9212 (N_9212,N_7081,N_8149);
nor U9213 (N_9213,N_8395,N_7449);
nand U9214 (N_9214,N_8276,N_7241);
and U9215 (N_9215,N_7909,N_8809);
nand U9216 (N_9216,N_7632,N_8429);
nor U9217 (N_9217,N_7195,N_7479);
nand U9218 (N_9218,N_6933,N_8184);
and U9219 (N_9219,N_7442,N_8810);
nand U9220 (N_9220,N_7969,N_6388);
and U9221 (N_9221,N_6702,N_8728);
nor U9222 (N_9222,N_7417,N_6092);
nand U9223 (N_9223,N_6277,N_6965);
or U9224 (N_9224,N_8642,N_7749);
and U9225 (N_9225,N_7698,N_7252);
and U9226 (N_9226,N_7743,N_6172);
and U9227 (N_9227,N_7074,N_7535);
nor U9228 (N_9228,N_6638,N_8378);
or U9229 (N_9229,N_6619,N_6081);
nand U9230 (N_9230,N_7448,N_7306);
and U9231 (N_9231,N_8590,N_8793);
nand U9232 (N_9232,N_8816,N_8437);
and U9233 (N_9233,N_7811,N_6778);
and U9234 (N_9234,N_8201,N_8464);
and U9235 (N_9235,N_6560,N_8092);
nand U9236 (N_9236,N_7980,N_7075);
and U9237 (N_9237,N_7469,N_7704);
and U9238 (N_9238,N_8676,N_8463);
or U9239 (N_9239,N_8444,N_8876);
nor U9240 (N_9240,N_8019,N_8266);
and U9241 (N_9241,N_6166,N_8140);
xnor U9242 (N_9242,N_6539,N_6235);
nor U9243 (N_9243,N_6022,N_8583);
or U9244 (N_9244,N_8371,N_7804);
nand U9245 (N_9245,N_6593,N_6188);
or U9246 (N_9246,N_7624,N_8945);
and U9247 (N_9247,N_8545,N_8499);
or U9248 (N_9248,N_8057,N_8254);
or U9249 (N_9249,N_7407,N_8426);
and U9250 (N_9250,N_8135,N_6655);
nor U9251 (N_9251,N_6036,N_8780);
nand U9252 (N_9252,N_6250,N_6305);
nor U9253 (N_9253,N_8954,N_7612);
xnor U9254 (N_9254,N_8883,N_7412);
xnor U9255 (N_9255,N_8800,N_7711);
nor U9256 (N_9256,N_8232,N_6108);
or U9257 (N_9257,N_6384,N_7028);
and U9258 (N_9258,N_7607,N_7790);
nor U9259 (N_9259,N_8247,N_7881);
and U9260 (N_9260,N_8027,N_6811);
and U9261 (N_9261,N_6984,N_6818);
and U9262 (N_9262,N_8689,N_7001);
nor U9263 (N_9263,N_6900,N_8687);
or U9264 (N_9264,N_8331,N_7794);
and U9265 (N_9265,N_6094,N_7024);
nor U9266 (N_9266,N_7299,N_8377);
or U9267 (N_9267,N_8046,N_6506);
nor U9268 (N_9268,N_6165,N_7805);
nand U9269 (N_9269,N_6985,N_8836);
or U9270 (N_9270,N_6162,N_8269);
xnor U9271 (N_9271,N_8543,N_8079);
nor U9272 (N_9272,N_7113,N_8237);
nor U9273 (N_9273,N_8474,N_7597);
nand U9274 (N_9274,N_6341,N_6993);
nand U9275 (N_9275,N_8603,N_6392);
nand U9276 (N_9276,N_6413,N_8907);
or U9277 (N_9277,N_6508,N_7331);
nor U9278 (N_9278,N_8120,N_7012);
and U9279 (N_9279,N_7609,N_6798);
and U9280 (N_9280,N_8572,N_8526);
nand U9281 (N_9281,N_7018,N_6043);
nand U9282 (N_9282,N_8913,N_6790);
nor U9283 (N_9283,N_7016,N_8875);
nand U9284 (N_9284,N_6570,N_8281);
nor U9285 (N_9285,N_8629,N_8105);
or U9286 (N_9286,N_6464,N_7411);
nand U9287 (N_9287,N_7725,N_6070);
and U9288 (N_9288,N_8013,N_7135);
or U9289 (N_9289,N_6998,N_8985);
nand U9290 (N_9290,N_7089,N_6003);
or U9291 (N_9291,N_7821,N_7147);
or U9292 (N_9292,N_7768,N_7766);
and U9293 (N_9293,N_7079,N_8082);
nor U9294 (N_9294,N_7486,N_8948);
and U9295 (N_9295,N_6994,N_6258);
and U9296 (N_9296,N_8402,N_6940);
nand U9297 (N_9297,N_7579,N_7705);
or U9298 (N_9298,N_7912,N_8471);
and U9299 (N_9299,N_7009,N_7325);
and U9300 (N_9300,N_7731,N_6098);
nor U9301 (N_9301,N_7002,N_8578);
or U9302 (N_9302,N_6694,N_6604);
and U9303 (N_9303,N_7150,N_7314);
or U9304 (N_9304,N_7019,N_7829);
and U9305 (N_9305,N_6817,N_7463);
nor U9306 (N_9306,N_8969,N_7675);
nor U9307 (N_9307,N_8960,N_7459);
nand U9308 (N_9308,N_7678,N_7703);
or U9309 (N_9309,N_7226,N_8797);
xnor U9310 (N_9310,N_6614,N_7233);
and U9311 (N_9311,N_7644,N_6995);
or U9312 (N_9312,N_7830,N_7575);
and U9313 (N_9313,N_6360,N_7342);
nor U9314 (N_9314,N_8712,N_6639);
nor U9315 (N_9315,N_6241,N_8344);
nor U9316 (N_9316,N_8196,N_6990);
nand U9317 (N_9317,N_6449,N_7655);
nor U9318 (N_9318,N_6581,N_6495);
or U9319 (N_9319,N_6792,N_7721);
and U9320 (N_9320,N_7733,N_6576);
and U9321 (N_9321,N_6552,N_7334);
nor U9322 (N_9322,N_8808,N_6516);
and U9323 (N_9323,N_7401,N_6307);
and U9324 (N_9324,N_7769,N_6009);
and U9325 (N_9325,N_6000,N_8398);
and U9326 (N_9326,N_7481,N_6118);
nand U9327 (N_9327,N_6720,N_8255);
and U9328 (N_9328,N_6059,N_6414);
and U9329 (N_9329,N_6119,N_7171);
xnor U9330 (N_9330,N_6819,N_7292);
or U9331 (N_9331,N_8576,N_8984);
and U9332 (N_9332,N_8477,N_6553);
nor U9333 (N_9333,N_7290,N_6967);
nor U9334 (N_9334,N_8513,N_6050);
and U9335 (N_9335,N_8319,N_7997);
nand U9336 (N_9336,N_6236,N_6278);
and U9337 (N_9337,N_8619,N_6611);
and U9338 (N_9338,N_8933,N_7103);
nand U9339 (N_9339,N_7210,N_6887);
and U9340 (N_9340,N_8261,N_7169);
nand U9341 (N_9341,N_8300,N_6773);
nand U9342 (N_9342,N_8866,N_7426);
and U9343 (N_9343,N_6244,N_7489);
nor U9344 (N_9344,N_6578,N_7416);
nor U9345 (N_9345,N_7377,N_6117);
nand U9346 (N_9346,N_7717,N_8900);
or U9347 (N_9347,N_7158,N_8874);
and U9348 (N_9348,N_8328,N_7659);
and U9349 (N_9349,N_8307,N_7906);
and U9350 (N_9350,N_8996,N_7163);
nor U9351 (N_9351,N_7496,N_7628);
nand U9352 (N_9352,N_7765,N_7880);
nand U9353 (N_9353,N_7670,N_7669);
or U9354 (N_9354,N_7585,N_7049);
or U9355 (N_9355,N_6661,N_6476);
xnor U9356 (N_9356,N_8760,N_7633);
nor U9357 (N_9357,N_6641,N_8720);
or U9358 (N_9358,N_8460,N_7550);
or U9359 (N_9359,N_7100,N_6726);
or U9360 (N_9360,N_8438,N_6606);
and U9361 (N_9361,N_8365,N_7787);
and U9362 (N_9362,N_8198,N_6185);
nor U9363 (N_9363,N_6721,N_8045);
nand U9364 (N_9364,N_6218,N_6575);
or U9365 (N_9365,N_6311,N_6213);
or U9366 (N_9366,N_6359,N_7435);
nor U9367 (N_9367,N_6946,N_6538);
nor U9368 (N_9368,N_6254,N_6409);
nor U9369 (N_9369,N_6458,N_7917);
nand U9370 (N_9370,N_8858,N_8842);
or U9371 (N_9371,N_7323,N_6753);
nor U9372 (N_9372,N_7257,N_6835);
or U9373 (N_9373,N_8535,N_7216);
nor U9374 (N_9374,N_7123,N_8770);
and U9375 (N_9375,N_7570,N_6845);
nand U9376 (N_9376,N_7728,N_7182);
or U9377 (N_9377,N_7510,N_8719);
and U9378 (N_9378,N_8708,N_8174);
xor U9379 (N_9379,N_8539,N_7419);
nor U9380 (N_9380,N_7820,N_8182);
nand U9381 (N_9381,N_7006,N_8299);
or U9382 (N_9382,N_6347,N_6627);
nor U9383 (N_9383,N_8077,N_8742);
and U9384 (N_9384,N_8384,N_7817);
nor U9385 (N_9385,N_8245,N_8259);
nand U9386 (N_9386,N_6324,N_8573);
or U9387 (N_9387,N_7537,N_6354);
nor U9388 (N_9388,N_6417,N_6759);
and U9389 (N_9389,N_8052,N_6787);
and U9390 (N_9390,N_7940,N_8738);
nand U9391 (N_9391,N_7198,N_6147);
nand U9392 (N_9392,N_8509,N_7958);
or U9393 (N_9393,N_8267,N_7896);
nand U9394 (N_9394,N_7789,N_6345);
nor U9395 (N_9395,N_8519,N_8979);
or U9396 (N_9396,N_7760,N_7128);
nand U9397 (N_9397,N_7211,N_6448);
nand U9398 (N_9398,N_6997,N_6594);
and U9399 (N_9399,N_8493,N_8531);
nand U9400 (N_9400,N_6757,N_8498);
nand U9401 (N_9401,N_8361,N_7924);
nand U9402 (N_9402,N_7138,N_7546);
nor U9403 (N_9403,N_6545,N_6482);
nor U9404 (N_9404,N_6740,N_8073);
nor U9405 (N_9405,N_6471,N_7175);
or U9406 (N_9406,N_8089,N_8733);
nand U9407 (N_9407,N_6535,N_7243);
nor U9408 (N_9408,N_8798,N_7951);
or U9409 (N_9409,N_7176,N_6437);
xor U9410 (N_9410,N_8541,N_7736);
nor U9411 (N_9411,N_8530,N_6536);
nand U9412 (N_9412,N_6067,N_6820);
or U9413 (N_9413,N_7533,N_6541);
nand U9414 (N_9414,N_6565,N_7304);
and U9415 (N_9415,N_7627,N_6828);
and U9416 (N_9416,N_7706,N_7737);
and U9417 (N_9417,N_7840,N_7160);
nand U9418 (N_9418,N_6116,N_6065);
or U9419 (N_9419,N_6743,N_6429);
and U9420 (N_9420,N_7751,N_8242);
or U9421 (N_9421,N_6202,N_7471);
or U9422 (N_9422,N_6222,N_8616);
nand U9423 (N_9423,N_8195,N_6629);
or U9424 (N_9424,N_7116,N_8621);
and U9425 (N_9425,N_8006,N_8909);
nor U9426 (N_9426,N_7038,N_7807);
or U9427 (N_9427,N_8011,N_6547);
and U9428 (N_9428,N_6352,N_6275);
nor U9429 (N_9429,N_6838,N_7430);
and U9430 (N_9430,N_7998,N_8515);
and U9431 (N_9431,N_6770,N_7988);
nor U9432 (N_9432,N_8840,N_6668);
and U9433 (N_9433,N_6355,N_7914);
and U9434 (N_9434,N_8562,N_7034);
nand U9435 (N_9435,N_8505,N_8412);
and U9436 (N_9436,N_7615,N_8446);
nand U9437 (N_9437,N_7047,N_6701);
and U9438 (N_9438,N_7302,N_7104);
and U9439 (N_9439,N_7063,N_8688);
and U9440 (N_9440,N_8326,N_6300);
nor U9441 (N_9441,N_6888,N_8016);
nand U9442 (N_9442,N_6806,N_8522);
or U9443 (N_9443,N_7156,N_7983);
and U9444 (N_9444,N_6762,N_7347);
nor U9445 (N_9445,N_6309,N_8246);
nor U9446 (N_9446,N_6031,N_7545);
nor U9447 (N_9447,N_8596,N_6530);
and U9448 (N_9448,N_7427,N_7686);
nor U9449 (N_9449,N_7359,N_6557);
or U9450 (N_9450,N_6867,N_7000);
and U9451 (N_9451,N_7457,N_6121);
or U9452 (N_9452,N_7010,N_7910);
nor U9453 (N_9453,N_8956,N_6408);
and U9454 (N_9454,N_7206,N_6462);
nor U9455 (N_9455,N_8406,N_8569);
nor U9456 (N_9456,N_7352,N_7576);
or U9457 (N_9457,N_8323,N_8443);
nand U9458 (N_9458,N_8898,N_7936);
and U9459 (N_9459,N_6461,N_6865);
nand U9460 (N_9460,N_7385,N_6816);
nand U9461 (N_9461,N_6503,N_7521);
and U9462 (N_9462,N_7167,N_8896);
or U9463 (N_9463,N_6164,N_8214);
or U9464 (N_9464,N_6969,N_7255);
and U9465 (N_9465,N_8668,N_8304);
and U9466 (N_9466,N_7693,N_6693);
and U9467 (N_9467,N_7273,N_6986);
nor U9468 (N_9468,N_8097,N_7295);
nor U9469 (N_9469,N_7078,N_7431);
and U9470 (N_9470,N_8623,N_6674);
or U9471 (N_9471,N_7358,N_8309);
nor U9472 (N_9472,N_7069,N_8986);
nor U9473 (N_9473,N_7467,N_6284);
nor U9474 (N_9474,N_8823,N_7055);
nor U9475 (N_9475,N_6518,N_6160);
or U9476 (N_9476,N_7491,N_8924);
nand U9477 (N_9477,N_7845,N_8141);
nand U9478 (N_9478,N_6737,N_6542);
and U9479 (N_9479,N_7168,N_7313);
or U9480 (N_9480,N_7697,N_6399);
or U9481 (N_9481,N_8670,N_6569);
or U9482 (N_9482,N_8947,N_7544);
or U9483 (N_9483,N_7099,N_7494);
and U9484 (N_9484,N_6167,N_8961);
nor U9485 (N_9485,N_6033,N_7738);
nor U9486 (N_9486,N_7524,N_7646);
or U9487 (N_9487,N_7761,N_8125);
or U9488 (N_9488,N_6191,N_8618);
nand U9489 (N_9489,N_7250,N_8396);
nor U9490 (N_9490,N_6574,N_6544);
or U9491 (N_9491,N_6151,N_8554);
nor U9492 (N_9492,N_7393,N_6517);
or U9493 (N_9493,N_6907,N_8265);
nor U9494 (N_9494,N_7658,N_6886);
and U9495 (N_9495,N_6469,N_6978);
nand U9496 (N_9496,N_6443,N_7932);
nor U9497 (N_9497,N_6975,N_8475);
nand U9498 (N_9498,N_8558,N_6259);
nand U9499 (N_9499,N_8054,N_8920);
nor U9500 (N_9500,N_7891,N_7841);
and U9501 (N_9501,N_8495,N_7536);
and U9502 (N_9502,N_7554,N_7872);
or U9503 (N_9503,N_7836,N_6103);
or U9504 (N_9504,N_8594,N_8830);
and U9505 (N_9505,N_7781,N_7716);
nor U9506 (N_9506,N_8308,N_7271);
and U9507 (N_9507,N_7453,N_7622);
and U9508 (N_9508,N_7476,N_7946);
nor U9509 (N_9509,N_6069,N_6852);
or U9510 (N_9510,N_8788,N_6531);
nor U9511 (N_9511,N_6217,N_8704);
xor U9512 (N_9512,N_6970,N_7788);
and U9513 (N_9513,N_7133,N_8262);
or U9514 (N_9514,N_6130,N_7797);
and U9515 (N_9515,N_6453,N_6230);
and U9516 (N_9516,N_7565,N_7185);
nand U9517 (N_9517,N_6180,N_7108);
or U9518 (N_9518,N_7610,N_6991);
or U9519 (N_9519,N_7353,N_6690);
xnor U9520 (N_9520,N_6955,N_8363);
or U9521 (N_9521,N_6874,N_7972);
nor U9522 (N_9522,N_8807,N_8752);
nor U9523 (N_9523,N_6268,N_6459);
or U9524 (N_9524,N_8278,N_6466);
nor U9525 (N_9525,N_6042,N_7631);
and U9526 (N_9526,N_6950,N_7558);
and U9527 (N_9527,N_8138,N_6633);
nor U9528 (N_9528,N_7525,N_6488);
and U9529 (N_9529,N_6338,N_6941);
or U9530 (N_9530,N_7943,N_8970);
and U9531 (N_9531,N_8508,N_8822);
or U9532 (N_9532,N_6631,N_7465);
nand U9533 (N_9533,N_8588,N_8358);
nand U9534 (N_9534,N_6851,N_6357);
and U9535 (N_9535,N_8133,N_6537);
nor U9536 (N_9536,N_8418,N_8673);
nor U9537 (N_9537,N_7986,N_7722);
nor U9538 (N_9538,N_6187,N_8018);
and U9539 (N_9539,N_6082,N_6463);
or U9540 (N_9540,N_8163,N_7137);
nor U9541 (N_9541,N_8356,N_6479);
and U9542 (N_9542,N_8655,N_7040);
or U9543 (N_9543,N_6358,N_8827);
or U9544 (N_9544,N_7149,N_8185);
nor U9545 (N_9545,N_7339,N_8383);
nand U9546 (N_9546,N_6722,N_6769);
or U9547 (N_9547,N_6326,N_8877);
nand U9548 (N_9548,N_6821,N_7520);
and U9549 (N_9549,N_6873,N_6760);
nand U9550 (N_9550,N_6292,N_6567);
and U9551 (N_9551,N_8124,N_6788);
and U9552 (N_9552,N_6018,N_6540);
and U9553 (N_9553,N_7517,N_7966);
nor U9554 (N_9554,N_8660,N_7231);
and U9555 (N_9555,N_7957,N_6029);
nand U9556 (N_9556,N_8812,N_6293);
and U9557 (N_9557,N_8677,N_7270);
nor U9558 (N_9558,N_8553,N_8648);
nor U9559 (N_9559,N_8683,N_7383);
nand U9560 (N_9560,N_8620,N_8713);
nand U9561 (N_9561,N_7317,N_6410);
nand U9562 (N_9562,N_7251,N_6138);
nor U9563 (N_9563,N_7224,N_8602);
nand U9564 (N_9564,N_6299,N_8496);
or U9565 (N_9565,N_8524,N_7191);
nor U9566 (N_9566,N_7086,N_8290);
or U9567 (N_9567,N_8362,N_6183);
xor U9568 (N_9568,N_7598,N_7180);
and U9569 (N_9569,N_7398,N_8661);
nor U9570 (N_9570,N_6749,N_6751);
and U9571 (N_9571,N_8928,N_8550);
nor U9572 (N_9572,N_7586,N_7652);
or U9573 (N_9573,N_6767,N_7037);
nor U9574 (N_9574,N_6472,N_6132);
nand U9575 (N_9575,N_6603,N_6703);
and U9576 (N_9576,N_6260,N_7350);
and U9577 (N_9577,N_8717,N_6666);
nor U9578 (N_9578,N_7025,N_7919);
or U9579 (N_9579,N_6366,N_8763);
nor U9580 (N_9580,N_6189,N_7327);
or U9581 (N_9581,N_8436,N_7204);
and U9582 (N_9582,N_8721,N_6905);
or U9583 (N_9583,N_6407,N_6455);
nand U9584 (N_9584,N_6379,N_7959);
nor U9585 (N_9585,N_6989,N_7838);
nor U9586 (N_9586,N_7124,N_6273);
or U9587 (N_9587,N_8108,N_8702);
and U9588 (N_9588,N_7949,N_7505);
or U9589 (N_9589,N_6446,N_7835);
or U9590 (N_9590,N_7614,N_6061);
and U9591 (N_9591,N_7567,N_7267);
or U9592 (N_9592,N_8459,N_8927);
nor U9593 (N_9593,N_8939,N_8889);
and U9594 (N_9594,N_6709,N_8536);
or U9595 (N_9595,N_6897,N_8186);
or U9596 (N_9596,N_6605,N_7183);
nand U9597 (N_9597,N_8975,N_8280);
or U9598 (N_9598,N_7572,N_8637);
nand U9599 (N_9599,N_7240,N_6382);
xor U9600 (N_9600,N_7621,N_6023);
or U9601 (N_9601,N_8454,N_8776);
nand U9602 (N_9602,N_6700,N_6109);
nand U9603 (N_9603,N_8868,N_6899);
and U9604 (N_9604,N_6571,N_6285);
and U9605 (N_9605,N_6295,N_7143);
and U9606 (N_9606,N_6698,N_8204);
nor U9607 (N_9607,N_7538,N_6086);
nor U9608 (N_9608,N_6714,N_7319);
or U9609 (N_9609,N_7826,N_8805);
xor U9610 (N_9610,N_6486,N_8202);
or U9611 (N_9611,N_7253,N_7968);
nor U9612 (N_9612,N_6712,N_8484);
and U9613 (N_9613,N_7714,N_7637);
and U9614 (N_9614,N_7653,N_7556);
and U9615 (N_9615,N_7897,N_6719);
or U9616 (N_9616,N_6590,N_7464);
nand U9617 (N_9617,N_6920,N_8605);
xor U9618 (N_9618,N_6227,N_6237);
nor U9619 (N_9619,N_7694,N_8575);
xor U9620 (N_9620,N_8861,N_7895);
nand U9621 (N_9621,N_6062,N_8250);
nand U9622 (N_9622,N_6750,N_8329);
nand U9623 (N_9623,N_8589,N_8357);
or U9624 (N_9624,N_6028,N_7630);
and U9625 (N_9625,N_6434,N_8041);
and U9626 (N_9626,N_7734,N_8769);
nand U9627 (N_9627,N_7762,N_8048);
and U9628 (N_9628,N_6296,N_6515);
and U9629 (N_9629,N_8183,N_7809);
or U9630 (N_9630,N_7053,N_8044);
or U9631 (N_9631,N_6736,N_7595);
nor U9632 (N_9632,N_6855,N_6842);
nor U9633 (N_9633,N_7956,N_7929);
or U9634 (N_9634,N_8360,N_7294);
nor U9635 (N_9635,N_6664,N_7814);
and U9636 (N_9636,N_8078,N_7890);
nand U9637 (N_9637,N_6279,N_6447);
xor U9638 (N_9638,N_7090,N_8447);
nand U9639 (N_9639,N_6234,N_6207);
or U9640 (N_9640,N_7723,N_8229);
and U9641 (N_9641,N_7003,N_8123);
nand U9642 (N_9642,N_8755,N_6400);
and U9643 (N_9643,N_8824,N_8559);
nor U9644 (N_9644,N_6981,N_6203);
and U9645 (N_9645,N_6454,N_6181);
or U9646 (N_9646,N_6157,N_6884);
or U9647 (N_9647,N_8571,N_7284);
nand U9648 (N_9648,N_7964,N_8392);
nand U9649 (N_9649,N_6681,N_7623);
xnor U9650 (N_9650,N_6208,N_8017);
and U9651 (N_9651,N_8959,N_7931);
xor U9652 (N_9652,N_7792,N_6583);
nor U9653 (N_9653,N_8216,N_8630);
xor U9654 (N_9654,N_8472,N_8962);
or U9655 (N_9655,N_6745,N_6021);
nand U9656 (N_9656,N_7582,N_8678);
nor U9657 (N_9657,N_7720,N_8479);
nand U9658 (N_9658,N_8624,N_6679);
nor U9659 (N_9659,N_7227,N_6524);
and U9660 (N_9660,N_7023,N_7710);
nor U9661 (N_9661,N_6528,N_6231);
and U9662 (N_9662,N_6425,N_6859);
nand U9663 (N_9663,N_6066,N_8083);
or U9664 (N_9664,N_8004,N_6927);
nor U9665 (N_9665,N_6956,N_8885);
and U9666 (N_9666,N_7862,N_7189);
and U9667 (N_9667,N_7239,N_6051);
nor U9668 (N_9668,N_8570,N_7030);
or U9669 (N_9669,N_8190,N_7497);
nor U9670 (N_9670,N_6190,N_6182);
xor U9671 (N_9671,N_6173,N_8864);
nor U9672 (N_9672,N_8893,N_7638);
and U9673 (N_9673,N_6304,N_7179);
nand U9674 (N_9674,N_6350,N_7395);
nand U9675 (N_9675,N_8455,N_7174);
or U9676 (N_9676,N_6573,N_6317);
or U9677 (N_9677,N_8942,N_8773);
and U9678 (N_9678,N_8416,N_7441);
and U9679 (N_9679,N_7217,N_7329);
and U9680 (N_9680,N_8485,N_6669);
and U9681 (N_9681,N_7907,N_8625);
nand U9682 (N_9682,N_8411,N_8096);
nand U9683 (N_9683,N_7437,N_8178);
and U9684 (N_9684,N_6725,N_7921);
nand U9685 (N_9685,N_7324,N_7926);
nor U9686 (N_9686,N_6198,N_8241);
nor U9687 (N_9687,N_7392,N_7054);
and U9688 (N_9688,N_7634,N_6796);
nor U9689 (N_9689,N_7683,N_8117);
nand U9690 (N_9690,N_8350,N_8646);
nand U9691 (N_9691,N_7283,N_6982);
nor U9692 (N_9692,N_8222,N_7864);
nor U9693 (N_9693,N_8468,N_8215);
or U9694 (N_9694,N_7663,N_6194);
and U9695 (N_9695,N_7853,N_8709);
or U9696 (N_9696,N_7004,N_6497);
nand U9697 (N_9697,N_7991,N_6142);
and U9698 (N_9698,N_6475,N_8566);
nand U9699 (N_9699,N_7266,N_7214);
and U9700 (N_9700,N_8549,N_8421);
and U9701 (N_9701,N_6146,N_7278);
or U9702 (N_9702,N_6074,N_8726);
or U9703 (N_9703,N_8318,N_8375);
and U9704 (N_9704,N_8516,N_7995);
and U9705 (N_9705,N_6416,N_8506);
and U9706 (N_9706,N_6777,N_7418);
nor U9707 (N_9707,N_6942,N_6220);
nand U9708 (N_9708,N_6763,N_6856);
nor U9709 (N_9709,N_6857,N_7856);
and U9710 (N_9710,N_7839,N_7553);
nor U9711 (N_9711,N_7732,N_6952);
and U9712 (N_9712,N_6356,N_6577);
and U9713 (N_9713,N_7166,N_8040);
nor U9714 (N_9714,N_6505,N_7747);
or U9715 (N_9715,N_6247,N_8234);
nand U9716 (N_9716,N_8343,N_8063);
nand U9717 (N_9717,N_8209,N_7254);
or U9718 (N_9718,N_8348,N_7490);
or U9719 (N_9719,N_7151,N_6781);
and U9720 (N_9720,N_7724,N_6156);
and U9721 (N_9721,N_8593,N_8068);
and U9722 (N_9722,N_7428,N_7776);
and U9723 (N_9723,N_6708,N_8285);
and U9724 (N_9724,N_6179,N_7677);
or U9725 (N_9725,N_6386,N_7234);
nor U9726 (N_9726,N_8652,N_7863);
or U9727 (N_9727,N_8586,N_8701);
nor U9728 (N_9728,N_8143,N_6159);
nand U9729 (N_9729,N_6848,N_7245);
or U9730 (N_9730,N_6689,N_6090);
xnor U9731 (N_9731,N_6834,N_7746);
nand U9732 (N_9732,N_8518,N_6972);
nor U9733 (N_9733,N_6136,N_8520);
nor U9734 (N_9734,N_8450,N_7483);
nand U9735 (N_9735,N_8601,N_7865);
and U9736 (N_9736,N_6936,N_8136);
and U9737 (N_9737,N_8316,N_6091);
nand U9738 (N_9738,N_8388,N_7287);
or U9739 (N_9739,N_8854,N_8203);
nand U9740 (N_9740,N_7785,N_8114);
and U9741 (N_9741,N_7315,N_8306);
nand U9742 (N_9742,N_8162,N_7232);
nor U9743 (N_9743,N_8860,N_6168);
or U9744 (N_9744,N_6937,N_6175);
xnor U9745 (N_9745,N_8666,N_8042);
or U9746 (N_9746,N_7316,N_6861);
or U9747 (N_9747,N_8374,N_8972);
and U9748 (N_9748,N_8943,N_8159);
nor U9749 (N_9749,N_7085,N_8152);
or U9750 (N_9750,N_8390,N_7365);
nand U9751 (N_9751,N_6520,N_6287);
and U9752 (N_9752,N_7911,N_8592);
nor U9753 (N_9753,N_6426,N_8950);
nand U9754 (N_9754,N_6137,N_8955);
and U9755 (N_9755,N_8905,N_7692);
nand U9756 (N_9756,N_7487,N_6197);
and U9757 (N_9757,N_8787,N_8949);
and U9758 (N_9758,N_8914,N_8937);
or U9759 (N_9759,N_6533,N_6196);
nand U9760 (N_9760,N_8385,N_6044);
nand U9761 (N_9761,N_8151,N_7275);
and U9762 (N_9762,N_6431,N_7551);
nand U9763 (N_9763,N_8754,N_7466);
nor U9764 (N_9764,N_7422,N_7188);
nor U9765 (N_9765,N_8434,N_7735);
or U9766 (N_9766,N_6860,N_7177);
nor U9767 (N_9767,N_8686,N_6114);
or U9768 (N_9768,N_8005,N_6487);
nor U9769 (N_9769,N_8613,N_6257);
and U9770 (N_9770,N_7795,N_8277);
nand U9771 (N_9771,N_8890,N_6113);
or U9772 (N_9772,N_6523,N_7913);
and U9773 (N_9773,N_8998,N_8349);
nor U9774 (N_9774,N_6272,N_6364);
nor U9775 (N_9775,N_6097,N_7461);
and U9776 (N_9776,N_7087,N_6344);
or U9777 (N_9777,N_8409,N_8494);
or U9778 (N_9778,N_6283,N_6862);
or U9779 (N_9779,N_7454,N_7380);
nand U9780 (N_9780,N_6363,N_6782);
nand U9781 (N_9781,N_8366,N_8074);
xor U9782 (N_9782,N_8381,N_6310);
nor U9783 (N_9783,N_7154,N_8901);
nor U9784 (N_9784,N_8380,N_8659);
or U9785 (N_9785,N_8109,N_7109);
and U9786 (N_9786,N_7539,N_8925);
nor U9787 (N_9787,N_8500,N_8367);
or U9788 (N_9788,N_7452,N_8181);
or U9789 (N_9789,N_7642,N_6068);
nand U9790 (N_9790,N_6158,N_7102);
and U9791 (N_9791,N_6930,N_7111);
nand U9792 (N_9792,N_7666,N_8700);
nor U9793 (N_9793,N_6550,N_6586);
nor U9794 (N_9794,N_8296,N_7065);
or U9795 (N_9795,N_6125,N_8103);
and U9796 (N_9796,N_8263,N_8387);
or U9797 (N_9797,N_8534,N_8191);
and U9798 (N_9798,N_6600,N_8512);
nor U9799 (N_9799,N_7573,N_7970);
nand U9800 (N_9800,N_7312,N_6687);
nor U9801 (N_9801,N_8744,N_8273);
xor U9802 (N_9802,N_6692,N_7594);
or U9803 (N_9803,N_7975,N_6648);
nor U9804 (N_9804,N_8220,N_6298);
nor U9805 (N_9805,N_6755,N_7056);
nand U9806 (N_9806,N_7406,N_8095);
nand U9807 (N_9807,N_8762,N_7918);
or U9808 (N_9808,N_6178,N_8789);
or U9809 (N_9809,N_7645,N_8879);
or U9810 (N_9810,N_6752,N_6824);
and U9811 (N_9811,N_8740,N_6149);
nor U9812 (N_9812,N_7945,N_6746);
nor U9813 (N_9813,N_8487,N_7190);
nand U9814 (N_9814,N_8091,N_7293);
and U9815 (N_9815,N_8002,N_7208);
nor U9816 (N_9816,N_8560,N_8230);
and U9817 (N_9817,N_8394,N_8139);
or U9818 (N_9818,N_8641,N_7939);
or U9819 (N_9819,N_6963,N_8790);
nand U9820 (N_9820,N_6613,N_7061);
or U9821 (N_9821,N_8260,N_7569);
nor U9822 (N_9822,N_7719,N_6131);
and U9823 (N_9823,N_8899,N_6823);
nand U9824 (N_9824,N_6992,N_6609);
nor U9825 (N_9825,N_8393,N_7591);
nand U9826 (N_9826,N_8288,N_6320);
nand U9827 (N_9827,N_6957,N_7298);
or U9828 (N_9828,N_6411,N_8710);
and U9829 (N_9829,N_7860,N_7346);
nand U9830 (N_9830,N_7244,N_8293);
nand U9831 (N_9831,N_8359,N_8916);
nor U9832 (N_9832,N_8376,N_6779);
nand U9833 (N_9833,N_7688,N_6483);
or U9834 (N_9834,N_8952,N_7894);
or U9835 (N_9835,N_7885,N_8851);
nand U9836 (N_9836,N_7207,N_6143);
and U9837 (N_9837,N_8353,N_8169);
or U9838 (N_9838,N_8944,N_6996);
nand U9839 (N_9839,N_6829,N_6349);
or U9840 (N_9840,N_8598,N_7484);
nand U9841 (N_9841,N_7067,N_7549);
nand U9842 (N_9842,N_7159,N_7480);
or U9843 (N_9843,N_6732,N_8112);
or U9844 (N_9844,N_7064,N_6678);
nand U9845 (N_9845,N_8622,N_7041);
nor U9846 (N_9846,N_6262,N_6562);
nand U9847 (N_9847,N_8497,N_6948);
or U9848 (N_9848,N_8654,N_8049);
nor U9849 (N_9849,N_8228,N_8130);
or U9850 (N_9850,N_7753,N_7806);
nor U9851 (N_9851,N_7541,N_7540);
nand U9852 (N_9852,N_8210,N_6110);
and U9853 (N_9853,N_8647,N_6089);
and U9854 (N_9854,N_8906,N_7515);
nor U9855 (N_9855,N_8767,N_8177);
nor U9856 (N_9856,N_8644,N_7635);
nand U9857 (N_9857,N_8989,N_8403);
nand U9858 (N_9858,N_6177,N_6063);
nor U9859 (N_9859,N_7265,N_7602);
nor U9860 (N_9860,N_8171,N_8069);
xnor U9861 (N_9861,N_6073,N_7808);
nor U9862 (N_9862,N_8119,N_6334);
nor U9863 (N_9863,N_7381,N_8736);
nor U9864 (N_9864,N_6913,N_7059);
and U9865 (N_9865,N_8249,N_6390);
or U9866 (N_9866,N_6822,N_7260);
or U9867 (N_9867,N_6489,N_8084);
nand U9868 (N_9868,N_8312,N_6561);
and U9869 (N_9869,N_8076,N_7774);
nand U9870 (N_9870,N_8145,N_6211);
nand U9871 (N_9871,N_6035,N_8897);
nand U9872 (N_9872,N_8026,N_7262);
and U9873 (N_9873,N_6744,N_8987);
nand U9874 (N_9874,N_6501,N_7402);
nand U9875 (N_9875,N_8415,N_6711);
or U9876 (N_9876,N_8226,N_6427);
nand U9877 (N_9877,N_7268,N_8564);
or U9878 (N_9878,N_6833,N_6731);
nand U9879 (N_9879,N_7752,N_8591);
or U9880 (N_9880,N_7888,N_7277);
and U9881 (N_9881,N_8225,N_7408);
nand U9882 (N_9882,N_6270,N_7552);
or U9883 (N_9883,N_8930,N_6199);
nand U9884 (N_9884,N_7667,N_8698);
and U9885 (N_9885,N_8275,N_8207);
nor U9886 (N_9886,N_7139,N_8964);
nand U9887 (N_9887,N_6328,N_8718);
or U9888 (N_9888,N_7303,N_8633);
nor U9889 (N_9889,N_8012,N_7145);
and U9890 (N_9890,N_7492,N_7095);
nand U9891 (N_9891,N_7042,N_6504);
or U9892 (N_9892,N_6657,N_6221);
nor U9893 (N_9893,N_6015,N_6011);
and U9894 (N_9894,N_8453,N_7288);
xor U9895 (N_9895,N_8146,N_7197);
and U9896 (N_9896,N_6155,N_7676);
nand U9897 (N_9897,N_6444,N_6048);
and U9898 (N_9898,N_6171,N_7110);
nand U9899 (N_9899,N_7247,N_8715);
nand U9900 (N_9900,N_7488,N_7165);
nor U9901 (N_9901,N_7639,N_7649);
or U9902 (N_9902,N_8457,N_7871);
nand U9903 (N_9903,N_8038,N_7360);
or U9904 (N_9904,N_6625,N_8771);
xor U9905 (N_9905,N_7222,N_7389);
nor U9906 (N_9906,N_6041,N_7928);
nor U9907 (N_9907,N_7599,N_7348);
nand U9908 (N_9908,N_8881,N_8611);
nand U9909 (N_9909,N_6789,N_8345);
nand U9910 (N_9910,N_6890,N_7574);
nor U9911 (N_9911,N_8772,N_6837);
nand U9912 (N_9912,N_8517,N_7194);
and U9913 (N_9913,N_6596,N_6134);
and U9914 (N_9914,N_6301,N_7513);
xor U9915 (N_9915,N_7982,N_7032);
nand U9916 (N_9916,N_6951,N_8803);
and U9917 (N_9917,N_7397,N_8238);
nand U9918 (N_9918,N_7855,N_8775);
nand U9919 (N_9919,N_8036,N_7202);
and U9920 (N_9920,N_7604,N_6926);
nand U9921 (N_9921,N_8051,N_8902);
nand U9922 (N_9922,N_7948,N_8007);
or U9923 (N_9923,N_7498,N_6120);
or U9924 (N_9924,N_7375,N_7297);
and U9925 (N_9925,N_7744,N_7802);
and U9926 (N_9926,N_8891,N_6373);
or U9927 (N_9927,N_7330,N_6511);
and U9928 (N_9928,N_6872,N_7528);
xor U9929 (N_9929,N_6543,N_8369);
nand U9930 (N_9930,N_7934,N_7228);
and U9931 (N_9931,N_8555,N_7778);
or U9932 (N_9932,N_8639,N_8681);
nand U9933 (N_9933,N_6017,N_7148);
and U9934 (N_9934,N_8626,N_8024);
or U9935 (N_9935,N_8291,N_8407);
nor U9936 (N_9936,N_7947,N_6111);
or U9937 (N_9937,N_8980,N_6983);
and U9938 (N_9938,N_8239,N_8819);
nand U9939 (N_9939,N_6673,N_6891);
nor U9940 (N_9940,N_6644,N_6621);
and U9941 (N_9941,N_8607,N_6102);
or U9942 (N_9942,N_8538,N_6435);
nor U9943 (N_9943,N_6465,N_6532);
or U9944 (N_9944,N_6925,N_8243);
and U9945 (N_9945,N_8604,N_7340);
or U9946 (N_9946,N_7269,N_7238);
and U9947 (N_9947,N_6319,N_8791);
or U9948 (N_9948,N_7376,N_7566);
nor U9949 (N_9949,N_7773,N_6525);
and U9950 (N_9950,N_7523,N_7071);
nand U9951 (N_9951,N_6595,N_6554);
and U9952 (N_9952,N_8895,N_7276);
or U9953 (N_9953,N_6020,N_8758);
or U9954 (N_9954,N_8179,N_7973);
and U9955 (N_9955,N_6494,N_6374);
nor U9956 (N_9956,N_8845,N_7242);
nand U9957 (N_9957,N_6478,N_6395);
or U9958 (N_9958,N_7636,N_7387);
nor U9959 (N_9959,N_7588,N_7601);
nand U9960 (N_9960,N_8992,N_8003);
or U9961 (N_9961,N_6598,N_8679);
nand U9962 (N_9962,N_6935,N_8050);
and U9963 (N_9963,N_6288,N_8483);
or U9964 (N_9964,N_8848,N_7870);
or U9965 (N_9965,N_8651,N_8533);
and U9966 (N_9966,N_8221,N_7230);
nor U9967 (N_9967,N_8213,N_7542);
nand U9968 (N_9968,N_6397,N_6423);
and U9969 (N_9969,N_6246,N_7851);
nor U9970 (N_9970,N_8053,N_8107);
nand U9971 (N_9971,N_8401,N_6923);
nor U9972 (N_9972,N_6914,N_7522);
nor U9973 (N_9973,N_8469,N_8608);
and U9974 (N_9974,N_8399,N_6076);
or U9975 (N_9975,N_8176,N_6441);
nor U9976 (N_9976,N_6432,N_6223);
or U9977 (N_9977,N_8236,N_8197);
nor U9978 (N_9978,N_8811,N_6599);
nand U9979 (N_9979,N_8058,N_8527);
or U9980 (N_9980,N_6212,N_6786);
nor U9981 (N_9981,N_6016,N_6420);
or U9982 (N_9982,N_6915,N_6406);
or U9983 (N_9983,N_6662,N_6002);
nand U9984 (N_9984,N_8922,N_8274);
and U9985 (N_9985,N_8634,N_8217);
or U9986 (N_9986,N_8995,N_6378);
nand U9987 (N_9987,N_8730,N_8692);
nor U9988 (N_9988,N_6047,N_6715);
or U9989 (N_9989,N_7842,N_8001);
or U9990 (N_9990,N_8043,N_7390);
and U9991 (N_9991,N_8514,N_8284);
or U9992 (N_9992,N_6348,N_6010);
nand U9993 (N_9993,N_8297,N_7263);
and U9994 (N_9994,N_6880,N_7134);
or U9995 (N_9995,N_8643,N_7699);
and U9996 (N_9996,N_8938,N_7665);
and U9997 (N_9997,N_7844,N_6800);
nand U9998 (N_9998,N_7584,N_8382);
or U9999 (N_9999,N_7904,N_7777);
or U10000 (N_10000,N_6452,N_7410);
nand U10001 (N_10001,N_8034,N_8849);
nand U10002 (N_10002,N_7967,N_6959);
nor U10003 (N_10003,N_7072,N_8166);
nand U10004 (N_10004,N_6336,N_6232);
or U10005 (N_10005,N_8030,N_8585);
or U10006 (N_10006,N_6184,N_8000);
and U10007 (N_10007,N_7289,N_6768);
or U10008 (N_10008,N_7530,N_7654);
nand U10009 (N_10009,N_8321,N_7898);
or U10010 (N_10010,N_6580,N_7578);
nor U10011 (N_10011,N_6012,N_7305);
nor U10012 (N_10012,N_8310,N_7285);
xnor U10013 (N_10013,N_8821,N_8354);
or U10014 (N_10014,N_7083,N_8482);
and U10015 (N_10015,N_6909,N_7848);
nand U10016 (N_10016,N_8867,N_8774);
or U10017 (N_10017,N_7662,N_6219);
nand U10018 (N_10018,N_7560,N_6507);
nand U10019 (N_10019,N_7989,N_8923);
nand U10020 (N_10020,N_8829,N_8649);
or U10021 (N_10021,N_8940,N_6369);
nor U10022 (N_10022,N_8705,N_7282);
or U10023 (N_10023,N_8172,N_8502);
nand U10024 (N_10024,N_7493,N_6422);
nand U10025 (N_10025,N_6724,N_7500);
nand U10026 (N_10026,N_7439,N_7112);
and U10027 (N_10027,N_6558,N_8287);
and U10028 (N_10028,N_7017,N_7527);
or U10029 (N_10029,N_6470,N_6318);
or U10030 (N_10030,N_8792,N_6245);
or U10031 (N_10031,N_8741,N_8667);
and U10032 (N_10032,N_6057,N_8311);
or U10033 (N_10033,N_7925,N_6825);
and U10034 (N_10034,N_8132,N_8584);
and U10035 (N_10035,N_8663,N_8101);
nand U10036 (N_10036,N_6780,N_8834);
nor U10037 (N_10037,N_6186,N_6836);
nand U10038 (N_10038,N_6696,N_6587);
and U10039 (N_10039,N_8338,N_6152);
nor U10040 (N_10040,N_8547,N_7608);
nand U10041 (N_10041,N_8684,N_6370);
nand U10042 (N_10042,N_8298,N_6302);
nor U10043 (N_10043,N_8504,N_8315);
nor U10044 (N_10044,N_8729,N_6024);
nor U10045 (N_10045,N_7643,N_6387);
nand U10046 (N_10046,N_8466,N_8645);
or U10047 (N_10047,N_6101,N_7068);
and U10048 (N_10048,N_8081,N_8115);
and U10049 (N_10049,N_7990,N_6396);
nand U10050 (N_10050,N_6659,N_8597);
or U10051 (N_10051,N_7157,N_8665);
nor U10052 (N_10052,N_8746,N_8750);
nand U10053 (N_10053,N_6988,N_6195);
or U10054 (N_10054,N_6027,N_7955);
nand U10055 (N_10055,N_6255,N_6733);
nand U10056 (N_10056,N_6308,N_7162);
and U10057 (N_10057,N_6335,N_6728);
or U10058 (N_10058,N_6954,N_7974);
and U10059 (N_10059,N_6799,N_8843);
nor U10060 (N_10060,N_6226,N_6144);
nand U10061 (N_10061,N_7460,N_8489);
or U10062 (N_10062,N_6739,N_7629);
xor U10063 (N_10063,N_6005,N_6660);
nor U10064 (N_10064,N_7120,N_6918);
and U10065 (N_10065,N_7759,N_8759);
or U10066 (N_10066,N_8264,N_8722);
nor U10067 (N_10067,N_8075,N_6870);
nand U10068 (N_10068,N_6947,N_6987);
and U10069 (N_10069,N_6026,N_7892);
nand U10070 (N_10070,N_8465,N_8244);
nand U10071 (N_10071,N_7121,N_8904);
and U10072 (N_10072,N_8693,N_6921);
nor U10073 (N_10073,N_8567,N_8070);
and U10074 (N_10074,N_6908,N_7859);
and U10075 (N_10075,N_6634,N_7937);
and U10076 (N_10076,N_8965,N_7779);
nor U10077 (N_10077,N_6436,N_6289);
and U10078 (N_10078,N_6079,N_6403);
nor U10079 (N_10079,N_7754,N_7119);
nand U10080 (N_10080,N_7953,N_6242);
nand U10081 (N_10081,N_7902,N_8958);
or U10082 (N_10082,N_8270,N_6481);
and U10083 (N_10083,N_8981,N_7984);
and U10084 (N_10084,N_6013,N_8111);
and U10085 (N_10085,N_8892,N_6650);
and U10086 (N_10086,N_8478,N_8224);
nand U10087 (N_10087,N_6672,N_7577);
or U10088 (N_10088,N_6126,N_8544);
nand U10089 (N_10089,N_8511,N_7679);
nand U10090 (N_10090,N_8982,N_7992);
nor U10091 (N_10091,N_7618,N_6106);
nor U10092 (N_10092,N_6514,N_6697);
or U10093 (N_10093,N_7126,N_6653);
nor U10094 (N_10094,N_8090,N_8339);
or U10095 (N_10095,N_7363,N_7828);
or U10096 (N_10096,N_8734,N_7048);
and U10097 (N_10097,N_6001,N_7846);
nand U10098 (N_10098,N_6622,N_6174);
and U10099 (N_10099,N_7506,N_6556);
nand U10100 (N_10100,N_8476,N_7482);
nand U10101 (N_10101,N_7587,N_7051);
nand U10102 (N_10102,N_7373,N_6252);
nor U10103 (N_10103,N_7186,N_7708);
or U10104 (N_10104,N_7664,N_6401);
nand U10105 (N_10105,N_8060,N_6903);
nand U10106 (N_10106,N_7045,N_7326);
xor U10107 (N_10107,N_8993,N_8292);
nand U10108 (N_10108,N_7404,N_6368);
and U10109 (N_10109,N_8749,N_6393);
or U10110 (N_10110,N_8831,N_7625);
xnor U10111 (N_10111,N_8161,N_6734);
nor U10112 (N_10112,N_7384,N_6663);
nand U10113 (N_10113,N_7977,N_8231);
and U10114 (N_10114,N_8971,N_7181);
nor U10115 (N_10115,N_8523,N_7672);
or U10116 (N_10116,N_7036,N_7874);
xnor U10117 (N_10117,N_6898,N_6894);
nand U10118 (N_10118,N_7458,N_6115);
nor U10119 (N_10119,N_7905,N_8137);
or U10120 (N_10120,N_8768,N_7433);
nor U10121 (N_10121,N_6123,N_8200);
or U10122 (N_10122,N_8432,N_8838);
nor U10123 (N_10123,N_8988,N_7962);
nor U10124 (N_10124,N_7354,N_6589);
and U10125 (N_10125,N_7509,N_6813);
nor U10126 (N_10126,N_6381,N_7478);
nand U10127 (N_10127,N_8397,N_6383);
and U10128 (N_10128,N_8548,N_8817);
or U10129 (N_10129,N_8028,N_7681);
nand U10130 (N_10130,N_8037,N_6928);
nand U10131 (N_10131,N_6522,N_8612);
nand U10132 (N_10132,N_7876,N_8946);
nor U10133 (N_10133,N_7343,N_6192);
and U10134 (N_10134,N_6846,N_8033);
nor U10135 (N_10135,N_8302,N_6014);
nand U10136 (N_10136,N_8456,N_6128);
and U10137 (N_10137,N_7044,N_7301);
and U10138 (N_10138,N_8888,N_8724);
nor U10139 (N_10139,N_6738,N_8064);
and U10140 (N_10140,N_6617,N_7344);
or U10141 (N_10141,N_7611,N_8192);
nor U10142 (N_10142,N_8976,N_8725);
nand U10143 (N_10143,N_7650,N_7503);
nor U10144 (N_10144,N_6124,N_8116);
nor U10145 (N_10145,N_8020,N_7803);
nand U10146 (N_10146,N_8563,N_6415);
or U10147 (N_10147,N_6685,N_8227);
and U10148 (N_10148,N_7170,N_6879);
nor U10149 (N_10149,N_8703,N_7261);
or U10150 (N_10150,N_7436,N_8818);
nor U10151 (N_10151,N_6249,N_8332);
nand U10152 (N_10152,N_7043,N_6019);
and U10153 (N_10153,N_7300,N_7685);
or U10154 (N_10154,N_8470,N_6682);
or U10155 (N_10155,N_6684,N_7280);
xnor U10156 (N_10156,N_8997,N_7824);
nor U10157 (N_10157,N_6313,N_7153);
and U10158 (N_10158,N_6405,N_6228);
nor U10159 (N_10159,N_6628,N_6643);
nand U10160 (N_10160,N_6200,N_7796);
nor U10161 (N_10161,N_7680,N_6647);
or U10162 (N_10162,N_6610,N_7626);
or U10163 (N_10163,N_7415,N_8631);
nand U10164 (N_10164,N_6052,N_8685);
nor U10165 (N_10165,N_8142,N_8449);
nand U10166 (N_10166,N_6747,N_7335);
nand U10167 (N_10167,N_7205,N_8164);
nor U10168 (N_10168,N_6251,N_7695);
and U10169 (N_10169,N_8283,N_8481);
nand U10170 (N_10170,N_6667,N_8653);
nor U10171 (N_10171,N_7729,N_7555);
and U10172 (N_10172,N_6096,N_7311);
and U10173 (N_10173,N_6748,N_8061);
nand U10174 (N_10174,N_6274,N_7345);
nor U10175 (N_10175,N_8794,N_6637);
or U10176 (N_10176,N_7414,N_8856);
and U10177 (N_10177,N_6771,N_8150);
nand U10178 (N_10178,N_6372,N_7473);
and U10179 (N_10179,N_6795,N_6093);
or U10180 (N_10180,N_8778,N_6699);
nor U10181 (N_10181,N_6843,N_7026);
xor U10182 (N_10182,N_6402,N_6337);
nand U10183 (N_10183,N_7993,N_6608);
and U10184 (N_10184,N_6783,N_7583);
nor U10185 (N_10185,N_7122,N_7922);
xor U10186 (N_10186,N_8066,N_7589);
nor U10187 (N_10187,N_8973,N_6083);
nand U10188 (N_10188,N_7715,N_8841);
or U10189 (N_10189,N_6100,N_8448);
nor U10190 (N_10190,N_7443,N_7745);
nor U10191 (N_10191,N_8256,N_7526);
and U10192 (N_10192,N_8552,N_6917);
and U10193 (N_10193,N_8820,N_7815);
or U10194 (N_10194,N_8873,N_7369);
or U10195 (N_10195,N_8869,N_7088);
and U10196 (N_10196,N_6421,N_8908);
and U10197 (N_10197,N_6618,N_7219);
and U10198 (N_10198,N_7434,N_8743);
nor U10199 (N_10199,N_6389,N_7822);
nand U10200 (N_10200,N_8855,N_6088);
nand U10201 (N_10201,N_8257,N_7847);
or U10202 (N_10202,N_7096,N_7106);
or U10203 (N_10203,N_6563,N_7115);
nand U10204 (N_10204,N_7378,N_6566);
or U10205 (N_10205,N_7866,N_8994);
nand U10206 (N_10206,N_8568,N_6492);
nand U10207 (N_10207,N_8313,N_6135);
or U10208 (N_10208,N_7548,N_8799);
nor U10209 (N_10209,N_6636,N_7883);
nor U10210 (N_10210,N_7617,N_6007);
nand U10211 (N_10211,N_8147,N_7409);
nor U10212 (N_10212,N_8408,N_7035);
or U10213 (N_10213,N_7996,N_8782);
or U10214 (N_10214,N_6030,N_8921);
nand U10215 (N_10215,N_6592,N_8211);
nand U10216 (N_10216,N_7903,N_8878);
and U10217 (N_10217,N_6809,N_8423);
xor U10218 (N_10218,N_8158,N_6491);
nand U10219 (N_10219,N_8170,N_6280);
nand U10220 (N_10220,N_6316,N_8690);
or U10221 (N_10221,N_6056,N_8532);
and U10222 (N_10222,N_6706,N_7031);
nor U10223 (N_10223,N_8031,N_7886);
nand U10224 (N_10224,N_7444,N_6670);
and U10225 (N_10225,N_7858,N_7660);
nor U10226 (N_10226,N_7272,N_8716);
and U10227 (N_10227,N_6049,N_8341);
nand U10228 (N_10228,N_6623,N_7093);
or U10229 (N_10229,N_7580,N_8706);
nor U10230 (N_10230,N_7141,N_8784);
nand U10231 (N_10231,N_7532,N_8727);
and U10232 (N_10232,N_7562,N_8325);
nand U10233 (N_10233,N_8887,N_6803);
nor U10234 (N_10234,N_7849,N_7050);
nand U10235 (N_10235,N_7229,N_6294);
xnor U10236 (N_10236,N_8106,N_7770);
nand U10237 (N_10237,N_8248,N_7367);
nand U10238 (N_10238,N_8556,N_6438);
and U10239 (N_10239,N_8424,N_8839);
or U10240 (N_10240,N_6325,N_6688);
xor U10241 (N_10241,N_8632,N_7336);
nand U10242 (N_10242,N_7130,N_6686);
or U10243 (N_10243,N_7107,N_8189);
nand U10244 (N_10244,N_7368,N_8853);
or U10245 (N_10245,N_8419,N_8233);
and U10246 (N_10246,N_6902,N_8540);
and U10247 (N_10247,N_6440,N_8461);
nand U10248 (N_10248,N_7899,N_7382);
or U10249 (N_10249,N_7136,N_6521);
nand U10250 (N_10250,N_7908,N_7199);
nor U10251 (N_10251,N_8751,N_6924);
and U10252 (N_10252,N_7495,N_8335);
or U10253 (N_10253,N_8966,N_7022);
or U10254 (N_10254,N_7619,N_7952);
nor U10255 (N_10255,N_8953,N_6391);
nor U10256 (N_10256,N_7742,N_8606);
or U10257 (N_10257,N_8144,N_8636);
and U10258 (N_10258,N_7543,N_7420);
xor U10259 (N_10259,N_7726,N_8580);
xor U10260 (N_10260,N_6312,N_7203);
and U10261 (N_10261,N_6980,N_6099);
nor U10262 (N_10262,N_6331,N_6869);
nand U10263 (N_10263,N_6306,N_6911);
or U10264 (N_10264,N_8015,N_8093);
and U10265 (N_10265,N_8327,N_8501);
nand U10266 (N_10266,N_7098,N_6680);
and U10267 (N_10267,N_7682,N_8029);
nor U10268 (N_10268,N_8442,N_6332);
nand U10269 (N_10269,N_8640,N_8694);
nand U10270 (N_10270,N_8102,N_6291);
or U10271 (N_10271,N_7518,N_7831);
or U10272 (N_10272,N_6375,N_7507);
or U10273 (N_10273,N_8173,N_7514);
or U10274 (N_10274,N_7318,N_7400);
nand U10275 (N_10275,N_8886,N_7477);
nor U10276 (N_10276,N_6385,N_6654);
nand U10277 (N_10277,N_8804,N_6238);
nor U10278 (N_10278,N_8761,N_8731);
nor U10279 (N_10279,N_6691,N_8503);
or U10280 (N_10280,N_6889,N_8342);
nor U10281 (N_10281,N_8153,N_8100);
or U10282 (N_10282,N_8745,N_6877);
nor U10283 (N_10283,N_8420,N_7307);
and U10284 (N_10284,N_7201,N_6805);
or U10285 (N_10285,N_6077,N_8193);
nor U10286 (N_10286,N_8188,N_6615);
or U10287 (N_10287,N_6412,N_8205);
nor U10288 (N_10288,N_8118,N_8167);
nand U10289 (N_10289,N_8175,N_7388);
nand U10290 (N_10290,N_6635,N_7605);
nand U10291 (N_10291,N_8148,N_6713);
and U10292 (N_10292,N_7833,N_8671);
nor U10293 (N_10293,N_7850,N_7568);
nor U10294 (N_10294,N_8301,N_6276);
and U10295 (N_10295,N_8088,N_8595);
nand U10296 (N_10296,N_8739,N_6866);
or U10297 (N_10297,N_6490,N_8669);
or U10298 (N_10298,N_8577,N_7741);
and U10299 (N_10299,N_8551,N_6754);
and U10300 (N_10300,N_6333,N_7950);
nor U10301 (N_10301,N_7873,N_6649);
or U10302 (N_10302,N_8833,N_6922);
and U10303 (N_10303,N_7581,N_8777);
nor U10304 (N_10304,N_8035,N_7976);
nand U10305 (N_10305,N_7274,N_7077);
nand U10306 (N_10306,N_6451,N_8857);
or U10307 (N_10307,N_8156,N_6080);
or U10308 (N_10308,N_8510,N_6551);
or U10309 (N_10309,N_6652,N_7445);
nor U10310 (N_10310,N_6224,N_7332);
nor U10311 (N_10311,N_6327,N_7712);
nor U10312 (N_10312,N_6968,N_7007);
xor U10313 (N_10313,N_8047,N_6060);
and U10314 (N_10314,N_6087,N_8430);
nor U10315 (N_10315,N_8427,N_6054);
nand U10316 (N_10316,N_8023,N_7008);
nand U10317 (N_10317,N_6105,N_7718);
or U10318 (N_10318,N_7101,N_8870);
and U10319 (N_10319,N_8748,N_6498);
nand U10320 (N_10320,N_6229,N_7700);
and U10321 (N_10321,N_6839,N_8977);
nand U10322 (N_10322,N_6710,N_7882);
nand U10323 (N_10323,N_8180,N_6127);
nor U10324 (N_10324,N_6323,N_7356);
or U10325 (N_10325,N_8695,N_6766);
or U10326 (N_10326,N_7613,N_7097);
nand U10327 (N_10327,N_6351,N_6353);
and U10328 (N_10328,N_7451,N_8871);
nand U10329 (N_10329,N_8208,N_8404);
and U10330 (N_10330,N_8452,N_7279);
and U10331 (N_10331,N_8846,N_8413);
nor U10332 (N_10332,N_7730,N_8865);
and U10333 (N_10333,N_7600,N_6468);
and U10334 (N_10334,N_6549,N_7547);
and U10335 (N_10335,N_7994,N_7485);
nand U10336 (N_10336,N_8911,N_6716);
and U10337 (N_10337,N_7640,N_8440);
and U10338 (N_10338,N_7281,N_7673);
xor U10339 (N_10339,N_6176,N_8847);
nor U10340 (N_10340,N_7707,N_6791);
or U10341 (N_10341,N_6814,N_7450);
and U10342 (N_10342,N_7349,N_6170);
and U10343 (N_10343,N_8067,N_8025);
nand U10344 (N_10344,N_7076,N_8126);
or U10345 (N_10345,N_8635,N_7771);
nand U10346 (N_10346,N_7772,N_6418);
nor U10347 (N_10347,N_8884,N_6499);
and U10348 (N_10348,N_6624,N_8735);
nor U10349 (N_10349,N_7200,N_6107);
nand U10350 (N_10350,N_7221,N_7259);
nor U10351 (N_10351,N_6008,N_8433);
and U10352 (N_10352,N_6032,N_6502);
nor U10353 (N_10353,N_8235,N_6474);
nand U10354 (N_10354,N_8936,N_6906);
xnor U10355 (N_10355,N_6640,N_7798);
xnor U10356 (N_10356,N_7696,N_8160);
nand U10357 (N_10357,N_8862,N_7775);
and U10358 (N_10358,N_8813,N_7596);
nand U10359 (N_10359,N_8525,N_7084);
and U10360 (N_10360,N_6085,N_8628);
nor U10361 (N_10361,N_7424,N_7033);
nor U10362 (N_10362,N_7938,N_8364);
nor U10363 (N_10363,N_7013,N_8587);
nand U10364 (N_10364,N_6584,N_6827);
and U10365 (N_10365,N_7499,N_6145);
or U10366 (N_10366,N_6612,N_7944);
nor U10367 (N_10367,N_8445,N_6433);
and U10368 (N_10368,N_8990,N_6875);
or U10369 (N_10369,N_8912,N_8187);
nand U10370 (N_10370,N_7889,N_7661);
nor U10371 (N_10371,N_6912,N_6046);
nor U10372 (N_10372,N_8753,N_8094);
and U10373 (N_10373,N_8756,N_8129);
nor U10374 (N_10374,N_8055,N_7161);
nand U10375 (N_10375,N_6588,N_6204);
and U10376 (N_10376,N_7534,N_6072);
or U10377 (N_10377,N_6239,N_8766);
nand U10378 (N_10378,N_6376,N_6999);
nand U10379 (N_10379,N_8121,N_6815);
and U10380 (N_10380,N_8537,N_7647);
nand U10381 (N_10381,N_8352,N_6876);
nand U10382 (N_10382,N_7184,N_6979);
and U10383 (N_10383,N_6977,N_8410);
xor U10384 (N_10384,N_7308,N_7867);
nor U10385 (N_10385,N_7758,N_6394);
nand U10386 (N_10386,N_7920,N_6718);
nand U10387 (N_10387,N_7142,N_8723);
or U10388 (N_10388,N_8707,N_7857);
and U10389 (N_10389,N_7603,N_7286);
nand U10390 (N_10390,N_8490,N_7531);
and U10391 (N_10391,N_7668,N_8664);
and U10392 (N_10392,N_7249,N_7501);
nor U10393 (N_10393,N_6321,N_7321);
nor U10394 (N_10394,N_8320,N_7333);
nand U10395 (N_10395,N_7590,N_6960);
and U10396 (N_10396,N_6579,N_7837);
nand U10397 (N_10397,N_8978,N_6801);
and U10398 (N_10398,N_6776,N_7783);
nand U10399 (N_10399,N_7933,N_8765);
nor U10400 (N_10400,N_6450,N_7868);
or U10401 (N_10401,N_7981,N_8286);
or U10402 (N_10402,N_8657,N_6804);
or U10403 (N_10403,N_8110,N_6267);
nand U10404 (N_10404,N_7971,N_7519);
and U10405 (N_10405,N_7173,N_8951);
and U10406 (N_10406,N_8340,N_7146);
nor U10407 (N_10407,N_7923,N_7066);
nand U10408 (N_10408,N_6025,N_6480);
nand U10409 (N_10409,N_6671,N_7193);
and U10410 (N_10410,N_7237,N_8289);
and U10411 (N_10411,N_7256,N_7508);
or U10412 (N_10412,N_6139,N_8935);
or U10413 (N_10413,N_6735,N_7900);
nor U10414 (N_10414,N_8128,N_7192);
nor U10415 (N_10415,N_6206,N_7472);
nor U10416 (N_10416,N_8917,N_6467);
nand U10417 (N_10417,N_6329,N_7291);
and U10418 (N_10418,N_8786,N_6885);
and U10419 (N_10419,N_6150,N_8650);
and U10420 (N_10420,N_7689,N_6895);
and U10421 (N_10421,N_7879,N_8542);
nand U10422 (N_10422,N_8253,N_6290);
nand U10423 (N_10423,N_6404,N_8796);
or U10424 (N_10424,N_8872,N_8324);
nand U10425 (N_10425,N_6695,N_8714);
nor U10426 (N_10426,N_7767,N_8521);
and U10427 (N_10427,N_8206,N_7786);
nand U10428 (N_10428,N_6729,N_7371);
or U10429 (N_10429,N_6271,N_6367);
nor U10430 (N_10430,N_8194,N_8439);
nor U10431 (N_10431,N_8672,N_6974);
or U10432 (N_10432,N_6730,N_8062);
or U10433 (N_10433,N_8737,N_7810);
or U10434 (N_10434,N_6095,N_7468);
nand U10435 (N_10435,N_7125,N_6129);
nor U10436 (N_10436,N_7987,N_7310);
or U10437 (N_10437,N_6658,N_6340);
nand U10438 (N_10438,N_7080,N_7561);
or U10439 (N_10439,N_8333,N_7021);
nand U10440 (N_10440,N_8059,N_8071);
or U10441 (N_10441,N_8154,N_6527);
nand U10442 (N_10442,N_6646,N_7446);
or U10443 (N_10443,N_7701,N_8422);
nand U10444 (N_10444,N_6330,N_7455);
nor U10445 (N_10445,N_8218,N_8252);
and U10446 (N_10446,N_6233,N_6473);
nand U10447 (N_10447,N_8932,N_7512);
and U10448 (N_10448,N_8974,N_8859);
nand U10449 (N_10449,N_6496,N_6209);
or U10450 (N_10450,N_6892,N_7784);
nor U10451 (N_10451,N_8983,N_8691);
and U10452 (N_10452,N_8852,N_7657);
nor U10453 (N_10453,N_6882,N_6315);
or U10454 (N_10454,N_6568,N_7258);
and U10455 (N_10455,N_7062,N_8462);
and U10456 (N_10456,N_6457,N_8546);
nand U10457 (N_10457,N_8305,N_6971);
and U10458 (N_10458,N_7671,N_6548);
nor U10459 (N_10459,N_8662,N_8272);
and U10460 (N_10460,N_6380,N_7755);
or U10461 (N_10461,N_8303,N_8336);
or U10462 (N_10462,N_6512,N_8957);
xor U10463 (N_10463,N_8968,N_6428);
and U10464 (N_10464,N_6485,N_7155);
nor U10465 (N_10465,N_7144,N_8405);
nor U10466 (N_10466,N_6210,N_6675);
nor U10467 (N_10467,N_7212,N_7516);
or U10468 (N_10468,N_7046,N_7825);
and U10469 (N_10469,N_6216,N_7073);
nor U10470 (N_10470,N_6758,N_8400);
nand U10471 (N_10471,N_7965,N_7164);
nor U10472 (N_10472,N_6161,N_8219);
or U10473 (N_10473,N_8279,N_8565);
and U10474 (N_10474,N_6303,N_8351);
or U10475 (N_10475,N_6812,N_6460);
and U10476 (N_10476,N_8330,N_7011);
and U10477 (N_10477,N_6371,N_6929);
or U10478 (N_10478,N_8282,N_6849);
or U10479 (N_10479,N_6248,N_7366);
nor U10480 (N_10480,N_8337,N_6263);
nor U10481 (N_10481,N_8600,N_7391);
or U10482 (N_10482,N_7827,N_6555);
or U10483 (N_10483,N_7127,N_7355);
nand U10484 (N_10484,N_6854,N_7960);
nor U10485 (N_10485,N_6361,N_6281);
and U10486 (N_10486,N_8697,N_6240);
xor U10487 (N_10487,N_7593,N_6585);
nor U10488 (N_10488,N_8009,N_6243);
nand U10489 (N_10489,N_7823,N_7394);
nand U10490 (N_10490,N_7429,N_8022);
or U10491 (N_10491,N_7196,N_6850);
nor U10492 (N_10492,N_7564,N_6342);
or U10493 (N_10493,N_7832,N_6078);
and U10494 (N_10494,N_7740,N_6973);
nor U10495 (N_10495,N_7264,N_6148);
nand U10496 (N_10496,N_8322,N_6904);
or U10497 (N_10497,N_8240,N_6774);
and U10498 (N_10498,N_8099,N_8334);
nand U10499 (N_10499,N_7854,N_7014);
and U10500 (N_10500,N_7970,N_8753);
or U10501 (N_10501,N_6829,N_7205);
and U10502 (N_10502,N_8320,N_6916);
or U10503 (N_10503,N_6575,N_6094);
and U10504 (N_10504,N_8790,N_8624);
nand U10505 (N_10505,N_7537,N_7843);
and U10506 (N_10506,N_8001,N_6179);
or U10507 (N_10507,N_8362,N_6285);
nand U10508 (N_10508,N_8153,N_8716);
and U10509 (N_10509,N_7713,N_8483);
or U10510 (N_10510,N_7432,N_8430);
or U10511 (N_10511,N_6696,N_8408);
or U10512 (N_10512,N_7665,N_6855);
and U10513 (N_10513,N_8492,N_6837);
or U10514 (N_10514,N_7752,N_7846);
or U10515 (N_10515,N_6174,N_8043);
and U10516 (N_10516,N_7696,N_7041);
nor U10517 (N_10517,N_8912,N_6550);
nor U10518 (N_10518,N_8906,N_8704);
nand U10519 (N_10519,N_6528,N_8512);
nand U10520 (N_10520,N_6155,N_6186);
nor U10521 (N_10521,N_8092,N_6329);
nor U10522 (N_10522,N_7487,N_8730);
and U10523 (N_10523,N_8345,N_8722);
and U10524 (N_10524,N_7821,N_6856);
nor U10525 (N_10525,N_6641,N_8164);
nor U10526 (N_10526,N_8992,N_8806);
and U10527 (N_10527,N_8806,N_8521);
nor U10528 (N_10528,N_8426,N_8830);
and U10529 (N_10529,N_7096,N_8185);
and U10530 (N_10530,N_6313,N_7417);
or U10531 (N_10531,N_7091,N_6348);
nand U10532 (N_10532,N_7188,N_8050);
or U10533 (N_10533,N_8294,N_8212);
and U10534 (N_10534,N_7895,N_6687);
nand U10535 (N_10535,N_8599,N_8832);
nor U10536 (N_10536,N_8709,N_7756);
and U10537 (N_10537,N_8622,N_7935);
and U10538 (N_10538,N_6538,N_8716);
nor U10539 (N_10539,N_7005,N_7183);
nor U10540 (N_10540,N_6444,N_8292);
nor U10541 (N_10541,N_8565,N_7014);
or U10542 (N_10542,N_7673,N_8602);
and U10543 (N_10543,N_8266,N_8900);
nor U10544 (N_10544,N_6900,N_7122);
or U10545 (N_10545,N_6555,N_7276);
and U10546 (N_10546,N_6970,N_8458);
nor U10547 (N_10547,N_7220,N_7482);
and U10548 (N_10548,N_7446,N_7559);
and U10549 (N_10549,N_6306,N_7197);
or U10550 (N_10550,N_8382,N_7095);
nand U10551 (N_10551,N_6677,N_8065);
or U10552 (N_10552,N_8693,N_6645);
or U10553 (N_10553,N_8274,N_8008);
nor U10554 (N_10554,N_6755,N_7542);
nand U10555 (N_10555,N_6895,N_8461);
or U10556 (N_10556,N_7031,N_7407);
nand U10557 (N_10557,N_7349,N_6648);
and U10558 (N_10558,N_7338,N_8642);
nor U10559 (N_10559,N_6247,N_8317);
and U10560 (N_10560,N_8563,N_6099);
nand U10561 (N_10561,N_8204,N_7832);
nand U10562 (N_10562,N_7147,N_7860);
nor U10563 (N_10563,N_7363,N_6313);
and U10564 (N_10564,N_8099,N_7094);
or U10565 (N_10565,N_7743,N_8871);
nor U10566 (N_10566,N_7476,N_8502);
or U10567 (N_10567,N_8179,N_6968);
and U10568 (N_10568,N_7375,N_6090);
or U10569 (N_10569,N_8545,N_6772);
and U10570 (N_10570,N_7661,N_7587);
or U10571 (N_10571,N_6446,N_8274);
or U10572 (N_10572,N_8912,N_8595);
nor U10573 (N_10573,N_8235,N_7050);
nand U10574 (N_10574,N_7892,N_8602);
and U10575 (N_10575,N_7116,N_6462);
and U10576 (N_10576,N_7543,N_8624);
nor U10577 (N_10577,N_7814,N_7323);
and U10578 (N_10578,N_6552,N_6753);
nand U10579 (N_10579,N_8798,N_8188);
nand U10580 (N_10580,N_6152,N_6647);
or U10581 (N_10581,N_7660,N_6865);
or U10582 (N_10582,N_7973,N_8499);
nor U10583 (N_10583,N_7216,N_6375);
or U10584 (N_10584,N_7372,N_7583);
nand U10585 (N_10585,N_8400,N_8919);
nand U10586 (N_10586,N_6532,N_8273);
and U10587 (N_10587,N_6835,N_7887);
or U10588 (N_10588,N_8929,N_7474);
or U10589 (N_10589,N_6508,N_8028);
and U10590 (N_10590,N_8993,N_7397);
nand U10591 (N_10591,N_8742,N_6018);
nand U10592 (N_10592,N_6763,N_8175);
nor U10593 (N_10593,N_7512,N_8966);
nand U10594 (N_10594,N_7235,N_7563);
nand U10595 (N_10595,N_7331,N_7903);
and U10596 (N_10596,N_6781,N_7773);
and U10597 (N_10597,N_8034,N_7378);
nand U10598 (N_10598,N_6187,N_6365);
and U10599 (N_10599,N_8628,N_6063);
or U10600 (N_10600,N_7146,N_7384);
or U10601 (N_10601,N_7931,N_8374);
nor U10602 (N_10602,N_6737,N_8493);
and U10603 (N_10603,N_7290,N_8092);
nor U10604 (N_10604,N_8222,N_8584);
and U10605 (N_10605,N_7800,N_6227);
and U10606 (N_10606,N_8089,N_7551);
and U10607 (N_10607,N_8509,N_8205);
xnor U10608 (N_10608,N_6128,N_8683);
and U10609 (N_10609,N_7143,N_6358);
or U10610 (N_10610,N_6267,N_6864);
and U10611 (N_10611,N_8337,N_7223);
nor U10612 (N_10612,N_8260,N_6181);
nor U10613 (N_10613,N_6007,N_7404);
nand U10614 (N_10614,N_7047,N_8760);
xnor U10615 (N_10615,N_6848,N_6569);
or U10616 (N_10616,N_6417,N_6362);
nand U10617 (N_10617,N_8016,N_8707);
nand U10618 (N_10618,N_6388,N_7290);
and U10619 (N_10619,N_6407,N_7953);
or U10620 (N_10620,N_8016,N_8334);
and U10621 (N_10621,N_6358,N_7249);
or U10622 (N_10622,N_6779,N_8338);
and U10623 (N_10623,N_8799,N_7468);
nand U10624 (N_10624,N_8083,N_7127);
nor U10625 (N_10625,N_6494,N_8754);
nand U10626 (N_10626,N_6391,N_7863);
or U10627 (N_10627,N_7362,N_8975);
and U10628 (N_10628,N_6839,N_6648);
and U10629 (N_10629,N_7211,N_7353);
and U10630 (N_10630,N_8011,N_8905);
or U10631 (N_10631,N_6319,N_6572);
and U10632 (N_10632,N_8982,N_7762);
nor U10633 (N_10633,N_8573,N_8210);
and U10634 (N_10634,N_6791,N_8119);
and U10635 (N_10635,N_7056,N_6049);
or U10636 (N_10636,N_6872,N_8243);
nand U10637 (N_10637,N_8251,N_8874);
nand U10638 (N_10638,N_7134,N_8745);
xnor U10639 (N_10639,N_7686,N_7951);
nor U10640 (N_10640,N_8283,N_7780);
and U10641 (N_10641,N_8878,N_6925);
or U10642 (N_10642,N_6047,N_6806);
and U10643 (N_10643,N_8816,N_6070);
and U10644 (N_10644,N_7847,N_7931);
or U10645 (N_10645,N_7847,N_8326);
nand U10646 (N_10646,N_8697,N_8325);
xor U10647 (N_10647,N_8615,N_7974);
nand U10648 (N_10648,N_6254,N_7402);
nor U10649 (N_10649,N_6983,N_8614);
and U10650 (N_10650,N_7167,N_8070);
and U10651 (N_10651,N_8944,N_8672);
xnor U10652 (N_10652,N_7334,N_8124);
nor U10653 (N_10653,N_8533,N_6457);
or U10654 (N_10654,N_8431,N_8486);
nor U10655 (N_10655,N_7598,N_6648);
or U10656 (N_10656,N_8332,N_6747);
nand U10657 (N_10657,N_7402,N_8476);
or U10658 (N_10658,N_6142,N_6784);
or U10659 (N_10659,N_8384,N_8093);
and U10660 (N_10660,N_8554,N_7023);
and U10661 (N_10661,N_8406,N_8319);
nor U10662 (N_10662,N_7826,N_8801);
nand U10663 (N_10663,N_8873,N_8617);
nor U10664 (N_10664,N_8815,N_8014);
nand U10665 (N_10665,N_8536,N_7757);
or U10666 (N_10666,N_6097,N_6556);
nand U10667 (N_10667,N_8391,N_6671);
or U10668 (N_10668,N_8751,N_7848);
nand U10669 (N_10669,N_6104,N_7004);
or U10670 (N_10670,N_6446,N_6839);
and U10671 (N_10671,N_6480,N_6720);
or U10672 (N_10672,N_6558,N_6085);
and U10673 (N_10673,N_8151,N_8500);
nand U10674 (N_10674,N_6521,N_7291);
or U10675 (N_10675,N_8812,N_7593);
or U10676 (N_10676,N_6030,N_8343);
nor U10677 (N_10677,N_6298,N_6944);
xor U10678 (N_10678,N_6949,N_8900);
nor U10679 (N_10679,N_6593,N_6918);
and U10680 (N_10680,N_6709,N_8202);
and U10681 (N_10681,N_8067,N_8298);
nand U10682 (N_10682,N_7628,N_6141);
and U10683 (N_10683,N_7643,N_8774);
and U10684 (N_10684,N_6242,N_7295);
nand U10685 (N_10685,N_6789,N_6484);
nor U10686 (N_10686,N_7245,N_6272);
and U10687 (N_10687,N_7820,N_8854);
nor U10688 (N_10688,N_6529,N_7361);
nand U10689 (N_10689,N_6837,N_7549);
nor U10690 (N_10690,N_6905,N_8038);
or U10691 (N_10691,N_8358,N_6236);
and U10692 (N_10692,N_7036,N_8968);
and U10693 (N_10693,N_8404,N_6831);
xor U10694 (N_10694,N_7229,N_8078);
and U10695 (N_10695,N_8767,N_7094);
nor U10696 (N_10696,N_6177,N_8061);
nand U10697 (N_10697,N_8097,N_7053);
nand U10698 (N_10698,N_8974,N_8739);
nand U10699 (N_10699,N_8716,N_8319);
and U10700 (N_10700,N_8263,N_7713);
nor U10701 (N_10701,N_6918,N_8704);
nor U10702 (N_10702,N_6151,N_6185);
nor U10703 (N_10703,N_6765,N_8455);
nor U10704 (N_10704,N_7955,N_8552);
and U10705 (N_10705,N_8447,N_7722);
nand U10706 (N_10706,N_8061,N_6451);
or U10707 (N_10707,N_8325,N_6919);
and U10708 (N_10708,N_8347,N_8976);
and U10709 (N_10709,N_7111,N_7358);
and U10710 (N_10710,N_7390,N_6572);
nand U10711 (N_10711,N_7335,N_7383);
and U10712 (N_10712,N_7373,N_7015);
or U10713 (N_10713,N_7124,N_7434);
nand U10714 (N_10714,N_8398,N_8238);
nor U10715 (N_10715,N_7337,N_8684);
or U10716 (N_10716,N_6707,N_7783);
and U10717 (N_10717,N_7251,N_6341);
nor U10718 (N_10718,N_8604,N_7460);
or U10719 (N_10719,N_7280,N_7272);
or U10720 (N_10720,N_6519,N_8902);
nor U10721 (N_10721,N_7056,N_6438);
nor U10722 (N_10722,N_7307,N_8077);
nor U10723 (N_10723,N_8129,N_6137);
nor U10724 (N_10724,N_7022,N_8727);
nor U10725 (N_10725,N_8655,N_7438);
and U10726 (N_10726,N_6420,N_8263);
nor U10727 (N_10727,N_6159,N_8924);
nand U10728 (N_10728,N_6923,N_7349);
nor U10729 (N_10729,N_7705,N_6563);
nand U10730 (N_10730,N_6873,N_7825);
and U10731 (N_10731,N_7182,N_6563);
xor U10732 (N_10732,N_6342,N_7602);
or U10733 (N_10733,N_6188,N_6343);
and U10734 (N_10734,N_6127,N_8799);
nand U10735 (N_10735,N_6417,N_7978);
nor U10736 (N_10736,N_8998,N_6518);
nor U10737 (N_10737,N_6671,N_7798);
nor U10738 (N_10738,N_8766,N_6829);
and U10739 (N_10739,N_7728,N_6456);
nor U10740 (N_10740,N_8764,N_8520);
and U10741 (N_10741,N_6833,N_8994);
nor U10742 (N_10742,N_7624,N_7857);
or U10743 (N_10743,N_6817,N_8150);
or U10744 (N_10744,N_6217,N_6277);
nor U10745 (N_10745,N_7033,N_8545);
and U10746 (N_10746,N_6808,N_6841);
nor U10747 (N_10747,N_7550,N_6002);
or U10748 (N_10748,N_8641,N_7894);
nand U10749 (N_10749,N_6047,N_7331);
nor U10750 (N_10750,N_6290,N_7177);
nor U10751 (N_10751,N_6452,N_8002);
and U10752 (N_10752,N_7828,N_7707);
nand U10753 (N_10753,N_6701,N_8101);
and U10754 (N_10754,N_6731,N_6216);
or U10755 (N_10755,N_8413,N_7927);
and U10756 (N_10756,N_7024,N_7004);
or U10757 (N_10757,N_7848,N_7792);
or U10758 (N_10758,N_8610,N_6286);
nand U10759 (N_10759,N_7605,N_8153);
or U10760 (N_10760,N_6127,N_6915);
or U10761 (N_10761,N_7993,N_8441);
and U10762 (N_10762,N_6526,N_8207);
or U10763 (N_10763,N_8085,N_8721);
or U10764 (N_10764,N_7641,N_7770);
or U10765 (N_10765,N_7396,N_8022);
and U10766 (N_10766,N_6483,N_6421);
nor U10767 (N_10767,N_6849,N_6644);
or U10768 (N_10768,N_7324,N_7447);
or U10769 (N_10769,N_7326,N_8508);
or U10770 (N_10770,N_6252,N_6498);
nor U10771 (N_10771,N_7168,N_6235);
nand U10772 (N_10772,N_7048,N_6727);
nand U10773 (N_10773,N_7423,N_6357);
or U10774 (N_10774,N_7974,N_8043);
and U10775 (N_10775,N_6312,N_8999);
nor U10776 (N_10776,N_7149,N_8389);
and U10777 (N_10777,N_7336,N_7319);
and U10778 (N_10778,N_8238,N_8468);
nor U10779 (N_10779,N_7940,N_6617);
and U10780 (N_10780,N_6322,N_7512);
xnor U10781 (N_10781,N_7642,N_8091);
nand U10782 (N_10782,N_7715,N_6300);
xor U10783 (N_10783,N_7092,N_6260);
nor U10784 (N_10784,N_6677,N_7294);
and U10785 (N_10785,N_7695,N_7343);
and U10786 (N_10786,N_6254,N_6219);
nand U10787 (N_10787,N_7666,N_6737);
nand U10788 (N_10788,N_7547,N_7272);
nand U10789 (N_10789,N_7199,N_6063);
nor U10790 (N_10790,N_8247,N_8921);
and U10791 (N_10791,N_6360,N_7307);
or U10792 (N_10792,N_8950,N_7250);
or U10793 (N_10793,N_7694,N_8264);
or U10794 (N_10794,N_6974,N_6961);
or U10795 (N_10795,N_8442,N_6760);
and U10796 (N_10796,N_7114,N_6154);
and U10797 (N_10797,N_7256,N_7453);
nor U10798 (N_10798,N_6785,N_8038);
or U10799 (N_10799,N_6195,N_6092);
or U10800 (N_10800,N_6436,N_7839);
nand U10801 (N_10801,N_6273,N_6484);
or U10802 (N_10802,N_6849,N_8459);
nand U10803 (N_10803,N_7821,N_6977);
nand U10804 (N_10804,N_6329,N_6995);
or U10805 (N_10805,N_7816,N_7933);
nor U10806 (N_10806,N_8129,N_6902);
or U10807 (N_10807,N_8520,N_6377);
or U10808 (N_10808,N_6475,N_6482);
and U10809 (N_10809,N_6033,N_6153);
or U10810 (N_10810,N_8141,N_6147);
and U10811 (N_10811,N_8335,N_8762);
and U10812 (N_10812,N_7029,N_6780);
or U10813 (N_10813,N_8264,N_8199);
and U10814 (N_10814,N_7459,N_7426);
or U10815 (N_10815,N_8090,N_6001);
nand U10816 (N_10816,N_8317,N_6348);
xor U10817 (N_10817,N_6246,N_8642);
and U10818 (N_10818,N_6737,N_6036);
nand U10819 (N_10819,N_6734,N_7810);
or U10820 (N_10820,N_7213,N_8072);
or U10821 (N_10821,N_6367,N_8710);
nor U10822 (N_10822,N_7747,N_6476);
nor U10823 (N_10823,N_8624,N_8153);
and U10824 (N_10824,N_6024,N_7260);
and U10825 (N_10825,N_8185,N_6772);
and U10826 (N_10826,N_7911,N_7909);
and U10827 (N_10827,N_7715,N_8589);
nor U10828 (N_10828,N_8997,N_6192);
nand U10829 (N_10829,N_8189,N_8906);
or U10830 (N_10830,N_6534,N_8172);
nor U10831 (N_10831,N_6308,N_8344);
and U10832 (N_10832,N_7422,N_8096);
nand U10833 (N_10833,N_7709,N_7073);
and U10834 (N_10834,N_6632,N_8132);
and U10835 (N_10835,N_6802,N_6107);
nand U10836 (N_10836,N_7175,N_7848);
nor U10837 (N_10837,N_8235,N_7450);
nand U10838 (N_10838,N_6627,N_6057);
nor U10839 (N_10839,N_8146,N_7504);
and U10840 (N_10840,N_6187,N_6293);
nor U10841 (N_10841,N_8526,N_7092);
or U10842 (N_10842,N_7082,N_8529);
or U10843 (N_10843,N_7063,N_6600);
or U10844 (N_10844,N_7356,N_6814);
xor U10845 (N_10845,N_7589,N_7328);
nor U10846 (N_10846,N_7133,N_7239);
nand U10847 (N_10847,N_6146,N_7386);
nor U10848 (N_10848,N_7799,N_6529);
and U10849 (N_10849,N_8760,N_6878);
or U10850 (N_10850,N_8498,N_6504);
and U10851 (N_10851,N_6986,N_7619);
and U10852 (N_10852,N_8289,N_8631);
or U10853 (N_10853,N_6357,N_8305);
or U10854 (N_10854,N_8548,N_6054);
nor U10855 (N_10855,N_8390,N_6797);
or U10856 (N_10856,N_6109,N_7855);
and U10857 (N_10857,N_8241,N_7847);
nor U10858 (N_10858,N_8373,N_6047);
or U10859 (N_10859,N_8948,N_8079);
xor U10860 (N_10860,N_6579,N_7256);
nor U10861 (N_10861,N_8421,N_8418);
or U10862 (N_10862,N_6869,N_7458);
nand U10863 (N_10863,N_6215,N_6965);
xnor U10864 (N_10864,N_8865,N_7469);
nand U10865 (N_10865,N_7608,N_8585);
or U10866 (N_10866,N_8790,N_8465);
and U10867 (N_10867,N_6782,N_6410);
or U10868 (N_10868,N_6582,N_6604);
nor U10869 (N_10869,N_6386,N_8648);
and U10870 (N_10870,N_8461,N_8457);
or U10871 (N_10871,N_6593,N_6023);
and U10872 (N_10872,N_7846,N_7436);
and U10873 (N_10873,N_8404,N_8414);
or U10874 (N_10874,N_7496,N_8360);
or U10875 (N_10875,N_8044,N_7641);
nand U10876 (N_10876,N_7869,N_7658);
and U10877 (N_10877,N_7236,N_6653);
and U10878 (N_10878,N_8386,N_7288);
and U10879 (N_10879,N_6730,N_6592);
or U10880 (N_10880,N_8546,N_8311);
nor U10881 (N_10881,N_6326,N_6369);
or U10882 (N_10882,N_8026,N_6696);
nor U10883 (N_10883,N_6077,N_7590);
nor U10884 (N_10884,N_8156,N_7786);
nor U10885 (N_10885,N_8886,N_6709);
nand U10886 (N_10886,N_8108,N_8822);
nor U10887 (N_10887,N_8628,N_8681);
or U10888 (N_10888,N_7886,N_7386);
nand U10889 (N_10889,N_6792,N_6309);
xor U10890 (N_10890,N_7935,N_7575);
nor U10891 (N_10891,N_8676,N_7657);
nand U10892 (N_10892,N_6344,N_6998);
or U10893 (N_10893,N_8974,N_6243);
nor U10894 (N_10894,N_8178,N_6686);
and U10895 (N_10895,N_8518,N_8678);
nor U10896 (N_10896,N_6168,N_7490);
nand U10897 (N_10897,N_8316,N_7698);
nor U10898 (N_10898,N_7388,N_6839);
nor U10899 (N_10899,N_7042,N_7095);
and U10900 (N_10900,N_7816,N_6159);
or U10901 (N_10901,N_6551,N_7160);
nand U10902 (N_10902,N_6965,N_7058);
or U10903 (N_10903,N_8374,N_7044);
or U10904 (N_10904,N_8896,N_8586);
nand U10905 (N_10905,N_7614,N_8842);
nand U10906 (N_10906,N_7048,N_6347);
or U10907 (N_10907,N_7486,N_8681);
nor U10908 (N_10908,N_8853,N_7129);
nand U10909 (N_10909,N_7008,N_6264);
or U10910 (N_10910,N_8983,N_7731);
nor U10911 (N_10911,N_8984,N_8185);
nand U10912 (N_10912,N_7146,N_7425);
nand U10913 (N_10913,N_8743,N_6858);
nand U10914 (N_10914,N_7257,N_8855);
xor U10915 (N_10915,N_6960,N_8437);
xor U10916 (N_10916,N_8595,N_7371);
or U10917 (N_10917,N_8744,N_8456);
nor U10918 (N_10918,N_6058,N_6613);
and U10919 (N_10919,N_7247,N_7178);
or U10920 (N_10920,N_7926,N_8462);
or U10921 (N_10921,N_6684,N_8721);
or U10922 (N_10922,N_7528,N_7452);
and U10923 (N_10923,N_6974,N_8620);
nand U10924 (N_10924,N_7488,N_8077);
nor U10925 (N_10925,N_7191,N_7601);
nand U10926 (N_10926,N_6979,N_7802);
nand U10927 (N_10927,N_8738,N_6781);
nor U10928 (N_10928,N_8755,N_8049);
or U10929 (N_10929,N_6404,N_7697);
or U10930 (N_10930,N_8489,N_6273);
or U10931 (N_10931,N_7438,N_6945);
nor U10932 (N_10932,N_6531,N_6895);
or U10933 (N_10933,N_8855,N_7314);
xor U10934 (N_10934,N_8018,N_7666);
nand U10935 (N_10935,N_8788,N_7129);
nor U10936 (N_10936,N_7592,N_7142);
nor U10937 (N_10937,N_7789,N_7581);
nand U10938 (N_10938,N_8021,N_8318);
or U10939 (N_10939,N_8889,N_7668);
and U10940 (N_10940,N_6093,N_8517);
and U10941 (N_10941,N_8137,N_6846);
xor U10942 (N_10942,N_8251,N_6567);
nor U10943 (N_10943,N_6723,N_6980);
and U10944 (N_10944,N_8797,N_8682);
and U10945 (N_10945,N_7675,N_8275);
and U10946 (N_10946,N_8867,N_6855);
and U10947 (N_10947,N_6081,N_8648);
nor U10948 (N_10948,N_6134,N_7938);
xnor U10949 (N_10949,N_8362,N_7911);
and U10950 (N_10950,N_7534,N_7029);
xnor U10951 (N_10951,N_7471,N_7976);
and U10952 (N_10952,N_6423,N_7645);
and U10953 (N_10953,N_7476,N_6619);
nor U10954 (N_10954,N_6984,N_7843);
or U10955 (N_10955,N_7320,N_8752);
nor U10956 (N_10956,N_8890,N_8638);
or U10957 (N_10957,N_7338,N_7223);
nor U10958 (N_10958,N_6680,N_6228);
nor U10959 (N_10959,N_8692,N_7456);
or U10960 (N_10960,N_8240,N_8254);
nor U10961 (N_10961,N_8138,N_7320);
and U10962 (N_10962,N_6831,N_8704);
or U10963 (N_10963,N_7902,N_6906);
or U10964 (N_10964,N_6327,N_7965);
or U10965 (N_10965,N_6791,N_8853);
xnor U10966 (N_10966,N_8198,N_8116);
nor U10967 (N_10967,N_6232,N_6795);
or U10968 (N_10968,N_6633,N_8200);
nor U10969 (N_10969,N_6608,N_7632);
xor U10970 (N_10970,N_8943,N_6881);
and U10971 (N_10971,N_7662,N_6458);
or U10972 (N_10972,N_8116,N_8239);
nand U10973 (N_10973,N_6144,N_8773);
and U10974 (N_10974,N_6186,N_7772);
nor U10975 (N_10975,N_6359,N_7012);
or U10976 (N_10976,N_6170,N_8463);
nand U10977 (N_10977,N_8010,N_8662);
nand U10978 (N_10978,N_8863,N_6418);
or U10979 (N_10979,N_8386,N_7112);
or U10980 (N_10980,N_7785,N_6003);
or U10981 (N_10981,N_8303,N_6248);
nand U10982 (N_10982,N_8263,N_7896);
nor U10983 (N_10983,N_7909,N_7055);
nand U10984 (N_10984,N_8968,N_7349);
nor U10985 (N_10985,N_6381,N_6866);
nor U10986 (N_10986,N_8295,N_7202);
and U10987 (N_10987,N_6542,N_6901);
nand U10988 (N_10988,N_8211,N_6995);
or U10989 (N_10989,N_7920,N_6879);
and U10990 (N_10990,N_7871,N_8702);
nand U10991 (N_10991,N_8578,N_8101);
nand U10992 (N_10992,N_8425,N_6943);
and U10993 (N_10993,N_6853,N_6516);
nor U10994 (N_10994,N_7807,N_8174);
and U10995 (N_10995,N_8109,N_7516);
nand U10996 (N_10996,N_6974,N_8701);
or U10997 (N_10997,N_7712,N_7949);
nand U10998 (N_10998,N_7791,N_7493);
or U10999 (N_10999,N_7635,N_8423);
nor U11000 (N_11000,N_7435,N_6484);
and U11001 (N_11001,N_6001,N_6696);
nor U11002 (N_11002,N_6629,N_6390);
or U11003 (N_11003,N_8627,N_6223);
nand U11004 (N_11004,N_6146,N_6088);
or U11005 (N_11005,N_6405,N_7682);
nor U11006 (N_11006,N_6827,N_8717);
nand U11007 (N_11007,N_7552,N_8361);
and U11008 (N_11008,N_8392,N_6575);
or U11009 (N_11009,N_6300,N_6693);
nor U11010 (N_11010,N_6013,N_8995);
and U11011 (N_11011,N_6153,N_8349);
nand U11012 (N_11012,N_7598,N_6774);
nand U11013 (N_11013,N_8984,N_8197);
or U11014 (N_11014,N_6399,N_7316);
or U11015 (N_11015,N_8007,N_7925);
nand U11016 (N_11016,N_7038,N_7382);
nand U11017 (N_11017,N_8296,N_8753);
nor U11018 (N_11018,N_6028,N_8041);
and U11019 (N_11019,N_6554,N_8909);
and U11020 (N_11020,N_7155,N_8445);
or U11021 (N_11021,N_7769,N_6760);
or U11022 (N_11022,N_7451,N_8189);
and U11023 (N_11023,N_6083,N_6680);
and U11024 (N_11024,N_7792,N_8550);
xor U11025 (N_11025,N_7876,N_7680);
and U11026 (N_11026,N_8338,N_8184);
nand U11027 (N_11027,N_6504,N_8405);
nand U11028 (N_11028,N_7973,N_6418);
and U11029 (N_11029,N_8382,N_6539);
nor U11030 (N_11030,N_8357,N_7582);
nand U11031 (N_11031,N_7166,N_7319);
and U11032 (N_11032,N_7388,N_7400);
and U11033 (N_11033,N_6288,N_6704);
xor U11034 (N_11034,N_6724,N_8843);
or U11035 (N_11035,N_6944,N_7356);
nor U11036 (N_11036,N_8596,N_6178);
and U11037 (N_11037,N_6321,N_7238);
nand U11038 (N_11038,N_8971,N_6242);
or U11039 (N_11039,N_6395,N_6433);
nand U11040 (N_11040,N_6340,N_8828);
or U11041 (N_11041,N_8632,N_6570);
or U11042 (N_11042,N_6162,N_8038);
nor U11043 (N_11043,N_8354,N_8456);
and U11044 (N_11044,N_7292,N_8356);
nand U11045 (N_11045,N_6285,N_7231);
nor U11046 (N_11046,N_8082,N_8694);
and U11047 (N_11047,N_6482,N_6204);
nand U11048 (N_11048,N_8680,N_7899);
nor U11049 (N_11049,N_7953,N_7060);
or U11050 (N_11050,N_8420,N_8343);
or U11051 (N_11051,N_7992,N_8312);
nor U11052 (N_11052,N_8195,N_7102);
or U11053 (N_11053,N_6395,N_8651);
nand U11054 (N_11054,N_8142,N_8012);
or U11055 (N_11055,N_6572,N_6507);
nor U11056 (N_11056,N_7479,N_7689);
nor U11057 (N_11057,N_7475,N_7675);
nor U11058 (N_11058,N_8793,N_6118);
nor U11059 (N_11059,N_8832,N_7068);
nand U11060 (N_11060,N_7382,N_7976);
nand U11061 (N_11061,N_7687,N_7928);
nand U11062 (N_11062,N_8147,N_6409);
or U11063 (N_11063,N_6388,N_8456);
and U11064 (N_11064,N_7473,N_7016);
and U11065 (N_11065,N_6780,N_6919);
nand U11066 (N_11066,N_6896,N_7400);
nand U11067 (N_11067,N_8234,N_7023);
or U11068 (N_11068,N_8057,N_6140);
or U11069 (N_11069,N_7402,N_8518);
or U11070 (N_11070,N_8276,N_7625);
nand U11071 (N_11071,N_7512,N_7669);
and U11072 (N_11072,N_8821,N_8157);
and U11073 (N_11073,N_6033,N_7944);
nor U11074 (N_11074,N_8464,N_6009);
nand U11075 (N_11075,N_6297,N_8735);
and U11076 (N_11076,N_6838,N_8961);
or U11077 (N_11077,N_7781,N_6794);
and U11078 (N_11078,N_8494,N_6922);
or U11079 (N_11079,N_7088,N_8710);
nand U11080 (N_11080,N_7543,N_7634);
nand U11081 (N_11081,N_6081,N_6042);
or U11082 (N_11082,N_8230,N_6941);
nand U11083 (N_11083,N_8699,N_8933);
and U11084 (N_11084,N_6570,N_7827);
and U11085 (N_11085,N_6743,N_8300);
and U11086 (N_11086,N_6193,N_6187);
and U11087 (N_11087,N_7338,N_8790);
xor U11088 (N_11088,N_6165,N_7668);
nand U11089 (N_11089,N_7052,N_8852);
and U11090 (N_11090,N_8242,N_7777);
nand U11091 (N_11091,N_6345,N_7543);
nand U11092 (N_11092,N_8368,N_8445);
or U11093 (N_11093,N_7813,N_6230);
and U11094 (N_11094,N_7195,N_6794);
nand U11095 (N_11095,N_8303,N_6665);
nor U11096 (N_11096,N_8362,N_6590);
xnor U11097 (N_11097,N_8751,N_7025);
or U11098 (N_11098,N_8491,N_7921);
nor U11099 (N_11099,N_8837,N_7337);
nand U11100 (N_11100,N_8185,N_7027);
nor U11101 (N_11101,N_7873,N_6868);
nor U11102 (N_11102,N_7952,N_7317);
nand U11103 (N_11103,N_6269,N_7441);
or U11104 (N_11104,N_6383,N_8494);
and U11105 (N_11105,N_6800,N_7219);
nor U11106 (N_11106,N_6580,N_7006);
or U11107 (N_11107,N_8340,N_6481);
and U11108 (N_11108,N_7304,N_7886);
nand U11109 (N_11109,N_6096,N_7090);
or U11110 (N_11110,N_8816,N_8496);
and U11111 (N_11111,N_7122,N_8943);
nand U11112 (N_11112,N_8927,N_7231);
nor U11113 (N_11113,N_7208,N_6047);
nor U11114 (N_11114,N_7915,N_6793);
nor U11115 (N_11115,N_8184,N_6913);
or U11116 (N_11116,N_8619,N_7053);
and U11117 (N_11117,N_6514,N_8189);
nand U11118 (N_11118,N_6727,N_7495);
and U11119 (N_11119,N_8677,N_6262);
nand U11120 (N_11120,N_8750,N_7905);
or U11121 (N_11121,N_7921,N_8703);
xor U11122 (N_11122,N_7253,N_8954);
and U11123 (N_11123,N_8991,N_6442);
or U11124 (N_11124,N_6416,N_7063);
nor U11125 (N_11125,N_8769,N_6232);
or U11126 (N_11126,N_7495,N_7071);
nor U11127 (N_11127,N_7109,N_6059);
nand U11128 (N_11128,N_8663,N_7778);
nor U11129 (N_11129,N_8519,N_7549);
or U11130 (N_11130,N_8028,N_7560);
nor U11131 (N_11131,N_6390,N_6162);
and U11132 (N_11132,N_6520,N_7970);
xor U11133 (N_11133,N_7561,N_6270);
and U11134 (N_11134,N_8331,N_6971);
nand U11135 (N_11135,N_7861,N_7783);
or U11136 (N_11136,N_6505,N_6870);
xnor U11137 (N_11137,N_7356,N_8808);
or U11138 (N_11138,N_8089,N_7348);
or U11139 (N_11139,N_7430,N_8302);
nor U11140 (N_11140,N_8725,N_7414);
nor U11141 (N_11141,N_7867,N_6239);
nand U11142 (N_11142,N_6970,N_8778);
nand U11143 (N_11143,N_6033,N_6734);
nand U11144 (N_11144,N_6967,N_8268);
and U11145 (N_11145,N_6659,N_8286);
or U11146 (N_11146,N_8188,N_6383);
and U11147 (N_11147,N_8636,N_6187);
and U11148 (N_11148,N_8682,N_8469);
nor U11149 (N_11149,N_7485,N_6587);
or U11150 (N_11150,N_6598,N_8106);
nor U11151 (N_11151,N_7047,N_7544);
or U11152 (N_11152,N_6361,N_8953);
and U11153 (N_11153,N_7052,N_7611);
nor U11154 (N_11154,N_6887,N_7076);
or U11155 (N_11155,N_8394,N_8664);
nor U11156 (N_11156,N_6211,N_6997);
nand U11157 (N_11157,N_6255,N_8356);
or U11158 (N_11158,N_8241,N_7857);
nor U11159 (N_11159,N_8791,N_6217);
nand U11160 (N_11160,N_6203,N_7531);
nor U11161 (N_11161,N_6889,N_6045);
nor U11162 (N_11162,N_8785,N_8839);
or U11163 (N_11163,N_7213,N_7423);
and U11164 (N_11164,N_6254,N_8415);
nand U11165 (N_11165,N_7608,N_7614);
and U11166 (N_11166,N_7762,N_8065);
and U11167 (N_11167,N_8367,N_6164);
nand U11168 (N_11168,N_7602,N_6283);
nor U11169 (N_11169,N_7674,N_6193);
nor U11170 (N_11170,N_6147,N_8626);
nand U11171 (N_11171,N_7288,N_7032);
or U11172 (N_11172,N_8886,N_7403);
and U11173 (N_11173,N_7629,N_7367);
and U11174 (N_11174,N_6132,N_6992);
nand U11175 (N_11175,N_7502,N_8688);
nor U11176 (N_11176,N_7209,N_8100);
nor U11177 (N_11177,N_7411,N_8087);
or U11178 (N_11178,N_8215,N_7267);
or U11179 (N_11179,N_8563,N_6239);
or U11180 (N_11180,N_7425,N_8960);
and U11181 (N_11181,N_6119,N_7849);
nor U11182 (N_11182,N_6432,N_8368);
nand U11183 (N_11183,N_7934,N_8193);
or U11184 (N_11184,N_6196,N_6123);
nor U11185 (N_11185,N_8202,N_7042);
and U11186 (N_11186,N_7372,N_6536);
nand U11187 (N_11187,N_8238,N_8196);
or U11188 (N_11188,N_8659,N_8641);
nand U11189 (N_11189,N_7085,N_7972);
xor U11190 (N_11190,N_6611,N_6244);
nor U11191 (N_11191,N_8603,N_6792);
or U11192 (N_11192,N_7056,N_8931);
and U11193 (N_11193,N_6051,N_8603);
or U11194 (N_11194,N_7719,N_7032);
and U11195 (N_11195,N_8171,N_6355);
nor U11196 (N_11196,N_7962,N_7958);
or U11197 (N_11197,N_6359,N_7287);
nor U11198 (N_11198,N_7195,N_7579);
nand U11199 (N_11199,N_8101,N_8251);
nor U11200 (N_11200,N_6243,N_7539);
nand U11201 (N_11201,N_6623,N_6738);
nand U11202 (N_11202,N_7199,N_8854);
or U11203 (N_11203,N_7613,N_8338);
or U11204 (N_11204,N_7946,N_8050);
nor U11205 (N_11205,N_6884,N_7628);
xnor U11206 (N_11206,N_6040,N_6414);
and U11207 (N_11207,N_8961,N_6380);
or U11208 (N_11208,N_8631,N_7523);
and U11209 (N_11209,N_7306,N_7323);
nor U11210 (N_11210,N_8656,N_8227);
nand U11211 (N_11211,N_7986,N_7480);
nand U11212 (N_11212,N_6091,N_8794);
or U11213 (N_11213,N_8183,N_6805);
nor U11214 (N_11214,N_8253,N_6822);
nand U11215 (N_11215,N_6493,N_6151);
nor U11216 (N_11216,N_6839,N_8648);
nand U11217 (N_11217,N_6577,N_7939);
and U11218 (N_11218,N_6035,N_6871);
and U11219 (N_11219,N_8701,N_6524);
and U11220 (N_11220,N_8957,N_6307);
nand U11221 (N_11221,N_6949,N_6557);
nand U11222 (N_11222,N_7472,N_7540);
nor U11223 (N_11223,N_6057,N_6302);
nand U11224 (N_11224,N_8456,N_8844);
nor U11225 (N_11225,N_6232,N_6161);
nand U11226 (N_11226,N_7873,N_7068);
and U11227 (N_11227,N_7388,N_6696);
nand U11228 (N_11228,N_6339,N_6822);
and U11229 (N_11229,N_6128,N_8917);
or U11230 (N_11230,N_6266,N_7982);
and U11231 (N_11231,N_6328,N_7413);
nand U11232 (N_11232,N_7427,N_8163);
and U11233 (N_11233,N_8725,N_7859);
or U11234 (N_11234,N_7578,N_8224);
or U11235 (N_11235,N_6462,N_8238);
nor U11236 (N_11236,N_8190,N_6488);
nand U11237 (N_11237,N_8622,N_6089);
nand U11238 (N_11238,N_8057,N_6010);
nand U11239 (N_11239,N_6455,N_8301);
nand U11240 (N_11240,N_7506,N_6951);
xnor U11241 (N_11241,N_6679,N_6566);
nand U11242 (N_11242,N_6201,N_7839);
nand U11243 (N_11243,N_8865,N_7875);
and U11244 (N_11244,N_6472,N_7330);
nand U11245 (N_11245,N_6792,N_8179);
nor U11246 (N_11246,N_6968,N_8472);
or U11247 (N_11247,N_8638,N_6650);
nor U11248 (N_11248,N_8560,N_6155);
nor U11249 (N_11249,N_8245,N_6023);
or U11250 (N_11250,N_8553,N_7953);
nor U11251 (N_11251,N_8843,N_8479);
nor U11252 (N_11252,N_7278,N_7966);
and U11253 (N_11253,N_8846,N_7378);
nor U11254 (N_11254,N_8738,N_7393);
and U11255 (N_11255,N_7359,N_8879);
or U11256 (N_11256,N_8882,N_8756);
nand U11257 (N_11257,N_6448,N_7201);
nor U11258 (N_11258,N_7122,N_8271);
nand U11259 (N_11259,N_6472,N_7621);
nand U11260 (N_11260,N_6036,N_8000);
nor U11261 (N_11261,N_7835,N_8450);
nand U11262 (N_11262,N_7819,N_7615);
or U11263 (N_11263,N_7219,N_7555);
nor U11264 (N_11264,N_7992,N_8231);
or U11265 (N_11265,N_8428,N_8441);
nor U11266 (N_11266,N_8883,N_6361);
nor U11267 (N_11267,N_7672,N_8250);
nand U11268 (N_11268,N_6175,N_7839);
nor U11269 (N_11269,N_8442,N_6529);
nor U11270 (N_11270,N_8790,N_8961);
or U11271 (N_11271,N_6137,N_8904);
nor U11272 (N_11272,N_6886,N_7046);
nand U11273 (N_11273,N_6377,N_6015);
or U11274 (N_11274,N_8956,N_7107);
nand U11275 (N_11275,N_7751,N_7245);
or U11276 (N_11276,N_8322,N_8467);
and U11277 (N_11277,N_7448,N_6865);
nand U11278 (N_11278,N_8440,N_6519);
and U11279 (N_11279,N_8847,N_6258);
nand U11280 (N_11280,N_6147,N_7301);
and U11281 (N_11281,N_6950,N_6288);
or U11282 (N_11282,N_8988,N_8437);
or U11283 (N_11283,N_6277,N_8740);
or U11284 (N_11284,N_8030,N_7015);
or U11285 (N_11285,N_7672,N_7054);
nand U11286 (N_11286,N_6409,N_7791);
xnor U11287 (N_11287,N_8136,N_7830);
nor U11288 (N_11288,N_6934,N_6085);
nand U11289 (N_11289,N_6902,N_8539);
or U11290 (N_11290,N_8193,N_6676);
or U11291 (N_11291,N_7975,N_7585);
xor U11292 (N_11292,N_8679,N_7784);
or U11293 (N_11293,N_7242,N_8623);
nor U11294 (N_11294,N_6575,N_7976);
nor U11295 (N_11295,N_6507,N_7889);
or U11296 (N_11296,N_8192,N_8049);
nand U11297 (N_11297,N_8843,N_6239);
nor U11298 (N_11298,N_6215,N_8457);
nor U11299 (N_11299,N_7665,N_8078);
or U11300 (N_11300,N_7801,N_8337);
and U11301 (N_11301,N_8382,N_6184);
and U11302 (N_11302,N_7353,N_8524);
nor U11303 (N_11303,N_8806,N_6846);
nand U11304 (N_11304,N_8184,N_8030);
or U11305 (N_11305,N_6879,N_7390);
nand U11306 (N_11306,N_7110,N_6474);
xor U11307 (N_11307,N_8388,N_6656);
or U11308 (N_11308,N_8975,N_7182);
nand U11309 (N_11309,N_6796,N_8019);
or U11310 (N_11310,N_7642,N_8028);
nor U11311 (N_11311,N_6894,N_8497);
and U11312 (N_11312,N_7145,N_7167);
and U11313 (N_11313,N_6997,N_8481);
nor U11314 (N_11314,N_8486,N_7456);
nand U11315 (N_11315,N_8822,N_6842);
nor U11316 (N_11316,N_8301,N_7060);
nand U11317 (N_11317,N_8174,N_6293);
nand U11318 (N_11318,N_7132,N_8824);
nor U11319 (N_11319,N_7617,N_7860);
or U11320 (N_11320,N_8183,N_8115);
nor U11321 (N_11321,N_6231,N_8540);
or U11322 (N_11322,N_7060,N_7820);
and U11323 (N_11323,N_8603,N_6271);
or U11324 (N_11324,N_6524,N_7619);
xnor U11325 (N_11325,N_8084,N_7067);
and U11326 (N_11326,N_8375,N_7466);
and U11327 (N_11327,N_6304,N_7512);
nor U11328 (N_11328,N_7712,N_7332);
nor U11329 (N_11329,N_7624,N_6837);
and U11330 (N_11330,N_8763,N_6369);
nor U11331 (N_11331,N_6516,N_7717);
nor U11332 (N_11332,N_7863,N_6714);
nor U11333 (N_11333,N_7110,N_8318);
or U11334 (N_11334,N_7841,N_7574);
and U11335 (N_11335,N_7412,N_8417);
and U11336 (N_11336,N_7165,N_7769);
nor U11337 (N_11337,N_8968,N_7940);
and U11338 (N_11338,N_7130,N_6605);
nand U11339 (N_11339,N_7324,N_6764);
and U11340 (N_11340,N_8359,N_7141);
or U11341 (N_11341,N_6484,N_8508);
nor U11342 (N_11342,N_8791,N_6853);
nand U11343 (N_11343,N_6645,N_6025);
or U11344 (N_11344,N_7311,N_8747);
xnor U11345 (N_11345,N_6966,N_8868);
and U11346 (N_11346,N_8579,N_7361);
nor U11347 (N_11347,N_6118,N_6836);
nor U11348 (N_11348,N_8996,N_6242);
or U11349 (N_11349,N_7157,N_6934);
or U11350 (N_11350,N_6646,N_8694);
or U11351 (N_11351,N_6871,N_7693);
xnor U11352 (N_11352,N_6251,N_6744);
and U11353 (N_11353,N_7571,N_6607);
and U11354 (N_11354,N_7891,N_8358);
nor U11355 (N_11355,N_8612,N_8757);
and U11356 (N_11356,N_6386,N_7297);
and U11357 (N_11357,N_7382,N_6422);
nand U11358 (N_11358,N_7661,N_6323);
and U11359 (N_11359,N_6004,N_6140);
nor U11360 (N_11360,N_6304,N_6329);
xnor U11361 (N_11361,N_6931,N_8094);
nor U11362 (N_11362,N_8775,N_7136);
and U11363 (N_11363,N_8270,N_6436);
nor U11364 (N_11364,N_6042,N_7849);
and U11365 (N_11365,N_6371,N_7568);
or U11366 (N_11366,N_8381,N_7606);
nand U11367 (N_11367,N_8437,N_8771);
or U11368 (N_11368,N_8000,N_7320);
or U11369 (N_11369,N_8894,N_7566);
or U11370 (N_11370,N_8760,N_6456);
or U11371 (N_11371,N_7682,N_8957);
nor U11372 (N_11372,N_7348,N_8127);
nor U11373 (N_11373,N_7889,N_6159);
nand U11374 (N_11374,N_7038,N_8331);
nand U11375 (N_11375,N_6702,N_7877);
nor U11376 (N_11376,N_6936,N_8004);
nand U11377 (N_11377,N_7062,N_7624);
or U11378 (N_11378,N_8912,N_7615);
nand U11379 (N_11379,N_7872,N_8451);
or U11380 (N_11380,N_8929,N_7248);
nor U11381 (N_11381,N_8410,N_7240);
nand U11382 (N_11382,N_6047,N_6736);
and U11383 (N_11383,N_6373,N_8545);
nand U11384 (N_11384,N_8247,N_8071);
or U11385 (N_11385,N_8980,N_8160);
nor U11386 (N_11386,N_6482,N_7760);
nand U11387 (N_11387,N_7474,N_7887);
nor U11388 (N_11388,N_8138,N_6841);
nand U11389 (N_11389,N_6867,N_6049);
nor U11390 (N_11390,N_7532,N_6649);
or U11391 (N_11391,N_6228,N_8887);
and U11392 (N_11392,N_7195,N_6107);
nor U11393 (N_11393,N_7155,N_8474);
nand U11394 (N_11394,N_6758,N_6900);
and U11395 (N_11395,N_7104,N_7726);
xnor U11396 (N_11396,N_8986,N_8392);
nand U11397 (N_11397,N_6699,N_8207);
and U11398 (N_11398,N_6236,N_6961);
and U11399 (N_11399,N_8559,N_6591);
or U11400 (N_11400,N_6715,N_6367);
nor U11401 (N_11401,N_6680,N_7404);
nand U11402 (N_11402,N_6089,N_6290);
nor U11403 (N_11403,N_7413,N_8084);
nor U11404 (N_11404,N_7748,N_7918);
nor U11405 (N_11405,N_7001,N_6050);
or U11406 (N_11406,N_7348,N_7088);
nor U11407 (N_11407,N_8981,N_7175);
and U11408 (N_11408,N_7310,N_8544);
nand U11409 (N_11409,N_6005,N_8190);
nor U11410 (N_11410,N_7580,N_7431);
or U11411 (N_11411,N_6703,N_6204);
nor U11412 (N_11412,N_6297,N_6821);
or U11413 (N_11413,N_7902,N_8755);
nor U11414 (N_11414,N_7369,N_8668);
and U11415 (N_11415,N_6862,N_8628);
nor U11416 (N_11416,N_6395,N_8390);
and U11417 (N_11417,N_6350,N_6230);
xnor U11418 (N_11418,N_8423,N_8152);
nand U11419 (N_11419,N_8634,N_6875);
and U11420 (N_11420,N_8681,N_7459);
nor U11421 (N_11421,N_7581,N_8289);
nor U11422 (N_11422,N_8738,N_8806);
xor U11423 (N_11423,N_8215,N_8922);
or U11424 (N_11424,N_8552,N_8343);
xor U11425 (N_11425,N_7457,N_7363);
nor U11426 (N_11426,N_8691,N_6852);
nor U11427 (N_11427,N_8026,N_8225);
or U11428 (N_11428,N_8842,N_6395);
or U11429 (N_11429,N_7408,N_8979);
and U11430 (N_11430,N_7284,N_7591);
nor U11431 (N_11431,N_7918,N_6659);
nor U11432 (N_11432,N_7706,N_7846);
nor U11433 (N_11433,N_8896,N_7888);
nor U11434 (N_11434,N_8715,N_6544);
nor U11435 (N_11435,N_6917,N_8351);
nor U11436 (N_11436,N_6707,N_7721);
and U11437 (N_11437,N_8176,N_6011);
nand U11438 (N_11438,N_6432,N_6717);
nand U11439 (N_11439,N_6616,N_8291);
nand U11440 (N_11440,N_8993,N_6897);
nor U11441 (N_11441,N_6158,N_8773);
or U11442 (N_11442,N_6722,N_8374);
nand U11443 (N_11443,N_8109,N_8541);
nand U11444 (N_11444,N_8106,N_7811);
and U11445 (N_11445,N_6459,N_8585);
nand U11446 (N_11446,N_8254,N_6321);
nand U11447 (N_11447,N_8629,N_6301);
nor U11448 (N_11448,N_6772,N_6695);
or U11449 (N_11449,N_6912,N_6896);
or U11450 (N_11450,N_8219,N_6686);
and U11451 (N_11451,N_8483,N_6970);
or U11452 (N_11452,N_6896,N_8925);
nand U11453 (N_11453,N_6803,N_8294);
or U11454 (N_11454,N_7139,N_8125);
and U11455 (N_11455,N_6787,N_6488);
and U11456 (N_11456,N_8106,N_7848);
nand U11457 (N_11457,N_7066,N_8806);
or U11458 (N_11458,N_6026,N_7379);
and U11459 (N_11459,N_7621,N_8036);
and U11460 (N_11460,N_7546,N_6393);
or U11461 (N_11461,N_7481,N_6253);
nor U11462 (N_11462,N_8123,N_8311);
or U11463 (N_11463,N_6517,N_7035);
and U11464 (N_11464,N_8274,N_7688);
nand U11465 (N_11465,N_7881,N_8776);
or U11466 (N_11466,N_8608,N_7508);
nand U11467 (N_11467,N_8569,N_8538);
nor U11468 (N_11468,N_8496,N_6256);
nor U11469 (N_11469,N_8630,N_8940);
nand U11470 (N_11470,N_6085,N_7416);
or U11471 (N_11471,N_7707,N_6140);
and U11472 (N_11472,N_7919,N_8320);
or U11473 (N_11473,N_8972,N_8732);
nor U11474 (N_11474,N_8290,N_8798);
and U11475 (N_11475,N_8195,N_8222);
nand U11476 (N_11476,N_7680,N_7985);
or U11477 (N_11477,N_6294,N_7808);
or U11478 (N_11478,N_8225,N_7592);
and U11479 (N_11479,N_8974,N_6829);
nor U11480 (N_11480,N_6193,N_8277);
nor U11481 (N_11481,N_6329,N_7111);
or U11482 (N_11482,N_6141,N_8173);
nand U11483 (N_11483,N_8058,N_8894);
nor U11484 (N_11484,N_6783,N_6594);
nor U11485 (N_11485,N_7948,N_7232);
or U11486 (N_11486,N_8437,N_6851);
nand U11487 (N_11487,N_8754,N_6976);
or U11488 (N_11488,N_7555,N_6858);
nor U11489 (N_11489,N_6019,N_6330);
nor U11490 (N_11490,N_7710,N_8400);
nor U11491 (N_11491,N_8784,N_7689);
nor U11492 (N_11492,N_8386,N_8888);
nand U11493 (N_11493,N_6520,N_7318);
and U11494 (N_11494,N_8249,N_8657);
nand U11495 (N_11495,N_7501,N_7498);
nor U11496 (N_11496,N_6465,N_7293);
nor U11497 (N_11497,N_6699,N_6371);
nand U11498 (N_11498,N_6565,N_7695);
nor U11499 (N_11499,N_7736,N_7764);
and U11500 (N_11500,N_6181,N_8643);
or U11501 (N_11501,N_6298,N_7546);
or U11502 (N_11502,N_7026,N_8786);
nor U11503 (N_11503,N_8857,N_8334);
nand U11504 (N_11504,N_7219,N_6074);
xnor U11505 (N_11505,N_8657,N_7390);
nor U11506 (N_11506,N_6376,N_8599);
and U11507 (N_11507,N_8867,N_8339);
or U11508 (N_11508,N_6742,N_7317);
or U11509 (N_11509,N_8799,N_7100);
and U11510 (N_11510,N_6158,N_6666);
and U11511 (N_11511,N_7742,N_8523);
or U11512 (N_11512,N_8641,N_7594);
and U11513 (N_11513,N_6804,N_8958);
and U11514 (N_11514,N_8214,N_8201);
nor U11515 (N_11515,N_8521,N_8109);
and U11516 (N_11516,N_6506,N_6618);
nand U11517 (N_11517,N_6152,N_7079);
or U11518 (N_11518,N_6879,N_6230);
and U11519 (N_11519,N_7726,N_6029);
xor U11520 (N_11520,N_6295,N_8040);
nand U11521 (N_11521,N_8837,N_7450);
nor U11522 (N_11522,N_6980,N_6546);
and U11523 (N_11523,N_8963,N_8590);
nor U11524 (N_11524,N_6120,N_8022);
nand U11525 (N_11525,N_8800,N_7444);
and U11526 (N_11526,N_7337,N_8053);
nand U11527 (N_11527,N_7487,N_6121);
or U11528 (N_11528,N_8958,N_6059);
and U11529 (N_11529,N_7357,N_7490);
and U11530 (N_11530,N_8756,N_7144);
nor U11531 (N_11531,N_7377,N_7148);
nand U11532 (N_11532,N_6282,N_8556);
and U11533 (N_11533,N_6176,N_7891);
and U11534 (N_11534,N_6950,N_8921);
and U11535 (N_11535,N_7157,N_8027);
nor U11536 (N_11536,N_7153,N_8965);
nor U11537 (N_11537,N_7617,N_8844);
nor U11538 (N_11538,N_7351,N_8139);
and U11539 (N_11539,N_8123,N_7315);
nand U11540 (N_11540,N_8639,N_6290);
nor U11541 (N_11541,N_6778,N_7581);
or U11542 (N_11542,N_6797,N_6701);
and U11543 (N_11543,N_7051,N_6393);
nor U11544 (N_11544,N_6266,N_6377);
or U11545 (N_11545,N_7915,N_8206);
nand U11546 (N_11546,N_7062,N_7712);
and U11547 (N_11547,N_8024,N_8035);
or U11548 (N_11548,N_6413,N_7898);
nand U11549 (N_11549,N_8667,N_8270);
nand U11550 (N_11550,N_7052,N_6210);
xor U11551 (N_11551,N_6530,N_6268);
and U11552 (N_11552,N_7646,N_6662);
or U11553 (N_11553,N_7068,N_6433);
nand U11554 (N_11554,N_7021,N_6589);
nor U11555 (N_11555,N_6278,N_8593);
or U11556 (N_11556,N_8024,N_7404);
and U11557 (N_11557,N_7114,N_6831);
nand U11558 (N_11558,N_8828,N_8800);
nand U11559 (N_11559,N_7979,N_7715);
or U11560 (N_11560,N_6033,N_8270);
nor U11561 (N_11561,N_6518,N_6901);
nor U11562 (N_11562,N_7926,N_6719);
and U11563 (N_11563,N_6538,N_6522);
nand U11564 (N_11564,N_8152,N_7240);
or U11565 (N_11565,N_7310,N_7133);
or U11566 (N_11566,N_7497,N_8903);
nand U11567 (N_11567,N_6400,N_6525);
nor U11568 (N_11568,N_6510,N_7512);
nor U11569 (N_11569,N_6909,N_7177);
nand U11570 (N_11570,N_6657,N_6140);
or U11571 (N_11571,N_7202,N_6453);
nand U11572 (N_11572,N_7575,N_7495);
or U11573 (N_11573,N_6414,N_7971);
nand U11574 (N_11574,N_8945,N_6377);
or U11575 (N_11575,N_7614,N_6462);
nand U11576 (N_11576,N_6976,N_6210);
and U11577 (N_11577,N_8849,N_7125);
xnor U11578 (N_11578,N_6573,N_7666);
nand U11579 (N_11579,N_6144,N_6098);
or U11580 (N_11580,N_6757,N_6649);
or U11581 (N_11581,N_6049,N_8687);
xor U11582 (N_11582,N_6250,N_7664);
and U11583 (N_11583,N_6785,N_7736);
and U11584 (N_11584,N_8289,N_8698);
or U11585 (N_11585,N_6600,N_8805);
nor U11586 (N_11586,N_8094,N_7667);
nand U11587 (N_11587,N_8943,N_6667);
nand U11588 (N_11588,N_8186,N_8463);
nor U11589 (N_11589,N_7989,N_7928);
or U11590 (N_11590,N_8006,N_6191);
or U11591 (N_11591,N_8979,N_7834);
or U11592 (N_11592,N_7060,N_6990);
and U11593 (N_11593,N_8044,N_8080);
and U11594 (N_11594,N_7813,N_6458);
and U11595 (N_11595,N_8998,N_7168);
or U11596 (N_11596,N_7033,N_8126);
and U11597 (N_11597,N_8675,N_8330);
and U11598 (N_11598,N_8231,N_7327);
and U11599 (N_11599,N_8054,N_7041);
nor U11600 (N_11600,N_7850,N_6449);
nor U11601 (N_11601,N_8413,N_8322);
and U11602 (N_11602,N_6752,N_8587);
nor U11603 (N_11603,N_6862,N_7933);
and U11604 (N_11604,N_6239,N_6192);
and U11605 (N_11605,N_7749,N_6253);
nor U11606 (N_11606,N_6509,N_7306);
and U11607 (N_11607,N_8932,N_8377);
nor U11608 (N_11608,N_8017,N_6432);
nor U11609 (N_11609,N_8911,N_7507);
nor U11610 (N_11610,N_7559,N_7093);
and U11611 (N_11611,N_8172,N_8632);
and U11612 (N_11612,N_8935,N_7768);
and U11613 (N_11613,N_7324,N_8563);
and U11614 (N_11614,N_7478,N_8472);
and U11615 (N_11615,N_7062,N_8907);
nand U11616 (N_11616,N_7059,N_7821);
or U11617 (N_11617,N_6848,N_6754);
nor U11618 (N_11618,N_6923,N_8706);
and U11619 (N_11619,N_7408,N_8919);
nand U11620 (N_11620,N_7497,N_7773);
and U11621 (N_11621,N_6851,N_7300);
nand U11622 (N_11622,N_8472,N_7146);
or U11623 (N_11623,N_7536,N_6999);
nor U11624 (N_11624,N_6003,N_7081);
nand U11625 (N_11625,N_6414,N_6949);
nand U11626 (N_11626,N_7291,N_8613);
and U11627 (N_11627,N_6283,N_7155);
nor U11628 (N_11628,N_6756,N_6753);
and U11629 (N_11629,N_6472,N_6945);
and U11630 (N_11630,N_8913,N_6387);
or U11631 (N_11631,N_8752,N_8473);
nand U11632 (N_11632,N_7983,N_6024);
nor U11633 (N_11633,N_7223,N_8050);
or U11634 (N_11634,N_6329,N_8927);
nand U11635 (N_11635,N_8094,N_6530);
nand U11636 (N_11636,N_8291,N_7554);
and U11637 (N_11637,N_8797,N_7801);
nor U11638 (N_11638,N_7636,N_6472);
nor U11639 (N_11639,N_7334,N_7743);
xor U11640 (N_11640,N_7181,N_7097);
nor U11641 (N_11641,N_8491,N_6632);
and U11642 (N_11642,N_8664,N_6489);
nand U11643 (N_11643,N_6351,N_6457);
and U11644 (N_11644,N_8707,N_7022);
or U11645 (N_11645,N_6686,N_7597);
nand U11646 (N_11646,N_6876,N_8398);
nand U11647 (N_11647,N_7921,N_8032);
nor U11648 (N_11648,N_6559,N_8071);
nor U11649 (N_11649,N_7959,N_8708);
nand U11650 (N_11650,N_7558,N_7636);
nand U11651 (N_11651,N_7415,N_6196);
nor U11652 (N_11652,N_6786,N_7526);
nand U11653 (N_11653,N_8558,N_8508);
or U11654 (N_11654,N_7705,N_7775);
xor U11655 (N_11655,N_8396,N_8025);
nor U11656 (N_11656,N_8445,N_8691);
nand U11657 (N_11657,N_8237,N_8414);
or U11658 (N_11658,N_8193,N_7664);
and U11659 (N_11659,N_7654,N_6431);
and U11660 (N_11660,N_6328,N_8945);
and U11661 (N_11661,N_7264,N_7046);
and U11662 (N_11662,N_7641,N_7719);
or U11663 (N_11663,N_8030,N_8765);
or U11664 (N_11664,N_8861,N_7947);
or U11665 (N_11665,N_8232,N_8695);
or U11666 (N_11666,N_7460,N_7003);
and U11667 (N_11667,N_8658,N_6372);
nor U11668 (N_11668,N_6192,N_6994);
nor U11669 (N_11669,N_8618,N_8463);
and U11670 (N_11670,N_7557,N_6517);
or U11671 (N_11671,N_8989,N_6690);
or U11672 (N_11672,N_6923,N_7595);
or U11673 (N_11673,N_7598,N_8936);
xnor U11674 (N_11674,N_8978,N_8352);
or U11675 (N_11675,N_6422,N_7362);
and U11676 (N_11676,N_6706,N_8076);
and U11677 (N_11677,N_7790,N_7304);
or U11678 (N_11678,N_7830,N_7312);
nor U11679 (N_11679,N_8820,N_8503);
nor U11680 (N_11680,N_6870,N_8044);
nand U11681 (N_11681,N_6872,N_8006);
or U11682 (N_11682,N_6565,N_8492);
or U11683 (N_11683,N_7036,N_6970);
nand U11684 (N_11684,N_6904,N_7715);
nor U11685 (N_11685,N_7075,N_6848);
and U11686 (N_11686,N_6948,N_6944);
nor U11687 (N_11687,N_6599,N_7635);
nand U11688 (N_11688,N_8226,N_7200);
nor U11689 (N_11689,N_8216,N_8153);
nand U11690 (N_11690,N_8938,N_6722);
or U11691 (N_11691,N_7967,N_6532);
nand U11692 (N_11692,N_8936,N_7804);
nor U11693 (N_11693,N_7976,N_8029);
nand U11694 (N_11694,N_6985,N_6473);
nand U11695 (N_11695,N_8434,N_6896);
nor U11696 (N_11696,N_8942,N_8948);
or U11697 (N_11697,N_6114,N_7903);
or U11698 (N_11698,N_7262,N_7870);
or U11699 (N_11699,N_7748,N_8650);
and U11700 (N_11700,N_8811,N_8479);
nand U11701 (N_11701,N_6828,N_8128);
or U11702 (N_11702,N_6121,N_8925);
or U11703 (N_11703,N_6308,N_7069);
or U11704 (N_11704,N_7558,N_8372);
nor U11705 (N_11705,N_6425,N_6172);
nor U11706 (N_11706,N_6108,N_6529);
xor U11707 (N_11707,N_7198,N_6123);
nor U11708 (N_11708,N_6409,N_6775);
nand U11709 (N_11709,N_8511,N_8839);
xor U11710 (N_11710,N_6627,N_7257);
nor U11711 (N_11711,N_7303,N_7399);
and U11712 (N_11712,N_6817,N_8524);
nor U11713 (N_11713,N_6530,N_7315);
xnor U11714 (N_11714,N_6821,N_7356);
xor U11715 (N_11715,N_7093,N_8143);
and U11716 (N_11716,N_8927,N_6036);
or U11717 (N_11717,N_6838,N_7347);
and U11718 (N_11718,N_8123,N_6940);
or U11719 (N_11719,N_7981,N_7274);
nor U11720 (N_11720,N_6298,N_8842);
nor U11721 (N_11721,N_6152,N_8467);
or U11722 (N_11722,N_6299,N_7660);
nand U11723 (N_11723,N_7022,N_7276);
nor U11724 (N_11724,N_8756,N_6229);
nand U11725 (N_11725,N_6693,N_6371);
nand U11726 (N_11726,N_8573,N_6395);
or U11727 (N_11727,N_8514,N_6452);
nor U11728 (N_11728,N_6012,N_7149);
or U11729 (N_11729,N_8813,N_7798);
nor U11730 (N_11730,N_7907,N_6615);
or U11731 (N_11731,N_8991,N_8711);
nor U11732 (N_11732,N_6943,N_7674);
and U11733 (N_11733,N_6169,N_6829);
nor U11734 (N_11734,N_7922,N_7932);
and U11735 (N_11735,N_8776,N_6433);
and U11736 (N_11736,N_8395,N_7596);
and U11737 (N_11737,N_7603,N_7738);
and U11738 (N_11738,N_7318,N_6672);
nand U11739 (N_11739,N_7463,N_6808);
nand U11740 (N_11740,N_8206,N_7152);
or U11741 (N_11741,N_8861,N_7171);
nand U11742 (N_11742,N_7305,N_6050);
nand U11743 (N_11743,N_6346,N_7294);
or U11744 (N_11744,N_6475,N_8105);
nor U11745 (N_11745,N_6198,N_8021);
nand U11746 (N_11746,N_6498,N_6230);
nor U11747 (N_11747,N_7447,N_8546);
nor U11748 (N_11748,N_6960,N_8976);
nor U11749 (N_11749,N_8434,N_6395);
or U11750 (N_11750,N_8052,N_7656);
nand U11751 (N_11751,N_7001,N_7179);
nand U11752 (N_11752,N_8562,N_6738);
and U11753 (N_11753,N_6857,N_7262);
nand U11754 (N_11754,N_7992,N_7674);
or U11755 (N_11755,N_8888,N_7294);
or U11756 (N_11756,N_6458,N_8430);
nor U11757 (N_11757,N_6552,N_6078);
and U11758 (N_11758,N_8015,N_6081);
or U11759 (N_11759,N_6051,N_8828);
or U11760 (N_11760,N_7676,N_6274);
or U11761 (N_11761,N_7910,N_8596);
nand U11762 (N_11762,N_8320,N_7687);
nor U11763 (N_11763,N_6728,N_6182);
nor U11764 (N_11764,N_7309,N_8166);
nand U11765 (N_11765,N_7112,N_8664);
and U11766 (N_11766,N_7815,N_8530);
and U11767 (N_11767,N_6795,N_6794);
and U11768 (N_11768,N_8018,N_8208);
nand U11769 (N_11769,N_7075,N_6937);
nor U11770 (N_11770,N_6319,N_7189);
or U11771 (N_11771,N_6123,N_6385);
nand U11772 (N_11772,N_7440,N_8070);
nand U11773 (N_11773,N_7687,N_6125);
or U11774 (N_11774,N_8892,N_6152);
xor U11775 (N_11775,N_6370,N_6557);
or U11776 (N_11776,N_6720,N_7931);
nand U11777 (N_11777,N_7992,N_7122);
or U11778 (N_11778,N_7920,N_6607);
nand U11779 (N_11779,N_7696,N_8498);
xnor U11780 (N_11780,N_7126,N_7946);
or U11781 (N_11781,N_7098,N_7035);
and U11782 (N_11782,N_7805,N_8235);
nand U11783 (N_11783,N_7637,N_6250);
nor U11784 (N_11784,N_7682,N_7027);
nand U11785 (N_11785,N_6058,N_7057);
or U11786 (N_11786,N_6161,N_6303);
or U11787 (N_11787,N_8077,N_6366);
or U11788 (N_11788,N_6755,N_8762);
nand U11789 (N_11789,N_8820,N_6364);
nand U11790 (N_11790,N_8403,N_6251);
and U11791 (N_11791,N_7409,N_8481);
and U11792 (N_11792,N_6785,N_6629);
or U11793 (N_11793,N_8078,N_6403);
or U11794 (N_11794,N_6991,N_8397);
nor U11795 (N_11795,N_8317,N_8748);
nand U11796 (N_11796,N_8787,N_8104);
and U11797 (N_11797,N_8095,N_6993);
and U11798 (N_11798,N_6082,N_8756);
and U11799 (N_11799,N_6864,N_8768);
or U11800 (N_11800,N_7492,N_8322);
nand U11801 (N_11801,N_6833,N_8283);
nand U11802 (N_11802,N_6806,N_8652);
nor U11803 (N_11803,N_6628,N_6004);
and U11804 (N_11804,N_6309,N_8135);
or U11805 (N_11805,N_7962,N_8555);
or U11806 (N_11806,N_6014,N_8311);
and U11807 (N_11807,N_7784,N_8387);
or U11808 (N_11808,N_8500,N_6533);
or U11809 (N_11809,N_7241,N_6635);
and U11810 (N_11810,N_7412,N_7899);
nand U11811 (N_11811,N_8187,N_7069);
or U11812 (N_11812,N_8088,N_7278);
and U11813 (N_11813,N_7752,N_7648);
or U11814 (N_11814,N_7888,N_6772);
or U11815 (N_11815,N_6530,N_8912);
and U11816 (N_11816,N_7072,N_7580);
nand U11817 (N_11817,N_8446,N_6028);
nand U11818 (N_11818,N_6977,N_7519);
nand U11819 (N_11819,N_8264,N_6286);
nor U11820 (N_11820,N_8302,N_6211);
xor U11821 (N_11821,N_8117,N_7240);
nand U11822 (N_11822,N_7963,N_8124);
or U11823 (N_11823,N_7353,N_6949);
xnor U11824 (N_11824,N_6523,N_7405);
or U11825 (N_11825,N_6584,N_8417);
or U11826 (N_11826,N_8273,N_7280);
or U11827 (N_11827,N_6779,N_7870);
or U11828 (N_11828,N_7376,N_6731);
nand U11829 (N_11829,N_8607,N_6848);
nand U11830 (N_11830,N_8577,N_6585);
or U11831 (N_11831,N_8182,N_7851);
nand U11832 (N_11832,N_7023,N_7334);
nand U11833 (N_11833,N_6342,N_7629);
and U11834 (N_11834,N_8070,N_6434);
or U11835 (N_11835,N_8284,N_6796);
nand U11836 (N_11836,N_8597,N_6510);
or U11837 (N_11837,N_6568,N_7730);
or U11838 (N_11838,N_6712,N_6129);
nand U11839 (N_11839,N_6078,N_8372);
nand U11840 (N_11840,N_8738,N_6885);
or U11841 (N_11841,N_8896,N_7696);
nand U11842 (N_11842,N_7868,N_6807);
and U11843 (N_11843,N_6523,N_6272);
nor U11844 (N_11844,N_6964,N_6649);
nor U11845 (N_11845,N_8836,N_6377);
or U11846 (N_11846,N_7625,N_6718);
xor U11847 (N_11847,N_6048,N_6165);
and U11848 (N_11848,N_7473,N_8550);
and U11849 (N_11849,N_8107,N_7960);
nand U11850 (N_11850,N_7691,N_8275);
and U11851 (N_11851,N_6868,N_8554);
and U11852 (N_11852,N_6725,N_8863);
and U11853 (N_11853,N_6508,N_8125);
or U11854 (N_11854,N_6847,N_8184);
nor U11855 (N_11855,N_7217,N_8195);
and U11856 (N_11856,N_8197,N_7458);
or U11857 (N_11857,N_8652,N_8659);
and U11858 (N_11858,N_8919,N_6947);
nor U11859 (N_11859,N_6055,N_6269);
nand U11860 (N_11860,N_8967,N_7921);
nor U11861 (N_11861,N_7582,N_7819);
nor U11862 (N_11862,N_8038,N_7906);
or U11863 (N_11863,N_6115,N_6790);
or U11864 (N_11864,N_7180,N_7479);
nand U11865 (N_11865,N_8299,N_8718);
nor U11866 (N_11866,N_7577,N_6151);
nand U11867 (N_11867,N_8540,N_7080);
nor U11868 (N_11868,N_7667,N_8557);
and U11869 (N_11869,N_6857,N_6600);
nor U11870 (N_11870,N_7329,N_7220);
nor U11871 (N_11871,N_8163,N_8468);
nand U11872 (N_11872,N_8597,N_6781);
and U11873 (N_11873,N_6248,N_6467);
or U11874 (N_11874,N_6588,N_6873);
and U11875 (N_11875,N_6707,N_7623);
nand U11876 (N_11876,N_6738,N_6716);
and U11877 (N_11877,N_6461,N_8557);
and U11878 (N_11878,N_7698,N_6513);
nand U11879 (N_11879,N_7508,N_7539);
and U11880 (N_11880,N_7350,N_7010);
and U11881 (N_11881,N_8960,N_6954);
nor U11882 (N_11882,N_7393,N_8121);
nand U11883 (N_11883,N_6467,N_7952);
nand U11884 (N_11884,N_8107,N_8868);
nor U11885 (N_11885,N_6464,N_6113);
or U11886 (N_11886,N_8251,N_8976);
or U11887 (N_11887,N_6254,N_6374);
or U11888 (N_11888,N_6790,N_8881);
or U11889 (N_11889,N_7345,N_8626);
or U11890 (N_11890,N_6952,N_6899);
nor U11891 (N_11891,N_6551,N_7749);
or U11892 (N_11892,N_6460,N_6349);
nor U11893 (N_11893,N_7208,N_7303);
nor U11894 (N_11894,N_8640,N_8946);
or U11895 (N_11895,N_7656,N_8965);
nand U11896 (N_11896,N_7234,N_7216);
nor U11897 (N_11897,N_6445,N_6049);
and U11898 (N_11898,N_8879,N_8340);
or U11899 (N_11899,N_6840,N_6652);
and U11900 (N_11900,N_7953,N_6739);
or U11901 (N_11901,N_8425,N_6874);
and U11902 (N_11902,N_6230,N_8600);
and U11903 (N_11903,N_8053,N_7411);
and U11904 (N_11904,N_8852,N_6139);
nor U11905 (N_11905,N_7370,N_8256);
and U11906 (N_11906,N_6613,N_8666);
nand U11907 (N_11907,N_8838,N_7654);
nor U11908 (N_11908,N_6977,N_8241);
and U11909 (N_11909,N_8269,N_6493);
or U11910 (N_11910,N_6806,N_6840);
or U11911 (N_11911,N_7098,N_8914);
and U11912 (N_11912,N_8225,N_7032);
nand U11913 (N_11913,N_7138,N_6946);
and U11914 (N_11914,N_7684,N_7922);
or U11915 (N_11915,N_6526,N_7362);
nand U11916 (N_11916,N_7115,N_7224);
nand U11917 (N_11917,N_7301,N_8731);
or U11918 (N_11918,N_6347,N_8158);
nor U11919 (N_11919,N_6558,N_7653);
nand U11920 (N_11920,N_7448,N_6890);
nor U11921 (N_11921,N_8586,N_7540);
nor U11922 (N_11922,N_8705,N_7101);
and U11923 (N_11923,N_8378,N_7164);
and U11924 (N_11924,N_8483,N_7211);
and U11925 (N_11925,N_8982,N_8713);
nand U11926 (N_11926,N_7365,N_8653);
and U11927 (N_11927,N_8881,N_7303);
or U11928 (N_11928,N_8041,N_6611);
or U11929 (N_11929,N_6296,N_7763);
nor U11930 (N_11930,N_6469,N_7524);
nand U11931 (N_11931,N_8956,N_7959);
nand U11932 (N_11932,N_8238,N_8038);
or U11933 (N_11933,N_7167,N_8655);
nand U11934 (N_11934,N_6093,N_8989);
or U11935 (N_11935,N_7652,N_6504);
or U11936 (N_11936,N_8369,N_8482);
nor U11937 (N_11937,N_8812,N_6390);
and U11938 (N_11938,N_6562,N_8865);
nand U11939 (N_11939,N_6120,N_8445);
nor U11940 (N_11940,N_6454,N_7709);
nand U11941 (N_11941,N_6708,N_8512);
and U11942 (N_11942,N_7905,N_7897);
nand U11943 (N_11943,N_7617,N_7186);
or U11944 (N_11944,N_7716,N_7398);
nand U11945 (N_11945,N_6207,N_7504);
nand U11946 (N_11946,N_7683,N_7443);
nor U11947 (N_11947,N_6319,N_7241);
or U11948 (N_11948,N_6425,N_8201);
or U11949 (N_11949,N_8672,N_6421);
xor U11950 (N_11950,N_8464,N_7406);
and U11951 (N_11951,N_8695,N_6741);
xor U11952 (N_11952,N_7955,N_8175);
or U11953 (N_11953,N_6845,N_6930);
or U11954 (N_11954,N_6644,N_8040);
and U11955 (N_11955,N_8150,N_6504);
nor U11956 (N_11956,N_7317,N_8451);
nor U11957 (N_11957,N_8874,N_6986);
nor U11958 (N_11958,N_8389,N_8132);
and U11959 (N_11959,N_8842,N_6796);
nand U11960 (N_11960,N_6478,N_8006);
or U11961 (N_11961,N_6045,N_8159);
nand U11962 (N_11962,N_7811,N_6337);
nand U11963 (N_11963,N_6578,N_8482);
nand U11964 (N_11964,N_7169,N_7554);
and U11965 (N_11965,N_6842,N_7601);
nor U11966 (N_11966,N_8878,N_7419);
nand U11967 (N_11967,N_6933,N_6075);
or U11968 (N_11968,N_7808,N_7569);
and U11969 (N_11969,N_7217,N_8927);
or U11970 (N_11970,N_7476,N_8754);
nand U11971 (N_11971,N_6360,N_6372);
nand U11972 (N_11972,N_8166,N_6646);
nand U11973 (N_11973,N_6531,N_7202);
nor U11974 (N_11974,N_6002,N_6154);
or U11975 (N_11975,N_8192,N_8956);
nand U11976 (N_11976,N_7748,N_7615);
or U11977 (N_11977,N_8000,N_6387);
nand U11978 (N_11978,N_6385,N_6017);
nor U11979 (N_11979,N_6415,N_6168);
and U11980 (N_11980,N_8847,N_7909);
and U11981 (N_11981,N_6335,N_7957);
or U11982 (N_11982,N_8766,N_7932);
nand U11983 (N_11983,N_6984,N_6361);
nand U11984 (N_11984,N_6603,N_8668);
or U11985 (N_11985,N_6338,N_8147);
nand U11986 (N_11986,N_6171,N_8315);
and U11987 (N_11987,N_7723,N_6881);
and U11988 (N_11988,N_6394,N_8302);
nor U11989 (N_11989,N_6743,N_6337);
or U11990 (N_11990,N_8327,N_7009);
and U11991 (N_11991,N_8598,N_6079);
and U11992 (N_11992,N_6709,N_6656);
nor U11993 (N_11993,N_7457,N_8159);
nand U11994 (N_11994,N_7684,N_7893);
nand U11995 (N_11995,N_7856,N_8152);
nor U11996 (N_11996,N_8398,N_7628);
nor U11997 (N_11997,N_8938,N_6977);
and U11998 (N_11998,N_8744,N_7740);
and U11999 (N_11999,N_8104,N_6872);
nand U12000 (N_12000,N_9536,N_10586);
or U12001 (N_12001,N_10807,N_10222);
xor U12002 (N_12002,N_11967,N_9363);
nand U12003 (N_12003,N_9733,N_11240);
or U12004 (N_12004,N_9563,N_10069);
or U12005 (N_12005,N_11136,N_10072);
nor U12006 (N_12006,N_10535,N_9677);
nand U12007 (N_12007,N_10466,N_10071);
or U12008 (N_12008,N_11613,N_11480);
nand U12009 (N_12009,N_11339,N_11541);
nor U12010 (N_12010,N_11205,N_11599);
nand U12011 (N_12011,N_11884,N_9059);
nor U12012 (N_12012,N_9969,N_10711);
nand U12013 (N_12013,N_9071,N_10035);
or U12014 (N_12014,N_11002,N_9274);
or U12015 (N_12015,N_10785,N_11436);
or U12016 (N_12016,N_9655,N_11391);
nor U12017 (N_12017,N_9233,N_9523);
nor U12018 (N_12018,N_11686,N_10053);
and U12019 (N_12019,N_9282,N_11457);
nand U12020 (N_12020,N_11971,N_11807);
xnor U12021 (N_12021,N_11172,N_9076);
nand U12022 (N_12022,N_9954,N_10490);
or U12023 (N_12023,N_9322,N_11316);
nand U12024 (N_12024,N_9355,N_10361);
nand U12025 (N_12025,N_9179,N_9858);
and U12026 (N_12026,N_10600,N_10003);
or U12027 (N_12027,N_9125,N_9885);
nor U12028 (N_12028,N_11094,N_11337);
nand U12029 (N_12029,N_11673,N_9357);
nand U12030 (N_12030,N_11372,N_9814);
nor U12031 (N_12031,N_10285,N_9646);
and U12032 (N_12032,N_10126,N_9367);
xor U12033 (N_12033,N_9910,N_10210);
nor U12034 (N_12034,N_11351,N_10774);
or U12035 (N_12035,N_10217,N_11542);
and U12036 (N_12036,N_9765,N_11423);
and U12037 (N_12037,N_10160,N_9218);
nand U12038 (N_12038,N_10800,N_11593);
and U12039 (N_12039,N_9385,N_10742);
and U12040 (N_12040,N_11944,N_11727);
xor U12041 (N_12041,N_9764,N_10754);
and U12042 (N_12042,N_10067,N_10300);
nor U12043 (N_12043,N_9855,N_10993);
nand U12044 (N_12044,N_11640,N_9785);
or U12045 (N_12045,N_10756,N_11235);
and U12046 (N_12046,N_9590,N_9802);
nand U12047 (N_12047,N_10011,N_11748);
or U12048 (N_12048,N_9325,N_11112);
nand U12049 (N_12049,N_10396,N_10870);
nand U12050 (N_12050,N_11496,N_11888);
nand U12051 (N_12051,N_11620,N_11019);
nor U12052 (N_12052,N_11124,N_9628);
nor U12053 (N_12053,N_11553,N_11605);
nor U12054 (N_12054,N_9143,N_11607);
and U12055 (N_12055,N_10103,N_11459);
nand U12056 (N_12056,N_10965,N_11043);
nand U12057 (N_12057,N_9010,N_10178);
or U12058 (N_12058,N_9330,N_9888);
or U12059 (N_12059,N_11473,N_11466);
nor U12060 (N_12060,N_11144,N_10255);
nor U12061 (N_12061,N_9889,N_11030);
nor U12062 (N_12062,N_10647,N_9101);
or U12063 (N_12063,N_9253,N_11271);
or U12064 (N_12064,N_9611,N_10189);
and U12065 (N_12065,N_10463,N_11749);
nor U12066 (N_12066,N_9436,N_9130);
nor U12067 (N_12067,N_10359,N_11208);
nand U12068 (N_12068,N_10584,N_10683);
nor U12069 (N_12069,N_9745,N_10968);
and U12070 (N_12070,N_9631,N_10569);
or U12071 (N_12071,N_10141,N_10437);
nand U12072 (N_12072,N_11588,N_9196);
and U12073 (N_12073,N_11280,N_11292);
or U12074 (N_12074,N_11058,N_11489);
or U12075 (N_12075,N_9629,N_9776);
and U12076 (N_12076,N_11129,N_9600);
and U12077 (N_12077,N_9548,N_9392);
or U12078 (N_12078,N_9752,N_11806);
and U12079 (N_12079,N_11910,N_11196);
nand U12080 (N_12080,N_10699,N_9916);
or U12081 (N_12081,N_11564,N_9002);
or U12082 (N_12082,N_10493,N_11609);
nor U12083 (N_12083,N_10532,N_11074);
and U12084 (N_12084,N_10525,N_9252);
nor U12085 (N_12085,N_10575,N_9505);
nand U12086 (N_12086,N_9890,N_9199);
nand U12087 (N_12087,N_10935,N_11085);
nand U12088 (N_12088,N_9727,N_10081);
or U12089 (N_12089,N_10770,N_11691);
or U12090 (N_12090,N_11777,N_9486);
nor U12091 (N_12091,N_10290,N_9000);
or U12092 (N_12092,N_9801,N_10723);
and U12093 (N_12093,N_10443,N_9580);
or U12094 (N_12094,N_11226,N_10410);
or U12095 (N_12095,N_11476,N_11049);
xor U12096 (N_12096,N_11031,N_10385);
or U12097 (N_12097,N_11090,N_9359);
nor U12098 (N_12098,N_9375,N_11601);
and U12099 (N_12099,N_10083,N_11092);
nand U12100 (N_12100,N_9024,N_11732);
nand U12101 (N_12101,N_9191,N_10401);
and U12102 (N_12102,N_9659,N_11799);
nor U12103 (N_12103,N_9576,N_11930);
and U12104 (N_12104,N_11695,N_11922);
and U12105 (N_12105,N_10658,N_9861);
and U12106 (N_12106,N_9566,N_10029);
and U12107 (N_12107,N_10079,N_11080);
nor U12108 (N_12108,N_10681,N_10345);
or U12109 (N_12109,N_10737,N_10619);
nor U12110 (N_12110,N_11573,N_11176);
nor U12111 (N_12111,N_10892,N_11356);
nor U12112 (N_12112,N_11320,N_9517);
or U12113 (N_12113,N_9379,N_10981);
nor U12114 (N_12114,N_10707,N_10393);
nand U12115 (N_12115,N_10452,N_11314);
or U12116 (N_12116,N_11540,N_9031);
nor U12117 (N_12117,N_10641,N_9763);
nor U12118 (N_12118,N_10732,N_11750);
and U12119 (N_12119,N_9453,N_10571);
or U12120 (N_12120,N_10115,N_10592);
nand U12121 (N_12121,N_9133,N_10540);
or U12122 (N_12122,N_9609,N_10709);
nand U12123 (N_12123,N_10340,N_9020);
nand U12124 (N_12124,N_11919,N_10082);
or U12125 (N_12125,N_9264,N_10191);
nor U12126 (N_12126,N_9042,N_11441);
and U12127 (N_12127,N_10219,N_10866);
and U12128 (N_12128,N_11228,N_9216);
nor U12129 (N_12129,N_9481,N_11409);
nor U12130 (N_12130,N_10594,N_10549);
or U12131 (N_12131,N_10492,N_9533);
or U12132 (N_12132,N_10613,N_11253);
nand U12133 (N_12133,N_10779,N_9524);
and U12134 (N_12134,N_11858,N_9415);
and U12135 (N_12135,N_9963,N_10105);
nand U12136 (N_12136,N_11417,N_10025);
and U12137 (N_12137,N_11986,N_11159);
and U12138 (N_12138,N_10762,N_9480);
nor U12139 (N_12139,N_9650,N_11317);
nor U12140 (N_12140,N_9177,N_10016);
and U12141 (N_12141,N_9729,N_9873);
nand U12142 (N_12142,N_10916,N_11629);
nor U12143 (N_12143,N_9894,N_9632);
nor U12144 (N_12144,N_9660,N_10153);
nand U12145 (N_12145,N_9388,N_11632);
nand U12146 (N_12146,N_9913,N_10766);
and U12147 (N_12147,N_9248,N_9777);
xor U12148 (N_12148,N_11891,N_11330);
and U12149 (N_12149,N_10901,N_10114);
or U12150 (N_12150,N_10799,N_11187);
and U12151 (N_12151,N_10314,N_9146);
nor U12152 (N_12152,N_9514,N_10582);
or U12153 (N_12153,N_10132,N_11761);
nand U12154 (N_12154,N_10564,N_9074);
nor U12155 (N_12155,N_10252,N_10206);
nand U12156 (N_12156,N_11188,N_11942);
nor U12157 (N_12157,N_9872,N_11532);
or U12158 (N_12158,N_10491,N_11957);
xor U12159 (N_12159,N_11261,N_10043);
and U12160 (N_12160,N_10000,N_11946);
and U12161 (N_12161,N_10167,N_11778);
nor U12162 (N_12162,N_9394,N_9903);
nor U12163 (N_12163,N_11538,N_9842);
nor U12164 (N_12164,N_11341,N_11225);
nor U12165 (N_12165,N_11635,N_9255);
or U12166 (N_12166,N_9122,N_11108);
and U12167 (N_12167,N_11072,N_9259);
nor U12168 (N_12168,N_10070,N_10119);
nand U12169 (N_12169,N_9382,N_9766);
and U12170 (N_12170,N_10581,N_9791);
and U12171 (N_12171,N_9658,N_9625);
or U12172 (N_12172,N_11513,N_11837);
nand U12173 (N_12173,N_10323,N_11230);
nand U12174 (N_12174,N_11081,N_10448);
nand U12175 (N_12175,N_10149,N_10286);
nand U12176 (N_12176,N_10986,N_10041);
and U12177 (N_12177,N_10104,N_11012);
nand U12178 (N_12178,N_9689,N_9131);
nand U12179 (N_12179,N_11477,N_9892);
nand U12180 (N_12180,N_11907,N_9180);
and U12181 (N_12181,N_11528,N_10434);
nand U12182 (N_12182,N_11497,N_11373);
and U12183 (N_12183,N_10238,N_10997);
nand U12184 (N_12184,N_9877,N_11863);
or U12185 (N_12185,N_9500,N_10695);
nand U12186 (N_12186,N_9579,N_11796);
and U12187 (N_12187,N_10169,N_9732);
xor U12188 (N_12188,N_11652,N_9778);
and U12189 (N_12189,N_9174,N_10265);
nand U12190 (N_12190,N_11527,N_10527);
nor U12191 (N_12191,N_10453,N_9340);
nor U12192 (N_12192,N_11997,N_11410);
and U12193 (N_12193,N_11823,N_10636);
nor U12194 (N_12194,N_9077,N_11547);
nor U12195 (N_12195,N_10529,N_11260);
xor U12196 (N_12196,N_10100,N_10567);
and U12197 (N_12197,N_10258,N_10377);
nor U12198 (N_12198,N_11435,N_11213);
or U12199 (N_12199,N_9746,N_10203);
and U12200 (N_12200,N_10608,N_10364);
and U12201 (N_12201,N_11034,N_9879);
and U12202 (N_12202,N_10825,N_9613);
and U12203 (N_12203,N_10291,N_11862);
and U12204 (N_12204,N_10806,N_11518);
nor U12205 (N_12205,N_10601,N_10667);
nor U12206 (N_12206,N_9499,N_9496);
nor U12207 (N_12207,N_11303,N_9428);
xnor U12208 (N_12208,N_9598,N_10269);
or U12209 (N_12209,N_11171,N_10812);
and U12210 (N_12210,N_11523,N_9370);
or U12211 (N_12211,N_9951,N_10894);
nor U12212 (N_12212,N_11089,N_10014);
and U12213 (N_12213,N_11835,N_9742);
nand U12214 (N_12214,N_11560,N_10363);
nor U12215 (N_12215,N_9046,N_11234);
and U12216 (N_12216,N_10308,N_11396);
nor U12217 (N_12217,N_10531,N_9837);
nand U12218 (N_12218,N_11050,N_9210);
nand U12219 (N_12219,N_9704,N_10118);
and U12220 (N_12220,N_9671,N_9456);
or U12221 (N_12221,N_10485,N_9782);
nand U12222 (N_12222,N_10157,N_10470);
nor U12223 (N_12223,N_10175,N_11883);
nand U12224 (N_12224,N_9294,N_10316);
nor U12225 (N_12225,N_10346,N_10885);
or U12226 (N_12226,N_10591,N_11247);
or U12227 (N_12227,N_10024,N_10205);
nand U12228 (N_12228,N_11654,N_9896);
nor U12229 (N_12229,N_9984,N_9289);
nand U12230 (N_12230,N_9054,N_11965);
nor U12231 (N_12231,N_11326,N_11504);
nor U12232 (N_12232,N_11263,N_10524);
nand U12233 (N_12233,N_9051,N_11057);
nand U12234 (N_12234,N_10403,N_9229);
nor U12235 (N_12235,N_11054,N_10729);
nor U12236 (N_12236,N_9828,N_11684);
nand U12237 (N_12237,N_9056,N_11309);
xor U12238 (N_12238,N_11246,N_10772);
xor U12239 (N_12239,N_9217,N_10851);
nand U12240 (N_12240,N_11825,N_10579);
or U12241 (N_12241,N_11066,N_9265);
and U12242 (N_12242,N_10568,N_11596);
or U12243 (N_12243,N_10760,N_11747);
or U12244 (N_12244,N_9959,N_10058);
or U12245 (N_12245,N_11220,N_11842);
xor U12246 (N_12246,N_10449,N_11118);
and U12247 (N_12247,N_10486,N_9323);
or U12248 (N_12248,N_10302,N_11832);
nand U12249 (N_12249,N_11038,N_9129);
nor U12250 (N_12250,N_10367,N_10649);
or U12251 (N_12251,N_9041,N_10356);
or U12252 (N_12252,N_10122,N_10947);
nor U12253 (N_12253,N_10478,N_9883);
nor U12254 (N_12254,N_10268,N_9213);
nor U12255 (N_12255,N_10243,N_9932);
or U12256 (N_12256,N_11252,N_9830);
or U12257 (N_12257,N_10875,N_11589);
nor U12258 (N_12258,N_9315,N_10963);
and U12259 (N_12259,N_11617,N_11389);
nand U12260 (N_12260,N_9736,N_11313);
and U12261 (N_12261,N_10390,N_9539);
and U12262 (N_12262,N_11487,N_9308);
and U12263 (N_12263,N_10873,N_9559);
nand U12264 (N_12264,N_11053,N_11828);
nor U12265 (N_12265,N_11296,N_10288);
nor U12266 (N_12266,N_11819,N_11539);
nor U12267 (N_12267,N_9412,N_9943);
nor U12268 (N_12268,N_10099,N_10921);
nand U12269 (N_12269,N_10696,N_10976);
nor U12270 (N_12270,N_11614,N_10609);
nand U12271 (N_12271,N_11402,N_10065);
and U12272 (N_12272,N_10506,N_11723);
or U12273 (N_12273,N_9098,N_10773);
or U12274 (N_12274,N_11682,N_9997);
and U12275 (N_12275,N_11088,N_10859);
nor U12276 (N_12276,N_9283,N_10253);
nor U12277 (N_12277,N_9540,N_10689);
nand U12278 (N_12278,N_11281,N_10398);
nor U12279 (N_12279,N_9201,N_11503);
nor U12280 (N_12280,N_9343,N_11388);
nor U12281 (N_12281,N_10778,N_10653);
and U12282 (N_12282,N_10545,N_11522);
nand U12283 (N_12283,N_10295,N_9808);
or U12284 (N_12284,N_11264,N_9942);
or U12285 (N_12285,N_10144,N_10956);
or U12286 (N_12286,N_11386,N_11975);
nand U12287 (N_12287,N_9527,N_10933);
nor U12288 (N_12288,N_9497,N_11960);
nand U12289 (N_12289,N_10417,N_11788);
nor U12290 (N_12290,N_10309,N_10795);
or U12291 (N_12291,N_11414,N_11624);
and U12292 (N_12292,N_11745,N_9623);
or U12293 (N_12293,N_9586,N_10161);
nand U12294 (N_12294,N_11287,N_10526);
nor U12295 (N_12295,N_9687,N_9982);
nand U12296 (N_12296,N_10847,N_11751);
xnor U12297 (N_12297,N_11404,N_11288);
or U12298 (N_12298,N_11525,N_11040);
and U12299 (N_12299,N_11420,N_11084);
and U12300 (N_12300,N_10106,N_11675);
nand U12301 (N_12301,N_10728,N_9464);
and U12302 (N_12302,N_9716,N_10412);
nand U12303 (N_12303,N_10315,N_10757);
nand U12304 (N_12304,N_9543,N_11157);
or U12305 (N_12305,N_11904,N_10007);
nor U12306 (N_12306,N_9400,N_11821);
and U12307 (N_12307,N_11025,N_9106);
nand U12308 (N_12308,N_11880,N_11511);
and U12309 (N_12309,N_9028,N_9862);
nor U12310 (N_12310,N_9164,N_9794);
nand U12311 (N_12311,N_10990,N_11935);
or U12312 (N_12312,N_10702,N_11437);
nand U12313 (N_12313,N_10242,N_11375);
nand U12314 (N_12314,N_9319,N_11071);
or U12315 (N_12315,N_9637,N_9402);
or U12316 (N_12316,N_11254,N_11174);
nand U12317 (N_12317,N_11135,N_11802);
and U12318 (N_12318,N_9748,N_11087);
or U12319 (N_12319,N_9925,N_9905);
or U12320 (N_12320,N_10121,N_9413);
nor U12321 (N_12321,N_10143,N_11371);
and U12322 (N_12322,N_11991,N_9787);
nor U12323 (N_12323,N_11818,N_9409);
nand U12324 (N_12324,N_11270,N_10158);
and U12325 (N_12325,N_10063,N_10578);
and U12326 (N_12326,N_11067,N_9332);
nand U12327 (N_12327,N_10184,N_10631);
or U12328 (N_12328,N_9240,N_9171);
or U12329 (N_12329,N_10354,N_10155);
or U12330 (N_12330,N_9572,N_10088);
nand U12331 (N_12331,N_9163,N_9354);
or U12332 (N_12332,N_9907,N_9361);
nand U12333 (N_12333,N_9991,N_11906);
or U12334 (N_12334,N_9336,N_10022);
nand U12335 (N_12335,N_9437,N_10967);
nand U12336 (N_12336,N_11585,N_9928);
nand U12337 (N_12337,N_9914,N_9055);
or U12338 (N_12338,N_11036,N_9757);
nor U12339 (N_12339,N_9234,N_9734);
nor U12340 (N_12340,N_10945,N_11978);
and U12341 (N_12341,N_10218,N_10911);
nand U12342 (N_12342,N_9263,N_11328);
and U12343 (N_12343,N_9546,N_9104);
or U12344 (N_12344,N_11203,N_11923);
and U12345 (N_12345,N_9714,N_11011);
and U12346 (N_12346,N_11696,N_11364);
and U12347 (N_12347,N_9703,N_11145);
or U12348 (N_12348,N_9696,N_10661);
or U12349 (N_12349,N_11964,N_11063);
nand U12350 (N_12350,N_10339,N_9569);
or U12351 (N_12351,N_10538,N_11469);
xor U12352 (N_12352,N_10111,N_9169);
and U12353 (N_12353,N_11676,N_10301);
xor U12354 (N_12354,N_9147,N_9845);
nor U12355 (N_12355,N_9657,N_9422);
and U12356 (N_12356,N_9601,N_10198);
or U12357 (N_12357,N_10329,N_9878);
and U12358 (N_12358,N_10441,N_10381);
or U12359 (N_12359,N_11576,N_10426);
nand U12360 (N_12360,N_11524,N_11434);
and U12361 (N_12361,N_11794,N_10256);
nor U12362 (N_12362,N_11035,N_9421);
or U12363 (N_12363,N_9467,N_10908);
or U12364 (N_12364,N_9225,N_11168);
xor U12365 (N_12365,N_10960,N_11559);
and U12366 (N_12366,N_11507,N_10201);
and U12367 (N_12367,N_10985,N_9882);
nor U12368 (N_12368,N_11981,N_11005);
nor U12369 (N_12369,N_11915,N_9811);
nand U12370 (N_12370,N_10305,N_11376);
nor U12371 (N_12371,N_11853,N_9377);
nor U12372 (N_12372,N_11537,N_10332);
or U12373 (N_12373,N_11619,N_9908);
nor U12374 (N_12374,N_9521,N_10239);
or U12375 (N_12375,N_9909,N_11175);
nor U12376 (N_12376,N_9710,N_11413);
or U12377 (N_12377,N_9346,N_10277);
and U12378 (N_12378,N_11241,N_10101);
nand U12379 (N_12379,N_10321,N_11349);
nand U12380 (N_12380,N_10783,N_9328);
nand U12381 (N_12381,N_10042,N_10131);
nand U12382 (N_12382,N_9498,N_10429);
nand U12383 (N_12383,N_10726,N_9661);
and U12384 (N_12384,N_9023,N_9432);
or U12385 (N_12385,N_11618,N_11392);
and U12386 (N_12386,N_9544,N_10775);
nand U12387 (N_12387,N_10303,N_9478);
xor U12388 (N_12388,N_11905,N_11211);
nor U12389 (N_12389,N_9522,N_11369);
nand U12390 (N_12390,N_10620,N_11579);
or U12391 (N_12391,N_10949,N_11284);
and U12392 (N_12392,N_10900,N_11984);
nand U12393 (N_12393,N_10299,N_10618);
nor U12394 (N_12394,N_11911,N_10194);
or U12395 (N_12395,N_11913,N_10971);
nand U12396 (N_12396,N_9620,N_9508);
nand U12397 (N_12397,N_9119,N_9839);
nand U12398 (N_12398,N_10557,N_9475);
and U12399 (N_12399,N_10261,N_9013);
nor U12400 (N_12400,N_11003,N_11563);
nor U12401 (N_12401,N_10599,N_11784);
and U12402 (N_12402,N_10026,N_9973);
or U12403 (N_12403,N_10379,N_9256);
and U12404 (N_12404,N_10606,N_9009);
xnor U12405 (N_12405,N_9519,N_9720);
or U12406 (N_12406,N_10580,N_10755);
or U12407 (N_12407,N_10460,N_10741);
nand U12408 (N_12408,N_9605,N_11200);
nand U12409 (N_12409,N_10270,N_9649);
nand U12410 (N_12410,N_11338,N_11325);
xor U12411 (N_12411,N_10980,N_10336);
nor U12412 (N_12412,N_9534,N_10045);
nand U12413 (N_12413,N_9961,N_9309);
and U12414 (N_12414,N_9455,N_10510);
nand U12415 (N_12415,N_9953,N_9485);
nor U12416 (N_12416,N_9737,N_9468);
nor U12417 (N_12417,N_11992,N_11626);
and U12418 (N_12418,N_9178,N_11179);
nand U12419 (N_12419,N_10259,N_9927);
and U12420 (N_12420,N_9474,N_10054);
nand U12421 (N_12421,N_11555,N_9805);
nor U12422 (N_12422,N_11015,N_10895);
or U12423 (N_12423,N_9881,N_10701);
and U12424 (N_12424,N_10061,N_10929);
and U12425 (N_12425,N_10684,N_9454);
and U12426 (N_12426,N_9445,N_9859);
and U12427 (N_12427,N_11561,N_9416);
or U12428 (N_12428,N_10744,N_11401);
and U12429 (N_12429,N_10803,N_11610);
and U12430 (N_12430,N_10322,N_9109);
nand U12431 (N_12431,N_11804,N_10245);
and U12432 (N_12432,N_11584,N_9281);
and U12433 (N_12433,N_9458,N_9369);
or U12434 (N_12434,N_10123,N_11348);
or U12435 (N_12435,N_9335,N_9887);
xnor U12436 (N_12436,N_11440,N_10794);
and U12437 (N_12437,N_9097,N_9441);
and U12438 (N_12438,N_10232,N_11896);
nand U12439 (N_12439,N_11422,N_11277);
nand U12440 (N_12440,N_10874,N_11156);
nor U12441 (N_12441,N_9817,N_10366);
and U12442 (N_12442,N_9026,N_10734);
nor U12443 (N_12443,N_11709,N_9139);
nand U12444 (N_12444,N_9744,N_9080);
and U12445 (N_12445,N_11123,N_10865);
nor U12446 (N_12446,N_11494,N_11845);
and U12447 (N_12447,N_10767,N_11482);
or U12448 (N_12448,N_11447,N_9086);
and U12449 (N_12449,N_11082,N_10113);
nor U12450 (N_12450,N_10920,N_9946);
and U12451 (N_12451,N_10550,N_11329);
nand U12452 (N_12452,N_9081,N_10743);
nor U12453 (N_12453,N_11882,N_9803);
nand U12454 (N_12454,N_10846,N_11552);
nand U12455 (N_12455,N_9922,N_10673);
or U12456 (N_12456,N_11140,N_9140);
nor U12457 (N_12457,N_11486,N_10626);
nor U12458 (N_12458,N_9681,N_9254);
and U12459 (N_12459,N_10988,N_9017);
xor U12460 (N_12460,N_10512,N_9034);
nor U12461 (N_12461,N_10904,N_9089);
and U12462 (N_12462,N_9078,N_11976);
or U12463 (N_12463,N_11458,N_9112);
nor U12464 (N_12464,N_9001,N_11731);
nand U12465 (N_12465,N_11546,N_11289);
and U12466 (N_12466,N_10882,N_11568);
and U12467 (N_12467,N_11790,N_10128);
or U12468 (N_12468,N_10602,N_10440);
or U12469 (N_12469,N_10343,N_9271);
or U12470 (N_12470,N_10629,N_10724);
or U12471 (N_12471,N_11917,N_9075);
xnor U12472 (N_12472,N_10712,N_9607);
nor U12473 (N_12473,N_11945,N_11014);
nor U12474 (N_12474,N_11892,N_10502);
nor U12475 (N_12475,N_9672,N_11024);
nand U12476 (N_12476,N_9575,N_9529);
and U12477 (N_12477,N_9556,N_11683);
and U12478 (N_12478,N_10224,N_11562);
nor U12479 (N_12479,N_10116,N_10202);
nand U12480 (N_12480,N_9525,N_11644);
nor U12481 (N_12481,N_9484,N_10630);
nor U12482 (N_12482,N_10891,N_9700);
and U12483 (N_12483,N_11468,N_11519);
nor U12484 (N_12484,N_10461,N_9768);
or U12485 (N_12485,N_11041,N_11061);
nand U12486 (N_12486,N_10547,N_9507);
and U12487 (N_12487,N_11740,N_11856);
nor U12488 (N_12488,N_10279,N_11233);
nand U12489 (N_12489,N_9829,N_9347);
nor U12490 (N_12490,N_9707,N_11471);
nor U12491 (N_12491,N_11841,N_11204);
and U12492 (N_12492,N_9049,N_9220);
nor U12493 (N_12493,N_10501,N_9636);
or U12494 (N_12494,N_9815,N_9435);
and U12495 (N_12495,N_11724,N_10969);
nand U12496 (N_12496,N_11638,N_9935);
or U12497 (N_12497,N_11051,N_11502);
or U12498 (N_12498,N_11004,N_9528);
nor U12499 (N_12499,N_9504,N_10853);
nand U12500 (N_12500,N_11711,N_10562);
or U12501 (N_12501,N_10907,N_10170);
nand U12502 (N_12502,N_11700,N_9985);
nor U12503 (N_12503,N_9709,N_11362);
and U12504 (N_12504,N_11521,N_9401);
or U12505 (N_12505,N_10324,N_11429);
and U12506 (N_12506,N_9186,N_11941);
nor U12507 (N_12507,N_11427,N_10974);
nor U12508 (N_12508,N_11558,N_9393);
nor U12509 (N_12509,N_11718,N_9790);
or U12510 (N_12510,N_9476,N_11595);
and U12511 (N_12511,N_11954,N_10397);
and U12512 (N_12512,N_9772,N_10241);
nor U12513 (N_12513,N_9115,N_11826);
or U12514 (N_12514,N_10955,N_9465);
nor U12515 (N_12515,N_10341,N_11977);
nor U12516 (N_12516,N_11671,N_11467);
nor U12517 (N_12517,N_10903,N_9770);
nand U12518 (N_12518,N_9286,N_10181);
nand U12519 (N_12519,N_11190,N_11746);
nor U12520 (N_12520,N_9380,N_10708);
nand U12521 (N_12521,N_9151,N_10899);
and U12522 (N_12522,N_11193,N_10481);
and U12523 (N_12523,N_9144,N_11592);
or U12524 (N_12524,N_9564,N_9667);
and U12525 (N_12525,N_10992,N_10662);
and U12526 (N_12526,N_10573,N_10214);
or U12527 (N_12527,N_9249,N_9717);
nor U12528 (N_12528,N_9693,N_11186);
nor U12529 (N_12529,N_10639,N_10306);
xor U12530 (N_12530,N_11472,N_9461);
and U12531 (N_12531,N_10273,N_11065);
nor U12532 (N_12532,N_10686,N_11126);
or U12533 (N_12533,N_9065,N_9162);
nand U12534 (N_12534,N_10298,N_11194);
nand U12535 (N_12535,N_9293,N_11551);
nand U12536 (N_12536,N_11658,N_11022);
nor U12537 (N_12537,N_11571,N_9821);
nand U12538 (N_12538,N_10559,N_10934);
nor U12539 (N_12539,N_9944,N_11814);
or U12540 (N_12540,N_9452,N_9719);
nand U12541 (N_12541,N_10694,N_10978);
nor U12542 (N_12542,N_10798,N_9320);
nor U12543 (N_12543,N_9278,N_10972);
nand U12544 (N_12544,N_11499,N_10498);
or U12545 (N_12545,N_10693,N_9503);
nor U12546 (N_12546,N_11258,N_9082);
nor U12547 (N_12547,N_9135,N_9015);
nor U12548 (N_12548,N_9236,N_11810);
nand U12549 (N_12549,N_9756,N_9571);
nand U12550 (N_12550,N_9691,N_10625);
nand U12551 (N_12551,N_10634,N_9275);
nand U12552 (N_12552,N_9970,N_11771);
nand U12553 (N_12553,N_11446,N_9627);
or U12554 (N_12554,N_11192,N_9867);
and U12555 (N_12555,N_9103,N_11007);
and U12556 (N_12556,N_11498,N_10479);
or U12557 (N_12557,N_9653,N_10802);
nand U12558 (N_12558,N_10522,N_10715);
and U12559 (N_12559,N_9176,N_9697);
nand U12560 (N_12560,N_11479,N_11239);
and U12561 (N_12561,N_9429,N_11178);
and U12562 (N_12562,N_10304,N_11045);
and U12563 (N_12563,N_11781,N_10617);
and U12564 (N_12564,N_10771,N_11827);
nor U12565 (N_12565,N_11443,N_10952);
or U12566 (N_12566,N_11893,N_11465);
xnor U12567 (N_12567,N_9530,N_9918);
nand U12568 (N_12568,N_9462,N_11295);
nor U12569 (N_12569,N_9033,N_11150);
xnor U12570 (N_12570,N_10665,N_9136);
nand U12571 (N_12571,N_11243,N_10943);
xor U12572 (N_12572,N_10623,N_10801);
and U12573 (N_12573,N_10165,N_11820);
or U12574 (N_12574,N_11431,N_9188);
nor U12575 (N_12575,N_11475,N_11969);
and U12576 (N_12576,N_10360,N_11298);
and U12577 (N_12577,N_9141,N_9442);
or U12578 (N_12578,N_9762,N_10505);
nor U12579 (N_12579,N_11426,N_9390);
and U12580 (N_12580,N_11353,N_10721);
xnor U12581 (N_12581,N_11754,N_11567);
and U12582 (N_12582,N_9550,N_10635);
nand U12583 (N_12583,N_9060,N_10380);
or U12584 (N_12584,N_10910,N_10796);
and U12585 (N_12585,N_9223,N_11886);
nand U12586 (N_12586,N_10247,N_11358);
and U12587 (N_12587,N_9302,N_11073);
nor U12588 (N_12588,N_9156,N_9084);
and U12589 (N_12589,N_10156,N_9874);
and U12590 (N_12590,N_11849,N_9850);
and U12591 (N_12591,N_10091,N_11844);
nand U12592 (N_12592,N_11674,N_10432);
nand U12593 (N_12593,N_10520,N_10428);
nand U12594 (N_12594,N_9612,N_9383);
nand U12595 (N_12595,N_11714,N_11379);
nand U12596 (N_12596,N_11079,N_10476);
nor U12597 (N_12597,N_9224,N_11813);
or U12598 (N_12598,N_9092,N_9818);
nand U12599 (N_12599,N_9663,N_11685);
and U12600 (N_12600,N_11667,N_11237);
nand U12601 (N_12601,N_11989,N_9868);
nand U12602 (N_12602,N_9352,N_10221);
nor U12603 (N_12603,N_10928,N_9721);
or U12604 (N_12604,N_11438,N_10148);
nand U12605 (N_12605,N_10678,N_9535);
nand U12606 (N_12606,N_10484,N_11508);
nor U12607 (N_12607,N_9834,N_9864);
and U12608 (N_12608,N_9057,N_9952);
nor U12609 (N_12609,N_10719,N_10832);
and U12610 (N_12610,N_11999,N_10480);
or U12611 (N_12611,N_10318,N_11765);
nor U12612 (N_12612,N_9972,N_11775);
or U12613 (N_12613,N_10836,N_11953);
or U12614 (N_12614,N_9644,N_11877);
nand U12615 (N_12615,N_9823,N_11831);
and U12616 (N_12616,N_11972,N_9920);
and U12617 (N_12617,N_11864,N_9538);
and U12618 (N_12618,N_10674,N_11860);
or U12619 (N_12619,N_11077,N_10337);
or U12620 (N_12620,N_10597,N_10643);
and U12621 (N_12621,N_11661,N_9495);
and U12622 (N_12622,N_11310,N_11008);
nand U12623 (N_12623,N_11481,N_11286);
nand U12624 (N_12624,N_11817,N_11822);
nand U12625 (N_12625,N_10951,N_10705);
nor U12626 (N_12626,N_10488,N_11594);
nand U12627 (N_12627,N_10312,N_11603);
and U12628 (N_12628,N_10375,N_11980);
nor U12629 (N_12629,N_10563,N_11808);
nor U12630 (N_12630,N_10738,N_11324);
or U12631 (N_12631,N_9381,N_10459);
nand U12632 (N_12632,N_11432,N_10552);
or U12633 (N_12633,N_11994,N_10319);
nand U12634 (N_12634,N_10835,N_10052);
or U12635 (N_12635,N_10930,N_10566);
xnor U12636 (N_12636,N_11897,N_10445);
or U12637 (N_12637,N_11780,N_11433);
nand U12638 (N_12638,N_11055,N_9209);
or U12639 (N_12639,N_11461,N_10508);
xor U12640 (N_12640,N_9227,N_10706);
and U12641 (N_12641,N_11838,N_10444);
or U12642 (N_12642,N_9638,N_9974);
nand U12643 (N_12643,N_11006,N_9239);
or U12644 (N_12644,N_9652,N_10296);
nand U12645 (N_12645,N_11664,N_11962);
nand U12646 (N_12646,N_10248,N_11142);
or U12647 (N_12647,N_9280,N_10112);
or U12648 (N_12648,N_10333,N_9300);
nand U12649 (N_12649,N_10196,N_10038);
and U12650 (N_12650,N_10235,N_9978);
nor U12651 (N_12651,N_9152,N_10005);
nand U12652 (N_12652,N_11924,N_11939);
and U12653 (N_12653,N_9313,N_10495);
and U12654 (N_12654,N_11268,N_9595);
or U12655 (N_12655,N_11526,N_11411);
nand U12656 (N_12656,N_10439,N_11753);
nand U12657 (N_12657,N_9809,N_11580);
or U12658 (N_12658,N_11650,N_11951);
nand U12659 (N_12659,N_9725,N_11106);
nor U12660 (N_12660,N_9553,N_9202);
nor U12661 (N_12661,N_11026,N_9244);
and U12662 (N_12662,N_9898,N_11424);
and U12663 (N_12663,N_9993,N_11565);
nand U12664 (N_12664,N_11165,N_9599);
nand U12665 (N_12665,N_9250,N_11660);
nor U12666 (N_12666,N_9683,N_11215);
or U12667 (N_12667,N_10863,N_11017);
nand U12668 (N_12668,N_10047,N_10937);
nor U12669 (N_12669,N_10136,N_9880);
nand U12670 (N_12670,N_9198,N_10108);
and U12671 (N_12671,N_9342,N_11987);
or U12672 (N_12672,N_9424,N_10034);
nor U12673 (N_12673,N_9775,N_11306);
nand U12674 (N_12674,N_11550,N_10320);
nand U12675 (N_12675,N_11631,N_11042);
nand U12676 (N_12676,N_10477,N_9622);
nor U12677 (N_12677,N_11737,N_11321);
and U12678 (N_12678,N_11350,N_11415);
nand U12679 (N_12679,N_9444,N_10850);
and U12680 (N_12680,N_10809,N_9287);
and U12681 (N_12681,N_11444,N_9079);
nand U12682 (N_12682,N_11517,N_11151);
and U12683 (N_12683,N_9915,N_10096);
nor U12684 (N_12684,N_9558,N_9306);
nor U12685 (N_12685,N_10879,N_10176);
nor U12686 (N_12686,N_9288,N_10861);
nand U12687 (N_12687,N_9314,N_9852);
nor U12688 (N_12688,N_9899,N_11291);
or U12689 (N_12689,N_11127,N_9781);
or U12690 (N_12690,N_11717,N_11183);
and U12691 (N_12691,N_11332,N_10828);
or U12692 (N_12692,N_9155,N_11416);
and U12693 (N_12693,N_11574,N_10753);
nand U12694 (N_12694,N_9986,N_9822);
or U12695 (N_12695,N_11219,N_9698);
nor U12696 (N_12696,N_9948,N_9088);
nor U12697 (N_12697,N_9376,N_9870);
or U12698 (N_12698,N_11693,N_9053);
or U12699 (N_12699,N_11672,N_9741);
nand U12700 (N_12700,N_10236,N_10447);
nand U12701 (N_12701,N_10489,N_9585);
or U12702 (N_12702,N_9773,N_10284);
or U12703 (N_12703,N_11716,N_11920);
or U12704 (N_12704,N_11943,N_10994);
or U12705 (N_12705,N_10659,N_9933);
and U12706 (N_12706,N_9205,N_9578);
nand U12707 (N_12707,N_9792,N_9257);
nor U12708 (N_12708,N_10890,N_11335);
or U12709 (N_12709,N_9187,N_10276);
and U12710 (N_12710,N_10097,N_10867);
nand U12711 (N_12711,N_9482,N_11143);
nor U12712 (N_12712,N_11227,N_9573);
nand U12713 (N_12713,N_11816,N_11566);
nor U12714 (N_12714,N_11662,N_9616);
or U12715 (N_12715,N_11657,N_9305);
nor U12716 (N_12716,N_9168,N_10257);
or U12717 (N_12717,N_10792,N_9127);
and U12718 (N_12718,N_10675,N_9771);
nor U12719 (N_12719,N_10098,N_10877);
xor U12720 (N_12720,N_9457,N_10260);
nand U12721 (N_12721,N_10691,N_11250);
and U12722 (N_12722,N_9971,N_11448);
xor U12723 (N_12723,N_10946,N_10787);
nand U12724 (N_12724,N_9759,N_11642);
and U12725 (N_12725,N_10926,N_10209);
nor U12726 (N_12726,N_11236,N_10399);
nand U12727 (N_12727,N_11855,N_11846);
nand U12728 (N_12728,N_10162,N_11901);
nand U12729 (N_12729,N_9581,N_10788);
nor U12730 (N_12730,N_9906,N_11738);
nor U12731 (N_12731,N_11119,N_10127);
nor U12732 (N_12732,N_10593,N_9296);
nand U12733 (N_12733,N_11602,N_10632);
or U12734 (N_12734,N_11583,N_11643);
nand U12735 (N_12735,N_11133,N_10811);
and U12736 (N_12736,N_10858,N_9532);
xor U12737 (N_12737,N_11493,N_9405);
or U12738 (N_12738,N_10180,N_9675);
nor U12739 (N_12739,N_9979,N_10095);
or U12740 (N_12740,N_9848,N_9583);
nor U12741 (N_12741,N_9856,N_11009);
nor U12742 (N_12742,N_10970,N_10731);
or U12743 (N_12743,N_10019,N_9512);
nor U12744 (N_12744,N_9064,N_9194);
and U12745 (N_12745,N_10769,N_10164);
or U12746 (N_12746,N_10373,N_10614);
nor U12747 (N_12747,N_11634,N_10676);
nor U12748 (N_12748,N_11697,N_9329);
nand U12749 (N_12749,N_10791,N_11070);
and U12750 (N_12750,N_9463,N_9321);
nor U12751 (N_12751,N_10605,N_9836);
xor U12752 (N_12752,N_9349,N_11340);
and U12753 (N_12753,N_11857,N_10425);
or U12754 (N_12754,N_10735,N_9154);
nor U12755 (N_12755,N_10213,N_9515);
nand U12756 (N_12756,N_11963,N_11269);
or U12757 (N_12757,N_10818,N_10962);
xnor U12758 (N_12758,N_10685,N_10843);
nand U12759 (N_12759,N_10465,N_9027);
nor U12760 (N_12760,N_9269,N_11044);
nand U12761 (N_12761,N_11979,N_10372);
or U12762 (N_12762,N_11646,N_9159);
and U12763 (N_12763,N_11774,N_9806);
nand U12764 (N_12764,N_9371,N_9341);
or U12765 (N_12765,N_10588,N_9594);
nand U12766 (N_12766,N_10917,N_9955);
and U12767 (N_12767,N_10414,N_9712);
and U12768 (N_12768,N_10395,N_11290);
nand U12769 (N_12769,N_10500,N_10925);
and U12770 (N_12770,N_9726,N_9551);
nand U12771 (N_12771,N_10177,N_10249);
and U12772 (N_12772,N_9708,N_11959);
xnor U12773 (N_12773,N_9395,N_9316);
and U12774 (N_12774,N_11056,N_9626);
nand U12775 (N_12775,N_11556,N_10752);
or U12776 (N_12776,N_9312,N_10326);
and U12777 (N_12777,N_9506,N_9364);
nand U12778 (N_12778,N_10725,N_9665);
nor U12779 (N_12779,N_10130,N_11209);
and U12780 (N_12780,N_10814,N_9753);
and U12781 (N_12781,N_10621,N_9668);
nor U12782 (N_12782,N_11052,N_10880);
nand U12783 (N_12783,N_9266,N_11868);
and U12784 (N_12784,N_11786,N_9930);
or U12785 (N_12785,N_9560,N_9195);
and U12786 (N_12786,N_9987,N_11029);
or U12787 (N_12787,N_11195,N_10468);
and U12788 (N_12788,N_11095,N_9891);
or U12789 (N_12789,N_10871,N_11741);
and U12790 (N_12790,N_10826,N_9807);
nor U12791 (N_12791,N_10824,N_11097);
and U12792 (N_12792,N_10062,N_11633);
nor U12793 (N_12793,N_10740,N_9547);
nor U12794 (N_12794,N_10124,N_10415);
nor U12795 (N_12795,N_11229,N_11948);
nor U12796 (N_12796,N_9926,N_9414);
nand U12797 (N_12797,N_10615,N_9344);
and U12798 (N_12798,N_9584,N_10384);
nand U12799 (N_12799,N_10964,N_10307);
or U12800 (N_12800,N_11681,N_10442);
and U12801 (N_12801,N_9399,N_10745);
and U12802 (N_12802,N_11866,N_9876);
nor U12803 (N_12803,N_11308,N_11463);
nand U12804 (N_12804,N_10147,N_11879);
nand U12805 (N_12805,N_11116,N_9443);
and U12806 (N_12806,N_9235,N_9574);
and U12807 (N_12807,N_9608,N_10152);
or U12808 (N_12808,N_10710,N_10852);
or U12809 (N_12809,N_11125,N_10869);
nor U12810 (N_12810,N_11582,N_10515);
nor U12811 (N_12811,N_11060,N_9960);
xnor U12812 (N_12812,N_10228,N_10183);
and U12813 (N_12813,N_11743,N_10854);
and U12814 (N_12814,N_11692,N_10950);
xor U12815 (N_12815,N_9843,N_9284);
nand U12816 (N_12816,N_11739,N_9285);
nor U12817 (N_12817,N_11406,N_11850);
nand U12818 (N_12818,N_9360,N_11251);
nor U12819 (N_12819,N_11721,N_11783);
nor U12820 (N_12820,N_11212,N_11154);
nor U12821 (N_12821,N_10135,N_10446);
or U12822 (N_12822,N_10382,N_11713);
and U12823 (N_12823,N_10310,N_9005);
or U12824 (N_12824,N_9114,N_9783);
nand U12825 (N_12825,N_10017,N_11952);
nand U12826 (N_12826,N_9541,N_11450);
and U12827 (N_12827,N_11791,N_9116);
xnor U12828 (N_12828,N_11591,N_9110);
or U12829 (N_12829,N_10915,N_10120);
xor U12830 (N_12830,N_11859,N_11093);
xor U12831 (N_12831,N_11995,N_9113);
nand U12832 (N_12832,N_10838,N_11158);
nand U12833 (N_12833,N_9664,N_9501);
xnor U12834 (N_12834,N_11742,N_9863);
nor U12835 (N_12835,N_11867,N_10897);
xor U12836 (N_12836,N_9797,N_11304);
or U12837 (N_12837,N_11678,N_10031);
nor U12838 (N_12838,N_9813,N_11840);
and U12839 (N_12839,N_10289,N_10688);
nor U12840 (N_12840,N_9483,N_10110);
nand U12841 (N_12841,N_10427,N_9810);
and U12842 (N_12842,N_9670,N_9980);
nor U12843 (N_12843,N_10645,N_10086);
and U12844 (N_12844,N_11985,N_9731);
nor U12845 (N_12845,N_10066,N_9949);
and U12846 (N_12846,N_10431,N_10138);
nand U12847 (N_12847,N_10827,N_10474);
or U12848 (N_12848,N_9520,N_9921);
nor U12849 (N_12849,N_9094,N_10350);
or U12850 (N_12850,N_11800,N_11898);
and U12851 (N_12851,N_11354,N_9222);
nor U12852 (N_12852,N_11453,N_9430);
nor U12853 (N_12853,N_10020,N_10404);
or U12854 (N_12854,N_10936,N_11274);
nor U12855 (N_12855,N_9934,N_9231);
and U12856 (N_12856,N_10642,N_9680);
xor U12857 (N_12857,N_9107,N_10651);
nand U12858 (N_12858,N_11961,N_10887);
nand U12859 (N_12859,N_9126,N_9091);
or U12860 (N_12860,N_9157,N_10487);
or U12861 (N_12861,N_11367,N_9016);
or U12862 (N_12862,N_10680,N_11322);
or U12863 (N_12863,N_9743,N_11873);
or U12864 (N_12864,N_9100,N_11782);
or U12865 (N_12865,N_10516,N_10570);
nor U12866 (N_12866,N_11223,N_9450);
or U12867 (N_12867,N_10358,N_11854);
nor U12868 (N_12868,N_10961,N_9642);
xnor U12869 (N_12869,N_11789,N_11557);
nor U12870 (N_12870,N_9471,N_9214);
nor U12871 (N_12871,N_11059,N_10407);
nor U12872 (N_12872,N_10454,N_9230);
or U12873 (N_12873,N_10953,N_10784);
nand U12874 (N_12874,N_9011,N_10654);
nor U12875 (N_12875,N_10387,N_11232);
or U12876 (N_12876,N_9964,N_9121);
nand U12877 (N_12877,N_9685,N_9433);
or U12878 (N_12878,N_10244,N_9749);
or U12879 (N_12879,N_11412,N_9337);
nand U12880 (N_12880,N_10266,N_9841);
or U12881 (N_12881,N_11608,N_10223);
nor U12882 (N_12882,N_10028,N_9869);
and U12883 (N_12883,N_10664,N_11875);
or U12884 (N_12884,N_9592,N_10834);
and U12885 (N_12885,N_11276,N_9243);
nand U12886 (N_12886,N_9844,N_11871);
and U12887 (N_12887,N_11347,N_10750);
xor U12888 (N_12888,N_10537,N_10023);
nor U12889 (N_12889,N_10938,N_10262);
nand U12890 (N_12890,N_11449,N_10671);
and U12891 (N_12891,N_11656,N_9715);
nor U12892 (N_12892,N_11506,N_11615);
or U12893 (N_12893,N_9582,N_10616);
and U12894 (N_12894,N_9602,N_10499);
or U12895 (N_12895,N_10560,N_9795);
xnor U12896 (N_12896,N_10881,N_10055);
or U12897 (N_12897,N_10954,N_9470);
and U12898 (N_12898,N_10528,N_9203);
or U12899 (N_12899,N_11757,N_9021);
nand U12900 (N_12900,N_11534,N_9241);
or U12901 (N_12901,N_10497,N_10857);
xnor U12902 (N_12902,N_11408,N_11470);
nand U12903 (N_12903,N_10690,N_9246);
and U12904 (N_12904,N_11928,N_10758);
nor U12905 (N_12905,N_11177,N_10033);
or U12906 (N_12906,N_10650,N_11032);
or U12907 (N_12907,N_9831,N_9153);
nor U12908 (N_12908,N_10451,N_9819);
nor U12909 (N_12909,N_11983,N_10713);
and U12910 (N_12910,N_10328,N_9070);
nor U12911 (N_12911,N_9045,N_11021);
or U12912 (N_12912,N_9857,N_9706);
nor U12913 (N_12913,N_10902,N_9489);
or U12914 (N_12914,N_11319,N_11302);
nor U12915 (N_12915,N_9029,N_10692);
nand U12916 (N_12916,N_10044,N_9780);
or U12917 (N_12917,N_10166,N_10009);
and U12918 (N_12918,N_10918,N_11331);
and U12919 (N_12919,N_10374,N_10064);
and U12920 (N_12920,N_9798,N_10089);
nor U12921 (N_12921,N_10278,N_11653);
nor U12922 (N_12922,N_10173,N_11889);
nand U12923 (N_12923,N_11970,N_10888);
or U12924 (N_12924,N_10996,N_9148);
and U12925 (N_12925,N_9410,N_11918);
or U12926 (N_12926,N_11839,N_11020);
nor U12927 (N_12927,N_11137,N_9567);
and U12928 (N_12928,N_10913,N_10565);
or U12929 (N_12929,N_9181,N_11852);
nor U12930 (N_12930,N_9679,N_11266);
nor U12931 (N_12931,N_9299,N_11315);
nand U12932 (N_12932,N_11166,N_11570);
nor U12933 (N_12933,N_10893,N_10494);
or U12934 (N_12934,N_9958,N_9832);
nor U12935 (N_12935,N_9272,N_9804);
or U12936 (N_12936,N_9448,N_9150);
or U12937 (N_12937,N_9052,N_9095);
nand U12938 (N_12938,N_10142,N_11430);
or U12939 (N_12939,N_11869,N_10819);
and U12940 (N_12940,N_9761,N_11509);
and U12941 (N_12941,N_10780,N_11162);
nor U12942 (N_12942,N_11836,N_11037);
and U12943 (N_12943,N_10909,N_11809);
or U12944 (N_12944,N_11812,N_9386);
and U12945 (N_12945,N_9651,N_9279);
and U12946 (N_12946,N_9800,N_9338);
or U12947 (N_12947,N_11805,N_10093);
nor U12948 (N_12948,N_11763,N_9030);
or U12949 (N_12949,N_11881,N_11238);
or U12950 (N_12950,N_11708,N_11442);
and U12951 (N_12951,N_11612,N_9981);
or U12952 (N_12952,N_10975,N_11147);
nand U12953 (N_12953,N_11587,N_10841);
nand U12954 (N_12954,N_9886,N_11163);
nor U12955 (N_12955,N_11874,N_11138);
nand U12956 (N_12956,N_9273,N_11533);
and U12957 (N_12957,N_10250,N_10117);
or U12958 (N_12958,N_11403,N_9173);
nand U12959 (N_12959,N_9722,N_10195);
or U12960 (N_12960,N_9820,N_9492);
and U12961 (N_12961,N_10125,N_10233);
and U12962 (N_12962,N_9039,N_10402);
or U12963 (N_12963,N_10006,N_9303);
and U12964 (N_12964,N_10612,N_9902);
nand U12965 (N_12965,N_10583,N_9940);
nand U12966 (N_12966,N_10436,N_10231);
nand U12967 (N_12967,N_9884,N_10862);
nand U12968 (N_12968,N_9366,N_10720);
or U12969 (N_12969,N_10906,N_11380);
or U12970 (N_12970,N_10746,N_10073);
and U12971 (N_12971,N_10751,N_9617);
nand U12972 (N_12972,N_11834,N_9643);
and U12973 (N_12973,N_10422,N_11083);
or U12974 (N_12974,N_10733,N_9090);
nor U12975 (N_12975,N_10002,N_10987);
nor U12976 (N_12976,N_10462,N_10855);
nor U12977 (N_12977,N_9134,N_10627);
and U12978 (N_12978,N_10932,N_11621);
nand U12979 (N_12979,N_11327,N_9192);
and U12980 (N_12980,N_9469,N_9799);
or U12981 (N_12981,N_11405,N_10193);
or U12982 (N_12982,N_10134,N_11460);
nor U12983 (N_12983,N_11648,N_11378);
nor U12984 (N_12984,N_10577,N_9317);
nand U12985 (N_12985,N_11181,N_9516);
nor U12986 (N_12986,N_10856,N_10553);
or U12987 (N_12987,N_10813,N_11776);
or U12988 (N_12988,N_10542,N_9977);
and U12989 (N_12989,N_11100,N_10607);
nor U12990 (N_12990,N_11767,N_9614);
nand U12991 (N_12991,N_9304,N_9656);
xor U12992 (N_12992,N_9490,N_10351);
nand U12993 (N_12993,N_9447,N_10327);
or U12994 (N_12994,N_10471,N_9919);
and U12995 (N_12995,N_10482,N_11398);
xor U12996 (N_12996,N_10283,N_11216);
and U12997 (N_12997,N_9062,N_11702);
or U12998 (N_12998,N_11569,N_9406);
and U12999 (N_12999,N_11586,N_11764);
and U13000 (N_13000,N_10473,N_11993);
and U13001 (N_13001,N_11101,N_10698);
nor U13002 (N_13002,N_9295,N_9326);
nand U13003 (N_13003,N_9165,N_11912);
nor U13004 (N_13004,N_9111,N_11224);
nor U13005 (N_13005,N_10056,N_9728);
and U13006 (N_13006,N_11670,N_9846);
nand U13007 (N_13007,N_10297,N_11755);
and U13008 (N_13008,N_11199,N_11824);
or U13009 (N_13009,N_11189,N_10611);
nand U13010 (N_13010,N_9004,N_9397);
or U13011 (N_13011,N_9211,N_9513);
nand U13012 (N_13012,N_9408,N_9692);
xor U13013 (N_13013,N_10556,N_10763);
nand U13014 (N_13014,N_9228,N_10883);
nand U13015 (N_13015,N_11134,N_11600);
and U13016 (N_13016,N_11344,N_10199);
or U13017 (N_13017,N_10405,N_11770);
or U13018 (N_13018,N_9740,N_11529);
nor U13019 (N_13019,N_10842,N_9853);
and U13020 (N_13020,N_10898,N_10805);
nor U13021 (N_13021,N_9040,N_9183);
nor U13022 (N_13022,N_10386,N_10816);
nand U13023 (N_13023,N_9789,N_11990);
nand U13024 (N_13024,N_10876,N_11885);
or U13025 (N_13025,N_10927,N_9358);
nand U13026 (N_13026,N_10657,N_10371);
nor U13027 (N_13027,N_11666,N_10820);
or U13028 (N_13028,N_9724,N_11167);
or U13029 (N_13029,N_9937,N_9840);
and U13030 (N_13030,N_9093,N_11359);
nand U13031 (N_13031,N_9048,N_9640);
or U13032 (N_13032,N_10246,N_9537);
nor U13033 (N_13033,N_9924,N_11334);
and U13034 (N_13034,N_9267,N_11120);
nor U13035 (N_13035,N_11478,N_10076);
and U13036 (N_13036,N_11647,N_9676);
or U13037 (N_13037,N_10418,N_11278);
nand U13038 (N_13038,N_9509,N_10884);
nor U13039 (N_13039,N_9419,N_10644);
and U13040 (N_13040,N_11104,N_11830);
or U13041 (N_13041,N_10018,N_11578);
or U13042 (N_13042,N_10190,N_10001);
nor U13043 (N_13043,N_11221,N_9705);
nor U13044 (N_13044,N_11098,N_9407);
or U13045 (N_13045,N_10227,N_11152);
nor U13046 (N_13046,N_11210,N_9431);
xor U13047 (N_13047,N_10610,N_9603);
nor U13048 (N_13048,N_10682,N_11343);
and U13049 (N_13049,N_10652,N_11352);
nand U13050 (N_13050,N_10450,N_11000);
nand U13051 (N_13051,N_11611,N_10628);
nor U13052 (N_13052,N_10982,N_10137);
and U13053 (N_13053,N_9466,N_10589);
and U13054 (N_13054,N_11217,N_11180);
nand U13055 (N_13055,N_9170,N_10504);
nor U13056 (N_13056,N_10469,N_11514);
nand U13057 (N_13057,N_9568,N_11275);
nand U13058 (N_13058,N_9096,N_11018);
or U13059 (N_13059,N_10914,N_11169);
and U13060 (N_13060,N_11707,N_10886);
nor U13061 (N_13061,N_10905,N_9378);
and U13062 (N_13062,N_10730,N_11606);
or U13063 (N_13063,N_9438,N_9477);
and U13064 (N_13064,N_10739,N_9035);
nor U13065 (N_13065,N_11797,N_9812);
or U13066 (N_13066,N_9145,N_11793);
and U13067 (N_13067,N_11730,N_9161);
and U13068 (N_13068,N_11028,N_10511);
and U13069 (N_13069,N_10598,N_9389);
or U13070 (N_13070,N_10254,N_9365);
nand U13071 (N_13071,N_9893,N_11581);
or U13072 (N_13072,N_11301,N_9423);
or U13073 (N_13073,N_10078,N_9618);
and U13074 (N_13074,N_9426,N_11956);
and U13075 (N_13075,N_10844,N_11762);
and U13076 (N_13076,N_9063,N_10840);
and U13077 (N_13077,N_9487,N_10423);
xor U13078 (N_13078,N_9396,N_11407);
nand U13079 (N_13079,N_9221,N_9518);
nand U13080 (N_13080,N_11900,N_9105);
and U13081 (N_13081,N_10313,N_11773);
nor U13082 (N_13082,N_11815,N_10507);
nand U13083 (N_13083,N_11694,N_11894);
nor U13084 (N_13084,N_10150,N_11257);
and U13085 (N_13085,N_11787,N_11548);
and U13086 (N_13086,N_10368,N_11929);
nor U13087 (N_13087,N_9142,N_9190);
or U13088 (N_13088,N_10878,N_10534);
nor U13089 (N_13089,N_10551,N_10923);
nor U13090 (N_13090,N_10274,N_9247);
nor U13091 (N_13091,N_10240,N_11848);
nand U13092 (N_13092,N_11111,N_10378);
and U13093 (N_13093,N_10077,N_9167);
nor U13094 (N_13094,N_10554,N_11366);
nor U13095 (N_13095,N_9911,N_9356);
nor U13096 (N_13096,N_9755,N_11360);
xnor U13097 (N_13097,N_11307,N_11387);
nor U13098 (N_13098,N_10979,N_11572);
or U13099 (N_13099,N_10924,N_9073);
or U13100 (N_13100,N_10208,N_11760);
or U13101 (N_13101,N_11047,N_11428);
nor U13102 (N_13102,N_10829,N_10817);
nor U13103 (N_13103,N_9132,N_9037);
nand U13104 (N_13104,N_9261,N_10074);
or U13105 (N_13105,N_11068,N_10226);
nand U13106 (N_13106,N_11109,N_11010);
nor U13107 (N_13107,N_11113,N_9895);
xor U13108 (N_13108,N_11998,N_10638);
nand U13109 (N_13109,N_10747,N_9014);
and U13110 (N_13110,N_10595,N_9068);
xnor U13111 (N_13111,N_9860,N_10347);
nor U13112 (N_13112,N_9182,N_10518);
or U13113 (N_13113,N_9420,N_9301);
nand U13114 (N_13114,N_10797,N_9975);
and U13115 (N_13115,N_10084,N_9333);
nand U13116 (N_13116,N_11974,N_10420);
nand U13117 (N_13117,N_10860,N_10187);
nand U13118 (N_13118,N_9374,N_10868);
nand U13119 (N_13119,N_11938,N_11305);
nor U13120 (N_13120,N_10831,N_11734);
or U13121 (N_13121,N_9411,N_11439);
nand U13122 (N_13122,N_9268,N_11419);
nand U13123 (N_13123,N_11690,N_10021);
or U13124 (N_13124,N_11492,N_11099);
and U13125 (N_13125,N_10311,N_9449);
nor U13126 (N_13126,N_10513,N_9897);
nor U13127 (N_13127,N_9999,N_9635);
or U13128 (N_13128,N_9245,N_11445);
xnor U13129 (N_13129,N_9043,N_11197);
and U13130 (N_13130,N_10761,N_9619);
nand U13131 (N_13131,N_9270,N_10736);
nand U13132 (N_13132,N_11333,N_11549);
and U13133 (N_13133,N_10438,N_10548);
and U13134 (N_13134,N_9784,N_11146);
nor U13135 (N_13135,N_9158,N_9493);
nand U13136 (N_13136,N_11688,N_11927);
and U13137 (N_13137,N_10777,N_11377);
or U13138 (N_13138,N_9639,N_11779);
or U13139 (N_13139,N_10670,N_10230);
and U13140 (N_13140,N_11530,N_11577);
and U13141 (N_13141,N_9022,N_10456);
nand U13142 (N_13142,N_10656,N_9149);
and U13143 (N_13143,N_9941,N_10163);
nand U13144 (N_13144,N_9237,N_10185);
and U13145 (N_13145,N_9666,N_11792);
nand U13146 (N_13146,N_9739,N_10748);
or U13147 (N_13147,N_11202,N_10912);
nand U13148 (N_13148,N_9007,N_9615);
and U13149 (N_13149,N_11153,N_9427);
nand U13150 (N_13150,N_10212,N_10251);
or U13151 (N_13151,N_9593,N_9479);
and U13152 (N_13152,N_11207,N_9562);
and U13153 (N_13153,N_11198,N_11604);
or U13154 (N_13154,N_11039,N_11091);
nand U13155 (N_13155,N_9606,N_10267);
nor U13156 (N_13156,N_10503,N_9947);
and U13157 (N_13157,N_10509,N_9912);
or U13158 (N_13158,N_11536,N_10049);
nand U13159 (N_13159,N_10718,N_11400);
nand U13160 (N_13160,N_11768,N_10821);
and U13161 (N_13161,N_9318,N_11346);
xnor U13162 (N_13162,N_11218,N_10388);
nand U13163 (N_13163,N_11733,N_9936);
nor U13164 (N_13164,N_10633,N_11575);
xnor U13165 (N_13165,N_11890,N_9827);
or U13166 (N_13166,N_9215,N_11023);
nor U13167 (N_13167,N_9083,N_9008);
xor U13168 (N_13168,N_9998,N_11130);
and U13169 (N_13169,N_10325,N_11214);
nand U13170 (N_13170,N_9990,N_11752);
or U13171 (N_13171,N_11103,N_9362);
nand U13172 (N_13172,N_11679,N_10211);
or U13173 (N_13173,N_11117,N_10338);
nor U13174 (N_13174,N_11715,N_9038);
and U13175 (N_13175,N_11283,N_9682);
and U13176 (N_13176,N_11937,N_9589);
nand U13177 (N_13177,N_9387,N_10159);
nor U13178 (N_13178,N_11501,N_10669);
and U13179 (N_13179,N_9124,N_11191);
or U13180 (N_13180,N_10416,N_11947);
or U13181 (N_13181,N_10392,N_10941);
and U13182 (N_13182,N_10576,N_10411);
nand U13183 (N_13183,N_11384,N_11545);
nand U13184 (N_13184,N_11636,N_9204);
and U13185 (N_13185,N_10107,N_10815);
nand U13186 (N_13186,N_11637,N_10759);
nand U13187 (N_13187,N_11735,N_11833);
or U13188 (N_13188,N_11870,N_10475);
nor U13189 (N_13189,N_10154,N_10186);
xnor U13190 (N_13190,N_10370,N_9996);
and U13191 (N_13191,N_10048,N_9555);
or U13192 (N_13192,N_9939,N_10409);
and U13193 (N_13193,N_9310,N_10558);
or U13194 (N_13194,N_9793,N_10075);
nand U13195 (N_13195,N_11932,N_10646);
nand U13196 (N_13196,N_11698,N_10833);
and U13197 (N_13197,N_11669,N_9128);
xor U13198 (N_13198,N_10555,N_9166);
nand U13199 (N_13199,N_11311,N_11395);
and U13200 (N_13200,N_9018,N_9648);
or U13201 (N_13201,N_10027,N_9067);
or U13202 (N_13202,N_10192,N_10433);
nand U13203 (N_13203,N_10587,N_11484);
and U13204 (N_13204,N_10391,N_11623);
xnor U13205 (N_13205,N_10808,N_9751);
or U13206 (N_13206,N_9292,N_9061);
or U13207 (N_13207,N_10353,N_11452);
nand U13208 (N_13208,N_9418,N_10015);
and U13209 (N_13209,N_10837,N_10330);
or U13210 (N_13210,N_9373,N_9750);
and U13211 (N_13211,N_10419,N_11756);
and U13212 (N_13212,N_11899,N_11064);
and U13213 (N_13213,N_11272,N_11222);
and U13214 (N_13214,N_11201,N_11027);
and U13215 (N_13215,N_10768,N_10050);
nor U13216 (N_13216,N_11132,N_11185);
nand U13217 (N_13217,N_11374,N_11914);
and U13218 (N_13218,N_9769,N_11803);
nor U13219 (N_13219,N_10984,N_10280);
nor U13220 (N_13220,N_11936,N_9262);
nor U13221 (N_13221,N_11267,N_9117);
nor U13222 (N_13222,N_9348,N_9604);
nor U13223 (N_13223,N_9172,N_10464);
or U13224 (N_13224,N_9587,N_9866);
nand U13225 (N_13225,N_11299,N_9904);
or U13226 (N_13226,N_11390,N_9345);
nor U13227 (N_13227,N_11908,N_9277);
and U13228 (N_13228,N_9066,N_10090);
and U13229 (N_13229,N_11323,N_11639);
and U13230 (N_13230,N_9699,N_9917);
nand U13231 (N_13231,N_11342,N_11982);
nor U13232 (N_13232,N_11865,N_11046);
nand U13233 (N_13233,N_10789,N_10216);
nor U13234 (N_13234,N_10225,N_10714);
or U13235 (N_13235,N_10944,N_10727);
or U13236 (N_13236,N_9591,N_9391);
or U13237 (N_13237,N_11139,N_10483);
and U13238 (N_13238,N_11722,N_10355);
and U13239 (N_13239,N_9747,N_10080);
nor U13240 (N_13240,N_11988,N_9208);
and U13241 (N_13241,N_10948,N_10389);
nor U13242 (N_13242,N_10544,N_11096);
or U13243 (N_13243,N_10983,N_10896);
nor U13244 (N_13244,N_10030,N_10704);
xnor U13245 (N_13245,N_9718,N_9531);
or U13246 (N_13246,N_10037,N_11294);
and U13247 (N_13247,N_10369,N_11393);
and U13248 (N_13248,N_9641,N_9502);
or U13249 (N_13249,N_11622,N_10957);
xnor U13250 (N_13250,N_9875,N_9003);
or U13251 (N_13251,N_9334,N_9695);
or U13252 (N_13252,N_10603,N_11363);
nor U13253 (N_13253,N_11282,N_11076);
and U13254 (N_13254,N_9327,N_11418);
nand U13255 (N_13255,N_9353,N_10672);
or U13256 (N_13256,N_9339,N_10294);
and U13257 (N_13257,N_9298,N_10810);
or U13258 (N_13258,N_10039,N_11628);
nand U13259 (N_13259,N_10458,N_11590);
nor U13260 (N_13260,N_9219,N_9956);
and U13261 (N_13261,N_10546,N_9901);
nand U13262 (N_13262,N_11285,N_10958);
or U13263 (N_13263,N_9425,N_11772);
or U13264 (N_13264,N_11505,N_11062);
nor U13265 (N_13265,N_9758,N_9945);
nand U13266 (N_13266,N_11365,N_11249);
nor U13267 (N_13267,N_10640,N_10129);
or U13268 (N_13268,N_10991,N_10059);
or U13269 (N_13269,N_9983,N_9184);
nand U13270 (N_13270,N_9398,N_10776);
or U13271 (N_13271,N_11451,N_11535);
and U13272 (N_13272,N_9735,N_9120);
nor U13273 (N_13273,N_11078,N_11544);
nand U13274 (N_13274,N_10999,N_10102);
nor U13275 (N_13275,N_11244,N_10845);
or U13276 (N_13276,N_11495,N_11958);
and U13277 (N_13277,N_10648,N_10220);
or U13278 (N_13278,N_10051,N_11382);
and U13279 (N_13279,N_10663,N_10036);
and U13280 (N_13280,N_10966,N_11649);
xnor U13281 (N_13281,N_11114,N_9662);
nand U13282 (N_13282,N_11454,N_11627);
and U13283 (N_13283,N_11847,N_11491);
or U13284 (N_13284,N_11483,N_11488);
nand U13285 (N_13285,N_10057,N_11490);
nand U13286 (N_13286,N_10287,N_10782);
nand U13287 (N_13287,N_11141,N_11625);
xnor U13288 (N_13288,N_10749,N_11520);
and U13289 (N_13289,N_9633,N_9047);
nor U13290 (N_13290,N_9440,N_9796);
or U13291 (N_13291,N_10561,N_10765);
nand U13292 (N_13292,N_11725,N_10087);
or U13293 (N_13293,N_11512,N_9674);
or U13294 (N_13294,N_10171,N_9694);
or U13295 (N_13295,N_9565,N_11843);
nand U13296 (N_13296,N_9597,N_9669);
and U13297 (N_13297,N_11712,N_9526);
or U13298 (N_13298,N_9621,N_11949);
nor U13299 (N_13299,N_10362,N_9966);
and U13300 (N_13300,N_9511,N_9950);
and U13301 (N_13301,N_9962,N_11231);
and U13302 (N_13302,N_11801,N_9647);
nor U13303 (N_13303,N_9238,N_10517);
or U13304 (N_13304,N_11394,N_11245);
or U13305 (N_13305,N_10094,N_10848);
nand U13306 (N_13306,N_11102,N_11704);
and U13307 (N_13307,N_9542,N_11598);
or U13308 (N_13308,N_11149,N_11131);
nand U13309 (N_13309,N_10514,N_11001);
nor U13310 (N_13310,N_10679,N_10722);
nor U13311 (N_13311,N_10533,N_11273);
and U13312 (N_13312,N_10068,N_9311);
nand U13313 (N_13313,N_11630,N_11170);
nor U13314 (N_13314,N_9788,N_10179);
or U13315 (N_13315,N_11689,N_11720);
and U13316 (N_13316,N_11048,N_9570);
or U13317 (N_13317,N_10008,N_10293);
nand U13318 (N_13318,N_10543,N_11641);
and U13319 (N_13319,N_9417,N_11383);
nor U13320 (N_13320,N_10942,N_10010);
nand U13321 (N_13321,N_10703,N_11300);
and U13322 (N_13322,N_11677,N_9929);
and U13323 (N_13323,N_10668,N_9711);
and U13324 (N_13324,N_9988,N_9723);
nor U13325 (N_13325,N_11421,N_9654);
xnor U13326 (N_13326,N_9197,N_11110);
or U13327 (N_13327,N_9610,N_11851);
nor U13328 (N_13328,N_10264,N_10292);
or U13329 (N_13329,N_9472,N_10700);
or U13330 (N_13330,N_10365,N_11013);
or U13331 (N_13331,N_11934,N_9491);
or U13332 (N_13332,N_9865,N_11255);
nand U13333 (N_13333,N_10973,N_11385);
nor U13334 (N_13334,N_10139,N_11462);
or U13335 (N_13335,N_11184,N_9767);
nand U13336 (N_13336,N_9085,N_9351);
and U13337 (N_13337,N_11921,N_10472);
nand U13338 (N_13338,N_11926,N_11798);
nor U13339 (N_13339,N_9854,N_11399);
or U13340 (N_13340,N_9849,N_9577);
or U13341 (N_13341,N_10939,N_10622);
nor U13342 (N_13342,N_11456,N_10585);
nand U13343 (N_13343,N_9160,N_10092);
nand U13344 (N_13344,N_11069,N_9058);
nand U13345 (N_13345,N_11996,N_11357);
or U13346 (N_13346,N_11265,N_9688);
nor U13347 (N_13347,N_9403,N_11759);
or U13348 (N_13348,N_9251,N_11909);
nor U13349 (N_13349,N_9686,N_10331);
xor U13350 (N_13350,N_10234,N_10572);
xnor U13351 (N_13351,N_10272,N_10467);
or U13352 (N_13352,N_11785,N_11164);
and U13353 (N_13353,N_10660,N_9087);
or U13354 (N_13354,N_9102,N_11259);
xor U13355 (N_13355,N_11173,N_9630);
or U13356 (N_13356,N_9588,N_10521);
nand U13357 (N_13357,N_11729,N_10687);
nor U13358 (N_13358,N_10455,N_11312);
nor U13359 (N_13359,N_11861,N_9976);
and U13360 (N_13360,N_11903,N_9307);
nor U13361 (N_13361,N_9290,N_11680);
nand U13362 (N_13362,N_11086,N_9025);
or U13363 (N_13363,N_9549,N_10237);
nor U13364 (N_13364,N_9368,N_11148);
nor U13365 (N_13365,N_9738,N_10317);
or U13366 (N_13366,N_9754,N_9965);
or U13367 (N_13367,N_9824,N_9069);
nor U13368 (N_13368,N_9099,N_10146);
nand U13369 (N_13369,N_11318,N_10666);
nor U13370 (N_13370,N_9036,N_11500);
nand U13371 (N_13371,N_9968,N_9957);
and U13372 (N_13372,N_10200,N_11033);
and U13373 (N_13373,N_9260,N_9331);
xor U13374 (N_13374,N_9938,N_10940);
or U13375 (N_13375,N_9189,N_10624);
nor U13376 (N_13376,N_9851,N_9372);
or U13377 (N_13377,N_9995,N_11878);
and U13378 (N_13378,N_9779,N_9634);
nor U13379 (N_13379,N_10998,N_9596);
nor U13380 (N_13380,N_9645,N_10830);
and U13381 (N_13381,N_11485,N_10839);
or U13382 (N_13382,N_11705,N_9137);
and U13383 (N_13383,N_10864,N_9108);
nor U13384 (N_13384,N_11248,N_11663);
nor U13385 (N_13385,N_10931,N_11651);
and U13386 (N_13386,N_9816,N_11474);
nor U13387 (N_13387,N_10229,N_11726);
nand U13388 (N_13388,N_10421,N_9193);
nor U13389 (N_13389,N_9989,N_11531);
nand U13390 (N_13390,N_9384,N_9297);
nor U13391 (N_13391,N_11701,N_9006);
or U13392 (N_13392,N_11925,N_11361);
nor U13393 (N_13393,N_9072,N_9258);
and U13394 (N_13394,N_11706,N_9494);
nor U13395 (N_13395,N_10168,N_10151);
nand U13396 (N_13396,N_10872,N_11370);
and U13397 (N_13397,N_9673,N_9324);
and U13398 (N_13398,N_10032,N_11425);
nand U13399 (N_13399,N_10182,N_10716);
and U13400 (N_13400,N_10406,N_9557);
xnor U13401 (N_13401,N_11703,N_10085);
or U13402 (N_13402,N_10889,N_10281);
nor U13403 (N_13403,N_9510,N_9473);
nor U13404 (N_13404,N_9838,N_10536);
nand U13405 (N_13405,N_11940,N_11687);
xor U13406 (N_13406,N_10334,N_10655);
nand U13407 (N_13407,N_9774,N_10344);
and U13408 (N_13408,N_11355,N_10496);
or U13409 (N_13409,N_11182,N_9404);
nor U13410 (N_13410,N_10424,N_11256);
nand U13411 (N_13411,N_10637,N_9451);
or U13412 (N_13412,N_10574,N_9434);
or U13413 (N_13413,N_11297,N_10004);
or U13414 (N_13414,N_11155,N_9012);
xor U13415 (N_13415,N_9994,N_11655);
nand U13416 (N_13416,N_10060,N_10989);
xnor U13417 (N_13417,N_9701,N_10352);
nor U13418 (N_13418,N_11616,N_9923);
and U13419 (N_13419,N_9044,N_9847);
xor U13420 (N_13420,N_10207,N_9992);
or U13421 (N_13421,N_9900,N_11242);
nand U13422 (N_13422,N_9554,N_11728);
nor U13423 (N_13423,N_10697,N_9678);
nor U13424 (N_13424,N_10335,N_10604);
and U13425 (N_13425,N_11121,N_10413);
or U13426 (N_13426,N_11515,N_10435);
nor U13427 (N_13427,N_9760,N_10046);
or U13428 (N_13428,N_11161,N_9175);
or U13429 (N_13429,N_10764,N_11345);
or U13430 (N_13430,N_9200,N_10539);
nand U13431 (N_13431,N_11968,N_10790);
nor U13432 (N_13432,N_11206,N_11455);
or U13433 (N_13433,N_11769,N_9545);
nor U13434 (N_13434,N_9019,N_10977);
and U13435 (N_13435,N_9561,N_11336);
nor U13436 (N_13436,N_10717,N_10215);
nor U13437 (N_13437,N_9032,N_11543);
nand U13438 (N_13438,N_11128,N_10282);
nor U13439 (N_13439,N_9350,N_11829);
nor U13440 (N_13440,N_10457,N_11160);
and U13441 (N_13441,N_9967,N_11916);
or U13442 (N_13442,N_9488,N_10786);
and U13443 (N_13443,N_10408,N_11107);
nand U13444 (N_13444,N_11645,N_10188);
nand U13445 (N_13445,N_10271,N_10357);
and U13446 (N_13446,N_9826,N_9871);
and U13447 (N_13447,N_11516,N_11665);
or U13448 (N_13448,N_11811,N_10394);
or U13449 (N_13449,N_9931,N_10995);
nand U13450 (N_13450,N_9459,N_10823);
or U13451 (N_13451,N_10174,N_9242);
or U13452 (N_13452,N_10400,N_11510);
or U13453 (N_13453,N_9050,N_10349);
nand U13454 (N_13454,N_10172,N_10519);
or U13455 (N_13455,N_11597,N_10804);
nor U13456 (N_13456,N_9460,N_11955);
or U13457 (N_13457,N_10430,N_9276);
or U13458 (N_13458,N_10677,N_9291);
nor U13459 (N_13459,N_9212,N_10342);
and U13460 (N_13460,N_11758,N_9786);
nand U13461 (N_13461,N_11876,N_11075);
xnor U13462 (N_13462,N_10012,N_10793);
nor U13463 (N_13463,N_9835,N_11872);
nor U13464 (N_13464,N_10541,N_11105);
nand U13465 (N_13465,N_10523,N_9730);
nor U13466 (N_13466,N_10040,N_11554);
nor U13467 (N_13467,N_9123,N_11887);
nand U13468 (N_13468,N_9138,N_9207);
nand U13469 (N_13469,N_10013,N_9713);
xor U13470 (N_13470,N_11744,N_9552);
nand U13471 (N_13471,N_11262,N_9702);
nor U13472 (N_13472,N_11710,N_11293);
nor U13473 (N_13473,N_11973,N_9690);
and U13474 (N_13474,N_9825,N_10133);
nand U13475 (N_13475,N_11397,N_10781);
or U13476 (N_13476,N_11464,N_11719);
nor U13477 (N_13477,N_10275,N_10959);
nand U13478 (N_13478,N_11902,N_10109);
nand U13479 (N_13479,N_9833,N_11668);
nor U13480 (N_13480,N_9439,N_11699);
nand U13481 (N_13481,N_11766,N_10263);
or U13482 (N_13482,N_10197,N_11122);
and U13483 (N_13483,N_10140,N_9684);
nand U13484 (N_13484,N_9206,N_10383);
nand U13485 (N_13485,N_9624,N_9185);
nand U13486 (N_13486,N_9232,N_11016);
or U13487 (N_13487,N_11659,N_11931);
nand U13488 (N_13488,N_10348,N_11795);
nor U13489 (N_13489,N_10204,N_11279);
nor U13490 (N_13490,N_11368,N_11115);
nor U13491 (N_13491,N_11933,N_10145);
or U13492 (N_13492,N_10919,N_11895);
and U13493 (N_13493,N_11381,N_10596);
nor U13494 (N_13494,N_9118,N_11966);
and U13495 (N_13495,N_10849,N_10590);
or U13496 (N_13496,N_9446,N_10376);
or U13497 (N_13497,N_9226,N_10922);
or U13498 (N_13498,N_10530,N_11736);
nor U13499 (N_13499,N_11950,N_10822);
nand U13500 (N_13500,N_9567,N_9680);
or U13501 (N_13501,N_9703,N_11978);
and U13502 (N_13502,N_11633,N_10647);
nor U13503 (N_13503,N_10912,N_11235);
nand U13504 (N_13504,N_11058,N_11134);
xnor U13505 (N_13505,N_11359,N_10791);
or U13506 (N_13506,N_10003,N_10328);
or U13507 (N_13507,N_11517,N_10407);
or U13508 (N_13508,N_10359,N_11990);
or U13509 (N_13509,N_11635,N_11873);
nand U13510 (N_13510,N_9704,N_9701);
nor U13511 (N_13511,N_9718,N_11680);
nand U13512 (N_13512,N_9859,N_9186);
nor U13513 (N_13513,N_10198,N_10927);
nand U13514 (N_13514,N_9851,N_10249);
nand U13515 (N_13515,N_9809,N_11262);
or U13516 (N_13516,N_9241,N_11388);
or U13517 (N_13517,N_9450,N_11509);
or U13518 (N_13518,N_9268,N_11276);
and U13519 (N_13519,N_11379,N_9137);
and U13520 (N_13520,N_11796,N_9117);
nand U13521 (N_13521,N_10423,N_11938);
and U13522 (N_13522,N_9549,N_11307);
xnor U13523 (N_13523,N_11482,N_9025);
or U13524 (N_13524,N_11098,N_10093);
nor U13525 (N_13525,N_11005,N_10516);
or U13526 (N_13526,N_10999,N_10527);
nand U13527 (N_13527,N_11214,N_10312);
nand U13528 (N_13528,N_9097,N_9758);
or U13529 (N_13529,N_11434,N_11923);
nor U13530 (N_13530,N_10936,N_9371);
nand U13531 (N_13531,N_11087,N_10541);
nor U13532 (N_13532,N_10440,N_10279);
or U13533 (N_13533,N_11505,N_10770);
nor U13534 (N_13534,N_11478,N_9207);
nand U13535 (N_13535,N_11572,N_11262);
or U13536 (N_13536,N_11013,N_10894);
or U13537 (N_13537,N_11157,N_9341);
nand U13538 (N_13538,N_11085,N_11754);
nand U13539 (N_13539,N_9864,N_10980);
and U13540 (N_13540,N_11419,N_10688);
nor U13541 (N_13541,N_11187,N_10962);
nand U13542 (N_13542,N_10099,N_11194);
nand U13543 (N_13543,N_10821,N_10528);
and U13544 (N_13544,N_10671,N_9630);
or U13545 (N_13545,N_10599,N_9036);
or U13546 (N_13546,N_11779,N_9569);
and U13547 (N_13547,N_11499,N_9820);
or U13548 (N_13548,N_10474,N_9535);
and U13549 (N_13549,N_11093,N_9653);
and U13550 (N_13550,N_10075,N_9325);
nand U13551 (N_13551,N_11497,N_10505);
nor U13552 (N_13552,N_10938,N_9257);
and U13553 (N_13553,N_10252,N_10697);
or U13554 (N_13554,N_11268,N_9385);
nand U13555 (N_13555,N_10767,N_9727);
or U13556 (N_13556,N_10885,N_10461);
nand U13557 (N_13557,N_10864,N_11085);
and U13558 (N_13558,N_11258,N_9371);
nand U13559 (N_13559,N_9314,N_11890);
or U13560 (N_13560,N_11608,N_11012);
nor U13561 (N_13561,N_11083,N_10806);
nand U13562 (N_13562,N_10700,N_10671);
or U13563 (N_13563,N_10690,N_11609);
and U13564 (N_13564,N_11966,N_9449);
and U13565 (N_13565,N_10557,N_10359);
or U13566 (N_13566,N_10341,N_10982);
nor U13567 (N_13567,N_10666,N_9041);
nand U13568 (N_13568,N_9185,N_10401);
and U13569 (N_13569,N_11487,N_10317);
or U13570 (N_13570,N_10223,N_10965);
nand U13571 (N_13571,N_10850,N_11488);
nor U13572 (N_13572,N_11944,N_10335);
nor U13573 (N_13573,N_11050,N_9010);
nand U13574 (N_13574,N_11226,N_11532);
and U13575 (N_13575,N_9477,N_11508);
or U13576 (N_13576,N_9880,N_9774);
or U13577 (N_13577,N_10602,N_10166);
and U13578 (N_13578,N_11237,N_9390);
and U13579 (N_13579,N_11444,N_10078);
xnor U13580 (N_13580,N_10766,N_11665);
or U13581 (N_13581,N_10393,N_9225);
nand U13582 (N_13582,N_9133,N_9201);
nor U13583 (N_13583,N_9892,N_10310);
and U13584 (N_13584,N_9467,N_10216);
nand U13585 (N_13585,N_9703,N_10671);
or U13586 (N_13586,N_10372,N_9615);
nand U13587 (N_13587,N_9142,N_9912);
nand U13588 (N_13588,N_9861,N_9088);
nand U13589 (N_13589,N_10102,N_9158);
nand U13590 (N_13590,N_9084,N_9637);
or U13591 (N_13591,N_11168,N_9145);
and U13592 (N_13592,N_10347,N_10925);
and U13593 (N_13593,N_9000,N_11395);
and U13594 (N_13594,N_9787,N_10698);
or U13595 (N_13595,N_11665,N_11304);
nor U13596 (N_13596,N_11626,N_10774);
or U13597 (N_13597,N_9188,N_11440);
xor U13598 (N_13598,N_9124,N_9562);
nand U13599 (N_13599,N_9902,N_11471);
nor U13600 (N_13600,N_9921,N_9750);
and U13601 (N_13601,N_9821,N_9766);
or U13602 (N_13602,N_10549,N_10378);
xnor U13603 (N_13603,N_9470,N_10299);
nor U13604 (N_13604,N_9193,N_9917);
nor U13605 (N_13605,N_9069,N_11587);
nand U13606 (N_13606,N_10074,N_10973);
or U13607 (N_13607,N_11088,N_10048);
or U13608 (N_13608,N_9270,N_11179);
nor U13609 (N_13609,N_10024,N_10599);
and U13610 (N_13610,N_11801,N_11287);
nand U13611 (N_13611,N_10235,N_10253);
and U13612 (N_13612,N_9856,N_11300);
nor U13613 (N_13613,N_9331,N_10435);
nand U13614 (N_13614,N_9159,N_10151);
nor U13615 (N_13615,N_9745,N_10894);
nor U13616 (N_13616,N_11314,N_9881);
xor U13617 (N_13617,N_11067,N_10976);
or U13618 (N_13618,N_9215,N_9428);
and U13619 (N_13619,N_11562,N_11637);
xor U13620 (N_13620,N_11499,N_10356);
or U13621 (N_13621,N_9239,N_10973);
nand U13622 (N_13622,N_9054,N_10469);
xnor U13623 (N_13623,N_10704,N_10185);
or U13624 (N_13624,N_11221,N_9843);
and U13625 (N_13625,N_11837,N_11728);
xor U13626 (N_13626,N_11698,N_11173);
or U13627 (N_13627,N_11098,N_9090);
nor U13628 (N_13628,N_10218,N_9994);
nand U13629 (N_13629,N_10837,N_9638);
and U13630 (N_13630,N_10011,N_10837);
nor U13631 (N_13631,N_9485,N_11874);
or U13632 (N_13632,N_10173,N_9035);
and U13633 (N_13633,N_9696,N_10731);
nor U13634 (N_13634,N_10181,N_9660);
nand U13635 (N_13635,N_11444,N_9458);
or U13636 (N_13636,N_11826,N_11518);
and U13637 (N_13637,N_9310,N_9181);
nor U13638 (N_13638,N_10527,N_10301);
and U13639 (N_13639,N_10547,N_11718);
nand U13640 (N_13640,N_9380,N_11859);
and U13641 (N_13641,N_9144,N_9396);
nand U13642 (N_13642,N_11368,N_9310);
and U13643 (N_13643,N_9646,N_9754);
and U13644 (N_13644,N_11489,N_10394);
nand U13645 (N_13645,N_10565,N_9378);
or U13646 (N_13646,N_9953,N_10185);
or U13647 (N_13647,N_9874,N_9520);
nor U13648 (N_13648,N_11397,N_9760);
and U13649 (N_13649,N_10583,N_9391);
or U13650 (N_13650,N_10834,N_10520);
xor U13651 (N_13651,N_11537,N_11897);
nor U13652 (N_13652,N_9822,N_9654);
or U13653 (N_13653,N_9521,N_10687);
xnor U13654 (N_13654,N_11550,N_9517);
nand U13655 (N_13655,N_11706,N_10261);
and U13656 (N_13656,N_9674,N_11395);
and U13657 (N_13657,N_11412,N_11045);
nand U13658 (N_13658,N_11783,N_11367);
nand U13659 (N_13659,N_11157,N_10898);
nor U13660 (N_13660,N_9233,N_9353);
nand U13661 (N_13661,N_10840,N_9035);
nor U13662 (N_13662,N_11153,N_9061);
or U13663 (N_13663,N_10351,N_11295);
or U13664 (N_13664,N_10326,N_11973);
or U13665 (N_13665,N_10873,N_9776);
and U13666 (N_13666,N_9300,N_11294);
nand U13667 (N_13667,N_10156,N_9064);
nand U13668 (N_13668,N_9992,N_11217);
nor U13669 (N_13669,N_10544,N_11228);
and U13670 (N_13670,N_11776,N_9846);
or U13671 (N_13671,N_10235,N_10794);
nand U13672 (N_13672,N_10112,N_10088);
xor U13673 (N_13673,N_11589,N_11650);
nor U13674 (N_13674,N_10400,N_11573);
and U13675 (N_13675,N_9916,N_11028);
nor U13676 (N_13676,N_9899,N_11030);
or U13677 (N_13677,N_9209,N_9687);
and U13678 (N_13678,N_11479,N_9476);
and U13679 (N_13679,N_9009,N_11659);
nor U13680 (N_13680,N_11472,N_10941);
and U13681 (N_13681,N_11829,N_11340);
nor U13682 (N_13682,N_9443,N_9565);
nor U13683 (N_13683,N_11604,N_10385);
and U13684 (N_13684,N_9916,N_11242);
or U13685 (N_13685,N_11265,N_11190);
or U13686 (N_13686,N_10035,N_10564);
nor U13687 (N_13687,N_10093,N_10340);
and U13688 (N_13688,N_11268,N_11085);
or U13689 (N_13689,N_10900,N_11351);
nor U13690 (N_13690,N_10512,N_11066);
nand U13691 (N_13691,N_9456,N_11237);
and U13692 (N_13692,N_9598,N_9348);
or U13693 (N_13693,N_11965,N_10480);
nor U13694 (N_13694,N_9171,N_11589);
nor U13695 (N_13695,N_9626,N_10484);
nand U13696 (N_13696,N_9861,N_11256);
nand U13697 (N_13697,N_9156,N_10075);
or U13698 (N_13698,N_9849,N_9732);
nor U13699 (N_13699,N_10104,N_10137);
nand U13700 (N_13700,N_10207,N_10325);
nor U13701 (N_13701,N_10347,N_10516);
nand U13702 (N_13702,N_10301,N_10733);
nand U13703 (N_13703,N_10818,N_11760);
and U13704 (N_13704,N_10625,N_9910);
nand U13705 (N_13705,N_9512,N_10113);
xnor U13706 (N_13706,N_9689,N_9714);
nor U13707 (N_13707,N_10112,N_11774);
nor U13708 (N_13708,N_11050,N_11873);
nand U13709 (N_13709,N_9633,N_9916);
and U13710 (N_13710,N_10360,N_11340);
and U13711 (N_13711,N_9241,N_10490);
nand U13712 (N_13712,N_10703,N_10616);
nand U13713 (N_13713,N_9541,N_11352);
nand U13714 (N_13714,N_10386,N_10840);
or U13715 (N_13715,N_11501,N_11980);
and U13716 (N_13716,N_9507,N_10020);
nor U13717 (N_13717,N_9479,N_11576);
and U13718 (N_13718,N_11213,N_11714);
nand U13719 (N_13719,N_9473,N_9657);
nand U13720 (N_13720,N_9585,N_9379);
and U13721 (N_13721,N_11878,N_10319);
and U13722 (N_13722,N_11956,N_10139);
nor U13723 (N_13723,N_10879,N_9355);
nand U13724 (N_13724,N_10798,N_9998);
nand U13725 (N_13725,N_11012,N_9978);
nand U13726 (N_13726,N_9556,N_10344);
or U13727 (N_13727,N_10460,N_11135);
or U13728 (N_13728,N_9820,N_10078);
nand U13729 (N_13729,N_11474,N_10695);
and U13730 (N_13730,N_11899,N_11259);
or U13731 (N_13731,N_11364,N_11235);
and U13732 (N_13732,N_10555,N_9918);
or U13733 (N_13733,N_10298,N_10523);
nand U13734 (N_13734,N_11046,N_9407);
nor U13735 (N_13735,N_11937,N_11061);
nand U13736 (N_13736,N_9648,N_9651);
nand U13737 (N_13737,N_11153,N_11879);
nand U13738 (N_13738,N_10968,N_11131);
and U13739 (N_13739,N_11790,N_9767);
nor U13740 (N_13740,N_10726,N_10800);
nand U13741 (N_13741,N_9001,N_10932);
nor U13742 (N_13742,N_9744,N_9882);
or U13743 (N_13743,N_9213,N_11165);
or U13744 (N_13744,N_10922,N_11636);
nand U13745 (N_13745,N_10280,N_10114);
nand U13746 (N_13746,N_11423,N_10364);
nand U13747 (N_13747,N_9948,N_11855);
or U13748 (N_13748,N_11740,N_9308);
or U13749 (N_13749,N_11759,N_9265);
or U13750 (N_13750,N_9516,N_9242);
and U13751 (N_13751,N_11965,N_11798);
or U13752 (N_13752,N_9372,N_11949);
nand U13753 (N_13753,N_9235,N_9730);
nand U13754 (N_13754,N_10323,N_10580);
xor U13755 (N_13755,N_11732,N_9087);
nand U13756 (N_13756,N_10414,N_11189);
and U13757 (N_13757,N_11784,N_11611);
or U13758 (N_13758,N_9505,N_9583);
or U13759 (N_13759,N_11357,N_11223);
or U13760 (N_13760,N_9589,N_9137);
nand U13761 (N_13761,N_9161,N_9733);
nand U13762 (N_13762,N_9143,N_9931);
nand U13763 (N_13763,N_10750,N_10890);
nand U13764 (N_13764,N_10977,N_11120);
nand U13765 (N_13765,N_11942,N_10986);
nor U13766 (N_13766,N_11312,N_10656);
nand U13767 (N_13767,N_10265,N_10750);
and U13768 (N_13768,N_10511,N_11904);
or U13769 (N_13769,N_10555,N_11223);
and U13770 (N_13770,N_11443,N_9893);
and U13771 (N_13771,N_10794,N_10022);
and U13772 (N_13772,N_10357,N_9143);
nor U13773 (N_13773,N_9262,N_9358);
and U13774 (N_13774,N_11713,N_9115);
or U13775 (N_13775,N_10368,N_9213);
and U13776 (N_13776,N_9576,N_10130);
and U13777 (N_13777,N_11235,N_10625);
and U13778 (N_13778,N_11360,N_10566);
or U13779 (N_13779,N_10459,N_11672);
nor U13780 (N_13780,N_10134,N_10910);
nand U13781 (N_13781,N_9164,N_9573);
and U13782 (N_13782,N_11195,N_11896);
and U13783 (N_13783,N_11973,N_9194);
or U13784 (N_13784,N_10135,N_11457);
or U13785 (N_13785,N_9052,N_10852);
or U13786 (N_13786,N_10335,N_10141);
and U13787 (N_13787,N_11610,N_9261);
or U13788 (N_13788,N_11201,N_11660);
nand U13789 (N_13789,N_10879,N_9299);
xor U13790 (N_13790,N_10662,N_11717);
nor U13791 (N_13791,N_11611,N_9475);
or U13792 (N_13792,N_10034,N_9486);
nor U13793 (N_13793,N_11616,N_9472);
or U13794 (N_13794,N_10231,N_11323);
or U13795 (N_13795,N_10902,N_11571);
nand U13796 (N_13796,N_10606,N_11608);
or U13797 (N_13797,N_10604,N_9419);
or U13798 (N_13798,N_9438,N_11879);
or U13799 (N_13799,N_11869,N_11808);
and U13800 (N_13800,N_11007,N_10070);
or U13801 (N_13801,N_11218,N_9497);
and U13802 (N_13802,N_11827,N_9731);
or U13803 (N_13803,N_9974,N_11707);
or U13804 (N_13804,N_9155,N_10763);
or U13805 (N_13805,N_10322,N_9700);
nand U13806 (N_13806,N_10178,N_9772);
nor U13807 (N_13807,N_10180,N_9730);
or U13808 (N_13808,N_10927,N_10539);
or U13809 (N_13809,N_9197,N_11069);
or U13810 (N_13810,N_10365,N_9608);
nor U13811 (N_13811,N_9664,N_10008);
and U13812 (N_13812,N_11874,N_9738);
nand U13813 (N_13813,N_9839,N_11179);
xnor U13814 (N_13814,N_9184,N_11964);
nor U13815 (N_13815,N_9211,N_9202);
nor U13816 (N_13816,N_10051,N_10154);
and U13817 (N_13817,N_10900,N_11771);
and U13818 (N_13818,N_9119,N_10351);
nor U13819 (N_13819,N_10465,N_10646);
and U13820 (N_13820,N_11575,N_9882);
nand U13821 (N_13821,N_9004,N_9365);
nor U13822 (N_13822,N_9005,N_11907);
or U13823 (N_13823,N_11694,N_10223);
nand U13824 (N_13824,N_9110,N_10186);
and U13825 (N_13825,N_9921,N_9530);
and U13826 (N_13826,N_10671,N_10418);
nor U13827 (N_13827,N_10218,N_11289);
or U13828 (N_13828,N_10206,N_10975);
nor U13829 (N_13829,N_9742,N_10654);
nand U13830 (N_13830,N_11552,N_11471);
nand U13831 (N_13831,N_11669,N_10981);
or U13832 (N_13832,N_10623,N_9356);
nor U13833 (N_13833,N_9250,N_9256);
nor U13834 (N_13834,N_10044,N_10264);
xor U13835 (N_13835,N_9774,N_11140);
nand U13836 (N_13836,N_11916,N_9503);
nand U13837 (N_13837,N_9962,N_9854);
nand U13838 (N_13838,N_9002,N_11834);
nand U13839 (N_13839,N_9321,N_10252);
nor U13840 (N_13840,N_11810,N_9990);
and U13841 (N_13841,N_11384,N_11634);
nor U13842 (N_13842,N_10750,N_11403);
or U13843 (N_13843,N_10194,N_10702);
and U13844 (N_13844,N_9915,N_11821);
nor U13845 (N_13845,N_9250,N_11723);
or U13846 (N_13846,N_11850,N_11367);
and U13847 (N_13847,N_9344,N_11142);
or U13848 (N_13848,N_10732,N_9362);
and U13849 (N_13849,N_10635,N_10036);
and U13850 (N_13850,N_10514,N_11675);
and U13851 (N_13851,N_9842,N_11353);
and U13852 (N_13852,N_10653,N_9821);
and U13853 (N_13853,N_9046,N_11649);
or U13854 (N_13854,N_11575,N_9378);
and U13855 (N_13855,N_9408,N_11559);
and U13856 (N_13856,N_11749,N_10292);
and U13857 (N_13857,N_10452,N_10681);
nand U13858 (N_13858,N_9546,N_9906);
or U13859 (N_13859,N_10019,N_11694);
nand U13860 (N_13860,N_10992,N_9593);
or U13861 (N_13861,N_10587,N_10316);
nand U13862 (N_13862,N_10475,N_10523);
or U13863 (N_13863,N_10889,N_9617);
or U13864 (N_13864,N_9078,N_11613);
nand U13865 (N_13865,N_11877,N_9904);
and U13866 (N_13866,N_10563,N_9232);
and U13867 (N_13867,N_9250,N_11907);
nor U13868 (N_13868,N_9342,N_11966);
nand U13869 (N_13869,N_10152,N_9872);
and U13870 (N_13870,N_10227,N_9138);
or U13871 (N_13871,N_11776,N_10688);
or U13872 (N_13872,N_9348,N_10727);
nand U13873 (N_13873,N_11461,N_10618);
or U13874 (N_13874,N_9701,N_10520);
nand U13875 (N_13875,N_11558,N_10420);
or U13876 (N_13876,N_11619,N_11386);
or U13877 (N_13877,N_9379,N_9325);
nor U13878 (N_13878,N_11321,N_11041);
nor U13879 (N_13879,N_9364,N_11491);
nor U13880 (N_13880,N_11312,N_10880);
nor U13881 (N_13881,N_9821,N_10687);
nor U13882 (N_13882,N_10692,N_11359);
nand U13883 (N_13883,N_10145,N_11784);
nand U13884 (N_13884,N_11003,N_11858);
and U13885 (N_13885,N_10242,N_10904);
and U13886 (N_13886,N_10410,N_11428);
nand U13887 (N_13887,N_11667,N_9581);
xor U13888 (N_13888,N_11101,N_10022);
or U13889 (N_13889,N_10091,N_10073);
and U13890 (N_13890,N_9677,N_11525);
nor U13891 (N_13891,N_11556,N_9683);
nand U13892 (N_13892,N_11165,N_10880);
and U13893 (N_13893,N_10534,N_10763);
and U13894 (N_13894,N_9066,N_10415);
or U13895 (N_13895,N_11157,N_10705);
nor U13896 (N_13896,N_10264,N_10755);
xnor U13897 (N_13897,N_11272,N_9537);
nor U13898 (N_13898,N_11586,N_11972);
nand U13899 (N_13899,N_11588,N_11632);
nor U13900 (N_13900,N_10201,N_9477);
and U13901 (N_13901,N_9631,N_11615);
nand U13902 (N_13902,N_10970,N_10271);
nor U13903 (N_13903,N_9234,N_11108);
or U13904 (N_13904,N_9503,N_9780);
or U13905 (N_13905,N_11009,N_11558);
nor U13906 (N_13906,N_11198,N_10227);
nand U13907 (N_13907,N_11343,N_11925);
nor U13908 (N_13908,N_10867,N_10664);
nor U13909 (N_13909,N_10579,N_11621);
nand U13910 (N_13910,N_9736,N_11024);
nand U13911 (N_13911,N_11168,N_10296);
nand U13912 (N_13912,N_11243,N_11351);
and U13913 (N_13913,N_10956,N_9309);
or U13914 (N_13914,N_10372,N_11876);
xor U13915 (N_13915,N_9834,N_9373);
and U13916 (N_13916,N_9606,N_10857);
or U13917 (N_13917,N_9334,N_10212);
and U13918 (N_13918,N_10775,N_9745);
nand U13919 (N_13919,N_9268,N_9084);
nor U13920 (N_13920,N_10301,N_9207);
or U13921 (N_13921,N_10956,N_10785);
or U13922 (N_13922,N_11260,N_9985);
or U13923 (N_13923,N_10926,N_11923);
and U13924 (N_13924,N_11513,N_11519);
and U13925 (N_13925,N_9882,N_9424);
and U13926 (N_13926,N_10502,N_9681);
nor U13927 (N_13927,N_11002,N_9675);
nand U13928 (N_13928,N_11781,N_11561);
or U13929 (N_13929,N_10179,N_9211);
and U13930 (N_13930,N_9742,N_10982);
or U13931 (N_13931,N_10957,N_11325);
or U13932 (N_13932,N_9060,N_11063);
nand U13933 (N_13933,N_10527,N_11882);
or U13934 (N_13934,N_11265,N_11883);
nor U13935 (N_13935,N_10327,N_11945);
or U13936 (N_13936,N_10699,N_10239);
nor U13937 (N_13937,N_10500,N_11855);
nor U13938 (N_13938,N_10465,N_11784);
nand U13939 (N_13939,N_10927,N_10476);
nand U13940 (N_13940,N_10113,N_11672);
or U13941 (N_13941,N_9317,N_9505);
nor U13942 (N_13942,N_10647,N_11994);
nor U13943 (N_13943,N_9406,N_9922);
nand U13944 (N_13944,N_11469,N_9097);
nor U13945 (N_13945,N_10385,N_11780);
and U13946 (N_13946,N_11950,N_9273);
or U13947 (N_13947,N_10925,N_11679);
xnor U13948 (N_13948,N_11789,N_9863);
and U13949 (N_13949,N_9773,N_9929);
nor U13950 (N_13950,N_9445,N_11396);
nor U13951 (N_13951,N_9142,N_9839);
or U13952 (N_13952,N_9987,N_10170);
and U13953 (N_13953,N_10202,N_11593);
or U13954 (N_13954,N_10861,N_10006);
nor U13955 (N_13955,N_10258,N_11915);
nand U13956 (N_13956,N_9034,N_9487);
nor U13957 (N_13957,N_9801,N_10992);
or U13958 (N_13958,N_9096,N_10772);
nand U13959 (N_13959,N_11045,N_9977);
or U13960 (N_13960,N_11392,N_11008);
or U13961 (N_13961,N_9496,N_9575);
nand U13962 (N_13962,N_11072,N_11877);
or U13963 (N_13963,N_11196,N_9980);
nor U13964 (N_13964,N_10347,N_9251);
and U13965 (N_13965,N_11421,N_11434);
nand U13966 (N_13966,N_11679,N_10074);
nand U13967 (N_13967,N_11947,N_10931);
and U13968 (N_13968,N_9525,N_11469);
nand U13969 (N_13969,N_10025,N_11095);
nor U13970 (N_13970,N_9071,N_9096);
nor U13971 (N_13971,N_10224,N_11576);
nand U13972 (N_13972,N_9764,N_11064);
and U13973 (N_13973,N_11055,N_10685);
and U13974 (N_13974,N_9092,N_10491);
or U13975 (N_13975,N_9926,N_10885);
nand U13976 (N_13976,N_11447,N_11882);
or U13977 (N_13977,N_11383,N_11253);
nor U13978 (N_13978,N_11167,N_10154);
nor U13979 (N_13979,N_9705,N_10945);
nor U13980 (N_13980,N_11177,N_11765);
and U13981 (N_13981,N_11530,N_9233);
nor U13982 (N_13982,N_9257,N_11122);
nand U13983 (N_13983,N_10978,N_11221);
and U13984 (N_13984,N_10776,N_9913);
and U13985 (N_13985,N_9205,N_10613);
nor U13986 (N_13986,N_9203,N_11798);
nand U13987 (N_13987,N_10219,N_9847);
nand U13988 (N_13988,N_10695,N_11497);
nand U13989 (N_13989,N_11852,N_11390);
nand U13990 (N_13990,N_11970,N_9016);
nor U13991 (N_13991,N_10637,N_9628);
xor U13992 (N_13992,N_11547,N_9348);
or U13993 (N_13993,N_9936,N_10855);
nand U13994 (N_13994,N_9285,N_9078);
or U13995 (N_13995,N_10085,N_10600);
nor U13996 (N_13996,N_11398,N_9741);
nor U13997 (N_13997,N_9042,N_9909);
or U13998 (N_13998,N_10364,N_11164);
nor U13999 (N_13999,N_11318,N_10515);
xor U14000 (N_14000,N_9737,N_9311);
nor U14001 (N_14001,N_11229,N_10657);
and U14002 (N_14002,N_11198,N_11156);
or U14003 (N_14003,N_10575,N_9798);
or U14004 (N_14004,N_9736,N_10495);
or U14005 (N_14005,N_9200,N_9935);
and U14006 (N_14006,N_9174,N_9492);
and U14007 (N_14007,N_11047,N_10036);
nor U14008 (N_14008,N_9453,N_9175);
and U14009 (N_14009,N_11487,N_9439);
nor U14010 (N_14010,N_9988,N_11453);
nor U14011 (N_14011,N_11429,N_9966);
nand U14012 (N_14012,N_9499,N_10088);
or U14013 (N_14013,N_9500,N_10675);
nand U14014 (N_14014,N_11836,N_11163);
and U14015 (N_14015,N_9479,N_9619);
nor U14016 (N_14016,N_11988,N_11693);
or U14017 (N_14017,N_11144,N_10874);
and U14018 (N_14018,N_9531,N_9241);
nand U14019 (N_14019,N_9783,N_9375);
or U14020 (N_14020,N_9385,N_10739);
and U14021 (N_14021,N_11780,N_10416);
nor U14022 (N_14022,N_9582,N_9654);
and U14023 (N_14023,N_11344,N_11609);
nor U14024 (N_14024,N_9619,N_11544);
nand U14025 (N_14025,N_9368,N_10335);
nor U14026 (N_14026,N_10885,N_9218);
or U14027 (N_14027,N_11383,N_11483);
nor U14028 (N_14028,N_10943,N_9484);
and U14029 (N_14029,N_9188,N_9173);
nor U14030 (N_14030,N_10602,N_9562);
or U14031 (N_14031,N_10586,N_9934);
and U14032 (N_14032,N_9929,N_10095);
nor U14033 (N_14033,N_9156,N_9063);
and U14034 (N_14034,N_9277,N_9902);
nor U14035 (N_14035,N_10158,N_10649);
nor U14036 (N_14036,N_11079,N_9630);
nand U14037 (N_14037,N_9750,N_11880);
nor U14038 (N_14038,N_9825,N_9072);
nand U14039 (N_14039,N_9578,N_9374);
or U14040 (N_14040,N_9157,N_10358);
nor U14041 (N_14041,N_9288,N_9002);
nor U14042 (N_14042,N_11316,N_11680);
or U14043 (N_14043,N_10345,N_10013);
xor U14044 (N_14044,N_11287,N_11439);
or U14045 (N_14045,N_11917,N_11023);
nand U14046 (N_14046,N_9721,N_9914);
nand U14047 (N_14047,N_11400,N_9180);
and U14048 (N_14048,N_9671,N_10535);
and U14049 (N_14049,N_10183,N_9491);
nor U14050 (N_14050,N_11418,N_9824);
nand U14051 (N_14051,N_9869,N_10267);
and U14052 (N_14052,N_10008,N_10072);
nor U14053 (N_14053,N_9439,N_9058);
or U14054 (N_14054,N_9880,N_11939);
nor U14055 (N_14055,N_9173,N_9353);
or U14056 (N_14056,N_9119,N_10988);
nor U14057 (N_14057,N_11462,N_9248);
nor U14058 (N_14058,N_10384,N_9736);
nor U14059 (N_14059,N_10099,N_9722);
nor U14060 (N_14060,N_10059,N_10031);
or U14061 (N_14061,N_10844,N_10223);
nor U14062 (N_14062,N_11187,N_10540);
or U14063 (N_14063,N_11115,N_11682);
or U14064 (N_14064,N_9733,N_11029);
or U14065 (N_14065,N_11636,N_10950);
or U14066 (N_14066,N_10221,N_10076);
nor U14067 (N_14067,N_11783,N_11976);
and U14068 (N_14068,N_10442,N_9308);
nor U14069 (N_14069,N_9378,N_10328);
or U14070 (N_14070,N_9190,N_9388);
nand U14071 (N_14071,N_11792,N_10566);
or U14072 (N_14072,N_9434,N_11415);
nand U14073 (N_14073,N_9939,N_9532);
and U14074 (N_14074,N_11073,N_10944);
nand U14075 (N_14075,N_10605,N_10853);
and U14076 (N_14076,N_11843,N_10267);
or U14077 (N_14077,N_11594,N_11774);
nand U14078 (N_14078,N_10509,N_9932);
nor U14079 (N_14079,N_11827,N_11104);
nand U14080 (N_14080,N_9230,N_11173);
nand U14081 (N_14081,N_11224,N_9465);
nand U14082 (N_14082,N_11722,N_10396);
nand U14083 (N_14083,N_9531,N_9164);
nor U14084 (N_14084,N_11055,N_10013);
nand U14085 (N_14085,N_11464,N_9809);
nand U14086 (N_14086,N_9832,N_11522);
nand U14087 (N_14087,N_11805,N_11016);
or U14088 (N_14088,N_9541,N_11205);
nand U14089 (N_14089,N_11362,N_10613);
nand U14090 (N_14090,N_9111,N_10216);
nor U14091 (N_14091,N_10588,N_9641);
nand U14092 (N_14092,N_9434,N_11424);
or U14093 (N_14093,N_10524,N_10201);
nand U14094 (N_14094,N_11687,N_9811);
or U14095 (N_14095,N_10780,N_11287);
nand U14096 (N_14096,N_11481,N_11085);
and U14097 (N_14097,N_11887,N_11876);
nand U14098 (N_14098,N_9058,N_10126);
and U14099 (N_14099,N_9570,N_10407);
nor U14100 (N_14100,N_9076,N_10234);
and U14101 (N_14101,N_11408,N_10189);
or U14102 (N_14102,N_10620,N_9915);
nor U14103 (N_14103,N_11290,N_9971);
and U14104 (N_14104,N_11226,N_11006);
nor U14105 (N_14105,N_10361,N_10458);
nor U14106 (N_14106,N_10284,N_9221);
nor U14107 (N_14107,N_11131,N_11144);
and U14108 (N_14108,N_11087,N_11688);
nand U14109 (N_14109,N_11988,N_10964);
nor U14110 (N_14110,N_10405,N_10245);
nand U14111 (N_14111,N_10840,N_10173);
or U14112 (N_14112,N_10299,N_11946);
xnor U14113 (N_14113,N_10605,N_9869);
nor U14114 (N_14114,N_9625,N_11949);
nand U14115 (N_14115,N_10809,N_9243);
nand U14116 (N_14116,N_9451,N_11843);
nand U14117 (N_14117,N_11779,N_11553);
nor U14118 (N_14118,N_10321,N_9050);
and U14119 (N_14119,N_10031,N_11778);
or U14120 (N_14120,N_10027,N_11989);
and U14121 (N_14121,N_9669,N_11869);
or U14122 (N_14122,N_10491,N_10510);
and U14123 (N_14123,N_9137,N_9906);
and U14124 (N_14124,N_10680,N_10737);
or U14125 (N_14125,N_9859,N_10669);
and U14126 (N_14126,N_11093,N_11626);
nand U14127 (N_14127,N_10176,N_9191);
nor U14128 (N_14128,N_9724,N_11687);
nor U14129 (N_14129,N_9573,N_9122);
or U14130 (N_14130,N_10808,N_11109);
and U14131 (N_14131,N_10145,N_10418);
and U14132 (N_14132,N_9588,N_10972);
or U14133 (N_14133,N_9462,N_11035);
or U14134 (N_14134,N_9025,N_9270);
or U14135 (N_14135,N_11470,N_10737);
nand U14136 (N_14136,N_10754,N_10594);
nor U14137 (N_14137,N_11486,N_11730);
nor U14138 (N_14138,N_11856,N_11598);
or U14139 (N_14139,N_9676,N_10307);
nor U14140 (N_14140,N_9184,N_11623);
or U14141 (N_14141,N_11272,N_11399);
or U14142 (N_14142,N_11297,N_10832);
nor U14143 (N_14143,N_11999,N_9652);
nor U14144 (N_14144,N_10911,N_11187);
and U14145 (N_14145,N_10507,N_10773);
nand U14146 (N_14146,N_11917,N_11815);
and U14147 (N_14147,N_11665,N_9845);
nor U14148 (N_14148,N_9185,N_9298);
or U14149 (N_14149,N_10948,N_11523);
and U14150 (N_14150,N_10602,N_11106);
nand U14151 (N_14151,N_9491,N_11896);
xnor U14152 (N_14152,N_9241,N_9110);
and U14153 (N_14153,N_9286,N_9583);
nand U14154 (N_14154,N_10581,N_9516);
and U14155 (N_14155,N_11667,N_11483);
nand U14156 (N_14156,N_9533,N_9323);
nand U14157 (N_14157,N_9638,N_9264);
nor U14158 (N_14158,N_10132,N_11935);
or U14159 (N_14159,N_10745,N_10330);
and U14160 (N_14160,N_10154,N_11719);
and U14161 (N_14161,N_11074,N_10529);
nand U14162 (N_14162,N_10882,N_11868);
nand U14163 (N_14163,N_11687,N_10685);
and U14164 (N_14164,N_9875,N_9810);
or U14165 (N_14165,N_9205,N_9585);
and U14166 (N_14166,N_9595,N_10062);
nor U14167 (N_14167,N_10816,N_10201);
or U14168 (N_14168,N_9018,N_9550);
nand U14169 (N_14169,N_9696,N_9308);
or U14170 (N_14170,N_10343,N_10021);
or U14171 (N_14171,N_10860,N_9457);
and U14172 (N_14172,N_10306,N_9875);
or U14173 (N_14173,N_10460,N_11230);
nand U14174 (N_14174,N_10074,N_11994);
nor U14175 (N_14175,N_11470,N_9327);
and U14176 (N_14176,N_11679,N_9033);
nand U14177 (N_14177,N_11880,N_11485);
or U14178 (N_14178,N_10803,N_10583);
and U14179 (N_14179,N_9772,N_11393);
nand U14180 (N_14180,N_11899,N_9805);
or U14181 (N_14181,N_10188,N_11526);
nor U14182 (N_14182,N_11458,N_11213);
xnor U14183 (N_14183,N_9978,N_9697);
or U14184 (N_14184,N_10450,N_10423);
nor U14185 (N_14185,N_11258,N_9528);
or U14186 (N_14186,N_10201,N_10539);
and U14187 (N_14187,N_10577,N_9177);
or U14188 (N_14188,N_11512,N_9716);
xor U14189 (N_14189,N_10832,N_11034);
nor U14190 (N_14190,N_11948,N_10388);
and U14191 (N_14191,N_10716,N_11345);
nand U14192 (N_14192,N_9987,N_11329);
and U14193 (N_14193,N_11785,N_10519);
and U14194 (N_14194,N_10573,N_10899);
and U14195 (N_14195,N_10929,N_10976);
or U14196 (N_14196,N_11487,N_9903);
nor U14197 (N_14197,N_9043,N_9755);
or U14198 (N_14198,N_11642,N_9557);
nor U14199 (N_14199,N_11227,N_9805);
nor U14200 (N_14200,N_10277,N_9625);
and U14201 (N_14201,N_11366,N_9471);
nand U14202 (N_14202,N_10114,N_9151);
nor U14203 (N_14203,N_10207,N_11193);
and U14204 (N_14204,N_10767,N_11767);
or U14205 (N_14205,N_9048,N_10247);
and U14206 (N_14206,N_9644,N_9001);
and U14207 (N_14207,N_10789,N_10396);
nor U14208 (N_14208,N_11945,N_9376);
and U14209 (N_14209,N_9085,N_10103);
nand U14210 (N_14210,N_10448,N_10171);
nand U14211 (N_14211,N_10768,N_11900);
nand U14212 (N_14212,N_9869,N_9010);
and U14213 (N_14213,N_9585,N_9061);
or U14214 (N_14214,N_11352,N_10592);
or U14215 (N_14215,N_11825,N_10394);
nand U14216 (N_14216,N_10928,N_11569);
xor U14217 (N_14217,N_9768,N_11366);
and U14218 (N_14218,N_9433,N_11612);
nor U14219 (N_14219,N_11646,N_9924);
nor U14220 (N_14220,N_10229,N_9784);
nand U14221 (N_14221,N_9075,N_9791);
or U14222 (N_14222,N_10739,N_10473);
xnor U14223 (N_14223,N_11441,N_10629);
nor U14224 (N_14224,N_10937,N_11564);
nand U14225 (N_14225,N_11026,N_11513);
nand U14226 (N_14226,N_11515,N_11930);
nand U14227 (N_14227,N_9308,N_11771);
and U14228 (N_14228,N_9175,N_11384);
nor U14229 (N_14229,N_11319,N_9227);
nor U14230 (N_14230,N_10227,N_9983);
nor U14231 (N_14231,N_10660,N_10682);
or U14232 (N_14232,N_11275,N_9658);
nand U14233 (N_14233,N_9932,N_9928);
or U14234 (N_14234,N_11478,N_9570);
nand U14235 (N_14235,N_10828,N_10664);
nand U14236 (N_14236,N_9609,N_11274);
nor U14237 (N_14237,N_11371,N_9969);
nand U14238 (N_14238,N_9668,N_10265);
or U14239 (N_14239,N_10659,N_9081);
or U14240 (N_14240,N_9604,N_11741);
nor U14241 (N_14241,N_11989,N_11637);
nor U14242 (N_14242,N_9306,N_11776);
or U14243 (N_14243,N_11126,N_9753);
nor U14244 (N_14244,N_11221,N_9678);
and U14245 (N_14245,N_11089,N_10539);
nand U14246 (N_14246,N_9718,N_9457);
or U14247 (N_14247,N_9530,N_9207);
or U14248 (N_14248,N_9977,N_11478);
and U14249 (N_14249,N_9994,N_11218);
nand U14250 (N_14250,N_10520,N_9966);
and U14251 (N_14251,N_11926,N_11328);
nand U14252 (N_14252,N_11224,N_10077);
nor U14253 (N_14253,N_9800,N_11703);
and U14254 (N_14254,N_9495,N_10988);
or U14255 (N_14255,N_11855,N_10716);
or U14256 (N_14256,N_10436,N_11055);
nor U14257 (N_14257,N_11766,N_10052);
nand U14258 (N_14258,N_10680,N_10855);
nand U14259 (N_14259,N_9373,N_10888);
or U14260 (N_14260,N_10487,N_11965);
nor U14261 (N_14261,N_9389,N_9149);
and U14262 (N_14262,N_9869,N_10985);
xor U14263 (N_14263,N_11993,N_10005);
and U14264 (N_14264,N_11912,N_10895);
nand U14265 (N_14265,N_9310,N_10398);
or U14266 (N_14266,N_10789,N_10189);
nor U14267 (N_14267,N_11016,N_10344);
and U14268 (N_14268,N_9293,N_11165);
nor U14269 (N_14269,N_11236,N_11315);
nand U14270 (N_14270,N_10591,N_10141);
xor U14271 (N_14271,N_11691,N_9767);
nand U14272 (N_14272,N_9559,N_9122);
or U14273 (N_14273,N_11310,N_10571);
or U14274 (N_14274,N_9257,N_11159);
or U14275 (N_14275,N_10264,N_10384);
nor U14276 (N_14276,N_9863,N_11992);
nor U14277 (N_14277,N_9127,N_10363);
nand U14278 (N_14278,N_9481,N_10012);
nor U14279 (N_14279,N_11178,N_11116);
or U14280 (N_14280,N_10517,N_9380);
nor U14281 (N_14281,N_10853,N_11698);
or U14282 (N_14282,N_9518,N_11613);
or U14283 (N_14283,N_10408,N_11603);
or U14284 (N_14284,N_11811,N_10822);
or U14285 (N_14285,N_11383,N_10649);
nor U14286 (N_14286,N_11849,N_11235);
nor U14287 (N_14287,N_11689,N_10204);
xor U14288 (N_14288,N_9828,N_11018);
nand U14289 (N_14289,N_9910,N_11805);
or U14290 (N_14290,N_11781,N_10431);
and U14291 (N_14291,N_11131,N_11374);
nand U14292 (N_14292,N_10109,N_9262);
nand U14293 (N_14293,N_10020,N_9456);
nand U14294 (N_14294,N_10160,N_11428);
nand U14295 (N_14295,N_11375,N_9994);
or U14296 (N_14296,N_9668,N_11632);
nand U14297 (N_14297,N_11931,N_9311);
nand U14298 (N_14298,N_9142,N_11560);
or U14299 (N_14299,N_11178,N_9391);
and U14300 (N_14300,N_11043,N_10433);
xor U14301 (N_14301,N_9389,N_9494);
nand U14302 (N_14302,N_9190,N_10346);
nor U14303 (N_14303,N_11982,N_9459);
and U14304 (N_14304,N_9063,N_11916);
nand U14305 (N_14305,N_11979,N_9523);
and U14306 (N_14306,N_11048,N_11099);
and U14307 (N_14307,N_11591,N_10559);
or U14308 (N_14308,N_10308,N_10897);
nand U14309 (N_14309,N_10276,N_11882);
or U14310 (N_14310,N_9931,N_10616);
nand U14311 (N_14311,N_11358,N_10201);
nor U14312 (N_14312,N_11825,N_11495);
nor U14313 (N_14313,N_11510,N_11332);
nor U14314 (N_14314,N_11627,N_11476);
nor U14315 (N_14315,N_11787,N_11461);
and U14316 (N_14316,N_9183,N_11520);
and U14317 (N_14317,N_11895,N_11465);
xnor U14318 (N_14318,N_10344,N_10252);
nand U14319 (N_14319,N_11416,N_11777);
and U14320 (N_14320,N_9466,N_10461);
nor U14321 (N_14321,N_11835,N_11558);
or U14322 (N_14322,N_10149,N_9686);
or U14323 (N_14323,N_10745,N_9389);
or U14324 (N_14324,N_10961,N_10092);
or U14325 (N_14325,N_11114,N_11280);
nand U14326 (N_14326,N_11576,N_9264);
or U14327 (N_14327,N_11430,N_11802);
nor U14328 (N_14328,N_10371,N_10142);
or U14329 (N_14329,N_9455,N_11627);
nor U14330 (N_14330,N_11643,N_10730);
or U14331 (N_14331,N_9618,N_9074);
and U14332 (N_14332,N_9344,N_11952);
or U14333 (N_14333,N_9148,N_11821);
xor U14334 (N_14334,N_11165,N_10267);
and U14335 (N_14335,N_11371,N_10273);
nand U14336 (N_14336,N_9882,N_11590);
nand U14337 (N_14337,N_9011,N_11895);
nor U14338 (N_14338,N_9323,N_11682);
and U14339 (N_14339,N_9856,N_11585);
xnor U14340 (N_14340,N_11257,N_11819);
or U14341 (N_14341,N_11551,N_9190);
nor U14342 (N_14342,N_10292,N_9292);
nor U14343 (N_14343,N_11716,N_9124);
or U14344 (N_14344,N_11942,N_10407);
or U14345 (N_14345,N_9413,N_9480);
nand U14346 (N_14346,N_9832,N_11961);
and U14347 (N_14347,N_10548,N_11230);
and U14348 (N_14348,N_9497,N_9288);
or U14349 (N_14349,N_11615,N_11327);
nor U14350 (N_14350,N_10637,N_10287);
nand U14351 (N_14351,N_11904,N_9770);
and U14352 (N_14352,N_10438,N_9445);
and U14353 (N_14353,N_11940,N_9089);
or U14354 (N_14354,N_9397,N_9411);
nor U14355 (N_14355,N_10827,N_10991);
or U14356 (N_14356,N_10443,N_10484);
nand U14357 (N_14357,N_10497,N_10783);
and U14358 (N_14358,N_9434,N_10284);
or U14359 (N_14359,N_11818,N_10400);
nand U14360 (N_14360,N_10650,N_11615);
or U14361 (N_14361,N_10280,N_9410);
nand U14362 (N_14362,N_11905,N_10194);
nand U14363 (N_14363,N_10299,N_11916);
or U14364 (N_14364,N_11808,N_11948);
nand U14365 (N_14365,N_9614,N_11084);
nand U14366 (N_14366,N_10758,N_10402);
and U14367 (N_14367,N_11232,N_11997);
or U14368 (N_14368,N_9779,N_11696);
or U14369 (N_14369,N_9853,N_10038);
and U14370 (N_14370,N_10665,N_11927);
nor U14371 (N_14371,N_9379,N_9454);
nor U14372 (N_14372,N_10623,N_10700);
nor U14373 (N_14373,N_9795,N_11038);
and U14374 (N_14374,N_9360,N_9268);
or U14375 (N_14375,N_9883,N_10567);
and U14376 (N_14376,N_11544,N_10014);
nand U14377 (N_14377,N_9717,N_11942);
nor U14378 (N_14378,N_9710,N_10919);
and U14379 (N_14379,N_10097,N_10992);
or U14380 (N_14380,N_11791,N_9173);
or U14381 (N_14381,N_11418,N_9021);
and U14382 (N_14382,N_9771,N_11374);
nor U14383 (N_14383,N_9223,N_9249);
nor U14384 (N_14384,N_10891,N_9156);
nand U14385 (N_14385,N_11111,N_10900);
nor U14386 (N_14386,N_11552,N_9455);
and U14387 (N_14387,N_10830,N_10514);
or U14388 (N_14388,N_9490,N_9936);
xnor U14389 (N_14389,N_10869,N_11984);
and U14390 (N_14390,N_9437,N_9249);
nor U14391 (N_14391,N_11233,N_9387);
nor U14392 (N_14392,N_9516,N_10662);
or U14393 (N_14393,N_11613,N_11270);
nor U14394 (N_14394,N_11038,N_9699);
nor U14395 (N_14395,N_11324,N_10237);
nand U14396 (N_14396,N_9856,N_9364);
and U14397 (N_14397,N_10006,N_11815);
nor U14398 (N_14398,N_10607,N_10436);
or U14399 (N_14399,N_10592,N_9562);
nor U14400 (N_14400,N_9075,N_10021);
and U14401 (N_14401,N_10393,N_11982);
nor U14402 (N_14402,N_11699,N_10170);
and U14403 (N_14403,N_11908,N_11310);
or U14404 (N_14404,N_11994,N_9966);
nand U14405 (N_14405,N_10968,N_10937);
nor U14406 (N_14406,N_10288,N_10797);
nand U14407 (N_14407,N_11019,N_9788);
and U14408 (N_14408,N_11450,N_10451);
nor U14409 (N_14409,N_10671,N_9642);
and U14410 (N_14410,N_9573,N_10610);
or U14411 (N_14411,N_10393,N_9341);
and U14412 (N_14412,N_11319,N_9185);
or U14413 (N_14413,N_9024,N_9812);
or U14414 (N_14414,N_9293,N_11715);
or U14415 (N_14415,N_11681,N_9748);
or U14416 (N_14416,N_11988,N_10643);
or U14417 (N_14417,N_11644,N_10178);
nand U14418 (N_14418,N_9309,N_10552);
nand U14419 (N_14419,N_11798,N_9689);
nand U14420 (N_14420,N_11918,N_9974);
and U14421 (N_14421,N_10503,N_10570);
or U14422 (N_14422,N_11287,N_11859);
and U14423 (N_14423,N_9009,N_11031);
and U14424 (N_14424,N_10004,N_9564);
or U14425 (N_14425,N_10386,N_11872);
nor U14426 (N_14426,N_10795,N_10681);
or U14427 (N_14427,N_10069,N_9439);
and U14428 (N_14428,N_9795,N_9801);
and U14429 (N_14429,N_9293,N_10281);
nor U14430 (N_14430,N_10390,N_10840);
or U14431 (N_14431,N_10215,N_10511);
nand U14432 (N_14432,N_9088,N_9575);
or U14433 (N_14433,N_11837,N_10307);
or U14434 (N_14434,N_10982,N_9910);
and U14435 (N_14435,N_9310,N_11082);
xor U14436 (N_14436,N_11786,N_9150);
or U14437 (N_14437,N_10812,N_9563);
nand U14438 (N_14438,N_11333,N_10453);
nor U14439 (N_14439,N_10577,N_11595);
nand U14440 (N_14440,N_9956,N_10842);
and U14441 (N_14441,N_9286,N_9532);
nand U14442 (N_14442,N_10308,N_9838);
nor U14443 (N_14443,N_10404,N_11706);
xor U14444 (N_14444,N_10108,N_11085);
or U14445 (N_14445,N_10691,N_10677);
or U14446 (N_14446,N_11265,N_9687);
and U14447 (N_14447,N_9760,N_11924);
and U14448 (N_14448,N_10413,N_9532);
or U14449 (N_14449,N_10978,N_9715);
or U14450 (N_14450,N_11084,N_9067);
or U14451 (N_14451,N_11415,N_11313);
or U14452 (N_14452,N_10458,N_11463);
and U14453 (N_14453,N_11110,N_9590);
and U14454 (N_14454,N_10542,N_9592);
nor U14455 (N_14455,N_9751,N_11645);
or U14456 (N_14456,N_9970,N_10802);
and U14457 (N_14457,N_11149,N_9291);
or U14458 (N_14458,N_9455,N_11655);
nor U14459 (N_14459,N_10152,N_9751);
and U14460 (N_14460,N_10389,N_11824);
nor U14461 (N_14461,N_11960,N_11821);
nand U14462 (N_14462,N_10201,N_9546);
or U14463 (N_14463,N_10931,N_9126);
nand U14464 (N_14464,N_10565,N_11426);
or U14465 (N_14465,N_10737,N_10279);
or U14466 (N_14466,N_9222,N_11705);
xnor U14467 (N_14467,N_11181,N_9263);
xnor U14468 (N_14468,N_9658,N_10190);
and U14469 (N_14469,N_9416,N_11617);
and U14470 (N_14470,N_11067,N_10926);
xnor U14471 (N_14471,N_9931,N_11326);
or U14472 (N_14472,N_9124,N_11776);
nand U14473 (N_14473,N_9769,N_9520);
nand U14474 (N_14474,N_11710,N_10337);
nand U14475 (N_14475,N_9891,N_11878);
nor U14476 (N_14476,N_11894,N_9519);
or U14477 (N_14477,N_10938,N_11588);
or U14478 (N_14478,N_9564,N_11762);
nand U14479 (N_14479,N_11142,N_9637);
and U14480 (N_14480,N_11974,N_11057);
nor U14481 (N_14481,N_9960,N_10742);
nor U14482 (N_14482,N_9390,N_10219);
and U14483 (N_14483,N_11357,N_10360);
nor U14484 (N_14484,N_9769,N_10355);
and U14485 (N_14485,N_11740,N_10831);
or U14486 (N_14486,N_11260,N_9405);
or U14487 (N_14487,N_9763,N_10037);
or U14488 (N_14488,N_10217,N_10660);
nand U14489 (N_14489,N_9637,N_10891);
nand U14490 (N_14490,N_9861,N_11537);
or U14491 (N_14491,N_9933,N_11953);
nand U14492 (N_14492,N_9961,N_9402);
xnor U14493 (N_14493,N_11531,N_10604);
nor U14494 (N_14494,N_11964,N_10305);
and U14495 (N_14495,N_11190,N_10722);
xor U14496 (N_14496,N_11493,N_9221);
and U14497 (N_14497,N_10738,N_10906);
nand U14498 (N_14498,N_9541,N_9942);
or U14499 (N_14499,N_10414,N_10439);
and U14500 (N_14500,N_9981,N_9301);
and U14501 (N_14501,N_9733,N_10963);
and U14502 (N_14502,N_11105,N_11116);
nand U14503 (N_14503,N_9099,N_11511);
nor U14504 (N_14504,N_10257,N_10546);
nor U14505 (N_14505,N_9806,N_10481);
or U14506 (N_14506,N_11496,N_9971);
or U14507 (N_14507,N_9325,N_11025);
and U14508 (N_14508,N_11742,N_9079);
nand U14509 (N_14509,N_11923,N_9176);
nor U14510 (N_14510,N_10108,N_11161);
and U14511 (N_14511,N_10766,N_9003);
nand U14512 (N_14512,N_11831,N_10959);
nand U14513 (N_14513,N_10346,N_10068);
nand U14514 (N_14514,N_9251,N_11055);
nand U14515 (N_14515,N_11131,N_9327);
and U14516 (N_14516,N_9737,N_11656);
nor U14517 (N_14517,N_9176,N_11424);
or U14518 (N_14518,N_9769,N_11175);
and U14519 (N_14519,N_11082,N_9263);
nand U14520 (N_14520,N_9963,N_11807);
or U14521 (N_14521,N_9793,N_10268);
nand U14522 (N_14522,N_11271,N_11063);
or U14523 (N_14523,N_9603,N_9300);
nand U14524 (N_14524,N_10938,N_11870);
nor U14525 (N_14525,N_9186,N_10366);
and U14526 (N_14526,N_11578,N_10446);
nor U14527 (N_14527,N_10148,N_9424);
nand U14528 (N_14528,N_10949,N_11789);
nand U14529 (N_14529,N_9480,N_10391);
nor U14530 (N_14530,N_9345,N_10481);
nand U14531 (N_14531,N_11360,N_11607);
or U14532 (N_14532,N_10874,N_10636);
and U14533 (N_14533,N_9999,N_10840);
nor U14534 (N_14534,N_11300,N_10097);
nand U14535 (N_14535,N_9786,N_11277);
nand U14536 (N_14536,N_11652,N_11303);
nand U14537 (N_14537,N_9249,N_9268);
and U14538 (N_14538,N_10225,N_10917);
or U14539 (N_14539,N_10471,N_9058);
or U14540 (N_14540,N_9410,N_9243);
nor U14541 (N_14541,N_10634,N_11003);
or U14542 (N_14542,N_10420,N_11550);
or U14543 (N_14543,N_9051,N_11496);
and U14544 (N_14544,N_11297,N_11510);
or U14545 (N_14545,N_10417,N_9756);
or U14546 (N_14546,N_10705,N_10635);
nand U14547 (N_14547,N_11114,N_10664);
and U14548 (N_14548,N_10993,N_11672);
or U14549 (N_14549,N_9320,N_9474);
and U14550 (N_14550,N_10023,N_9619);
and U14551 (N_14551,N_10233,N_11157);
nor U14552 (N_14552,N_11545,N_11981);
or U14553 (N_14553,N_9564,N_9209);
nand U14554 (N_14554,N_10730,N_9300);
nor U14555 (N_14555,N_9003,N_11143);
or U14556 (N_14556,N_11330,N_9871);
or U14557 (N_14557,N_10468,N_9710);
or U14558 (N_14558,N_11493,N_11337);
nand U14559 (N_14559,N_10215,N_11766);
nand U14560 (N_14560,N_11522,N_9434);
and U14561 (N_14561,N_10634,N_9277);
and U14562 (N_14562,N_10885,N_11414);
and U14563 (N_14563,N_11407,N_11952);
xnor U14564 (N_14564,N_9241,N_10058);
nand U14565 (N_14565,N_9940,N_10394);
and U14566 (N_14566,N_11706,N_10457);
and U14567 (N_14567,N_10253,N_11551);
or U14568 (N_14568,N_10515,N_10560);
or U14569 (N_14569,N_9837,N_9032);
and U14570 (N_14570,N_11930,N_10570);
nand U14571 (N_14571,N_10702,N_9090);
nand U14572 (N_14572,N_10522,N_11541);
or U14573 (N_14573,N_9402,N_10930);
nor U14574 (N_14574,N_9309,N_10297);
nor U14575 (N_14575,N_9623,N_9542);
and U14576 (N_14576,N_10501,N_11711);
nor U14577 (N_14577,N_11340,N_11318);
nor U14578 (N_14578,N_11181,N_10404);
or U14579 (N_14579,N_9853,N_10190);
nand U14580 (N_14580,N_9566,N_9365);
nor U14581 (N_14581,N_11271,N_11192);
or U14582 (N_14582,N_11949,N_11148);
nor U14583 (N_14583,N_9308,N_9369);
nand U14584 (N_14584,N_10018,N_9221);
nor U14585 (N_14585,N_9109,N_9174);
and U14586 (N_14586,N_9204,N_11500);
and U14587 (N_14587,N_9160,N_9688);
nor U14588 (N_14588,N_9100,N_11180);
or U14589 (N_14589,N_10267,N_9202);
or U14590 (N_14590,N_9155,N_11985);
and U14591 (N_14591,N_9356,N_11067);
or U14592 (N_14592,N_9244,N_10900);
and U14593 (N_14593,N_9433,N_11540);
and U14594 (N_14594,N_9258,N_10569);
nor U14595 (N_14595,N_9028,N_11257);
or U14596 (N_14596,N_10265,N_10402);
nor U14597 (N_14597,N_11292,N_10533);
nor U14598 (N_14598,N_11715,N_9332);
and U14599 (N_14599,N_11676,N_10803);
nor U14600 (N_14600,N_10580,N_11047);
xor U14601 (N_14601,N_10860,N_11687);
nand U14602 (N_14602,N_10417,N_9979);
nand U14603 (N_14603,N_9466,N_10973);
or U14604 (N_14604,N_11470,N_10684);
nand U14605 (N_14605,N_10751,N_11711);
or U14606 (N_14606,N_11226,N_9276);
nor U14607 (N_14607,N_9584,N_11002);
xnor U14608 (N_14608,N_11354,N_9216);
nand U14609 (N_14609,N_10850,N_11484);
and U14610 (N_14610,N_9230,N_9823);
or U14611 (N_14611,N_11183,N_9033);
nand U14612 (N_14612,N_11933,N_9336);
or U14613 (N_14613,N_9433,N_10324);
or U14614 (N_14614,N_10978,N_10104);
nor U14615 (N_14615,N_11929,N_11855);
nor U14616 (N_14616,N_9015,N_10885);
nor U14617 (N_14617,N_10870,N_10070);
nand U14618 (N_14618,N_10714,N_10026);
or U14619 (N_14619,N_11934,N_11771);
nor U14620 (N_14620,N_11948,N_9387);
nand U14621 (N_14621,N_11799,N_11832);
nor U14622 (N_14622,N_9089,N_10895);
nor U14623 (N_14623,N_10068,N_10598);
or U14624 (N_14624,N_10236,N_11810);
and U14625 (N_14625,N_10288,N_11831);
nor U14626 (N_14626,N_11090,N_9007);
and U14627 (N_14627,N_10644,N_11179);
or U14628 (N_14628,N_10782,N_9668);
nor U14629 (N_14629,N_9532,N_10657);
and U14630 (N_14630,N_11684,N_9239);
nand U14631 (N_14631,N_11101,N_11715);
nand U14632 (N_14632,N_9313,N_10502);
nor U14633 (N_14633,N_11982,N_11811);
and U14634 (N_14634,N_10708,N_11248);
or U14635 (N_14635,N_9052,N_11311);
or U14636 (N_14636,N_11476,N_11135);
or U14637 (N_14637,N_9864,N_11565);
nand U14638 (N_14638,N_10654,N_11082);
or U14639 (N_14639,N_11266,N_11451);
and U14640 (N_14640,N_11467,N_11464);
nand U14641 (N_14641,N_10858,N_9523);
and U14642 (N_14642,N_10252,N_11254);
nand U14643 (N_14643,N_10507,N_10417);
nand U14644 (N_14644,N_9529,N_10153);
or U14645 (N_14645,N_10837,N_9531);
nand U14646 (N_14646,N_10304,N_10485);
xnor U14647 (N_14647,N_9583,N_10007);
nand U14648 (N_14648,N_11424,N_11560);
and U14649 (N_14649,N_11634,N_11516);
nor U14650 (N_14650,N_9333,N_10015);
nor U14651 (N_14651,N_9623,N_10655);
nand U14652 (N_14652,N_10030,N_9619);
and U14653 (N_14653,N_11545,N_11964);
nor U14654 (N_14654,N_10444,N_10999);
and U14655 (N_14655,N_9275,N_9963);
and U14656 (N_14656,N_9767,N_10588);
nand U14657 (N_14657,N_11560,N_11531);
and U14658 (N_14658,N_9463,N_9751);
and U14659 (N_14659,N_9766,N_9104);
and U14660 (N_14660,N_10203,N_11567);
or U14661 (N_14661,N_9758,N_11773);
and U14662 (N_14662,N_10659,N_10798);
nand U14663 (N_14663,N_10497,N_9806);
nand U14664 (N_14664,N_10563,N_11813);
or U14665 (N_14665,N_11028,N_11376);
nand U14666 (N_14666,N_11388,N_9989);
and U14667 (N_14667,N_11320,N_9816);
or U14668 (N_14668,N_9216,N_9080);
nand U14669 (N_14669,N_9041,N_11101);
or U14670 (N_14670,N_10238,N_9040);
nor U14671 (N_14671,N_11742,N_9442);
nor U14672 (N_14672,N_10771,N_11923);
nor U14673 (N_14673,N_11818,N_9969);
and U14674 (N_14674,N_11544,N_11065);
or U14675 (N_14675,N_9176,N_10016);
or U14676 (N_14676,N_9554,N_10505);
or U14677 (N_14677,N_10859,N_11351);
and U14678 (N_14678,N_9648,N_11598);
or U14679 (N_14679,N_10728,N_9860);
xor U14680 (N_14680,N_9759,N_9980);
or U14681 (N_14681,N_11281,N_11886);
nor U14682 (N_14682,N_9581,N_10986);
nand U14683 (N_14683,N_11071,N_11065);
nor U14684 (N_14684,N_10365,N_9404);
or U14685 (N_14685,N_9938,N_9122);
and U14686 (N_14686,N_9165,N_11948);
and U14687 (N_14687,N_11767,N_11645);
and U14688 (N_14688,N_10591,N_11500);
nand U14689 (N_14689,N_11439,N_9504);
or U14690 (N_14690,N_9889,N_9409);
or U14691 (N_14691,N_11955,N_11499);
or U14692 (N_14692,N_10741,N_9127);
or U14693 (N_14693,N_10250,N_10928);
and U14694 (N_14694,N_9041,N_11614);
or U14695 (N_14695,N_11243,N_9903);
nor U14696 (N_14696,N_9688,N_9955);
nor U14697 (N_14697,N_10163,N_9863);
or U14698 (N_14698,N_10364,N_10365);
nor U14699 (N_14699,N_11814,N_11687);
or U14700 (N_14700,N_9877,N_10394);
or U14701 (N_14701,N_11997,N_10999);
nor U14702 (N_14702,N_11824,N_10984);
nand U14703 (N_14703,N_10488,N_9368);
nor U14704 (N_14704,N_11249,N_9312);
nor U14705 (N_14705,N_9378,N_10019);
nor U14706 (N_14706,N_9887,N_10062);
nand U14707 (N_14707,N_10060,N_10681);
and U14708 (N_14708,N_11747,N_11713);
and U14709 (N_14709,N_10965,N_11093);
nand U14710 (N_14710,N_9679,N_10992);
nor U14711 (N_14711,N_10785,N_9989);
and U14712 (N_14712,N_10757,N_10506);
nand U14713 (N_14713,N_10853,N_10965);
or U14714 (N_14714,N_11751,N_11323);
nand U14715 (N_14715,N_10320,N_9644);
nor U14716 (N_14716,N_11951,N_9775);
nor U14717 (N_14717,N_10930,N_10016);
nand U14718 (N_14718,N_10494,N_11311);
nor U14719 (N_14719,N_9664,N_10952);
xnor U14720 (N_14720,N_9217,N_9552);
nand U14721 (N_14721,N_11519,N_10135);
and U14722 (N_14722,N_10365,N_9300);
nand U14723 (N_14723,N_10480,N_10437);
or U14724 (N_14724,N_10308,N_11557);
nor U14725 (N_14725,N_10880,N_10392);
and U14726 (N_14726,N_11789,N_10349);
nand U14727 (N_14727,N_11154,N_9891);
and U14728 (N_14728,N_10394,N_11325);
or U14729 (N_14729,N_10846,N_9649);
and U14730 (N_14730,N_9226,N_9749);
or U14731 (N_14731,N_10002,N_10613);
and U14732 (N_14732,N_10762,N_10355);
and U14733 (N_14733,N_11314,N_11075);
nor U14734 (N_14734,N_10862,N_11634);
and U14735 (N_14735,N_11704,N_10082);
or U14736 (N_14736,N_10999,N_10169);
or U14737 (N_14737,N_10037,N_11345);
or U14738 (N_14738,N_9200,N_11146);
nor U14739 (N_14739,N_9108,N_10320);
nor U14740 (N_14740,N_10799,N_9413);
and U14741 (N_14741,N_10019,N_10693);
xor U14742 (N_14742,N_11738,N_11765);
nand U14743 (N_14743,N_9589,N_11209);
nand U14744 (N_14744,N_10025,N_10018);
or U14745 (N_14745,N_10227,N_10816);
nor U14746 (N_14746,N_11856,N_10460);
and U14747 (N_14747,N_11426,N_11706);
and U14748 (N_14748,N_11858,N_9811);
nand U14749 (N_14749,N_9493,N_11167);
or U14750 (N_14750,N_10768,N_11680);
or U14751 (N_14751,N_9379,N_11418);
nor U14752 (N_14752,N_11763,N_9143);
xnor U14753 (N_14753,N_11482,N_9010);
nand U14754 (N_14754,N_9688,N_10764);
and U14755 (N_14755,N_11546,N_11029);
or U14756 (N_14756,N_11715,N_11671);
nand U14757 (N_14757,N_10323,N_9736);
and U14758 (N_14758,N_9978,N_10361);
or U14759 (N_14759,N_10760,N_9202);
and U14760 (N_14760,N_10169,N_10743);
nor U14761 (N_14761,N_9359,N_10551);
and U14762 (N_14762,N_10218,N_9976);
and U14763 (N_14763,N_9191,N_10815);
and U14764 (N_14764,N_11912,N_11005);
nor U14765 (N_14765,N_10972,N_9576);
nand U14766 (N_14766,N_10647,N_9099);
nor U14767 (N_14767,N_11159,N_11561);
nand U14768 (N_14768,N_11808,N_9467);
nor U14769 (N_14769,N_11000,N_9012);
nand U14770 (N_14770,N_10462,N_9470);
nand U14771 (N_14771,N_10509,N_9941);
or U14772 (N_14772,N_10086,N_10224);
and U14773 (N_14773,N_9865,N_10491);
nand U14774 (N_14774,N_9521,N_11553);
nor U14775 (N_14775,N_10965,N_11692);
and U14776 (N_14776,N_10772,N_9792);
nor U14777 (N_14777,N_10336,N_11697);
and U14778 (N_14778,N_11315,N_10688);
and U14779 (N_14779,N_11035,N_10889);
or U14780 (N_14780,N_10861,N_11696);
nor U14781 (N_14781,N_11556,N_10939);
or U14782 (N_14782,N_11948,N_10277);
and U14783 (N_14783,N_9442,N_10210);
nor U14784 (N_14784,N_9282,N_11961);
nor U14785 (N_14785,N_9715,N_11108);
nand U14786 (N_14786,N_9068,N_9441);
and U14787 (N_14787,N_11486,N_10482);
nand U14788 (N_14788,N_11136,N_11035);
or U14789 (N_14789,N_11110,N_10627);
nor U14790 (N_14790,N_10782,N_10619);
nand U14791 (N_14791,N_11619,N_10500);
nand U14792 (N_14792,N_9896,N_10291);
nor U14793 (N_14793,N_11159,N_11359);
or U14794 (N_14794,N_11080,N_11018);
and U14795 (N_14795,N_10714,N_10538);
and U14796 (N_14796,N_9436,N_11932);
and U14797 (N_14797,N_10753,N_9344);
or U14798 (N_14798,N_11792,N_10274);
or U14799 (N_14799,N_9301,N_11579);
nor U14800 (N_14800,N_11884,N_10462);
xor U14801 (N_14801,N_9395,N_11425);
xor U14802 (N_14802,N_9724,N_11575);
xnor U14803 (N_14803,N_11763,N_11542);
nand U14804 (N_14804,N_11804,N_10402);
nor U14805 (N_14805,N_11324,N_11019);
or U14806 (N_14806,N_11453,N_11705);
and U14807 (N_14807,N_11672,N_11276);
or U14808 (N_14808,N_9842,N_11676);
nor U14809 (N_14809,N_10865,N_11766);
and U14810 (N_14810,N_9444,N_9655);
or U14811 (N_14811,N_9443,N_11276);
or U14812 (N_14812,N_9487,N_9319);
nand U14813 (N_14813,N_11400,N_9056);
and U14814 (N_14814,N_9678,N_10463);
or U14815 (N_14815,N_11250,N_11159);
and U14816 (N_14816,N_11225,N_11723);
or U14817 (N_14817,N_9535,N_11179);
or U14818 (N_14818,N_10271,N_10569);
nor U14819 (N_14819,N_9440,N_10899);
nand U14820 (N_14820,N_9332,N_9346);
and U14821 (N_14821,N_9504,N_10761);
and U14822 (N_14822,N_10210,N_11947);
nand U14823 (N_14823,N_10119,N_10633);
nand U14824 (N_14824,N_10575,N_10201);
nor U14825 (N_14825,N_10234,N_9192);
and U14826 (N_14826,N_11253,N_9708);
nand U14827 (N_14827,N_10933,N_10456);
xnor U14828 (N_14828,N_11550,N_9246);
nand U14829 (N_14829,N_10485,N_10188);
nor U14830 (N_14830,N_10655,N_9706);
nor U14831 (N_14831,N_10911,N_10293);
and U14832 (N_14832,N_11412,N_11725);
nand U14833 (N_14833,N_11409,N_10326);
or U14834 (N_14834,N_11148,N_10546);
nor U14835 (N_14835,N_9857,N_11905);
nand U14836 (N_14836,N_10615,N_9288);
or U14837 (N_14837,N_9224,N_10118);
and U14838 (N_14838,N_10250,N_10469);
nor U14839 (N_14839,N_10725,N_9393);
or U14840 (N_14840,N_9422,N_10278);
nor U14841 (N_14841,N_9066,N_9811);
or U14842 (N_14842,N_9296,N_9111);
nand U14843 (N_14843,N_11284,N_11888);
and U14844 (N_14844,N_11231,N_11698);
or U14845 (N_14845,N_10327,N_9403);
or U14846 (N_14846,N_11015,N_11192);
or U14847 (N_14847,N_11520,N_11254);
nor U14848 (N_14848,N_11269,N_11230);
and U14849 (N_14849,N_9135,N_9171);
and U14850 (N_14850,N_9428,N_11696);
nand U14851 (N_14851,N_10674,N_11327);
nand U14852 (N_14852,N_11465,N_11700);
nor U14853 (N_14853,N_10159,N_10990);
and U14854 (N_14854,N_9451,N_11156);
xnor U14855 (N_14855,N_9438,N_9076);
nand U14856 (N_14856,N_11377,N_11040);
nand U14857 (N_14857,N_11721,N_9225);
nor U14858 (N_14858,N_10374,N_10542);
nand U14859 (N_14859,N_9573,N_9089);
nor U14860 (N_14860,N_11156,N_10058);
or U14861 (N_14861,N_11198,N_10742);
or U14862 (N_14862,N_9165,N_10853);
nor U14863 (N_14863,N_9286,N_11538);
or U14864 (N_14864,N_10389,N_9175);
and U14865 (N_14865,N_10429,N_10970);
or U14866 (N_14866,N_11852,N_10698);
nor U14867 (N_14867,N_9269,N_9245);
and U14868 (N_14868,N_11126,N_10057);
xnor U14869 (N_14869,N_9226,N_9230);
or U14870 (N_14870,N_9778,N_11317);
or U14871 (N_14871,N_11021,N_10924);
nand U14872 (N_14872,N_9369,N_10146);
and U14873 (N_14873,N_11935,N_11590);
nand U14874 (N_14874,N_11935,N_10254);
nand U14875 (N_14875,N_9076,N_11137);
nand U14876 (N_14876,N_9069,N_11723);
nor U14877 (N_14877,N_9254,N_9528);
xnor U14878 (N_14878,N_9748,N_11951);
and U14879 (N_14879,N_9643,N_11954);
nor U14880 (N_14880,N_10365,N_11659);
or U14881 (N_14881,N_9965,N_9646);
or U14882 (N_14882,N_9886,N_11270);
or U14883 (N_14883,N_11305,N_11753);
nor U14884 (N_14884,N_9234,N_11217);
and U14885 (N_14885,N_9856,N_10149);
nor U14886 (N_14886,N_9445,N_9235);
and U14887 (N_14887,N_11714,N_11127);
and U14888 (N_14888,N_9502,N_9874);
and U14889 (N_14889,N_9269,N_9209);
and U14890 (N_14890,N_10251,N_11200);
and U14891 (N_14891,N_11441,N_10900);
and U14892 (N_14892,N_11615,N_11229);
nor U14893 (N_14893,N_11223,N_11547);
nand U14894 (N_14894,N_11488,N_11000);
or U14895 (N_14895,N_9465,N_10464);
nor U14896 (N_14896,N_9235,N_11065);
nand U14897 (N_14897,N_10053,N_11463);
or U14898 (N_14898,N_10153,N_10453);
or U14899 (N_14899,N_10351,N_11083);
or U14900 (N_14900,N_9307,N_9705);
and U14901 (N_14901,N_11064,N_9781);
nor U14902 (N_14902,N_11552,N_11418);
xnor U14903 (N_14903,N_10853,N_11746);
nor U14904 (N_14904,N_10009,N_11034);
nand U14905 (N_14905,N_10838,N_10001);
and U14906 (N_14906,N_11777,N_11848);
nor U14907 (N_14907,N_11007,N_10746);
or U14908 (N_14908,N_9770,N_11286);
or U14909 (N_14909,N_9025,N_11655);
and U14910 (N_14910,N_9742,N_11813);
and U14911 (N_14911,N_11283,N_9604);
nor U14912 (N_14912,N_9066,N_10693);
or U14913 (N_14913,N_11833,N_11869);
nor U14914 (N_14914,N_9318,N_10322);
or U14915 (N_14915,N_11272,N_9634);
nand U14916 (N_14916,N_9253,N_11443);
nor U14917 (N_14917,N_9670,N_11479);
or U14918 (N_14918,N_9074,N_9332);
and U14919 (N_14919,N_9097,N_9113);
nor U14920 (N_14920,N_10085,N_9429);
or U14921 (N_14921,N_10888,N_10246);
or U14922 (N_14922,N_10805,N_9615);
or U14923 (N_14923,N_10507,N_9670);
xnor U14924 (N_14924,N_11806,N_11869);
or U14925 (N_14925,N_9143,N_11718);
nor U14926 (N_14926,N_9370,N_11934);
or U14927 (N_14927,N_10312,N_9636);
nor U14928 (N_14928,N_9561,N_9861);
nand U14929 (N_14929,N_10918,N_10282);
and U14930 (N_14930,N_11151,N_11508);
nor U14931 (N_14931,N_11687,N_9481);
nand U14932 (N_14932,N_11990,N_9421);
or U14933 (N_14933,N_10283,N_9050);
or U14934 (N_14934,N_10041,N_9943);
or U14935 (N_14935,N_10159,N_10940);
or U14936 (N_14936,N_11919,N_9637);
and U14937 (N_14937,N_9127,N_11444);
or U14938 (N_14938,N_9636,N_11933);
or U14939 (N_14939,N_10412,N_9029);
nand U14940 (N_14940,N_10114,N_10862);
xnor U14941 (N_14941,N_10362,N_10810);
and U14942 (N_14942,N_10075,N_9811);
or U14943 (N_14943,N_9618,N_11151);
or U14944 (N_14944,N_9333,N_11524);
or U14945 (N_14945,N_9985,N_9120);
and U14946 (N_14946,N_9196,N_10717);
and U14947 (N_14947,N_11732,N_9448);
nor U14948 (N_14948,N_10971,N_9924);
or U14949 (N_14949,N_11898,N_11876);
or U14950 (N_14950,N_11262,N_11581);
nor U14951 (N_14951,N_11515,N_9848);
nand U14952 (N_14952,N_11623,N_10789);
and U14953 (N_14953,N_10936,N_9744);
nand U14954 (N_14954,N_9848,N_10924);
or U14955 (N_14955,N_11449,N_10357);
and U14956 (N_14956,N_11516,N_9609);
nand U14957 (N_14957,N_9542,N_9439);
and U14958 (N_14958,N_11632,N_9315);
nor U14959 (N_14959,N_9568,N_9364);
or U14960 (N_14960,N_10869,N_11328);
or U14961 (N_14961,N_10127,N_11301);
nor U14962 (N_14962,N_9841,N_11368);
nor U14963 (N_14963,N_11243,N_9708);
and U14964 (N_14964,N_10338,N_11789);
or U14965 (N_14965,N_11901,N_10100);
nor U14966 (N_14966,N_9401,N_11456);
nand U14967 (N_14967,N_9206,N_9773);
or U14968 (N_14968,N_11771,N_11924);
and U14969 (N_14969,N_9275,N_10815);
nor U14970 (N_14970,N_11293,N_9897);
or U14971 (N_14971,N_9496,N_9587);
nor U14972 (N_14972,N_10411,N_9400);
nor U14973 (N_14973,N_10345,N_11753);
xnor U14974 (N_14974,N_9616,N_11265);
and U14975 (N_14975,N_10199,N_9573);
nor U14976 (N_14976,N_9016,N_11242);
nand U14977 (N_14977,N_10572,N_9630);
xnor U14978 (N_14978,N_11432,N_11174);
and U14979 (N_14979,N_11621,N_10460);
nor U14980 (N_14980,N_10690,N_10019);
xnor U14981 (N_14981,N_10062,N_10387);
or U14982 (N_14982,N_10024,N_9019);
and U14983 (N_14983,N_11638,N_10800);
nand U14984 (N_14984,N_11101,N_11723);
or U14985 (N_14985,N_10066,N_11239);
nor U14986 (N_14986,N_9164,N_9249);
and U14987 (N_14987,N_10003,N_9821);
nor U14988 (N_14988,N_11966,N_11293);
or U14989 (N_14989,N_9231,N_9406);
nand U14990 (N_14990,N_11185,N_9128);
nand U14991 (N_14991,N_9271,N_9724);
and U14992 (N_14992,N_9781,N_9847);
and U14993 (N_14993,N_11393,N_11827);
and U14994 (N_14994,N_10841,N_11722);
and U14995 (N_14995,N_9974,N_10162);
or U14996 (N_14996,N_9228,N_10212);
nor U14997 (N_14997,N_10757,N_9065);
or U14998 (N_14998,N_10736,N_10466);
or U14999 (N_14999,N_11340,N_9927);
and UO_0 (O_0,N_13508,N_13601);
nand UO_1 (O_1,N_12726,N_13185);
and UO_2 (O_2,N_13400,N_14419);
and UO_3 (O_3,N_13740,N_14175);
and UO_4 (O_4,N_12385,N_12227);
and UO_5 (O_5,N_14490,N_12874);
or UO_6 (O_6,N_13478,N_14340);
xor UO_7 (O_7,N_12959,N_14066);
nor UO_8 (O_8,N_12200,N_13383);
nand UO_9 (O_9,N_14257,N_14583);
nand UO_10 (O_10,N_14142,N_14268);
nor UO_11 (O_11,N_13916,N_13472);
nor UO_12 (O_12,N_14761,N_13694);
and UO_13 (O_13,N_12443,N_14668);
or UO_14 (O_14,N_14516,N_14284);
nor UO_15 (O_15,N_14594,N_12677);
or UO_16 (O_16,N_14520,N_14446);
or UO_17 (O_17,N_13109,N_13064);
and UO_18 (O_18,N_12649,N_12722);
and UO_19 (O_19,N_14343,N_14805);
or UO_20 (O_20,N_12226,N_12168);
or UO_21 (O_21,N_12557,N_13489);
nand UO_22 (O_22,N_13161,N_14772);
or UO_23 (O_23,N_13720,N_12803);
and UO_24 (O_24,N_12373,N_13053);
nand UO_25 (O_25,N_13116,N_14041);
or UO_26 (O_26,N_14973,N_12841);
nor UO_27 (O_27,N_14881,N_12009);
and UO_28 (O_28,N_14060,N_12580);
and UO_29 (O_29,N_14466,N_13816);
nand UO_30 (O_30,N_13594,N_13349);
nand UO_31 (O_31,N_13429,N_14991);
nor UO_32 (O_32,N_14531,N_13487);
nor UO_33 (O_33,N_14480,N_12126);
nor UO_34 (O_34,N_14487,N_14905);
or UO_35 (O_35,N_14322,N_14467);
nand UO_36 (O_36,N_12669,N_13335);
and UO_37 (O_37,N_13492,N_14997);
nand UO_38 (O_38,N_13453,N_14204);
or UO_39 (O_39,N_12053,N_12732);
and UO_40 (O_40,N_12564,N_14510);
nor UO_41 (O_41,N_13742,N_12727);
nand UO_42 (O_42,N_14471,N_13401);
and UO_43 (O_43,N_13954,N_12575);
nor UO_44 (O_44,N_14933,N_14248);
nor UO_45 (O_45,N_13074,N_14442);
and UO_46 (O_46,N_14802,N_14554);
and UO_47 (O_47,N_13680,N_12056);
or UO_48 (O_48,N_12461,N_14553);
nand UO_49 (O_49,N_13113,N_12509);
and UO_50 (O_50,N_12081,N_13577);
nand UO_51 (O_51,N_14454,N_12246);
and UO_52 (O_52,N_12869,N_13463);
nor UO_53 (O_53,N_12277,N_13094);
or UO_54 (O_54,N_14300,N_13785);
nor UO_55 (O_55,N_13348,N_12138);
or UO_56 (O_56,N_13067,N_13904);
nor UO_57 (O_57,N_14792,N_12505);
and UO_58 (O_58,N_13805,N_13768);
or UO_59 (O_59,N_14261,N_13448);
and UO_60 (O_60,N_14896,N_12272);
or UO_61 (O_61,N_12328,N_14193);
nor UO_62 (O_62,N_13485,N_14517);
nor UO_63 (O_63,N_12660,N_13329);
nand UO_64 (O_64,N_14716,N_12264);
nand UO_65 (O_65,N_13332,N_12670);
or UO_66 (O_66,N_12771,N_13422);
and UO_67 (O_67,N_13530,N_12755);
nor UO_68 (O_68,N_13264,N_12667);
xor UO_69 (O_69,N_14938,N_13043);
nand UO_70 (O_70,N_13470,N_13156);
or UO_71 (O_71,N_14366,N_14036);
xor UO_72 (O_72,N_12173,N_13419);
and UO_73 (O_73,N_13011,N_13249);
nor UO_74 (O_74,N_14230,N_12178);
nor UO_75 (O_75,N_12000,N_13208);
xnor UO_76 (O_76,N_14396,N_13174);
or UO_77 (O_77,N_14316,N_14870);
nor UO_78 (O_78,N_14711,N_13518);
or UO_79 (O_79,N_12571,N_13178);
and UO_80 (O_80,N_14379,N_14647);
nand UO_81 (O_81,N_14131,N_14281);
nand UO_82 (O_82,N_12257,N_12599);
nor UO_83 (O_83,N_13410,N_14535);
and UO_84 (O_84,N_12230,N_14106);
nand UO_85 (O_85,N_13803,N_14810);
nand UO_86 (O_86,N_14608,N_13862);
nor UO_87 (O_87,N_13793,N_12772);
and UO_88 (O_88,N_12080,N_13613);
nand UO_89 (O_89,N_12513,N_12543);
and UO_90 (O_90,N_13901,N_14470);
or UO_91 (O_91,N_14108,N_12531);
and UO_92 (O_92,N_12118,N_14122);
nor UO_93 (O_93,N_14236,N_12866);
nor UO_94 (O_94,N_13922,N_12100);
and UO_95 (O_95,N_12703,N_13093);
nor UO_96 (O_96,N_12371,N_14964);
or UO_97 (O_97,N_13034,N_14035);
nand UO_98 (O_98,N_12560,N_13750);
or UO_99 (O_99,N_14341,N_14544);
nor UO_100 (O_100,N_13950,N_14127);
nor UO_101 (O_101,N_14519,N_13173);
nor UO_102 (O_102,N_12642,N_13447);
nand UO_103 (O_103,N_13184,N_14026);
or UO_104 (O_104,N_14523,N_14542);
or UO_105 (O_105,N_13291,N_12165);
xor UO_106 (O_106,N_13960,N_13866);
or UO_107 (O_107,N_14853,N_14468);
nand UO_108 (O_108,N_14347,N_13566);
xor UO_109 (O_109,N_12838,N_13764);
or UO_110 (O_110,N_12937,N_12967);
nor UO_111 (O_111,N_14655,N_13426);
and UO_112 (O_112,N_14688,N_12343);
nor UO_113 (O_113,N_14364,N_13058);
xnor UO_114 (O_114,N_13369,N_13195);
or UO_115 (O_115,N_13341,N_13942);
or UO_116 (O_116,N_14021,N_13548);
and UO_117 (O_117,N_13851,N_12210);
or UO_118 (O_118,N_13714,N_12525);
nand UO_119 (O_119,N_14776,N_14426);
nand UO_120 (O_120,N_13236,N_13271);
nand UO_121 (O_121,N_13997,N_12068);
and UO_122 (O_122,N_12262,N_14497);
nand UO_123 (O_123,N_12457,N_12060);
or UO_124 (O_124,N_14774,N_13837);
nand UO_125 (O_125,N_13843,N_13060);
or UO_126 (O_126,N_12087,N_14430);
xor UO_127 (O_127,N_13656,N_14930);
or UO_128 (O_128,N_13819,N_12375);
and UO_129 (O_129,N_14040,N_13118);
nor UO_130 (O_130,N_13700,N_14049);
nand UO_131 (O_131,N_12673,N_13358);
nor UO_132 (O_132,N_14264,N_13936);
and UO_133 (O_133,N_13800,N_13239);
xor UO_134 (O_134,N_14047,N_13153);
or UO_135 (O_135,N_14837,N_13428);
or UO_136 (O_136,N_12406,N_14894);
nor UO_137 (O_137,N_13956,N_14725);
nor UO_138 (O_138,N_13534,N_13567);
nor UO_139 (O_139,N_14346,N_14053);
or UO_140 (O_140,N_14639,N_14765);
nor UO_141 (O_141,N_13649,N_14505);
or UO_142 (O_142,N_12043,N_13145);
and UO_143 (O_143,N_14023,N_14589);
and UO_144 (O_144,N_14694,N_12032);
nand UO_145 (O_145,N_13874,N_12347);
and UO_146 (O_146,N_14547,N_13591);
or UO_147 (O_147,N_12439,N_12256);
nand UO_148 (O_148,N_14697,N_14701);
nand UO_149 (O_149,N_14692,N_13931);
nor UO_150 (O_150,N_12931,N_12441);
xnor UO_151 (O_151,N_12867,N_12985);
or UO_152 (O_152,N_14179,N_14579);
and UO_153 (O_153,N_12573,N_13587);
nor UO_154 (O_154,N_13845,N_13664);
nand UO_155 (O_155,N_13215,N_14481);
nand UO_156 (O_156,N_13917,N_12326);
or UO_157 (O_157,N_12176,N_14390);
or UO_158 (O_158,N_13037,N_14435);
nand UO_159 (O_159,N_13861,N_12893);
nand UO_160 (O_160,N_14820,N_14581);
xnor UO_161 (O_161,N_14676,N_13023);
or UO_162 (O_162,N_14144,N_14325);
and UO_163 (O_163,N_12212,N_13085);
nor UO_164 (O_164,N_14819,N_14929);
or UO_165 (O_165,N_14491,N_14141);
or UO_166 (O_166,N_13607,N_12903);
and UO_167 (O_167,N_14158,N_13939);
or UO_168 (O_168,N_13048,N_14251);
nor UO_169 (O_169,N_14287,N_14199);
nand UO_170 (O_170,N_14840,N_13268);
nor UO_171 (O_171,N_13451,N_14643);
or UO_172 (O_172,N_13616,N_14726);
or UO_173 (O_173,N_14500,N_13375);
or UO_174 (O_174,N_12983,N_12284);
nor UO_175 (O_175,N_12036,N_12739);
nand UO_176 (O_176,N_13965,N_13540);
nor UO_177 (O_177,N_13437,N_13842);
xnor UO_178 (O_178,N_12045,N_12179);
nor UO_179 (O_179,N_13407,N_14154);
or UO_180 (O_180,N_14139,N_13600);
nor UO_181 (O_181,N_12276,N_13284);
and UO_182 (O_182,N_14094,N_12136);
nand UO_183 (O_183,N_13771,N_13985);
nand UO_184 (O_184,N_12236,N_12777);
nor UO_185 (O_185,N_14615,N_13898);
nand UO_186 (O_186,N_14641,N_14684);
or UO_187 (O_187,N_14232,N_13844);
xnor UO_188 (O_188,N_13497,N_13265);
and UO_189 (O_189,N_13026,N_14404);
nor UO_190 (O_190,N_12492,N_12533);
or UO_191 (O_191,N_12241,N_13392);
xor UO_192 (O_192,N_12940,N_13275);
or UO_193 (O_193,N_13903,N_14133);
nor UO_194 (O_194,N_13491,N_12161);
and UO_195 (O_195,N_13435,N_14514);
nor UO_196 (O_196,N_14784,N_12494);
xnor UO_197 (O_197,N_14195,N_13339);
nor UO_198 (O_198,N_12481,N_13707);
nand UO_199 (O_199,N_12871,N_12460);
nand UO_200 (O_200,N_12656,N_12684);
or UO_201 (O_201,N_12002,N_12027);
nand UO_202 (O_202,N_13233,N_13306);
nor UO_203 (O_203,N_13242,N_13498);
or UO_204 (O_204,N_12719,N_14174);
nand UO_205 (O_205,N_14999,N_13505);
and UO_206 (O_206,N_13726,N_13083);
or UO_207 (O_207,N_13780,N_14648);
nor UO_208 (O_208,N_12590,N_13370);
or UO_209 (O_209,N_14080,N_14713);
nor UO_210 (O_210,N_12380,N_13504);
nor UO_211 (O_211,N_12714,N_12381);
nand UO_212 (O_212,N_12191,N_14475);
nand UO_213 (O_213,N_12711,N_12263);
and UO_214 (O_214,N_12736,N_12828);
nand UO_215 (O_215,N_14971,N_14636);
or UO_216 (O_216,N_14767,N_12994);
nor UO_217 (O_217,N_13240,N_14890);
nand UO_218 (O_218,N_12709,N_14646);
xor UO_219 (O_219,N_13609,N_14951);
nand UO_220 (O_220,N_13499,N_13888);
nand UO_221 (O_221,N_12506,N_12405);
and UO_222 (O_222,N_14027,N_14134);
nand UO_223 (O_223,N_13692,N_14226);
nor UO_224 (O_224,N_12998,N_12142);
xnor UO_225 (O_225,N_13517,N_14223);
or UO_226 (O_226,N_14576,N_12244);
and UO_227 (O_227,N_12394,N_13608);
nand UO_228 (O_228,N_12909,N_12631);
nor UO_229 (O_229,N_12745,N_14886);
nand UO_230 (O_230,N_13519,N_13944);
nand UO_231 (O_231,N_13999,N_14085);
nand UO_232 (O_232,N_13605,N_14758);
and UO_233 (O_233,N_12540,N_13475);
nand UO_234 (O_234,N_13933,N_12744);
or UO_235 (O_235,N_13218,N_13163);
or UO_236 (O_236,N_13795,N_14897);
and UO_237 (O_237,N_14351,N_14671);
nand UO_238 (O_238,N_14869,N_13162);
and UO_239 (O_239,N_14683,N_13364);
nor UO_240 (O_240,N_12497,N_14486);
and UO_241 (O_241,N_14735,N_13635);
nor UO_242 (O_242,N_14795,N_13913);
or UO_243 (O_243,N_12929,N_13243);
nand UO_244 (O_244,N_14799,N_12872);
and UO_245 (O_245,N_13814,N_14652);
and UO_246 (O_246,N_13543,N_14062);
nand UO_247 (O_247,N_14415,N_13107);
and UO_248 (O_248,N_14729,N_12830);
or UO_249 (O_249,N_14391,N_12288);
or UO_250 (O_250,N_12616,N_13736);
nand UO_251 (O_251,N_13398,N_14348);
nand UO_252 (O_252,N_13103,N_13296);
and UO_253 (O_253,N_14588,N_14455);
and UO_254 (O_254,N_12603,N_12912);
or UO_255 (O_255,N_12435,N_12170);
nor UO_256 (O_256,N_14440,N_12362);
nand UO_257 (O_257,N_14303,N_13235);
and UO_258 (O_258,N_12942,N_13059);
and UO_259 (O_259,N_14368,N_12758);
nand UO_260 (O_260,N_12213,N_12005);
nand UO_261 (O_261,N_12201,N_14654);
nand UO_262 (O_262,N_12153,N_12993);
nand UO_263 (O_263,N_14358,N_13981);
nand UO_264 (O_264,N_13911,N_13953);
nand UO_265 (O_265,N_13586,N_13386);
nand UO_266 (O_266,N_12379,N_12717);
nor UO_267 (O_267,N_14871,N_13870);
and UO_268 (O_268,N_13778,N_13579);
nand UO_269 (O_269,N_13821,N_14690);
nor UO_270 (O_270,N_12418,N_12401);
nand UO_271 (O_271,N_12333,N_12376);
nand UO_272 (O_272,N_14184,N_13512);
nor UO_273 (O_273,N_14039,N_13687);
and UO_274 (O_274,N_14393,N_14731);
nand UO_275 (O_275,N_14914,N_14704);
nand UO_276 (O_276,N_12427,N_13248);
nor UO_277 (O_277,N_14273,N_13467);
and UO_278 (O_278,N_14533,N_14521);
nand UO_279 (O_279,N_14902,N_12408);
or UO_280 (O_280,N_14329,N_13886);
or UO_281 (O_281,N_13295,N_14425);
nand UO_282 (O_282,N_12663,N_13998);
or UO_283 (O_283,N_13310,N_14986);
nor UO_284 (O_284,N_14388,N_14022);
or UO_285 (O_285,N_13142,N_14278);
or UO_286 (O_286,N_12521,N_13996);
and UO_287 (O_287,N_12555,N_12860);
nand UO_288 (O_288,N_14687,N_13387);
nor UO_289 (O_289,N_14384,N_14561);
or UO_290 (O_290,N_13990,N_12955);
xor UO_291 (O_291,N_14374,N_12747);
nor UO_292 (O_292,N_13979,N_13167);
nor UO_293 (O_293,N_12514,N_14317);
nand UO_294 (O_294,N_12280,N_14186);
or UO_295 (O_295,N_14335,N_14715);
or UO_296 (O_296,N_14167,N_13462);
nand UO_297 (O_297,N_14823,N_14605);
nand UO_298 (O_298,N_13501,N_12857);
and UO_299 (O_299,N_13257,N_13464);
and UO_300 (O_300,N_14843,N_13183);
and UO_301 (O_301,N_12339,N_13217);
nand UO_302 (O_302,N_14439,N_13188);
nand UO_303 (O_303,N_12639,N_14734);
nand UO_304 (O_304,N_12643,N_14038);
nand UO_305 (O_305,N_14365,N_14436);
nand UO_306 (O_306,N_12329,N_12437);
nor UO_307 (O_307,N_12104,N_13413);
and UO_308 (O_308,N_13164,N_13147);
and UO_309 (O_309,N_13572,N_14740);
nor UO_310 (O_310,N_13958,N_12250);
and UO_311 (O_311,N_13802,N_12655);
and UO_312 (O_312,N_13787,N_12067);
nand UO_313 (O_313,N_14188,N_14441);
nand UO_314 (O_314,N_14105,N_12783);
or UO_315 (O_315,N_14925,N_13820);
or UO_316 (O_316,N_13513,N_13791);
nand UO_317 (O_317,N_14698,N_13158);
or UO_318 (O_318,N_12614,N_13896);
and UO_319 (O_319,N_12785,N_14507);
or UO_320 (O_320,N_12342,N_13561);
nand UO_321 (O_321,N_13166,N_12957);
or UO_322 (O_322,N_12410,N_14798);
xor UO_323 (O_323,N_12759,N_12735);
nor UO_324 (O_324,N_12977,N_14791);
nand UO_325 (O_325,N_12944,N_12778);
nand UO_326 (O_326,N_13366,N_14363);
nor UO_327 (O_327,N_14912,N_14399);
or UO_328 (O_328,N_12799,N_14781);
xnor UO_329 (O_329,N_13385,N_12354);
and UO_330 (O_330,N_13100,N_12470);
or UO_331 (O_331,N_12116,N_13697);
nor UO_332 (O_332,N_13266,N_14292);
nor UO_333 (O_333,N_12287,N_14889);
nand UO_334 (O_334,N_14246,N_12887);
or UO_335 (O_335,N_14756,N_13945);
nor UO_336 (O_336,N_12878,N_12600);
and UO_337 (O_337,N_12355,N_13938);
nor UO_338 (O_338,N_12834,N_12050);
or UO_339 (O_339,N_14849,N_13495);
nand UO_340 (O_340,N_12148,N_14460);
and UO_341 (O_341,N_12928,N_12038);
or UO_342 (O_342,N_12596,N_14445);
and UO_343 (O_343,N_12240,N_14686);
or UO_344 (O_344,N_14201,N_12751);
and UO_345 (O_345,N_14631,N_12692);
and UO_346 (O_346,N_14736,N_13054);
nand UO_347 (O_347,N_13086,N_12242);
nand UO_348 (O_348,N_12987,N_13568);
nand UO_349 (O_349,N_14738,N_12042);
or UO_350 (O_350,N_14679,N_13947);
nor UO_351 (O_351,N_12552,N_14381);
nand UO_352 (O_352,N_12279,N_13927);
and UO_353 (O_353,N_12905,N_12659);
nand UO_354 (O_354,N_12260,N_13702);
nand UO_355 (O_355,N_12760,N_13671);
nor UO_356 (O_356,N_14337,N_12247);
nor UO_357 (O_357,N_13804,N_12364);
nor UO_358 (O_358,N_13294,N_12473);
and UO_359 (O_359,N_13441,N_13450);
nor UO_360 (O_360,N_12205,N_12197);
nand UO_361 (O_361,N_14113,N_13655);
nor UO_362 (O_362,N_12044,N_14276);
nand UO_363 (O_363,N_12224,N_12054);
or UO_364 (O_364,N_13432,N_12147);
nand UO_365 (O_365,N_12255,N_12899);
nand UO_366 (O_366,N_14623,N_13779);
and UO_367 (O_367,N_13615,N_14800);
or UO_368 (O_368,N_12693,N_12723);
or UO_369 (O_369,N_13891,N_14259);
or UO_370 (O_370,N_14007,N_14543);
xnor UO_371 (O_371,N_12423,N_14691);
nand UO_372 (O_372,N_14386,N_12465);
nor UO_373 (O_373,N_12559,N_12298);
nand UO_374 (O_374,N_13703,N_13932);
or UO_375 (O_375,N_12843,N_12119);
or UO_376 (O_376,N_13200,N_14006);
nand UO_377 (O_377,N_12487,N_14985);
or UO_378 (O_378,N_12071,N_13810);
and UO_379 (O_379,N_14045,N_12243);
or UO_380 (O_380,N_14663,N_14147);
and UO_381 (O_381,N_12661,N_12793);
xor UO_382 (O_382,N_14712,N_13289);
nor UO_383 (O_383,N_14002,N_12219);
or UO_384 (O_384,N_14383,N_13777);
and UO_385 (O_385,N_12795,N_14747);
or UO_386 (O_386,N_13123,N_12110);
or UO_387 (O_387,N_13095,N_13262);
nand UO_388 (O_388,N_13313,N_12382);
and UO_389 (O_389,N_13739,N_14089);
or UO_390 (O_390,N_13075,N_14954);
nand UO_391 (O_391,N_12077,N_13807);
nand UO_392 (O_392,N_12203,N_12416);
and UO_393 (O_393,N_12627,N_13603);
or UO_394 (O_394,N_14827,N_14478);
or UO_395 (O_395,N_13368,N_13974);
nor UO_396 (O_396,N_13005,N_14307);
or UO_397 (O_397,N_13893,N_12891);
nand UO_398 (O_398,N_13693,N_13550);
nand UO_399 (O_399,N_14215,N_13602);
or UO_400 (O_400,N_14857,N_13066);
xor UO_401 (O_401,N_14220,N_13670);
or UO_402 (O_402,N_12155,N_14005);
nand UO_403 (O_403,N_13957,N_12705);
nand UO_404 (O_404,N_13277,N_12906);
nor UO_405 (O_405,N_12114,N_12158);
nand UO_406 (O_406,N_12062,N_13246);
nor UO_407 (O_407,N_14197,N_13225);
or UO_408 (O_408,N_14557,N_13770);
or UO_409 (O_409,N_12344,N_13120);
nor UO_410 (O_410,N_13300,N_13651);
nand UO_411 (O_411,N_13399,N_14610);
or UO_412 (O_412,N_13000,N_14330);
and UO_413 (O_413,N_13592,N_12628);
nor UO_414 (O_414,N_12558,N_13897);
or UO_415 (O_415,N_13376,N_13772);
nand UO_416 (O_416,N_13824,N_12391);
nand UO_417 (O_417,N_14670,N_14666);
and UO_418 (O_418,N_14067,N_13681);
and UO_419 (O_419,N_14262,N_14550);
nor UO_420 (O_420,N_12489,N_14515);
and UO_421 (O_421,N_13630,N_13102);
and UO_422 (O_422,N_14214,N_13551);
and UO_423 (O_423,N_12716,N_14082);
or UO_424 (O_424,N_12790,N_13180);
and UO_425 (O_425,N_12051,N_12292);
nor UO_426 (O_426,N_12794,N_13261);
nand UO_427 (O_427,N_13612,N_12327);
nand UO_428 (O_428,N_12432,N_13654);
or UO_429 (O_429,N_14096,N_14757);
nor UO_430 (O_430,N_13207,N_13055);
and UO_431 (O_431,N_12688,N_13506);
and UO_432 (O_432,N_12098,N_14057);
or UO_433 (O_433,N_14656,N_13659);
nor UO_434 (O_434,N_12082,N_14888);
nor UO_435 (O_435,N_13558,N_13536);
nand UO_436 (O_436,N_14129,N_14077);
nand UO_437 (O_437,N_13645,N_14995);
nand UO_438 (O_438,N_13080,N_12637);
nand UO_439 (O_439,N_12006,N_13646);
nor UO_440 (O_440,N_14242,N_13767);
nand UO_441 (O_441,N_12577,N_14218);
and UO_442 (O_442,N_14593,N_12935);
or UO_443 (O_443,N_14956,N_14224);
and UO_444 (O_444,N_13581,N_12356);
nand UO_445 (O_445,N_13863,N_14875);
and UO_446 (O_446,N_14739,N_13553);
nor UO_447 (O_447,N_13781,N_13696);
nor UO_448 (O_448,N_13042,N_14046);
nand UO_449 (O_449,N_12650,N_12781);
nand UO_450 (O_450,N_13869,N_12295);
nand UO_451 (O_451,N_14482,N_14402);
or UO_452 (O_452,N_13477,N_14372);
nor UO_453 (O_453,N_12107,N_13347);
nor UO_454 (O_454,N_14707,N_12387);
nor UO_455 (O_455,N_14586,N_14311);
nor UO_456 (O_456,N_12207,N_14858);
and UO_457 (O_457,N_13232,N_14209);
or UO_458 (O_458,N_13502,N_12096);
nor UO_459 (O_459,N_14097,N_12169);
or UO_460 (O_460,N_12787,N_13854);
and UO_461 (O_461,N_14042,N_13827);
or UO_462 (O_462,N_13117,N_14164);
nor UO_463 (O_463,N_12598,N_14314);
or UO_464 (O_464,N_12947,N_13087);
and UO_465 (O_465,N_12145,N_12945);
xnor UO_466 (O_466,N_14653,N_14528);
or UO_467 (O_467,N_13730,N_14710);
xor UO_468 (O_468,N_13391,N_14008);
and UO_469 (O_469,N_12109,N_14649);
or UO_470 (O_470,N_12039,N_12350);
nor UO_471 (O_471,N_13483,N_13624);
nand UO_472 (O_472,N_13878,N_13639);
or UO_473 (O_473,N_14153,N_12562);
nand UO_474 (O_474,N_13476,N_13937);
nor UO_475 (O_475,N_13390,N_12018);
and UO_476 (O_476,N_14941,N_12607);
or UO_477 (O_477,N_12971,N_12517);
nand UO_478 (O_478,N_14103,N_13443);
and UO_479 (O_479,N_13454,N_12166);
or UO_480 (O_480,N_14948,N_13292);
nand UO_481 (O_481,N_13662,N_12784);
nand UO_482 (O_482,N_14068,N_14614);
nand UO_483 (O_483,N_14650,N_13337);
nand UO_484 (O_484,N_14705,N_13830);
nor UO_485 (O_485,N_12800,N_13350);
and UO_486 (O_486,N_12337,N_14009);
and UO_487 (O_487,N_13713,N_13663);
and UO_488 (O_488,N_14783,N_14887);
and UO_489 (O_489,N_14872,N_14422);
nand UO_490 (O_490,N_12812,N_14969);
and UO_491 (O_491,N_14968,N_13509);
nor UO_492 (O_492,N_14024,N_13856);
and UO_493 (O_493,N_13411,N_12933);
nor UO_494 (O_494,N_13675,N_13983);
or UO_495 (O_495,N_12398,N_13748);
and UO_496 (O_496,N_14350,N_12992);
nor UO_497 (O_497,N_12613,N_14847);
nor UO_498 (O_498,N_13395,N_12188);
nor UO_499 (O_499,N_14534,N_14779);
and UO_500 (O_500,N_14635,N_12234);
and UO_501 (O_501,N_14228,N_13440);
nand UO_502 (O_502,N_12697,N_12503);
or UO_503 (O_503,N_12454,N_13077);
xor UO_504 (O_504,N_13970,N_13461);
or UO_505 (O_505,N_14745,N_12402);
or UO_506 (O_506,N_12816,N_12676);
nand UO_507 (O_507,N_13338,N_12894);
or UO_508 (O_508,N_13220,N_13542);
and UO_509 (O_509,N_13653,N_12261);
nor UO_510 (O_510,N_13007,N_14908);
or UO_511 (O_511,N_12130,N_14258);
nor UO_512 (O_512,N_13421,N_12433);
nand UO_513 (O_513,N_13811,N_13204);
xor UO_514 (O_514,N_14616,N_14825);
nor UO_515 (O_515,N_14574,N_12882);
or UO_516 (O_516,N_12445,N_14157);
nor UO_517 (O_517,N_13929,N_14862);
nor UO_518 (O_518,N_14904,N_13001);
and UO_519 (O_519,N_13761,N_14892);
nand UO_520 (O_520,N_13797,N_14659);
and UO_521 (O_521,N_13589,N_12282);
nor UO_522 (O_522,N_13479,N_12835);
nand UO_523 (O_523,N_14634,N_14293);
nor UO_524 (O_524,N_14879,N_14861);
nor UO_525 (O_525,N_14628,N_13210);
or UO_526 (O_526,N_14876,N_14052);
nand UO_527 (O_527,N_13588,N_14205);
or UO_528 (O_528,N_12694,N_13179);
and UO_529 (O_529,N_12647,N_13324);
nor UO_530 (O_530,N_14953,N_13241);
or UO_531 (O_531,N_12567,N_13144);
nor UO_532 (O_532,N_12546,N_12753);
nand UO_533 (O_533,N_13885,N_14187);
nor UO_534 (O_534,N_12544,N_12464);
and UO_535 (O_535,N_14434,N_12831);
or UO_536 (O_536,N_13331,N_14824);
nand UO_537 (O_537,N_13480,N_14667);
and UO_538 (O_538,N_14423,N_13170);
and UO_539 (O_539,N_13297,N_14746);
and UO_540 (O_540,N_12490,N_14560);
nand UO_541 (O_541,N_14485,N_13621);
and UO_542 (O_542,N_12273,N_14416);
nand UO_543 (O_543,N_13444,N_13151);
nor UO_544 (O_544,N_13890,N_12491);
nor UO_545 (O_545,N_12315,N_12388);
nor UO_546 (O_546,N_13190,N_14200);
nand UO_547 (O_547,N_12780,N_13424);
xnor UO_548 (O_548,N_12725,N_13755);
or UO_549 (O_549,N_13127,N_12156);
nor UO_550 (O_550,N_13817,N_14702);
nor UO_551 (O_551,N_14398,N_14360);
and UO_552 (O_552,N_13719,N_12017);
and UO_553 (O_553,N_14181,N_13209);
nand UO_554 (O_554,N_13667,N_13027);
nor UO_555 (O_555,N_14816,N_14112);
nor UO_556 (O_556,N_12908,N_13689);
nor UO_557 (O_557,N_13633,N_12442);
or UO_558 (O_558,N_12696,N_12357);
or UO_559 (O_559,N_13643,N_12604);
and UO_560 (O_560,N_13315,N_12099);
xor UO_561 (O_561,N_12447,N_14163);
or UO_562 (O_562,N_14728,N_14575);
nand UO_563 (O_563,N_12591,N_14371);
nand UO_564 (O_564,N_13063,N_12073);
nor UO_565 (O_565,N_14165,N_12845);
nor UO_566 (O_566,N_12349,N_12296);
and UO_567 (O_567,N_14484,N_13871);
and UO_568 (O_568,N_13484,N_12449);
xnor UO_569 (O_569,N_12782,N_14462);
nand UO_570 (O_570,N_12302,N_14238);
or UO_571 (O_571,N_13177,N_13333);
or UO_572 (O_572,N_12766,N_12254);
nand UO_573 (O_573,N_14289,N_12952);
nor UO_574 (O_574,N_14962,N_12563);
or UO_575 (O_575,N_14945,N_14952);
or UO_576 (O_576,N_13914,N_13794);
or UO_577 (O_577,N_12680,N_12029);
or UO_578 (O_578,N_12713,N_13101);
or UO_579 (O_579,N_12047,N_13019);
xor UO_580 (O_580,N_12589,N_12475);
and UO_581 (O_581,N_13836,N_12536);
or UO_582 (O_582,N_12022,N_12369);
and UO_583 (O_583,N_12194,N_14506);
and UO_584 (O_584,N_14864,N_12761);
nand UO_585 (O_585,N_13528,N_14362);
or UO_586 (O_586,N_13815,N_12938);
nand UO_587 (O_587,N_12426,N_12063);
or UO_588 (O_588,N_13507,N_13557);
nand UO_589 (O_589,N_12779,N_13674);
or UO_590 (O_590,N_14940,N_14766);
nand UO_591 (O_591,N_12728,N_13614);
nor UO_592 (O_592,N_12704,N_13971);
or UO_593 (O_593,N_14540,N_12707);
nor UO_594 (O_594,N_14240,N_12979);
or UO_595 (O_595,N_12896,N_14695);
or UO_596 (O_596,N_12174,N_12710);
and UO_597 (O_597,N_14935,N_14806);
nand UO_598 (O_598,N_12184,N_14277);
or UO_599 (O_599,N_13786,N_12595);
and UO_600 (O_600,N_12500,N_12646);
or UO_601 (O_601,N_14095,N_13039);
nand UO_602 (O_602,N_14562,N_12059);
and UO_603 (O_603,N_13318,N_14611);
or UO_604 (O_604,N_12682,N_12877);
or UO_605 (O_605,N_12910,N_12113);
nor UO_606 (O_606,N_14380,N_12982);
nor UO_607 (O_607,N_13988,N_12004);
or UO_608 (O_608,N_13160,N_13330);
or UO_609 (O_609,N_13909,N_12367);
or UO_610 (O_610,N_12496,N_12448);
and UO_611 (O_611,N_14015,N_14247);
and UO_612 (O_612,N_12175,N_13013);
and UO_613 (O_613,N_12915,N_14974);
nand UO_614 (O_614,N_12537,N_13855);
and UO_615 (O_615,N_12876,N_13731);
nor UO_616 (O_616,N_14432,N_13481);
nor UO_617 (O_617,N_12888,N_12654);
nand UO_618 (O_618,N_14294,N_12055);
nor UO_619 (O_619,N_12664,N_12917);
and UO_620 (O_620,N_13935,N_12995);
or UO_621 (O_621,N_14111,N_12024);
or UO_622 (O_622,N_14996,N_14793);
xor UO_623 (O_623,N_12314,N_14936);
and UO_624 (O_624,N_14458,N_12545);
and UO_625 (O_625,N_12615,N_12958);
nand UO_626 (O_626,N_13831,N_14489);
nor UO_627 (O_627,N_14310,N_13322);
nor UO_628 (O_628,N_13991,N_12392);
and UO_629 (O_629,N_13171,N_12844);
nor UO_630 (O_630,N_12765,N_12875);
nand UO_631 (O_631,N_12702,N_12088);
nand UO_632 (O_632,N_12786,N_14272);
nand UO_633 (O_633,N_13915,N_12214);
and UO_634 (O_634,N_12415,N_14034);
nor UO_635 (O_635,N_13631,N_13022);
nand UO_636 (O_636,N_12927,N_14966);
and UO_637 (O_637,N_12085,N_12608);
nand UO_638 (O_638,N_14385,N_12346);
and UO_639 (O_639,N_13418,N_13606);
nand UO_640 (O_640,N_14877,N_13446);
nand UO_641 (O_641,N_14651,N_14114);
or UO_642 (O_642,N_12934,N_13743);
nand UO_643 (O_643,N_12281,N_14509);
nand UO_644 (O_644,N_13282,N_14620);
and UO_645 (O_645,N_12515,N_14998);
and UO_646 (O_646,N_12417,N_14504);
or UO_647 (O_647,N_13115,N_13255);
and UO_648 (O_648,N_14219,N_13883);
or UO_649 (O_649,N_12320,N_13425);
xnor UO_650 (O_650,N_13363,N_13423);
and UO_651 (O_651,N_12960,N_13584);
or UO_652 (O_652,N_12969,N_14090);
or UO_653 (O_653,N_13197,N_13049);
nand UO_654 (O_654,N_13666,N_12671);
or UO_655 (O_655,N_12507,N_12274);
nor UO_656 (O_656,N_13925,N_14444);
or UO_657 (O_657,N_13850,N_12269);
and UO_658 (O_658,N_12037,N_12268);
xnor UO_659 (O_659,N_12335,N_14602);
nand UO_660 (O_660,N_13202,N_12101);
and UO_661 (O_661,N_13216,N_14963);
or UO_662 (O_662,N_14312,N_12079);
nand UO_663 (O_663,N_12954,N_12012);
nor UO_664 (O_664,N_14183,N_13076);
or UO_665 (O_665,N_12420,N_12832);
or UO_666 (O_666,N_14477,N_12127);
and UO_667 (O_667,N_12078,N_12820);
nor UO_668 (O_668,N_13525,N_13445);
nand UO_669 (O_669,N_13134,N_12015);
and UO_670 (O_670,N_12294,N_12019);
nor UO_671 (O_671,N_12996,N_14582);
and UO_672 (O_672,N_13038,N_12978);
nand UO_673 (O_673,N_14770,N_14555);
and UO_674 (O_674,N_14375,N_14569);
nand UO_675 (O_675,N_12547,N_14749);
xor UO_676 (O_676,N_13575,N_12452);
nand UO_677 (O_677,N_14541,N_12825);
or UO_678 (O_678,N_14148,N_13014);
or UO_679 (O_679,N_12499,N_14092);
nor UO_680 (O_680,N_14189,N_14866);
xnor UO_681 (O_681,N_13751,N_14429);
and UO_682 (O_682,N_14304,N_13154);
and UO_683 (O_683,N_13279,N_12228);
and UO_684 (O_684,N_12626,N_12084);
and UO_685 (O_685,N_12290,N_14797);
or UO_686 (O_686,N_13175,N_14156);
nor UO_687 (O_687,N_13046,N_12400);
nor UO_688 (O_688,N_14627,N_12411);
or UO_689 (O_689,N_14173,N_14661);
or UO_690 (O_690,N_12132,N_13303);
or UO_691 (O_691,N_14916,N_13775);
nor UO_692 (O_692,N_12146,N_12115);
or UO_693 (O_693,N_12623,N_13493);
nand UO_694 (O_694,N_14678,N_14672);
nand UO_695 (O_695,N_12149,N_13879);
and UO_696 (O_696,N_13968,N_12007);
or UO_697 (O_697,N_12516,N_14059);
or UO_698 (O_698,N_14658,N_12363);
or UO_699 (O_699,N_13471,N_14978);
or UO_700 (O_700,N_14400,N_14269);
and UO_701 (O_701,N_14091,N_12121);
or UO_702 (O_702,N_13756,N_14961);
or UO_703 (O_703,N_13286,N_13826);
nor UO_704 (O_704,N_12629,N_12466);
nor UO_705 (O_705,N_13222,N_13230);
nor UO_706 (O_706,N_12592,N_13378);
and UO_707 (O_707,N_14830,N_12477);
nor UO_708 (O_708,N_14580,N_13377);
xor UO_709 (O_709,N_14891,N_13884);
or UO_710 (O_710,N_12202,N_13882);
or UO_711 (O_711,N_14377,N_14882);
nor UO_712 (O_712,N_13353,N_13902);
and UO_713 (O_713,N_14043,N_14920);
nor UO_714 (O_714,N_13978,N_14578);
or UO_715 (O_715,N_12943,N_12579);
and UO_716 (O_716,N_12897,N_13486);
nand UO_717 (O_717,N_13365,N_14609);
nand UO_718 (O_718,N_13907,N_13533);
xnor UO_719 (O_719,N_12440,N_13808);
nand UO_720 (O_720,N_13140,N_13585);
nor UO_721 (O_721,N_13618,N_12808);
and UO_722 (O_722,N_13848,N_12640);
and UO_723 (O_723,N_12805,N_13047);
or UO_724 (O_724,N_13361,N_12283);
or UO_725 (O_725,N_13964,N_13698);
and UO_726 (O_726,N_12570,N_13009);
or UO_727 (O_727,N_12021,N_14984);
nand UO_728 (O_728,N_14548,N_12472);
nand UO_729 (O_729,N_14321,N_14016);
nand UO_730 (O_730,N_12890,N_14000);
or UO_731 (O_731,N_14075,N_14135);
nand UO_732 (O_732,N_14832,N_13521);
nor UO_733 (O_733,N_12948,N_13090);
nor UO_734 (O_734,N_14202,N_12819);
nand UO_735 (O_735,N_13072,N_14977);
nor UO_736 (O_736,N_13404,N_14677);
nand UO_737 (O_737,N_12699,N_14983);
or UO_738 (O_738,N_13473,N_14178);
or UO_739 (O_739,N_12013,N_14570);
and UO_740 (O_740,N_14789,N_14433);
nor UO_741 (O_741,N_13632,N_14566);
or UO_742 (O_742,N_14191,N_12980);
nand UO_743 (O_743,N_12455,N_12583);
or UO_744 (O_744,N_14498,N_12403);
and UO_745 (O_745,N_14353,N_14527);
and UO_746 (O_746,N_13789,N_14170);
nand UO_747 (O_747,N_14545,N_13229);
or UO_748 (O_748,N_12431,N_14706);
nand UO_749 (O_749,N_13371,N_12941);
nand UO_750 (O_750,N_12253,N_12066);
nor UO_751 (O_751,N_12767,N_13057);
nand UO_752 (O_752,N_13695,N_14235);
nor UO_753 (O_753,N_14093,N_14612);
nor UO_754 (O_754,N_13198,N_12189);
xor UO_755 (O_755,N_14965,N_14010);
nor UO_756 (O_756,N_12518,N_12824);
nand UO_757 (O_757,N_12456,N_13343);
and UO_758 (O_758,N_12361,N_12569);
nand UO_759 (O_759,N_13910,N_13346);
or UO_760 (O_760,N_12706,N_13766);
and UO_761 (O_761,N_13955,N_13625);
nand UO_762 (O_762,N_13912,N_12990);
nor UO_763 (O_763,N_14033,N_13619);
nand UO_764 (O_764,N_14055,N_14856);
nor UO_765 (O_765,N_12868,N_14003);
nand UO_766 (O_766,N_13565,N_12129);
nor UO_767 (O_767,N_12209,N_13833);
nand UO_768 (O_768,N_14502,N_14937);
nand UO_769 (O_769,N_14564,N_13710);
nand UO_770 (O_770,N_13427,N_14567);
or UO_771 (O_771,N_12386,N_14417);
nand UO_772 (O_772,N_13071,N_13254);
and UO_773 (O_773,N_12167,N_14742);
xor UO_774 (O_774,N_12069,N_12192);
nand UO_775 (O_775,N_14821,N_12864);
nand UO_776 (O_776,N_14839,N_14291);
nand UO_777 (O_777,N_12792,N_13628);
nand UO_778 (O_778,N_12511,N_14116);
nor UO_779 (O_779,N_14143,N_14285);
nand UO_780 (O_780,N_14539,N_13003);
and UO_781 (O_781,N_14483,N_12186);
xor UO_782 (O_782,N_14140,N_14884);
or UO_783 (O_783,N_13949,N_14622);
and UO_784 (O_784,N_14525,N_12904);
nand UO_785 (O_785,N_13984,N_14048);
nand UO_786 (O_786,N_14804,N_14993);
and UO_787 (O_787,N_14336,N_13665);
and UO_788 (O_788,N_14459,N_13760);
nand UO_789 (O_789,N_14573,N_14333);
nand UO_790 (O_790,N_14079,N_12665);
nor UO_791 (O_791,N_12317,N_13706);
nand UO_792 (O_792,N_14600,N_13203);
and UO_793 (O_793,N_13420,N_12072);
nand UO_794 (O_794,N_14982,N_12923);
and UO_795 (O_795,N_13868,N_14414);
and UO_796 (O_796,N_12675,N_12150);
or UO_797 (O_797,N_14326,N_14780);
and UO_798 (O_798,N_12715,N_12479);
or UO_799 (O_799,N_12862,N_14376);
nor UO_800 (O_800,N_13205,N_13576);
or UO_801 (O_801,N_12731,N_12421);
nand UO_802 (O_802,N_13281,N_13012);
nor UO_803 (O_803,N_14645,N_13564);
nor UO_804 (O_804,N_13677,N_14980);
xnor UO_805 (O_805,N_13835,N_13157);
nand UO_806 (O_806,N_12348,N_12397);
or UO_807 (O_807,N_14878,N_13627);
nor UO_808 (O_808,N_12097,N_12806);
or UO_809 (O_809,N_13834,N_12687);
nand UO_810 (O_810,N_12164,N_13309);
nor UO_811 (O_811,N_13288,N_12467);
nor UO_812 (O_812,N_12572,N_14771);
nand UO_813 (O_813,N_12028,N_12809);
or UO_814 (O_814,N_14124,N_14401);
and UO_815 (O_815,N_12316,N_13769);
nor UO_816 (O_816,N_14813,N_12484);
and UO_817 (O_817,N_14743,N_12483);
or UO_818 (O_818,N_12873,N_12094);
nand UO_819 (O_819,N_12459,N_14762);
or UO_820 (O_820,N_14243,N_12309);
and UO_821 (O_821,N_12645,N_14473);
or UO_822 (O_822,N_12360,N_13078);
nand UO_823 (O_823,N_12574,N_12691);
xor UO_824 (O_824,N_12565,N_13788);
nand UO_825 (O_825,N_14412,N_13029);
nand UO_826 (O_826,N_13299,N_14182);
or UO_827 (O_827,N_12622,N_14513);
or UO_828 (O_828,N_13244,N_12925);
and UO_829 (O_829,N_13524,N_12690);
or UO_830 (O_830,N_13159,N_14718);
nand UO_831 (O_831,N_14286,N_12474);
or UO_832 (O_832,N_14835,N_14822);
nand UO_833 (O_833,N_12249,N_12404);
nand UO_834 (O_834,N_12504,N_14029);
xnor UO_835 (O_835,N_13818,N_13717);
nand UO_836 (O_836,N_12389,N_13017);
xnor UO_837 (O_837,N_13276,N_14254);
or UO_838 (O_838,N_12601,N_12738);
and UO_839 (O_839,N_13930,N_13622);
and UO_840 (O_840,N_13599,N_14464);
or UO_841 (O_841,N_14606,N_14120);
and UO_842 (O_842,N_13563,N_13832);
and UO_843 (O_843,N_12252,N_13373);
or UO_844 (O_844,N_12974,N_12542);
nor UO_845 (O_845,N_14865,N_12453);
nor UO_846 (O_846,N_14549,N_14596);
nor UO_847 (O_847,N_14947,N_13596);
and UO_848 (O_848,N_14449,N_14270);
nor UO_849 (O_849,N_14838,N_12493);
nor UO_850 (O_850,N_12089,N_12076);
and UO_851 (O_851,N_12788,N_12151);
or UO_852 (O_852,N_13881,N_13033);
nor UO_853 (O_853,N_14076,N_13774);
nor UO_854 (O_854,N_12217,N_14102);
nand UO_855 (O_855,N_13298,N_12303);
nand UO_856 (O_856,N_12424,N_12522);
nand UO_857 (O_857,N_13194,N_13723);
nand UO_858 (O_858,N_13040,N_14512);
or UO_859 (O_859,N_14298,N_14975);
nor UO_860 (O_860,N_13908,N_12856);
or UO_861 (O_861,N_14976,N_12962);
and UO_862 (O_862,N_12235,N_13214);
nand UO_863 (O_863,N_14395,N_12366);
nor UO_864 (O_864,N_12351,N_14913);
and UO_865 (O_865,N_12729,N_12413);
nor UO_866 (O_866,N_13516,N_12251);
or UO_867 (O_867,N_14488,N_13384);
and UO_868 (O_868,N_14241,N_14944);
nand UO_869 (O_869,N_12981,N_12332);
and UO_870 (O_870,N_13133,N_13578);
nor UO_871 (O_871,N_14411,N_12539);
or UO_872 (O_872,N_12134,N_12434);
xnor UO_873 (O_873,N_14722,N_14216);
and UO_874 (O_874,N_13701,N_14452);
or UO_875 (O_875,N_13105,N_12850);
or UO_876 (O_876,N_14389,N_14394);
nand UO_877 (O_877,N_14137,N_12102);
nand UO_878 (O_878,N_12773,N_13652);
nand UO_879 (O_879,N_12139,N_13403);
nand UO_880 (O_880,N_13138,N_13468);
and UO_881 (O_881,N_13712,N_14297);
nor UO_882 (O_882,N_13699,N_13351);
or UO_883 (O_883,N_13784,N_13859);
and UO_884 (O_884,N_12916,N_14696);
nand UO_885 (O_885,N_14493,N_12365);
and UO_886 (O_886,N_14324,N_12721);
or UO_887 (O_887,N_13015,N_13121);
nand UO_888 (O_888,N_13928,N_12818);
nor UO_889 (O_889,N_12074,N_14907);
nand UO_890 (O_890,N_12695,N_12229);
nor UO_891 (O_891,N_13511,N_13598);
nand UO_892 (O_892,N_12880,N_13079);
or UO_893 (O_893,N_13381,N_12140);
or UO_894 (O_894,N_12086,N_12157);
or UO_895 (O_895,N_12633,N_12526);
or UO_896 (O_896,N_13394,N_12587);
or UO_897 (O_897,N_14267,N_13008);
nor UO_898 (O_898,N_14565,N_12815);
or UO_899 (O_899,N_13452,N_12641);
nand UO_900 (O_900,N_13219,N_13389);
nor UO_901 (O_901,N_13062,N_12297);
nor UO_902 (O_902,N_13570,N_13126);
nor UO_903 (O_903,N_12508,N_14410);
nor UO_904 (O_904,N_13051,N_14162);
or UO_905 (O_905,N_12124,N_14161);
nor UO_906 (O_906,N_12605,N_13466);
nand UO_907 (O_907,N_13196,N_14900);
nor UO_908 (O_908,N_12774,N_12859);
or UO_909 (O_909,N_12154,N_14168);
and UO_910 (O_910,N_14664,N_14901);
and UO_911 (O_911,N_14128,N_14708);
or UO_912 (O_912,N_12429,N_12425);
nor UO_913 (O_913,N_13304,N_14196);
and UO_914 (O_914,N_12757,N_13141);
or UO_915 (O_915,N_14342,N_13515);
nand UO_916 (O_916,N_12482,N_12141);
and UO_917 (O_917,N_12162,N_13853);
and UO_918 (O_918,N_12638,N_14051);
nand UO_919 (O_919,N_13237,N_14989);
nand UO_920 (O_920,N_12117,N_13972);
or UO_921 (O_921,N_12090,N_14828);
nand UO_922 (O_922,N_12377,N_13110);
nand UO_923 (O_923,N_14946,N_12610);
and UO_924 (O_924,N_13285,N_13206);
nand UO_925 (O_925,N_14260,N_13951);
nor UO_926 (O_926,N_13962,N_12105);
and UO_927 (O_927,N_12683,N_12480);
and UO_928 (O_928,N_13457,N_13280);
xnor UO_929 (O_929,N_13535,N_14176);
nor UO_930 (O_930,N_13641,N_12428);
nor UO_931 (O_931,N_14932,N_14760);
and UO_932 (O_932,N_13016,N_13966);
or UO_933 (O_933,N_13412,N_13221);
or UO_934 (O_934,N_14637,N_13626);
nor UO_935 (O_935,N_14714,N_14004);
nand UO_936 (O_936,N_14854,N_13860);
or UO_937 (O_937,N_13176,N_13531);
or UO_938 (O_938,N_13181,N_13571);
nand UO_939 (O_939,N_12976,N_14501);
xnor UO_940 (O_940,N_14851,N_13099);
or UO_941 (O_941,N_12914,N_14803);
or UO_942 (O_942,N_12512,N_14211);
nand UO_943 (O_943,N_13876,N_12125);
nor UO_944 (O_944,N_12120,N_13212);
nor UO_945 (O_945,N_14149,N_14585);
nand UO_946 (O_946,N_14601,N_13434);
and UO_947 (O_947,N_12681,N_12823);
xnor UO_948 (O_948,N_13308,N_12259);
or UO_949 (O_949,N_12285,N_14926);
and UO_950 (O_950,N_13119,N_13582);
or UO_951 (O_951,N_14253,N_12884);
nand UO_952 (O_952,N_12895,N_13604);
or UO_953 (O_953,N_13752,N_13069);
nand UO_954 (O_954,N_14222,N_14536);
and UO_955 (O_955,N_14359,N_13961);
nor UO_956 (O_956,N_14190,N_12144);
nor UO_957 (O_957,N_13131,N_14069);
or UO_958 (O_958,N_13500,N_13494);
nand UO_959 (O_959,N_13488,N_13857);
or UO_960 (O_960,N_12223,N_12922);
nand UO_961 (O_961,N_12553,N_14809);
nor UO_962 (O_962,N_14787,N_12821);
nor UO_963 (O_963,N_12848,N_12847);
nand UO_964 (O_964,N_13382,N_13963);
nand UO_965 (O_965,N_14794,N_12898);
or UO_966 (O_966,N_14591,N_12023);
or UO_967 (O_967,N_12737,N_14597);
nand UO_968 (O_968,N_12291,N_14640);
nand UO_969 (O_969,N_13715,N_12951);
nand UO_970 (O_970,N_12584,N_13986);
nand UO_971 (O_971,N_14915,N_13541);
nor UO_972 (O_972,N_14424,N_13746);
or UO_973 (O_973,N_14074,N_12634);
and UO_974 (O_974,N_12190,N_14117);
or UO_975 (O_975,N_12885,N_13924);
or UO_976 (O_976,N_14463,N_14237);
or UO_977 (O_977,N_13503,N_12137);
and UO_978 (O_978,N_14960,N_14867);
nor UO_979 (O_979,N_13560,N_12458);
or UO_980 (O_980,N_14373,N_14406);
nor UO_981 (O_981,N_13617,N_12801);
nand UO_982 (O_982,N_14949,N_13545);
nand UO_983 (O_983,N_14456,N_13969);
nor UO_984 (O_984,N_13732,N_14088);
nor UO_985 (O_985,N_14917,N_12672);
nand UO_986 (O_986,N_14850,N_13065);
and UO_987 (O_987,N_12111,N_12463);
and UO_988 (O_988,N_13089,N_13091);
and UO_989 (O_989,N_13340,N_13554);
or UO_990 (O_990,N_12308,N_13684);
or UO_991 (O_991,N_12215,N_14171);
nand UO_992 (O_992,N_14083,N_14842);
nand UO_993 (O_993,N_13537,N_13894);
or UO_994 (O_994,N_12674,N_12529);
nor UO_995 (O_995,N_12135,N_12797);
or UO_996 (O_996,N_12016,N_14808);
nor UO_997 (O_997,N_13595,N_13150);
and UO_998 (O_998,N_12468,N_13992);
nor UO_999 (O_999,N_13552,N_13192);
nor UO_1000 (O_1000,N_13465,N_12550);
nand UO_1001 (O_1001,N_12334,N_12065);
nor UO_1002 (O_1002,N_12854,N_12762);
nor UO_1003 (O_1003,N_14538,N_12331);
nand UO_1004 (O_1004,N_14790,N_13549);
nand UO_1005 (O_1005,N_13439,N_14217);
nand UO_1006 (O_1006,N_14332,N_12701);
and UO_1007 (O_1007,N_13562,N_13729);
nand UO_1008 (O_1008,N_13438,N_14212);
nor UO_1009 (O_1009,N_13458,N_13290);
and UO_1010 (O_1010,N_13690,N_13642);
nor UO_1011 (O_1011,N_12092,N_14019);
and UO_1012 (O_1012,N_12307,N_12180);
nand UO_1013 (O_1013,N_13669,N_13325);
nor UO_1014 (O_1014,N_14841,N_12865);
xnor UO_1015 (O_1015,N_14572,N_13092);
xor UO_1016 (O_1016,N_14556,N_13187);
or UO_1017 (O_1017,N_14331,N_14495);
and UO_1018 (O_1018,N_12624,N_12502);
or UO_1019 (O_1019,N_12310,N_14657);
nand UO_1020 (O_1020,N_13367,N_12436);
and UO_1021 (O_1021,N_14918,N_14479);
or UO_1022 (O_1022,N_13191,N_13301);
nand UO_1023 (O_1023,N_12886,N_12752);
and UO_1024 (O_1024,N_13456,N_12814);
and UO_1025 (O_1025,N_13926,N_13809);
or UO_1026 (O_1026,N_12187,N_13056);
or UO_1027 (O_1027,N_12407,N_13305);
or UO_1028 (O_1028,N_13959,N_12769);
and UO_1029 (O_1029,N_12048,N_14618);
or UO_1030 (O_1030,N_12033,N_12330);
nand UO_1031 (O_1031,N_13527,N_12889);
or UO_1032 (O_1032,N_14306,N_14338);
nor UO_1033 (O_1033,N_12390,N_14689);
and UO_1034 (O_1034,N_14680,N_12106);
nor UO_1035 (O_1035,N_14058,N_12034);
nand UO_1036 (O_1036,N_12430,N_12399);
nor UO_1037 (O_1037,N_13782,N_13685);
nand UO_1038 (O_1038,N_13749,N_13096);
and UO_1039 (O_1039,N_12305,N_12763);
nor UO_1040 (O_1040,N_13490,N_14957);
nor UO_1041 (O_1041,N_14895,N_14431);
nor UO_1042 (O_1042,N_12939,N_14037);
or UO_1043 (O_1043,N_13887,N_13112);
and UO_1044 (O_1044,N_12965,N_12510);
or UO_1045 (O_1045,N_14958,N_13149);
nand UO_1046 (O_1046,N_12968,N_13326);
and UO_1047 (O_1047,N_14308,N_13111);
nand UO_1048 (O_1048,N_13036,N_13716);
xnor UO_1049 (O_1049,N_13122,N_14249);
or UO_1050 (O_1050,N_13829,N_14450);
xnor UO_1051 (O_1051,N_12750,N_14361);
or UO_1052 (O_1052,N_13683,N_13574);
or UO_1053 (O_1053,N_14138,N_13773);
nand UO_1054 (O_1054,N_12775,N_13647);
nand UO_1055 (O_1055,N_14221,N_13061);
and UO_1056 (O_1056,N_14563,N_12532);
and UO_1057 (O_1057,N_14014,N_13414);
nand UO_1058 (O_1058,N_12014,N_14768);
and UO_1059 (O_1059,N_14121,N_14207);
or UO_1060 (O_1060,N_14409,N_14552);
or UO_1061 (O_1061,N_12741,N_14320);
or UO_1062 (O_1062,N_14924,N_13678);
nor UO_1063 (O_1063,N_12266,N_13379);
or UO_1064 (O_1064,N_12057,N_13640);
nor UO_1065 (O_1065,N_14846,N_12840);
xor UO_1066 (O_1066,N_13899,N_13356);
or UO_1067 (O_1067,N_14522,N_14155);
and UO_1068 (O_1068,N_14624,N_12049);
or UO_1069 (O_1069,N_12444,N_12743);
and UO_1070 (O_1070,N_12956,N_14868);
nand UO_1071 (O_1071,N_14457,N_12620);
nand UO_1072 (O_1072,N_13258,N_14244);
or UO_1073 (O_1073,N_14427,N_13547);
and UO_1074 (O_1074,N_14208,N_14499);
or UO_1075 (O_1075,N_14327,N_13031);
nand UO_1076 (O_1076,N_13128,N_14438);
and UO_1077 (O_1077,N_14972,N_14065);
and UO_1078 (O_1078,N_13973,N_14250);
or UO_1079 (O_1079,N_14629,N_12700);
nor UO_1080 (O_1080,N_13251,N_13302);
and UO_1081 (O_1081,N_13852,N_12833);
or UO_1082 (O_1082,N_13273,N_14551);
and UO_1083 (O_1083,N_14387,N_12008);
and UO_1084 (O_1084,N_12644,N_12177);
xor UO_1085 (O_1085,N_12216,N_12679);
nor UO_1086 (O_1086,N_13812,N_12900);
nor UO_1087 (O_1087,N_12988,N_14227);
or UO_1088 (O_1088,N_13035,N_13657);
and UO_1089 (O_1089,N_14873,N_13919);
or UO_1090 (O_1090,N_13256,N_13738);
and UO_1091 (O_1091,N_12160,N_13776);
and UO_1092 (O_1092,N_12756,N_14334);
nor UO_1093 (O_1093,N_12520,N_13253);
nand UO_1094 (O_1094,N_14192,N_12606);
nor UO_1095 (O_1095,N_12973,N_12582);
nand UO_1096 (O_1096,N_12374,N_13753);
and UO_1097 (O_1097,N_13436,N_12770);
or UO_1098 (O_1098,N_12534,N_14469);
nand UO_1099 (O_1099,N_12378,N_12218);
nor UO_1100 (O_1100,N_13482,N_13082);
nand UO_1101 (O_1101,N_13354,N_13155);
nor UO_1102 (O_1102,N_12653,N_14934);
nor UO_1103 (O_1103,N_14437,N_12001);
and UO_1104 (O_1104,N_12498,N_14018);
or UO_1105 (O_1105,N_13682,N_12708);
and UO_1106 (O_1106,N_14323,N_13193);
or UO_1107 (O_1107,N_13106,N_14378);
nor UO_1108 (O_1108,N_13357,N_13114);
and UO_1109 (O_1109,N_14370,N_14064);
nor UO_1110 (O_1110,N_14465,N_13199);
or UO_1111 (O_1111,N_14844,N_14883);
nor UO_1112 (O_1112,N_14172,N_14524);
nand UO_1113 (O_1113,N_13088,N_14855);
nor UO_1114 (O_1114,N_12519,N_12395);
nand UO_1115 (O_1115,N_12538,N_14328);
and UO_1116 (O_1116,N_13880,N_13224);
or UO_1117 (O_1117,N_13104,N_14118);
nand UO_1118 (O_1118,N_14811,N_12181);
nor UO_1119 (O_1119,N_12293,N_14662);
nand UO_1120 (O_1120,N_14107,N_14030);
and UO_1121 (O_1121,N_12554,N_13526);
and UO_1122 (O_1122,N_12341,N_14721);
and UO_1123 (O_1123,N_13686,N_14319);
nand UO_1124 (O_1124,N_14081,N_13269);
nor UO_1125 (O_1125,N_13522,N_13806);
or UO_1126 (O_1126,N_12040,N_14349);
or UO_1127 (O_1127,N_12313,N_14669);
nand UO_1128 (O_1128,N_12352,N_14598);
or UO_1129 (O_1129,N_14693,N_12245);
nor UO_1130 (O_1130,N_13312,N_13858);
and UO_1131 (O_1131,N_12275,N_13182);
nand UO_1132 (O_1132,N_13741,N_14318);
and UO_1133 (O_1133,N_14169,N_13323);
nand UO_1134 (O_1134,N_12222,N_12796);
or UO_1135 (O_1135,N_12648,N_12198);
or UO_1136 (O_1136,N_12312,N_13374);
nand UO_1137 (O_1137,N_12299,N_13918);
nor UO_1138 (O_1138,N_13977,N_12919);
nor UO_1139 (O_1139,N_12237,N_14723);
nand UO_1140 (O_1140,N_13704,N_12524);
nand UO_1141 (O_1141,N_14955,N_12478);
nand UO_1142 (O_1142,N_12997,N_14665);
or UO_1143 (O_1143,N_14786,N_14782);
nand UO_1144 (O_1144,N_14730,N_12839);
and UO_1145 (O_1145,N_13041,N_13538);
nand UO_1146 (O_1146,N_13734,N_12271);
nand UO_1147 (O_1147,N_14020,N_14265);
nor UO_1148 (O_1148,N_13146,N_14290);
or UO_1149 (O_1149,N_13980,N_13052);
nor UO_1150 (O_1150,N_13799,N_13721);
or UO_1151 (O_1151,N_12011,N_14927);
nand UO_1152 (O_1152,N_13865,N_12966);
or UO_1153 (O_1153,N_12734,N_13745);
nand UO_1154 (O_1154,N_12949,N_13744);
and UO_1155 (O_1155,N_12238,N_14603);
nor UO_1156 (O_1156,N_14356,N_14011);
nor UO_1157 (O_1157,N_14778,N_14732);
and UO_1158 (O_1158,N_12811,N_12541);
nor UO_1159 (O_1159,N_14305,N_12133);
nor UO_1160 (O_1160,N_14568,N_12211);
nand UO_1161 (O_1161,N_13081,N_13733);
nand UO_1162 (O_1162,N_13660,N_12635);
nand UO_1163 (O_1163,N_13610,N_13252);
nor UO_1164 (O_1164,N_13272,N_14587);
or UO_1165 (O_1165,N_12485,N_13045);
nand UO_1166 (O_1166,N_14903,N_14369);
nor UO_1167 (O_1167,N_14675,N_12946);
and UO_1168 (O_1168,N_12907,N_12193);
nor UO_1169 (O_1169,N_13555,N_14185);
nor UO_1170 (O_1170,N_13611,N_13278);
or UO_1171 (O_1171,N_14132,N_12849);
nand UO_1172 (O_1172,N_14263,N_14644);
or UO_1173 (O_1173,N_12446,N_12301);
nand UO_1174 (O_1174,N_12321,N_12409);
nand UO_1175 (O_1175,N_12206,N_12093);
nor UO_1176 (O_1176,N_12289,N_12999);
nand UO_1177 (O_1177,N_12611,N_12754);
and UO_1178 (O_1178,N_13152,N_14617);
and UO_1179 (O_1179,N_12632,N_12451);
nor UO_1180 (O_1180,N_12340,N_12926);
and UO_1181 (O_1181,N_14180,N_14255);
or UO_1182 (O_1182,N_13759,N_13165);
or UO_1183 (O_1183,N_13661,N_14421);
nor UO_1184 (O_1184,N_13975,N_14812);
and UO_1185 (O_1185,N_14633,N_14301);
and UO_1186 (O_1186,N_14339,N_14213);
and UO_1187 (O_1187,N_13597,N_14256);
or UO_1188 (O_1188,N_13725,N_12804);
nor UO_1189 (O_1189,N_14518,N_13593);
nand UO_1190 (O_1190,N_13765,N_13474);
nand UO_1191 (O_1191,N_12712,N_13449);
nor UO_1192 (O_1192,N_14911,N_13825);
or UO_1193 (O_1193,N_14733,N_14453);
and UO_1194 (O_1194,N_14054,N_14100);
and UO_1195 (O_1195,N_12822,N_13442);
nor UO_1196 (O_1196,N_13136,N_13867);
or UO_1197 (O_1197,N_14418,N_13989);
nor UO_1198 (O_1198,N_12286,N_14345);
and UO_1199 (O_1199,N_13532,N_13336);
nand UO_1200 (O_1200,N_13025,N_13397);
and UO_1201 (O_1201,N_13415,N_14225);
or UO_1202 (O_1202,N_13650,N_12304);
or UO_1203 (O_1203,N_13270,N_12486);
nand UO_1204 (O_1204,N_14831,N_14119);
and UO_1205 (O_1205,N_14150,N_13362);
nor UO_1206 (O_1206,N_12581,N_12984);
nor UO_1207 (O_1207,N_13510,N_13847);
nand UO_1208 (O_1208,N_14296,N_12528);
nand UO_1209 (O_1209,N_14206,N_14474);
and UO_1210 (O_1210,N_13274,N_12810);
nor UO_1211 (O_1211,N_13319,N_12185);
xnor UO_1212 (O_1212,N_12652,N_14859);
nor UO_1213 (O_1213,N_12476,N_14769);
nand UO_1214 (O_1214,N_13287,N_14621);
and UO_1215 (O_1215,N_12163,N_13583);
nand UO_1216 (O_1216,N_13097,N_12619);
or UO_1217 (O_1217,N_14759,N_14885);
nand UO_1218 (O_1218,N_12221,N_14709);
nor UO_1219 (O_1219,N_13727,N_12852);
or UO_1220 (O_1220,N_13946,N_14408);
or UO_1221 (O_1221,N_14104,N_14939);
nand UO_1222 (O_1222,N_12566,N_13873);
nor UO_1223 (O_1223,N_13872,N_14177);
and UO_1224 (O_1224,N_13688,N_13864);
and UO_1225 (O_1225,N_12182,N_14357);
and UO_1226 (O_1226,N_12863,N_13201);
nand UO_1227 (O_1227,N_14893,N_13044);
and UO_1228 (O_1228,N_12666,N_12842);
or UO_1229 (O_1229,N_12578,N_14674);
and UO_1230 (O_1230,N_13402,N_12131);
and UO_1231 (O_1231,N_13728,N_14595);
nand UO_1232 (O_1232,N_13982,N_14072);
and UO_1233 (O_1233,N_12593,N_14084);
or UO_1234 (O_1234,N_14352,N_12462);
and UO_1235 (O_1235,N_12196,N_14397);
nor UO_1236 (O_1236,N_14282,N_12064);
nor UO_1237 (O_1237,N_12901,N_13148);
nor UO_1238 (O_1238,N_13629,N_12970);
or UO_1239 (O_1239,N_12239,N_14744);
nand UO_1240 (O_1240,N_12108,N_13839);
or UO_1241 (O_1241,N_12950,N_12265);
nor UO_1242 (O_1242,N_12870,N_14642);
nand UO_1243 (O_1243,N_14044,N_14921);
nand UO_1244 (O_1244,N_12748,N_14829);
and UO_1245 (O_1245,N_12594,N_13223);
and UO_1246 (O_1246,N_13556,N_13875);
nor UO_1247 (O_1247,N_14125,N_12911);
nand UO_1248 (O_1248,N_13823,N_14987);
or UO_1249 (O_1249,N_13590,N_12618);
or UO_1250 (O_1250,N_12851,N_12258);
nor UO_1251 (O_1251,N_13417,N_12358);
and UO_1252 (O_1252,N_13125,N_12768);
or UO_1253 (O_1253,N_12143,N_12829);
or UO_1254 (O_1254,N_12920,N_13186);
or UO_1255 (O_1255,N_14231,N_14834);
nand UO_1256 (O_1256,N_13130,N_13711);
nor UO_1257 (O_1257,N_13293,N_14280);
xor UO_1258 (O_1258,N_14992,N_12220);
and UO_1259 (O_1259,N_13021,N_13994);
or UO_1260 (O_1260,N_13987,N_14013);
nor UO_1261 (O_1261,N_14428,N_14315);
or UO_1262 (O_1262,N_12061,N_13006);
nand UO_1263 (O_1263,N_14472,N_13658);
nor UO_1264 (O_1264,N_14355,N_13637);
nor UO_1265 (O_1265,N_13143,N_12030);
and UO_1266 (O_1266,N_12384,N_13636);
nand UO_1267 (O_1267,N_12733,N_13623);
nor UO_1268 (O_1268,N_12913,N_12123);
nand UO_1269 (O_1269,N_14028,N_13737);
nand UO_1270 (O_1270,N_13460,N_13469);
nor UO_1271 (O_1271,N_14775,N_12685);
or UO_1272 (O_1272,N_12225,N_12930);
and UO_1273 (O_1273,N_14050,N_12172);
nand UO_1274 (O_1274,N_14063,N_13523);
or UO_1275 (O_1275,N_14990,N_12902);
and UO_1276 (O_1276,N_13024,N_13238);
nor UO_1277 (O_1277,N_13757,N_14880);
and UO_1278 (O_1278,N_12651,N_12450);
or UO_1279 (O_1279,N_12195,N_12396);
and UO_1280 (O_1280,N_12469,N_14492);
and UO_1281 (O_1281,N_14271,N_14239);
nor UO_1282 (O_1282,N_13546,N_13213);
or UO_1283 (O_1283,N_12052,N_13259);
nor UO_1284 (O_1284,N_14198,N_13352);
and UO_1285 (O_1285,N_13838,N_13250);
nor UO_1286 (O_1286,N_13792,N_13388);
nor UO_1287 (O_1287,N_12306,N_14123);
and UO_1288 (O_1288,N_12881,N_14720);
nor UO_1289 (O_1289,N_13137,N_13393);
or UO_1290 (O_1290,N_13108,N_12746);
or UO_1291 (O_1291,N_14750,N_14511);
and UO_1292 (O_1292,N_14099,N_13430);
and UO_1293 (O_1293,N_12070,N_14748);
nand UO_1294 (O_1294,N_14012,N_13676);
and UO_1295 (O_1295,N_13307,N_12232);
or UO_1296 (O_1296,N_12720,N_12678);
or UO_1297 (O_1297,N_13892,N_12324);
or UO_1298 (O_1298,N_12171,N_14931);
and UO_1299 (O_1299,N_14344,N_14673);
nor UO_1300 (O_1300,N_12548,N_14494);
and UO_1301 (O_1301,N_14136,N_12932);
and UO_1302 (O_1302,N_12609,N_12311);
and UO_1303 (O_1303,N_14087,N_12597);
or UO_1304 (O_1304,N_14194,N_14910);
nand UO_1305 (O_1305,N_13520,N_13763);
or UO_1306 (O_1306,N_12414,N_12826);
and UO_1307 (O_1307,N_13514,N_13050);
and UO_1308 (O_1308,N_13169,N_12422);
or UO_1309 (O_1309,N_13644,N_14592);
nand UO_1310 (O_1310,N_14274,N_13317);
or UO_1311 (O_1311,N_14302,N_13995);
or UO_1312 (O_1312,N_12791,N_12083);
or UO_1313 (O_1313,N_14476,N_12742);
nor UO_1314 (O_1314,N_12718,N_14354);
nand UO_1315 (O_1315,N_14160,N_14078);
or UO_1316 (O_1316,N_14252,N_12658);
or UO_1317 (O_1317,N_14848,N_14660);
or UO_1318 (O_1318,N_14275,N_13943);
and UO_1319 (O_1319,N_13648,N_14210);
nor UO_1320 (O_1320,N_14309,N_12370);
and UO_1321 (O_1321,N_14988,N_13895);
xor UO_1322 (O_1322,N_12152,N_12495);
and UO_1323 (O_1323,N_14874,N_12025);
nor UO_1324 (O_1324,N_14503,N_14532);
nand UO_1325 (O_1325,N_14919,N_12003);
nor UO_1326 (O_1326,N_12095,N_14826);
or UO_1327 (O_1327,N_12986,N_14928);
or UO_1328 (O_1328,N_14785,N_12527);
and UO_1329 (O_1329,N_13211,N_13559);
nor UO_1330 (O_1330,N_14098,N_13539);
nor UO_1331 (O_1331,N_13018,N_13189);
nor UO_1332 (O_1332,N_12556,N_14801);
nor UO_1333 (O_1333,N_13889,N_12549);
nor UO_1334 (O_1334,N_14443,N_13359);
nor UO_1335 (O_1335,N_12336,N_13360);
or UO_1336 (O_1336,N_14571,N_14001);
nor UO_1337 (O_1337,N_12602,N_12419);
nand UO_1338 (O_1338,N_13691,N_13822);
nor UO_1339 (O_1339,N_14719,N_12183);
nand UO_1340 (O_1340,N_14942,N_14245);
nand UO_1341 (O_1341,N_12588,N_14817);
and UO_1342 (O_1342,N_13673,N_12586);
nand UO_1343 (O_1343,N_13380,N_12488);
and UO_1344 (O_1344,N_14833,N_14836);
and UO_1345 (O_1345,N_14906,N_13431);
xnor UO_1346 (O_1346,N_12686,N_13372);
or UO_1347 (O_1347,N_13569,N_14923);
and UO_1348 (O_1348,N_13002,N_14496);
and UO_1349 (O_1349,N_12668,N_12412);
and UO_1350 (O_1350,N_13139,N_12359);
and UO_1351 (O_1351,N_14777,N_13529);
or UO_1352 (O_1352,N_14420,N_14681);
nand UO_1353 (O_1353,N_13234,N_13020);
or UO_1354 (O_1354,N_13396,N_14126);
nand UO_1355 (O_1355,N_13405,N_13920);
xor UO_1356 (O_1356,N_14392,N_14530);
or UO_1357 (O_1357,N_12438,N_14299);
nand UO_1358 (O_1358,N_14382,N_13672);
nor UO_1359 (O_1359,N_14922,N_13228);
nand UO_1360 (O_1360,N_12046,N_12026);
and UO_1361 (O_1361,N_14796,N_14753);
or UO_1362 (O_1362,N_14145,N_12091);
and UO_1363 (O_1363,N_14508,N_14626);
and UO_1364 (O_1364,N_12010,N_14685);
or UO_1365 (O_1365,N_14071,N_12989);
or UO_1366 (O_1366,N_13722,N_14451);
nor UO_1367 (O_1367,N_12827,N_12325);
nor UO_1368 (O_1368,N_12159,N_12749);
nand UO_1369 (O_1369,N_13952,N_12551);
nor UO_1370 (O_1370,N_13344,N_12858);
or UO_1371 (O_1371,N_12662,N_14546);
or UO_1372 (O_1372,N_14056,N_13758);
or UO_1373 (O_1373,N_12368,N_13073);
nor UO_1374 (O_1374,N_14313,N_13226);
nor UO_1375 (O_1375,N_13231,N_13408);
or UO_1376 (O_1376,N_12918,N_13124);
or UO_1377 (O_1377,N_14061,N_14741);
or UO_1378 (O_1378,N_13032,N_12322);
xor UO_1379 (O_1379,N_12963,N_13634);
and UO_1380 (O_1380,N_14101,N_13409);
or UO_1381 (O_1381,N_12103,N_14283);
nor UO_1382 (O_1382,N_13709,N_13923);
or UO_1383 (O_1383,N_13267,N_13580);
and UO_1384 (O_1384,N_14943,N_12836);
and UO_1385 (O_1385,N_12393,N_14818);
or UO_1386 (O_1386,N_12323,N_12267);
nand UO_1387 (O_1387,N_14367,N_12617);
or UO_1388 (O_1388,N_12625,N_13028);
nor UO_1389 (O_1389,N_13416,N_13790);
nand UO_1390 (O_1390,N_12199,N_13010);
and UO_1391 (O_1391,N_14638,N_13314);
nor UO_1392 (O_1392,N_13084,N_14086);
nor UO_1393 (O_1393,N_12802,N_13948);
and UO_1394 (O_1394,N_14070,N_14109);
or UO_1395 (O_1395,N_12846,N_12657);
nor UO_1396 (O_1396,N_12855,N_12319);
or UO_1397 (O_1397,N_12058,N_13921);
or UO_1398 (O_1398,N_14017,N_12798);
nand UO_1399 (O_1399,N_14558,N_12112);
nand UO_1400 (O_1400,N_12991,N_12961);
nor UO_1401 (O_1401,N_13877,N_13993);
and UO_1402 (O_1402,N_14607,N_12208);
nor UO_1403 (O_1403,N_14994,N_12278);
and UO_1404 (O_1404,N_13841,N_12730);
nor UO_1405 (O_1405,N_12523,N_13355);
nand UO_1406 (O_1406,N_14613,N_12204);
or UO_1407 (O_1407,N_13724,N_14970);
and UO_1408 (O_1408,N_13679,N_14950);
nor UO_1409 (O_1409,N_13247,N_12807);
nand UO_1410 (O_1410,N_14755,N_12300);
nand UO_1411 (O_1411,N_14166,N_13762);
and UO_1412 (O_1412,N_14979,N_13068);
or UO_1413 (O_1413,N_14967,N_14737);
and UO_1414 (O_1414,N_12879,N_12471);
and UO_1415 (O_1415,N_14751,N_13004);
or UO_1416 (O_1416,N_14130,N_13135);
nor UO_1417 (O_1417,N_14682,N_14604);
nor UO_1418 (O_1418,N_12740,N_14234);
nor UO_1419 (O_1419,N_12345,N_13132);
nor UO_1420 (O_1420,N_12861,N_14754);
nor UO_1421 (O_1421,N_12924,N_13327);
nand UO_1422 (O_1422,N_14559,N_14860);
nand UO_1423 (O_1423,N_12953,N_12338);
or UO_1424 (O_1424,N_14152,N_12530);
and UO_1425 (O_1425,N_13263,N_13747);
nand UO_1426 (O_1426,N_12353,N_13708);
nand UO_1427 (O_1427,N_14814,N_14909);
nand UO_1428 (O_1428,N_13668,N_12075);
nand UO_1429 (O_1429,N_14526,N_13934);
nand UO_1430 (O_1430,N_13801,N_12248);
or UO_1431 (O_1431,N_12231,N_13334);
or UO_1432 (O_1432,N_13098,N_13940);
nor UO_1433 (O_1433,N_13321,N_13311);
and UO_1434 (O_1434,N_12789,N_13245);
and UO_1435 (O_1435,N_14577,N_12535);
and UO_1436 (O_1436,N_13320,N_14073);
nor UO_1437 (O_1437,N_13227,N_12921);
nor UO_1438 (O_1438,N_14724,N_14229);
nor UO_1439 (O_1439,N_13941,N_14699);
and UO_1440 (O_1440,N_13813,N_14863);
and UO_1441 (O_1441,N_12764,N_14405);
and UO_1442 (O_1442,N_12041,N_12837);
and UO_1443 (O_1443,N_14407,N_12612);
and UO_1444 (O_1444,N_14773,N_13070);
and UO_1445 (O_1445,N_14288,N_14413);
nor UO_1446 (O_1446,N_14203,N_14852);
nand UO_1447 (O_1447,N_13906,N_14279);
or UO_1448 (O_1448,N_14630,N_13840);
nor UO_1449 (O_1449,N_13455,N_13976);
nor UO_1450 (O_1450,N_12383,N_12724);
nor UO_1451 (O_1451,N_13783,N_12501);
or UO_1452 (O_1452,N_13030,N_13260);
nand UO_1453 (O_1453,N_12630,N_13316);
or UO_1454 (O_1454,N_12975,N_12576);
nand UO_1455 (O_1455,N_13905,N_12233);
or UO_1456 (O_1456,N_13754,N_13172);
nor UO_1457 (O_1457,N_14764,N_13620);
nor UO_1458 (O_1458,N_12972,N_12936);
and UO_1459 (O_1459,N_14529,N_14110);
nand UO_1460 (O_1460,N_13900,N_14700);
or UO_1461 (O_1461,N_14632,N_13496);
nor UO_1462 (O_1462,N_12817,N_14703);
nand UO_1463 (O_1463,N_12031,N_14537);
nor UO_1464 (O_1464,N_14763,N_14752);
and UO_1465 (O_1465,N_13846,N_14266);
nand UO_1466 (O_1466,N_14146,N_14590);
or UO_1467 (O_1467,N_14899,N_12035);
or UO_1468 (O_1468,N_14461,N_12318);
nor UO_1469 (O_1469,N_14447,N_12020);
xor UO_1470 (O_1470,N_14233,N_14159);
or UO_1471 (O_1471,N_13328,N_13798);
nand UO_1472 (O_1472,N_14448,N_12270);
nor UO_1473 (O_1473,N_12561,N_14032);
or UO_1474 (O_1474,N_13283,N_13638);
nand UO_1475 (O_1475,N_12853,N_12636);
nor UO_1476 (O_1476,N_14031,N_14403);
or UO_1477 (O_1477,N_14717,N_12883);
nand UO_1478 (O_1478,N_12689,N_12698);
nand UO_1479 (O_1479,N_13168,N_13459);
nand UO_1480 (O_1480,N_12621,N_12964);
and UO_1481 (O_1481,N_14025,N_12122);
and UO_1482 (O_1482,N_13129,N_14619);
nand UO_1483 (O_1483,N_12568,N_12813);
and UO_1484 (O_1484,N_12776,N_14898);
nand UO_1485 (O_1485,N_14599,N_14788);
nor UO_1486 (O_1486,N_14151,N_13849);
nand UO_1487 (O_1487,N_13718,N_13406);
or UO_1488 (O_1488,N_14727,N_13433);
nor UO_1489 (O_1489,N_14625,N_14845);
nand UO_1490 (O_1490,N_13342,N_13573);
nor UO_1491 (O_1491,N_13828,N_12128);
and UO_1492 (O_1492,N_13345,N_13796);
nand UO_1493 (O_1493,N_13705,N_14815);
nor UO_1494 (O_1494,N_13544,N_13735);
or UO_1495 (O_1495,N_13967,N_12892);
xor UO_1496 (O_1496,N_14807,N_14295);
nor UO_1497 (O_1497,N_14584,N_14115);
nand UO_1498 (O_1498,N_12585,N_14981);
nand UO_1499 (O_1499,N_12372,N_14959);
nand UO_1500 (O_1500,N_13044,N_13872);
or UO_1501 (O_1501,N_12077,N_14093);
xor UO_1502 (O_1502,N_14713,N_12142);
nor UO_1503 (O_1503,N_14002,N_14052);
or UO_1504 (O_1504,N_12884,N_12011);
or UO_1505 (O_1505,N_12154,N_12333);
and UO_1506 (O_1506,N_14234,N_13148);
and UO_1507 (O_1507,N_12035,N_12133);
nor UO_1508 (O_1508,N_13677,N_12484);
nand UO_1509 (O_1509,N_13467,N_12286);
nand UO_1510 (O_1510,N_12352,N_14592);
nor UO_1511 (O_1511,N_13377,N_14011);
and UO_1512 (O_1512,N_14720,N_13322);
or UO_1513 (O_1513,N_13859,N_12152);
nor UO_1514 (O_1514,N_12004,N_14499);
or UO_1515 (O_1515,N_13040,N_14568);
and UO_1516 (O_1516,N_13729,N_12856);
nor UO_1517 (O_1517,N_12138,N_14822);
nand UO_1518 (O_1518,N_13442,N_12566);
and UO_1519 (O_1519,N_14462,N_14755);
and UO_1520 (O_1520,N_13414,N_14083);
or UO_1521 (O_1521,N_13584,N_14004);
and UO_1522 (O_1522,N_12997,N_13370);
or UO_1523 (O_1523,N_14912,N_13554);
xnor UO_1524 (O_1524,N_14241,N_12732);
nand UO_1525 (O_1525,N_14670,N_13639);
nand UO_1526 (O_1526,N_13812,N_13171);
nor UO_1527 (O_1527,N_13093,N_14215);
or UO_1528 (O_1528,N_13562,N_12266);
or UO_1529 (O_1529,N_12799,N_13691);
or UO_1530 (O_1530,N_13353,N_13966);
and UO_1531 (O_1531,N_12498,N_14601);
nand UO_1532 (O_1532,N_13168,N_14784);
and UO_1533 (O_1533,N_13778,N_12655);
nor UO_1534 (O_1534,N_12964,N_14074);
and UO_1535 (O_1535,N_13678,N_12236);
and UO_1536 (O_1536,N_13719,N_14405);
and UO_1537 (O_1537,N_13998,N_12005);
and UO_1538 (O_1538,N_14382,N_13729);
and UO_1539 (O_1539,N_12891,N_14890);
nand UO_1540 (O_1540,N_14303,N_14009);
and UO_1541 (O_1541,N_12513,N_13079);
and UO_1542 (O_1542,N_14308,N_13879);
xnor UO_1543 (O_1543,N_12058,N_14388);
or UO_1544 (O_1544,N_12061,N_12906);
nor UO_1545 (O_1545,N_12129,N_13041);
and UO_1546 (O_1546,N_12523,N_13959);
and UO_1547 (O_1547,N_13528,N_13781);
nand UO_1548 (O_1548,N_12540,N_14822);
nand UO_1549 (O_1549,N_14511,N_12474);
nand UO_1550 (O_1550,N_13946,N_12871);
nand UO_1551 (O_1551,N_14846,N_13693);
nor UO_1552 (O_1552,N_13976,N_14375);
nor UO_1553 (O_1553,N_13203,N_14855);
nor UO_1554 (O_1554,N_13438,N_13872);
nand UO_1555 (O_1555,N_14030,N_12890);
nor UO_1556 (O_1556,N_13697,N_14551);
nor UO_1557 (O_1557,N_14373,N_14316);
nor UO_1558 (O_1558,N_12550,N_12444);
nand UO_1559 (O_1559,N_14481,N_14424);
nand UO_1560 (O_1560,N_14816,N_13143);
nor UO_1561 (O_1561,N_13086,N_14601);
and UO_1562 (O_1562,N_12027,N_13112);
and UO_1563 (O_1563,N_14606,N_14771);
or UO_1564 (O_1564,N_13628,N_13949);
nor UO_1565 (O_1565,N_12462,N_12651);
nor UO_1566 (O_1566,N_12166,N_13690);
and UO_1567 (O_1567,N_13911,N_14777);
nor UO_1568 (O_1568,N_12433,N_13993);
nor UO_1569 (O_1569,N_14673,N_13234);
and UO_1570 (O_1570,N_13499,N_14715);
and UO_1571 (O_1571,N_12957,N_12509);
or UO_1572 (O_1572,N_13647,N_12698);
or UO_1573 (O_1573,N_14533,N_12044);
nand UO_1574 (O_1574,N_12415,N_14269);
nor UO_1575 (O_1575,N_12123,N_12653);
or UO_1576 (O_1576,N_14998,N_13790);
or UO_1577 (O_1577,N_12132,N_13607);
nor UO_1578 (O_1578,N_13484,N_14849);
or UO_1579 (O_1579,N_12735,N_13077);
nand UO_1580 (O_1580,N_12487,N_12796);
and UO_1581 (O_1581,N_12374,N_14105);
nand UO_1582 (O_1582,N_12439,N_13215);
nor UO_1583 (O_1583,N_13215,N_14683);
nor UO_1584 (O_1584,N_13960,N_13789);
nand UO_1585 (O_1585,N_14005,N_12325);
or UO_1586 (O_1586,N_13940,N_12740);
nand UO_1587 (O_1587,N_12348,N_12696);
or UO_1588 (O_1588,N_14192,N_14053);
or UO_1589 (O_1589,N_13679,N_13121);
nor UO_1590 (O_1590,N_14823,N_13463);
and UO_1591 (O_1591,N_14931,N_13299);
or UO_1592 (O_1592,N_13778,N_14319);
nand UO_1593 (O_1593,N_12209,N_13809);
or UO_1594 (O_1594,N_14701,N_12300);
nor UO_1595 (O_1595,N_14725,N_12226);
nor UO_1596 (O_1596,N_13764,N_12902);
nor UO_1597 (O_1597,N_14522,N_12013);
nand UO_1598 (O_1598,N_12689,N_14278);
nor UO_1599 (O_1599,N_14922,N_12214);
nand UO_1600 (O_1600,N_12365,N_13042);
or UO_1601 (O_1601,N_13848,N_14867);
nand UO_1602 (O_1602,N_14221,N_14310);
nor UO_1603 (O_1603,N_13192,N_12607);
and UO_1604 (O_1604,N_14783,N_12263);
nor UO_1605 (O_1605,N_12688,N_13242);
xor UO_1606 (O_1606,N_14382,N_12630);
and UO_1607 (O_1607,N_12587,N_12032);
nand UO_1608 (O_1608,N_13362,N_14082);
nand UO_1609 (O_1609,N_14122,N_12687);
nor UO_1610 (O_1610,N_12017,N_13087);
nand UO_1611 (O_1611,N_14924,N_12281);
and UO_1612 (O_1612,N_14464,N_12532);
nand UO_1613 (O_1613,N_12420,N_13326);
nor UO_1614 (O_1614,N_13270,N_13298);
or UO_1615 (O_1615,N_13811,N_13665);
nor UO_1616 (O_1616,N_13741,N_13904);
nand UO_1617 (O_1617,N_12797,N_14526);
nor UO_1618 (O_1618,N_13139,N_13926);
nand UO_1619 (O_1619,N_14326,N_14594);
nor UO_1620 (O_1620,N_14319,N_13381);
and UO_1621 (O_1621,N_12593,N_13365);
or UO_1622 (O_1622,N_12625,N_12920);
or UO_1623 (O_1623,N_14431,N_14199);
and UO_1624 (O_1624,N_14114,N_12665);
and UO_1625 (O_1625,N_13405,N_12869);
or UO_1626 (O_1626,N_13457,N_13503);
and UO_1627 (O_1627,N_14163,N_13936);
or UO_1628 (O_1628,N_12315,N_14491);
or UO_1629 (O_1629,N_13813,N_12055);
nand UO_1630 (O_1630,N_13183,N_14808);
or UO_1631 (O_1631,N_12721,N_14847);
xnor UO_1632 (O_1632,N_14563,N_12858);
xnor UO_1633 (O_1633,N_13398,N_14044);
nand UO_1634 (O_1634,N_12908,N_14138);
or UO_1635 (O_1635,N_13047,N_14319);
or UO_1636 (O_1636,N_14119,N_13660);
or UO_1637 (O_1637,N_12880,N_13874);
xor UO_1638 (O_1638,N_13150,N_12012);
or UO_1639 (O_1639,N_13632,N_12757);
or UO_1640 (O_1640,N_13033,N_13265);
or UO_1641 (O_1641,N_14251,N_13801);
and UO_1642 (O_1642,N_12241,N_12148);
nand UO_1643 (O_1643,N_12465,N_12979);
nand UO_1644 (O_1644,N_14236,N_13179);
or UO_1645 (O_1645,N_14783,N_12826);
nand UO_1646 (O_1646,N_14344,N_12974);
nor UO_1647 (O_1647,N_12414,N_13940);
nand UO_1648 (O_1648,N_12783,N_12446);
nor UO_1649 (O_1649,N_12212,N_13530);
nor UO_1650 (O_1650,N_13241,N_12006);
and UO_1651 (O_1651,N_12053,N_13520);
or UO_1652 (O_1652,N_13411,N_14458);
or UO_1653 (O_1653,N_13294,N_13905);
nand UO_1654 (O_1654,N_13080,N_14568);
nor UO_1655 (O_1655,N_13787,N_13655);
nor UO_1656 (O_1656,N_14858,N_13141);
or UO_1657 (O_1657,N_12243,N_12005);
or UO_1658 (O_1658,N_13416,N_12902);
and UO_1659 (O_1659,N_14755,N_13384);
or UO_1660 (O_1660,N_12182,N_13442);
and UO_1661 (O_1661,N_13586,N_13336);
or UO_1662 (O_1662,N_14593,N_12511);
or UO_1663 (O_1663,N_12346,N_14870);
or UO_1664 (O_1664,N_14226,N_12901);
nor UO_1665 (O_1665,N_13261,N_13686);
or UO_1666 (O_1666,N_13681,N_13367);
nor UO_1667 (O_1667,N_12709,N_12109);
nor UO_1668 (O_1668,N_14324,N_14571);
or UO_1669 (O_1669,N_13927,N_12289);
or UO_1670 (O_1670,N_12371,N_12067);
nor UO_1671 (O_1671,N_12359,N_13484);
nand UO_1672 (O_1672,N_13989,N_14625);
nand UO_1673 (O_1673,N_13860,N_14380);
or UO_1674 (O_1674,N_14229,N_13085);
or UO_1675 (O_1675,N_13835,N_13533);
nand UO_1676 (O_1676,N_14673,N_12972);
and UO_1677 (O_1677,N_12902,N_14836);
nand UO_1678 (O_1678,N_14054,N_12267);
or UO_1679 (O_1679,N_12637,N_13480);
and UO_1680 (O_1680,N_14393,N_14511);
nand UO_1681 (O_1681,N_13537,N_14067);
nand UO_1682 (O_1682,N_12389,N_12570);
and UO_1683 (O_1683,N_12956,N_12938);
nand UO_1684 (O_1684,N_12988,N_13650);
or UO_1685 (O_1685,N_14649,N_14195);
or UO_1686 (O_1686,N_14792,N_14636);
and UO_1687 (O_1687,N_13655,N_12233);
and UO_1688 (O_1688,N_12068,N_13762);
nand UO_1689 (O_1689,N_14223,N_14437);
nor UO_1690 (O_1690,N_14964,N_12779);
nor UO_1691 (O_1691,N_14361,N_14656);
or UO_1692 (O_1692,N_13689,N_12189);
and UO_1693 (O_1693,N_13309,N_14962);
nor UO_1694 (O_1694,N_13293,N_13863);
nor UO_1695 (O_1695,N_14605,N_12909);
nand UO_1696 (O_1696,N_14073,N_14765);
xnor UO_1697 (O_1697,N_12575,N_14118);
or UO_1698 (O_1698,N_14241,N_13085);
and UO_1699 (O_1699,N_13184,N_13800);
nand UO_1700 (O_1700,N_12727,N_12470);
and UO_1701 (O_1701,N_14119,N_13222);
nor UO_1702 (O_1702,N_14466,N_13759);
and UO_1703 (O_1703,N_13161,N_13216);
nor UO_1704 (O_1704,N_12586,N_13373);
nor UO_1705 (O_1705,N_14874,N_14811);
nor UO_1706 (O_1706,N_13708,N_12059);
or UO_1707 (O_1707,N_13081,N_14129);
or UO_1708 (O_1708,N_13564,N_13004);
nor UO_1709 (O_1709,N_14343,N_14728);
nand UO_1710 (O_1710,N_13295,N_14961);
or UO_1711 (O_1711,N_14948,N_13884);
nand UO_1712 (O_1712,N_12466,N_13867);
xnor UO_1713 (O_1713,N_12167,N_13726);
nand UO_1714 (O_1714,N_14497,N_13759);
or UO_1715 (O_1715,N_14901,N_14696);
or UO_1716 (O_1716,N_12476,N_13063);
or UO_1717 (O_1717,N_12589,N_12825);
nor UO_1718 (O_1718,N_12308,N_14732);
nand UO_1719 (O_1719,N_12064,N_14642);
nand UO_1720 (O_1720,N_12934,N_12624);
or UO_1721 (O_1721,N_12646,N_12229);
nand UO_1722 (O_1722,N_14408,N_14572);
nor UO_1723 (O_1723,N_14148,N_12244);
nand UO_1724 (O_1724,N_13390,N_14464);
and UO_1725 (O_1725,N_12888,N_14034);
xnor UO_1726 (O_1726,N_13738,N_14134);
or UO_1727 (O_1727,N_13826,N_13787);
or UO_1728 (O_1728,N_14400,N_13303);
nand UO_1729 (O_1729,N_13693,N_13858);
and UO_1730 (O_1730,N_14140,N_12946);
or UO_1731 (O_1731,N_14332,N_13235);
or UO_1732 (O_1732,N_14639,N_13507);
and UO_1733 (O_1733,N_13253,N_13632);
or UO_1734 (O_1734,N_12858,N_13507);
and UO_1735 (O_1735,N_12063,N_12120);
and UO_1736 (O_1736,N_12628,N_13273);
or UO_1737 (O_1737,N_14947,N_12743);
and UO_1738 (O_1738,N_12040,N_13159);
and UO_1739 (O_1739,N_12205,N_12454);
or UO_1740 (O_1740,N_14471,N_13161);
or UO_1741 (O_1741,N_13824,N_13984);
and UO_1742 (O_1742,N_12969,N_13266);
nor UO_1743 (O_1743,N_14114,N_13620);
nand UO_1744 (O_1744,N_13937,N_13822);
or UO_1745 (O_1745,N_13306,N_14996);
xor UO_1746 (O_1746,N_12722,N_12929);
nor UO_1747 (O_1747,N_14579,N_14943);
nor UO_1748 (O_1748,N_14915,N_13180);
and UO_1749 (O_1749,N_14242,N_12988);
and UO_1750 (O_1750,N_14411,N_14783);
or UO_1751 (O_1751,N_13838,N_13496);
or UO_1752 (O_1752,N_13492,N_13395);
and UO_1753 (O_1753,N_14739,N_14634);
and UO_1754 (O_1754,N_13168,N_14622);
or UO_1755 (O_1755,N_12520,N_13583);
and UO_1756 (O_1756,N_13530,N_13578);
nor UO_1757 (O_1757,N_12083,N_12087);
nor UO_1758 (O_1758,N_14342,N_14264);
and UO_1759 (O_1759,N_12457,N_13599);
or UO_1760 (O_1760,N_13490,N_14318);
nand UO_1761 (O_1761,N_12411,N_13128);
and UO_1762 (O_1762,N_13661,N_12724);
nand UO_1763 (O_1763,N_14291,N_12810);
and UO_1764 (O_1764,N_13386,N_12559);
nand UO_1765 (O_1765,N_13283,N_14014);
nand UO_1766 (O_1766,N_12933,N_12792);
nor UO_1767 (O_1767,N_14081,N_12321);
nor UO_1768 (O_1768,N_14284,N_14276);
and UO_1769 (O_1769,N_13077,N_12858);
nor UO_1770 (O_1770,N_14947,N_12399);
xnor UO_1771 (O_1771,N_14282,N_14577);
or UO_1772 (O_1772,N_12793,N_12381);
and UO_1773 (O_1773,N_13631,N_12496);
nand UO_1774 (O_1774,N_13755,N_14390);
nor UO_1775 (O_1775,N_13612,N_14824);
and UO_1776 (O_1776,N_12249,N_14729);
nor UO_1777 (O_1777,N_14002,N_14391);
and UO_1778 (O_1778,N_12332,N_14089);
nand UO_1779 (O_1779,N_12702,N_12848);
nand UO_1780 (O_1780,N_13139,N_13863);
nor UO_1781 (O_1781,N_13183,N_14127);
nor UO_1782 (O_1782,N_14005,N_12816);
nor UO_1783 (O_1783,N_14382,N_13577);
nand UO_1784 (O_1784,N_13576,N_12434);
nand UO_1785 (O_1785,N_12198,N_13073);
nor UO_1786 (O_1786,N_12691,N_13606);
and UO_1787 (O_1787,N_12722,N_12265);
nand UO_1788 (O_1788,N_13309,N_14050);
nand UO_1789 (O_1789,N_13431,N_12052);
nor UO_1790 (O_1790,N_12877,N_12625);
nand UO_1791 (O_1791,N_14753,N_12085);
or UO_1792 (O_1792,N_12492,N_12489);
nor UO_1793 (O_1793,N_12109,N_12065);
or UO_1794 (O_1794,N_12221,N_13355);
and UO_1795 (O_1795,N_13643,N_12070);
or UO_1796 (O_1796,N_14578,N_12248);
or UO_1797 (O_1797,N_13627,N_14917);
nand UO_1798 (O_1798,N_13755,N_13212);
or UO_1799 (O_1799,N_14442,N_14295);
or UO_1800 (O_1800,N_12560,N_13244);
nand UO_1801 (O_1801,N_13419,N_13464);
and UO_1802 (O_1802,N_12777,N_13318);
nand UO_1803 (O_1803,N_13616,N_13582);
or UO_1804 (O_1804,N_14142,N_14462);
and UO_1805 (O_1805,N_14255,N_13610);
and UO_1806 (O_1806,N_14331,N_12478);
nand UO_1807 (O_1807,N_14427,N_13195);
nand UO_1808 (O_1808,N_14495,N_12091);
or UO_1809 (O_1809,N_14485,N_14643);
or UO_1810 (O_1810,N_12307,N_12864);
nor UO_1811 (O_1811,N_14179,N_12219);
nor UO_1812 (O_1812,N_12657,N_12341);
nand UO_1813 (O_1813,N_14993,N_13195);
and UO_1814 (O_1814,N_12090,N_13573);
and UO_1815 (O_1815,N_14779,N_13022);
and UO_1816 (O_1816,N_12394,N_12496);
or UO_1817 (O_1817,N_13450,N_12241);
nor UO_1818 (O_1818,N_13519,N_13277);
nor UO_1819 (O_1819,N_12884,N_14668);
or UO_1820 (O_1820,N_13040,N_14449);
xor UO_1821 (O_1821,N_14622,N_13654);
nand UO_1822 (O_1822,N_12148,N_12871);
and UO_1823 (O_1823,N_14942,N_14798);
nand UO_1824 (O_1824,N_13419,N_14349);
and UO_1825 (O_1825,N_14595,N_14840);
nand UO_1826 (O_1826,N_12071,N_14299);
and UO_1827 (O_1827,N_12657,N_12976);
or UO_1828 (O_1828,N_14555,N_13565);
nor UO_1829 (O_1829,N_14546,N_12754);
nand UO_1830 (O_1830,N_13113,N_14710);
or UO_1831 (O_1831,N_13503,N_13179);
nand UO_1832 (O_1832,N_14961,N_12207);
or UO_1833 (O_1833,N_14647,N_13679);
and UO_1834 (O_1834,N_14657,N_14270);
and UO_1835 (O_1835,N_14073,N_12852);
or UO_1836 (O_1836,N_13867,N_13763);
or UO_1837 (O_1837,N_12888,N_12311);
and UO_1838 (O_1838,N_14394,N_12305);
and UO_1839 (O_1839,N_12752,N_12902);
nand UO_1840 (O_1840,N_12737,N_14981);
or UO_1841 (O_1841,N_14841,N_14160);
nand UO_1842 (O_1842,N_14236,N_13817);
nand UO_1843 (O_1843,N_12300,N_13472);
nand UO_1844 (O_1844,N_13417,N_13957);
and UO_1845 (O_1845,N_13364,N_12879);
nand UO_1846 (O_1846,N_13556,N_14021);
nor UO_1847 (O_1847,N_13282,N_13083);
or UO_1848 (O_1848,N_13546,N_12025);
xnor UO_1849 (O_1849,N_14678,N_14577);
nand UO_1850 (O_1850,N_14373,N_14759);
nand UO_1851 (O_1851,N_14083,N_12631);
or UO_1852 (O_1852,N_13857,N_12140);
or UO_1853 (O_1853,N_13032,N_12771);
nor UO_1854 (O_1854,N_12959,N_13234);
nand UO_1855 (O_1855,N_12882,N_13949);
and UO_1856 (O_1856,N_12982,N_12406);
and UO_1857 (O_1857,N_13828,N_13499);
and UO_1858 (O_1858,N_12313,N_12949);
and UO_1859 (O_1859,N_13179,N_14917);
and UO_1860 (O_1860,N_12300,N_13213);
and UO_1861 (O_1861,N_13959,N_14150);
and UO_1862 (O_1862,N_12492,N_14355);
or UO_1863 (O_1863,N_13367,N_14633);
nand UO_1864 (O_1864,N_12533,N_12439);
and UO_1865 (O_1865,N_14639,N_14264);
nand UO_1866 (O_1866,N_12957,N_13808);
or UO_1867 (O_1867,N_13588,N_13511);
nor UO_1868 (O_1868,N_13424,N_14321);
and UO_1869 (O_1869,N_13704,N_14805);
nor UO_1870 (O_1870,N_13442,N_12697);
or UO_1871 (O_1871,N_13930,N_13459);
and UO_1872 (O_1872,N_14782,N_12374);
nor UO_1873 (O_1873,N_14080,N_12687);
nor UO_1874 (O_1874,N_13441,N_14189);
nand UO_1875 (O_1875,N_12631,N_14629);
and UO_1876 (O_1876,N_14527,N_13895);
or UO_1877 (O_1877,N_13471,N_13196);
and UO_1878 (O_1878,N_13077,N_12231);
nor UO_1879 (O_1879,N_12983,N_12839);
nor UO_1880 (O_1880,N_12251,N_14118);
nand UO_1881 (O_1881,N_12817,N_12973);
or UO_1882 (O_1882,N_14968,N_13354);
nand UO_1883 (O_1883,N_12289,N_13528);
and UO_1884 (O_1884,N_12067,N_13975);
nor UO_1885 (O_1885,N_12313,N_14161);
nand UO_1886 (O_1886,N_14789,N_12431);
and UO_1887 (O_1887,N_14427,N_13218);
or UO_1888 (O_1888,N_14821,N_14384);
or UO_1889 (O_1889,N_12491,N_13749);
nand UO_1890 (O_1890,N_12084,N_12673);
or UO_1891 (O_1891,N_12175,N_12161);
nand UO_1892 (O_1892,N_13820,N_14184);
nand UO_1893 (O_1893,N_12253,N_13021);
nand UO_1894 (O_1894,N_13019,N_13767);
or UO_1895 (O_1895,N_14913,N_14358);
and UO_1896 (O_1896,N_12562,N_14828);
nand UO_1897 (O_1897,N_13556,N_12731);
nand UO_1898 (O_1898,N_14611,N_14839);
nor UO_1899 (O_1899,N_13525,N_14511);
or UO_1900 (O_1900,N_13254,N_12249);
and UO_1901 (O_1901,N_13641,N_14773);
and UO_1902 (O_1902,N_14674,N_13801);
nand UO_1903 (O_1903,N_13772,N_14535);
or UO_1904 (O_1904,N_12024,N_12020);
or UO_1905 (O_1905,N_13360,N_13147);
nand UO_1906 (O_1906,N_14888,N_14855);
or UO_1907 (O_1907,N_12328,N_12504);
and UO_1908 (O_1908,N_12918,N_13211);
or UO_1909 (O_1909,N_14045,N_14455);
nor UO_1910 (O_1910,N_14166,N_14825);
nand UO_1911 (O_1911,N_14406,N_14930);
or UO_1912 (O_1912,N_14128,N_12898);
nor UO_1913 (O_1913,N_13084,N_13798);
or UO_1914 (O_1914,N_14924,N_12130);
nand UO_1915 (O_1915,N_12821,N_13778);
nor UO_1916 (O_1916,N_12492,N_13201);
and UO_1917 (O_1917,N_12809,N_13519);
nor UO_1918 (O_1918,N_14108,N_14257);
and UO_1919 (O_1919,N_13661,N_13092);
nand UO_1920 (O_1920,N_14331,N_13320);
nor UO_1921 (O_1921,N_12651,N_12618);
and UO_1922 (O_1922,N_13564,N_14044);
or UO_1923 (O_1923,N_13946,N_12624);
nand UO_1924 (O_1924,N_12485,N_14387);
or UO_1925 (O_1925,N_14239,N_13677);
or UO_1926 (O_1926,N_14342,N_12376);
or UO_1927 (O_1927,N_12792,N_12828);
nand UO_1928 (O_1928,N_14628,N_12655);
or UO_1929 (O_1929,N_13463,N_13329);
or UO_1930 (O_1930,N_12204,N_13669);
or UO_1931 (O_1931,N_12337,N_14954);
and UO_1932 (O_1932,N_12562,N_13358);
or UO_1933 (O_1933,N_13273,N_12915);
nor UO_1934 (O_1934,N_12812,N_13331);
nor UO_1935 (O_1935,N_13614,N_12986);
nand UO_1936 (O_1936,N_14789,N_12132);
or UO_1937 (O_1937,N_13831,N_12051);
nand UO_1938 (O_1938,N_14195,N_14596);
or UO_1939 (O_1939,N_12149,N_14621);
or UO_1940 (O_1940,N_14226,N_13077);
and UO_1941 (O_1941,N_13456,N_12575);
or UO_1942 (O_1942,N_12918,N_12783);
nand UO_1943 (O_1943,N_14210,N_13921);
or UO_1944 (O_1944,N_13570,N_12215);
and UO_1945 (O_1945,N_13805,N_13252);
nand UO_1946 (O_1946,N_13036,N_14891);
nand UO_1947 (O_1947,N_12447,N_14580);
or UO_1948 (O_1948,N_12492,N_12911);
or UO_1949 (O_1949,N_13558,N_14055);
nor UO_1950 (O_1950,N_12826,N_12487);
nand UO_1951 (O_1951,N_13076,N_14481);
nor UO_1952 (O_1952,N_13965,N_13719);
nand UO_1953 (O_1953,N_12793,N_14678);
nor UO_1954 (O_1954,N_14846,N_14273);
and UO_1955 (O_1955,N_14172,N_13147);
nor UO_1956 (O_1956,N_12020,N_13514);
or UO_1957 (O_1957,N_14312,N_13738);
nor UO_1958 (O_1958,N_12929,N_13350);
nor UO_1959 (O_1959,N_12219,N_12046);
and UO_1960 (O_1960,N_14366,N_14320);
and UO_1961 (O_1961,N_13461,N_14703);
nand UO_1962 (O_1962,N_12167,N_14330);
and UO_1963 (O_1963,N_14590,N_14016);
nand UO_1964 (O_1964,N_12929,N_12988);
or UO_1965 (O_1965,N_13087,N_14852);
or UO_1966 (O_1966,N_14595,N_14545);
and UO_1967 (O_1967,N_13664,N_13358);
xnor UO_1968 (O_1968,N_12312,N_13452);
nand UO_1969 (O_1969,N_13056,N_12391);
and UO_1970 (O_1970,N_14298,N_13876);
or UO_1971 (O_1971,N_12694,N_14335);
nand UO_1972 (O_1972,N_12274,N_12349);
nand UO_1973 (O_1973,N_14253,N_14310);
or UO_1974 (O_1974,N_13140,N_12962);
or UO_1975 (O_1975,N_12609,N_12423);
nor UO_1976 (O_1976,N_14497,N_13311);
nor UO_1977 (O_1977,N_13792,N_14810);
or UO_1978 (O_1978,N_12464,N_13396);
nand UO_1979 (O_1979,N_12504,N_14253);
nor UO_1980 (O_1980,N_13229,N_12501);
or UO_1981 (O_1981,N_14589,N_14294);
nand UO_1982 (O_1982,N_12183,N_12380);
nor UO_1983 (O_1983,N_13945,N_14340);
nor UO_1984 (O_1984,N_12354,N_14927);
nand UO_1985 (O_1985,N_13332,N_12645);
nand UO_1986 (O_1986,N_12041,N_14362);
and UO_1987 (O_1987,N_13055,N_13700);
nand UO_1988 (O_1988,N_13649,N_12748);
and UO_1989 (O_1989,N_14734,N_13212);
or UO_1990 (O_1990,N_12359,N_13399);
and UO_1991 (O_1991,N_14945,N_13131);
nand UO_1992 (O_1992,N_14874,N_14624);
nand UO_1993 (O_1993,N_14157,N_14159);
or UO_1994 (O_1994,N_14912,N_13192);
or UO_1995 (O_1995,N_13403,N_14908);
or UO_1996 (O_1996,N_14387,N_14911);
nor UO_1997 (O_1997,N_12312,N_13078);
nand UO_1998 (O_1998,N_14943,N_13266);
nor UO_1999 (O_1999,N_13586,N_14272);
endmodule