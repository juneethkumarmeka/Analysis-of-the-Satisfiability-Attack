module basic_1000_10000_1500_5_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_645,In_27);
nand U1 (N_1,In_804,In_278);
nand U2 (N_2,In_785,In_157);
nand U3 (N_3,In_184,In_255);
xor U4 (N_4,In_663,In_810);
nand U5 (N_5,In_846,In_742);
or U6 (N_6,In_658,In_973);
or U7 (N_7,In_272,In_829);
nand U8 (N_8,In_240,In_215);
nor U9 (N_9,In_35,In_950);
nor U10 (N_10,In_895,In_511);
and U11 (N_11,In_28,In_869);
nor U12 (N_12,In_942,In_294);
and U13 (N_13,In_794,In_261);
or U14 (N_14,In_33,In_669);
nand U15 (N_15,In_126,In_552);
nand U16 (N_16,In_471,In_466);
xnor U17 (N_17,In_981,In_15);
nor U18 (N_18,In_628,In_695);
nor U19 (N_19,In_750,In_102);
or U20 (N_20,In_17,In_745);
or U21 (N_21,In_786,In_237);
and U22 (N_22,In_822,In_39);
or U23 (N_23,In_44,In_680);
nand U24 (N_24,In_925,In_806);
nor U25 (N_25,In_916,In_905);
nor U26 (N_26,In_470,In_932);
nand U27 (N_27,In_716,In_53);
nand U28 (N_28,In_660,In_775);
nand U29 (N_29,In_275,In_351);
nor U30 (N_30,In_2,In_540);
nor U31 (N_31,In_762,In_222);
or U32 (N_32,In_591,In_779);
nand U33 (N_33,In_383,In_343);
or U34 (N_34,In_207,In_103);
or U35 (N_35,In_839,In_418);
or U36 (N_36,In_861,In_149);
nand U37 (N_37,In_532,In_163);
and U38 (N_38,In_263,In_605);
nor U39 (N_39,In_162,In_451);
and U40 (N_40,In_681,In_880);
and U41 (N_41,In_167,In_654);
or U42 (N_42,In_731,In_459);
or U43 (N_43,In_623,In_583);
or U44 (N_44,In_177,In_141);
nor U45 (N_45,In_937,In_843);
nor U46 (N_46,In_409,In_210);
or U47 (N_47,In_691,In_347);
or U48 (N_48,In_575,In_600);
nand U49 (N_49,In_538,In_514);
nor U50 (N_50,In_195,In_649);
and U51 (N_51,In_143,In_170);
nand U52 (N_52,In_465,In_105);
nand U53 (N_53,In_907,In_978);
and U54 (N_54,In_273,In_760);
and U55 (N_55,In_257,In_225);
or U56 (N_56,In_190,In_235);
nand U57 (N_57,In_624,In_239);
or U58 (N_58,In_543,In_191);
nand U59 (N_59,In_642,In_979);
and U60 (N_60,In_404,In_578);
xor U61 (N_61,In_783,In_574);
nor U62 (N_62,In_118,In_693);
and U63 (N_63,In_446,In_971);
nand U64 (N_64,In_307,In_0);
nand U65 (N_65,In_124,In_262);
and U66 (N_66,In_411,In_290);
and U67 (N_67,In_644,In_831);
or U68 (N_68,In_968,In_49);
nor U69 (N_69,In_505,In_635);
and U70 (N_70,In_919,In_121);
and U71 (N_71,In_595,In_65);
and U72 (N_72,In_111,In_677);
nand U73 (N_73,In_253,In_882);
nor U74 (N_74,In_577,In_276);
nand U75 (N_75,In_723,In_245);
or U76 (N_76,In_668,In_733);
or U77 (N_77,In_117,In_798);
nand U78 (N_78,In_369,In_682);
and U79 (N_79,In_868,In_867);
or U80 (N_80,In_939,In_833);
or U81 (N_81,In_771,In_803);
nand U82 (N_82,In_483,In_544);
nand U83 (N_83,In_581,In_510);
xnor U84 (N_84,In_468,In_325);
or U85 (N_85,In_728,In_489);
nand U86 (N_86,In_836,In_828);
nor U87 (N_87,In_479,In_431);
and U88 (N_88,In_440,In_554);
and U89 (N_89,In_396,In_493);
nor U90 (N_90,In_76,In_259);
and U91 (N_91,In_961,In_453);
and U92 (N_92,In_333,In_758);
nand U93 (N_93,In_346,In_722);
and U94 (N_94,In_309,In_40);
and U95 (N_95,In_280,In_789);
nor U96 (N_96,In_650,In_855);
and U97 (N_97,In_85,In_726);
nand U98 (N_98,In_107,In_952);
nor U99 (N_99,In_221,In_58);
or U100 (N_100,In_740,In_558);
and U101 (N_101,In_41,In_587);
nor U102 (N_102,In_11,In_871);
or U103 (N_103,In_189,In_454);
and U104 (N_104,In_357,In_705);
nor U105 (N_105,In_93,In_429);
or U106 (N_106,In_533,In_82);
nor U107 (N_107,In_365,In_529);
nand U108 (N_108,In_179,In_50);
or U109 (N_109,In_169,In_975);
and U110 (N_110,In_761,In_321);
or U111 (N_111,In_70,In_81);
nor U112 (N_112,In_661,In_603);
nand U113 (N_113,In_934,In_29);
nor U114 (N_114,In_545,In_592);
nor U115 (N_115,In_136,In_497);
and U116 (N_116,In_774,In_980);
and U117 (N_117,In_714,In_550);
or U118 (N_118,In_735,In_830);
nand U119 (N_119,In_399,In_612);
nor U120 (N_120,In_232,In_795);
or U121 (N_121,In_75,In_675);
nor U122 (N_122,In_371,In_182);
nand U123 (N_123,In_64,In_559);
nand U124 (N_124,In_523,In_66);
and U125 (N_125,In_525,In_341);
nor U126 (N_126,In_990,In_426);
xnor U127 (N_127,In_956,In_913);
nor U128 (N_128,In_361,In_911);
nand U129 (N_129,In_556,In_865);
nor U130 (N_130,In_817,In_436);
nor U131 (N_131,In_98,In_209);
nand U132 (N_132,In_339,In_110);
and U133 (N_133,In_776,In_873);
or U134 (N_134,In_694,In_992);
nor U135 (N_135,In_244,In_224);
nor U136 (N_136,In_18,In_666);
nor U137 (N_137,In_667,In_501);
and U138 (N_138,In_204,In_57);
nand U139 (N_139,In_770,In_355);
nand U140 (N_140,In_260,In_349);
nand U141 (N_141,In_315,In_945);
nor U142 (N_142,In_203,In_314);
and U143 (N_143,In_100,In_123);
or U144 (N_144,In_683,In_665);
xnor U145 (N_145,In_6,In_432);
nand U146 (N_146,In_879,In_460);
nor U147 (N_147,In_99,In_264);
and U148 (N_148,In_922,In_74);
and U149 (N_149,In_702,In_757);
nand U150 (N_150,In_211,In_270);
xor U151 (N_151,In_590,In_25);
nand U152 (N_152,In_94,In_381);
nor U153 (N_153,In_329,In_258);
and U154 (N_154,In_46,In_318);
nand U155 (N_155,In_827,In_863);
nand U156 (N_156,In_909,In_250);
and U157 (N_157,In_252,In_763);
nand U158 (N_158,In_697,In_542);
nor U159 (N_159,In_427,In_674);
or U160 (N_160,In_385,In_188);
nor U161 (N_161,In_551,In_9);
nand U162 (N_162,In_958,In_287);
nor U163 (N_163,In_151,In_21);
nor U164 (N_164,In_138,In_363);
or U165 (N_165,In_319,In_613);
nor U166 (N_166,In_793,In_130);
nor U167 (N_167,In_637,In_573);
or U168 (N_168,In_967,In_970);
nand U169 (N_169,In_180,In_835);
and U170 (N_170,In_298,In_653);
nor U171 (N_171,In_249,In_236);
and U172 (N_172,In_36,In_455);
nor U173 (N_173,In_824,In_502);
or U174 (N_174,In_481,In_320);
and U175 (N_175,In_288,In_24);
nand U176 (N_176,In_92,In_500);
or U177 (N_177,In_384,In_947);
or U178 (N_178,In_615,In_238);
or U179 (N_179,In_362,In_567);
or U180 (N_180,In_562,In_535);
nor U181 (N_181,In_488,In_487);
nand U182 (N_182,In_335,In_708);
nor U183 (N_183,In_208,In_128);
or U184 (N_184,In_580,In_368);
and U185 (N_185,In_62,In_622);
nor U186 (N_186,In_571,In_302);
or U187 (N_187,In_696,In_837);
and U188 (N_188,In_988,In_434);
nor U189 (N_189,In_698,In_484);
nor U190 (N_190,In_800,In_498);
and U191 (N_191,In_389,In_313);
or U192 (N_192,In_638,In_673);
and U193 (N_193,In_570,In_738);
nor U194 (N_194,In_308,In_269);
nand U195 (N_195,In_926,In_917);
or U196 (N_196,In_206,In_639);
or U197 (N_197,In_557,In_423);
nand U198 (N_198,In_334,In_568);
nand U199 (N_199,In_965,In_146);
nand U200 (N_200,In_393,In_936);
and U201 (N_201,In_183,In_812);
or U202 (N_202,In_340,In_614);
nor U203 (N_203,In_68,In_657);
nor U204 (N_204,In_796,In_651);
and U205 (N_205,In_688,In_175);
nor U206 (N_206,In_386,In_876);
nor U207 (N_207,In_864,In_854);
or U208 (N_208,In_946,In_524);
or U209 (N_209,In_89,In_825);
and U210 (N_210,In_555,In_491);
and U211 (N_211,In_312,In_150);
and U212 (N_212,In_442,In_108);
nor U213 (N_213,In_194,In_553);
and U214 (N_214,In_494,In_664);
and U215 (N_215,In_405,In_626);
nand U216 (N_216,In_91,In_202);
nand U217 (N_217,In_720,In_986);
or U218 (N_218,In_930,In_220);
nand U219 (N_219,In_621,In_63);
nand U220 (N_220,In_912,In_417);
nand U221 (N_221,In_569,In_515);
or U222 (N_222,In_690,In_743);
nand U223 (N_223,In_546,In_684);
or U224 (N_224,In_116,In_845);
or U225 (N_225,In_809,In_801);
nand U226 (N_226,In_853,In_754);
nand U227 (N_227,In_3,In_5);
or U228 (N_228,In_154,In_920);
or U229 (N_229,In_344,In_749);
nand U230 (N_230,In_462,In_306);
nand U231 (N_231,In_375,In_267);
nand U232 (N_232,In_181,In_407);
and U233 (N_233,In_327,In_242);
and U234 (N_234,In_671,In_509);
xnor U235 (N_235,In_474,In_142);
nor U236 (N_236,In_984,In_139);
xor U237 (N_237,In_633,In_802);
and U238 (N_238,In_486,In_160);
and U239 (N_239,In_449,In_84);
xnor U240 (N_240,In_337,In_928);
nor U241 (N_241,In_316,In_838);
and U242 (N_242,In_715,In_23);
and U243 (N_243,In_610,In_566);
nand U244 (N_244,In_200,In_201);
nand U245 (N_245,In_710,In_929);
nor U246 (N_246,In_292,In_480);
and U247 (N_247,In_692,In_799);
or U248 (N_248,In_137,In_286);
or U249 (N_249,In_174,In_834);
nor U250 (N_250,In_26,In_528);
nand U251 (N_251,In_890,In_406);
nor U252 (N_252,In_229,In_403);
and U253 (N_253,In_73,In_7);
and U254 (N_254,In_301,In_935);
nor U255 (N_255,In_214,In_281);
nor U256 (N_256,In_915,In_322);
xor U257 (N_257,In_437,In_901);
or U258 (N_258,In_45,In_59);
and U259 (N_259,In_37,In_963);
nand U260 (N_260,In_104,In_114);
and U261 (N_261,In_373,In_601);
nor U262 (N_262,In_790,In_408);
nand U263 (N_263,In_972,In_12);
nand U264 (N_264,In_711,In_140);
nand U265 (N_265,In_908,In_428);
and U266 (N_266,In_818,In_900);
nor U267 (N_267,In_196,In_55);
nand U268 (N_268,In_452,In_823);
nor U269 (N_269,In_461,In_976);
xnor U270 (N_270,In_456,In_1);
and U271 (N_271,In_994,In_561);
nor U272 (N_272,In_955,In_560);
and U273 (N_273,In_883,In_655);
xor U274 (N_274,In_629,In_927);
and U275 (N_275,In_966,In_858);
or U276 (N_276,In_862,In_526);
and U277 (N_277,In_739,In_377);
nor U278 (N_278,In_473,In_767);
nor U279 (N_279,In_962,In_844);
xnor U280 (N_280,In_80,In_69);
nand U281 (N_281,In_951,In_889);
nor U282 (N_282,In_134,In_997);
nor U283 (N_283,In_888,In_941);
nor U284 (N_284,In_378,In_8);
nor U285 (N_285,In_413,In_495);
nor U286 (N_286,In_672,In_820);
nand U287 (N_287,In_791,In_685);
nand U288 (N_288,In_331,In_686);
nand U289 (N_289,In_477,In_506);
xnor U290 (N_290,In_198,In_960);
nor U291 (N_291,In_747,In_875);
nand U292 (N_292,In_957,In_185);
or U293 (N_293,In_367,In_507);
nor U294 (N_294,In_416,In_51);
nand U295 (N_295,In_458,In_447);
or U296 (N_296,In_857,In_866);
nor U297 (N_297,In_689,In_326);
or U298 (N_298,In_643,In_152);
and U299 (N_299,In_819,In_166);
nor U300 (N_300,In_983,In_608);
or U301 (N_301,In_585,In_811);
and U302 (N_302,In_508,In_54);
nand U303 (N_303,In_527,In_119);
nand U304 (N_304,In_401,In_282);
nor U305 (N_305,In_77,In_289);
nor U306 (N_306,In_34,In_106);
nor U307 (N_307,In_759,In_332);
nor U308 (N_308,In_390,In_734);
and U309 (N_309,In_303,In_380);
or U310 (N_310,In_792,In_849);
nor U311 (N_311,In_707,In_859);
nor U312 (N_312,In_372,In_268);
nand U313 (N_313,In_522,In_701);
nor U314 (N_314,In_234,In_548);
nand U315 (N_315,In_159,In_353);
nor U316 (N_316,In_778,In_415);
and U317 (N_317,In_226,In_620);
nand U318 (N_318,In_874,In_4);
or U319 (N_319,In_475,In_959);
or U320 (N_320,In_704,In_359);
nor U321 (N_321,In_618,In_512);
and U322 (N_322,In_247,In_631);
and U323 (N_323,In_476,In_16);
nor U324 (N_324,In_72,In_354);
or U325 (N_325,In_485,In_850);
or U326 (N_326,In_814,In_88);
and U327 (N_327,In_444,In_732);
or U328 (N_328,In_109,In_158);
nor U329 (N_329,In_549,In_679);
or U330 (N_330,In_599,In_852);
nor U331 (N_331,In_254,In_582);
nand U332 (N_332,In_899,In_165);
and U333 (N_333,In_821,In_464);
or U334 (N_334,In_218,In_22);
nand U335 (N_335,In_921,In_903);
or U336 (N_336,In_518,In_816);
nor U337 (N_337,In_841,In_171);
nand U338 (N_338,In_872,In_145);
nand U339 (N_339,In_421,In_886);
nand U340 (N_340,In_588,In_719);
or U341 (N_341,In_898,In_617);
nand U342 (N_342,In_187,In_593);
nand U343 (N_343,In_212,In_517);
or U344 (N_344,In_777,In_634);
nor U345 (N_345,In_478,In_358);
nor U346 (N_346,In_176,In_893);
or U347 (N_347,In_297,In_519);
nand U348 (N_348,In_892,In_627);
nand U349 (N_349,In_96,In_987);
xor U350 (N_350,In_230,In_933);
nor U351 (N_351,In_42,In_414);
nor U352 (N_352,In_910,In_266);
or U353 (N_353,In_808,In_424);
and U354 (N_354,In_291,In_597);
and U355 (N_355,In_299,In_717);
nor U356 (N_356,In_199,In_95);
nand U357 (N_357,In_565,In_311);
nand U358 (N_358,In_989,In_161);
nor U359 (N_359,In_317,In_641);
nor U360 (N_360,In_410,In_376);
and U361 (N_361,In_67,In_305);
and U362 (N_362,In_700,In_769);
or U363 (N_363,In_310,In_382);
nand U364 (N_364,In_135,In_241);
nor U365 (N_365,In_216,In_61);
and U366 (N_366,In_894,In_101);
or U367 (N_367,In_931,In_178);
nor U368 (N_368,In_576,In_445);
nand U369 (N_369,In_729,In_30);
or U370 (N_370,In_656,In_205);
or U371 (N_371,In_632,In_129);
nor U372 (N_372,In_125,In_284);
and U373 (N_373,In_787,In_164);
nand U374 (N_374,In_231,In_646);
nand U375 (N_375,In_744,In_388);
nor U376 (N_376,In_330,In_884);
and U377 (N_377,In_586,In_147);
and U378 (N_378,In_847,In_725);
or U379 (N_379,In_496,In_718);
or U380 (N_380,In_596,In_400);
nor U381 (N_381,In_482,In_13);
nand U382 (N_382,In_441,In_896);
nor U383 (N_383,In_860,In_217);
nand U384 (N_384,In_438,In_56);
and U385 (N_385,In_598,In_492);
nand U386 (N_386,In_906,In_395);
or U387 (N_387,In_87,In_534);
nand U388 (N_388,In_589,In_513);
or U389 (N_389,In_594,In_856);
xor U390 (N_390,In_248,In_885);
nand U391 (N_391,In_848,In_998);
nand U392 (N_392,In_379,In_897);
nor U393 (N_393,In_788,In_625);
nand U394 (N_394,In_328,In_746);
or U395 (N_395,In_472,In_541);
nand U396 (N_396,In_826,In_619);
nand U397 (N_397,In_293,In_914);
or U398 (N_398,In_47,In_724);
or U399 (N_399,In_425,In_766);
nor U400 (N_400,In_748,In_607);
nor U401 (N_401,In_611,In_213);
xnor U402 (N_402,In_342,In_122);
or U403 (N_403,In_851,In_536);
nor U404 (N_404,In_904,In_435);
nor U405 (N_405,In_228,In_324);
nor U406 (N_406,In_647,In_153);
or U407 (N_407,In_348,In_422);
and U408 (N_408,In_797,In_842);
and U409 (N_409,In_687,In_420);
nor U410 (N_410,In_999,In_606);
nand U411 (N_411,In_659,In_48);
nand U412 (N_412,In_448,In_949);
xnor U413 (N_413,In_113,In_345);
or U414 (N_414,In_737,In_572);
and U415 (N_415,In_520,In_304);
nor U416 (N_416,In_784,In_991);
nor U417 (N_417,In_350,In_944);
and U418 (N_418,In_878,In_516);
and U419 (N_419,In_374,In_172);
and U420 (N_420,In_20,In_394);
and U421 (N_421,In_948,In_265);
and U422 (N_422,In_392,In_636);
nand U423 (N_423,In_813,In_387);
xnor U424 (N_424,In_336,In_450);
nor U425 (N_425,In_279,In_877);
nor U426 (N_426,In_223,In_736);
nor U427 (N_427,In_364,In_168);
nor U428 (N_428,In_870,In_765);
or U429 (N_429,In_727,In_300);
nor U430 (N_430,In_186,In_887);
or U431 (N_431,In_969,In_918);
or U432 (N_432,In_283,In_370);
or U433 (N_433,In_902,In_982);
and U434 (N_434,In_243,In_755);
or U435 (N_435,In_90,In_277);
and U436 (N_436,In_564,In_173);
or U437 (N_437,In_227,In_547);
and U438 (N_438,In_832,In_954);
or U439 (N_439,In_32,In_721);
and U440 (N_440,In_132,In_753);
nand U441 (N_441,In_219,In_996);
and U442 (N_442,In_953,In_14);
or U443 (N_443,In_499,In_604);
nand U444 (N_444,In_805,In_974);
or U445 (N_445,In_338,In_251);
nand U446 (N_446,In_768,In_352);
nor U447 (N_447,In_881,In_193);
xor U448 (N_448,In_148,In_616);
nor U449 (N_449,In_10,In_756);
nor U450 (N_450,In_156,In_670);
nor U451 (N_451,In_43,In_120);
nand U452 (N_452,In_530,In_430);
and U453 (N_453,In_412,In_133);
and U454 (N_454,In_891,In_295);
and U455 (N_455,In_964,In_246);
or U456 (N_456,In_741,In_60);
or U457 (N_457,In_31,In_433);
nand U458 (N_458,In_602,In_467);
and U459 (N_459,In_678,In_563);
or U460 (N_460,In_155,In_19);
and U461 (N_461,In_943,In_97);
nor U462 (N_462,In_706,In_764);
or U463 (N_463,In_938,In_995);
nand U464 (N_464,In_630,In_127);
or U465 (N_465,In_807,In_233);
nor U466 (N_466,In_391,In_38);
and U467 (N_467,In_131,In_985);
and U468 (N_468,In_356,In_52);
nand U469 (N_469,In_504,In_285);
nand U470 (N_470,In_752,In_923);
xnor U471 (N_471,In_662,In_579);
nand U472 (N_472,In_86,In_197);
or U473 (N_473,In_503,In_115);
and U474 (N_474,In_402,In_521);
nand U475 (N_475,In_730,In_144);
or U476 (N_476,In_703,In_709);
nor U477 (N_477,In_782,In_398);
nor U478 (N_478,In_457,In_751);
nor U479 (N_479,In_924,In_772);
or U480 (N_480,In_78,In_443);
nand U481 (N_481,In_323,In_439);
and U482 (N_482,In_584,In_71);
nor U483 (N_483,In_296,In_463);
nand U484 (N_484,In_699,In_648);
nand U485 (N_485,In_79,In_840);
nor U486 (N_486,In_609,In_713);
nand U487 (N_487,In_781,In_490);
nor U488 (N_488,In_397,In_360);
xnor U489 (N_489,In_112,In_815);
nand U490 (N_490,In_274,In_773);
nor U491 (N_491,In_676,In_993);
and U492 (N_492,In_712,In_977);
nand U493 (N_493,In_640,In_256);
nand U494 (N_494,In_531,In_537);
nor U495 (N_495,In_940,In_780);
nand U496 (N_496,In_539,In_192);
nor U497 (N_497,In_419,In_366);
or U498 (N_498,In_83,In_469);
nand U499 (N_499,In_271,In_652);
nor U500 (N_500,In_61,In_46);
and U501 (N_501,In_511,In_189);
nor U502 (N_502,In_772,In_49);
or U503 (N_503,In_271,In_57);
and U504 (N_504,In_376,In_165);
and U505 (N_505,In_775,In_883);
nor U506 (N_506,In_698,In_656);
or U507 (N_507,In_840,In_673);
nand U508 (N_508,In_370,In_138);
nand U509 (N_509,In_55,In_217);
or U510 (N_510,In_521,In_443);
nand U511 (N_511,In_887,In_909);
or U512 (N_512,In_884,In_55);
or U513 (N_513,In_132,In_644);
nand U514 (N_514,In_853,In_342);
and U515 (N_515,In_133,In_571);
nor U516 (N_516,In_390,In_91);
or U517 (N_517,In_37,In_604);
nor U518 (N_518,In_563,In_928);
nor U519 (N_519,In_527,In_958);
nor U520 (N_520,In_665,In_216);
nand U521 (N_521,In_463,In_282);
nand U522 (N_522,In_941,In_189);
and U523 (N_523,In_535,In_19);
or U524 (N_524,In_947,In_963);
nand U525 (N_525,In_862,In_712);
xor U526 (N_526,In_579,In_362);
and U527 (N_527,In_686,In_684);
xor U528 (N_528,In_611,In_563);
nor U529 (N_529,In_699,In_501);
nand U530 (N_530,In_261,In_109);
and U531 (N_531,In_678,In_478);
and U532 (N_532,In_808,In_222);
nand U533 (N_533,In_556,In_535);
nor U534 (N_534,In_757,In_552);
and U535 (N_535,In_650,In_380);
or U536 (N_536,In_698,In_939);
nor U537 (N_537,In_254,In_372);
or U538 (N_538,In_348,In_274);
or U539 (N_539,In_458,In_951);
xor U540 (N_540,In_757,In_902);
and U541 (N_541,In_289,In_348);
nand U542 (N_542,In_921,In_716);
xor U543 (N_543,In_58,In_614);
nor U544 (N_544,In_354,In_788);
nor U545 (N_545,In_705,In_120);
nor U546 (N_546,In_113,In_508);
nand U547 (N_547,In_179,In_227);
or U548 (N_548,In_692,In_195);
nor U549 (N_549,In_440,In_483);
nor U550 (N_550,In_348,In_832);
and U551 (N_551,In_280,In_340);
nand U552 (N_552,In_571,In_934);
or U553 (N_553,In_761,In_189);
nand U554 (N_554,In_847,In_643);
nor U555 (N_555,In_156,In_920);
nand U556 (N_556,In_328,In_545);
and U557 (N_557,In_995,In_587);
nand U558 (N_558,In_460,In_548);
nor U559 (N_559,In_711,In_554);
and U560 (N_560,In_379,In_38);
or U561 (N_561,In_759,In_93);
nor U562 (N_562,In_772,In_330);
nor U563 (N_563,In_615,In_402);
nand U564 (N_564,In_918,In_163);
or U565 (N_565,In_47,In_692);
or U566 (N_566,In_953,In_330);
nor U567 (N_567,In_905,In_770);
nor U568 (N_568,In_509,In_3);
or U569 (N_569,In_307,In_846);
nor U570 (N_570,In_133,In_687);
nand U571 (N_571,In_747,In_787);
xnor U572 (N_572,In_461,In_767);
nor U573 (N_573,In_333,In_608);
nor U574 (N_574,In_212,In_226);
or U575 (N_575,In_900,In_65);
nand U576 (N_576,In_131,In_457);
nor U577 (N_577,In_764,In_169);
and U578 (N_578,In_388,In_112);
xnor U579 (N_579,In_173,In_428);
nor U580 (N_580,In_922,In_11);
or U581 (N_581,In_417,In_178);
or U582 (N_582,In_157,In_16);
nand U583 (N_583,In_95,In_897);
and U584 (N_584,In_915,In_433);
or U585 (N_585,In_326,In_927);
or U586 (N_586,In_400,In_672);
or U587 (N_587,In_286,In_279);
nand U588 (N_588,In_808,In_507);
and U589 (N_589,In_577,In_449);
or U590 (N_590,In_586,In_941);
and U591 (N_591,In_641,In_13);
or U592 (N_592,In_672,In_537);
and U593 (N_593,In_821,In_55);
or U594 (N_594,In_299,In_576);
and U595 (N_595,In_668,In_163);
or U596 (N_596,In_987,In_461);
or U597 (N_597,In_915,In_628);
nor U598 (N_598,In_450,In_653);
nor U599 (N_599,In_950,In_349);
nand U600 (N_600,In_186,In_160);
or U601 (N_601,In_152,In_54);
xor U602 (N_602,In_135,In_643);
nor U603 (N_603,In_819,In_566);
and U604 (N_604,In_79,In_241);
nand U605 (N_605,In_391,In_97);
or U606 (N_606,In_357,In_944);
nand U607 (N_607,In_532,In_579);
nor U608 (N_608,In_972,In_407);
nor U609 (N_609,In_283,In_32);
and U610 (N_610,In_684,In_455);
or U611 (N_611,In_753,In_735);
and U612 (N_612,In_473,In_415);
and U613 (N_613,In_651,In_492);
and U614 (N_614,In_362,In_648);
and U615 (N_615,In_607,In_806);
nor U616 (N_616,In_824,In_458);
and U617 (N_617,In_325,In_729);
nand U618 (N_618,In_864,In_904);
nand U619 (N_619,In_787,In_580);
nor U620 (N_620,In_280,In_292);
nand U621 (N_621,In_731,In_615);
nand U622 (N_622,In_426,In_214);
nand U623 (N_623,In_778,In_85);
or U624 (N_624,In_377,In_980);
nor U625 (N_625,In_144,In_462);
nor U626 (N_626,In_646,In_684);
nand U627 (N_627,In_216,In_131);
or U628 (N_628,In_893,In_630);
nand U629 (N_629,In_638,In_399);
and U630 (N_630,In_960,In_253);
nor U631 (N_631,In_804,In_837);
or U632 (N_632,In_927,In_430);
or U633 (N_633,In_71,In_168);
nand U634 (N_634,In_667,In_341);
and U635 (N_635,In_275,In_731);
nand U636 (N_636,In_920,In_273);
and U637 (N_637,In_572,In_407);
nor U638 (N_638,In_764,In_522);
or U639 (N_639,In_949,In_170);
nand U640 (N_640,In_325,In_731);
or U641 (N_641,In_829,In_837);
nor U642 (N_642,In_234,In_840);
or U643 (N_643,In_237,In_980);
nand U644 (N_644,In_253,In_3);
and U645 (N_645,In_281,In_334);
nand U646 (N_646,In_869,In_418);
nand U647 (N_647,In_977,In_507);
and U648 (N_648,In_489,In_547);
nand U649 (N_649,In_317,In_370);
or U650 (N_650,In_337,In_250);
nand U651 (N_651,In_556,In_965);
and U652 (N_652,In_737,In_808);
or U653 (N_653,In_413,In_740);
and U654 (N_654,In_633,In_21);
and U655 (N_655,In_727,In_712);
nand U656 (N_656,In_712,In_898);
or U657 (N_657,In_622,In_865);
nand U658 (N_658,In_542,In_956);
or U659 (N_659,In_913,In_403);
and U660 (N_660,In_224,In_146);
nor U661 (N_661,In_927,In_29);
and U662 (N_662,In_544,In_912);
nor U663 (N_663,In_17,In_230);
nor U664 (N_664,In_95,In_761);
nor U665 (N_665,In_235,In_254);
nand U666 (N_666,In_474,In_233);
nor U667 (N_667,In_865,In_947);
or U668 (N_668,In_546,In_542);
nor U669 (N_669,In_680,In_375);
or U670 (N_670,In_372,In_452);
nand U671 (N_671,In_549,In_475);
nand U672 (N_672,In_325,In_862);
nor U673 (N_673,In_733,In_734);
or U674 (N_674,In_6,In_559);
and U675 (N_675,In_401,In_555);
nor U676 (N_676,In_128,In_190);
nor U677 (N_677,In_228,In_590);
or U678 (N_678,In_41,In_547);
and U679 (N_679,In_99,In_936);
nor U680 (N_680,In_802,In_932);
and U681 (N_681,In_796,In_946);
and U682 (N_682,In_620,In_184);
or U683 (N_683,In_22,In_976);
nand U684 (N_684,In_222,In_829);
or U685 (N_685,In_753,In_359);
or U686 (N_686,In_170,In_481);
nor U687 (N_687,In_250,In_66);
nor U688 (N_688,In_157,In_912);
or U689 (N_689,In_247,In_595);
nor U690 (N_690,In_52,In_967);
and U691 (N_691,In_550,In_523);
nand U692 (N_692,In_899,In_632);
nor U693 (N_693,In_146,In_386);
xnor U694 (N_694,In_646,In_595);
xnor U695 (N_695,In_202,In_979);
xor U696 (N_696,In_52,In_188);
or U697 (N_697,In_139,In_608);
nor U698 (N_698,In_31,In_922);
or U699 (N_699,In_400,In_514);
or U700 (N_700,In_863,In_857);
xnor U701 (N_701,In_776,In_314);
and U702 (N_702,In_798,In_988);
nand U703 (N_703,In_167,In_861);
xor U704 (N_704,In_990,In_703);
nor U705 (N_705,In_568,In_724);
nand U706 (N_706,In_545,In_392);
nor U707 (N_707,In_392,In_156);
and U708 (N_708,In_311,In_974);
and U709 (N_709,In_997,In_989);
or U710 (N_710,In_308,In_192);
and U711 (N_711,In_55,In_458);
and U712 (N_712,In_292,In_144);
nand U713 (N_713,In_46,In_704);
nor U714 (N_714,In_862,In_201);
nor U715 (N_715,In_72,In_703);
nand U716 (N_716,In_789,In_349);
and U717 (N_717,In_111,In_435);
xor U718 (N_718,In_143,In_129);
and U719 (N_719,In_468,In_459);
nor U720 (N_720,In_566,In_991);
or U721 (N_721,In_103,In_634);
nand U722 (N_722,In_986,In_321);
or U723 (N_723,In_269,In_154);
and U724 (N_724,In_468,In_485);
and U725 (N_725,In_713,In_62);
xnor U726 (N_726,In_314,In_480);
or U727 (N_727,In_150,In_890);
nand U728 (N_728,In_661,In_534);
and U729 (N_729,In_789,In_735);
or U730 (N_730,In_460,In_315);
and U731 (N_731,In_794,In_506);
nor U732 (N_732,In_565,In_10);
and U733 (N_733,In_246,In_24);
and U734 (N_734,In_461,In_712);
and U735 (N_735,In_853,In_388);
xor U736 (N_736,In_124,In_694);
and U737 (N_737,In_687,In_478);
or U738 (N_738,In_983,In_932);
nand U739 (N_739,In_870,In_237);
and U740 (N_740,In_187,In_431);
or U741 (N_741,In_324,In_249);
or U742 (N_742,In_755,In_840);
nand U743 (N_743,In_952,In_4);
nand U744 (N_744,In_8,In_978);
nor U745 (N_745,In_368,In_485);
and U746 (N_746,In_741,In_229);
nor U747 (N_747,In_117,In_824);
or U748 (N_748,In_287,In_380);
nand U749 (N_749,In_734,In_276);
nor U750 (N_750,In_774,In_773);
or U751 (N_751,In_929,In_146);
nand U752 (N_752,In_612,In_982);
nand U753 (N_753,In_394,In_954);
nor U754 (N_754,In_335,In_686);
nand U755 (N_755,In_733,In_356);
or U756 (N_756,In_354,In_883);
nand U757 (N_757,In_0,In_126);
nor U758 (N_758,In_943,In_634);
nand U759 (N_759,In_549,In_241);
or U760 (N_760,In_759,In_123);
nand U761 (N_761,In_406,In_872);
and U762 (N_762,In_718,In_896);
nor U763 (N_763,In_387,In_868);
nand U764 (N_764,In_696,In_966);
and U765 (N_765,In_407,In_630);
xnor U766 (N_766,In_443,In_223);
and U767 (N_767,In_715,In_759);
nor U768 (N_768,In_652,In_396);
nor U769 (N_769,In_809,In_228);
nor U770 (N_770,In_32,In_606);
nor U771 (N_771,In_398,In_926);
nor U772 (N_772,In_857,In_781);
and U773 (N_773,In_248,In_117);
or U774 (N_774,In_217,In_40);
and U775 (N_775,In_138,In_486);
and U776 (N_776,In_894,In_414);
nand U777 (N_777,In_97,In_961);
nand U778 (N_778,In_884,In_768);
and U779 (N_779,In_165,In_688);
and U780 (N_780,In_326,In_864);
and U781 (N_781,In_827,In_961);
nor U782 (N_782,In_471,In_151);
nor U783 (N_783,In_774,In_629);
and U784 (N_784,In_381,In_910);
and U785 (N_785,In_347,In_238);
nor U786 (N_786,In_114,In_536);
nand U787 (N_787,In_159,In_148);
nor U788 (N_788,In_298,In_905);
nor U789 (N_789,In_839,In_582);
nor U790 (N_790,In_816,In_683);
or U791 (N_791,In_205,In_406);
or U792 (N_792,In_952,In_299);
nor U793 (N_793,In_981,In_452);
or U794 (N_794,In_690,In_983);
or U795 (N_795,In_938,In_390);
and U796 (N_796,In_604,In_837);
and U797 (N_797,In_543,In_944);
nand U798 (N_798,In_572,In_515);
and U799 (N_799,In_606,In_601);
nor U800 (N_800,In_105,In_710);
or U801 (N_801,In_539,In_283);
nor U802 (N_802,In_37,In_862);
nand U803 (N_803,In_950,In_632);
or U804 (N_804,In_831,In_952);
or U805 (N_805,In_243,In_57);
nor U806 (N_806,In_768,In_623);
and U807 (N_807,In_777,In_617);
nand U808 (N_808,In_462,In_68);
and U809 (N_809,In_746,In_421);
or U810 (N_810,In_941,In_133);
nor U811 (N_811,In_330,In_615);
and U812 (N_812,In_90,In_717);
nor U813 (N_813,In_199,In_311);
nor U814 (N_814,In_508,In_804);
nor U815 (N_815,In_342,In_140);
and U816 (N_816,In_867,In_612);
or U817 (N_817,In_50,In_934);
nand U818 (N_818,In_859,In_335);
xnor U819 (N_819,In_499,In_59);
nand U820 (N_820,In_670,In_184);
nor U821 (N_821,In_561,In_839);
xnor U822 (N_822,In_469,In_466);
and U823 (N_823,In_333,In_165);
and U824 (N_824,In_722,In_514);
and U825 (N_825,In_823,In_566);
nand U826 (N_826,In_146,In_413);
and U827 (N_827,In_688,In_128);
and U828 (N_828,In_195,In_521);
or U829 (N_829,In_795,In_831);
xor U830 (N_830,In_114,In_425);
and U831 (N_831,In_335,In_74);
or U832 (N_832,In_604,In_934);
xnor U833 (N_833,In_418,In_331);
nand U834 (N_834,In_329,In_987);
or U835 (N_835,In_740,In_64);
nand U836 (N_836,In_562,In_350);
and U837 (N_837,In_257,In_446);
or U838 (N_838,In_679,In_926);
nand U839 (N_839,In_534,In_829);
or U840 (N_840,In_580,In_435);
nand U841 (N_841,In_935,In_173);
or U842 (N_842,In_17,In_630);
or U843 (N_843,In_758,In_365);
or U844 (N_844,In_998,In_805);
xnor U845 (N_845,In_683,In_227);
nor U846 (N_846,In_419,In_438);
nand U847 (N_847,In_392,In_663);
nand U848 (N_848,In_821,In_804);
or U849 (N_849,In_109,In_840);
and U850 (N_850,In_693,In_373);
or U851 (N_851,In_584,In_570);
nand U852 (N_852,In_533,In_928);
or U853 (N_853,In_786,In_969);
or U854 (N_854,In_458,In_753);
or U855 (N_855,In_966,In_606);
nand U856 (N_856,In_977,In_699);
or U857 (N_857,In_972,In_988);
nor U858 (N_858,In_470,In_795);
nor U859 (N_859,In_288,In_705);
nand U860 (N_860,In_112,In_469);
and U861 (N_861,In_272,In_884);
nor U862 (N_862,In_276,In_37);
nand U863 (N_863,In_505,In_937);
nand U864 (N_864,In_777,In_778);
and U865 (N_865,In_684,In_447);
nor U866 (N_866,In_410,In_161);
nor U867 (N_867,In_913,In_257);
or U868 (N_868,In_930,In_826);
and U869 (N_869,In_652,In_842);
xnor U870 (N_870,In_539,In_822);
nor U871 (N_871,In_647,In_497);
nor U872 (N_872,In_490,In_926);
nor U873 (N_873,In_244,In_400);
nand U874 (N_874,In_205,In_574);
nand U875 (N_875,In_987,In_4);
nor U876 (N_876,In_752,In_601);
or U877 (N_877,In_759,In_328);
or U878 (N_878,In_971,In_781);
nor U879 (N_879,In_899,In_652);
and U880 (N_880,In_70,In_587);
nand U881 (N_881,In_104,In_82);
and U882 (N_882,In_426,In_736);
and U883 (N_883,In_748,In_423);
nand U884 (N_884,In_622,In_502);
nor U885 (N_885,In_658,In_801);
nor U886 (N_886,In_584,In_722);
nand U887 (N_887,In_634,In_384);
nand U888 (N_888,In_40,In_500);
or U889 (N_889,In_888,In_262);
or U890 (N_890,In_801,In_611);
nand U891 (N_891,In_856,In_236);
nand U892 (N_892,In_781,In_725);
nor U893 (N_893,In_773,In_557);
nor U894 (N_894,In_59,In_660);
nor U895 (N_895,In_871,In_878);
nor U896 (N_896,In_914,In_52);
nor U897 (N_897,In_202,In_436);
nor U898 (N_898,In_491,In_479);
or U899 (N_899,In_594,In_242);
nand U900 (N_900,In_660,In_701);
nand U901 (N_901,In_78,In_201);
or U902 (N_902,In_215,In_737);
nand U903 (N_903,In_281,In_168);
nand U904 (N_904,In_83,In_493);
nand U905 (N_905,In_20,In_638);
nor U906 (N_906,In_523,In_855);
nor U907 (N_907,In_786,In_100);
and U908 (N_908,In_385,In_591);
nor U909 (N_909,In_423,In_928);
and U910 (N_910,In_967,In_888);
nor U911 (N_911,In_450,In_111);
or U912 (N_912,In_413,In_777);
and U913 (N_913,In_28,In_998);
nand U914 (N_914,In_104,In_116);
nand U915 (N_915,In_423,In_923);
nor U916 (N_916,In_142,In_314);
nand U917 (N_917,In_844,In_35);
and U918 (N_918,In_73,In_443);
nor U919 (N_919,In_11,In_256);
nor U920 (N_920,In_528,In_735);
or U921 (N_921,In_935,In_54);
nor U922 (N_922,In_476,In_764);
and U923 (N_923,In_641,In_928);
and U924 (N_924,In_824,In_329);
nor U925 (N_925,In_350,In_143);
nand U926 (N_926,In_781,In_999);
nor U927 (N_927,In_213,In_210);
and U928 (N_928,In_311,In_445);
and U929 (N_929,In_552,In_771);
nor U930 (N_930,In_634,In_189);
and U931 (N_931,In_904,In_428);
nand U932 (N_932,In_743,In_670);
or U933 (N_933,In_622,In_40);
and U934 (N_934,In_564,In_489);
nand U935 (N_935,In_88,In_563);
or U936 (N_936,In_392,In_396);
and U937 (N_937,In_438,In_280);
and U938 (N_938,In_905,In_394);
nand U939 (N_939,In_307,In_693);
xor U940 (N_940,In_484,In_380);
and U941 (N_941,In_429,In_112);
nor U942 (N_942,In_124,In_222);
nand U943 (N_943,In_541,In_836);
nor U944 (N_944,In_372,In_21);
or U945 (N_945,In_896,In_839);
nand U946 (N_946,In_246,In_706);
nand U947 (N_947,In_200,In_732);
nor U948 (N_948,In_615,In_877);
nand U949 (N_949,In_129,In_691);
nand U950 (N_950,In_574,In_998);
nor U951 (N_951,In_428,In_303);
and U952 (N_952,In_727,In_235);
nor U953 (N_953,In_302,In_204);
and U954 (N_954,In_360,In_65);
nand U955 (N_955,In_597,In_330);
or U956 (N_956,In_847,In_325);
or U957 (N_957,In_59,In_802);
and U958 (N_958,In_26,In_671);
and U959 (N_959,In_60,In_818);
or U960 (N_960,In_633,In_360);
nor U961 (N_961,In_848,In_628);
or U962 (N_962,In_982,In_85);
nand U963 (N_963,In_443,In_430);
and U964 (N_964,In_402,In_377);
nand U965 (N_965,In_9,In_368);
or U966 (N_966,In_576,In_895);
nand U967 (N_967,In_26,In_257);
or U968 (N_968,In_187,In_280);
or U969 (N_969,In_25,In_173);
or U970 (N_970,In_784,In_378);
nand U971 (N_971,In_257,In_319);
and U972 (N_972,In_31,In_437);
and U973 (N_973,In_619,In_175);
or U974 (N_974,In_908,In_528);
or U975 (N_975,In_383,In_310);
nand U976 (N_976,In_989,In_896);
and U977 (N_977,In_155,In_816);
and U978 (N_978,In_917,In_344);
nor U979 (N_979,In_835,In_266);
nand U980 (N_980,In_171,In_235);
and U981 (N_981,In_628,In_437);
nor U982 (N_982,In_893,In_362);
or U983 (N_983,In_814,In_2);
and U984 (N_984,In_438,In_342);
nor U985 (N_985,In_91,In_469);
or U986 (N_986,In_702,In_423);
nor U987 (N_987,In_793,In_205);
and U988 (N_988,In_608,In_960);
nor U989 (N_989,In_964,In_87);
nor U990 (N_990,In_961,In_294);
and U991 (N_991,In_555,In_311);
nor U992 (N_992,In_925,In_742);
nor U993 (N_993,In_362,In_809);
nor U994 (N_994,In_908,In_809);
nor U995 (N_995,In_787,In_153);
nand U996 (N_996,In_606,In_931);
or U997 (N_997,In_183,In_490);
nor U998 (N_998,In_396,In_784);
nand U999 (N_999,In_993,In_592);
nor U1000 (N_1000,In_158,In_196);
nand U1001 (N_1001,In_228,In_275);
and U1002 (N_1002,In_407,In_61);
or U1003 (N_1003,In_122,In_603);
or U1004 (N_1004,In_485,In_186);
nand U1005 (N_1005,In_42,In_512);
and U1006 (N_1006,In_854,In_459);
nand U1007 (N_1007,In_315,In_975);
nand U1008 (N_1008,In_625,In_584);
or U1009 (N_1009,In_409,In_159);
nand U1010 (N_1010,In_241,In_645);
nor U1011 (N_1011,In_669,In_84);
nand U1012 (N_1012,In_93,In_551);
or U1013 (N_1013,In_566,In_554);
nand U1014 (N_1014,In_934,In_242);
or U1015 (N_1015,In_177,In_117);
nor U1016 (N_1016,In_49,In_738);
nand U1017 (N_1017,In_717,In_875);
nor U1018 (N_1018,In_846,In_449);
nor U1019 (N_1019,In_512,In_835);
and U1020 (N_1020,In_431,In_995);
or U1021 (N_1021,In_609,In_541);
or U1022 (N_1022,In_738,In_290);
nor U1023 (N_1023,In_415,In_625);
nor U1024 (N_1024,In_51,In_617);
nand U1025 (N_1025,In_205,In_315);
nand U1026 (N_1026,In_682,In_160);
nor U1027 (N_1027,In_256,In_451);
xor U1028 (N_1028,In_137,In_269);
nand U1029 (N_1029,In_381,In_830);
nor U1030 (N_1030,In_564,In_417);
or U1031 (N_1031,In_450,In_994);
and U1032 (N_1032,In_14,In_574);
and U1033 (N_1033,In_419,In_148);
nor U1034 (N_1034,In_586,In_971);
xor U1035 (N_1035,In_733,In_438);
and U1036 (N_1036,In_521,In_880);
or U1037 (N_1037,In_101,In_656);
nand U1038 (N_1038,In_850,In_89);
and U1039 (N_1039,In_679,In_580);
and U1040 (N_1040,In_263,In_754);
and U1041 (N_1041,In_367,In_222);
or U1042 (N_1042,In_17,In_697);
nor U1043 (N_1043,In_716,In_130);
nand U1044 (N_1044,In_31,In_6);
and U1045 (N_1045,In_414,In_886);
and U1046 (N_1046,In_518,In_761);
and U1047 (N_1047,In_174,In_374);
nand U1048 (N_1048,In_31,In_617);
and U1049 (N_1049,In_720,In_450);
nor U1050 (N_1050,In_119,In_920);
nor U1051 (N_1051,In_769,In_308);
nand U1052 (N_1052,In_941,In_222);
and U1053 (N_1053,In_171,In_665);
and U1054 (N_1054,In_875,In_954);
nand U1055 (N_1055,In_415,In_103);
or U1056 (N_1056,In_202,In_9);
and U1057 (N_1057,In_785,In_434);
nor U1058 (N_1058,In_804,In_428);
or U1059 (N_1059,In_166,In_45);
or U1060 (N_1060,In_889,In_311);
nand U1061 (N_1061,In_105,In_884);
nor U1062 (N_1062,In_210,In_844);
or U1063 (N_1063,In_530,In_57);
and U1064 (N_1064,In_745,In_402);
nand U1065 (N_1065,In_620,In_155);
or U1066 (N_1066,In_513,In_719);
nor U1067 (N_1067,In_728,In_712);
nand U1068 (N_1068,In_86,In_733);
nor U1069 (N_1069,In_73,In_986);
or U1070 (N_1070,In_856,In_746);
and U1071 (N_1071,In_724,In_511);
or U1072 (N_1072,In_198,In_38);
and U1073 (N_1073,In_536,In_104);
and U1074 (N_1074,In_511,In_920);
nor U1075 (N_1075,In_323,In_471);
or U1076 (N_1076,In_572,In_360);
and U1077 (N_1077,In_752,In_794);
nand U1078 (N_1078,In_28,In_614);
nand U1079 (N_1079,In_897,In_152);
nor U1080 (N_1080,In_847,In_628);
nand U1081 (N_1081,In_321,In_477);
or U1082 (N_1082,In_17,In_953);
nor U1083 (N_1083,In_789,In_61);
or U1084 (N_1084,In_712,In_806);
nor U1085 (N_1085,In_553,In_433);
and U1086 (N_1086,In_179,In_352);
nand U1087 (N_1087,In_630,In_92);
nand U1088 (N_1088,In_671,In_537);
and U1089 (N_1089,In_676,In_70);
or U1090 (N_1090,In_120,In_754);
nor U1091 (N_1091,In_495,In_699);
and U1092 (N_1092,In_739,In_454);
and U1093 (N_1093,In_518,In_389);
and U1094 (N_1094,In_541,In_736);
and U1095 (N_1095,In_48,In_59);
nand U1096 (N_1096,In_300,In_958);
nand U1097 (N_1097,In_301,In_796);
and U1098 (N_1098,In_721,In_656);
or U1099 (N_1099,In_971,In_434);
and U1100 (N_1100,In_340,In_862);
nand U1101 (N_1101,In_450,In_138);
nand U1102 (N_1102,In_511,In_93);
and U1103 (N_1103,In_739,In_714);
or U1104 (N_1104,In_411,In_561);
nor U1105 (N_1105,In_6,In_226);
nand U1106 (N_1106,In_290,In_52);
xnor U1107 (N_1107,In_721,In_44);
and U1108 (N_1108,In_595,In_121);
nand U1109 (N_1109,In_951,In_948);
nor U1110 (N_1110,In_243,In_191);
or U1111 (N_1111,In_376,In_79);
nand U1112 (N_1112,In_900,In_312);
and U1113 (N_1113,In_62,In_278);
nand U1114 (N_1114,In_514,In_667);
and U1115 (N_1115,In_882,In_982);
and U1116 (N_1116,In_183,In_164);
nor U1117 (N_1117,In_533,In_72);
nand U1118 (N_1118,In_792,In_654);
nand U1119 (N_1119,In_564,In_726);
nand U1120 (N_1120,In_641,In_793);
and U1121 (N_1121,In_556,In_995);
nand U1122 (N_1122,In_451,In_693);
and U1123 (N_1123,In_723,In_670);
xnor U1124 (N_1124,In_158,In_581);
or U1125 (N_1125,In_561,In_590);
nand U1126 (N_1126,In_871,In_514);
nand U1127 (N_1127,In_923,In_603);
or U1128 (N_1128,In_854,In_327);
nand U1129 (N_1129,In_579,In_674);
and U1130 (N_1130,In_51,In_584);
nor U1131 (N_1131,In_896,In_220);
or U1132 (N_1132,In_33,In_4);
nor U1133 (N_1133,In_570,In_330);
and U1134 (N_1134,In_194,In_786);
nor U1135 (N_1135,In_439,In_897);
or U1136 (N_1136,In_578,In_685);
or U1137 (N_1137,In_195,In_107);
or U1138 (N_1138,In_860,In_696);
nor U1139 (N_1139,In_358,In_915);
and U1140 (N_1140,In_739,In_655);
nand U1141 (N_1141,In_491,In_327);
xor U1142 (N_1142,In_665,In_397);
nand U1143 (N_1143,In_687,In_622);
and U1144 (N_1144,In_172,In_222);
nor U1145 (N_1145,In_738,In_123);
nand U1146 (N_1146,In_884,In_67);
nor U1147 (N_1147,In_848,In_236);
and U1148 (N_1148,In_664,In_514);
nand U1149 (N_1149,In_806,In_542);
and U1150 (N_1150,In_38,In_676);
or U1151 (N_1151,In_932,In_892);
nand U1152 (N_1152,In_694,In_193);
or U1153 (N_1153,In_325,In_674);
nor U1154 (N_1154,In_65,In_48);
nand U1155 (N_1155,In_380,In_156);
nor U1156 (N_1156,In_701,In_436);
and U1157 (N_1157,In_550,In_292);
or U1158 (N_1158,In_717,In_946);
nor U1159 (N_1159,In_883,In_383);
or U1160 (N_1160,In_227,In_50);
and U1161 (N_1161,In_697,In_427);
and U1162 (N_1162,In_280,In_131);
nand U1163 (N_1163,In_830,In_351);
xnor U1164 (N_1164,In_648,In_754);
and U1165 (N_1165,In_855,In_752);
nor U1166 (N_1166,In_872,In_527);
or U1167 (N_1167,In_996,In_431);
nand U1168 (N_1168,In_23,In_999);
nor U1169 (N_1169,In_629,In_591);
nor U1170 (N_1170,In_636,In_849);
nand U1171 (N_1171,In_651,In_403);
nor U1172 (N_1172,In_357,In_432);
nor U1173 (N_1173,In_217,In_728);
nor U1174 (N_1174,In_247,In_390);
and U1175 (N_1175,In_727,In_221);
or U1176 (N_1176,In_678,In_220);
and U1177 (N_1177,In_64,In_860);
and U1178 (N_1178,In_920,In_533);
or U1179 (N_1179,In_204,In_426);
and U1180 (N_1180,In_480,In_913);
nor U1181 (N_1181,In_605,In_535);
nor U1182 (N_1182,In_269,In_279);
nand U1183 (N_1183,In_534,In_232);
or U1184 (N_1184,In_890,In_636);
or U1185 (N_1185,In_634,In_871);
nor U1186 (N_1186,In_247,In_839);
nand U1187 (N_1187,In_362,In_304);
nor U1188 (N_1188,In_28,In_246);
nand U1189 (N_1189,In_194,In_992);
nand U1190 (N_1190,In_514,In_467);
nor U1191 (N_1191,In_197,In_50);
nor U1192 (N_1192,In_793,In_729);
xor U1193 (N_1193,In_721,In_175);
or U1194 (N_1194,In_820,In_921);
nor U1195 (N_1195,In_839,In_713);
nor U1196 (N_1196,In_486,In_696);
and U1197 (N_1197,In_928,In_365);
or U1198 (N_1198,In_190,In_454);
nor U1199 (N_1199,In_19,In_150);
or U1200 (N_1200,In_387,In_99);
nand U1201 (N_1201,In_457,In_58);
or U1202 (N_1202,In_969,In_70);
or U1203 (N_1203,In_710,In_553);
nand U1204 (N_1204,In_138,In_22);
nor U1205 (N_1205,In_916,In_191);
and U1206 (N_1206,In_827,In_833);
nor U1207 (N_1207,In_117,In_10);
or U1208 (N_1208,In_336,In_8);
nor U1209 (N_1209,In_820,In_432);
nand U1210 (N_1210,In_781,In_840);
nor U1211 (N_1211,In_57,In_630);
or U1212 (N_1212,In_839,In_47);
nand U1213 (N_1213,In_266,In_333);
nand U1214 (N_1214,In_163,In_332);
and U1215 (N_1215,In_930,In_979);
and U1216 (N_1216,In_320,In_632);
nand U1217 (N_1217,In_779,In_942);
and U1218 (N_1218,In_520,In_998);
nor U1219 (N_1219,In_142,In_962);
and U1220 (N_1220,In_306,In_375);
nor U1221 (N_1221,In_916,In_177);
nor U1222 (N_1222,In_765,In_246);
and U1223 (N_1223,In_502,In_503);
nor U1224 (N_1224,In_592,In_401);
nor U1225 (N_1225,In_953,In_748);
nand U1226 (N_1226,In_896,In_760);
nand U1227 (N_1227,In_313,In_378);
nand U1228 (N_1228,In_367,In_624);
nor U1229 (N_1229,In_413,In_501);
and U1230 (N_1230,In_559,In_317);
nor U1231 (N_1231,In_861,In_380);
nand U1232 (N_1232,In_476,In_788);
nor U1233 (N_1233,In_734,In_273);
and U1234 (N_1234,In_714,In_557);
or U1235 (N_1235,In_337,In_678);
nor U1236 (N_1236,In_139,In_813);
nor U1237 (N_1237,In_328,In_756);
nand U1238 (N_1238,In_860,In_261);
or U1239 (N_1239,In_960,In_270);
and U1240 (N_1240,In_424,In_824);
or U1241 (N_1241,In_75,In_917);
nand U1242 (N_1242,In_833,In_349);
nand U1243 (N_1243,In_484,In_758);
nor U1244 (N_1244,In_940,In_357);
or U1245 (N_1245,In_550,In_254);
or U1246 (N_1246,In_807,In_39);
or U1247 (N_1247,In_97,In_823);
or U1248 (N_1248,In_515,In_989);
or U1249 (N_1249,In_247,In_774);
nand U1250 (N_1250,In_702,In_128);
nor U1251 (N_1251,In_22,In_922);
or U1252 (N_1252,In_522,In_945);
nand U1253 (N_1253,In_68,In_455);
nor U1254 (N_1254,In_105,In_390);
or U1255 (N_1255,In_396,In_437);
and U1256 (N_1256,In_410,In_901);
nand U1257 (N_1257,In_302,In_234);
and U1258 (N_1258,In_319,In_630);
and U1259 (N_1259,In_899,In_355);
or U1260 (N_1260,In_770,In_622);
and U1261 (N_1261,In_890,In_8);
or U1262 (N_1262,In_754,In_954);
nand U1263 (N_1263,In_553,In_871);
and U1264 (N_1264,In_727,In_511);
nor U1265 (N_1265,In_302,In_15);
nand U1266 (N_1266,In_156,In_326);
nand U1267 (N_1267,In_385,In_356);
or U1268 (N_1268,In_932,In_474);
or U1269 (N_1269,In_119,In_581);
and U1270 (N_1270,In_755,In_409);
or U1271 (N_1271,In_469,In_262);
nand U1272 (N_1272,In_232,In_370);
xnor U1273 (N_1273,In_98,In_545);
nand U1274 (N_1274,In_143,In_332);
or U1275 (N_1275,In_325,In_827);
nand U1276 (N_1276,In_806,In_672);
and U1277 (N_1277,In_944,In_235);
and U1278 (N_1278,In_62,In_488);
or U1279 (N_1279,In_829,In_939);
nand U1280 (N_1280,In_789,In_484);
and U1281 (N_1281,In_655,In_433);
and U1282 (N_1282,In_93,In_422);
nor U1283 (N_1283,In_809,In_529);
and U1284 (N_1284,In_331,In_361);
nor U1285 (N_1285,In_803,In_512);
and U1286 (N_1286,In_73,In_141);
nor U1287 (N_1287,In_855,In_432);
nor U1288 (N_1288,In_11,In_497);
nor U1289 (N_1289,In_633,In_699);
nand U1290 (N_1290,In_861,In_571);
nor U1291 (N_1291,In_211,In_992);
nand U1292 (N_1292,In_527,In_303);
or U1293 (N_1293,In_440,In_148);
or U1294 (N_1294,In_776,In_3);
nor U1295 (N_1295,In_475,In_258);
and U1296 (N_1296,In_969,In_348);
nor U1297 (N_1297,In_177,In_732);
nand U1298 (N_1298,In_576,In_682);
xnor U1299 (N_1299,In_810,In_94);
nand U1300 (N_1300,In_654,In_426);
xnor U1301 (N_1301,In_177,In_160);
nor U1302 (N_1302,In_164,In_397);
nor U1303 (N_1303,In_160,In_369);
nand U1304 (N_1304,In_755,In_514);
nor U1305 (N_1305,In_559,In_809);
nand U1306 (N_1306,In_589,In_173);
and U1307 (N_1307,In_840,In_287);
nand U1308 (N_1308,In_645,In_510);
or U1309 (N_1309,In_185,In_751);
and U1310 (N_1310,In_24,In_162);
and U1311 (N_1311,In_955,In_454);
nand U1312 (N_1312,In_813,In_53);
and U1313 (N_1313,In_635,In_745);
nor U1314 (N_1314,In_739,In_266);
xor U1315 (N_1315,In_236,In_776);
or U1316 (N_1316,In_392,In_637);
and U1317 (N_1317,In_891,In_637);
nand U1318 (N_1318,In_461,In_649);
nand U1319 (N_1319,In_333,In_706);
and U1320 (N_1320,In_539,In_740);
nor U1321 (N_1321,In_582,In_833);
nor U1322 (N_1322,In_514,In_224);
and U1323 (N_1323,In_622,In_608);
nor U1324 (N_1324,In_525,In_803);
and U1325 (N_1325,In_751,In_551);
nor U1326 (N_1326,In_487,In_417);
nor U1327 (N_1327,In_895,In_878);
nor U1328 (N_1328,In_643,In_301);
nor U1329 (N_1329,In_519,In_44);
or U1330 (N_1330,In_537,In_618);
or U1331 (N_1331,In_664,In_946);
xnor U1332 (N_1332,In_913,In_838);
and U1333 (N_1333,In_356,In_679);
nand U1334 (N_1334,In_371,In_664);
and U1335 (N_1335,In_108,In_387);
nor U1336 (N_1336,In_322,In_554);
nand U1337 (N_1337,In_807,In_791);
and U1338 (N_1338,In_956,In_759);
or U1339 (N_1339,In_991,In_479);
nand U1340 (N_1340,In_634,In_768);
nor U1341 (N_1341,In_328,In_444);
nand U1342 (N_1342,In_358,In_888);
nand U1343 (N_1343,In_876,In_561);
nor U1344 (N_1344,In_70,In_445);
and U1345 (N_1345,In_440,In_912);
nand U1346 (N_1346,In_832,In_26);
or U1347 (N_1347,In_589,In_409);
nand U1348 (N_1348,In_139,In_973);
nor U1349 (N_1349,In_407,In_80);
nor U1350 (N_1350,In_476,In_464);
or U1351 (N_1351,In_862,In_448);
nand U1352 (N_1352,In_759,In_115);
nand U1353 (N_1353,In_444,In_456);
or U1354 (N_1354,In_621,In_198);
or U1355 (N_1355,In_620,In_618);
and U1356 (N_1356,In_367,In_602);
nor U1357 (N_1357,In_515,In_182);
nor U1358 (N_1358,In_765,In_495);
or U1359 (N_1359,In_193,In_142);
nor U1360 (N_1360,In_530,In_626);
and U1361 (N_1361,In_92,In_403);
or U1362 (N_1362,In_71,In_870);
xnor U1363 (N_1363,In_487,In_183);
or U1364 (N_1364,In_792,In_668);
or U1365 (N_1365,In_345,In_198);
and U1366 (N_1366,In_427,In_443);
or U1367 (N_1367,In_776,In_108);
or U1368 (N_1368,In_537,In_344);
nand U1369 (N_1369,In_201,In_514);
nand U1370 (N_1370,In_787,In_659);
nor U1371 (N_1371,In_60,In_180);
or U1372 (N_1372,In_890,In_786);
or U1373 (N_1373,In_32,In_854);
or U1374 (N_1374,In_750,In_494);
and U1375 (N_1375,In_978,In_639);
nand U1376 (N_1376,In_308,In_974);
nand U1377 (N_1377,In_111,In_441);
nor U1378 (N_1378,In_211,In_218);
or U1379 (N_1379,In_613,In_637);
and U1380 (N_1380,In_706,In_956);
nand U1381 (N_1381,In_812,In_961);
nor U1382 (N_1382,In_842,In_383);
nor U1383 (N_1383,In_737,In_296);
and U1384 (N_1384,In_725,In_41);
and U1385 (N_1385,In_902,In_479);
nor U1386 (N_1386,In_252,In_743);
nand U1387 (N_1387,In_676,In_880);
nor U1388 (N_1388,In_37,In_541);
nand U1389 (N_1389,In_671,In_973);
and U1390 (N_1390,In_732,In_269);
nand U1391 (N_1391,In_121,In_614);
or U1392 (N_1392,In_410,In_534);
or U1393 (N_1393,In_45,In_208);
and U1394 (N_1394,In_913,In_589);
or U1395 (N_1395,In_35,In_568);
and U1396 (N_1396,In_307,In_857);
xor U1397 (N_1397,In_391,In_341);
nor U1398 (N_1398,In_129,In_256);
nor U1399 (N_1399,In_188,In_612);
nor U1400 (N_1400,In_128,In_199);
nor U1401 (N_1401,In_766,In_358);
nor U1402 (N_1402,In_167,In_386);
and U1403 (N_1403,In_585,In_759);
or U1404 (N_1404,In_163,In_398);
or U1405 (N_1405,In_751,In_81);
nor U1406 (N_1406,In_230,In_332);
nor U1407 (N_1407,In_990,In_238);
or U1408 (N_1408,In_976,In_670);
nand U1409 (N_1409,In_124,In_558);
and U1410 (N_1410,In_954,In_717);
or U1411 (N_1411,In_74,In_28);
or U1412 (N_1412,In_534,In_82);
and U1413 (N_1413,In_423,In_353);
nand U1414 (N_1414,In_464,In_342);
nand U1415 (N_1415,In_843,In_692);
nand U1416 (N_1416,In_356,In_204);
nor U1417 (N_1417,In_506,In_722);
or U1418 (N_1418,In_458,In_492);
and U1419 (N_1419,In_838,In_587);
nor U1420 (N_1420,In_322,In_429);
nand U1421 (N_1421,In_491,In_5);
nand U1422 (N_1422,In_458,In_836);
or U1423 (N_1423,In_703,In_988);
nor U1424 (N_1424,In_952,In_371);
nor U1425 (N_1425,In_781,In_107);
nand U1426 (N_1426,In_802,In_43);
or U1427 (N_1427,In_629,In_8);
nand U1428 (N_1428,In_559,In_623);
nor U1429 (N_1429,In_344,In_472);
nand U1430 (N_1430,In_422,In_731);
and U1431 (N_1431,In_634,In_472);
or U1432 (N_1432,In_424,In_280);
and U1433 (N_1433,In_873,In_358);
nand U1434 (N_1434,In_659,In_928);
nor U1435 (N_1435,In_803,In_495);
and U1436 (N_1436,In_422,In_746);
and U1437 (N_1437,In_738,In_790);
and U1438 (N_1438,In_981,In_961);
nand U1439 (N_1439,In_448,In_761);
nand U1440 (N_1440,In_345,In_425);
and U1441 (N_1441,In_310,In_891);
and U1442 (N_1442,In_969,In_165);
nor U1443 (N_1443,In_420,In_938);
or U1444 (N_1444,In_817,In_912);
and U1445 (N_1445,In_118,In_500);
nand U1446 (N_1446,In_412,In_491);
and U1447 (N_1447,In_870,In_232);
and U1448 (N_1448,In_290,In_74);
nor U1449 (N_1449,In_954,In_101);
and U1450 (N_1450,In_427,In_23);
or U1451 (N_1451,In_163,In_620);
or U1452 (N_1452,In_666,In_393);
nor U1453 (N_1453,In_644,In_308);
nand U1454 (N_1454,In_503,In_988);
or U1455 (N_1455,In_131,In_984);
or U1456 (N_1456,In_583,In_335);
and U1457 (N_1457,In_371,In_141);
nor U1458 (N_1458,In_480,In_714);
or U1459 (N_1459,In_870,In_0);
and U1460 (N_1460,In_349,In_370);
nor U1461 (N_1461,In_240,In_49);
nor U1462 (N_1462,In_45,In_542);
or U1463 (N_1463,In_858,In_948);
and U1464 (N_1464,In_775,In_32);
nand U1465 (N_1465,In_118,In_727);
xnor U1466 (N_1466,In_5,In_852);
nand U1467 (N_1467,In_588,In_301);
xor U1468 (N_1468,In_84,In_973);
or U1469 (N_1469,In_248,In_6);
nand U1470 (N_1470,In_364,In_756);
xor U1471 (N_1471,In_116,In_50);
nor U1472 (N_1472,In_785,In_837);
and U1473 (N_1473,In_202,In_807);
nand U1474 (N_1474,In_904,In_759);
nand U1475 (N_1475,In_428,In_320);
and U1476 (N_1476,In_663,In_782);
nand U1477 (N_1477,In_192,In_161);
nand U1478 (N_1478,In_309,In_253);
nand U1479 (N_1479,In_930,In_678);
or U1480 (N_1480,In_401,In_939);
or U1481 (N_1481,In_79,In_143);
nand U1482 (N_1482,In_835,In_766);
nand U1483 (N_1483,In_691,In_196);
or U1484 (N_1484,In_188,In_540);
or U1485 (N_1485,In_85,In_754);
nor U1486 (N_1486,In_596,In_603);
and U1487 (N_1487,In_593,In_10);
or U1488 (N_1488,In_151,In_582);
nor U1489 (N_1489,In_825,In_785);
nand U1490 (N_1490,In_119,In_553);
xnor U1491 (N_1491,In_141,In_242);
nor U1492 (N_1492,In_326,In_178);
and U1493 (N_1493,In_76,In_998);
and U1494 (N_1494,In_726,In_455);
nor U1495 (N_1495,In_617,In_141);
nand U1496 (N_1496,In_187,In_216);
or U1497 (N_1497,In_98,In_716);
or U1498 (N_1498,In_496,In_180);
nand U1499 (N_1499,In_381,In_486);
nand U1500 (N_1500,In_89,In_989);
or U1501 (N_1501,In_543,In_211);
and U1502 (N_1502,In_299,In_30);
and U1503 (N_1503,In_456,In_260);
nor U1504 (N_1504,In_150,In_949);
and U1505 (N_1505,In_402,In_24);
nand U1506 (N_1506,In_641,In_985);
nand U1507 (N_1507,In_207,In_322);
and U1508 (N_1508,In_597,In_849);
nor U1509 (N_1509,In_458,In_594);
or U1510 (N_1510,In_147,In_165);
nand U1511 (N_1511,In_279,In_264);
nand U1512 (N_1512,In_892,In_173);
and U1513 (N_1513,In_388,In_770);
and U1514 (N_1514,In_579,In_851);
or U1515 (N_1515,In_20,In_92);
nor U1516 (N_1516,In_459,In_573);
nor U1517 (N_1517,In_521,In_747);
and U1518 (N_1518,In_720,In_109);
nand U1519 (N_1519,In_101,In_351);
or U1520 (N_1520,In_674,In_64);
nor U1521 (N_1521,In_824,In_234);
nor U1522 (N_1522,In_36,In_623);
nor U1523 (N_1523,In_408,In_300);
nand U1524 (N_1524,In_941,In_731);
and U1525 (N_1525,In_626,In_428);
nand U1526 (N_1526,In_737,In_35);
and U1527 (N_1527,In_597,In_550);
nand U1528 (N_1528,In_760,In_980);
or U1529 (N_1529,In_743,In_318);
and U1530 (N_1530,In_256,In_880);
nor U1531 (N_1531,In_188,In_171);
nor U1532 (N_1532,In_965,In_199);
and U1533 (N_1533,In_994,In_998);
or U1534 (N_1534,In_308,In_155);
or U1535 (N_1535,In_30,In_979);
and U1536 (N_1536,In_83,In_703);
nor U1537 (N_1537,In_546,In_97);
and U1538 (N_1538,In_603,In_38);
nor U1539 (N_1539,In_68,In_385);
or U1540 (N_1540,In_597,In_154);
nor U1541 (N_1541,In_561,In_758);
and U1542 (N_1542,In_232,In_358);
and U1543 (N_1543,In_232,In_424);
and U1544 (N_1544,In_850,In_456);
or U1545 (N_1545,In_578,In_462);
nor U1546 (N_1546,In_266,In_533);
and U1547 (N_1547,In_528,In_603);
nor U1548 (N_1548,In_936,In_451);
or U1549 (N_1549,In_830,In_255);
nor U1550 (N_1550,In_180,In_111);
nand U1551 (N_1551,In_941,In_239);
nand U1552 (N_1552,In_981,In_561);
nand U1553 (N_1553,In_425,In_250);
or U1554 (N_1554,In_820,In_994);
and U1555 (N_1555,In_115,In_996);
nor U1556 (N_1556,In_335,In_924);
nand U1557 (N_1557,In_126,In_239);
or U1558 (N_1558,In_103,In_270);
and U1559 (N_1559,In_552,In_484);
and U1560 (N_1560,In_431,In_567);
and U1561 (N_1561,In_975,In_333);
and U1562 (N_1562,In_90,In_831);
or U1563 (N_1563,In_253,In_911);
or U1564 (N_1564,In_741,In_341);
or U1565 (N_1565,In_231,In_379);
and U1566 (N_1566,In_498,In_513);
nand U1567 (N_1567,In_739,In_756);
nor U1568 (N_1568,In_754,In_21);
nor U1569 (N_1569,In_962,In_184);
nor U1570 (N_1570,In_252,In_166);
nor U1571 (N_1571,In_211,In_551);
xor U1572 (N_1572,In_409,In_548);
nor U1573 (N_1573,In_679,In_909);
xnor U1574 (N_1574,In_582,In_627);
nor U1575 (N_1575,In_842,In_536);
nor U1576 (N_1576,In_867,In_621);
nor U1577 (N_1577,In_577,In_877);
or U1578 (N_1578,In_939,In_295);
or U1579 (N_1579,In_453,In_784);
nor U1580 (N_1580,In_94,In_654);
nor U1581 (N_1581,In_866,In_334);
and U1582 (N_1582,In_464,In_238);
xor U1583 (N_1583,In_502,In_404);
nor U1584 (N_1584,In_968,In_61);
and U1585 (N_1585,In_411,In_927);
or U1586 (N_1586,In_699,In_115);
nor U1587 (N_1587,In_780,In_214);
nand U1588 (N_1588,In_266,In_677);
nand U1589 (N_1589,In_357,In_296);
and U1590 (N_1590,In_586,In_705);
nand U1591 (N_1591,In_866,In_657);
and U1592 (N_1592,In_557,In_659);
or U1593 (N_1593,In_837,In_30);
nor U1594 (N_1594,In_869,In_698);
nor U1595 (N_1595,In_284,In_116);
nand U1596 (N_1596,In_155,In_48);
nand U1597 (N_1597,In_596,In_707);
nor U1598 (N_1598,In_468,In_719);
nand U1599 (N_1599,In_525,In_275);
nand U1600 (N_1600,In_928,In_254);
and U1601 (N_1601,In_276,In_245);
or U1602 (N_1602,In_352,In_172);
nor U1603 (N_1603,In_941,In_464);
nand U1604 (N_1604,In_841,In_886);
nor U1605 (N_1605,In_103,In_828);
nand U1606 (N_1606,In_983,In_17);
nand U1607 (N_1607,In_474,In_588);
and U1608 (N_1608,In_923,In_698);
nand U1609 (N_1609,In_549,In_370);
nand U1610 (N_1610,In_767,In_551);
or U1611 (N_1611,In_545,In_31);
nand U1612 (N_1612,In_424,In_239);
or U1613 (N_1613,In_859,In_958);
nand U1614 (N_1614,In_537,In_842);
or U1615 (N_1615,In_586,In_998);
nor U1616 (N_1616,In_341,In_949);
nor U1617 (N_1617,In_823,In_881);
nand U1618 (N_1618,In_897,In_438);
nor U1619 (N_1619,In_218,In_584);
or U1620 (N_1620,In_895,In_253);
nor U1621 (N_1621,In_964,In_541);
and U1622 (N_1622,In_797,In_578);
or U1623 (N_1623,In_66,In_601);
or U1624 (N_1624,In_458,In_693);
and U1625 (N_1625,In_295,In_323);
nand U1626 (N_1626,In_623,In_26);
nor U1627 (N_1627,In_212,In_252);
nand U1628 (N_1628,In_517,In_488);
nor U1629 (N_1629,In_801,In_55);
and U1630 (N_1630,In_907,In_548);
nor U1631 (N_1631,In_171,In_868);
nand U1632 (N_1632,In_808,In_100);
nor U1633 (N_1633,In_130,In_291);
or U1634 (N_1634,In_173,In_702);
nand U1635 (N_1635,In_866,In_327);
and U1636 (N_1636,In_477,In_2);
nand U1637 (N_1637,In_357,In_186);
and U1638 (N_1638,In_748,In_419);
nand U1639 (N_1639,In_838,In_949);
nand U1640 (N_1640,In_262,In_514);
and U1641 (N_1641,In_486,In_291);
nand U1642 (N_1642,In_686,In_279);
nand U1643 (N_1643,In_355,In_835);
xnor U1644 (N_1644,In_697,In_181);
nand U1645 (N_1645,In_123,In_893);
or U1646 (N_1646,In_48,In_862);
and U1647 (N_1647,In_47,In_525);
nor U1648 (N_1648,In_866,In_494);
or U1649 (N_1649,In_466,In_129);
or U1650 (N_1650,In_746,In_630);
or U1651 (N_1651,In_710,In_315);
nor U1652 (N_1652,In_737,In_928);
or U1653 (N_1653,In_955,In_536);
and U1654 (N_1654,In_201,In_374);
and U1655 (N_1655,In_27,In_390);
or U1656 (N_1656,In_863,In_954);
or U1657 (N_1657,In_710,In_285);
nand U1658 (N_1658,In_709,In_933);
xnor U1659 (N_1659,In_758,In_895);
and U1660 (N_1660,In_242,In_632);
or U1661 (N_1661,In_47,In_42);
nand U1662 (N_1662,In_145,In_649);
nor U1663 (N_1663,In_979,In_613);
nor U1664 (N_1664,In_39,In_954);
and U1665 (N_1665,In_75,In_216);
and U1666 (N_1666,In_917,In_777);
nand U1667 (N_1667,In_506,In_689);
nand U1668 (N_1668,In_950,In_945);
or U1669 (N_1669,In_98,In_63);
nand U1670 (N_1670,In_92,In_517);
and U1671 (N_1671,In_485,In_224);
and U1672 (N_1672,In_26,In_295);
nor U1673 (N_1673,In_662,In_331);
nand U1674 (N_1674,In_690,In_349);
and U1675 (N_1675,In_378,In_403);
xnor U1676 (N_1676,In_711,In_455);
or U1677 (N_1677,In_451,In_897);
or U1678 (N_1678,In_331,In_63);
and U1679 (N_1679,In_643,In_935);
or U1680 (N_1680,In_286,In_363);
or U1681 (N_1681,In_892,In_494);
and U1682 (N_1682,In_71,In_983);
nor U1683 (N_1683,In_232,In_350);
nand U1684 (N_1684,In_9,In_49);
nand U1685 (N_1685,In_273,In_503);
nand U1686 (N_1686,In_978,In_945);
and U1687 (N_1687,In_2,In_302);
and U1688 (N_1688,In_760,In_453);
or U1689 (N_1689,In_858,In_854);
nor U1690 (N_1690,In_584,In_969);
and U1691 (N_1691,In_246,In_266);
and U1692 (N_1692,In_202,In_0);
or U1693 (N_1693,In_737,In_403);
xnor U1694 (N_1694,In_197,In_747);
nand U1695 (N_1695,In_460,In_499);
nor U1696 (N_1696,In_318,In_164);
or U1697 (N_1697,In_811,In_848);
or U1698 (N_1698,In_412,In_881);
or U1699 (N_1699,In_389,In_93);
nand U1700 (N_1700,In_743,In_424);
nand U1701 (N_1701,In_555,In_799);
nor U1702 (N_1702,In_103,In_137);
nand U1703 (N_1703,In_196,In_706);
nand U1704 (N_1704,In_545,In_922);
and U1705 (N_1705,In_706,In_653);
xor U1706 (N_1706,In_957,In_111);
or U1707 (N_1707,In_169,In_316);
nand U1708 (N_1708,In_65,In_104);
nand U1709 (N_1709,In_839,In_269);
and U1710 (N_1710,In_971,In_318);
and U1711 (N_1711,In_884,In_744);
and U1712 (N_1712,In_18,In_325);
and U1713 (N_1713,In_73,In_431);
nand U1714 (N_1714,In_210,In_780);
xor U1715 (N_1715,In_234,In_196);
nand U1716 (N_1716,In_688,In_787);
and U1717 (N_1717,In_515,In_174);
or U1718 (N_1718,In_911,In_197);
or U1719 (N_1719,In_125,In_745);
nor U1720 (N_1720,In_89,In_298);
nor U1721 (N_1721,In_515,In_213);
xor U1722 (N_1722,In_493,In_607);
nand U1723 (N_1723,In_580,In_677);
nor U1724 (N_1724,In_78,In_235);
nor U1725 (N_1725,In_679,In_117);
or U1726 (N_1726,In_166,In_15);
nand U1727 (N_1727,In_867,In_23);
nand U1728 (N_1728,In_571,In_18);
nand U1729 (N_1729,In_939,In_688);
and U1730 (N_1730,In_924,In_605);
or U1731 (N_1731,In_979,In_117);
or U1732 (N_1732,In_873,In_74);
and U1733 (N_1733,In_548,In_350);
nor U1734 (N_1734,In_494,In_877);
or U1735 (N_1735,In_935,In_427);
nor U1736 (N_1736,In_720,In_544);
and U1737 (N_1737,In_957,In_418);
or U1738 (N_1738,In_929,In_544);
nor U1739 (N_1739,In_487,In_191);
and U1740 (N_1740,In_687,In_91);
nor U1741 (N_1741,In_356,In_350);
nor U1742 (N_1742,In_872,In_590);
or U1743 (N_1743,In_650,In_765);
nor U1744 (N_1744,In_594,In_750);
or U1745 (N_1745,In_236,In_345);
and U1746 (N_1746,In_741,In_807);
and U1747 (N_1747,In_762,In_154);
nand U1748 (N_1748,In_178,In_5);
nor U1749 (N_1749,In_263,In_449);
or U1750 (N_1750,In_482,In_540);
or U1751 (N_1751,In_575,In_989);
or U1752 (N_1752,In_393,In_120);
or U1753 (N_1753,In_545,In_671);
nor U1754 (N_1754,In_141,In_555);
nor U1755 (N_1755,In_45,In_421);
nor U1756 (N_1756,In_437,In_670);
nor U1757 (N_1757,In_530,In_121);
nand U1758 (N_1758,In_684,In_976);
and U1759 (N_1759,In_921,In_625);
and U1760 (N_1760,In_0,In_298);
nand U1761 (N_1761,In_340,In_884);
nor U1762 (N_1762,In_9,In_130);
and U1763 (N_1763,In_941,In_672);
nor U1764 (N_1764,In_947,In_52);
or U1765 (N_1765,In_410,In_176);
nor U1766 (N_1766,In_10,In_172);
nand U1767 (N_1767,In_360,In_222);
and U1768 (N_1768,In_690,In_969);
and U1769 (N_1769,In_405,In_217);
nor U1770 (N_1770,In_657,In_946);
nand U1771 (N_1771,In_891,In_943);
or U1772 (N_1772,In_519,In_178);
and U1773 (N_1773,In_253,In_793);
and U1774 (N_1774,In_162,In_618);
or U1775 (N_1775,In_107,In_79);
nand U1776 (N_1776,In_400,In_120);
or U1777 (N_1777,In_462,In_470);
nor U1778 (N_1778,In_187,In_348);
nor U1779 (N_1779,In_405,In_678);
and U1780 (N_1780,In_652,In_94);
nor U1781 (N_1781,In_205,In_579);
or U1782 (N_1782,In_908,In_374);
and U1783 (N_1783,In_771,In_892);
nor U1784 (N_1784,In_807,In_507);
and U1785 (N_1785,In_804,In_381);
nand U1786 (N_1786,In_475,In_134);
nor U1787 (N_1787,In_53,In_989);
or U1788 (N_1788,In_603,In_508);
nor U1789 (N_1789,In_360,In_294);
nor U1790 (N_1790,In_650,In_659);
or U1791 (N_1791,In_742,In_883);
nor U1792 (N_1792,In_139,In_79);
or U1793 (N_1793,In_349,In_567);
nand U1794 (N_1794,In_909,In_822);
nand U1795 (N_1795,In_565,In_892);
and U1796 (N_1796,In_558,In_395);
nor U1797 (N_1797,In_487,In_795);
nor U1798 (N_1798,In_18,In_84);
or U1799 (N_1799,In_230,In_568);
nand U1800 (N_1800,In_451,In_687);
nand U1801 (N_1801,In_942,In_283);
and U1802 (N_1802,In_494,In_255);
and U1803 (N_1803,In_483,In_747);
nand U1804 (N_1804,In_812,In_958);
nand U1805 (N_1805,In_446,In_760);
nor U1806 (N_1806,In_986,In_68);
nand U1807 (N_1807,In_527,In_895);
and U1808 (N_1808,In_432,In_177);
or U1809 (N_1809,In_46,In_87);
nand U1810 (N_1810,In_406,In_783);
nand U1811 (N_1811,In_140,In_98);
or U1812 (N_1812,In_482,In_446);
or U1813 (N_1813,In_510,In_935);
and U1814 (N_1814,In_298,In_810);
or U1815 (N_1815,In_413,In_305);
and U1816 (N_1816,In_988,In_892);
nand U1817 (N_1817,In_747,In_675);
and U1818 (N_1818,In_523,In_474);
xnor U1819 (N_1819,In_425,In_555);
nand U1820 (N_1820,In_956,In_13);
or U1821 (N_1821,In_568,In_175);
nand U1822 (N_1822,In_935,In_236);
nand U1823 (N_1823,In_533,In_133);
nand U1824 (N_1824,In_860,In_988);
nor U1825 (N_1825,In_790,In_10);
nand U1826 (N_1826,In_985,In_906);
and U1827 (N_1827,In_848,In_903);
nor U1828 (N_1828,In_3,In_993);
and U1829 (N_1829,In_26,In_475);
nor U1830 (N_1830,In_29,In_884);
nor U1831 (N_1831,In_756,In_152);
nand U1832 (N_1832,In_450,In_74);
nor U1833 (N_1833,In_88,In_614);
nor U1834 (N_1834,In_558,In_426);
nor U1835 (N_1835,In_971,In_570);
and U1836 (N_1836,In_851,In_431);
nand U1837 (N_1837,In_13,In_496);
nand U1838 (N_1838,In_673,In_160);
or U1839 (N_1839,In_728,In_813);
nor U1840 (N_1840,In_944,In_125);
nor U1841 (N_1841,In_407,In_51);
or U1842 (N_1842,In_626,In_113);
or U1843 (N_1843,In_223,In_411);
or U1844 (N_1844,In_445,In_294);
or U1845 (N_1845,In_232,In_439);
nor U1846 (N_1846,In_410,In_618);
and U1847 (N_1847,In_296,In_824);
nor U1848 (N_1848,In_563,In_444);
nor U1849 (N_1849,In_418,In_309);
nor U1850 (N_1850,In_458,In_752);
or U1851 (N_1851,In_103,In_262);
nor U1852 (N_1852,In_894,In_701);
nor U1853 (N_1853,In_140,In_629);
and U1854 (N_1854,In_635,In_852);
nor U1855 (N_1855,In_722,In_46);
or U1856 (N_1856,In_105,In_709);
or U1857 (N_1857,In_590,In_252);
or U1858 (N_1858,In_436,In_593);
nand U1859 (N_1859,In_767,In_67);
and U1860 (N_1860,In_318,In_20);
and U1861 (N_1861,In_892,In_782);
nand U1862 (N_1862,In_865,In_900);
and U1863 (N_1863,In_579,In_145);
xnor U1864 (N_1864,In_121,In_763);
nor U1865 (N_1865,In_824,In_807);
nor U1866 (N_1866,In_109,In_628);
and U1867 (N_1867,In_867,In_88);
or U1868 (N_1868,In_180,In_378);
and U1869 (N_1869,In_9,In_134);
nor U1870 (N_1870,In_805,In_838);
nor U1871 (N_1871,In_307,In_385);
or U1872 (N_1872,In_776,In_505);
nor U1873 (N_1873,In_648,In_201);
and U1874 (N_1874,In_822,In_269);
or U1875 (N_1875,In_169,In_163);
nand U1876 (N_1876,In_640,In_149);
or U1877 (N_1877,In_669,In_125);
nor U1878 (N_1878,In_605,In_774);
nand U1879 (N_1879,In_348,In_415);
and U1880 (N_1880,In_720,In_527);
and U1881 (N_1881,In_67,In_521);
or U1882 (N_1882,In_276,In_332);
or U1883 (N_1883,In_397,In_41);
nand U1884 (N_1884,In_529,In_264);
or U1885 (N_1885,In_681,In_700);
and U1886 (N_1886,In_163,In_444);
and U1887 (N_1887,In_675,In_758);
and U1888 (N_1888,In_30,In_579);
or U1889 (N_1889,In_407,In_747);
nor U1890 (N_1890,In_499,In_321);
or U1891 (N_1891,In_944,In_410);
nor U1892 (N_1892,In_993,In_408);
nor U1893 (N_1893,In_561,In_602);
and U1894 (N_1894,In_17,In_725);
nand U1895 (N_1895,In_437,In_724);
or U1896 (N_1896,In_791,In_770);
nand U1897 (N_1897,In_158,In_833);
nand U1898 (N_1898,In_339,In_943);
and U1899 (N_1899,In_911,In_324);
nor U1900 (N_1900,In_864,In_535);
and U1901 (N_1901,In_101,In_559);
nor U1902 (N_1902,In_871,In_832);
nor U1903 (N_1903,In_189,In_140);
nor U1904 (N_1904,In_982,In_984);
and U1905 (N_1905,In_478,In_555);
nor U1906 (N_1906,In_435,In_881);
nor U1907 (N_1907,In_517,In_515);
xnor U1908 (N_1908,In_324,In_839);
nor U1909 (N_1909,In_189,In_570);
or U1910 (N_1910,In_994,In_560);
nor U1911 (N_1911,In_443,In_204);
nand U1912 (N_1912,In_679,In_369);
or U1913 (N_1913,In_423,In_560);
and U1914 (N_1914,In_792,In_483);
nand U1915 (N_1915,In_47,In_838);
or U1916 (N_1916,In_366,In_336);
and U1917 (N_1917,In_812,In_76);
and U1918 (N_1918,In_869,In_613);
or U1919 (N_1919,In_624,In_541);
nor U1920 (N_1920,In_429,In_5);
and U1921 (N_1921,In_150,In_279);
nor U1922 (N_1922,In_554,In_761);
or U1923 (N_1923,In_398,In_337);
nand U1924 (N_1924,In_351,In_748);
or U1925 (N_1925,In_105,In_857);
nor U1926 (N_1926,In_776,In_847);
nand U1927 (N_1927,In_505,In_502);
nand U1928 (N_1928,In_239,In_848);
and U1929 (N_1929,In_986,In_750);
or U1930 (N_1930,In_716,In_877);
and U1931 (N_1931,In_323,In_578);
or U1932 (N_1932,In_279,In_146);
or U1933 (N_1933,In_389,In_916);
nand U1934 (N_1934,In_24,In_96);
nor U1935 (N_1935,In_927,In_439);
and U1936 (N_1936,In_96,In_231);
nor U1937 (N_1937,In_342,In_767);
nand U1938 (N_1938,In_514,In_23);
nand U1939 (N_1939,In_462,In_333);
nor U1940 (N_1940,In_170,In_129);
or U1941 (N_1941,In_942,In_843);
and U1942 (N_1942,In_514,In_254);
nand U1943 (N_1943,In_798,In_330);
and U1944 (N_1944,In_878,In_533);
nand U1945 (N_1945,In_700,In_484);
and U1946 (N_1946,In_203,In_269);
nor U1947 (N_1947,In_591,In_976);
and U1948 (N_1948,In_955,In_318);
nor U1949 (N_1949,In_68,In_118);
nand U1950 (N_1950,In_755,In_428);
nand U1951 (N_1951,In_808,In_815);
or U1952 (N_1952,In_560,In_745);
nor U1953 (N_1953,In_570,In_646);
xnor U1954 (N_1954,In_252,In_303);
nor U1955 (N_1955,In_258,In_494);
nand U1956 (N_1956,In_988,In_697);
nor U1957 (N_1957,In_511,In_675);
nand U1958 (N_1958,In_430,In_489);
and U1959 (N_1959,In_26,In_900);
and U1960 (N_1960,In_271,In_520);
nor U1961 (N_1961,In_662,In_522);
nor U1962 (N_1962,In_513,In_862);
and U1963 (N_1963,In_411,In_937);
nor U1964 (N_1964,In_78,In_216);
nor U1965 (N_1965,In_473,In_802);
nand U1966 (N_1966,In_630,In_938);
and U1967 (N_1967,In_238,In_423);
nor U1968 (N_1968,In_54,In_332);
and U1969 (N_1969,In_252,In_568);
nor U1970 (N_1970,In_184,In_839);
nand U1971 (N_1971,In_47,In_9);
or U1972 (N_1972,In_38,In_181);
nor U1973 (N_1973,In_265,In_624);
or U1974 (N_1974,In_596,In_921);
nor U1975 (N_1975,In_6,In_709);
and U1976 (N_1976,In_394,In_729);
or U1977 (N_1977,In_329,In_122);
nand U1978 (N_1978,In_935,In_936);
nor U1979 (N_1979,In_941,In_656);
or U1980 (N_1980,In_66,In_431);
and U1981 (N_1981,In_962,In_0);
or U1982 (N_1982,In_979,In_521);
and U1983 (N_1983,In_947,In_103);
and U1984 (N_1984,In_588,In_271);
nor U1985 (N_1985,In_325,In_735);
and U1986 (N_1986,In_924,In_538);
and U1987 (N_1987,In_471,In_636);
or U1988 (N_1988,In_141,In_101);
nand U1989 (N_1989,In_79,In_227);
nor U1990 (N_1990,In_907,In_958);
nand U1991 (N_1991,In_388,In_349);
or U1992 (N_1992,In_415,In_22);
and U1993 (N_1993,In_522,In_960);
nand U1994 (N_1994,In_698,In_509);
and U1995 (N_1995,In_511,In_46);
and U1996 (N_1996,In_28,In_331);
or U1997 (N_1997,In_994,In_165);
or U1998 (N_1998,In_776,In_966);
nor U1999 (N_1999,In_803,In_515);
and U2000 (N_2000,N_522,N_1010);
and U2001 (N_2001,N_561,N_929);
nor U2002 (N_2002,N_1317,N_1568);
nor U2003 (N_2003,N_1822,N_1628);
nor U2004 (N_2004,N_1969,N_833);
nand U2005 (N_2005,N_219,N_50);
or U2006 (N_2006,N_1519,N_1300);
nor U2007 (N_2007,N_573,N_782);
and U2008 (N_2008,N_964,N_1600);
nor U2009 (N_2009,N_793,N_237);
nand U2010 (N_2010,N_1599,N_223);
nand U2011 (N_2011,N_424,N_334);
or U2012 (N_2012,N_416,N_1078);
and U2013 (N_2013,N_1182,N_1256);
and U2014 (N_2014,N_234,N_399);
nor U2015 (N_2015,N_1347,N_1412);
nand U2016 (N_2016,N_141,N_1803);
nor U2017 (N_2017,N_1198,N_972);
nor U2018 (N_2018,N_1899,N_1948);
or U2019 (N_2019,N_558,N_1479);
or U2020 (N_2020,N_643,N_1758);
nand U2021 (N_2021,N_1873,N_1745);
nand U2022 (N_2022,N_209,N_418);
and U2023 (N_2023,N_1666,N_878);
nand U2024 (N_2024,N_1016,N_825);
nor U2025 (N_2025,N_1001,N_42);
nand U2026 (N_2026,N_281,N_1856);
or U2027 (N_2027,N_195,N_1115);
nand U2028 (N_2028,N_730,N_282);
nor U2029 (N_2029,N_1794,N_846);
and U2030 (N_2030,N_1728,N_672);
nand U2031 (N_2031,N_1040,N_1447);
and U2032 (N_2032,N_284,N_227);
or U2033 (N_2033,N_1493,N_1104);
and U2034 (N_2034,N_688,N_707);
nand U2035 (N_2035,N_105,N_1153);
and U2036 (N_2036,N_1186,N_648);
or U2037 (N_2037,N_1397,N_395);
or U2038 (N_2038,N_687,N_104);
and U2039 (N_2039,N_1028,N_1158);
or U2040 (N_2040,N_1296,N_233);
nand U2041 (N_2041,N_1428,N_1625);
nand U2042 (N_2042,N_1357,N_852);
nor U2043 (N_2043,N_1420,N_1967);
or U2044 (N_2044,N_136,N_505);
or U2045 (N_2045,N_1301,N_254);
nor U2046 (N_2046,N_1272,N_1244);
and U2047 (N_2047,N_803,N_1175);
nand U2048 (N_2048,N_1473,N_1286);
nor U2049 (N_2049,N_269,N_1852);
nand U2050 (N_2050,N_723,N_287);
nor U2051 (N_2051,N_832,N_546);
or U2052 (N_2052,N_876,N_1498);
or U2053 (N_2053,N_1150,N_392);
nand U2054 (N_2054,N_1020,N_1726);
nand U2055 (N_2055,N_620,N_329);
and U2056 (N_2056,N_44,N_1680);
nor U2057 (N_2057,N_183,N_1553);
nor U2058 (N_2058,N_456,N_1570);
nor U2059 (N_2059,N_265,N_1316);
nor U2060 (N_2060,N_1635,N_952);
nand U2061 (N_2061,N_1349,N_693);
or U2062 (N_2062,N_677,N_544);
or U2063 (N_2063,N_1036,N_703);
or U2064 (N_2064,N_1389,N_719);
or U2065 (N_2065,N_1649,N_586);
and U2066 (N_2066,N_382,N_1499);
or U2067 (N_2067,N_1229,N_1114);
and U2068 (N_2068,N_201,N_1846);
and U2069 (N_2069,N_174,N_1631);
or U2070 (N_2070,N_1954,N_570);
nor U2071 (N_2071,N_829,N_1270);
nor U2072 (N_2072,N_20,N_1088);
nand U2073 (N_2073,N_1581,N_13);
nor U2074 (N_2074,N_1936,N_1064);
nor U2075 (N_2075,N_1667,N_486);
xor U2076 (N_2076,N_895,N_574);
nor U2077 (N_2077,N_1017,N_1613);
or U2078 (N_2078,N_1329,N_1864);
nor U2079 (N_2079,N_1754,N_1452);
nand U2080 (N_2080,N_1656,N_1056);
xor U2081 (N_2081,N_228,N_1964);
or U2082 (N_2082,N_515,N_649);
nand U2083 (N_2083,N_1273,N_795);
nor U2084 (N_2084,N_700,N_1509);
nor U2085 (N_2085,N_1465,N_1575);
nand U2086 (N_2086,N_1872,N_1627);
nor U2087 (N_2087,N_464,N_1266);
nor U2088 (N_2088,N_1384,N_423);
or U2089 (N_2089,N_1998,N_1468);
and U2090 (N_2090,N_1606,N_1097);
and U2091 (N_2091,N_1966,N_1436);
nand U2092 (N_2092,N_1845,N_651);
or U2093 (N_2093,N_1992,N_610);
nand U2094 (N_2094,N_1650,N_367);
nand U2095 (N_2095,N_1240,N_1083);
nor U2096 (N_2096,N_1518,N_1292);
and U2097 (N_2097,N_607,N_239);
or U2098 (N_2098,N_1454,N_684);
and U2099 (N_2099,N_405,N_1881);
nor U2100 (N_2100,N_583,N_1698);
nand U2101 (N_2101,N_1972,N_346);
nor U2102 (N_2102,N_1007,N_1193);
and U2103 (N_2103,N_998,N_1520);
and U2104 (N_2104,N_1477,N_664);
nor U2105 (N_2105,N_220,N_822);
xor U2106 (N_2106,N_824,N_1695);
nand U2107 (N_2107,N_954,N_580);
and U2108 (N_2108,N_200,N_1496);
nand U2109 (N_2109,N_937,N_1941);
and U2110 (N_2110,N_1180,N_814);
and U2111 (N_2111,N_1887,N_107);
nor U2112 (N_2112,N_283,N_1942);
nand U2113 (N_2113,N_407,N_735);
nand U2114 (N_2114,N_1179,N_1629);
nand U2115 (N_2115,N_1732,N_397);
nor U2116 (N_2116,N_1798,N_1209);
nor U2117 (N_2117,N_203,N_859);
nor U2118 (N_2118,N_1924,N_1602);
and U2119 (N_2119,N_461,N_617);
or U2120 (N_2120,N_1148,N_1206);
or U2121 (N_2121,N_1396,N_477);
nand U2122 (N_2122,N_678,N_1686);
or U2123 (N_2123,N_1101,N_1053);
and U2124 (N_2124,N_593,N_1343);
nor U2125 (N_2125,N_524,N_1279);
and U2126 (N_2126,N_1439,N_858);
nand U2127 (N_2127,N_670,N_1067);
and U2128 (N_2128,N_1879,N_1171);
nand U2129 (N_2129,N_1521,N_306);
or U2130 (N_2130,N_1713,N_1334);
and U2131 (N_2131,N_300,N_1855);
or U2132 (N_2132,N_1087,N_922);
and U2133 (N_2133,N_470,N_400);
nor U2134 (N_2134,N_1245,N_1000);
nand U2135 (N_2135,N_330,N_1424);
or U2136 (N_2136,N_404,N_1204);
and U2137 (N_2137,N_1061,N_62);
or U2138 (N_2138,N_1796,N_1931);
or U2139 (N_2139,N_1935,N_647);
and U2140 (N_2140,N_1988,N_32);
nand U2141 (N_2141,N_1912,N_1594);
or U2142 (N_2142,N_1634,N_1191);
or U2143 (N_2143,N_1073,N_454);
or U2144 (N_2144,N_1120,N_1251);
nor U2145 (N_2145,N_817,N_132);
or U2146 (N_2146,N_179,N_1095);
nand U2147 (N_2147,N_1320,N_96);
or U2148 (N_2148,N_1228,N_666);
and U2149 (N_2149,N_1643,N_799);
nand U2150 (N_2150,N_1042,N_1055);
nand U2151 (N_2151,N_1259,N_298);
and U2152 (N_2152,N_673,N_1973);
or U2153 (N_2153,N_857,N_913);
and U2154 (N_2154,N_836,N_997);
nor U2155 (N_2155,N_484,N_536);
and U2156 (N_2156,N_950,N_146);
or U2157 (N_2157,N_547,N_1504);
or U2158 (N_2158,N_1337,N_1841);
or U2159 (N_2159,N_542,N_1612);
nand U2160 (N_2160,N_1849,N_1395);
nand U2161 (N_2161,N_274,N_1417);
nor U2162 (N_2162,N_519,N_787);
nand U2163 (N_2163,N_376,N_1199);
and U2164 (N_2164,N_919,N_1348);
nand U2165 (N_2165,N_475,N_1837);
or U2166 (N_2166,N_609,N_907);
nor U2167 (N_2167,N_1587,N_71);
or U2168 (N_2168,N_981,N_77);
nor U2169 (N_2169,N_1003,N_927);
nand U2170 (N_2170,N_1891,N_1752);
nand U2171 (N_2171,N_206,N_1910);
nand U2172 (N_2172,N_1484,N_811);
and U2173 (N_2173,N_1611,N_1923);
nand U2174 (N_2174,N_956,N_35);
or U2175 (N_2175,N_1497,N_165);
nor U2176 (N_2176,N_1024,N_623);
nand U2177 (N_2177,N_439,N_601);
and U2178 (N_2178,N_226,N_1274);
and U2179 (N_2179,N_1840,N_285);
or U2180 (N_2180,N_675,N_493);
and U2181 (N_2181,N_756,N_1157);
nand U2182 (N_2182,N_1908,N_848);
nand U2183 (N_2183,N_68,N_1563);
or U2184 (N_2184,N_657,N_1748);
or U2185 (N_2185,N_821,N_626);
nor U2186 (N_2186,N_1930,N_387);
or U2187 (N_2187,N_358,N_1135);
or U2188 (N_2188,N_1419,N_313);
and U2189 (N_2189,N_152,N_1827);
nand U2190 (N_2190,N_885,N_340);
or U2191 (N_2191,N_1781,N_902);
nand U2192 (N_2192,N_1213,N_1647);
and U2193 (N_2193,N_1172,N_1838);
or U2194 (N_2194,N_1462,N_441);
nand U2195 (N_2195,N_1512,N_1543);
nand U2196 (N_2196,N_1940,N_886);
nand U2197 (N_2197,N_1770,N_1212);
and U2198 (N_2198,N_202,N_921);
or U2199 (N_2199,N_1381,N_745);
nor U2200 (N_2200,N_784,N_402);
nor U2201 (N_2201,N_541,N_1901);
or U2202 (N_2202,N_1922,N_1247);
or U2203 (N_2203,N_966,N_732);
nor U2204 (N_2204,N_936,N_1978);
and U2205 (N_2205,N_1729,N_1416);
nor U2206 (N_2206,N_1645,N_1608);
nor U2207 (N_2207,N_1778,N_1169);
nand U2208 (N_2208,N_1595,N_266);
or U2209 (N_2209,N_1684,N_496);
nor U2210 (N_2210,N_708,N_177);
nor U2211 (N_2211,N_1773,N_728);
and U2212 (N_2212,N_560,N_307);
nand U2213 (N_2213,N_1847,N_772);
and U2214 (N_2214,N_154,N_1878);
nand U2215 (N_2215,N_222,N_1641);
or U2216 (N_2216,N_299,N_1285);
xnor U2217 (N_2217,N_109,N_79);
or U2218 (N_2218,N_468,N_66);
nand U2219 (N_2219,N_1486,N_1832);
nor U2220 (N_2220,N_943,N_1690);
nand U2221 (N_2221,N_471,N_1775);
or U2222 (N_2222,N_24,N_888);
or U2223 (N_2223,N_1909,N_169);
nor U2224 (N_2224,N_1326,N_1839);
and U2225 (N_2225,N_1310,N_380);
or U2226 (N_2226,N_1687,N_633);
nand U2227 (N_2227,N_446,N_1124);
nor U2228 (N_2228,N_1203,N_479);
or U2229 (N_2229,N_1709,N_639);
or U2230 (N_2230,N_408,N_1038);
or U2231 (N_2231,N_1336,N_122);
or U2232 (N_2232,N_1471,N_1851);
and U2233 (N_2233,N_948,N_1724);
or U2234 (N_2234,N_842,N_1829);
and U2235 (N_2235,N_451,N_1380);
or U2236 (N_2236,N_590,N_738);
and U2237 (N_2237,N_1868,N_483);
and U2238 (N_2238,N_982,N_779);
nand U2239 (N_2239,N_995,N_1870);
and U2240 (N_2240,N_1346,N_1614);
nor U2241 (N_2241,N_1981,N_759);
nor U2242 (N_2242,N_820,N_722);
nor U2243 (N_2243,N_47,N_968);
nor U2244 (N_2244,N_1705,N_1844);
and U2245 (N_2245,N_1472,N_538);
and U2246 (N_2246,N_1507,N_1947);
nor U2247 (N_2247,N_1516,N_827);
xnor U2248 (N_2248,N_543,N_1305);
nand U2249 (N_2249,N_967,N_1975);
or U2250 (N_2250,N_1195,N_1815);
nor U2251 (N_2251,N_1315,N_1819);
nand U2252 (N_2252,N_379,N_767);
nand U2253 (N_2253,N_506,N_1534);
and U2254 (N_2254,N_11,N_1751);
nor U2255 (N_2255,N_1074,N_1820);
and U2256 (N_2256,N_54,N_473);
and U2257 (N_2257,N_260,N_602);
or U2258 (N_2258,N_1731,N_1955);
nor U2259 (N_2259,N_781,N_1574);
xor U2260 (N_2260,N_1707,N_83);
nor U2261 (N_2261,N_1181,N_1753);
and U2262 (N_2262,N_1077,N_157);
and U2263 (N_2263,N_1850,N_159);
nand U2264 (N_2264,N_1677,N_135);
nor U2265 (N_2265,N_689,N_305);
nor U2266 (N_2266,N_808,N_181);
and U2267 (N_2267,N_1584,N_1578);
nand U2268 (N_2268,N_1701,N_1685);
and U2269 (N_2269,N_115,N_765);
and U2270 (N_2270,N_1813,N_1413);
nor U2271 (N_2271,N_661,N_1692);
nand U2272 (N_2272,N_1159,N_1482);
nand U2273 (N_2273,N_1668,N_503);
xor U2274 (N_2274,N_1126,N_1694);
nand U2275 (N_2275,N_1399,N_45);
or U2276 (N_2276,N_1727,N_1354);
nor U2277 (N_2277,N_348,N_91);
nand U2278 (N_2278,N_501,N_749);
nand U2279 (N_2279,N_1322,N_1772);
or U2280 (N_2280,N_635,N_1716);
and U2281 (N_2281,N_775,N_143);
and U2282 (N_2282,N_51,N_216);
or U2283 (N_2283,N_1842,N_1934);
and U2284 (N_2284,N_628,N_869);
or U2285 (N_2285,N_1576,N_137);
nor U2286 (N_2286,N_448,N_1993);
or U2287 (N_2287,N_240,N_830);
nor U2288 (N_2288,N_1630,N_1363);
nor U2289 (N_2289,N_1019,N_1039);
or U2290 (N_2290,N_645,N_802);
nand U2291 (N_2291,N_1367,N_1928);
and U2292 (N_2292,N_1949,N_1387);
nor U2293 (N_2293,N_1639,N_447);
nand U2294 (N_2294,N_308,N_1052);
nand U2295 (N_2295,N_23,N_1081);
xnor U2296 (N_2296,N_410,N_78);
and U2297 (N_2297,N_839,N_1013);
and U2298 (N_2298,N_603,N_1757);
nor U2299 (N_2299,N_357,N_1792);
or U2300 (N_2300,N_1913,N_498);
or U2301 (N_2301,N_1513,N_1797);
nand U2302 (N_2302,N_1304,N_790);
nand U2303 (N_2303,N_1248,N_8);
nor U2304 (N_2304,N_1810,N_1289);
nand U2305 (N_2305,N_1253,N_1109);
and U2306 (N_2306,N_1071,N_315);
or U2307 (N_2307,N_1640,N_926);
or U2308 (N_2308,N_605,N_1489);
xnor U2309 (N_2309,N_816,N_419);
nor U2310 (N_2310,N_176,N_436);
and U2311 (N_2311,N_359,N_1123);
nor U2312 (N_2312,N_193,N_1886);
nor U2313 (N_2313,N_1092,N_1572);
or U2314 (N_2314,N_1549,N_1530);
nand U2315 (N_2315,N_396,N_840);
and U2316 (N_2316,N_375,N_740);
nor U2317 (N_2317,N_1332,N_1925);
nand U2318 (N_2318,N_750,N_806);
nand U2319 (N_2319,N_1173,N_931);
or U2320 (N_2320,N_123,N_253);
nand U2321 (N_2321,N_1569,N_559);
and U2322 (N_2322,N_7,N_642);
xor U2323 (N_2323,N_1485,N_1811);
or U2324 (N_2324,N_754,N_1165);
and U2325 (N_2325,N_1552,N_769);
nand U2326 (N_2326,N_1620,N_1108);
nand U2327 (N_2327,N_599,N_1638);
or U2328 (N_2328,N_705,N_249);
nand U2329 (N_2329,N_1113,N_482);
or U2330 (N_2330,N_1103,N_980);
nand U2331 (N_2331,N_1779,N_1721);
nand U2332 (N_2332,N_1571,N_1875);
nor U2333 (N_2333,N_747,N_1622);
or U2334 (N_2334,N_1566,N_6);
or U2335 (N_2335,N_1749,N_435);
and U2336 (N_2336,N_229,N_1529);
and U2337 (N_2337,N_81,N_894);
nand U2338 (N_2338,N_1808,N_1356);
and U2339 (N_2339,N_1062,N_398);
nor U2340 (N_2340,N_949,N_1335);
and U2341 (N_2341,N_514,N_1192);
nor U2342 (N_2342,N_1190,N_430);
nand U2343 (N_2343,N_99,N_494);
nor U2344 (N_2344,N_1795,N_1377);
xnor U2345 (N_2345,N_898,N_863);
nand U2346 (N_2346,N_472,N_679);
nand U2347 (N_2347,N_552,N_1980);
or U2348 (N_2348,N_213,N_1236);
nor U2349 (N_2349,N_1734,N_532);
or U2350 (N_2350,N_521,N_1756);
and U2351 (N_2351,N_1784,N_270);
or U2352 (N_2352,N_1926,N_131);
and U2353 (N_2353,N_403,N_916);
or U2354 (N_2354,N_1755,N_969);
and U2355 (N_2355,N_988,N_1110);
nor U2356 (N_2356,N_296,N_1596);
nor U2357 (N_2357,N_1111,N_1323);
or U2358 (N_2358,N_257,N_1425);
nand U2359 (N_2359,N_1807,N_1054);
nor U2360 (N_2360,N_890,N_1352);
or U2361 (N_2361,N_319,N_194);
nor U2362 (N_2362,N_95,N_530);
and U2363 (N_2363,N_1906,N_951);
or U2364 (N_2364,N_1715,N_1702);
nand U2365 (N_2365,N_40,N_1567);
nor U2366 (N_2366,N_721,N_1768);
and U2367 (N_2367,N_1565,N_211);
nand U2368 (N_2368,N_67,N_1505);
or U2369 (N_2369,N_1510,N_34);
nor U2370 (N_2370,N_720,N_406);
and U2371 (N_2371,N_581,N_1537);
nor U2372 (N_2372,N_867,N_545);
or U2373 (N_2373,N_1221,N_291);
and U2374 (N_2374,N_1459,N_17);
nor U2375 (N_2375,N_520,N_164);
nor U2376 (N_2376,N_2,N_490);
nand U2377 (N_2377,N_785,N_903);
and U2378 (N_2378,N_261,N_332);
and U2379 (N_2379,N_1362,N_333);
and U2380 (N_2380,N_467,N_854);
or U2381 (N_2381,N_338,N_844);
nor U2382 (N_2382,N_190,N_1122);
and U2383 (N_2383,N_1069,N_641);
nor U2384 (N_2384,N_1278,N_422);
nor U2385 (N_2385,N_459,N_810);
nor U2386 (N_2386,N_1682,N_163);
or U2387 (N_2387,N_1466,N_25);
nand U2388 (N_2388,N_1393,N_1943);
nand U2389 (N_2389,N_1607,N_1116);
nor U2390 (N_2390,N_27,N_1205);
nor U2391 (N_2391,N_771,N_1491);
nand U2392 (N_2392,N_1711,N_1670);
nand U2393 (N_2393,N_908,N_861);
nand U2394 (N_2394,N_1080,N_449);
or U2395 (N_2395,N_4,N_813);
nor U2396 (N_2396,N_336,N_1207);
nor U2397 (N_2397,N_1786,N_584);
nor U2398 (N_2398,N_262,N_741);
nand U2399 (N_2399,N_1874,N_1823);
or U2400 (N_2400,N_826,N_1591);
nand U2401 (N_2401,N_372,N_812);
and U2402 (N_2402,N_149,N_188);
and U2403 (N_2403,N_355,N_650);
nor U2404 (N_2404,N_696,N_102);
nor U2405 (N_2405,N_21,N_884);
xnor U2406 (N_2406,N_562,N_389);
xor U2407 (N_2407,N_204,N_1719);
nand U2408 (N_2408,N_1012,N_555);
or U2409 (N_2409,N_170,N_453);
and U2410 (N_2410,N_232,N_1117);
nor U2411 (N_2411,N_1456,N_381);
or U2412 (N_2412,N_1896,N_1324);
and U2413 (N_2413,N_1252,N_1968);
or U2414 (N_2414,N_932,N_130);
and U2415 (N_2415,N_61,N_934);
nand U2416 (N_2416,N_1771,N_101);
nor U2417 (N_2417,N_1100,N_278);
nor U2418 (N_2418,N_729,N_1603);
or U2419 (N_2419,N_1072,N_1438);
or U2420 (N_2420,N_1446,N_1583);
and U2421 (N_2421,N_1284,N_1956);
nand U2422 (N_2422,N_1342,N_1293);
nand U2423 (N_2423,N_1234,N_778);
nor U2424 (N_2424,N_915,N_856);
or U2425 (N_2425,N_991,N_866);
and U2426 (N_2426,N_377,N_1133);
nor U2427 (N_2427,N_1714,N_985);
and U2428 (N_2428,N_710,N_798);
nand U2429 (N_2429,N_725,N_1525);
nand U2430 (N_2430,N_928,N_535);
or U2431 (N_2431,N_365,N_1235);
nand U2432 (N_2432,N_1201,N_84);
or U2433 (N_2433,N_69,N_853);
or U2434 (N_2434,N_704,N_629);
nor U2435 (N_2435,N_1535,N_1360);
nand U2436 (N_2436,N_1366,N_258);
and U2437 (N_2437,N_1619,N_302);
and U2438 (N_2438,N_1994,N_205);
nand U2439 (N_2439,N_489,N_1657);
or U2440 (N_2440,N_187,N_342);
or U2441 (N_2441,N_1254,N_1589);
and U2442 (N_2442,N_1933,N_1556);
nand U2443 (N_2443,N_1880,N_556);
nor U2444 (N_2444,N_356,N_273);
or U2445 (N_2445,N_1524,N_763);
or U2446 (N_2446,N_1962,N_843);
nor U2447 (N_2447,N_1021,N_871);
nand U2448 (N_2448,N_549,N_1060);
and U2449 (N_2449,N_1105,N_1761);
and U2450 (N_2450,N_1050,N_774);
nand U2451 (N_2451,N_1089,N_1210);
or U2452 (N_2452,N_636,N_576);
nor U2453 (N_2453,N_469,N_529);
nor U2454 (N_2454,N_151,N_807);
and U2455 (N_2455,N_1762,N_1742);
and U2456 (N_2456,N_1735,N_1929);
nand U2457 (N_2457,N_1979,N_1548);
and U2458 (N_2458,N_1090,N_1411);
nand U2459 (N_2459,N_663,N_1573);
and U2460 (N_2460,N_5,N_668);
nand U2461 (N_2461,N_1358,N_1805);
nor U2462 (N_2462,N_697,N_1211);
nor U2463 (N_2463,N_10,N_414);
nor U2464 (N_2464,N_1665,N_488);
nor U2465 (N_2465,N_1562,N_1951);
and U2466 (N_2466,N_975,N_1299);
or U2467 (N_2467,N_1268,N_480);
xor U2468 (N_2468,N_75,N_445);
or U2469 (N_2469,N_1066,N_1269);
and U2470 (N_2470,N_371,N_1545);
nand U2471 (N_2471,N_322,N_1453);
xnor U2472 (N_2472,N_39,N_1281);
and U2473 (N_2473,N_337,N_933);
or U2474 (N_2474,N_1131,N_714);
or U2475 (N_2475,N_343,N_724);
nor U2476 (N_2476,N_706,N_587);
nand U2477 (N_2477,N_133,N_1672);
nor U2478 (N_2478,N_199,N_637);
nor U2479 (N_2479,N_1134,N_823);
and U2480 (N_2480,N_912,N_373);
and U2481 (N_2481,N_1463,N_318);
or U2482 (N_2482,N_1338,N_996);
nand U2483 (N_2483,N_776,N_533);
or U2484 (N_2484,N_321,N_1263);
or U2485 (N_2485,N_1290,N_1750);
or U2486 (N_2486,N_1894,N_386);
nand U2487 (N_2487,N_1693,N_1196);
nor U2488 (N_2488,N_1809,N_1409);
or U2489 (N_2489,N_457,N_1231);
and U2490 (N_2490,N_1659,N_1238);
and U2491 (N_2491,N_660,N_1508);
and U2492 (N_2492,N_1740,N_1517);
nor U2493 (N_2493,N_275,N_1458);
nand U2494 (N_2494,N_1154,N_748);
and U2495 (N_2495,N_654,N_691);
nor U2496 (N_2496,N_1185,N_1262);
nand U2497 (N_2497,N_1370,N_1882);
nor U2498 (N_2498,N_1433,N_320);
or U2499 (N_2499,N_680,N_147);
nor U2500 (N_2500,N_214,N_1006);
nand U2501 (N_2501,N_1788,N_572);
nand U2502 (N_2502,N_1558,N_106);
nor U2503 (N_2503,N_914,N_986);
nor U2504 (N_2504,N_841,N_736);
nor U2505 (N_2505,N_1350,N_652);
and U2506 (N_2506,N_160,N_786);
nor U2507 (N_2507,N_1557,N_98);
nor U2508 (N_2508,N_597,N_344);
or U2509 (N_2509,N_1156,N_874);
or U2510 (N_2510,N_1364,N_1893);
and U2511 (N_2511,N_29,N_990);
or U2512 (N_2512,N_1739,N_1586);
nor U2513 (N_2513,N_1369,N_74);
xor U2514 (N_2514,N_301,N_280);
and U2515 (N_2515,N_481,N_1085);
and U2516 (N_2516,N_849,N_244);
nand U2517 (N_2517,N_977,N_1722);
xor U2518 (N_2518,N_1623,N_292);
nor U2519 (N_2519,N_658,N_930);
nor U2520 (N_2520,N_19,N_800);
nand U2521 (N_2521,N_412,N_429);
or U2522 (N_2522,N_1946,N_1533);
nor U2523 (N_2523,N_1442,N_1903);
and U2524 (N_2524,N_310,N_1265);
nand U2525 (N_2525,N_1125,N_1730);
nand U2526 (N_2526,N_766,N_312);
xor U2527 (N_2527,N_1976,N_1325);
nand U2528 (N_2528,N_111,N_1303);
or U2529 (N_2529,N_1560,N_1610);
nand U2530 (N_2530,N_293,N_113);
and U2531 (N_2531,N_575,N_1624);
and U2532 (N_2532,N_1637,N_247);
nand U2533 (N_2533,N_994,N_1282);
nand U2534 (N_2534,N_279,N_1676);
and U2535 (N_2535,N_1239,N_1511);
or U2536 (N_2536,N_374,N_773);
or U2537 (N_2537,N_1255,N_1218);
and U2538 (N_2538,N_460,N_116);
and U2539 (N_2539,N_794,N_1200);
or U2540 (N_2540,N_1653,N_182);
nor U2541 (N_2541,N_923,N_1541);
and U2542 (N_2542,N_819,N_1174);
nand U2543 (N_2543,N_804,N_837);
nor U2544 (N_2544,N_550,N_432);
or U2545 (N_2545,N_121,N_134);
nor U2546 (N_2546,N_618,N_744);
and U2547 (N_2547,N_277,N_1374);
and U2548 (N_2548,N_420,N_1233);
nor U2549 (N_2549,N_1791,N_578);
nand U2550 (N_2550,N_604,N_1461);
or U2551 (N_2551,N_1522,N_57);
and U2552 (N_2552,N_655,N_1242);
and U2553 (N_2553,N_1155,N_1961);
or U2554 (N_2554,N_491,N_289);
and U2555 (N_2555,N_142,N_1971);
xnor U2556 (N_2556,N_526,N_119);
nand U2557 (N_2557,N_370,N_674);
nand U2558 (N_2558,N_797,N_198);
or U2559 (N_2559,N_1331,N_476);
nor U2560 (N_2560,N_1059,N_192);
nand U2561 (N_2561,N_15,N_1488);
and U2562 (N_2562,N_1857,N_60);
nor U2563 (N_2563,N_1214,N_695);
or U2564 (N_2564,N_564,N_1536);
or U2565 (N_2565,N_128,N_125);
xnor U2566 (N_2566,N_897,N_1076);
or U2567 (N_2567,N_155,N_1002);
nor U2568 (N_2568,N_516,N_1223);
nor U2569 (N_2569,N_751,N_1464);
and U2570 (N_2570,N_591,N_1889);
nor U2571 (N_2571,N_1683,N_973);
or U2572 (N_2572,N_939,N_1814);
and U2573 (N_2573,N_443,N_1490);
or U2574 (N_2574,N_1478,N_1696);
nand U2575 (N_2575,N_1662,N_1306);
nand U2576 (N_2576,N_510,N_1152);
nor U2577 (N_2577,N_1361,N_828);
and U2578 (N_2578,N_770,N_1093);
nand U2579 (N_2579,N_1267,N_504);
and U2580 (N_2580,N_56,N_883);
nand U2581 (N_2581,N_1700,N_1999);
xor U2582 (N_2582,N_369,N_139);
nand U2583 (N_2583,N_1098,N_701);
and U2584 (N_2584,N_539,N_53);
or U2585 (N_2585,N_690,N_1869);
or U2586 (N_2586,N_621,N_1022);
nor U2587 (N_2587,N_1294,N_1806);
nor U2588 (N_2588,N_245,N_920);
or U2589 (N_2589,N_1450,N_1183);
nor U2590 (N_2590,N_1767,N_945);
nor U2591 (N_2591,N_1802,N_613);
nand U2592 (N_2592,N_345,N_1658);
xor U2593 (N_2593,N_1044,N_1960);
nor U2594 (N_2594,N_1445,N_120);
nor U2595 (N_2595,N_172,N_1648);
nand U2596 (N_2596,N_924,N_567);
or U2597 (N_2597,N_537,N_248);
nand U2598 (N_2598,N_585,N_1070);
nand U2599 (N_2599,N_983,N_1532);
or U2600 (N_2600,N_1547,N_1031);
or U2601 (N_2601,N_1011,N_1515);
and U2602 (N_2602,N_1318,N_1219);
nor U2603 (N_2603,N_1633,N_733);
or U2604 (N_2604,N_1144,N_1664);
or U2605 (N_2605,N_1481,N_1388);
or U2606 (N_2606,N_791,N_215);
and U2607 (N_2607,N_297,N_1644);
nand U2608 (N_2608,N_1222,N_440);
and U2609 (N_2609,N_126,N_1243);
and U2610 (N_2610,N_350,N_1215);
nor U2611 (N_2611,N_1905,N_1220);
and U2612 (N_2612,N_1585,N_1743);
and U2613 (N_2613,N_612,N_394);
or U2614 (N_2614,N_792,N_509);
or U2615 (N_2615,N_566,N_1249);
and U2616 (N_2616,N_124,N_1136);
and U2617 (N_2617,N_415,N_1333);
nor U2618 (N_2618,N_1793,N_1014);
nor U2619 (N_2619,N_433,N_1291);
nand U2620 (N_2620,N_1400,N_1843);
or U2621 (N_2621,N_1883,N_731);
nor U2622 (N_2622,N_117,N_1476);
or U2623 (N_2623,N_127,N_1043);
nor U2624 (N_2624,N_150,N_317);
or U2625 (N_2625,N_780,N_1495);
nand U2626 (N_2626,N_1260,N_1440);
nor U2627 (N_2627,N_1871,N_528);
or U2628 (N_2628,N_757,N_255);
or U2629 (N_2629,N_746,N_1443);
or U2630 (N_2630,N_1577,N_1385);
and U2631 (N_2631,N_881,N_557);
nor U2632 (N_2632,N_1738,N_1455);
and U2633 (N_2633,N_1818,N_1588);
nand U2634 (N_2634,N_1593,N_1965);
or U2635 (N_2635,N_761,N_1984);
or U2636 (N_2636,N_1084,N_1160);
nand U2637 (N_2637,N_963,N_1187);
xor U2638 (N_2638,N_1378,N_1386);
and U2639 (N_2639,N_1121,N_1651);
nor U2640 (N_2640,N_1783,N_891);
or U2641 (N_2641,N_1995,N_1669);
and U2642 (N_2642,N_709,N_999);
nand U2643 (N_2643,N_563,N_845);
nand U2644 (N_2644,N_1164,N_940);
nand U2645 (N_2645,N_877,N_702);
nor U2646 (N_2646,N_427,N_1327);
nor U2647 (N_2647,N_1405,N_1957);
nand U2648 (N_2648,N_1918,N_667);
nand U2649 (N_2649,N_892,N_391);
and U2650 (N_2650,N_1137,N_1733);
nor U2651 (N_2651,N_156,N_1319);
nand U2652 (N_2652,N_743,N_90);
nor U2653 (N_2653,N_264,N_421);
nand U2654 (N_2654,N_1202,N_683);
and U2655 (N_2655,N_1661,N_1932);
nor U2656 (N_2656,N_1427,N_108);
nor U2657 (N_2657,N_1224,N_873);
and U2658 (N_2658,N_1765,N_1704);
nor U2659 (N_2659,N_855,N_1769);
and U2660 (N_2660,N_531,N_1710);
nor U2661 (N_2661,N_1514,N_686);
nand U2662 (N_2662,N_384,N_1283);
and U2663 (N_2663,N_1825,N_38);
nor U2664 (N_2664,N_272,N_1652);
or U2665 (N_2665,N_1119,N_947);
nor U2666 (N_2666,N_1106,N_1776);
or U2667 (N_2667,N_455,N_85);
and U2668 (N_2668,N_271,N_989);
nor U2669 (N_2669,N_987,N_1139);
and U2670 (N_2670,N_970,N_1474);
and U2671 (N_2671,N_218,N_1703);
or U2672 (N_2672,N_627,N_1208);
xnor U2673 (N_2673,N_167,N_777);
or U2674 (N_2674,N_946,N_882);
and U2675 (N_2675,N_250,N_716);
or U2676 (N_2676,N_1777,N_1312);
nor U2677 (N_2677,N_1920,N_1018);
or U2678 (N_2678,N_1888,N_1604);
or U2679 (N_2679,N_175,N_1986);
and U2680 (N_2680,N_335,N_1163);
xnor U2681 (N_2681,N_1816,N_1673);
or U2682 (N_2682,N_252,N_669);
or U2683 (N_2683,N_1937,N_1339);
nand U2684 (N_2684,N_401,N_487);
and U2685 (N_2685,N_1441,N_1344);
or U2686 (N_2686,N_1678,N_1787);
or U2687 (N_2687,N_717,N_1764);
and U2688 (N_2688,N_86,N_815);
xnor U2689 (N_2689,N_1741,N_1225);
xor U2690 (N_2690,N_1009,N_1712);
nor U2691 (N_2691,N_646,N_1161);
nand U2692 (N_2692,N_63,N_378);
or U2693 (N_2693,N_268,N_862);
nor U2694 (N_2694,N_1746,N_632);
and U2695 (N_2695,N_1835,N_1782);
and U2696 (N_2696,N_362,N_755);
and U2697 (N_2697,N_1034,N_178);
and U2698 (N_2698,N_1130,N_1004);
or U2699 (N_2699,N_595,N_737);
nand U2700 (N_2700,N_889,N_1128);
nor U2701 (N_2701,N_1708,N_1720);
nor U2702 (N_2702,N_1884,N_1298);
or U2703 (N_2703,N_1029,N_0);
and U2704 (N_2704,N_1538,N_474);
or U2705 (N_2705,N_551,N_52);
and U2706 (N_2706,N_1916,N_805);
nor U2707 (N_2707,N_437,N_630);
nand U2708 (N_2708,N_1426,N_1030);
xnor U2709 (N_2709,N_1328,N_640);
and U2710 (N_2710,N_571,N_1390);
or U2711 (N_2711,N_1048,N_1939);
nor U2712 (N_2712,N_1531,N_185);
and U2713 (N_2713,N_1876,N_1280);
nor U2714 (N_2714,N_681,N_1636);
and U2715 (N_2715,N_1178,N_80);
nand U2716 (N_2716,N_354,N_1475);
and U2717 (N_2717,N_1434,N_752);
nand U2718 (N_2718,N_1848,N_1615);
nand U2719 (N_2719,N_512,N_511);
nand U2720 (N_2720,N_1457,N_393);
nand U2721 (N_2721,N_1470,N_565);
nand U2722 (N_2722,N_88,N_339);
nand U2723 (N_2723,N_1094,N_622);
nor U2724 (N_2724,N_1983,N_267);
nor U2725 (N_2725,N_148,N_835);
and U2726 (N_2726,N_1421,N_1129);
and U2727 (N_2727,N_1141,N_962);
nand U2728 (N_2728,N_1096,N_1373);
xor U2729 (N_2729,N_758,N_1170);
or U2730 (N_2730,N_100,N_1246);
and U2731 (N_2731,N_788,N_1271);
and U2732 (N_2732,N_1597,N_1145);
and U2733 (N_2733,N_1675,N_413);
or U2734 (N_2734,N_955,N_495);
nor U2735 (N_2735,N_715,N_251);
xnor U2736 (N_2736,N_1854,N_917);
nand U2737 (N_2737,N_1311,N_1448);
nor U2738 (N_2738,N_850,N_1877);
and U2739 (N_2739,N_168,N_1166);
nand U2740 (N_2740,N_1744,N_899);
xnor U2741 (N_2741,N_93,N_608);
nor U2742 (N_2742,N_140,N_290);
and U2743 (N_2743,N_1,N_783);
nor U2744 (N_2744,N_309,N_331);
and U2745 (N_2745,N_1919,N_55);
or U2746 (N_2746,N_974,N_1826);
or U2747 (N_2747,N_230,N_1528);
and U2748 (N_2748,N_644,N_1550);
nand U2749 (N_2749,N_235,N_1341);
or U2750 (N_2750,N_409,N_692);
and U2751 (N_2751,N_525,N_295);
and U2752 (N_2752,N_1789,N_1330);
or U2753 (N_2753,N_712,N_1379);
or U2754 (N_2754,N_796,N_31);
nand U2755 (N_2755,N_1671,N_1904);
nor U2756 (N_2756,N_993,N_97);
xnor U2757 (N_2757,N_1184,N_941);
nand U2758 (N_2758,N_1642,N_1351);
xnor U2759 (N_2759,N_1063,N_698);
and U2760 (N_2760,N_1898,N_341);
or U2761 (N_2761,N_1483,N_129);
and U2762 (N_2762,N_492,N_327);
nand U2763 (N_2763,N_611,N_1345);
and U2764 (N_2764,N_1970,N_513);
and U2765 (N_2765,N_221,N_600);
nand U2766 (N_2766,N_485,N_789);
nor U2767 (N_2767,N_1102,N_764);
nand U2768 (N_2768,N_1035,N_450);
nor U2769 (N_2769,N_1944,N_1655);
nor U2770 (N_2770,N_1435,N_1314);
or U2771 (N_2771,N_880,N_1812);
or U2772 (N_2772,N_1057,N_1288);
and U2773 (N_2773,N_1853,N_212);
nand U2774 (N_2774,N_659,N_1355);
nand U2775 (N_2775,N_1147,N_64);
and U2776 (N_2776,N_1277,N_1974);
xnor U2777 (N_2777,N_893,N_1307);
and U2778 (N_2778,N_363,N_1799);
nor U2779 (N_2779,N_1406,N_82);
and U2780 (N_2780,N_1834,N_1414);
nand U2781 (N_2781,N_887,N_360);
nand U2782 (N_2782,N_1551,N_314);
and U2783 (N_2783,N_65,N_166);
and U2784 (N_2784,N_753,N_1836);
or U2785 (N_2785,N_103,N_1688);
nor U2786 (N_2786,N_1747,N_992);
and U2787 (N_2787,N_1691,N_1359);
and U2788 (N_2788,N_554,N_1917);
and U2789 (N_2789,N_1865,N_161);
and U2790 (N_2790,N_1099,N_1674);
nor U2791 (N_2791,N_1449,N_818);
and U2792 (N_2792,N_1501,N_231);
and U2793 (N_2793,N_462,N_1991);
nor U2794 (N_2794,N_383,N_1774);
or U2795 (N_2795,N_699,N_1365);
and U2796 (N_2796,N_1950,N_1860);
nor U2797 (N_2797,N_548,N_534);
or U2798 (N_2798,N_1005,N_870);
nand U2799 (N_2799,N_1506,N_909);
and U2800 (N_2800,N_711,N_1392);
and U2801 (N_2801,N_323,N_1008);
nor U2802 (N_2802,N_41,N_1142);
and U2803 (N_2803,N_1663,N_259);
or U2804 (N_2804,N_1621,N_1086);
nor U2805 (N_2805,N_263,N_1216);
or U2806 (N_2806,N_760,N_1276);
or U2807 (N_2807,N_1194,N_1025);
or U2808 (N_2808,N_1544,N_1915);
or U2809 (N_2809,N_1540,N_1927);
and U2810 (N_2810,N_294,N_1555);
nand U2811 (N_2811,N_118,N_1759);
nor U2812 (N_2812,N_351,N_1188);
nor U2813 (N_2813,N_1467,N_1403);
nor U2814 (N_2814,N_1885,N_1127);
and U2815 (N_2815,N_682,N_326);
or U2816 (N_2816,N_1480,N_153);
or U2817 (N_2817,N_22,N_1717);
xor U2818 (N_2818,N_868,N_1353);
nor U2819 (N_2819,N_971,N_1911);
and U2820 (N_2820,N_1261,N_1554);
nor U2821 (N_2821,N_502,N_1725);
nor U2822 (N_2822,N_1391,N_463);
nand U2823 (N_2823,N_353,N_18);
nand U2824 (N_2824,N_596,N_59);
or U2825 (N_2825,N_1902,N_1831);
nor U2826 (N_2826,N_246,N_1895);
and U2827 (N_2827,N_851,N_1859);
nor U2828 (N_2828,N_1697,N_1217);
nor U2829 (N_2829,N_979,N_624);
and U2830 (N_2830,N_1033,N_217);
nand U2831 (N_2831,N_582,N_910);
nor U2832 (N_2832,N_112,N_197);
nand U2833 (N_2833,N_1699,N_466);
nand U2834 (N_2834,N_568,N_452);
or U2835 (N_2835,N_1582,N_1681);
nor U2836 (N_2836,N_37,N_70);
nor U2837 (N_2837,N_304,N_28);
and U2838 (N_2838,N_1821,N_1500);
nor U2839 (N_2839,N_1065,N_58);
and U2840 (N_2840,N_1410,N_1945);
and U2841 (N_2841,N_92,N_236);
and U2842 (N_2842,N_1907,N_834);
and U2843 (N_2843,N_1494,N_965);
nor U2844 (N_2844,N_1398,N_207);
or U2845 (N_2845,N_1046,N_1437);
or U2846 (N_2846,N_417,N_653);
or U2847 (N_2847,N_114,N_1914);
or U2848 (N_2848,N_1646,N_1723);
xor U2849 (N_2849,N_243,N_1023);
nor U2850 (N_2850,N_1977,N_631);
and U2851 (N_2851,N_30,N_1626);
and U2852 (N_2852,N_171,N_1997);
nand U2853 (N_2853,N_48,N_1250);
or U2854 (N_2854,N_26,N_1866);
nor U2855 (N_2855,N_676,N_347);
and U2856 (N_2856,N_935,N_1737);
xnor U2857 (N_2857,N_1780,N_76);
or U2858 (N_2858,N_1503,N_1230);
or U2859 (N_2859,N_1407,N_1817);
or U2860 (N_2860,N_1601,N_36);
nor U2861 (N_2861,N_276,N_1592);
and U2862 (N_2862,N_896,N_1858);
nand U2863 (N_2863,N_523,N_458);
nand U2864 (N_2864,N_1963,N_1580);
nor U2865 (N_2865,N_606,N_1985);
nor U2866 (N_2866,N_1897,N_598);
nand U2867 (N_2867,N_368,N_1689);
nor U2868 (N_2868,N_1590,N_1718);
nand U2869 (N_2869,N_1041,N_1958);
or U2870 (N_2870,N_656,N_49);
nand U2871 (N_2871,N_875,N_210);
and U2872 (N_2872,N_1579,N_1295);
or U2873 (N_2873,N_1058,N_958);
or U2874 (N_2874,N_517,N_904);
nand U2875 (N_2875,N_1830,N_1189);
or U2876 (N_2876,N_1408,N_390);
xnor U2877 (N_2877,N_1460,N_1237);
nand U2878 (N_2878,N_901,N_1952);
and U2879 (N_2879,N_225,N_589);
nor U2880 (N_2880,N_1368,N_1151);
or U2881 (N_2881,N_1953,N_518);
and U2882 (N_2882,N_1900,N_1559);
or U2883 (N_2883,N_1546,N_508);
nor U2884 (N_2884,N_1143,N_425);
nand U2885 (N_2885,N_1313,N_1785);
nor U2886 (N_2886,N_1132,N_918);
and U2887 (N_2887,N_1989,N_1800);
nand U2888 (N_2888,N_72,N_241);
nor U2889 (N_2889,N_43,N_553);
nor U2890 (N_2890,N_864,N_1679);
nand U2891 (N_2891,N_1258,N_242);
nand U2892 (N_2892,N_1469,N_162);
and U2893 (N_2893,N_957,N_625);
nand U2894 (N_2894,N_911,N_1015);
or U2895 (N_2895,N_594,N_1492);
nor U2896 (N_2896,N_619,N_1618);
and U2897 (N_2897,N_1138,N_1079);
nand U2898 (N_2898,N_1890,N_426);
nand U2899 (N_2899,N_442,N_1632);
nor U2900 (N_2900,N_577,N_1340);
and U2901 (N_2901,N_1140,N_110);
nor U2902 (N_2902,N_1921,N_1422);
nor U2903 (N_2903,N_762,N_73);
xor U2904 (N_2904,N_1047,N_809);
or U2905 (N_2905,N_1394,N_1564);
or U2906 (N_2906,N_1027,N_1862);
nor U2907 (N_2907,N_1026,N_1068);
and U2908 (N_2908,N_14,N_592);
xor U2909 (N_2909,N_1539,N_286);
and U2910 (N_2910,N_1371,N_1107);
nor U2911 (N_2911,N_1241,N_1146);
or U2912 (N_2912,N_1616,N_1444);
nor U2913 (N_2913,N_1418,N_1082);
xor U2914 (N_2914,N_801,N_434);
and U2915 (N_2915,N_311,N_665);
nor U2916 (N_2916,N_94,N_444);
and U2917 (N_2917,N_616,N_1197);
and U2918 (N_2918,N_173,N_1760);
nor U2919 (N_2919,N_847,N_288);
or U2920 (N_2920,N_860,N_1861);
or U2921 (N_2921,N_1987,N_1938);
and U2922 (N_2922,N_364,N_1432);
nor U2923 (N_2923,N_540,N_944);
and U2924 (N_2924,N_385,N_1598);
or U2925 (N_2925,N_879,N_184);
nor U2926 (N_2926,N_1302,N_1415);
and U2927 (N_2927,N_1561,N_1232);
nor U2928 (N_2928,N_734,N_615);
and U2929 (N_2929,N_1487,N_1959);
or U2930 (N_2930,N_726,N_138);
or U2931 (N_2931,N_1431,N_497);
and U2932 (N_2932,N_1402,N_1112);
and U2933 (N_2933,N_1051,N_1264);
and U2934 (N_2934,N_191,N_180);
and U2935 (N_2935,N_1526,N_1892);
or U2936 (N_2936,N_1654,N_960);
nor U2937 (N_2937,N_1660,N_189);
nand U2938 (N_2938,N_186,N_1168);
nor U2939 (N_2939,N_1297,N_12);
nand U2940 (N_2940,N_1275,N_1451);
nand U2941 (N_2941,N_1801,N_1226);
and U2942 (N_2942,N_1118,N_349);
or U2943 (N_2943,N_1401,N_961);
and U2944 (N_2944,N_1736,N_1804);
nor U2945 (N_2945,N_1982,N_1766);
nand U2946 (N_2946,N_316,N_588);
or U2947 (N_2947,N_499,N_1091);
and U2948 (N_2948,N_1617,N_838);
or U2949 (N_2949,N_1372,N_634);
nand U2950 (N_2950,N_1828,N_388);
or U2951 (N_2951,N_1383,N_1833);
or U2952 (N_2952,N_1149,N_33);
and U2953 (N_2953,N_1605,N_361);
nor U2954 (N_2954,N_1075,N_900);
nor U2955 (N_2955,N_145,N_89);
or U2956 (N_2956,N_1706,N_1037);
or U2957 (N_2957,N_942,N_144);
and U2958 (N_2958,N_718,N_16);
or U2959 (N_2959,N_938,N_1609);
nand U2960 (N_2960,N_465,N_500);
nand U2961 (N_2961,N_742,N_1032);
or U2962 (N_2962,N_739,N_3);
nand U2963 (N_2963,N_579,N_953);
and U2964 (N_2964,N_224,N_1542);
and U2965 (N_2965,N_569,N_431);
nor U2966 (N_2966,N_906,N_976);
and U2967 (N_2967,N_638,N_1527);
and U2968 (N_2968,N_1996,N_1867);
or U2969 (N_2969,N_713,N_1790);
nand U2970 (N_2970,N_1423,N_1176);
and U2971 (N_2971,N_1162,N_984);
nor U2972 (N_2972,N_303,N_1763);
nor U2973 (N_2973,N_1824,N_1404);
or U2974 (N_2974,N_87,N_1045);
or U2975 (N_2975,N_196,N_614);
nand U2976 (N_2976,N_478,N_662);
and U2977 (N_2977,N_905,N_325);
and U2978 (N_2978,N_685,N_256);
nor U2979 (N_2979,N_1309,N_1502);
nand U2980 (N_2980,N_1167,N_831);
and U2981 (N_2981,N_527,N_1227);
nor U2982 (N_2982,N_1375,N_1429);
nor U2983 (N_2983,N_324,N_158);
and U2984 (N_2984,N_1990,N_9);
nand U2985 (N_2985,N_872,N_428);
and U2986 (N_2986,N_208,N_1177);
and U2987 (N_2987,N_238,N_1523);
nor U2988 (N_2988,N_1321,N_865);
nand U2989 (N_2989,N_1287,N_727);
nor U2990 (N_2990,N_1376,N_1863);
and U2991 (N_2991,N_1308,N_411);
and U2992 (N_2992,N_1257,N_1382);
nand U2993 (N_2993,N_366,N_959);
or U2994 (N_2994,N_978,N_671);
and U2995 (N_2995,N_438,N_507);
and U2996 (N_2996,N_46,N_768);
nor U2997 (N_2997,N_352,N_1430);
nand U2998 (N_2998,N_1049,N_328);
nand U2999 (N_2999,N_925,N_694);
or U3000 (N_3000,N_1188,N_888);
or U3001 (N_3001,N_374,N_131);
or U3002 (N_3002,N_545,N_57);
nor U3003 (N_3003,N_1151,N_1463);
nor U3004 (N_3004,N_1388,N_963);
nand U3005 (N_3005,N_576,N_1838);
or U3006 (N_3006,N_936,N_354);
nor U3007 (N_3007,N_115,N_233);
nor U3008 (N_3008,N_250,N_672);
nand U3009 (N_3009,N_1208,N_164);
nand U3010 (N_3010,N_857,N_1019);
nor U3011 (N_3011,N_1144,N_17);
nor U3012 (N_3012,N_1470,N_551);
nor U3013 (N_3013,N_1717,N_1351);
nand U3014 (N_3014,N_318,N_713);
and U3015 (N_3015,N_917,N_709);
and U3016 (N_3016,N_1114,N_27);
nor U3017 (N_3017,N_1282,N_220);
or U3018 (N_3018,N_1873,N_480);
nand U3019 (N_3019,N_1462,N_1746);
or U3020 (N_3020,N_1223,N_1963);
or U3021 (N_3021,N_533,N_691);
nand U3022 (N_3022,N_1683,N_1247);
and U3023 (N_3023,N_1306,N_1448);
and U3024 (N_3024,N_506,N_1559);
or U3025 (N_3025,N_1662,N_21);
or U3026 (N_3026,N_1794,N_1524);
and U3027 (N_3027,N_353,N_1776);
nand U3028 (N_3028,N_603,N_175);
or U3029 (N_3029,N_1969,N_354);
nand U3030 (N_3030,N_1119,N_694);
nand U3031 (N_3031,N_1083,N_1732);
nand U3032 (N_3032,N_1518,N_1545);
and U3033 (N_3033,N_1594,N_592);
nor U3034 (N_3034,N_1734,N_315);
and U3035 (N_3035,N_1323,N_63);
and U3036 (N_3036,N_120,N_482);
nor U3037 (N_3037,N_20,N_526);
nand U3038 (N_3038,N_1838,N_914);
or U3039 (N_3039,N_156,N_864);
nor U3040 (N_3040,N_1482,N_50);
and U3041 (N_3041,N_893,N_1567);
or U3042 (N_3042,N_1250,N_1577);
or U3043 (N_3043,N_1255,N_1544);
nor U3044 (N_3044,N_1500,N_74);
nand U3045 (N_3045,N_186,N_1189);
and U3046 (N_3046,N_265,N_334);
or U3047 (N_3047,N_844,N_1545);
xnor U3048 (N_3048,N_905,N_538);
or U3049 (N_3049,N_314,N_27);
xnor U3050 (N_3050,N_1836,N_1652);
nand U3051 (N_3051,N_336,N_1466);
and U3052 (N_3052,N_1457,N_92);
and U3053 (N_3053,N_321,N_1331);
nor U3054 (N_3054,N_1588,N_1103);
nor U3055 (N_3055,N_1822,N_1808);
nand U3056 (N_3056,N_293,N_360);
nor U3057 (N_3057,N_615,N_1238);
and U3058 (N_3058,N_299,N_1334);
or U3059 (N_3059,N_539,N_1891);
and U3060 (N_3060,N_1419,N_1508);
nand U3061 (N_3061,N_246,N_32);
nand U3062 (N_3062,N_1570,N_432);
or U3063 (N_3063,N_1543,N_1175);
or U3064 (N_3064,N_1010,N_838);
or U3065 (N_3065,N_1264,N_257);
nand U3066 (N_3066,N_384,N_350);
nand U3067 (N_3067,N_1875,N_141);
and U3068 (N_3068,N_1889,N_555);
or U3069 (N_3069,N_50,N_1570);
nor U3070 (N_3070,N_1988,N_588);
nor U3071 (N_3071,N_1298,N_1220);
and U3072 (N_3072,N_1269,N_680);
or U3073 (N_3073,N_1862,N_883);
xnor U3074 (N_3074,N_553,N_478);
or U3075 (N_3075,N_1072,N_149);
or U3076 (N_3076,N_1772,N_123);
or U3077 (N_3077,N_442,N_1345);
or U3078 (N_3078,N_1304,N_943);
or U3079 (N_3079,N_417,N_286);
and U3080 (N_3080,N_1879,N_476);
and U3081 (N_3081,N_366,N_881);
nand U3082 (N_3082,N_1764,N_1884);
or U3083 (N_3083,N_1870,N_1896);
nor U3084 (N_3084,N_1547,N_1348);
xor U3085 (N_3085,N_624,N_1817);
nand U3086 (N_3086,N_1851,N_308);
or U3087 (N_3087,N_1100,N_646);
and U3088 (N_3088,N_598,N_69);
nand U3089 (N_3089,N_1471,N_656);
nand U3090 (N_3090,N_215,N_1353);
nand U3091 (N_3091,N_701,N_1827);
nand U3092 (N_3092,N_1449,N_964);
nand U3093 (N_3093,N_797,N_1783);
nand U3094 (N_3094,N_1336,N_197);
nand U3095 (N_3095,N_600,N_1456);
or U3096 (N_3096,N_259,N_1659);
or U3097 (N_3097,N_609,N_967);
or U3098 (N_3098,N_1020,N_118);
nand U3099 (N_3099,N_1457,N_137);
or U3100 (N_3100,N_206,N_1524);
nor U3101 (N_3101,N_1116,N_1253);
nand U3102 (N_3102,N_1254,N_1690);
or U3103 (N_3103,N_1614,N_429);
and U3104 (N_3104,N_1725,N_1267);
nor U3105 (N_3105,N_1338,N_649);
nand U3106 (N_3106,N_1506,N_593);
nand U3107 (N_3107,N_571,N_1606);
and U3108 (N_3108,N_270,N_273);
and U3109 (N_3109,N_1948,N_349);
nor U3110 (N_3110,N_1448,N_1595);
xnor U3111 (N_3111,N_1929,N_1743);
nor U3112 (N_3112,N_659,N_1529);
and U3113 (N_3113,N_1617,N_1906);
or U3114 (N_3114,N_304,N_839);
nand U3115 (N_3115,N_395,N_1034);
or U3116 (N_3116,N_1158,N_1075);
or U3117 (N_3117,N_225,N_1813);
or U3118 (N_3118,N_1670,N_1852);
and U3119 (N_3119,N_1515,N_1154);
or U3120 (N_3120,N_970,N_250);
and U3121 (N_3121,N_1921,N_442);
nand U3122 (N_3122,N_1367,N_1314);
nor U3123 (N_3123,N_871,N_338);
or U3124 (N_3124,N_1239,N_691);
nor U3125 (N_3125,N_1653,N_589);
xor U3126 (N_3126,N_1068,N_695);
and U3127 (N_3127,N_100,N_1737);
or U3128 (N_3128,N_774,N_195);
nand U3129 (N_3129,N_1958,N_194);
or U3130 (N_3130,N_393,N_1872);
and U3131 (N_3131,N_1673,N_1908);
and U3132 (N_3132,N_120,N_1965);
nand U3133 (N_3133,N_1964,N_1459);
nor U3134 (N_3134,N_171,N_1693);
nand U3135 (N_3135,N_1793,N_518);
or U3136 (N_3136,N_660,N_1635);
nand U3137 (N_3137,N_960,N_1531);
nand U3138 (N_3138,N_307,N_930);
or U3139 (N_3139,N_1300,N_897);
and U3140 (N_3140,N_1063,N_656);
or U3141 (N_3141,N_1864,N_805);
and U3142 (N_3142,N_1996,N_774);
nor U3143 (N_3143,N_604,N_1733);
and U3144 (N_3144,N_88,N_1048);
nor U3145 (N_3145,N_1349,N_559);
or U3146 (N_3146,N_1830,N_1302);
or U3147 (N_3147,N_1662,N_1409);
nor U3148 (N_3148,N_1298,N_1143);
or U3149 (N_3149,N_582,N_1403);
and U3150 (N_3150,N_1476,N_978);
nand U3151 (N_3151,N_1559,N_679);
nor U3152 (N_3152,N_866,N_525);
or U3153 (N_3153,N_1793,N_581);
nand U3154 (N_3154,N_1350,N_1155);
xor U3155 (N_3155,N_1162,N_1577);
nand U3156 (N_3156,N_220,N_1020);
and U3157 (N_3157,N_1027,N_553);
or U3158 (N_3158,N_37,N_1460);
nand U3159 (N_3159,N_1646,N_1814);
nor U3160 (N_3160,N_131,N_92);
and U3161 (N_3161,N_304,N_928);
nand U3162 (N_3162,N_1198,N_289);
or U3163 (N_3163,N_1732,N_655);
or U3164 (N_3164,N_521,N_1787);
nor U3165 (N_3165,N_628,N_440);
or U3166 (N_3166,N_145,N_1896);
or U3167 (N_3167,N_1096,N_1800);
nor U3168 (N_3168,N_1099,N_413);
or U3169 (N_3169,N_864,N_495);
or U3170 (N_3170,N_479,N_519);
xnor U3171 (N_3171,N_1652,N_204);
nor U3172 (N_3172,N_610,N_765);
and U3173 (N_3173,N_1607,N_79);
and U3174 (N_3174,N_1268,N_160);
and U3175 (N_3175,N_435,N_604);
or U3176 (N_3176,N_942,N_537);
nand U3177 (N_3177,N_562,N_43);
nand U3178 (N_3178,N_1022,N_409);
nand U3179 (N_3179,N_958,N_126);
or U3180 (N_3180,N_740,N_1901);
nand U3181 (N_3181,N_1032,N_521);
or U3182 (N_3182,N_1544,N_470);
nand U3183 (N_3183,N_1903,N_1449);
or U3184 (N_3184,N_268,N_755);
nor U3185 (N_3185,N_1557,N_440);
nor U3186 (N_3186,N_879,N_1467);
and U3187 (N_3187,N_708,N_1210);
xor U3188 (N_3188,N_1916,N_402);
nand U3189 (N_3189,N_1021,N_300);
and U3190 (N_3190,N_637,N_830);
nand U3191 (N_3191,N_457,N_1573);
nor U3192 (N_3192,N_556,N_316);
or U3193 (N_3193,N_336,N_833);
nand U3194 (N_3194,N_1001,N_235);
nor U3195 (N_3195,N_153,N_8);
or U3196 (N_3196,N_796,N_396);
nand U3197 (N_3197,N_497,N_1969);
nand U3198 (N_3198,N_1335,N_1074);
nor U3199 (N_3199,N_787,N_279);
nand U3200 (N_3200,N_1451,N_1861);
and U3201 (N_3201,N_1963,N_1782);
or U3202 (N_3202,N_1310,N_854);
and U3203 (N_3203,N_1780,N_872);
nor U3204 (N_3204,N_539,N_797);
nor U3205 (N_3205,N_1994,N_123);
nor U3206 (N_3206,N_1943,N_590);
and U3207 (N_3207,N_352,N_1794);
or U3208 (N_3208,N_400,N_1955);
or U3209 (N_3209,N_351,N_1781);
or U3210 (N_3210,N_1199,N_857);
and U3211 (N_3211,N_1651,N_1978);
nand U3212 (N_3212,N_1286,N_230);
nor U3213 (N_3213,N_1103,N_72);
nand U3214 (N_3214,N_941,N_809);
or U3215 (N_3215,N_783,N_1187);
nor U3216 (N_3216,N_970,N_237);
nand U3217 (N_3217,N_1276,N_50);
or U3218 (N_3218,N_1181,N_1167);
nor U3219 (N_3219,N_299,N_521);
nand U3220 (N_3220,N_1605,N_839);
nand U3221 (N_3221,N_1237,N_1901);
nor U3222 (N_3222,N_123,N_1479);
nor U3223 (N_3223,N_495,N_725);
nand U3224 (N_3224,N_1319,N_7);
nor U3225 (N_3225,N_203,N_827);
or U3226 (N_3226,N_1535,N_788);
nand U3227 (N_3227,N_514,N_401);
nand U3228 (N_3228,N_1072,N_232);
nor U3229 (N_3229,N_572,N_1846);
nor U3230 (N_3230,N_52,N_864);
nand U3231 (N_3231,N_1647,N_917);
or U3232 (N_3232,N_427,N_287);
nand U3233 (N_3233,N_965,N_1650);
nor U3234 (N_3234,N_84,N_1470);
nand U3235 (N_3235,N_682,N_373);
nand U3236 (N_3236,N_1059,N_1331);
nand U3237 (N_3237,N_228,N_1804);
nand U3238 (N_3238,N_434,N_1054);
and U3239 (N_3239,N_534,N_663);
nand U3240 (N_3240,N_1439,N_824);
and U3241 (N_3241,N_1646,N_1238);
and U3242 (N_3242,N_1254,N_622);
and U3243 (N_3243,N_889,N_1485);
or U3244 (N_3244,N_1040,N_1690);
nor U3245 (N_3245,N_1196,N_1467);
or U3246 (N_3246,N_1622,N_1467);
nand U3247 (N_3247,N_1033,N_1401);
nand U3248 (N_3248,N_1441,N_1342);
and U3249 (N_3249,N_240,N_1840);
nand U3250 (N_3250,N_386,N_651);
nor U3251 (N_3251,N_411,N_983);
nor U3252 (N_3252,N_1740,N_600);
and U3253 (N_3253,N_1108,N_1402);
nand U3254 (N_3254,N_1445,N_1607);
nand U3255 (N_3255,N_1229,N_38);
nor U3256 (N_3256,N_718,N_1206);
nor U3257 (N_3257,N_727,N_408);
or U3258 (N_3258,N_1730,N_1686);
xor U3259 (N_3259,N_158,N_1367);
and U3260 (N_3260,N_1217,N_1342);
and U3261 (N_3261,N_1247,N_797);
or U3262 (N_3262,N_682,N_937);
xnor U3263 (N_3263,N_519,N_1980);
or U3264 (N_3264,N_1851,N_1419);
and U3265 (N_3265,N_193,N_600);
and U3266 (N_3266,N_74,N_527);
and U3267 (N_3267,N_571,N_1145);
nor U3268 (N_3268,N_1710,N_1909);
or U3269 (N_3269,N_1976,N_162);
nor U3270 (N_3270,N_1753,N_1670);
or U3271 (N_3271,N_1508,N_919);
or U3272 (N_3272,N_745,N_951);
nand U3273 (N_3273,N_640,N_232);
and U3274 (N_3274,N_717,N_267);
and U3275 (N_3275,N_465,N_1053);
and U3276 (N_3276,N_512,N_341);
or U3277 (N_3277,N_714,N_1087);
nand U3278 (N_3278,N_45,N_1549);
nand U3279 (N_3279,N_1032,N_1675);
or U3280 (N_3280,N_1550,N_678);
nand U3281 (N_3281,N_1236,N_761);
nand U3282 (N_3282,N_1001,N_809);
or U3283 (N_3283,N_1496,N_1346);
or U3284 (N_3284,N_1863,N_844);
and U3285 (N_3285,N_1631,N_851);
and U3286 (N_3286,N_1548,N_1215);
nor U3287 (N_3287,N_273,N_495);
or U3288 (N_3288,N_1786,N_837);
and U3289 (N_3289,N_1704,N_161);
and U3290 (N_3290,N_1350,N_556);
and U3291 (N_3291,N_1095,N_971);
nor U3292 (N_3292,N_563,N_1789);
nor U3293 (N_3293,N_369,N_215);
nand U3294 (N_3294,N_1293,N_268);
nand U3295 (N_3295,N_802,N_954);
nor U3296 (N_3296,N_1466,N_763);
nand U3297 (N_3297,N_736,N_399);
nand U3298 (N_3298,N_1794,N_456);
nand U3299 (N_3299,N_423,N_922);
nor U3300 (N_3300,N_1295,N_652);
or U3301 (N_3301,N_1404,N_1652);
and U3302 (N_3302,N_696,N_1648);
nand U3303 (N_3303,N_163,N_1855);
or U3304 (N_3304,N_722,N_919);
and U3305 (N_3305,N_631,N_957);
or U3306 (N_3306,N_1472,N_745);
nand U3307 (N_3307,N_1832,N_488);
nor U3308 (N_3308,N_84,N_1946);
or U3309 (N_3309,N_126,N_1303);
nor U3310 (N_3310,N_289,N_1390);
nand U3311 (N_3311,N_1993,N_1559);
nor U3312 (N_3312,N_357,N_1311);
nor U3313 (N_3313,N_1829,N_1631);
and U3314 (N_3314,N_861,N_1361);
and U3315 (N_3315,N_1938,N_1689);
or U3316 (N_3316,N_1719,N_1519);
nor U3317 (N_3317,N_1687,N_438);
nand U3318 (N_3318,N_1027,N_1726);
or U3319 (N_3319,N_1698,N_1781);
nand U3320 (N_3320,N_1514,N_1321);
or U3321 (N_3321,N_1267,N_136);
nor U3322 (N_3322,N_39,N_733);
xor U3323 (N_3323,N_1458,N_1309);
nand U3324 (N_3324,N_149,N_479);
and U3325 (N_3325,N_938,N_48);
and U3326 (N_3326,N_575,N_1410);
xnor U3327 (N_3327,N_240,N_1437);
and U3328 (N_3328,N_395,N_1703);
and U3329 (N_3329,N_1389,N_530);
or U3330 (N_3330,N_1672,N_867);
or U3331 (N_3331,N_787,N_193);
nand U3332 (N_3332,N_1597,N_1656);
xnor U3333 (N_3333,N_631,N_1020);
nor U3334 (N_3334,N_1500,N_1056);
or U3335 (N_3335,N_848,N_769);
or U3336 (N_3336,N_672,N_1582);
nand U3337 (N_3337,N_1185,N_1493);
nor U3338 (N_3338,N_527,N_1562);
and U3339 (N_3339,N_38,N_1748);
or U3340 (N_3340,N_591,N_821);
or U3341 (N_3341,N_935,N_182);
and U3342 (N_3342,N_43,N_1583);
nand U3343 (N_3343,N_1442,N_1705);
nor U3344 (N_3344,N_1615,N_514);
nand U3345 (N_3345,N_491,N_1395);
nand U3346 (N_3346,N_1984,N_1734);
nor U3347 (N_3347,N_991,N_673);
nand U3348 (N_3348,N_1803,N_688);
nor U3349 (N_3349,N_1766,N_1602);
and U3350 (N_3350,N_854,N_131);
and U3351 (N_3351,N_1195,N_1953);
nand U3352 (N_3352,N_204,N_616);
or U3353 (N_3353,N_1215,N_740);
or U3354 (N_3354,N_324,N_746);
nand U3355 (N_3355,N_1477,N_530);
or U3356 (N_3356,N_1182,N_192);
or U3357 (N_3357,N_899,N_703);
or U3358 (N_3358,N_783,N_1469);
or U3359 (N_3359,N_1555,N_1824);
or U3360 (N_3360,N_1918,N_762);
or U3361 (N_3361,N_132,N_268);
nand U3362 (N_3362,N_1935,N_1328);
nand U3363 (N_3363,N_1445,N_1369);
xnor U3364 (N_3364,N_547,N_769);
nand U3365 (N_3365,N_624,N_115);
nand U3366 (N_3366,N_312,N_384);
xor U3367 (N_3367,N_1316,N_1010);
nand U3368 (N_3368,N_851,N_1185);
or U3369 (N_3369,N_350,N_50);
nor U3370 (N_3370,N_1507,N_1124);
and U3371 (N_3371,N_1595,N_1287);
or U3372 (N_3372,N_753,N_605);
or U3373 (N_3373,N_244,N_1879);
nand U3374 (N_3374,N_613,N_730);
nand U3375 (N_3375,N_914,N_1581);
xor U3376 (N_3376,N_1924,N_1537);
and U3377 (N_3377,N_569,N_1000);
or U3378 (N_3378,N_1498,N_1286);
nor U3379 (N_3379,N_764,N_1651);
or U3380 (N_3380,N_1626,N_438);
and U3381 (N_3381,N_229,N_1886);
nor U3382 (N_3382,N_1316,N_779);
nand U3383 (N_3383,N_94,N_1833);
nor U3384 (N_3384,N_403,N_1854);
and U3385 (N_3385,N_1451,N_1979);
xor U3386 (N_3386,N_564,N_1271);
or U3387 (N_3387,N_503,N_806);
or U3388 (N_3388,N_1974,N_204);
nand U3389 (N_3389,N_1342,N_1847);
or U3390 (N_3390,N_1603,N_41);
nor U3391 (N_3391,N_1382,N_1952);
nor U3392 (N_3392,N_671,N_71);
nand U3393 (N_3393,N_592,N_46);
nand U3394 (N_3394,N_1648,N_1364);
and U3395 (N_3395,N_1995,N_926);
and U3396 (N_3396,N_1567,N_1993);
or U3397 (N_3397,N_421,N_854);
or U3398 (N_3398,N_1271,N_1135);
and U3399 (N_3399,N_100,N_168);
or U3400 (N_3400,N_365,N_1224);
nor U3401 (N_3401,N_740,N_548);
and U3402 (N_3402,N_641,N_676);
or U3403 (N_3403,N_292,N_571);
nor U3404 (N_3404,N_223,N_649);
or U3405 (N_3405,N_1773,N_1892);
and U3406 (N_3406,N_1384,N_1187);
and U3407 (N_3407,N_1091,N_1342);
and U3408 (N_3408,N_707,N_51);
or U3409 (N_3409,N_1827,N_1098);
nor U3410 (N_3410,N_1981,N_607);
and U3411 (N_3411,N_1299,N_94);
nor U3412 (N_3412,N_1308,N_132);
nor U3413 (N_3413,N_885,N_79);
nand U3414 (N_3414,N_342,N_963);
or U3415 (N_3415,N_1619,N_453);
or U3416 (N_3416,N_1091,N_1353);
or U3417 (N_3417,N_1902,N_528);
nor U3418 (N_3418,N_245,N_1239);
nand U3419 (N_3419,N_646,N_1911);
nor U3420 (N_3420,N_1156,N_1855);
nor U3421 (N_3421,N_1375,N_985);
and U3422 (N_3422,N_1659,N_483);
or U3423 (N_3423,N_863,N_1519);
nand U3424 (N_3424,N_856,N_1611);
and U3425 (N_3425,N_1346,N_327);
and U3426 (N_3426,N_1790,N_1753);
and U3427 (N_3427,N_1271,N_511);
nor U3428 (N_3428,N_1119,N_1714);
or U3429 (N_3429,N_898,N_952);
and U3430 (N_3430,N_1000,N_1582);
nand U3431 (N_3431,N_1763,N_280);
and U3432 (N_3432,N_246,N_1978);
and U3433 (N_3433,N_344,N_1056);
nor U3434 (N_3434,N_1100,N_1316);
nor U3435 (N_3435,N_552,N_99);
or U3436 (N_3436,N_1068,N_1394);
and U3437 (N_3437,N_1302,N_228);
nor U3438 (N_3438,N_771,N_1291);
and U3439 (N_3439,N_1049,N_5);
and U3440 (N_3440,N_179,N_1701);
nand U3441 (N_3441,N_816,N_146);
nand U3442 (N_3442,N_1552,N_559);
or U3443 (N_3443,N_974,N_552);
nand U3444 (N_3444,N_1573,N_816);
nand U3445 (N_3445,N_657,N_1034);
nand U3446 (N_3446,N_273,N_362);
nand U3447 (N_3447,N_1910,N_709);
and U3448 (N_3448,N_608,N_1209);
or U3449 (N_3449,N_130,N_1619);
or U3450 (N_3450,N_1932,N_1148);
and U3451 (N_3451,N_1073,N_78);
nor U3452 (N_3452,N_1539,N_129);
and U3453 (N_3453,N_1957,N_448);
or U3454 (N_3454,N_196,N_1376);
and U3455 (N_3455,N_876,N_1792);
nand U3456 (N_3456,N_177,N_207);
nor U3457 (N_3457,N_973,N_841);
nand U3458 (N_3458,N_671,N_1516);
nand U3459 (N_3459,N_110,N_199);
and U3460 (N_3460,N_1526,N_295);
nor U3461 (N_3461,N_414,N_399);
nand U3462 (N_3462,N_806,N_1958);
and U3463 (N_3463,N_1691,N_100);
and U3464 (N_3464,N_296,N_364);
and U3465 (N_3465,N_271,N_1713);
and U3466 (N_3466,N_1615,N_1632);
nand U3467 (N_3467,N_1185,N_1652);
and U3468 (N_3468,N_724,N_1687);
nand U3469 (N_3469,N_263,N_926);
or U3470 (N_3470,N_1087,N_65);
xor U3471 (N_3471,N_401,N_405);
or U3472 (N_3472,N_1694,N_1759);
or U3473 (N_3473,N_616,N_1286);
nand U3474 (N_3474,N_381,N_1230);
nand U3475 (N_3475,N_1206,N_1594);
or U3476 (N_3476,N_1036,N_1468);
and U3477 (N_3477,N_22,N_1551);
and U3478 (N_3478,N_1620,N_253);
nor U3479 (N_3479,N_740,N_818);
or U3480 (N_3480,N_224,N_598);
nor U3481 (N_3481,N_1612,N_1738);
nor U3482 (N_3482,N_688,N_776);
and U3483 (N_3483,N_1877,N_936);
and U3484 (N_3484,N_1689,N_794);
or U3485 (N_3485,N_935,N_51);
or U3486 (N_3486,N_1994,N_1397);
nor U3487 (N_3487,N_473,N_262);
xor U3488 (N_3488,N_1198,N_1821);
or U3489 (N_3489,N_1124,N_207);
or U3490 (N_3490,N_1841,N_631);
nor U3491 (N_3491,N_1687,N_380);
nand U3492 (N_3492,N_860,N_133);
nand U3493 (N_3493,N_1087,N_603);
nor U3494 (N_3494,N_718,N_285);
and U3495 (N_3495,N_209,N_1187);
nor U3496 (N_3496,N_1468,N_1943);
nor U3497 (N_3497,N_1268,N_13);
nand U3498 (N_3498,N_9,N_1971);
nor U3499 (N_3499,N_685,N_1114);
nor U3500 (N_3500,N_1490,N_1605);
nor U3501 (N_3501,N_474,N_1530);
nand U3502 (N_3502,N_80,N_1418);
or U3503 (N_3503,N_1233,N_871);
nor U3504 (N_3504,N_1644,N_1358);
or U3505 (N_3505,N_492,N_1945);
or U3506 (N_3506,N_1031,N_175);
and U3507 (N_3507,N_1107,N_225);
nor U3508 (N_3508,N_1971,N_383);
xnor U3509 (N_3509,N_584,N_922);
nand U3510 (N_3510,N_378,N_884);
nand U3511 (N_3511,N_1386,N_1142);
nand U3512 (N_3512,N_1943,N_68);
nand U3513 (N_3513,N_51,N_119);
or U3514 (N_3514,N_1689,N_995);
or U3515 (N_3515,N_742,N_1386);
nor U3516 (N_3516,N_1280,N_244);
xnor U3517 (N_3517,N_57,N_1419);
and U3518 (N_3518,N_273,N_1400);
nor U3519 (N_3519,N_1938,N_640);
and U3520 (N_3520,N_1003,N_1758);
and U3521 (N_3521,N_1144,N_1003);
nand U3522 (N_3522,N_43,N_841);
nand U3523 (N_3523,N_1711,N_792);
nor U3524 (N_3524,N_1724,N_1707);
and U3525 (N_3525,N_1878,N_1314);
nor U3526 (N_3526,N_1528,N_1842);
and U3527 (N_3527,N_1774,N_1843);
nand U3528 (N_3528,N_1145,N_461);
or U3529 (N_3529,N_1712,N_297);
nor U3530 (N_3530,N_1287,N_1853);
or U3531 (N_3531,N_1189,N_1611);
nand U3532 (N_3532,N_214,N_1339);
nand U3533 (N_3533,N_578,N_105);
or U3534 (N_3534,N_1859,N_203);
nand U3535 (N_3535,N_653,N_1471);
or U3536 (N_3536,N_1882,N_328);
or U3537 (N_3537,N_1720,N_109);
or U3538 (N_3538,N_1059,N_1344);
nor U3539 (N_3539,N_651,N_1618);
nand U3540 (N_3540,N_199,N_1509);
nand U3541 (N_3541,N_236,N_1034);
and U3542 (N_3542,N_512,N_1977);
nor U3543 (N_3543,N_1311,N_566);
and U3544 (N_3544,N_1634,N_716);
and U3545 (N_3545,N_790,N_1484);
nand U3546 (N_3546,N_1117,N_1933);
nand U3547 (N_3547,N_152,N_37);
and U3548 (N_3548,N_157,N_1107);
nand U3549 (N_3549,N_929,N_1234);
and U3550 (N_3550,N_952,N_244);
and U3551 (N_3551,N_1394,N_580);
nor U3552 (N_3552,N_299,N_1116);
and U3553 (N_3553,N_301,N_521);
and U3554 (N_3554,N_1729,N_1412);
and U3555 (N_3555,N_1556,N_599);
nand U3556 (N_3556,N_441,N_588);
or U3557 (N_3557,N_997,N_1767);
nor U3558 (N_3558,N_430,N_1466);
nor U3559 (N_3559,N_1173,N_115);
nand U3560 (N_3560,N_763,N_1080);
and U3561 (N_3561,N_1350,N_1636);
nor U3562 (N_3562,N_527,N_975);
or U3563 (N_3563,N_269,N_1068);
nand U3564 (N_3564,N_1570,N_1210);
and U3565 (N_3565,N_82,N_547);
or U3566 (N_3566,N_714,N_1848);
nor U3567 (N_3567,N_137,N_983);
or U3568 (N_3568,N_535,N_1718);
and U3569 (N_3569,N_1426,N_1614);
and U3570 (N_3570,N_1390,N_754);
or U3571 (N_3571,N_1506,N_1810);
and U3572 (N_3572,N_1856,N_623);
nand U3573 (N_3573,N_778,N_1065);
nand U3574 (N_3574,N_1450,N_1887);
nor U3575 (N_3575,N_1515,N_441);
nand U3576 (N_3576,N_718,N_670);
and U3577 (N_3577,N_1178,N_204);
or U3578 (N_3578,N_341,N_1534);
nand U3579 (N_3579,N_1649,N_1042);
and U3580 (N_3580,N_150,N_855);
and U3581 (N_3581,N_1807,N_1119);
nand U3582 (N_3582,N_270,N_324);
or U3583 (N_3583,N_69,N_1891);
nand U3584 (N_3584,N_204,N_187);
or U3585 (N_3585,N_303,N_1134);
nand U3586 (N_3586,N_220,N_978);
nand U3587 (N_3587,N_742,N_383);
or U3588 (N_3588,N_39,N_268);
and U3589 (N_3589,N_931,N_421);
nand U3590 (N_3590,N_1799,N_820);
and U3591 (N_3591,N_1488,N_554);
nand U3592 (N_3592,N_483,N_524);
nor U3593 (N_3593,N_30,N_120);
or U3594 (N_3594,N_1560,N_1414);
and U3595 (N_3595,N_496,N_451);
nand U3596 (N_3596,N_1246,N_729);
and U3597 (N_3597,N_63,N_153);
and U3598 (N_3598,N_1611,N_1289);
nand U3599 (N_3599,N_1881,N_383);
or U3600 (N_3600,N_1446,N_1753);
or U3601 (N_3601,N_1220,N_1473);
nor U3602 (N_3602,N_1995,N_1463);
nor U3603 (N_3603,N_615,N_1892);
and U3604 (N_3604,N_1621,N_248);
and U3605 (N_3605,N_424,N_970);
and U3606 (N_3606,N_584,N_413);
or U3607 (N_3607,N_346,N_1778);
nor U3608 (N_3608,N_537,N_1797);
or U3609 (N_3609,N_853,N_1237);
nand U3610 (N_3610,N_66,N_107);
nor U3611 (N_3611,N_1822,N_1755);
and U3612 (N_3612,N_930,N_826);
and U3613 (N_3613,N_1605,N_585);
or U3614 (N_3614,N_63,N_515);
nor U3615 (N_3615,N_732,N_802);
xnor U3616 (N_3616,N_837,N_1904);
nand U3617 (N_3617,N_565,N_1376);
nand U3618 (N_3618,N_1665,N_315);
nor U3619 (N_3619,N_1386,N_489);
nor U3620 (N_3620,N_418,N_1394);
nand U3621 (N_3621,N_998,N_1595);
and U3622 (N_3622,N_1268,N_434);
nor U3623 (N_3623,N_1559,N_798);
nand U3624 (N_3624,N_894,N_1014);
or U3625 (N_3625,N_467,N_1414);
or U3626 (N_3626,N_927,N_1686);
and U3627 (N_3627,N_855,N_322);
nor U3628 (N_3628,N_1822,N_1383);
and U3629 (N_3629,N_34,N_542);
or U3630 (N_3630,N_345,N_494);
nor U3631 (N_3631,N_130,N_1898);
nand U3632 (N_3632,N_1120,N_600);
and U3633 (N_3633,N_719,N_1529);
nand U3634 (N_3634,N_1508,N_516);
and U3635 (N_3635,N_761,N_10);
and U3636 (N_3636,N_1800,N_867);
and U3637 (N_3637,N_1901,N_544);
and U3638 (N_3638,N_1473,N_560);
nor U3639 (N_3639,N_44,N_283);
nand U3640 (N_3640,N_734,N_852);
or U3641 (N_3641,N_539,N_1366);
and U3642 (N_3642,N_4,N_96);
nor U3643 (N_3643,N_1336,N_1596);
nor U3644 (N_3644,N_537,N_638);
nand U3645 (N_3645,N_1700,N_1569);
nand U3646 (N_3646,N_476,N_769);
nand U3647 (N_3647,N_907,N_332);
or U3648 (N_3648,N_1809,N_20);
or U3649 (N_3649,N_1374,N_1129);
nor U3650 (N_3650,N_1762,N_1100);
or U3651 (N_3651,N_1639,N_1496);
nand U3652 (N_3652,N_1017,N_797);
nand U3653 (N_3653,N_652,N_1924);
and U3654 (N_3654,N_11,N_1008);
nor U3655 (N_3655,N_1216,N_1661);
nor U3656 (N_3656,N_697,N_594);
nand U3657 (N_3657,N_1652,N_1415);
nand U3658 (N_3658,N_39,N_685);
or U3659 (N_3659,N_1152,N_1547);
and U3660 (N_3660,N_1299,N_719);
and U3661 (N_3661,N_1012,N_344);
and U3662 (N_3662,N_1139,N_413);
nand U3663 (N_3663,N_901,N_1254);
or U3664 (N_3664,N_148,N_1655);
nor U3665 (N_3665,N_1841,N_1311);
or U3666 (N_3666,N_1921,N_586);
nand U3667 (N_3667,N_578,N_403);
nor U3668 (N_3668,N_1675,N_1521);
and U3669 (N_3669,N_506,N_275);
or U3670 (N_3670,N_1324,N_570);
and U3671 (N_3671,N_577,N_1787);
nand U3672 (N_3672,N_1447,N_1809);
nor U3673 (N_3673,N_1842,N_1105);
or U3674 (N_3674,N_1464,N_1169);
and U3675 (N_3675,N_744,N_484);
nand U3676 (N_3676,N_1132,N_1268);
nor U3677 (N_3677,N_1336,N_560);
nand U3678 (N_3678,N_1652,N_791);
nand U3679 (N_3679,N_853,N_983);
or U3680 (N_3680,N_262,N_933);
nand U3681 (N_3681,N_1694,N_186);
and U3682 (N_3682,N_374,N_629);
and U3683 (N_3683,N_522,N_967);
and U3684 (N_3684,N_1160,N_870);
nand U3685 (N_3685,N_1917,N_1986);
nand U3686 (N_3686,N_331,N_512);
and U3687 (N_3687,N_984,N_1971);
nand U3688 (N_3688,N_1,N_1143);
or U3689 (N_3689,N_1565,N_930);
nand U3690 (N_3690,N_1362,N_299);
or U3691 (N_3691,N_11,N_1208);
or U3692 (N_3692,N_955,N_153);
nand U3693 (N_3693,N_702,N_407);
nor U3694 (N_3694,N_854,N_708);
and U3695 (N_3695,N_788,N_190);
and U3696 (N_3696,N_535,N_69);
or U3697 (N_3697,N_809,N_1206);
and U3698 (N_3698,N_157,N_724);
xnor U3699 (N_3699,N_750,N_374);
nor U3700 (N_3700,N_372,N_1792);
nor U3701 (N_3701,N_392,N_451);
and U3702 (N_3702,N_116,N_21);
nand U3703 (N_3703,N_1583,N_1059);
nand U3704 (N_3704,N_278,N_1776);
and U3705 (N_3705,N_596,N_904);
or U3706 (N_3706,N_1071,N_151);
or U3707 (N_3707,N_1864,N_707);
or U3708 (N_3708,N_140,N_826);
and U3709 (N_3709,N_1683,N_1731);
nor U3710 (N_3710,N_1813,N_885);
nor U3711 (N_3711,N_1814,N_1109);
nor U3712 (N_3712,N_1814,N_1566);
or U3713 (N_3713,N_912,N_313);
nand U3714 (N_3714,N_1987,N_60);
nor U3715 (N_3715,N_964,N_1129);
or U3716 (N_3716,N_1386,N_1415);
xnor U3717 (N_3717,N_941,N_603);
nor U3718 (N_3718,N_1564,N_56);
and U3719 (N_3719,N_1388,N_1102);
nand U3720 (N_3720,N_1156,N_4);
or U3721 (N_3721,N_289,N_805);
or U3722 (N_3722,N_1908,N_1730);
nor U3723 (N_3723,N_427,N_547);
nor U3724 (N_3724,N_321,N_135);
or U3725 (N_3725,N_1411,N_1113);
nand U3726 (N_3726,N_973,N_313);
nor U3727 (N_3727,N_921,N_836);
and U3728 (N_3728,N_1527,N_767);
or U3729 (N_3729,N_417,N_1704);
nor U3730 (N_3730,N_1316,N_990);
and U3731 (N_3731,N_1034,N_1250);
and U3732 (N_3732,N_1045,N_641);
or U3733 (N_3733,N_717,N_1202);
xnor U3734 (N_3734,N_932,N_1969);
or U3735 (N_3735,N_939,N_217);
and U3736 (N_3736,N_753,N_1999);
nand U3737 (N_3737,N_706,N_894);
and U3738 (N_3738,N_655,N_1392);
nand U3739 (N_3739,N_388,N_605);
and U3740 (N_3740,N_1976,N_1410);
nand U3741 (N_3741,N_1863,N_579);
or U3742 (N_3742,N_1058,N_1123);
nor U3743 (N_3743,N_1797,N_1471);
nand U3744 (N_3744,N_1359,N_277);
nand U3745 (N_3745,N_1056,N_1600);
nor U3746 (N_3746,N_1300,N_1243);
nand U3747 (N_3747,N_1356,N_1108);
or U3748 (N_3748,N_363,N_1554);
and U3749 (N_3749,N_807,N_1730);
or U3750 (N_3750,N_1549,N_325);
nor U3751 (N_3751,N_772,N_1323);
xor U3752 (N_3752,N_1462,N_201);
nor U3753 (N_3753,N_990,N_252);
and U3754 (N_3754,N_167,N_612);
and U3755 (N_3755,N_1464,N_469);
nand U3756 (N_3756,N_174,N_822);
or U3757 (N_3757,N_1875,N_1894);
and U3758 (N_3758,N_80,N_490);
or U3759 (N_3759,N_1798,N_1382);
or U3760 (N_3760,N_598,N_1911);
and U3761 (N_3761,N_1357,N_1244);
nand U3762 (N_3762,N_1371,N_1872);
or U3763 (N_3763,N_752,N_1127);
and U3764 (N_3764,N_508,N_984);
nand U3765 (N_3765,N_249,N_197);
and U3766 (N_3766,N_529,N_59);
and U3767 (N_3767,N_1226,N_796);
and U3768 (N_3768,N_152,N_759);
nand U3769 (N_3769,N_1503,N_11);
or U3770 (N_3770,N_901,N_1010);
nor U3771 (N_3771,N_518,N_169);
nor U3772 (N_3772,N_1277,N_504);
or U3773 (N_3773,N_489,N_1284);
xnor U3774 (N_3774,N_902,N_1009);
xnor U3775 (N_3775,N_1668,N_829);
nand U3776 (N_3776,N_851,N_648);
and U3777 (N_3777,N_491,N_1925);
nand U3778 (N_3778,N_1420,N_1934);
and U3779 (N_3779,N_414,N_1021);
nor U3780 (N_3780,N_813,N_1714);
nand U3781 (N_3781,N_1323,N_1084);
nand U3782 (N_3782,N_455,N_1614);
xnor U3783 (N_3783,N_70,N_933);
and U3784 (N_3784,N_604,N_1180);
nor U3785 (N_3785,N_1976,N_229);
nor U3786 (N_3786,N_1341,N_665);
nand U3787 (N_3787,N_1022,N_589);
nand U3788 (N_3788,N_725,N_486);
and U3789 (N_3789,N_1421,N_1887);
or U3790 (N_3790,N_1458,N_219);
nand U3791 (N_3791,N_1299,N_747);
nand U3792 (N_3792,N_1011,N_179);
nor U3793 (N_3793,N_175,N_927);
and U3794 (N_3794,N_1715,N_532);
and U3795 (N_3795,N_1881,N_538);
and U3796 (N_3796,N_600,N_1970);
nand U3797 (N_3797,N_1073,N_1374);
and U3798 (N_3798,N_255,N_1170);
nand U3799 (N_3799,N_1543,N_182);
and U3800 (N_3800,N_1102,N_37);
and U3801 (N_3801,N_240,N_198);
and U3802 (N_3802,N_91,N_1183);
nor U3803 (N_3803,N_1860,N_1294);
and U3804 (N_3804,N_268,N_1071);
or U3805 (N_3805,N_1038,N_1220);
or U3806 (N_3806,N_132,N_867);
and U3807 (N_3807,N_1837,N_312);
or U3808 (N_3808,N_19,N_591);
nor U3809 (N_3809,N_70,N_97);
and U3810 (N_3810,N_893,N_33);
or U3811 (N_3811,N_1199,N_349);
or U3812 (N_3812,N_541,N_1507);
nand U3813 (N_3813,N_1692,N_751);
nor U3814 (N_3814,N_384,N_995);
and U3815 (N_3815,N_1820,N_1270);
nor U3816 (N_3816,N_331,N_1424);
or U3817 (N_3817,N_400,N_1984);
and U3818 (N_3818,N_835,N_1198);
nor U3819 (N_3819,N_821,N_951);
nand U3820 (N_3820,N_1522,N_1986);
nand U3821 (N_3821,N_631,N_611);
or U3822 (N_3822,N_1575,N_1193);
nor U3823 (N_3823,N_462,N_716);
nand U3824 (N_3824,N_1357,N_332);
and U3825 (N_3825,N_636,N_268);
nor U3826 (N_3826,N_48,N_1048);
or U3827 (N_3827,N_974,N_1441);
and U3828 (N_3828,N_1556,N_531);
xnor U3829 (N_3829,N_1939,N_1459);
and U3830 (N_3830,N_1322,N_691);
or U3831 (N_3831,N_1604,N_282);
xor U3832 (N_3832,N_948,N_1013);
or U3833 (N_3833,N_275,N_953);
or U3834 (N_3834,N_804,N_1551);
xor U3835 (N_3835,N_1193,N_1802);
nor U3836 (N_3836,N_1364,N_1953);
and U3837 (N_3837,N_995,N_603);
nand U3838 (N_3838,N_472,N_313);
and U3839 (N_3839,N_1623,N_227);
nand U3840 (N_3840,N_133,N_1475);
nand U3841 (N_3841,N_1266,N_1443);
nand U3842 (N_3842,N_1525,N_1167);
nand U3843 (N_3843,N_1066,N_373);
and U3844 (N_3844,N_380,N_1510);
and U3845 (N_3845,N_389,N_595);
xnor U3846 (N_3846,N_1642,N_956);
nand U3847 (N_3847,N_1950,N_1768);
nand U3848 (N_3848,N_262,N_939);
nor U3849 (N_3849,N_835,N_875);
nand U3850 (N_3850,N_411,N_197);
nand U3851 (N_3851,N_1581,N_973);
nand U3852 (N_3852,N_1387,N_126);
xnor U3853 (N_3853,N_300,N_720);
or U3854 (N_3854,N_95,N_1116);
nor U3855 (N_3855,N_673,N_644);
nand U3856 (N_3856,N_682,N_1603);
nand U3857 (N_3857,N_1573,N_25);
or U3858 (N_3858,N_807,N_993);
and U3859 (N_3859,N_1281,N_683);
or U3860 (N_3860,N_595,N_1168);
or U3861 (N_3861,N_200,N_1385);
nor U3862 (N_3862,N_1085,N_1511);
and U3863 (N_3863,N_702,N_74);
nor U3864 (N_3864,N_866,N_1522);
and U3865 (N_3865,N_1760,N_743);
nand U3866 (N_3866,N_495,N_1294);
and U3867 (N_3867,N_568,N_446);
or U3868 (N_3868,N_133,N_863);
and U3869 (N_3869,N_889,N_1626);
or U3870 (N_3870,N_944,N_775);
or U3871 (N_3871,N_1231,N_1914);
nand U3872 (N_3872,N_1166,N_816);
nand U3873 (N_3873,N_842,N_139);
or U3874 (N_3874,N_14,N_880);
or U3875 (N_3875,N_1603,N_1374);
nand U3876 (N_3876,N_1947,N_1809);
and U3877 (N_3877,N_79,N_351);
and U3878 (N_3878,N_1283,N_1110);
and U3879 (N_3879,N_1599,N_844);
nor U3880 (N_3880,N_1232,N_760);
nor U3881 (N_3881,N_1563,N_814);
nand U3882 (N_3882,N_1839,N_1537);
or U3883 (N_3883,N_1337,N_32);
and U3884 (N_3884,N_752,N_579);
xor U3885 (N_3885,N_1841,N_1216);
xnor U3886 (N_3886,N_588,N_475);
nand U3887 (N_3887,N_512,N_983);
and U3888 (N_3888,N_619,N_1621);
nor U3889 (N_3889,N_1022,N_1760);
or U3890 (N_3890,N_88,N_1828);
or U3891 (N_3891,N_432,N_1295);
and U3892 (N_3892,N_1135,N_960);
or U3893 (N_3893,N_1470,N_574);
or U3894 (N_3894,N_599,N_1213);
and U3895 (N_3895,N_1592,N_1560);
xor U3896 (N_3896,N_1138,N_486);
or U3897 (N_3897,N_1394,N_1150);
nand U3898 (N_3898,N_1966,N_299);
nor U3899 (N_3899,N_1596,N_782);
and U3900 (N_3900,N_661,N_1164);
and U3901 (N_3901,N_101,N_1732);
nor U3902 (N_3902,N_1076,N_681);
and U3903 (N_3903,N_1544,N_499);
and U3904 (N_3904,N_1283,N_984);
nand U3905 (N_3905,N_1102,N_1085);
or U3906 (N_3906,N_1177,N_1119);
or U3907 (N_3907,N_1735,N_1652);
nand U3908 (N_3908,N_262,N_1430);
nor U3909 (N_3909,N_1298,N_1788);
or U3910 (N_3910,N_961,N_745);
or U3911 (N_3911,N_32,N_1639);
or U3912 (N_3912,N_139,N_1387);
xnor U3913 (N_3913,N_863,N_1419);
or U3914 (N_3914,N_29,N_1744);
or U3915 (N_3915,N_830,N_948);
nor U3916 (N_3916,N_1933,N_1730);
xnor U3917 (N_3917,N_929,N_934);
nand U3918 (N_3918,N_555,N_977);
or U3919 (N_3919,N_23,N_149);
or U3920 (N_3920,N_1383,N_1370);
and U3921 (N_3921,N_417,N_1691);
or U3922 (N_3922,N_1910,N_570);
or U3923 (N_3923,N_346,N_1438);
or U3924 (N_3924,N_339,N_224);
nand U3925 (N_3925,N_57,N_944);
and U3926 (N_3926,N_31,N_1939);
and U3927 (N_3927,N_1793,N_1883);
nor U3928 (N_3928,N_44,N_1686);
nand U3929 (N_3929,N_1531,N_1375);
nor U3930 (N_3930,N_1677,N_1242);
nor U3931 (N_3931,N_121,N_1772);
nor U3932 (N_3932,N_787,N_1561);
and U3933 (N_3933,N_1985,N_1674);
and U3934 (N_3934,N_376,N_722);
and U3935 (N_3935,N_606,N_13);
nor U3936 (N_3936,N_512,N_1487);
or U3937 (N_3937,N_1217,N_1657);
and U3938 (N_3938,N_1135,N_1829);
nor U3939 (N_3939,N_895,N_755);
nand U3940 (N_3940,N_736,N_1065);
or U3941 (N_3941,N_1260,N_1919);
xnor U3942 (N_3942,N_236,N_39);
or U3943 (N_3943,N_736,N_207);
nor U3944 (N_3944,N_1488,N_1524);
nor U3945 (N_3945,N_985,N_450);
nand U3946 (N_3946,N_767,N_1830);
nand U3947 (N_3947,N_781,N_544);
or U3948 (N_3948,N_1914,N_500);
or U3949 (N_3949,N_106,N_595);
nand U3950 (N_3950,N_370,N_869);
and U3951 (N_3951,N_1024,N_463);
nand U3952 (N_3952,N_1822,N_819);
or U3953 (N_3953,N_1695,N_1916);
xnor U3954 (N_3954,N_157,N_243);
xnor U3955 (N_3955,N_1903,N_866);
or U3956 (N_3956,N_1814,N_1623);
and U3957 (N_3957,N_345,N_1937);
or U3958 (N_3958,N_786,N_254);
or U3959 (N_3959,N_429,N_1611);
nor U3960 (N_3960,N_1028,N_1639);
nor U3961 (N_3961,N_813,N_1651);
nor U3962 (N_3962,N_1073,N_1772);
and U3963 (N_3963,N_958,N_1685);
nand U3964 (N_3964,N_789,N_1470);
nand U3965 (N_3965,N_1659,N_1398);
and U3966 (N_3966,N_1671,N_795);
nor U3967 (N_3967,N_1584,N_295);
and U3968 (N_3968,N_1879,N_1901);
or U3969 (N_3969,N_1617,N_360);
nand U3970 (N_3970,N_1432,N_444);
or U3971 (N_3971,N_1019,N_291);
or U3972 (N_3972,N_1225,N_1497);
or U3973 (N_3973,N_1755,N_701);
and U3974 (N_3974,N_152,N_1639);
nand U3975 (N_3975,N_1877,N_969);
nand U3976 (N_3976,N_1872,N_1174);
and U3977 (N_3977,N_1288,N_348);
nand U3978 (N_3978,N_776,N_1723);
nor U3979 (N_3979,N_1189,N_1947);
or U3980 (N_3980,N_163,N_1742);
and U3981 (N_3981,N_757,N_992);
nand U3982 (N_3982,N_877,N_333);
or U3983 (N_3983,N_1205,N_1657);
nand U3984 (N_3984,N_793,N_280);
or U3985 (N_3985,N_224,N_64);
xnor U3986 (N_3986,N_518,N_600);
and U3987 (N_3987,N_835,N_419);
xor U3988 (N_3988,N_1818,N_1318);
and U3989 (N_3989,N_595,N_1395);
nor U3990 (N_3990,N_215,N_377);
and U3991 (N_3991,N_13,N_1669);
nor U3992 (N_3992,N_545,N_404);
nor U3993 (N_3993,N_666,N_1072);
nor U3994 (N_3994,N_1848,N_1606);
and U3995 (N_3995,N_685,N_822);
nand U3996 (N_3996,N_1149,N_223);
and U3997 (N_3997,N_456,N_735);
nand U3998 (N_3998,N_498,N_787);
nand U3999 (N_3999,N_1153,N_470);
and U4000 (N_4000,N_3833,N_3506);
nand U4001 (N_4001,N_3403,N_3661);
and U4002 (N_4002,N_2399,N_2927);
nand U4003 (N_4003,N_3832,N_2631);
and U4004 (N_4004,N_2165,N_3110);
nor U4005 (N_4005,N_3617,N_2202);
or U4006 (N_4006,N_2650,N_3858);
nor U4007 (N_4007,N_2586,N_3412);
or U4008 (N_4008,N_2201,N_2323);
or U4009 (N_4009,N_3411,N_3247);
and U4010 (N_4010,N_3364,N_3990);
nor U4011 (N_4011,N_3086,N_3480);
xnor U4012 (N_4012,N_2815,N_3509);
or U4013 (N_4013,N_2733,N_3267);
or U4014 (N_4014,N_3492,N_3393);
and U4015 (N_4015,N_3375,N_3866);
and U4016 (N_4016,N_3437,N_2732);
nor U4017 (N_4017,N_2736,N_3056);
and U4018 (N_4018,N_2960,N_3141);
nand U4019 (N_4019,N_3225,N_2488);
or U4020 (N_4020,N_3652,N_3494);
nand U4021 (N_4021,N_2497,N_2729);
or U4022 (N_4022,N_3200,N_3031);
nor U4023 (N_4023,N_3326,N_2826);
and U4024 (N_4024,N_2671,N_2577);
and U4025 (N_4025,N_3486,N_2528);
or U4026 (N_4026,N_3242,N_2821);
nand U4027 (N_4027,N_2331,N_2299);
and U4028 (N_4028,N_2391,N_3429);
or U4029 (N_4029,N_2524,N_3721);
or U4030 (N_4030,N_2773,N_2931);
xor U4031 (N_4031,N_3266,N_2963);
or U4032 (N_4032,N_2914,N_2805);
nor U4033 (N_4033,N_3102,N_2980);
nand U4034 (N_4034,N_2272,N_2315);
or U4035 (N_4035,N_3515,N_2120);
and U4036 (N_4036,N_3954,N_3557);
or U4037 (N_4037,N_2382,N_2464);
nor U4038 (N_4038,N_3419,N_2264);
nor U4039 (N_4039,N_2039,N_3612);
and U4040 (N_4040,N_3005,N_3907);
nor U4041 (N_4041,N_3383,N_3132);
nor U4042 (N_4042,N_2471,N_2626);
nor U4043 (N_4043,N_3618,N_2988);
nor U4044 (N_4044,N_3452,N_2329);
nand U4045 (N_4045,N_2769,N_3381);
or U4046 (N_4046,N_3867,N_2747);
or U4047 (N_4047,N_2590,N_3021);
nand U4048 (N_4048,N_3626,N_2661);
or U4049 (N_4049,N_2993,N_3294);
or U4050 (N_4050,N_3896,N_3302);
nor U4051 (N_4051,N_3666,N_2684);
and U4052 (N_4052,N_3569,N_2418);
and U4053 (N_4053,N_2564,N_2069);
and U4054 (N_4054,N_3087,N_3959);
nor U4055 (N_4055,N_3685,N_2830);
and U4056 (N_4056,N_2891,N_3507);
nor U4057 (N_4057,N_3933,N_2699);
and U4058 (N_4058,N_2047,N_2258);
nor U4059 (N_4059,N_3669,N_3877);
nand U4060 (N_4060,N_2324,N_2808);
and U4061 (N_4061,N_2137,N_2919);
or U4062 (N_4062,N_3085,N_2900);
and U4063 (N_4063,N_3045,N_2597);
or U4064 (N_4064,N_3170,N_3344);
or U4065 (N_4065,N_3033,N_2036);
or U4066 (N_4066,N_3694,N_2726);
and U4067 (N_4067,N_2390,N_2744);
and U4068 (N_4068,N_3746,N_3373);
and U4069 (N_4069,N_2345,N_3377);
and U4070 (N_4070,N_3939,N_3516);
or U4071 (N_4071,N_3036,N_2628);
nor U4072 (N_4072,N_3614,N_3476);
nor U4073 (N_4073,N_2281,N_2761);
and U4074 (N_4074,N_3121,N_3065);
nor U4075 (N_4075,N_3236,N_2740);
nor U4076 (N_4076,N_3823,N_2774);
nand U4077 (N_4077,N_3317,N_3495);
and U4078 (N_4078,N_3001,N_3589);
and U4079 (N_4079,N_2354,N_2175);
nand U4080 (N_4080,N_2063,N_2673);
nand U4081 (N_4081,N_2288,N_2799);
nor U4082 (N_4082,N_2298,N_2909);
nor U4083 (N_4083,N_3020,N_2804);
nor U4084 (N_4084,N_2300,N_3642);
nand U4085 (N_4085,N_2516,N_2833);
nor U4086 (N_4086,N_3223,N_3425);
and U4087 (N_4087,N_2782,N_3625);
and U4088 (N_4088,N_3578,N_2886);
xor U4089 (N_4089,N_2797,N_3632);
or U4090 (N_4090,N_3927,N_2320);
nand U4091 (N_4091,N_2430,N_3489);
nand U4092 (N_4092,N_3248,N_3016);
and U4093 (N_4093,N_2468,N_2579);
nor U4094 (N_4094,N_3865,N_3211);
or U4095 (N_4095,N_3988,N_2713);
nand U4096 (N_4096,N_2049,N_2776);
nor U4097 (N_4097,N_3035,N_2177);
and U4098 (N_4098,N_3991,N_2231);
and U4099 (N_4099,N_2241,N_3719);
or U4100 (N_4100,N_3816,N_3011);
nand U4101 (N_4101,N_3303,N_2601);
and U4102 (N_4102,N_2618,N_2883);
nand U4103 (N_4103,N_3118,N_2584);
nor U4104 (N_4104,N_3128,N_3930);
nor U4105 (N_4105,N_2238,N_2448);
and U4106 (N_4106,N_3052,N_2071);
or U4107 (N_4107,N_3924,N_3096);
nor U4108 (N_4108,N_2563,N_2690);
and U4109 (N_4109,N_3705,N_2373);
or U4110 (N_4110,N_3722,N_3095);
nand U4111 (N_4111,N_3590,N_3504);
and U4112 (N_4112,N_2494,N_2734);
and U4113 (N_4113,N_2982,N_2932);
and U4114 (N_4114,N_3050,N_2630);
or U4115 (N_4115,N_3280,N_3708);
or U4116 (N_4116,N_3586,N_2881);
or U4117 (N_4117,N_2917,N_2949);
nor U4118 (N_4118,N_3799,N_3432);
or U4119 (N_4119,N_2170,N_2279);
nor U4120 (N_4120,N_3842,N_2944);
or U4121 (N_4121,N_3921,N_2540);
nor U4122 (N_4122,N_2283,N_2921);
nand U4123 (N_4123,N_2542,N_2719);
nor U4124 (N_4124,N_3100,N_3973);
or U4125 (N_4125,N_2578,N_2495);
nand U4126 (N_4126,N_3461,N_2169);
nand U4127 (N_4127,N_2306,N_2290);
nand U4128 (N_4128,N_3581,N_3026);
nand U4129 (N_4129,N_2447,N_2603);
nand U4130 (N_4130,N_3671,N_3931);
and U4131 (N_4131,N_2951,N_2152);
nor U4132 (N_4132,N_2655,N_2820);
nor U4133 (N_4133,N_3374,N_2029);
or U4134 (N_4134,N_3341,N_3623);
or U4135 (N_4135,N_2191,N_2543);
or U4136 (N_4136,N_3658,N_2217);
and U4137 (N_4137,N_3598,N_2180);
nand U4138 (N_4138,N_3464,N_2859);
nor U4139 (N_4139,N_3633,N_2860);
or U4140 (N_4140,N_3218,N_3090);
or U4141 (N_4141,N_2537,N_2515);
nand U4142 (N_4142,N_3354,N_2666);
or U4143 (N_4143,N_3868,N_2259);
nor U4144 (N_4144,N_2520,N_3295);
or U4145 (N_4145,N_2487,N_3079);
nand U4146 (N_4146,N_2562,N_2714);
or U4147 (N_4147,N_3171,N_2941);
nor U4148 (N_4148,N_2853,N_3693);
nor U4149 (N_4149,N_2884,N_3998);
or U4150 (N_4150,N_2222,N_3160);
nor U4151 (N_4151,N_2293,N_2888);
nand U4152 (N_4152,N_2307,N_3822);
nand U4153 (N_4153,N_3336,N_2212);
or U4154 (N_4154,N_3664,N_2312);
nand U4155 (N_4155,N_3308,N_2095);
and U4156 (N_4156,N_3539,N_2897);
or U4157 (N_4157,N_3217,N_2636);
nand U4158 (N_4158,N_2512,N_2925);
nor U4159 (N_4159,N_2576,N_2055);
nand U4160 (N_4160,N_2768,N_2359);
nor U4161 (N_4161,N_2702,N_3893);
nor U4162 (N_4162,N_3695,N_2803);
or U4163 (N_4163,N_2349,N_3212);
or U4164 (N_4164,N_2139,N_3980);
or U4165 (N_4165,N_3238,N_2013);
nand U4166 (N_4166,N_3108,N_3596);
nand U4167 (N_4167,N_3156,N_2529);
nor U4168 (N_4168,N_3335,N_3207);
nand U4169 (N_4169,N_2214,N_2841);
and U4170 (N_4170,N_2068,N_3416);
nand U4171 (N_4171,N_3152,N_2829);
or U4172 (N_4172,N_3150,N_3301);
or U4173 (N_4173,N_3653,N_3901);
or U4174 (N_4174,N_3176,N_2580);
nor U4175 (N_4175,N_3819,N_3526);
nand U4176 (N_4176,N_3811,N_3628);
nand U4177 (N_4177,N_2566,N_3024);
nor U4178 (N_4178,N_3583,N_2026);
nor U4179 (N_4179,N_3550,N_2270);
nand U4180 (N_4180,N_2381,N_3448);
nor U4181 (N_4181,N_2425,N_3760);
xor U4182 (N_4182,N_3709,N_2374);
nand U4183 (N_4183,N_2965,N_2970);
nand U4184 (N_4184,N_3874,N_3870);
nor U4185 (N_4185,N_2412,N_2966);
and U4186 (N_4186,N_3838,N_2454);
or U4187 (N_4187,N_2544,N_3735);
and U4188 (N_4188,N_2715,N_2637);
nor U4189 (N_4189,N_3305,N_2445);
nor U4190 (N_4190,N_2764,N_2301);
and U4191 (N_4191,N_2469,N_2278);
nand U4192 (N_4192,N_3343,N_3478);
nor U4193 (N_4193,N_3491,N_2717);
and U4194 (N_4194,N_3820,N_3183);
nor U4195 (N_4195,N_3275,N_3967);
nand U4196 (N_4196,N_3027,N_3668);
nand U4197 (N_4197,N_3051,N_3208);
or U4198 (N_4198,N_3906,N_3213);
and U4199 (N_4199,N_2898,N_3109);
nor U4200 (N_4200,N_2878,N_3396);
nor U4201 (N_4201,N_2405,N_2422);
and U4202 (N_4202,N_2784,N_3792);
or U4203 (N_4203,N_2854,N_3349);
nand U4204 (N_4204,N_3384,N_3477);
nand U4205 (N_4205,N_3070,N_2882);
or U4206 (N_4206,N_3852,N_3358);
nand U4207 (N_4207,N_3046,N_3787);
nor U4208 (N_4208,N_3240,N_2572);
or U4209 (N_4209,N_2148,N_3388);
nand U4210 (N_4210,N_2535,N_2971);
nand U4211 (N_4211,N_2824,N_3075);
nor U4212 (N_4212,N_2844,N_3984);
nor U4213 (N_4213,N_3941,N_2800);
or U4214 (N_4214,N_2151,N_3631);
xnor U4215 (N_4215,N_3235,N_3264);
nor U4216 (N_4216,N_2989,N_3957);
or U4217 (N_4217,N_3184,N_3844);
nor U4218 (N_4218,N_3473,N_2130);
and U4219 (N_4219,N_2123,N_3487);
nor U4220 (N_4220,N_3450,N_2073);
nand U4221 (N_4221,N_3646,N_2956);
nand U4222 (N_4222,N_3788,N_3985);
nand U4223 (N_4223,N_2632,N_2649);
nor U4224 (N_4224,N_2806,N_2114);
or U4225 (N_4225,N_3995,N_3689);
and U4226 (N_4226,N_3513,N_2718);
nand U4227 (N_4227,N_2765,N_3078);
xnor U4228 (N_4228,N_3688,N_2081);
nor U4229 (N_4229,N_3201,N_2340);
and U4230 (N_4230,N_3511,N_3701);
nand U4231 (N_4231,N_3284,N_2505);
nand U4232 (N_4232,N_2807,N_2369);
and U4233 (N_4233,N_2195,N_2858);
nor U4234 (N_4234,N_2140,N_2097);
and U4235 (N_4235,N_3363,N_2362);
nand U4236 (N_4236,N_3112,N_3433);
or U4237 (N_4237,N_3334,N_3361);
and U4238 (N_4238,N_3770,N_2001);
or U4239 (N_4239,N_2035,N_2093);
nor U4240 (N_4240,N_3360,N_3185);
nor U4241 (N_4241,N_2924,N_3714);
nor U4242 (N_4242,N_3179,N_3214);
nor U4243 (N_4243,N_2530,N_2823);
or U4244 (N_4244,N_3889,N_2334);
or U4245 (N_4245,N_3910,N_2875);
nor U4246 (N_4246,N_2675,N_2048);
nand U4247 (N_4247,N_3791,N_3287);
nor U4248 (N_4248,N_2504,N_3420);
nand U4249 (N_4249,N_2861,N_2203);
nand U4250 (N_4250,N_3474,N_2478);
xnor U4251 (N_4251,N_2078,N_3863);
nor U4252 (N_4252,N_3042,N_3565);
nand U4253 (N_4253,N_2190,N_3699);
nor U4254 (N_4254,N_2781,N_2969);
or U4255 (N_4255,N_3622,N_3271);
nor U4256 (N_4256,N_2134,N_2427);
nor U4257 (N_4257,N_3890,N_2146);
or U4258 (N_4258,N_2538,N_3062);
or U4259 (N_4259,N_2604,N_2701);
and U4260 (N_4260,N_3814,N_2770);
and U4261 (N_4261,N_2356,N_3736);
or U4262 (N_4262,N_2674,N_2045);
nor U4263 (N_4263,N_3470,N_3008);
nor U4264 (N_4264,N_3857,N_2363);
nor U4265 (N_4265,N_3879,N_2635);
nor U4266 (N_4266,N_2365,N_3643);
nor U4267 (N_4267,N_2102,N_2556);
nor U4268 (N_4268,N_3327,N_2871);
and U4269 (N_4269,N_3014,N_2974);
nor U4270 (N_4270,N_2113,N_3728);
and U4271 (N_4271,N_2500,N_3840);
nand U4272 (N_4272,N_2263,N_2218);
or U4273 (N_4273,N_2642,N_2163);
or U4274 (N_4274,N_2547,N_3165);
nor U4275 (N_4275,N_3398,N_2756);
and U4276 (N_4276,N_2711,N_2694);
nor U4277 (N_4277,N_3724,N_3665);
or U4278 (N_4278,N_3274,N_3366);
or U4279 (N_4279,N_3734,N_3672);
nand U4280 (N_4280,N_3945,N_3925);
xor U4281 (N_4281,N_3825,N_3543);
or U4282 (N_4282,N_2759,N_3488);
nor U4283 (N_4283,N_2825,N_3257);
nor U4284 (N_4284,N_3084,N_3723);
nand U4285 (N_4285,N_3754,N_2125);
nand U4286 (N_4286,N_2678,N_3902);
nor U4287 (N_4287,N_2171,N_3594);
nand U4288 (N_4288,N_3338,N_3517);
or U4289 (N_4289,N_3315,N_3683);
and U4290 (N_4290,N_3936,N_3580);
nand U4291 (N_4291,N_2533,N_3356);
and U4292 (N_4292,N_3193,N_2025);
nand U4293 (N_4293,N_2271,N_3029);
or U4294 (N_4294,N_2051,N_2470);
nor U4295 (N_4295,N_3177,N_2183);
nand U4296 (N_4296,N_2004,N_3993);
nand U4297 (N_4297,N_2607,N_3399);
nand U4298 (N_4298,N_2745,N_2229);
nor U4299 (N_4299,N_3861,N_2157);
and U4300 (N_4300,N_3169,N_2907);
or U4301 (N_4301,N_3704,N_2930);
and U4302 (N_4302,N_2124,N_3233);
nand U4303 (N_4303,N_3055,N_2978);
or U4304 (N_4304,N_3106,N_3752);
or U4305 (N_4305,N_2997,N_2173);
nand U4306 (N_4306,N_3424,N_2091);
or U4307 (N_4307,N_3376,N_2582);
and U4308 (N_4308,N_3122,N_3831);
nor U4309 (N_4309,N_3808,N_3706);
nor U4310 (N_4310,N_2789,N_2905);
nor U4311 (N_4311,N_3094,N_2952);
nor U4312 (N_4312,N_3892,N_3219);
and U4313 (N_4313,N_3932,N_3717);
or U4314 (N_4314,N_3940,N_2786);
nor U4315 (N_4315,N_2459,N_2379);
or U4316 (N_4316,N_3154,N_2467);
nor U4317 (N_4317,N_2274,N_2431);
nand U4318 (N_4318,N_3687,N_2233);
or U4319 (N_4319,N_3234,N_3944);
or U4320 (N_4320,N_2981,N_2156);
and U4321 (N_4321,N_2172,N_2778);
nor U4322 (N_4322,N_2458,N_3009);
or U4323 (N_4323,N_2519,N_3764);
and U4324 (N_4324,N_2780,N_2939);
nand U4325 (N_4325,N_2126,N_2251);
or U4326 (N_4326,N_3853,N_3611);
nor U4327 (N_4327,N_3057,N_3149);
xor U4328 (N_4328,N_2292,N_2903);
nand U4329 (N_4329,N_3362,N_3216);
nor U4330 (N_4330,N_3255,N_3083);
or U4331 (N_4331,N_2273,N_2634);
or U4332 (N_4332,N_3455,N_2041);
and U4333 (N_4333,N_2444,N_3883);
or U4334 (N_4334,N_3410,N_2602);
nor U4335 (N_4335,N_3732,N_3987);
and U4336 (N_4336,N_2145,N_3028);
nand U4337 (N_4337,N_2794,N_2498);
or U4338 (N_4338,N_2936,N_3847);
nand U4339 (N_4339,N_2044,N_3283);
nor U4340 (N_4340,N_2600,N_2613);
or U4341 (N_4341,N_3544,N_2567);
nor U4342 (N_4342,N_3430,N_2685);
and U4343 (N_4343,N_3250,N_3147);
and U4344 (N_4344,N_3649,N_2249);
nor U4345 (N_4345,N_2926,N_3192);
nor U4346 (N_4346,N_3813,N_3597);
nand U4347 (N_4347,N_3585,N_3684);
nor U4348 (N_4348,N_2252,N_2648);
or U4349 (N_4349,N_3204,N_3786);
or U4350 (N_4350,N_2902,N_2302);
nor U4351 (N_4351,N_2625,N_2842);
or U4352 (N_4352,N_2698,N_3568);
nand U4353 (N_4353,N_2593,N_2216);
or U4354 (N_4354,N_3347,N_3224);
and U4355 (N_4355,N_3835,N_2096);
xnor U4356 (N_4356,N_3807,N_2333);
nor U4357 (N_4357,N_3215,N_2378);
or U4358 (N_4358,N_2309,N_3809);
nand U4359 (N_4359,N_2940,N_3675);
nor U4360 (N_4360,N_3548,N_2380);
nand U4361 (N_4361,N_2182,N_3686);
or U4362 (N_4362,N_3750,N_3174);
nand U4363 (N_4363,N_2289,N_2449);
nor U4364 (N_4364,N_2228,N_3908);
or U4365 (N_4365,N_3414,N_2511);
nor U4366 (N_4366,N_3928,N_2121);
or U4367 (N_4367,N_2060,N_2099);
or U4368 (N_4368,N_2708,N_2396);
or U4369 (N_4369,N_2973,N_2938);
nor U4370 (N_4370,N_3560,N_2811);
nand U4371 (N_4371,N_2551,N_3960);
and U4372 (N_4372,N_3292,N_3917);
nor U4373 (N_4373,N_3202,N_3116);
nor U4374 (N_4374,N_2461,N_2539);
xnor U4375 (N_4375,N_2680,N_2667);
nand U4376 (N_4376,N_3210,N_2366);
nor U4377 (N_4377,N_3875,N_2042);
nand U4378 (N_4378,N_3634,N_3145);
or U4379 (N_4379,N_2052,N_2583);
nand U4380 (N_4380,N_3641,N_3573);
nand U4381 (N_4381,N_2703,N_3905);
xor U4382 (N_4382,N_2338,N_3876);
and U4383 (N_4383,N_3880,N_3558);
or U4384 (N_4384,N_3860,N_3089);
or U4385 (N_4385,N_2235,N_3781);
or U4386 (N_4386,N_2462,N_3196);
or U4387 (N_4387,N_3309,N_2611);
nor U4388 (N_4388,N_2640,N_3319);
or U4389 (N_4389,N_2599,N_2452);
and U4390 (N_4390,N_3365,N_2856);
nand U4391 (N_4391,N_3926,N_3447);
or U4392 (N_4392,N_2456,N_2007);
nor U4393 (N_4393,N_2596,N_2850);
nand U4394 (N_4394,N_3038,N_3310);
nor U4395 (N_4395,N_2420,N_2392);
nor U4396 (N_4396,N_2809,N_3333);
xor U4397 (N_4397,N_2994,N_2879);
nand U4398 (N_4398,N_3244,N_3804);
and U4399 (N_4399,N_2508,N_3584);
nand U4400 (N_4400,N_3797,N_3350);
nor U4401 (N_4401,N_2406,N_2463);
nor U4402 (N_4402,N_3790,N_2594);
nor U4403 (N_4403,N_2348,N_3012);
nand U4404 (N_4404,N_2686,N_3126);
nand U4405 (N_4405,N_2296,N_2387);
or U4406 (N_4406,N_2408,N_2466);
nor U4407 (N_4407,N_3453,N_3140);
nor U4408 (N_4408,N_3826,N_3041);
and U4409 (N_4409,N_2737,N_3537);
nor U4410 (N_4410,N_2168,N_3405);
and U4411 (N_4411,N_3670,N_3348);
nand U4412 (N_4412,N_3776,N_3794);
and U4413 (N_4413,N_2090,N_2061);
nor U4414 (N_4414,N_3189,N_2915);
nand U4415 (N_4415,N_3800,N_3963);
nand U4416 (N_4416,N_2706,N_3745);
nor U4417 (N_4417,N_2245,N_2083);
nor U4418 (N_4418,N_3340,N_3953);
or U4419 (N_4419,N_3994,N_2864);
nor U4420 (N_4420,N_2972,N_2793);
nor U4421 (N_4421,N_2442,N_3166);
nor U4422 (N_4422,N_3703,N_3976);
nor U4423 (N_4423,N_3965,N_3692);
nor U4424 (N_4424,N_2654,N_2766);
nand U4425 (N_4425,N_2242,N_3961);
or U4426 (N_4426,N_3167,N_2199);
and U4427 (N_4427,N_2038,N_2336);
or U4428 (N_4428,N_2394,N_3519);
nor U4429 (N_4429,N_2877,N_2870);
or U4430 (N_4430,N_2481,N_2246);
and U4431 (N_4431,N_3390,N_3047);
nand U4432 (N_4432,N_3369,N_2187);
nand U4433 (N_4433,N_3682,N_2008);
or U4434 (N_4434,N_2370,N_3277);
and U4435 (N_4435,N_2890,N_2922);
or U4436 (N_4436,N_3259,N_2018);
nor U4437 (N_4437,N_2403,N_3113);
or U4438 (N_4438,N_2028,N_3923);
nand U4439 (N_4439,N_3730,N_3739);
nor U4440 (N_4440,N_3601,N_2371);
or U4441 (N_4441,N_2906,N_2436);
nor U4442 (N_4442,N_2499,N_3602);
or U4443 (N_4443,N_2419,N_2265);
xor U4444 (N_4444,N_3720,N_2257);
and U4445 (N_4445,N_2200,N_2484);
and U4446 (N_4446,N_3575,N_3949);
or U4447 (N_4447,N_2196,N_2904);
nor U4448 (N_4448,N_3552,N_2122);
and U4449 (N_4449,N_2958,N_3093);
xor U4450 (N_4450,N_3273,N_3357);
or U4451 (N_4451,N_3966,N_2928);
nand U4452 (N_4452,N_3468,N_3843);
nand U4453 (N_4453,N_3712,N_3608);
nand U4454 (N_4454,N_2771,N_2372);
or U4455 (N_4455,N_3391,N_3158);
nor U4456 (N_4456,N_3541,N_3559);
and U4457 (N_4457,N_2709,N_2020);
and U4458 (N_4458,N_3269,N_2284);
or U4459 (N_4459,N_3496,N_3332);
nor U4460 (N_4460,N_2536,N_3836);
nand U4461 (N_4461,N_2046,N_2389);
nand U4462 (N_4462,N_2087,N_2351);
nor U4463 (N_4463,N_2098,N_3784);
and U4464 (N_4464,N_2950,N_3545);
or U4465 (N_4465,N_3845,N_2388);
nand U4466 (N_4466,N_2852,N_3636);
or U4467 (N_4467,N_2943,N_2477);
and U4468 (N_4468,N_3119,N_3593);
or U4469 (N_4469,N_2691,N_2094);
and U4470 (N_4470,N_2992,N_3900);
nor U4471 (N_4471,N_2076,N_2064);
nand U4472 (N_4472,N_3522,N_2953);
and U4473 (N_4473,N_3131,N_2656);
nand U4474 (N_4474,N_3520,N_2085);
nor U4475 (N_4475,N_3493,N_3841);
and U4476 (N_4476,N_3740,N_3574);
or U4477 (N_4477,N_2082,N_3479);
xor U4478 (N_4478,N_2801,N_3293);
or U4479 (N_4479,N_3025,N_2266);
or U4480 (N_4480,N_2189,N_2268);
and U4481 (N_4481,N_3549,N_2983);
and U4482 (N_4482,N_2166,N_2440);
nand U4483 (N_4483,N_2617,N_3197);
and U4484 (N_4484,N_2946,N_3426);
or U4485 (N_4485,N_3785,N_3107);
nand U4486 (N_4486,N_2798,N_2568);
nand U4487 (N_4487,N_2553,N_2619);
or U4488 (N_4488,N_2731,N_2043);
or U4489 (N_4489,N_3251,N_3818);
and U4490 (N_4490,N_3570,N_2310);
nand U4491 (N_4491,N_3318,N_3422);
nor U4492 (N_4492,N_2460,N_2627);
or U4493 (N_4493,N_3345,N_2426);
and U4494 (N_4494,N_2465,N_2104);
and U4495 (N_4495,N_3645,N_2814);
and U4496 (N_4496,N_3178,N_3935);
or U4497 (N_4497,N_3471,N_3439);
nor U4498 (N_4498,N_3249,N_2569);
xnor U4499 (N_4499,N_2605,N_3762);
xor U4500 (N_4500,N_3263,N_2155);
nand U4501 (N_4501,N_3591,N_3180);
nor U4502 (N_4502,N_3015,N_3465);
or U4503 (N_4503,N_3501,N_3142);
and U4504 (N_4504,N_3049,N_2006);
xnor U4505 (N_4505,N_2342,N_2070);
nand U4506 (N_4506,N_3472,N_2506);
and U4507 (N_4507,N_2239,N_2574);
nor U4508 (N_4508,N_3871,N_2862);
or U4509 (N_4509,N_2210,N_2984);
and U4510 (N_4510,N_2521,N_3904);
nand U4511 (N_4511,N_2688,N_2510);
nand U4512 (N_4512,N_3182,N_2414);
nand U4513 (N_4513,N_3624,N_3992);
nand U4514 (N_4514,N_2434,N_2643);
nand U4515 (N_4515,N_3700,N_2400);
nand U4516 (N_4516,N_2110,N_2062);
nand U4517 (N_4517,N_3938,N_3518);
and U4518 (N_4518,N_3629,N_2021);
and U4519 (N_4519,N_3555,N_3291);
nor U4520 (N_4520,N_2722,N_2552);
nand U4521 (N_4521,N_3530,N_3322);
and U4522 (N_4522,N_2050,N_3698);
xnor U4523 (N_4523,N_3187,N_3418);
or U4524 (N_4524,N_3483,N_2480);
nand U4525 (N_4525,N_3503,N_3285);
or U4526 (N_4526,N_3314,N_2092);
nor U4527 (N_4527,N_2610,N_3894);
nor U4528 (N_4528,N_2260,N_2479);
nor U4529 (N_4529,N_3307,N_2541);
or U4530 (N_4530,N_3229,N_3000);
nor U4531 (N_4531,N_2705,N_3253);
nor U4532 (N_4532,N_2103,N_2154);
nor U4533 (N_4533,N_2423,N_3017);
or U4534 (N_4534,N_3856,N_2409);
or U4535 (N_4535,N_2220,N_2916);
and U4536 (N_4536,N_3442,N_2303);
nor U4537 (N_4537,N_2913,N_2023);
or U4538 (N_4538,N_3986,N_2570);
nand U4539 (N_4539,N_3497,N_3386);
nor U4540 (N_4540,N_3330,N_2346);
nand U4541 (N_4541,N_2855,N_2030);
or U4542 (N_4542,N_2294,N_3796);
or U4543 (N_4543,N_3312,N_2995);
or U4544 (N_4544,N_2325,N_2127);
nand U4545 (N_4545,N_2428,N_2571);
nor U4546 (N_4546,N_2660,N_2056);
and U4547 (N_4547,N_3531,N_2355);
nand U4548 (N_4548,N_2933,N_2188);
and U4549 (N_4549,N_3245,N_2697);
nand U4550 (N_4550,N_2308,N_3916);
nor U4551 (N_4551,N_2827,N_3427);
and U4552 (N_4552,N_3532,N_2194);
or U4553 (N_4553,N_3756,N_3789);
or U4554 (N_4554,N_2818,N_2838);
nand U4555 (N_4555,N_2313,N_3114);
or U4556 (N_4556,N_2244,N_3929);
nor U4557 (N_4557,N_3321,N_2153);
and U4558 (N_4558,N_3098,N_3408);
or U4559 (N_4559,N_3716,N_2591);
nand U4560 (N_4560,N_3621,N_2136);
nand U4561 (N_4561,N_3895,N_3690);
and U4562 (N_4562,N_2384,N_3230);
and U4563 (N_4563,N_2311,N_3656);
or U4564 (N_4564,N_3485,N_3638);
or U4565 (N_4565,N_3793,N_3869);
and U4566 (N_4566,N_3677,N_3097);
and U4567 (N_4567,N_3246,N_3778);
or U4568 (N_4568,N_3252,N_2573);
or U4569 (N_4569,N_2176,N_2053);
and U4570 (N_4570,N_2402,N_2910);
or U4571 (N_4571,N_3974,N_2866);
and U4572 (N_4572,N_3592,N_2185);
nor U4573 (N_4573,N_2534,N_3385);
or U4574 (N_4574,N_2084,N_3449);
nand U4575 (N_4575,N_2261,N_2158);
and U4576 (N_4576,N_2286,N_2977);
nor U4577 (N_4577,N_3821,N_2262);
nor U4578 (N_4578,N_2672,N_3782);
or U4579 (N_4579,N_2011,N_3738);
or U4580 (N_4580,N_3130,N_3872);
xor U4581 (N_4581,N_2150,N_2695);
and U4582 (N_4582,N_3605,N_3220);
and U4583 (N_4583,N_2646,N_2383);
nand U4584 (N_4584,N_3859,N_2851);
nor U4585 (N_4585,N_3286,N_3538);
or U4586 (N_4586,N_3616,N_3395);
and U4587 (N_4587,N_2790,N_3337);
nor U4588 (N_4588,N_3101,N_3711);
nand U4589 (N_4589,N_3535,N_2142);
and U4590 (N_4590,N_3175,N_3798);
nand U4591 (N_4591,N_2357,N_2234);
nand U4592 (N_4592,N_3839,N_3136);
nor U4593 (N_4593,N_2657,N_3221);
nand U4594 (N_4594,N_2624,N_3898);
nor U4595 (N_4595,N_3678,N_2587);
and U4596 (N_4596,N_2753,N_3946);
nand U4597 (N_4597,N_2507,N_2638);
nor U4598 (N_4598,N_2285,N_3498);
nor U4599 (N_4599,N_2869,N_2561);
nand U4600 (N_4600,N_3968,N_3133);
nor U4601 (N_4601,N_2716,N_3371);
and U4602 (N_4602,N_3299,N_2280);
nand U4603 (N_4603,N_2446,N_2438);
nor U4604 (N_4604,N_2012,N_3757);
xor U4605 (N_4605,N_2339,N_2620);
or U4606 (N_4606,N_3667,N_3571);
or U4607 (N_4607,N_3887,N_2397);
nand U4608 (N_4608,N_3120,N_2100);
nor U4609 (N_4609,N_3815,N_3718);
nand U4610 (N_4610,N_3352,N_2295);
xnor U4611 (N_4611,N_3576,N_2645);
nand U4612 (N_4612,N_3002,N_3710);
nand U4613 (N_4613,N_3956,N_3368);
or U4614 (N_4614,N_2208,N_3209);
nand U4615 (N_4615,N_2230,N_2352);
nor U4616 (N_4616,N_2128,N_3702);
or U4617 (N_4617,N_2531,N_2920);
nand U4618 (N_4618,N_3969,N_2670);
and U4619 (N_4619,N_3650,N_2792);
or U4620 (N_4620,N_3378,N_2232);
or U4621 (N_4621,N_2948,N_2129);
xor U4622 (N_4622,N_3855,N_3268);
nor U4623 (N_4623,N_3725,N_2876);
or U4624 (N_4624,N_3256,N_2964);
or U4625 (N_4625,N_2040,N_3587);
and U4626 (N_4626,N_3076,N_3144);
nor U4627 (N_4627,N_2297,N_3884);
or U4628 (N_4628,N_2178,N_3775);
and U4629 (N_4629,N_2282,N_2682);
nor U4630 (N_4630,N_3074,N_2174);
or U4631 (N_4631,N_2887,N_3475);
nor U4632 (N_4632,N_3137,N_3276);
and U4633 (N_4633,N_2079,N_3032);
nor U4634 (N_4634,N_3502,N_2557);
or U4635 (N_4635,N_2704,N_3331);
and U4636 (N_4636,N_3289,N_2857);
and U4637 (N_4637,N_3726,N_3769);
nand U4638 (N_4638,N_3674,N_3655);
and U4639 (N_4639,N_2501,N_2664);
nand U4640 (N_4640,N_2621,N_2712);
nand U4641 (N_4641,N_2401,N_3713);
or U4642 (N_4642,N_3346,N_3691);
xor U4643 (N_4643,N_2589,N_2115);
nor U4644 (N_4644,N_3124,N_2696);
and U4645 (N_4645,N_3443,N_2318);
and U4646 (N_4646,N_3523,N_2132);
or U4647 (N_4647,N_2341,N_3022);
nand U4648 (N_4648,N_3060,N_2663);
or U4649 (N_4649,N_3588,N_3546);
or U4650 (N_4650,N_2817,N_2433);
xor U4651 (N_4651,N_3304,N_2754);
nor U4652 (N_4652,N_3606,N_2967);
nand U4653 (N_4653,N_2361,N_2548);
and U4654 (N_4654,N_2889,N_3771);
nor U4655 (N_4655,N_2138,N_3139);
nor U4656 (N_4656,N_2892,N_3802);
and U4657 (N_4657,N_3742,N_2668);
nand U4658 (N_4658,N_2911,N_3155);
or U4659 (N_4659,N_3068,N_3996);
or U4660 (N_4660,N_2019,N_3173);
nor U4661 (N_4661,N_3948,N_3972);
and U4662 (N_4662,N_3630,N_2893);
or U4663 (N_4663,N_2237,N_3500);
and U4664 (N_4664,N_2316,N_2874);
and U4665 (N_4665,N_2247,N_2681);
nand U4666 (N_4666,N_2559,N_2918);
nor U4667 (N_4667,N_3261,N_3380);
and U4668 (N_4668,N_3010,N_3510);
nand U4669 (N_4669,N_3663,N_2901);
and U4670 (N_4670,N_2912,N_2942);
and U4671 (N_4671,N_3635,N_2376);
and U4672 (N_4672,N_3370,N_2377);
and U4673 (N_4673,N_3505,N_3743);
nor U4674 (N_4674,N_2255,N_2022);
nand U4675 (N_4675,N_2608,N_2692);
nand U4676 (N_4676,N_3765,N_3599);
xor U4677 (N_4677,N_3647,N_2725);
nand U4678 (N_4678,N_3324,N_3862);
nand U4679 (N_4679,N_2161,N_3899);
or U4680 (N_4680,N_3463,N_3064);
nor U4681 (N_4681,N_3146,N_2837);
or U4682 (N_4682,N_2476,N_2088);
nor U4683 (N_4683,N_3950,N_2337);
nor U4684 (N_4684,N_2791,N_3850);
nand U4685 (N_4685,N_2863,N_2116);
or U4686 (N_4686,N_2819,N_2276);
nand U4687 (N_4687,N_2491,N_3059);
or U4688 (N_4688,N_3977,N_2908);
nand U4689 (N_4689,N_2211,N_2527);
or U4690 (N_4690,N_2606,N_2836);
xor U4691 (N_4691,N_2089,N_2206);
or U4692 (N_4692,N_2846,N_2828);
nor U4693 (N_4693,N_3129,N_2080);
and U4694 (N_4694,N_2344,N_2490);
nand U4695 (N_4695,N_2758,N_3763);
and U4696 (N_4696,N_2755,N_2204);
nor U4697 (N_4697,N_3044,N_3680);
or U4698 (N_4698,N_2482,N_3607);
nand U4699 (N_4699,N_2721,N_2750);
or U4700 (N_4700,N_3707,N_3143);
nor U4701 (N_4701,N_3897,N_3903);
nand U4702 (N_4702,N_3351,N_2133);
nand U4703 (N_4703,N_2895,N_3837);
nor U4704 (N_4704,N_2275,N_3556);
and U4705 (N_4705,N_3007,N_2330);
nand U4706 (N_4706,N_3159,N_2937);
or U4707 (N_4707,N_3003,N_3148);
and U4708 (N_4708,N_3508,N_3190);
nand U4709 (N_4709,N_2147,N_2439);
or U4710 (N_4710,N_2954,N_3610);
or U4711 (N_4711,N_3157,N_3077);
nand U4712 (N_4712,N_3227,N_2609);
and U4713 (N_4713,N_3812,N_2435);
nor U4714 (N_4714,N_2167,N_2353);
nor U4715 (N_4715,N_3536,N_2872);
nand U4716 (N_4716,N_3226,N_2945);
and U4717 (N_4717,N_2457,N_3296);
nand U4718 (N_4718,N_3529,N_2112);
or U4719 (N_4719,N_3013,N_2785);
nor U4720 (N_4720,N_3272,N_2739);
or U4721 (N_4721,N_2687,N_2549);
and U4722 (N_4722,N_2896,N_2957);
nor U4723 (N_4723,N_2291,N_3400);
and U4724 (N_4724,N_3441,N_2513);
or U4725 (N_4725,N_3563,N_3228);
or U4726 (N_4726,N_3848,N_2343);
or U4727 (N_4727,N_3423,N_3172);
nand U4728 (N_4728,N_2332,N_3080);
and U4729 (N_4729,N_2935,N_3397);
xnor U4730 (N_4730,N_3194,N_3777);
and U4731 (N_4731,N_2287,N_3943);
nand U4732 (N_4732,N_2653,N_2117);
and U4733 (N_4733,N_2525,N_2652);
nand U4734 (N_4734,N_2135,N_2417);
nor U4735 (N_4735,N_2748,N_3533);
nor U4736 (N_4736,N_2990,N_2727);
nor U4737 (N_4737,N_2424,N_2746);
and U4738 (N_4738,N_2033,N_3458);
and U4739 (N_4739,N_2350,N_2243);
nand U4740 (N_4740,N_3955,N_3191);
nor U4741 (N_4741,N_3199,N_3195);
or U4742 (N_4742,N_2248,N_3846);
nor U4743 (N_4743,N_2075,N_2735);
nor U4744 (N_4744,N_3751,N_3952);
and U4745 (N_4745,N_3091,N_2059);
nand U4746 (N_4746,N_2867,N_2304);
or U4747 (N_4747,N_2588,N_2658);
nor U4748 (N_4748,N_3482,N_2847);
nand U4749 (N_4749,N_3824,N_3744);
nor U4750 (N_4750,N_3749,N_2186);
or U4751 (N_4751,N_2532,N_2003);
or U4752 (N_4752,N_2779,N_2575);
nand U4753 (N_4753,N_2014,N_2641);
and U4754 (N_4754,N_3134,N_3609);
and U4755 (N_4755,N_2555,N_3092);
and U4756 (N_4756,N_3406,N_2101);
nand U4757 (N_4757,N_3979,N_2616);
nand U4758 (N_4758,N_3265,N_2107);
nor U4759 (N_4759,N_2775,N_3942);
nand U4760 (N_4760,N_2796,N_3830);
nor U4761 (N_4761,N_3058,N_2009);
and U4762 (N_4762,N_3919,N_3072);
nor U4763 (N_4763,N_3282,N_3881);
and U4764 (N_4764,N_3081,N_2741);
nand U4765 (N_4765,N_3413,N_3780);
nor U4766 (N_4766,N_2253,N_2899);
nand U4767 (N_4767,N_2873,N_3161);
or U4768 (N_4768,N_3297,N_3451);
and U4769 (N_4769,N_3767,N_2450);
and U4770 (N_4770,N_3524,N_3827);
and U4771 (N_4771,N_2141,N_3577);
and U4772 (N_4772,N_2565,N_2546);
or U4773 (N_4773,N_3579,N_2581);
nor U4774 (N_4774,N_3766,N_3640);
xnor U4775 (N_4775,N_3151,N_3528);
and U4776 (N_4776,N_3715,N_3311);
nand U4777 (N_4777,N_3239,N_3562);
nor U4778 (N_4778,N_3915,N_3127);
or U4779 (N_4779,N_2179,N_3436);
and U4780 (N_4780,N_2453,N_3404);
xnor U4781 (N_4781,N_2947,N_3342);
or U4782 (N_4782,N_3662,N_2326);
or U4783 (N_4783,N_2822,N_2795);
or U4784 (N_4784,N_3382,N_3099);
nand U4785 (N_4785,N_3203,N_3648);
or U4786 (N_4786,N_2831,N_3660);
and U4787 (N_4787,N_3755,N_2615);
nor U4788 (N_4788,N_2360,N_3627);
nand U4789 (N_4789,N_3731,N_2955);
nand U4790 (N_4790,N_3054,N_2209);
nor U4791 (N_4791,N_2550,N_2514);
nor U4792 (N_4792,N_2037,N_3982);
nor U4793 (N_4793,N_2522,N_2254);
nand U4794 (N_4794,N_3753,N_3039);
and U4795 (N_4795,N_3205,N_2413);
nor U4796 (N_4796,N_2031,N_2256);
nor U4797 (N_4797,N_3547,N_2455);
nand U4798 (N_4798,N_2986,N_2086);
nand U4799 (N_4799,N_2629,N_2119);
or U4800 (N_4800,N_3019,N_3372);
nor U4801 (N_4801,N_3997,N_2197);
and U4802 (N_4802,N_2959,N_3759);
or U4803 (N_4803,N_3359,N_2192);
nor U4804 (N_4804,N_3909,N_2227);
and U4805 (N_4805,N_2659,N_2010);
nor U4806 (N_4806,N_2728,N_3198);
or U4807 (N_4807,N_3367,N_3911);
nand U4808 (N_4808,N_2393,N_2720);
nand U4809 (N_4809,N_3104,N_3023);
and U4810 (N_4810,N_2441,N_2109);
nand U4811 (N_4811,N_3920,N_3164);
and U4812 (N_4812,N_3459,N_2027);
or U4813 (N_4813,N_2560,N_3066);
nor U4814 (N_4814,N_3888,N_2224);
and U4815 (N_4815,N_2496,N_3768);
and U4816 (N_4816,N_3600,N_2585);
nor U4817 (N_4817,N_3290,N_2730);
nand U4818 (N_4818,N_2016,N_3603);
or U4819 (N_4819,N_2923,N_3355);
and U4820 (N_4820,N_3854,N_3758);
nand U4821 (N_4821,N_3389,N_3981);
and U4822 (N_4822,N_2662,N_3181);
nand U4823 (N_4823,N_3328,N_3849);
nor U4824 (N_4824,N_2757,N_2429);
xnor U4825 (N_4825,N_2375,N_2364);
or U4826 (N_4826,N_2398,N_3554);
and U4827 (N_4827,N_3748,N_3402);
nand U4828 (N_4828,N_2976,N_3975);
nor U4829 (N_4829,N_3329,N_2848);
nand U4830 (N_4830,N_3540,N_2410);
or U4831 (N_4831,N_3456,N_3073);
nor U4832 (N_4832,N_2077,N_3913);
nand U4833 (N_4833,N_2404,N_2105);
and U4834 (N_4834,N_3834,N_2015);
nor U4835 (N_4835,N_2517,N_2223);
or U4836 (N_4836,N_3697,N_2407);
and U4837 (N_4837,N_2683,N_2437);
or U4838 (N_4838,N_2305,N_2317);
nor U4839 (N_4839,N_2767,N_2812);
nor U4840 (N_4840,N_2639,N_3222);
or U4841 (N_4841,N_2749,N_2198);
or U4842 (N_4842,N_2034,N_3962);
or U4843 (N_4843,N_2267,N_2679);
and U4844 (N_4844,N_2689,N_3481);
nand U4845 (N_4845,N_2319,N_2225);
nand U4846 (N_4846,N_3882,N_3551);
and U4847 (N_4847,N_3644,N_3258);
and U4848 (N_4848,N_3278,N_2724);
and U4849 (N_4849,N_2693,N_3288);
nor U4850 (N_4850,N_3043,N_3444);
and U4851 (N_4851,N_2999,N_3409);
or U4852 (N_4852,N_2751,N_3279);
nand U4853 (N_4853,N_3978,N_3886);
xor U4854 (N_4854,N_3281,N_3951);
or U4855 (N_4855,N_2111,N_2762);
nor U4856 (N_4856,N_3803,N_2108);
nor U4857 (N_4857,N_2816,N_2160);
nor U4858 (N_4858,N_3421,N_3030);
nor U4859 (N_4859,N_2386,N_2677);
nor U4860 (N_4860,N_2024,N_2451);
and U4861 (N_4861,N_3805,N_2143);
nor U4862 (N_4862,N_3125,N_2385);
or U4863 (N_4863,N_2213,N_2647);
xnor U4864 (N_4864,N_2277,N_3428);
nand U4865 (N_4865,N_3417,N_2486);
nand U4866 (N_4866,N_2633,N_3958);
nor U4867 (N_4867,N_2066,N_3851);
nand U4868 (N_4868,N_3434,N_2322);
nand U4869 (N_4869,N_3115,N_3004);
and U4870 (N_4870,N_2106,N_2968);
and U4871 (N_4871,N_3937,N_2777);
nor U4872 (N_4872,N_3934,N_3407);
nor U4873 (N_4873,N_2554,N_3553);
or U4874 (N_4874,N_2065,N_3254);
nor U4875 (N_4875,N_3300,N_2763);
nand U4876 (N_4876,N_2669,N_3168);
and U4877 (N_4877,N_3082,N_2998);
nand U4878 (N_4878,N_3772,N_3741);
nor U4879 (N_4879,N_2032,N_2219);
or U4880 (N_4880,N_3040,N_2164);
nor U4881 (N_4881,N_3446,N_2240);
nand U4882 (N_4882,N_3435,N_3679);
and U4883 (N_4883,N_2215,N_3262);
and U4884 (N_4884,N_2005,N_3162);
nand U4885 (N_4885,N_2207,N_3572);
nor U4886 (N_4886,N_2118,N_2367);
xnor U4887 (N_4887,N_3457,N_2368);
nand U4888 (N_4888,N_2493,N_2492);
nand U4889 (N_4889,N_2676,N_3306);
or U4890 (N_4890,N_3313,N_3681);
nor U4891 (N_4891,N_3206,N_2987);
or U4892 (N_4892,N_3037,N_3620);
nand U4893 (N_4893,N_3445,N_3795);
nor U4894 (N_4894,N_2996,N_2880);
or U4895 (N_4895,N_2184,N_3138);
and U4896 (N_4896,N_3088,N_2416);
and U4897 (N_4897,N_2868,N_3914);
or U4898 (N_4898,N_3779,N_3320);
and U4899 (N_4899,N_2849,N_2000);
or U4900 (N_4900,N_3512,N_3063);
nor U4901 (N_4901,N_3817,N_2835);
nor U4902 (N_4902,N_2250,N_3654);
or U4903 (N_4903,N_2328,N_3071);
nand U4904 (N_4904,N_2509,N_2595);
nor U4905 (N_4905,N_2788,N_3123);
nor U4906 (N_4906,N_2226,N_3323);
nand U4907 (N_4907,N_3729,N_3696);
nand U4908 (N_4908,N_3514,N_2162);
nand U4909 (N_4909,N_3053,N_3260);
and U4910 (N_4910,N_2411,N_3619);
nor U4911 (N_4911,N_3801,N_3983);
nor U4912 (N_4912,N_2144,N_3048);
nor U4913 (N_4913,N_2934,N_2485);
nand U4914 (N_4914,N_3659,N_3111);
nor U4915 (N_4915,N_2985,N_3657);
nor U4916 (N_4916,N_3462,N_2975);
or U4917 (N_4917,N_3392,N_2205);
nor U4918 (N_4918,N_3231,N_3918);
or U4919 (N_4919,N_2700,N_2236);
nand U4920 (N_4920,N_2810,N_3431);
or U4921 (N_4921,N_2738,N_2483);
or U4922 (N_4922,N_2503,N_3810);
nor U4923 (N_4923,N_3466,N_2991);
xor U4924 (N_4924,N_2489,N_3947);
or U4925 (N_4925,N_3971,N_2526);
nor U4926 (N_4926,N_3637,N_2644);
nor U4927 (N_4927,N_3401,N_2839);
nand U4928 (N_4928,N_2592,N_3467);
and U4929 (N_4929,N_2181,N_2979);
nand U4930 (N_4930,N_3490,N_3604);
nand U4931 (N_4931,N_2347,N_3460);
nor U4932 (N_4932,N_3298,N_3440);
and U4933 (N_4933,N_2845,N_2614);
nor U4934 (N_4934,N_2327,N_3773);
or U4935 (N_4935,N_2269,N_3243);
nand U4936 (N_4936,N_3885,N_3878);
nor U4937 (N_4937,N_3469,N_3829);
and U4938 (N_4938,N_3567,N_2421);
nand U4939 (N_4939,N_2074,N_3163);
or U4940 (N_4940,N_2783,N_3999);
and U4941 (N_4941,N_3747,N_2335);
nor U4942 (N_4942,N_2894,N_3566);
or U4943 (N_4943,N_2813,N_3774);
or U4944 (N_4944,N_2057,N_2502);
and U4945 (N_4945,N_3676,N_3018);
nand U4946 (N_4946,N_2961,N_3527);
nor U4947 (N_4947,N_2131,N_2221);
and U4948 (N_4948,N_3484,N_3270);
nor U4949 (N_4949,N_2523,N_3454);
or U4950 (N_4950,N_2612,N_3499);
or U4951 (N_4951,N_3105,N_2787);
and U4952 (N_4952,N_3615,N_3534);
nand U4953 (N_4953,N_3521,N_2072);
nand U4954 (N_4954,N_3034,N_3186);
nand U4955 (N_4955,N_2772,N_2432);
or U4956 (N_4956,N_3964,N_2358);
xnor U4957 (N_4957,N_2802,N_3783);
or U4958 (N_4958,N_3989,N_3061);
nand U4959 (N_4959,N_2017,N_3525);
nor U4960 (N_4960,N_2622,N_3806);
or U4961 (N_4961,N_3006,N_2598);
nand U4962 (N_4962,N_2752,N_3241);
and U4963 (N_4963,N_3912,N_2474);
nor U4964 (N_4964,N_2545,N_3415);
xnor U4965 (N_4965,N_2623,N_2002);
xor U4966 (N_4966,N_3613,N_3117);
or U4967 (N_4967,N_2760,N_2742);
nor U4968 (N_4968,N_2193,N_2067);
and U4969 (N_4969,N_3316,N_3864);
nand U4970 (N_4970,N_2843,N_3232);
nand U4971 (N_4971,N_3237,N_2472);
or U4972 (N_4972,N_2473,N_3067);
nor U4973 (N_4973,N_3651,N_3727);
or U4974 (N_4974,N_2321,N_2651);
or U4975 (N_4975,N_3325,N_3153);
nor U4976 (N_4976,N_2743,N_2518);
nand U4977 (N_4977,N_3639,N_2665);
or U4978 (N_4978,N_2149,N_3103);
or U4979 (N_4979,N_3582,N_2962);
or U4980 (N_4980,N_3891,N_3188);
and U4981 (N_4981,N_2865,N_2710);
or U4982 (N_4982,N_3438,N_2885);
xnor U4983 (N_4983,N_3564,N_3394);
nand U4984 (N_4984,N_2840,N_3828);
nor U4985 (N_4985,N_2707,N_2415);
or U4986 (N_4986,N_2058,N_3561);
nor U4987 (N_4987,N_2834,N_2395);
nor U4988 (N_4988,N_3135,N_2832);
and U4989 (N_4989,N_3353,N_2929);
nor U4990 (N_4990,N_3387,N_2558);
and U4991 (N_4991,N_3069,N_3737);
or U4992 (N_4992,N_2723,N_2159);
nor U4993 (N_4993,N_3970,N_2475);
and U4994 (N_4994,N_2443,N_3761);
and U4995 (N_4995,N_3673,N_3379);
nor U4996 (N_4996,N_3542,N_2314);
or U4997 (N_4997,N_3733,N_3595);
or U4998 (N_4998,N_2054,N_3339);
and U4999 (N_4999,N_3873,N_3922);
and U5000 (N_5000,N_2161,N_3061);
and U5001 (N_5001,N_3085,N_3354);
nor U5002 (N_5002,N_3053,N_2451);
or U5003 (N_5003,N_3726,N_3974);
or U5004 (N_5004,N_3558,N_3718);
nand U5005 (N_5005,N_2957,N_3155);
and U5006 (N_5006,N_3030,N_3899);
nand U5007 (N_5007,N_2185,N_2848);
or U5008 (N_5008,N_2459,N_3569);
nor U5009 (N_5009,N_2309,N_2490);
and U5010 (N_5010,N_2835,N_2222);
and U5011 (N_5011,N_2465,N_3827);
nor U5012 (N_5012,N_2452,N_3477);
and U5013 (N_5013,N_2840,N_3423);
or U5014 (N_5014,N_2137,N_2219);
nand U5015 (N_5015,N_3363,N_2920);
and U5016 (N_5016,N_3168,N_2730);
and U5017 (N_5017,N_2646,N_2327);
nor U5018 (N_5018,N_2124,N_2389);
and U5019 (N_5019,N_2275,N_2574);
or U5020 (N_5020,N_3468,N_3682);
and U5021 (N_5021,N_2862,N_2119);
and U5022 (N_5022,N_2744,N_2623);
nor U5023 (N_5023,N_3531,N_2474);
nor U5024 (N_5024,N_3182,N_3684);
or U5025 (N_5025,N_2413,N_3911);
nor U5026 (N_5026,N_2929,N_3184);
nor U5027 (N_5027,N_3817,N_2864);
nand U5028 (N_5028,N_2315,N_2243);
nor U5029 (N_5029,N_3273,N_3055);
nor U5030 (N_5030,N_3027,N_2701);
or U5031 (N_5031,N_3154,N_3041);
nor U5032 (N_5032,N_3914,N_2700);
nor U5033 (N_5033,N_2970,N_3798);
nand U5034 (N_5034,N_3467,N_2079);
nor U5035 (N_5035,N_2430,N_2299);
nor U5036 (N_5036,N_3857,N_2811);
and U5037 (N_5037,N_3600,N_2588);
nand U5038 (N_5038,N_3157,N_2512);
nor U5039 (N_5039,N_3648,N_3798);
or U5040 (N_5040,N_2419,N_2728);
and U5041 (N_5041,N_3269,N_2792);
or U5042 (N_5042,N_2624,N_3091);
nor U5043 (N_5043,N_2722,N_2799);
or U5044 (N_5044,N_2632,N_2071);
xor U5045 (N_5045,N_3610,N_2575);
or U5046 (N_5046,N_2807,N_2064);
and U5047 (N_5047,N_3311,N_3817);
nor U5048 (N_5048,N_2359,N_2713);
nor U5049 (N_5049,N_2290,N_3443);
nor U5050 (N_5050,N_2496,N_2648);
and U5051 (N_5051,N_2833,N_3003);
nor U5052 (N_5052,N_3739,N_3309);
or U5053 (N_5053,N_2249,N_3713);
and U5054 (N_5054,N_2704,N_3656);
and U5055 (N_5055,N_3480,N_2955);
nand U5056 (N_5056,N_2984,N_2322);
nand U5057 (N_5057,N_2478,N_3514);
and U5058 (N_5058,N_2565,N_2278);
nor U5059 (N_5059,N_2539,N_2410);
nand U5060 (N_5060,N_3863,N_2449);
and U5061 (N_5061,N_3384,N_2287);
nor U5062 (N_5062,N_3047,N_2657);
or U5063 (N_5063,N_3367,N_2274);
and U5064 (N_5064,N_3678,N_2790);
and U5065 (N_5065,N_2081,N_3731);
nor U5066 (N_5066,N_2689,N_3389);
nor U5067 (N_5067,N_3768,N_3524);
nand U5068 (N_5068,N_3724,N_3837);
or U5069 (N_5069,N_3938,N_3595);
or U5070 (N_5070,N_2538,N_3218);
and U5071 (N_5071,N_2734,N_2045);
nand U5072 (N_5072,N_2331,N_2177);
and U5073 (N_5073,N_3449,N_2362);
and U5074 (N_5074,N_2611,N_3592);
and U5075 (N_5075,N_2598,N_2686);
nor U5076 (N_5076,N_2349,N_3579);
nor U5077 (N_5077,N_3510,N_3995);
or U5078 (N_5078,N_3836,N_2442);
nand U5079 (N_5079,N_2343,N_2787);
or U5080 (N_5080,N_3581,N_3531);
or U5081 (N_5081,N_2821,N_3744);
and U5082 (N_5082,N_2014,N_3691);
nand U5083 (N_5083,N_2944,N_2441);
or U5084 (N_5084,N_3756,N_3444);
nand U5085 (N_5085,N_2935,N_3462);
nor U5086 (N_5086,N_2682,N_3295);
or U5087 (N_5087,N_2497,N_3477);
nor U5088 (N_5088,N_2652,N_2917);
xnor U5089 (N_5089,N_2688,N_2189);
nor U5090 (N_5090,N_3465,N_3757);
or U5091 (N_5091,N_3957,N_3653);
or U5092 (N_5092,N_2919,N_3349);
nand U5093 (N_5093,N_3967,N_3470);
nand U5094 (N_5094,N_3907,N_2642);
and U5095 (N_5095,N_3835,N_3808);
nor U5096 (N_5096,N_3619,N_3880);
nor U5097 (N_5097,N_3004,N_2610);
nor U5098 (N_5098,N_3307,N_3749);
nor U5099 (N_5099,N_2856,N_2550);
and U5100 (N_5100,N_3954,N_2622);
nand U5101 (N_5101,N_2250,N_2304);
or U5102 (N_5102,N_3105,N_3622);
nand U5103 (N_5103,N_2617,N_3390);
and U5104 (N_5104,N_2739,N_3597);
nor U5105 (N_5105,N_3217,N_3767);
and U5106 (N_5106,N_2346,N_2960);
nor U5107 (N_5107,N_3356,N_2582);
nand U5108 (N_5108,N_2401,N_2046);
or U5109 (N_5109,N_2573,N_3342);
nor U5110 (N_5110,N_3728,N_3733);
or U5111 (N_5111,N_2786,N_2342);
nor U5112 (N_5112,N_2198,N_2595);
nor U5113 (N_5113,N_2732,N_3288);
and U5114 (N_5114,N_3053,N_3910);
nand U5115 (N_5115,N_3267,N_3993);
nor U5116 (N_5116,N_3893,N_3316);
nor U5117 (N_5117,N_3898,N_2234);
nor U5118 (N_5118,N_3429,N_2067);
and U5119 (N_5119,N_3187,N_2987);
nand U5120 (N_5120,N_2272,N_3025);
or U5121 (N_5121,N_3702,N_3455);
or U5122 (N_5122,N_3168,N_3319);
nor U5123 (N_5123,N_2989,N_2227);
or U5124 (N_5124,N_2148,N_2082);
nor U5125 (N_5125,N_2724,N_3551);
nor U5126 (N_5126,N_3068,N_2123);
nor U5127 (N_5127,N_2950,N_2727);
and U5128 (N_5128,N_2218,N_3534);
and U5129 (N_5129,N_2412,N_3669);
and U5130 (N_5130,N_2965,N_3843);
xor U5131 (N_5131,N_2258,N_2186);
nand U5132 (N_5132,N_2554,N_3732);
nand U5133 (N_5133,N_3029,N_2001);
and U5134 (N_5134,N_2687,N_3878);
nand U5135 (N_5135,N_3896,N_3177);
nor U5136 (N_5136,N_3693,N_2325);
or U5137 (N_5137,N_2462,N_3871);
nand U5138 (N_5138,N_3144,N_2541);
nor U5139 (N_5139,N_3846,N_2500);
nand U5140 (N_5140,N_3754,N_2205);
or U5141 (N_5141,N_3891,N_2129);
nand U5142 (N_5142,N_3530,N_2746);
or U5143 (N_5143,N_2296,N_3738);
nand U5144 (N_5144,N_3217,N_2146);
nor U5145 (N_5145,N_3502,N_3494);
nand U5146 (N_5146,N_2659,N_2885);
and U5147 (N_5147,N_2141,N_2635);
nand U5148 (N_5148,N_3849,N_2332);
or U5149 (N_5149,N_2457,N_2403);
and U5150 (N_5150,N_2258,N_2715);
nand U5151 (N_5151,N_2213,N_3130);
or U5152 (N_5152,N_2814,N_3622);
or U5153 (N_5153,N_2697,N_3444);
nand U5154 (N_5154,N_2420,N_3934);
and U5155 (N_5155,N_2576,N_3745);
or U5156 (N_5156,N_3932,N_2281);
or U5157 (N_5157,N_3069,N_3255);
and U5158 (N_5158,N_3510,N_2341);
and U5159 (N_5159,N_2152,N_3131);
or U5160 (N_5160,N_3663,N_3661);
nand U5161 (N_5161,N_3693,N_2026);
and U5162 (N_5162,N_3138,N_2943);
or U5163 (N_5163,N_3206,N_2465);
nor U5164 (N_5164,N_3334,N_3764);
nor U5165 (N_5165,N_3605,N_3313);
nand U5166 (N_5166,N_3592,N_3954);
nand U5167 (N_5167,N_3674,N_2773);
or U5168 (N_5168,N_3077,N_3429);
or U5169 (N_5169,N_3340,N_2804);
nor U5170 (N_5170,N_2388,N_3911);
or U5171 (N_5171,N_2933,N_2057);
nor U5172 (N_5172,N_2499,N_3210);
and U5173 (N_5173,N_2556,N_3947);
nor U5174 (N_5174,N_2155,N_2680);
or U5175 (N_5175,N_2885,N_2364);
nor U5176 (N_5176,N_2880,N_2648);
nor U5177 (N_5177,N_2149,N_3652);
and U5178 (N_5178,N_3427,N_3671);
nor U5179 (N_5179,N_2862,N_3193);
nand U5180 (N_5180,N_3354,N_2041);
and U5181 (N_5181,N_2416,N_3350);
nor U5182 (N_5182,N_3692,N_3453);
nor U5183 (N_5183,N_2498,N_2438);
nand U5184 (N_5184,N_2374,N_2945);
and U5185 (N_5185,N_2004,N_3349);
or U5186 (N_5186,N_3442,N_3406);
and U5187 (N_5187,N_3609,N_3113);
or U5188 (N_5188,N_2189,N_3248);
or U5189 (N_5189,N_2518,N_3749);
or U5190 (N_5190,N_3494,N_2275);
and U5191 (N_5191,N_2104,N_3008);
nand U5192 (N_5192,N_3187,N_3928);
nor U5193 (N_5193,N_3178,N_3590);
or U5194 (N_5194,N_3732,N_3301);
nor U5195 (N_5195,N_3823,N_3711);
xor U5196 (N_5196,N_3701,N_2551);
nor U5197 (N_5197,N_2477,N_2203);
or U5198 (N_5198,N_3739,N_3872);
nand U5199 (N_5199,N_3146,N_2080);
and U5200 (N_5200,N_2379,N_2188);
nor U5201 (N_5201,N_3803,N_3680);
and U5202 (N_5202,N_2106,N_2400);
or U5203 (N_5203,N_2169,N_3522);
xor U5204 (N_5204,N_2845,N_2928);
nor U5205 (N_5205,N_2647,N_2934);
nor U5206 (N_5206,N_2168,N_3978);
nor U5207 (N_5207,N_2739,N_3316);
or U5208 (N_5208,N_2053,N_2922);
nor U5209 (N_5209,N_3852,N_2688);
and U5210 (N_5210,N_2733,N_2143);
and U5211 (N_5211,N_3506,N_3701);
or U5212 (N_5212,N_3717,N_2835);
or U5213 (N_5213,N_2616,N_2686);
nor U5214 (N_5214,N_2742,N_3043);
and U5215 (N_5215,N_3541,N_3205);
or U5216 (N_5216,N_2265,N_3886);
nand U5217 (N_5217,N_3657,N_3737);
and U5218 (N_5218,N_3250,N_2498);
nand U5219 (N_5219,N_3721,N_2773);
nand U5220 (N_5220,N_3837,N_2632);
nand U5221 (N_5221,N_3828,N_3462);
and U5222 (N_5222,N_3417,N_2044);
nor U5223 (N_5223,N_3244,N_2936);
nor U5224 (N_5224,N_3926,N_3155);
and U5225 (N_5225,N_3944,N_3362);
nor U5226 (N_5226,N_2251,N_3523);
nor U5227 (N_5227,N_2364,N_3634);
nand U5228 (N_5228,N_3719,N_2573);
nand U5229 (N_5229,N_3786,N_3858);
xor U5230 (N_5230,N_3251,N_2039);
nor U5231 (N_5231,N_3372,N_3321);
nor U5232 (N_5232,N_2306,N_2897);
nand U5233 (N_5233,N_2693,N_2475);
nor U5234 (N_5234,N_3986,N_3293);
or U5235 (N_5235,N_2039,N_3452);
and U5236 (N_5236,N_2963,N_2910);
nand U5237 (N_5237,N_2486,N_2267);
or U5238 (N_5238,N_3236,N_3074);
nor U5239 (N_5239,N_3005,N_3771);
nor U5240 (N_5240,N_2776,N_3538);
and U5241 (N_5241,N_3992,N_3971);
and U5242 (N_5242,N_3226,N_3818);
nand U5243 (N_5243,N_3734,N_2680);
and U5244 (N_5244,N_3899,N_3012);
nand U5245 (N_5245,N_3870,N_2970);
or U5246 (N_5246,N_3577,N_2505);
nor U5247 (N_5247,N_3833,N_2617);
or U5248 (N_5248,N_2018,N_2033);
nand U5249 (N_5249,N_3972,N_3003);
nand U5250 (N_5250,N_3392,N_2782);
nand U5251 (N_5251,N_3103,N_3510);
and U5252 (N_5252,N_2799,N_2257);
or U5253 (N_5253,N_3681,N_3493);
nand U5254 (N_5254,N_2546,N_2124);
xnor U5255 (N_5255,N_2414,N_3787);
and U5256 (N_5256,N_2431,N_2825);
or U5257 (N_5257,N_3133,N_3566);
or U5258 (N_5258,N_2757,N_2324);
and U5259 (N_5259,N_2930,N_3270);
or U5260 (N_5260,N_2445,N_2722);
or U5261 (N_5261,N_2535,N_2790);
nand U5262 (N_5262,N_3627,N_2926);
and U5263 (N_5263,N_2295,N_3267);
nor U5264 (N_5264,N_3702,N_2906);
and U5265 (N_5265,N_3871,N_3006);
and U5266 (N_5266,N_3914,N_3253);
or U5267 (N_5267,N_2522,N_3526);
nand U5268 (N_5268,N_3548,N_2880);
or U5269 (N_5269,N_2249,N_2221);
nor U5270 (N_5270,N_2274,N_2127);
nand U5271 (N_5271,N_3697,N_3723);
or U5272 (N_5272,N_3299,N_2506);
or U5273 (N_5273,N_3083,N_2331);
or U5274 (N_5274,N_2814,N_2894);
xor U5275 (N_5275,N_3041,N_2064);
and U5276 (N_5276,N_2482,N_3699);
nor U5277 (N_5277,N_3767,N_2809);
and U5278 (N_5278,N_2958,N_2107);
and U5279 (N_5279,N_3039,N_3654);
or U5280 (N_5280,N_3578,N_2521);
and U5281 (N_5281,N_2771,N_3583);
nand U5282 (N_5282,N_2513,N_2040);
or U5283 (N_5283,N_3159,N_3036);
nor U5284 (N_5284,N_3340,N_2651);
nand U5285 (N_5285,N_2730,N_2472);
and U5286 (N_5286,N_3498,N_3581);
or U5287 (N_5287,N_3916,N_2888);
nor U5288 (N_5288,N_3907,N_2895);
and U5289 (N_5289,N_3701,N_2732);
nand U5290 (N_5290,N_2300,N_3010);
nand U5291 (N_5291,N_3202,N_2823);
or U5292 (N_5292,N_2242,N_2131);
or U5293 (N_5293,N_3248,N_3280);
xnor U5294 (N_5294,N_3364,N_3864);
and U5295 (N_5295,N_3230,N_3698);
nand U5296 (N_5296,N_2534,N_2754);
nand U5297 (N_5297,N_3429,N_2867);
and U5298 (N_5298,N_2351,N_2106);
or U5299 (N_5299,N_2306,N_2889);
or U5300 (N_5300,N_2091,N_3270);
or U5301 (N_5301,N_3830,N_2614);
nor U5302 (N_5302,N_3374,N_2613);
nand U5303 (N_5303,N_3610,N_2753);
nand U5304 (N_5304,N_2997,N_2934);
and U5305 (N_5305,N_3890,N_2104);
and U5306 (N_5306,N_3415,N_2301);
nand U5307 (N_5307,N_3210,N_3675);
nor U5308 (N_5308,N_2702,N_2355);
or U5309 (N_5309,N_3772,N_3904);
nor U5310 (N_5310,N_3130,N_2426);
nand U5311 (N_5311,N_2484,N_2135);
nor U5312 (N_5312,N_3642,N_3035);
and U5313 (N_5313,N_3081,N_3132);
and U5314 (N_5314,N_3116,N_3115);
nor U5315 (N_5315,N_3821,N_2658);
and U5316 (N_5316,N_3220,N_3469);
xor U5317 (N_5317,N_3493,N_3382);
nand U5318 (N_5318,N_3622,N_3881);
and U5319 (N_5319,N_2239,N_3171);
nand U5320 (N_5320,N_2780,N_2186);
or U5321 (N_5321,N_3170,N_2234);
and U5322 (N_5322,N_2699,N_2561);
nand U5323 (N_5323,N_3130,N_3754);
nor U5324 (N_5324,N_2391,N_3329);
or U5325 (N_5325,N_3595,N_3251);
xor U5326 (N_5326,N_3002,N_2368);
or U5327 (N_5327,N_3971,N_2815);
nand U5328 (N_5328,N_2590,N_3572);
nand U5329 (N_5329,N_2891,N_2493);
xnor U5330 (N_5330,N_3965,N_3105);
nor U5331 (N_5331,N_3976,N_2601);
and U5332 (N_5332,N_2725,N_2416);
or U5333 (N_5333,N_2014,N_2205);
or U5334 (N_5334,N_2899,N_3572);
and U5335 (N_5335,N_2811,N_3683);
nor U5336 (N_5336,N_2627,N_3919);
nor U5337 (N_5337,N_2161,N_2215);
nor U5338 (N_5338,N_3896,N_3698);
or U5339 (N_5339,N_2518,N_2419);
nand U5340 (N_5340,N_2099,N_3435);
or U5341 (N_5341,N_3972,N_3939);
and U5342 (N_5342,N_3067,N_3478);
or U5343 (N_5343,N_2936,N_3309);
and U5344 (N_5344,N_3680,N_3692);
and U5345 (N_5345,N_3396,N_2684);
nor U5346 (N_5346,N_3808,N_2138);
or U5347 (N_5347,N_3983,N_3991);
and U5348 (N_5348,N_2211,N_3250);
or U5349 (N_5349,N_3959,N_2225);
nand U5350 (N_5350,N_3316,N_2919);
and U5351 (N_5351,N_3351,N_3259);
and U5352 (N_5352,N_2101,N_3859);
or U5353 (N_5353,N_3688,N_3352);
nand U5354 (N_5354,N_3379,N_3098);
nor U5355 (N_5355,N_2794,N_2989);
and U5356 (N_5356,N_2097,N_3075);
nand U5357 (N_5357,N_3382,N_2323);
or U5358 (N_5358,N_2110,N_3827);
or U5359 (N_5359,N_2316,N_2058);
and U5360 (N_5360,N_2134,N_2591);
and U5361 (N_5361,N_2284,N_2667);
nor U5362 (N_5362,N_3366,N_3616);
and U5363 (N_5363,N_2630,N_2517);
or U5364 (N_5364,N_3576,N_3583);
nand U5365 (N_5365,N_2432,N_2203);
nor U5366 (N_5366,N_2749,N_3451);
or U5367 (N_5367,N_2146,N_3610);
nand U5368 (N_5368,N_3968,N_3058);
or U5369 (N_5369,N_3096,N_2424);
xnor U5370 (N_5370,N_2513,N_3337);
or U5371 (N_5371,N_2411,N_2143);
and U5372 (N_5372,N_2544,N_2566);
nand U5373 (N_5373,N_2029,N_3220);
nand U5374 (N_5374,N_2397,N_2776);
nor U5375 (N_5375,N_3966,N_2310);
or U5376 (N_5376,N_2270,N_3204);
and U5377 (N_5377,N_2405,N_3744);
nor U5378 (N_5378,N_2148,N_2964);
nor U5379 (N_5379,N_3847,N_3485);
or U5380 (N_5380,N_2704,N_2850);
or U5381 (N_5381,N_3147,N_3635);
or U5382 (N_5382,N_3722,N_2756);
nor U5383 (N_5383,N_3968,N_2226);
nand U5384 (N_5384,N_3586,N_3052);
nand U5385 (N_5385,N_3320,N_2344);
nand U5386 (N_5386,N_2902,N_3124);
or U5387 (N_5387,N_2795,N_2361);
nor U5388 (N_5388,N_2295,N_2309);
or U5389 (N_5389,N_2498,N_2152);
nand U5390 (N_5390,N_3502,N_3271);
and U5391 (N_5391,N_2830,N_3284);
or U5392 (N_5392,N_2533,N_2184);
nor U5393 (N_5393,N_3160,N_2039);
and U5394 (N_5394,N_3565,N_2693);
nand U5395 (N_5395,N_2679,N_3637);
nand U5396 (N_5396,N_2568,N_3038);
nand U5397 (N_5397,N_2576,N_3491);
nor U5398 (N_5398,N_3528,N_2180);
or U5399 (N_5399,N_2389,N_2645);
or U5400 (N_5400,N_3688,N_2226);
or U5401 (N_5401,N_3329,N_3346);
and U5402 (N_5402,N_2833,N_2830);
nor U5403 (N_5403,N_2392,N_3550);
nor U5404 (N_5404,N_2124,N_2642);
xnor U5405 (N_5405,N_2906,N_2677);
nand U5406 (N_5406,N_3312,N_2713);
or U5407 (N_5407,N_3764,N_3312);
and U5408 (N_5408,N_2697,N_2239);
or U5409 (N_5409,N_2902,N_2038);
and U5410 (N_5410,N_3307,N_2402);
and U5411 (N_5411,N_2042,N_3273);
nor U5412 (N_5412,N_3363,N_3728);
or U5413 (N_5413,N_3844,N_3745);
or U5414 (N_5414,N_2304,N_2042);
and U5415 (N_5415,N_2213,N_3122);
and U5416 (N_5416,N_3104,N_2223);
nand U5417 (N_5417,N_3249,N_3007);
nand U5418 (N_5418,N_2532,N_3669);
or U5419 (N_5419,N_3694,N_3501);
and U5420 (N_5420,N_2436,N_3353);
and U5421 (N_5421,N_3486,N_2796);
nand U5422 (N_5422,N_2533,N_3949);
nor U5423 (N_5423,N_2243,N_3657);
and U5424 (N_5424,N_2078,N_2790);
nor U5425 (N_5425,N_2623,N_3336);
nand U5426 (N_5426,N_3625,N_3766);
nand U5427 (N_5427,N_3793,N_2431);
or U5428 (N_5428,N_2662,N_3535);
or U5429 (N_5429,N_3414,N_3311);
nand U5430 (N_5430,N_2076,N_2942);
or U5431 (N_5431,N_3170,N_3868);
nor U5432 (N_5432,N_2043,N_3767);
nor U5433 (N_5433,N_3216,N_2266);
nor U5434 (N_5434,N_2816,N_2460);
or U5435 (N_5435,N_3701,N_2099);
nor U5436 (N_5436,N_2399,N_3520);
and U5437 (N_5437,N_2057,N_2149);
nand U5438 (N_5438,N_2926,N_2011);
and U5439 (N_5439,N_3617,N_2849);
nand U5440 (N_5440,N_3941,N_3682);
nand U5441 (N_5441,N_3059,N_2352);
nor U5442 (N_5442,N_3441,N_2444);
xnor U5443 (N_5443,N_2404,N_2198);
nor U5444 (N_5444,N_3119,N_3641);
nor U5445 (N_5445,N_3134,N_3031);
nor U5446 (N_5446,N_2495,N_2820);
nor U5447 (N_5447,N_2327,N_3371);
and U5448 (N_5448,N_3588,N_2111);
or U5449 (N_5449,N_3079,N_3482);
nor U5450 (N_5450,N_2337,N_3398);
and U5451 (N_5451,N_3141,N_2844);
nor U5452 (N_5452,N_2113,N_3598);
nand U5453 (N_5453,N_3014,N_2812);
and U5454 (N_5454,N_3098,N_3971);
nand U5455 (N_5455,N_3572,N_2963);
or U5456 (N_5456,N_2996,N_3106);
nor U5457 (N_5457,N_3170,N_3632);
and U5458 (N_5458,N_3599,N_3668);
nor U5459 (N_5459,N_3510,N_3210);
or U5460 (N_5460,N_3561,N_3275);
and U5461 (N_5461,N_3977,N_2081);
and U5462 (N_5462,N_2543,N_2528);
or U5463 (N_5463,N_2768,N_3423);
and U5464 (N_5464,N_3440,N_3575);
xor U5465 (N_5465,N_2923,N_3807);
and U5466 (N_5466,N_3272,N_3753);
or U5467 (N_5467,N_2166,N_3039);
or U5468 (N_5468,N_3744,N_2769);
and U5469 (N_5469,N_3450,N_2946);
or U5470 (N_5470,N_2516,N_2895);
nand U5471 (N_5471,N_3483,N_2141);
nor U5472 (N_5472,N_3819,N_2424);
nand U5473 (N_5473,N_2463,N_2867);
nor U5474 (N_5474,N_2223,N_2680);
and U5475 (N_5475,N_3149,N_3479);
nor U5476 (N_5476,N_3370,N_3056);
nor U5477 (N_5477,N_2040,N_3078);
nand U5478 (N_5478,N_3314,N_2771);
or U5479 (N_5479,N_3858,N_2106);
nor U5480 (N_5480,N_3040,N_2207);
nor U5481 (N_5481,N_3555,N_2776);
or U5482 (N_5482,N_2623,N_3407);
nand U5483 (N_5483,N_2760,N_2745);
or U5484 (N_5484,N_2981,N_2211);
or U5485 (N_5485,N_3887,N_3577);
nor U5486 (N_5486,N_2933,N_2647);
nand U5487 (N_5487,N_2383,N_2549);
nand U5488 (N_5488,N_2497,N_2629);
or U5489 (N_5489,N_3988,N_2091);
nand U5490 (N_5490,N_3193,N_3881);
or U5491 (N_5491,N_3516,N_3947);
nand U5492 (N_5492,N_3747,N_3559);
and U5493 (N_5493,N_3108,N_3256);
nand U5494 (N_5494,N_3026,N_3999);
and U5495 (N_5495,N_3557,N_2799);
nand U5496 (N_5496,N_2099,N_2771);
and U5497 (N_5497,N_3859,N_2838);
or U5498 (N_5498,N_2616,N_2051);
nand U5499 (N_5499,N_2751,N_2781);
nor U5500 (N_5500,N_2682,N_3401);
nand U5501 (N_5501,N_3792,N_2886);
nand U5502 (N_5502,N_2658,N_2146);
nor U5503 (N_5503,N_2330,N_3231);
and U5504 (N_5504,N_2854,N_3218);
or U5505 (N_5505,N_2030,N_3987);
and U5506 (N_5506,N_3961,N_2161);
nand U5507 (N_5507,N_2081,N_2680);
and U5508 (N_5508,N_2178,N_3841);
or U5509 (N_5509,N_2214,N_2395);
and U5510 (N_5510,N_2267,N_2187);
nand U5511 (N_5511,N_2522,N_2264);
nand U5512 (N_5512,N_3325,N_3618);
nor U5513 (N_5513,N_3701,N_2810);
and U5514 (N_5514,N_3241,N_3570);
nand U5515 (N_5515,N_2211,N_3581);
nor U5516 (N_5516,N_2185,N_2239);
nand U5517 (N_5517,N_3390,N_2291);
nor U5518 (N_5518,N_3834,N_3564);
nand U5519 (N_5519,N_2488,N_3030);
or U5520 (N_5520,N_2645,N_2098);
or U5521 (N_5521,N_3395,N_2267);
or U5522 (N_5522,N_2324,N_2242);
or U5523 (N_5523,N_3641,N_3409);
nand U5524 (N_5524,N_2716,N_3683);
nor U5525 (N_5525,N_3473,N_3772);
nor U5526 (N_5526,N_2183,N_2872);
nand U5527 (N_5527,N_2628,N_3998);
and U5528 (N_5528,N_3755,N_2167);
and U5529 (N_5529,N_3040,N_2263);
or U5530 (N_5530,N_3901,N_3252);
nand U5531 (N_5531,N_3487,N_3074);
nor U5532 (N_5532,N_2207,N_2613);
nand U5533 (N_5533,N_2102,N_2107);
and U5534 (N_5534,N_2015,N_2431);
and U5535 (N_5535,N_3662,N_3172);
nand U5536 (N_5536,N_3255,N_3431);
nor U5537 (N_5537,N_3040,N_2907);
or U5538 (N_5538,N_2135,N_3588);
and U5539 (N_5539,N_3889,N_3702);
and U5540 (N_5540,N_3602,N_2828);
nor U5541 (N_5541,N_2822,N_2939);
or U5542 (N_5542,N_3045,N_3752);
nand U5543 (N_5543,N_2236,N_2399);
or U5544 (N_5544,N_2124,N_3194);
or U5545 (N_5545,N_2721,N_2965);
xor U5546 (N_5546,N_2376,N_3539);
and U5547 (N_5547,N_2894,N_2506);
or U5548 (N_5548,N_2729,N_3296);
xor U5549 (N_5549,N_2181,N_3517);
nand U5550 (N_5550,N_3452,N_3646);
or U5551 (N_5551,N_2579,N_3188);
and U5552 (N_5552,N_3433,N_2846);
or U5553 (N_5553,N_3001,N_3006);
nand U5554 (N_5554,N_3922,N_3319);
and U5555 (N_5555,N_3371,N_3150);
or U5556 (N_5556,N_3244,N_3060);
and U5557 (N_5557,N_2086,N_2776);
or U5558 (N_5558,N_2759,N_2599);
nor U5559 (N_5559,N_3458,N_2013);
and U5560 (N_5560,N_3562,N_2032);
and U5561 (N_5561,N_3242,N_2103);
and U5562 (N_5562,N_3724,N_2449);
nand U5563 (N_5563,N_2221,N_2605);
nand U5564 (N_5564,N_2006,N_3651);
and U5565 (N_5565,N_3981,N_2488);
and U5566 (N_5566,N_3334,N_3705);
or U5567 (N_5567,N_2332,N_2249);
nor U5568 (N_5568,N_3026,N_2275);
or U5569 (N_5569,N_3958,N_3714);
or U5570 (N_5570,N_2564,N_3989);
and U5571 (N_5571,N_3693,N_3776);
nand U5572 (N_5572,N_2041,N_2853);
nand U5573 (N_5573,N_2983,N_3138);
and U5574 (N_5574,N_3463,N_2703);
and U5575 (N_5575,N_3490,N_3156);
nand U5576 (N_5576,N_3326,N_3933);
or U5577 (N_5577,N_3466,N_2646);
or U5578 (N_5578,N_3945,N_3738);
nand U5579 (N_5579,N_3400,N_3885);
or U5580 (N_5580,N_3911,N_3146);
and U5581 (N_5581,N_3142,N_2791);
nand U5582 (N_5582,N_2681,N_3958);
nand U5583 (N_5583,N_2940,N_3152);
or U5584 (N_5584,N_2526,N_3932);
nor U5585 (N_5585,N_2959,N_2605);
or U5586 (N_5586,N_2903,N_3596);
nand U5587 (N_5587,N_2064,N_3651);
and U5588 (N_5588,N_3405,N_2409);
nor U5589 (N_5589,N_3747,N_3695);
nand U5590 (N_5590,N_2046,N_2390);
nand U5591 (N_5591,N_3457,N_2793);
nor U5592 (N_5592,N_3218,N_2464);
nor U5593 (N_5593,N_2772,N_2351);
or U5594 (N_5594,N_3024,N_3141);
nand U5595 (N_5595,N_2382,N_3286);
and U5596 (N_5596,N_3198,N_3894);
nand U5597 (N_5597,N_3212,N_2897);
or U5598 (N_5598,N_3320,N_3687);
or U5599 (N_5599,N_2327,N_3296);
and U5600 (N_5600,N_2496,N_3522);
nand U5601 (N_5601,N_3214,N_3521);
and U5602 (N_5602,N_3059,N_2687);
and U5603 (N_5603,N_2065,N_3715);
nand U5604 (N_5604,N_2587,N_3982);
nand U5605 (N_5605,N_2116,N_3484);
nand U5606 (N_5606,N_2401,N_3461);
nand U5607 (N_5607,N_2352,N_2035);
or U5608 (N_5608,N_2039,N_3084);
or U5609 (N_5609,N_3367,N_3142);
and U5610 (N_5610,N_2661,N_3015);
nor U5611 (N_5611,N_2624,N_3710);
and U5612 (N_5612,N_3227,N_2288);
and U5613 (N_5613,N_3367,N_2177);
and U5614 (N_5614,N_2221,N_2034);
nand U5615 (N_5615,N_2241,N_2416);
and U5616 (N_5616,N_2158,N_3378);
nor U5617 (N_5617,N_3643,N_3455);
nor U5618 (N_5618,N_3740,N_3806);
or U5619 (N_5619,N_3966,N_2838);
nor U5620 (N_5620,N_3852,N_3159);
nand U5621 (N_5621,N_2163,N_2446);
nand U5622 (N_5622,N_2539,N_3371);
nor U5623 (N_5623,N_3329,N_3782);
or U5624 (N_5624,N_2730,N_2663);
and U5625 (N_5625,N_2258,N_3486);
nand U5626 (N_5626,N_2179,N_3960);
or U5627 (N_5627,N_2013,N_3239);
nor U5628 (N_5628,N_3164,N_3794);
nand U5629 (N_5629,N_2911,N_2097);
or U5630 (N_5630,N_3885,N_3800);
nand U5631 (N_5631,N_2868,N_3078);
and U5632 (N_5632,N_2404,N_3273);
and U5633 (N_5633,N_2026,N_3349);
and U5634 (N_5634,N_3711,N_2601);
nor U5635 (N_5635,N_2046,N_3269);
nor U5636 (N_5636,N_3395,N_2389);
or U5637 (N_5637,N_3640,N_2422);
or U5638 (N_5638,N_2749,N_3935);
or U5639 (N_5639,N_2166,N_2849);
nand U5640 (N_5640,N_3966,N_2878);
and U5641 (N_5641,N_2728,N_3863);
and U5642 (N_5642,N_3728,N_2844);
nand U5643 (N_5643,N_3861,N_2629);
and U5644 (N_5644,N_3092,N_3179);
nor U5645 (N_5645,N_3086,N_3522);
or U5646 (N_5646,N_3382,N_3221);
or U5647 (N_5647,N_3918,N_2246);
or U5648 (N_5648,N_2774,N_3271);
or U5649 (N_5649,N_2625,N_3085);
nand U5650 (N_5650,N_3455,N_3146);
nor U5651 (N_5651,N_3131,N_2778);
or U5652 (N_5652,N_3468,N_2354);
or U5653 (N_5653,N_3352,N_3914);
nor U5654 (N_5654,N_2897,N_3566);
and U5655 (N_5655,N_3477,N_2333);
or U5656 (N_5656,N_3638,N_3045);
and U5657 (N_5657,N_3346,N_2780);
nand U5658 (N_5658,N_2004,N_3754);
or U5659 (N_5659,N_3323,N_2922);
or U5660 (N_5660,N_2293,N_2802);
nand U5661 (N_5661,N_3087,N_2512);
or U5662 (N_5662,N_3280,N_2979);
and U5663 (N_5663,N_3415,N_3256);
or U5664 (N_5664,N_2926,N_3225);
nand U5665 (N_5665,N_3398,N_2995);
and U5666 (N_5666,N_2602,N_2657);
and U5667 (N_5667,N_3068,N_3785);
nand U5668 (N_5668,N_2479,N_2011);
nand U5669 (N_5669,N_3743,N_3436);
nor U5670 (N_5670,N_3014,N_3666);
or U5671 (N_5671,N_3231,N_2752);
xnor U5672 (N_5672,N_2082,N_3475);
and U5673 (N_5673,N_2772,N_2185);
or U5674 (N_5674,N_2960,N_3487);
and U5675 (N_5675,N_2870,N_3619);
or U5676 (N_5676,N_3757,N_3482);
or U5677 (N_5677,N_2647,N_2847);
or U5678 (N_5678,N_2905,N_2058);
or U5679 (N_5679,N_3036,N_2496);
nor U5680 (N_5680,N_2198,N_2693);
nand U5681 (N_5681,N_2392,N_2854);
or U5682 (N_5682,N_3890,N_3709);
nand U5683 (N_5683,N_2991,N_2890);
nor U5684 (N_5684,N_3234,N_3159);
and U5685 (N_5685,N_2429,N_3969);
nor U5686 (N_5686,N_3975,N_3851);
nor U5687 (N_5687,N_2378,N_3086);
and U5688 (N_5688,N_3232,N_2271);
nand U5689 (N_5689,N_2428,N_2137);
xor U5690 (N_5690,N_2445,N_2051);
and U5691 (N_5691,N_2154,N_3183);
or U5692 (N_5692,N_2614,N_2330);
and U5693 (N_5693,N_2729,N_2253);
xnor U5694 (N_5694,N_3144,N_2262);
nor U5695 (N_5695,N_3473,N_2568);
nand U5696 (N_5696,N_3390,N_2399);
and U5697 (N_5697,N_2429,N_2120);
or U5698 (N_5698,N_3987,N_2508);
nor U5699 (N_5699,N_3986,N_2693);
or U5700 (N_5700,N_3495,N_2646);
nand U5701 (N_5701,N_3133,N_2872);
or U5702 (N_5702,N_3924,N_3941);
or U5703 (N_5703,N_3340,N_3726);
nor U5704 (N_5704,N_3884,N_2383);
and U5705 (N_5705,N_3987,N_2733);
or U5706 (N_5706,N_2328,N_2135);
nand U5707 (N_5707,N_2253,N_3365);
nand U5708 (N_5708,N_3542,N_3097);
and U5709 (N_5709,N_2604,N_3891);
xor U5710 (N_5710,N_3261,N_2619);
nor U5711 (N_5711,N_2271,N_2554);
nand U5712 (N_5712,N_2048,N_2544);
nand U5713 (N_5713,N_2443,N_3369);
or U5714 (N_5714,N_3640,N_3350);
and U5715 (N_5715,N_2834,N_3248);
or U5716 (N_5716,N_2839,N_3955);
nand U5717 (N_5717,N_3668,N_3269);
nor U5718 (N_5718,N_2659,N_2588);
and U5719 (N_5719,N_3112,N_2005);
nand U5720 (N_5720,N_3821,N_2977);
and U5721 (N_5721,N_3727,N_3114);
nor U5722 (N_5722,N_3852,N_2792);
nor U5723 (N_5723,N_3359,N_2427);
nand U5724 (N_5724,N_2480,N_2981);
nor U5725 (N_5725,N_2409,N_2558);
nand U5726 (N_5726,N_3361,N_3080);
and U5727 (N_5727,N_3468,N_2868);
or U5728 (N_5728,N_3834,N_2735);
and U5729 (N_5729,N_2997,N_2974);
and U5730 (N_5730,N_2670,N_3108);
nand U5731 (N_5731,N_3870,N_3866);
and U5732 (N_5732,N_2192,N_3925);
nor U5733 (N_5733,N_3163,N_2629);
nand U5734 (N_5734,N_2387,N_2242);
nor U5735 (N_5735,N_3238,N_2513);
nand U5736 (N_5736,N_3303,N_2385);
nor U5737 (N_5737,N_3090,N_2993);
nor U5738 (N_5738,N_3004,N_2274);
nand U5739 (N_5739,N_2231,N_2512);
nor U5740 (N_5740,N_2798,N_2284);
or U5741 (N_5741,N_2235,N_2886);
nor U5742 (N_5742,N_2003,N_2266);
nor U5743 (N_5743,N_2937,N_3197);
and U5744 (N_5744,N_2864,N_3422);
or U5745 (N_5745,N_3681,N_3822);
xnor U5746 (N_5746,N_2617,N_3320);
or U5747 (N_5747,N_3974,N_3073);
nor U5748 (N_5748,N_2540,N_3404);
nor U5749 (N_5749,N_3489,N_2711);
and U5750 (N_5750,N_2196,N_2613);
nand U5751 (N_5751,N_2348,N_3528);
or U5752 (N_5752,N_3448,N_3368);
nor U5753 (N_5753,N_2093,N_2832);
xnor U5754 (N_5754,N_3577,N_3920);
and U5755 (N_5755,N_2770,N_2695);
and U5756 (N_5756,N_3454,N_3711);
nand U5757 (N_5757,N_2680,N_2897);
and U5758 (N_5758,N_2947,N_2780);
nor U5759 (N_5759,N_2412,N_3029);
nor U5760 (N_5760,N_3987,N_3503);
or U5761 (N_5761,N_2537,N_3875);
xor U5762 (N_5762,N_3037,N_3955);
or U5763 (N_5763,N_2934,N_3852);
and U5764 (N_5764,N_3118,N_3582);
nor U5765 (N_5765,N_2871,N_2710);
nand U5766 (N_5766,N_3540,N_2200);
nand U5767 (N_5767,N_3122,N_2336);
or U5768 (N_5768,N_2958,N_3433);
nand U5769 (N_5769,N_3641,N_3109);
nand U5770 (N_5770,N_3791,N_2300);
nand U5771 (N_5771,N_3436,N_3111);
and U5772 (N_5772,N_3542,N_3243);
nor U5773 (N_5773,N_2079,N_3155);
or U5774 (N_5774,N_3506,N_3065);
nor U5775 (N_5775,N_2969,N_2995);
nor U5776 (N_5776,N_2493,N_2106);
or U5777 (N_5777,N_2454,N_2376);
nor U5778 (N_5778,N_2330,N_3244);
or U5779 (N_5779,N_3947,N_3562);
nor U5780 (N_5780,N_2104,N_2112);
nor U5781 (N_5781,N_2818,N_2715);
or U5782 (N_5782,N_2180,N_2717);
and U5783 (N_5783,N_3434,N_3612);
or U5784 (N_5784,N_3606,N_3728);
nor U5785 (N_5785,N_3729,N_2075);
and U5786 (N_5786,N_3945,N_3404);
nand U5787 (N_5787,N_2547,N_3840);
nand U5788 (N_5788,N_3999,N_2839);
nand U5789 (N_5789,N_2290,N_2544);
and U5790 (N_5790,N_3243,N_2270);
nand U5791 (N_5791,N_3873,N_2349);
and U5792 (N_5792,N_3011,N_2859);
or U5793 (N_5793,N_3931,N_3433);
nor U5794 (N_5794,N_2509,N_3360);
nor U5795 (N_5795,N_3720,N_3669);
and U5796 (N_5796,N_2802,N_2663);
nor U5797 (N_5797,N_2483,N_2957);
nand U5798 (N_5798,N_3937,N_2468);
nand U5799 (N_5799,N_3252,N_2014);
and U5800 (N_5800,N_3538,N_3328);
and U5801 (N_5801,N_2636,N_2876);
or U5802 (N_5802,N_3201,N_2521);
or U5803 (N_5803,N_3430,N_2333);
nand U5804 (N_5804,N_3633,N_2082);
or U5805 (N_5805,N_3161,N_3855);
or U5806 (N_5806,N_2168,N_3417);
nand U5807 (N_5807,N_3940,N_3915);
nor U5808 (N_5808,N_2083,N_2608);
or U5809 (N_5809,N_2565,N_2455);
and U5810 (N_5810,N_3870,N_3958);
or U5811 (N_5811,N_2500,N_2770);
or U5812 (N_5812,N_2180,N_3851);
or U5813 (N_5813,N_2001,N_2971);
and U5814 (N_5814,N_3015,N_3008);
or U5815 (N_5815,N_3441,N_2241);
nor U5816 (N_5816,N_2107,N_2453);
or U5817 (N_5817,N_3585,N_2443);
and U5818 (N_5818,N_2484,N_2591);
nand U5819 (N_5819,N_2566,N_2247);
nand U5820 (N_5820,N_2024,N_3376);
xor U5821 (N_5821,N_2333,N_3150);
or U5822 (N_5822,N_3103,N_3880);
or U5823 (N_5823,N_2232,N_2015);
nor U5824 (N_5824,N_3356,N_3161);
or U5825 (N_5825,N_3778,N_2642);
or U5826 (N_5826,N_2770,N_2482);
nor U5827 (N_5827,N_3279,N_2260);
nor U5828 (N_5828,N_3351,N_2763);
xnor U5829 (N_5829,N_2238,N_2419);
or U5830 (N_5830,N_2495,N_3244);
or U5831 (N_5831,N_2316,N_3456);
and U5832 (N_5832,N_2546,N_3335);
nor U5833 (N_5833,N_3862,N_3231);
nor U5834 (N_5834,N_2082,N_3339);
or U5835 (N_5835,N_3838,N_3985);
or U5836 (N_5836,N_3045,N_2631);
nand U5837 (N_5837,N_2222,N_2081);
or U5838 (N_5838,N_2862,N_3782);
nand U5839 (N_5839,N_3190,N_2739);
nand U5840 (N_5840,N_3139,N_2767);
and U5841 (N_5841,N_3947,N_3344);
and U5842 (N_5842,N_2020,N_2037);
nand U5843 (N_5843,N_3860,N_2726);
and U5844 (N_5844,N_2733,N_2920);
or U5845 (N_5845,N_3850,N_3858);
nor U5846 (N_5846,N_3810,N_2294);
or U5847 (N_5847,N_3522,N_3519);
and U5848 (N_5848,N_2700,N_3138);
and U5849 (N_5849,N_3977,N_2037);
or U5850 (N_5850,N_3059,N_2782);
and U5851 (N_5851,N_2919,N_2400);
and U5852 (N_5852,N_2452,N_3915);
and U5853 (N_5853,N_3348,N_3565);
or U5854 (N_5854,N_2647,N_2673);
nand U5855 (N_5855,N_3557,N_3440);
nand U5856 (N_5856,N_3536,N_2472);
nor U5857 (N_5857,N_3554,N_3014);
and U5858 (N_5858,N_2938,N_3667);
or U5859 (N_5859,N_3341,N_3397);
nor U5860 (N_5860,N_2768,N_2473);
nor U5861 (N_5861,N_3502,N_3923);
nor U5862 (N_5862,N_3940,N_3164);
xnor U5863 (N_5863,N_3398,N_3251);
or U5864 (N_5864,N_3966,N_2134);
or U5865 (N_5865,N_3786,N_3737);
nor U5866 (N_5866,N_2603,N_3697);
nor U5867 (N_5867,N_2700,N_2051);
and U5868 (N_5868,N_2839,N_2661);
nor U5869 (N_5869,N_3712,N_3803);
nor U5870 (N_5870,N_3790,N_3886);
nor U5871 (N_5871,N_3848,N_3608);
or U5872 (N_5872,N_3201,N_3316);
and U5873 (N_5873,N_2580,N_3901);
or U5874 (N_5874,N_2657,N_3096);
nand U5875 (N_5875,N_3996,N_3124);
and U5876 (N_5876,N_2216,N_2388);
or U5877 (N_5877,N_2613,N_3626);
or U5878 (N_5878,N_3635,N_2001);
or U5879 (N_5879,N_2052,N_2768);
and U5880 (N_5880,N_3419,N_3193);
nand U5881 (N_5881,N_2793,N_2641);
and U5882 (N_5882,N_2535,N_3957);
and U5883 (N_5883,N_2700,N_2671);
nand U5884 (N_5884,N_2938,N_2726);
nand U5885 (N_5885,N_3298,N_3701);
nand U5886 (N_5886,N_3761,N_3149);
nor U5887 (N_5887,N_3729,N_3494);
nand U5888 (N_5888,N_3174,N_3818);
nor U5889 (N_5889,N_2582,N_2201);
nor U5890 (N_5890,N_3795,N_2188);
and U5891 (N_5891,N_3552,N_2864);
xnor U5892 (N_5892,N_2045,N_3349);
nand U5893 (N_5893,N_3049,N_2046);
nand U5894 (N_5894,N_2234,N_3252);
and U5895 (N_5895,N_2160,N_3325);
or U5896 (N_5896,N_3812,N_2877);
or U5897 (N_5897,N_3291,N_2208);
or U5898 (N_5898,N_3044,N_2055);
and U5899 (N_5899,N_3574,N_3412);
or U5900 (N_5900,N_3431,N_3251);
and U5901 (N_5901,N_2423,N_2087);
nor U5902 (N_5902,N_3338,N_2578);
nand U5903 (N_5903,N_3431,N_2838);
xor U5904 (N_5904,N_2261,N_2390);
nand U5905 (N_5905,N_2519,N_2437);
or U5906 (N_5906,N_2971,N_2089);
or U5907 (N_5907,N_3127,N_2743);
and U5908 (N_5908,N_3677,N_3583);
nor U5909 (N_5909,N_3302,N_3080);
nor U5910 (N_5910,N_3443,N_2761);
nor U5911 (N_5911,N_2303,N_2390);
nand U5912 (N_5912,N_3539,N_2490);
or U5913 (N_5913,N_2725,N_3813);
xnor U5914 (N_5914,N_2728,N_2544);
nand U5915 (N_5915,N_2385,N_2422);
and U5916 (N_5916,N_3586,N_3759);
and U5917 (N_5917,N_2261,N_3347);
and U5918 (N_5918,N_3485,N_2733);
nor U5919 (N_5919,N_2506,N_3560);
and U5920 (N_5920,N_2789,N_2892);
and U5921 (N_5921,N_3141,N_2744);
or U5922 (N_5922,N_2352,N_2554);
nor U5923 (N_5923,N_2169,N_3553);
and U5924 (N_5924,N_2076,N_3736);
nand U5925 (N_5925,N_2281,N_2119);
nand U5926 (N_5926,N_3466,N_2409);
nand U5927 (N_5927,N_2333,N_2561);
and U5928 (N_5928,N_3240,N_3421);
nand U5929 (N_5929,N_3002,N_3825);
nand U5930 (N_5930,N_2728,N_3699);
nand U5931 (N_5931,N_2563,N_2309);
or U5932 (N_5932,N_2856,N_2909);
and U5933 (N_5933,N_3206,N_2689);
nor U5934 (N_5934,N_2192,N_2823);
nor U5935 (N_5935,N_3114,N_3127);
nor U5936 (N_5936,N_2949,N_2729);
nor U5937 (N_5937,N_3640,N_3564);
and U5938 (N_5938,N_3607,N_2855);
nand U5939 (N_5939,N_3419,N_3517);
xnor U5940 (N_5940,N_2520,N_3634);
nor U5941 (N_5941,N_3109,N_3576);
and U5942 (N_5942,N_2817,N_3431);
or U5943 (N_5943,N_3708,N_2486);
nor U5944 (N_5944,N_2633,N_2556);
xnor U5945 (N_5945,N_3808,N_3322);
xor U5946 (N_5946,N_2513,N_3342);
nand U5947 (N_5947,N_2090,N_2413);
and U5948 (N_5948,N_2130,N_2904);
nand U5949 (N_5949,N_3436,N_2119);
nand U5950 (N_5950,N_2801,N_2348);
nor U5951 (N_5951,N_3734,N_2218);
or U5952 (N_5952,N_2433,N_3747);
nor U5953 (N_5953,N_3434,N_3606);
nand U5954 (N_5954,N_3177,N_2472);
nand U5955 (N_5955,N_3619,N_3892);
nor U5956 (N_5956,N_3444,N_2320);
nor U5957 (N_5957,N_3482,N_3456);
nand U5958 (N_5958,N_2329,N_3327);
and U5959 (N_5959,N_2102,N_2981);
and U5960 (N_5960,N_3075,N_2616);
nor U5961 (N_5961,N_2461,N_2371);
and U5962 (N_5962,N_3313,N_3042);
nor U5963 (N_5963,N_3043,N_3133);
nand U5964 (N_5964,N_3256,N_3571);
nand U5965 (N_5965,N_2063,N_3936);
or U5966 (N_5966,N_3163,N_3454);
and U5967 (N_5967,N_2025,N_2264);
and U5968 (N_5968,N_2473,N_3674);
and U5969 (N_5969,N_2249,N_2386);
and U5970 (N_5970,N_3687,N_2557);
or U5971 (N_5971,N_3375,N_2408);
nand U5972 (N_5972,N_2061,N_2878);
nor U5973 (N_5973,N_3549,N_3794);
or U5974 (N_5974,N_3567,N_2542);
nand U5975 (N_5975,N_3821,N_2021);
xor U5976 (N_5976,N_2924,N_3825);
and U5977 (N_5977,N_3041,N_2263);
nand U5978 (N_5978,N_3983,N_2258);
nand U5979 (N_5979,N_3330,N_2085);
nand U5980 (N_5980,N_3622,N_2064);
and U5981 (N_5981,N_2958,N_2154);
and U5982 (N_5982,N_3531,N_3331);
and U5983 (N_5983,N_2663,N_2075);
or U5984 (N_5984,N_2394,N_2258);
or U5985 (N_5985,N_2716,N_2890);
nor U5986 (N_5986,N_3347,N_2098);
or U5987 (N_5987,N_3166,N_3303);
and U5988 (N_5988,N_3894,N_3310);
nor U5989 (N_5989,N_2301,N_2127);
or U5990 (N_5990,N_2990,N_2408);
or U5991 (N_5991,N_3613,N_2204);
and U5992 (N_5992,N_3433,N_2446);
xor U5993 (N_5993,N_2265,N_3794);
nor U5994 (N_5994,N_3928,N_3726);
or U5995 (N_5995,N_3657,N_3146);
nor U5996 (N_5996,N_3499,N_2696);
and U5997 (N_5997,N_2686,N_3176);
and U5998 (N_5998,N_3592,N_3989);
nand U5999 (N_5999,N_2813,N_3714);
and U6000 (N_6000,N_5860,N_5543);
or U6001 (N_6001,N_5289,N_5343);
and U6002 (N_6002,N_5191,N_5951);
and U6003 (N_6003,N_4258,N_4180);
nand U6004 (N_6004,N_4315,N_5979);
or U6005 (N_6005,N_4555,N_4221);
nor U6006 (N_6006,N_5356,N_4954);
or U6007 (N_6007,N_5901,N_4909);
nor U6008 (N_6008,N_5863,N_5928);
nand U6009 (N_6009,N_4865,N_4862);
or U6010 (N_6010,N_4235,N_4592);
nand U6011 (N_6011,N_4553,N_5568);
nand U6012 (N_6012,N_4433,N_4847);
and U6013 (N_6013,N_4532,N_5910);
nor U6014 (N_6014,N_5023,N_4836);
and U6015 (N_6015,N_5763,N_5911);
xnor U6016 (N_6016,N_5809,N_5913);
and U6017 (N_6017,N_4947,N_4222);
nand U6018 (N_6018,N_4844,N_4062);
or U6019 (N_6019,N_4666,N_5485);
nor U6020 (N_6020,N_4458,N_5796);
xor U6021 (N_6021,N_4241,N_5790);
or U6022 (N_6022,N_4242,N_5243);
nand U6023 (N_6023,N_4394,N_4145);
xnor U6024 (N_6024,N_4245,N_4340);
nor U6025 (N_6025,N_4653,N_4013);
nor U6026 (N_6026,N_5434,N_5750);
and U6027 (N_6027,N_4372,N_4711);
or U6028 (N_6028,N_4169,N_4330);
and U6029 (N_6029,N_4705,N_4057);
or U6030 (N_6030,N_5521,N_5772);
and U6031 (N_6031,N_4318,N_5257);
or U6032 (N_6032,N_5031,N_4132);
nand U6033 (N_6033,N_4359,N_4485);
and U6034 (N_6034,N_4370,N_5037);
and U6035 (N_6035,N_4030,N_5898);
and U6036 (N_6036,N_4917,N_4515);
or U6037 (N_6037,N_5060,N_4595);
xor U6038 (N_6038,N_4938,N_5161);
and U6039 (N_6039,N_4829,N_5514);
and U6040 (N_6040,N_5725,N_5964);
nor U6041 (N_6041,N_4498,N_5841);
or U6042 (N_6042,N_5154,N_5696);
nand U6043 (N_6043,N_4767,N_5574);
nor U6044 (N_6044,N_4792,N_4183);
xnor U6045 (N_6045,N_4197,N_4546);
or U6046 (N_6046,N_5094,N_5525);
nor U6047 (N_6047,N_5312,N_5535);
nor U6048 (N_6048,N_5032,N_5739);
nor U6049 (N_6049,N_4682,N_5091);
or U6050 (N_6050,N_5275,N_5782);
nand U6051 (N_6051,N_4224,N_5516);
and U6052 (N_6052,N_4193,N_5666);
and U6053 (N_6053,N_5127,N_5384);
and U6054 (N_6054,N_5987,N_5217);
nand U6055 (N_6055,N_5152,N_5677);
xnor U6056 (N_6056,N_5184,N_4487);
nor U6057 (N_6057,N_4860,N_4200);
nand U6058 (N_6058,N_5416,N_4087);
and U6059 (N_6059,N_5661,N_4869);
nor U6060 (N_6060,N_5311,N_4150);
nand U6061 (N_6061,N_5998,N_5952);
nor U6062 (N_6062,N_5675,N_4575);
or U6063 (N_6063,N_4082,N_4143);
nor U6064 (N_6064,N_4730,N_5232);
nand U6065 (N_6065,N_5051,N_4760);
nand U6066 (N_6066,N_4067,N_4376);
nor U6067 (N_6067,N_4771,N_5728);
xor U6068 (N_6068,N_4078,N_5945);
nand U6069 (N_6069,N_4535,N_4616);
nand U6070 (N_6070,N_4636,N_4809);
nor U6071 (N_6071,N_4548,N_5837);
or U6072 (N_6072,N_5590,N_5242);
and U6073 (N_6073,N_4746,N_5269);
and U6074 (N_6074,N_5629,N_5102);
nor U6075 (N_6075,N_5918,N_4022);
or U6076 (N_6076,N_5764,N_5547);
nand U6077 (N_6077,N_4513,N_5592);
and U6078 (N_6078,N_4001,N_4483);
nand U6079 (N_6079,N_5749,N_5756);
nand U6080 (N_6080,N_5671,N_5271);
nand U6081 (N_6081,N_5062,N_5386);
nand U6082 (N_6082,N_5167,N_5417);
xor U6083 (N_6083,N_4131,N_4419);
xor U6084 (N_6084,N_5930,N_4605);
nor U6085 (N_6085,N_4570,N_4770);
nor U6086 (N_6086,N_4048,N_4630);
nand U6087 (N_6087,N_5787,N_4851);
nor U6088 (N_6088,N_5747,N_5720);
or U6089 (N_6089,N_5919,N_5971);
or U6090 (N_6090,N_5850,N_5385);
nor U6091 (N_6091,N_4945,N_5178);
nor U6092 (N_6092,N_5393,N_4294);
nand U6093 (N_6093,N_5105,N_4686);
nor U6094 (N_6094,N_5172,N_4953);
nor U6095 (N_6095,N_4644,N_4537);
nand U6096 (N_6096,N_4872,N_5812);
nand U6097 (N_6097,N_4657,N_5006);
and U6098 (N_6098,N_4218,N_5757);
or U6099 (N_6099,N_5294,N_5447);
nand U6100 (N_6100,N_4454,N_4597);
xnor U6101 (N_6101,N_4337,N_5843);
xnor U6102 (N_6102,N_4873,N_5323);
xnor U6103 (N_6103,N_5050,N_4698);
or U6104 (N_6104,N_5865,N_5745);
nor U6105 (N_6105,N_5231,N_5605);
or U6106 (N_6106,N_5025,N_4288);
and U6107 (N_6107,N_4501,N_5609);
or U6108 (N_6108,N_4772,N_5559);
xnor U6109 (N_6109,N_4503,N_4747);
and U6110 (N_6110,N_5528,N_4237);
nand U6111 (N_6111,N_5362,N_4021);
nand U6112 (N_6112,N_4144,N_5140);
nand U6113 (N_6113,N_4257,N_5679);
nand U6114 (N_6114,N_5372,N_5943);
or U6115 (N_6115,N_4940,N_5755);
nand U6116 (N_6116,N_5292,N_4684);
nand U6117 (N_6117,N_5807,N_4217);
nand U6118 (N_6118,N_5531,N_5098);
and U6119 (N_6119,N_4070,N_5880);
or U6120 (N_6120,N_4734,N_5299);
nor U6121 (N_6121,N_5821,N_5280);
nor U6122 (N_6122,N_4027,N_4750);
and U6123 (N_6123,N_4282,N_5282);
nand U6124 (N_6124,N_5538,N_4528);
and U6125 (N_6125,N_4065,N_5746);
nand U6126 (N_6126,N_4480,N_5578);
xnor U6127 (N_6127,N_4691,N_5293);
nor U6128 (N_6128,N_5955,N_4488);
nor U6129 (N_6129,N_4439,N_4960);
nand U6130 (N_6130,N_5001,N_4081);
nor U6131 (N_6131,N_5138,N_4898);
or U6132 (N_6132,N_4171,N_5460);
or U6133 (N_6133,N_4252,N_4277);
and U6134 (N_6134,N_5478,N_5129);
or U6135 (N_6135,N_4669,N_5148);
nor U6136 (N_6136,N_4739,N_5123);
and U6137 (N_6137,N_4588,N_5897);
or U6138 (N_6138,N_5683,N_4060);
or U6139 (N_6139,N_5741,N_5177);
and U6140 (N_6140,N_4357,N_5207);
or U6141 (N_6141,N_5237,N_4915);
and U6142 (N_6142,N_4789,N_5156);
nand U6143 (N_6143,N_4606,N_4253);
or U6144 (N_6144,N_4598,N_4331);
and U6145 (N_6145,N_5892,N_5501);
xor U6146 (N_6146,N_5228,N_5260);
nand U6147 (N_6147,N_4895,N_4857);
nor U6148 (N_6148,N_5249,N_5277);
or U6149 (N_6149,N_5017,N_5470);
and U6150 (N_6150,N_4828,N_4977);
and U6151 (N_6151,N_4525,N_4026);
nor U6152 (N_6152,N_5718,N_4929);
and U6153 (N_6153,N_4692,N_5014);
and U6154 (N_6154,N_4207,N_5404);
nor U6155 (N_6155,N_5084,N_5942);
and U6156 (N_6156,N_5099,N_5400);
and U6157 (N_6157,N_5097,N_4834);
and U6158 (N_6158,N_4516,N_4609);
or U6159 (N_6159,N_4325,N_4976);
nor U6160 (N_6160,N_4910,N_5043);
or U6161 (N_6161,N_5110,N_4924);
nand U6162 (N_6162,N_5168,N_5137);
or U6163 (N_6163,N_5296,N_4293);
or U6164 (N_6164,N_4071,N_4349);
nand U6165 (N_6165,N_4385,N_5413);
and U6166 (N_6166,N_5706,N_4538);
or U6167 (N_6167,N_4858,N_4648);
nand U6168 (N_6168,N_4335,N_4461);
nand U6169 (N_6169,N_5676,N_4264);
or U6170 (N_6170,N_5507,N_5702);
nand U6171 (N_6171,N_5786,N_4414);
nand U6172 (N_6172,N_5358,N_4974);
or U6173 (N_6173,N_4754,N_5414);
xnor U6174 (N_6174,N_5357,N_5007);
nand U6175 (N_6175,N_5151,N_5370);
nand U6176 (N_6176,N_5922,N_4526);
nor U6177 (N_6177,N_4391,N_4967);
xor U6178 (N_6178,N_4378,N_4901);
nor U6179 (N_6179,N_4761,N_5195);
nand U6180 (N_6180,N_4527,N_5585);
or U6181 (N_6181,N_5399,N_4107);
nor U6182 (N_6182,N_5854,N_4384);
or U6183 (N_6183,N_4499,N_4659);
nor U6184 (N_6184,N_4808,N_5618);
nor U6185 (N_6185,N_4326,N_4640);
or U6186 (N_6186,N_5405,N_5208);
nand U6187 (N_6187,N_4741,N_5363);
nor U6188 (N_6188,N_4662,N_5375);
and U6189 (N_6189,N_5831,N_5754);
nand U6190 (N_6190,N_4531,N_4854);
nand U6191 (N_6191,N_5803,N_5588);
nand U6192 (N_6192,N_4676,N_4032);
nor U6193 (N_6193,N_5496,N_4776);
or U6194 (N_6194,N_5354,N_5466);
nor U6195 (N_6195,N_5144,N_4208);
nor U6196 (N_6196,N_4382,N_4569);
nor U6197 (N_6197,N_4165,N_5817);
and U6198 (N_6198,N_5814,N_5233);
nor U6199 (N_6199,N_5864,N_4003);
nor U6200 (N_6200,N_4448,N_4113);
nor U6201 (N_6201,N_5111,N_4424);
and U6202 (N_6202,N_5201,N_4423);
and U6203 (N_6203,N_5638,N_4647);
nand U6204 (N_6204,N_5518,N_4817);
and U6205 (N_6205,N_5502,N_5439);
or U6206 (N_6206,N_4756,N_5853);
or U6207 (N_6207,N_4556,N_5934);
and U6208 (N_6208,N_4796,N_4846);
nor U6209 (N_6209,N_5488,N_5121);
and U6210 (N_6210,N_5779,N_4281);
nor U6211 (N_6211,N_4276,N_4261);
and U6212 (N_6212,N_5135,N_5164);
and U6213 (N_6213,N_4823,N_5455);
nor U6214 (N_6214,N_4395,N_5879);
or U6215 (N_6215,N_5010,N_4763);
nor U6216 (N_6216,N_4280,N_5364);
nand U6217 (N_6217,N_5956,N_5262);
or U6218 (N_6218,N_5020,N_5438);
or U6219 (N_6219,N_5132,N_5141);
and U6220 (N_6220,N_4352,N_5458);
or U6221 (N_6221,N_4742,N_5722);
nor U6222 (N_6222,N_5199,N_4008);
and U6223 (N_6223,N_4757,N_5183);
nand U6224 (N_6224,N_5691,N_4540);
nor U6225 (N_6225,N_4453,N_5421);
and U6226 (N_6226,N_4185,N_4184);
or U6227 (N_6227,N_5113,N_5092);
and U6228 (N_6228,N_5142,N_4274);
nor U6229 (N_6229,N_5089,N_5390);
and U6230 (N_6230,N_4520,N_5035);
nor U6231 (N_6231,N_4468,N_5347);
nor U6232 (N_6232,N_4043,N_5459);
xnor U6233 (N_6233,N_5244,N_5048);
nand U6234 (N_6234,N_4225,N_5895);
or U6235 (N_6235,N_5255,N_5622);
nor U6236 (N_6236,N_4627,N_5916);
and U6237 (N_6237,N_5729,N_4351);
and U6238 (N_6238,N_4713,N_4421);
nor U6239 (N_6239,N_4524,N_5371);
and U6240 (N_6240,N_5506,N_5068);
nor U6241 (N_6241,N_4130,N_5334);
xnor U6242 (N_6242,N_4700,N_5019);
nand U6243 (N_6243,N_4311,N_4289);
or U6244 (N_6244,N_5071,N_5200);
nand U6245 (N_6245,N_5862,N_4736);
or U6246 (N_6246,N_5038,N_4667);
nor U6247 (N_6247,N_4164,N_4016);
xnor U6248 (N_6248,N_4426,N_5561);
xnor U6249 (N_6249,N_4919,N_4024);
and U6250 (N_6250,N_4363,N_5569);
nand U6251 (N_6251,N_5418,N_4079);
nand U6252 (N_6252,N_5659,N_5811);
nand U6253 (N_6253,N_5155,N_5572);
and U6254 (N_6254,N_4220,N_5997);
nor U6255 (N_6255,N_5361,N_4913);
nand U6256 (N_6256,N_5326,N_4500);
nor U6257 (N_6257,N_4621,N_4589);
nand U6258 (N_6258,N_4308,N_5077);
nor U6259 (N_6259,N_4459,N_4434);
nand U6260 (N_6260,N_4074,N_4090);
nor U6261 (N_6261,N_5824,N_5925);
nor U6262 (N_6262,N_5229,N_4066);
or U6263 (N_6263,N_5454,N_4989);
nand U6264 (N_6264,N_4886,N_4018);
or U6265 (N_6265,N_5224,N_5285);
or U6266 (N_6266,N_4852,N_5662);
and U6267 (N_6267,N_5991,N_5833);
or U6268 (N_6268,N_5394,N_5214);
nand U6269 (N_6269,N_5461,N_5548);
and U6270 (N_6270,N_5192,N_5339);
or U6271 (N_6271,N_4802,N_4804);
nor U6272 (N_6272,N_4505,N_4701);
and U6273 (N_6273,N_5189,N_4558);
nand U6274 (N_6274,N_5594,N_4951);
or U6275 (N_6275,N_4878,N_4190);
nor U6276 (N_6276,N_5909,N_4464);
nand U6277 (N_6277,N_5623,N_4273);
nor U6278 (N_6278,N_4477,N_4342);
and U6279 (N_6279,N_4715,N_4830);
and U6280 (N_6280,N_4336,N_4455);
nor U6281 (N_6281,N_4702,N_4658);
nand U6282 (N_6282,N_5389,N_4722);
nor U6283 (N_6283,N_4029,N_5408);
nand U6284 (N_6284,N_5477,N_5036);
nand U6285 (N_6285,N_4663,N_4046);
nand U6286 (N_6286,N_4321,N_5867);
and U6287 (N_6287,N_5387,N_4853);
nor U6288 (N_6288,N_4914,N_5999);
nor U6289 (N_6289,N_5027,N_4995);
or U6290 (N_6290,N_4610,N_5655);
nand U6291 (N_6291,N_4568,N_5436);
nand U6292 (N_6292,N_5877,N_5567);
nand U6293 (N_6293,N_5171,N_4720);
nor U6294 (N_6294,N_4354,N_5963);
or U6295 (N_6295,N_4086,N_5090);
or U6296 (N_6296,N_5197,N_4660);
nor U6297 (N_6297,N_5883,N_4920);
or U6298 (N_6298,N_4213,N_5440);
or U6299 (N_6299,N_5643,N_5205);
and U6300 (N_6300,N_5773,N_4907);
nor U6301 (N_6301,N_4023,N_5975);
nor U6302 (N_6302,N_5522,N_4324);
or U6303 (N_6303,N_4814,N_4155);
and U6304 (N_6304,N_4894,N_5226);
and U6305 (N_6305,N_5861,N_5256);
nor U6306 (N_6306,N_5391,N_4069);
nor U6307 (N_6307,N_4020,N_5279);
nand U6308 (N_6308,N_5733,N_4380);
or U6309 (N_6309,N_5838,N_5815);
nor U6310 (N_6310,N_4752,N_5519);
or U6311 (N_6311,N_4406,N_4843);
or U6312 (N_6312,N_4803,N_5732);
and U6313 (N_6313,N_4076,N_5302);
and U6314 (N_6314,N_4706,N_4482);
and U6315 (N_6315,N_5926,N_4987);
or U6316 (N_6316,N_5713,N_5143);
or U6317 (N_6317,N_5120,N_5450);
nand U6318 (N_6318,N_5308,N_5818);
nand U6319 (N_6319,N_5544,N_4449);
nand U6320 (N_6320,N_5694,N_5960);
nand U6321 (N_6321,N_5063,N_5915);
and U6322 (N_6322,N_5211,N_5185);
nor U6323 (N_6323,N_4514,N_4496);
and U6324 (N_6324,N_4519,N_4051);
or U6325 (N_6325,N_5697,N_5044);
or U6326 (N_6326,N_5842,N_5301);
nand U6327 (N_6327,N_4017,N_4249);
and U6328 (N_6328,N_4083,N_5941);
nor U6329 (N_6329,N_5766,N_4036);
or U6330 (N_6330,N_5428,N_4937);
nor U6331 (N_6331,N_4397,N_5122);
nor U6332 (N_6332,N_4582,N_4045);
nor U6333 (N_6333,N_5731,N_4199);
and U6334 (N_6334,N_4148,N_4094);
nand U6335 (N_6335,N_4890,N_5834);
and U6336 (N_6336,N_5804,N_5619);
or U6337 (N_6337,N_4355,N_4968);
or U6338 (N_6338,N_4539,N_4782);
xnor U6339 (N_6339,N_4068,N_4306);
nand U6340 (N_6340,N_5734,N_4465);
nor U6341 (N_6341,N_4085,N_5087);
nand U6342 (N_6342,N_4191,N_4212);
and U6343 (N_6343,N_5735,N_4813);
and U6344 (N_6344,N_4432,N_5985);
nand U6345 (N_6345,N_5422,N_5753);
nand U6346 (N_6346,N_5489,N_4902);
or U6347 (N_6347,N_4248,N_4305);
xnor U6348 (N_6348,N_4728,N_5890);
or U6349 (N_6349,N_4687,N_4290);
or U6350 (N_6350,N_5562,N_4256);
or U6351 (N_6351,N_4826,N_4182);
nand U6352 (N_6352,N_4058,N_5680);
nor U6353 (N_6353,N_4329,N_4629);
xnor U6354 (N_6354,N_5587,N_4835);
nor U6355 (N_6355,N_4379,N_5510);
nor U6356 (N_6356,N_4447,N_4579);
nor U6357 (N_6357,N_5130,N_4810);
nor U6358 (N_6358,N_5527,N_5566);
nor U6359 (N_6359,N_5950,N_5188);
nand U6360 (N_6360,N_5730,N_4601);
nor U6361 (N_6361,N_5016,N_5822);
nor U6362 (N_6362,N_5774,N_4716);
nor U6363 (N_6363,N_4922,N_5026);
or U6364 (N_6364,N_5663,N_5480);
nor U6365 (N_6365,N_4301,N_5009);
nand U6366 (N_6366,N_5752,N_5712);
or U6367 (N_6367,N_4278,N_5775);
or U6368 (N_6368,N_5645,N_4775);
nand U6369 (N_6369,N_4504,N_5388);
or U6370 (N_6370,N_5223,N_4769);
and U6371 (N_6371,N_4059,N_5452);
and U6372 (N_6372,N_5075,N_5670);
nand U6373 (N_6373,N_4580,N_4204);
nand U6374 (N_6374,N_5632,N_4650);
nor U6375 (N_6375,N_4612,N_4061);
and U6376 (N_6376,N_4285,N_4822);
and U6377 (N_6377,N_4236,N_5689);
nand U6378 (N_6378,N_5541,N_5424);
and U6379 (N_6379,N_4973,N_5342);
nor U6380 (N_6380,N_4494,N_4560);
or U6381 (N_6381,N_4912,N_4972);
nor U6382 (N_6382,N_4645,N_5710);
and U6383 (N_6383,N_5235,N_5290);
nand U6384 (N_6384,N_5103,N_4908);
nor U6385 (N_6385,N_4512,N_4961);
nor U6386 (N_6386,N_4228,N_4773);
and U6387 (N_6387,N_4842,N_5291);
nand U6388 (N_6388,N_4201,N_4005);
nand U6389 (N_6389,N_4824,N_5626);
nor U6390 (N_6390,N_5855,N_5791);
and U6391 (N_6391,N_5258,N_4192);
nor U6392 (N_6392,N_4302,N_5473);
and U6393 (N_6393,N_5976,N_5236);
nand U6394 (N_6394,N_4127,N_5703);
nand U6395 (N_6395,N_5929,N_4269);
and U6396 (N_6396,N_4510,N_4602);
nand U6397 (N_6397,N_4405,N_4097);
and U6398 (N_6398,N_5820,N_4607);
or U6399 (N_6399,N_4347,N_4980);
or U6400 (N_6400,N_4467,N_5512);
and U6401 (N_6401,N_5604,N_4471);
and U6402 (N_6402,N_4719,N_4703);
and U6403 (N_6403,N_5012,N_5673);
nand U6404 (N_6404,N_5624,N_5553);
or U6405 (N_6405,N_5651,N_4371);
and U6406 (N_6406,N_5859,N_5250);
and U6407 (N_6407,N_5704,N_4251);
and U6408 (N_6408,N_5523,N_5685);
nor U6409 (N_6409,N_5771,N_4877);
or U6410 (N_6410,N_5715,N_4959);
nor U6411 (N_6411,N_5788,N_5314);
nor U6412 (N_6412,N_4833,N_4396);
and U6413 (N_6413,N_4966,N_5564);
nand U6414 (N_6414,N_5182,N_4014);
and U6415 (N_6415,N_5591,N_4375);
or U6416 (N_6416,N_5081,N_4797);
or U6417 (N_6417,N_5227,N_4751);
nand U6418 (N_6418,N_5029,N_5583);
nor U6419 (N_6419,N_5336,N_4619);
nand U6420 (N_6420,N_5225,N_4361);
nand U6421 (N_6421,N_4413,N_4096);
nand U6422 (N_6422,N_4105,N_4675);
or U6423 (N_6423,N_4103,N_5412);
and U6424 (N_6424,N_4056,N_5239);
nor U6425 (N_6425,N_4044,N_5064);
or U6426 (N_6426,N_5674,N_5170);
xnor U6427 (N_6427,N_5474,N_5642);
nor U6428 (N_6428,N_4656,N_5940);
nand U6429 (N_6429,N_4223,N_4339);
and U6430 (N_6430,N_5551,N_5065);
nand U6431 (N_6431,N_5410,N_4523);
nand U6432 (N_6432,N_5397,N_5810);
and U6433 (N_6433,N_5776,N_5497);
nand U6434 (N_6434,N_4718,N_5537);
nor U6435 (N_6435,N_5603,N_4587);
and U6436 (N_6436,N_4015,N_4267);
or U6437 (N_6437,N_5681,N_4350);
nor U6438 (N_6438,N_4317,N_4624);
or U6439 (N_6439,N_5797,N_5353);
and U6440 (N_6440,N_5581,N_4893);
nor U6441 (N_6441,N_4092,N_5778);
nor U6442 (N_6442,N_4615,N_5808);
and U6443 (N_6443,N_4709,N_5573);
and U6444 (N_6444,N_5905,N_4925);
and U6445 (N_6445,N_5316,N_5980);
or U6446 (N_6446,N_4904,N_4781);
nand U6447 (N_6447,N_5286,N_5265);
and U6448 (N_6448,N_4897,N_4296);
nor U6449 (N_6449,N_4508,N_4850);
and U6450 (N_6450,N_5443,N_5435);
nor U6451 (N_6451,N_4899,N_5816);
nor U6452 (N_6452,N_5669,N_4187);
nor U6453 (N_6453,N_5166,N_4572);
and U6454 (N_6454,N_5198,N_4870);
nand U6455 (N_6455,N_5515,N_5542);
and U6456 (N_6456,N_4944,N_4366);
or U6457 (N_6457,N_5767,N_4153);
nand U6458 (N_6458,N_5073,N_5259);
and U6459 (N_6459,N_4674,N_5457);
nor U6460 (N_6460,N_5139,N_4489);
xnor U6461 (N_6461,N_4472,N_5634);
nand U6462 (N_6462,N_5944,N_4456);
nand U6463 (N_6463,N_5484,N_5836);
xnor U6464 (N_6464,N_5355,N_4861);
or U6465 (N_6465,N_5599,N_4522);
nor U6466 (N_6466,N_4310,N_5882);
and U6467 (N_6467,N_5839,N_4827);
nand U6468 (N_6468,N_5106,N_5162);
nand U6469 (N_6469,N_4091,N_5636);
nand U6470 (N_6470,N_5917,N_5784);
nand U6471 (N_6471,N_4932,N_5490);
nand U6472 (N_6472,N_5829,N_4427);
nor U6473 (N_6473,N_5840,N_4479);
nor U6474 (N_6474,N_5801,N_4452);
or U6475 (N_6475,N_5639,N_4506);
and U6476 (N_6476,N_5303,N_5067);
and U6477 (N_6477,N_4664,N_5008);
or U6478 (N_6478,N_4883,N_5267);
and U6479 (N_6479,N_4620,N_5338);
and U6480 (N_6480,N_5194,N_4478);
nand U6481 (N_6481,N_4254,N_4215);
and U6482 (N_6482,N_4801,N_5554);
nor U6483 (N_6483,N_4383,N_4300);
and U6484 (N_6484,N_5401,N_5212);
nor U6485 (N_6485,N_5351,N_4177);
nor U6486 (N_6486,N_4216,N_5270);
nand U6487 (N_6487,N_4685,N_5133);
nor U6488 (N_6488,N_4287,N_5368);
or U6489 (N_6489,N_5692,N_4631);
or U6490 (N_6490,N_5494,N_4786);
nand U6491 (N_6491,N_5327,N_5830);
nor U6492 (N_6492,N_4839,N_5958);
nand U6493 (N_6493,N_5597,N_4743);
nor U6494 (N_6494,N_5360,N_4969);
nand U6495 (N_6495,N_4353,N_5613);
nor U6496 (N_6496,N_5319,N_5615);
nor U6497 (N_6497,N_5471,N_5481);
nand U6498 (N_6498,N_5973,N_5396);
nor U6499 (N_6499,N_5365,N_4677);
nor U6500 (N_6500,N_4481,N_4626);
nand U6501 (N_6501,N_4930,N_5295);
nand U6502 (N_6502,N_4881,N_5096);
nor U6503 (N_6503,N_4795,N_4322);
nor U6504 (N_6504,N_5658,N_5939);
or U6505 (N_6505,N_4299,N_5977);
and U6506 (N_6506,N_4259,N_4950);
nor U6507 (N_6507,N_5884,N_5086);
nand U6508 (N_6508,N_4807,N_4042);
or U6509 (N_6509,N_4748,N_4428);
or U6510 (N_6510,N_4279,N_4891);
xor U6511 (N_6511,N_5899,N_5344);
nor U6512 (N_6512,N_4307,N_5202);
nand U6513 (N_6513,N_5157,N_4033);
nand U6514 (N_6514,N_4988,N_4140);
and U6515 (N_6515,N_4812,N_5653);
or U6516 (N_6516,N_4753,N_4368);
or U6517 (N_6517,N_5264,N_5165);
nor U6518 (N_6518,N_4643,N_4412);
or U6519 (N_6519,N_5503,N_4497);
and U6520 (N_6520,N_4732,N_5274);
nor U6521 (N_6521,N_4965,N_4049);
nand U6522 (N_6522,N_5986,N_4726);
or U6523 (N_6523,N_4210,N_4816);
nor U6524 (N_6524,N_4911,N_5686);
nor U6525 (N_6525,N_4158,N_4275);
nor U6526 (N_6526,N_5959,N_4727);
and U6527 (N_6527,N_4838,N_4731);
nor U6528 (N_6528,N_4935,N_5946);
nor U6529 (N_6529,N_5215,N_4400);
nand U6530 (N_6530,N_4188,N_4004);
nand U6531 (N_6531,N_4955,N_4134);
nor U6532 (N_6532,N_5241,N_4006);
xor U6533 (N_6533,N_5546,N_5159);
nand U6534 (N_6534,N_5246,N_5533);
and U6535 (N_6535,N_4543,N_5931);
nor U6536 (N_6536,N_5665,N_4012);
nor U6537 (N_6537,N_5802,N_4167);
and U6538 (N_6538,N_5875,N_4613);
or U6539 (N_6539,N_5969,N_5711);
and U6540 (N_6540,N_4316,N_4997);
or U6541 (N_6541,N_5306,N_4295);
and U6542 (N_6542,N_4262,N_5762);
nand U6543 (N_6543,N_5617,N_5378);
or U6544 (N_6544,N_5254,N_4233);
nand U6545 (N_6545,N_5981,N_5876);
nor U6546 (N_6546,N_5770,N_5245);
nor U6547 (N_6547,N_4696,N_4655);
nand U6548 (N_6548,N_4749,N_5742);
and U6549 (N_6549,N_4205,N_5337);
or U6550 (N_6550,N_4100,N_5769);
or U6551 (N_6551,N_5793,N_4129);
nand U6552 (N_6552,N_4740,N_4896);
and U6553 (N_6553,N_4265,N_5990);
xor U6554 (N_6554,N_4639,N_4788);
and U6555 (N_6555,N_5359,N_4054);
or U6556 (N_6556,N_4557,N_4474);
nor U6557 (N_6557,N_5852,N_5621);
nand U6558 (N_6558,N_4981,N_5114);
nor U6559 (N_6559,N_4360,N_5751);
and U6560 (N_6560,N_5937,N_5805);
and U6561 (N_6561,N_5041,N_4388);
or U6562 (N_6562,N_4399,N_4122);
or U6563 (N_6563,N_4946,N_4401);
and U6564 (N_6564,N_5848,N_4047);
and U6565 (N_6565,N_5407,N_5018);
or U6566 (N_6566,N_4229,N_4931);
and U6567 (N_6567,N_4559,N_4116);
or U6568 (N_6568,N_5420,N_4476);
nor U6569 (N_6569,N_5719,N_4491);
and U6570 (N_6570,N_4203,N_4160);
and U6571 (N_6571,N_4840,N_5849);
or U6572 (N_6572,N_4614,N_4591);
and U6573 (N_6573,N_4707,N_4345);
nand U6574 (N_6574,N_5369,N_5332);
nor U6575 (N_6575,N_5529,N_5933);
nand U6576 (N_6576,N_5150,N_4928);
or U6577 (N_6577,N_5180,N_5571);
or U6578 (N_6578,N_4600,N_5687);
xor U6579 (N_6579,N_4563,N_5682);
nand U6580 (N_6580,N_5047,N_4984);
or U6581 (N_6581,N_4793,N_5717);
xor U6582 (N_6582,N_5423,N_4284);
nand U6583 (N_6583,N_5456,N_5924);
nor U6584 (N_6584,N_4466,N_4646);
and U6585 (N_6585,N_5698,N_4534);
nand U6586 (N_6586,N_4635,N_5500);
nor U6587 (N_6587,N_4072,N_5238);
nand U6588 (N_6588,N_5119,N_5953);
nand U6589 (N_6589,N_4695,N_4668);
or U6590 (N_6590,N_5690,N_5565);
xor U6591 (N_6591,N_5322,N_5426);
or U6592 (N_6592,N_5832,N_4683);
nand U6593 (N_6593,N_5589,N_5637);
nand U6594 (N_6594,N_5350,N_5555);
or U6595 (N_6595,N_4622,N_4247);
and U6596 (N_6596,N_4638,N_5688);
nor U6597 (N_6597,N_4346,N_5595);
nand U6598 (N_6598,N_5000,N_5644);
nand U6599 (N_6599,N_4712,N_5708);
nand U6600 (N_6600,N_4475,N_5181);
nand U6601 (N_6601,N_4670,N_4916);
or U6602 (N_6602,N_5486,N_5625);
nand U6603 (N_6603,N_5057,N_4025);
and U6604 (N_6604,N_5315,N_4312);
nand U6605 (N_6605,N_5136,N_4422);
nand U6606 (N_6606,N_5115,N_5580);
and U6607 (N_6607,N_5612,N_5376);
nor U6608 (N_6608,N_4549,N_4365);
or U6609 (N_6609,N_4882,N_4887);
or U6610 (N_6610,N_5857,N_5283);
xor U6611 (N_6611,N_5511,N_4429);
and U6612 (N_6612,N_4661,N_4874);
or U6613 (N_6613,N_5891,N_5116);
and U6614 (N_6614,N_5059,N_5045);
and U6615 (N_6615,N_5373,N_5954);
nor U6616 (N_6616,N_5147,N_5656);
nand U6617 (N_6617,N_4099,N_4445);
and U6618 (N_6618,N_4243,N_5556);
nor U6619 (N_6619,N_5957,N_5341);
xnor U6620 (N_6620,N_4971,N_4451);
xnor U6621 (N_6621,N_4063,N_4138);
or U6622 (N_6622,N_4170,N_4774);
nand U6623 (N_6623,N_4463,N_5995);
nor U6624 (N_6624,N_5970,N_5109);
and U6625 (N_6625,N_5607,N_5927);
nand U6626 (N_6626,N_5321,N_4785);
nor U6627 (N_6627,N_5046,N_4820);
nand U6628 (N_6628,N_5996,N_4871);
nor U6629 (N_6629,N_4035,N_4885);
nand U6630 (N_6630,N_5695,N_4864);
or U6631 (N_6631,N_5179,N_4625);
nand U6632 (N_6632,N_5499,N_5174);
or U6633 (N_6633,N_5881,N_4196);
or U6634 (N_6634,N_4958,N_4118);
nand U6635 (N_6635,N_5539,N_4509);
and U6636 (N_6636,N_5382,N_4146);
or U6637 (N_6637,N_5563,N_5190);
nor U6638 (N_6638,N_4356,N_5889);
or U6639 (N_6639,N_4876,N_4594);
and U6640 (N_6640,N_4800,N_4665);
nand U6641 (N_6641,N_5620,N_5825);
nand U6642 (N_6642,N_5904,N_4888);
and U6643 (N_6643,N_5463,N_4642);
nor U6644 (N_6644,N_5906,N_4328);
or U6645 (N_6645,N_4186,N_4441);
and U6646 (N_6646,N_5175,N_5726);
nand U6647 (N_6647,N_4777,N_5921);
nand U6648 (N_6648,N_4821,N_5348);
and U6649 (N_6649,N_5664,N_5908);
or U6650 (N_6650,N_4738,N_5220);
or U6651 (N_6651,N_4266,N_5472);
nor U6652 (N_6652,N_4900,N_5475);
nor U6653 (N_6653,N_5104,N_5600);
or U6654 (N_6654,N_4982,N_5380);
and U6655 (N_6655,N_5608,N_4291);
and U6656 (N_6656,N_4473,N_4128);
nand U6657 (N_6657,N_4162,N_4603);
and U6658 (N_6658,N_5284,N_5965);
or U6659 (N_6659,N_4604,N_4114);
and U6660 (N_6660,N_4206,N_5273);
or U6661 (N_6661,N_5549,N_5858);
and U6662 (N_6662,N_4338,N_5479);
or U6663 (N_6663,N_5509,N_5596);
or U6664 (N_6664,N_5487,N_4970);
and U6665 (N_6665,N_5495,N_5635);
or U6666 (N_6666,N_4762,N_4964);
nor U6667 (N_6667,N_4859,N_5684);
and U6668 (N_6668,N_4963,N_4334);
nor U6669 (N_6669,N_5403,N_5406);
xor U6670 (N_6670,N_5402,N_5252);
nor U6671 (N_6671,N_5800,N_5101);
nor U6672 (N_6672,N_4952,N_5545);
nand U6673 (N_6673,N_4486,N_5281);
or U6674 (N_6674,N_5992,N_4819);
and U6675 (N_6675,N_5983,N_4586);
nor U6676 (N_6676,N_5668,N_5799);
nor U6677 (N_6677,N_5768,N_5601);
and U6678 (N_6678,N_4596,N_4879);
and U6679 (N_6679,N_5219,N_5069);
nand U6680 (N_6680,N_5058,N_5602);
or U6681 (N_6681,N_4416,N_4780);
and U6682 (N_6682,N_5887,N_4219);
nand U6683 (N_6683,N_5033,N_4992);
nand U6684 (N_6684,N_5088,N_4080);
or U6685 (N_6685,N_4671,N_5869);
and U6686 (N_6686,N_5395,N_5693);
or U6687 (N_6687,N_4791,N_5744);
nor U6688 (N_6688,N_4028,N_4011);
nand U6689 (N_6689,N_5504,N_4652);
or U6690 (N_6690,N_4469,N_4120);
and U6691 (N_6691,N_4697,N_4689);
and U6692 (N_6692,N_5894,N_4462);
nand U6693 (N_6693,N_4431,N_5948);
and U6694 (N_6694,N_4943,N_5700);
and U6695 (N_6695,N_5309,N_4437);
and U6696 (N_6696,N_4381,N_5467);
or U6697 (N_6697,N_5074,N_5298);
nand U6698 (N_6698,N_5366,N_4617);
nor U6699 (N_6699,N_5039,N_5030);
nand U6700 (N_6700,N_5002,N_4101);
nor U6701 (N_6701,N_4694,N_4484);
and U6702 (N_6702,N_5330,N_4077);
nor U6703 (N_6703,N_4373,N_5630);
nor U6704 (N_6704,N_4717,N_5947);
nand U6705 (N_6705,N_5186,N_4855);
nor U6706 (N_6706,N_5445,N_5176);
nand U6707 (N_6707,N_5392,N_4927);
nor U6708 (N_6708,N_4457,N_5117);
nand U6709 (N_6709,N_5464,N_5021);
nor U6710 (N_6710,N_4126,N_5513);
nand U6711 (N_6711,N_4632,N_5491);
nand U6712 (N_6712,N_4152,N_4618);
and U6713 (N_6713,N_5844,N_5885);
nand U6714 (N_6714,N_5783,N_4398);
nand U6715 (N_6715,N_4768,N_4319);
nand U6716 (N_6716,N_5598,N_5451);
nand U6717 (N_6717,N_4034,N_4884);
or U6718 (N_6718,N_5896,N_5938);
nor U6719 (N_6719,N_4344,N_4189);
nand U6720 (N_6720,N_4978,N_4845);
nor U6721 (N_6721,N_5967,N_5251);
and U6722 (N_6722,N_4725,N_4124);
nor U6723 (N_6723,N_4163,N_4009);
nor U6724 (N_6724,N_5079,N_4435);
nand U6725 (N_6725,N_4690,N_5108);
and U6726 (N_6726,N_4848,N_4436);
or U6727 (N_6727,N_5304,N_4679);
nor U6728 (N_6728,N_4407,N_5118);
nor U6729 (N_6729,N_4417,N_5968);
and U6730 (N_6730,N_4404,N_5433);
or U6731 (N_6731,N_5483,N_4798);
and U6732 (N_6732,N_5640,N_4443);
and U6733 (N_6733,N_5806,N_5419);
xor U6734 (N_6734,N_4446,N_5276);
nand U6735 (N_6735,N_5203,N_5446);
and U6736 (N_6736,N_4765,N_4521);
or U6737 (N_6737,N_4343,N_4856);
or U6738 (N_6738,N_4031,N_4986);
nand U6739 (N_6739,N_5582,N_5213);
and U6740 (N_6740,N_5462,N_4142);
and U6741 (N_6741,N_5052,N_5210);
nand U6742 (N_6742,N_4172,N_4323);
or U6743 (N_6743,N_5886,N_4593);
nand U6744 (N_6744,N_5650,N_4533);
or U6745 (N_6745,N_4863,N_4849);
or U6746 (N_6746,N_4704,N_4562);
nor U6747 (N_6747,N_4393,N_4585);
nand U6748 (N_6748,N_4271,N_5085);
or U6749 (N_6749,N_4238,N_4806);
or U6750 (N_6750,N_4341,N_5907);
nor U6751 (N_6751,N_5724,N_4198);
nand U6752 (N_6752,N_5616,N_5701);
nor U6753 (N_6753,N_4584,N_5128);
or U6754 (N_6754,N_5013,N_4566);
nor U6755 (N_6755,N_4050,N_4374);
nor U6756 (N_6756,N_4409,N_4156);
or U6757 (N_6757,N_4460,N_4002);
nand U6758 (N_6758,N_5216,N_4744);
xor U6759 (N_6759,N_4298,N_4283);
nor U6760 (N_6760,N_4831,N_4389);
or U6761 (N_6761,N_5042,N_4983);
nor U6762 (N_6762,N_5610,N_5329);
nand U6763 (N_6763,N_4733,N_4415);
and U6764 (N_6764,N_5716,N_4866);
and U6765 (N_6765,N_4255,N_5145);
and U6766 (N_6766,N_4721,N_4420);
or U6767 (N_6767,N_5240,N_4109);
and U6768 (N_6768,N_4161,N_5415);
nand U6769 (N_6769,N_4745,N_5873);
or U6770 (N_6770,N_5667,N_4637);
nor U6771 (N_6771,N_4007,N_5349);
or U6772 (N_6772,N_5247,N_5878);
and U6773 (N_6773,N_5437,N_5431);
nor U6774 (N_6774,N_5520,N_4583);
xor U6775 (N_6775,N_4502,N_5517);
and U6776 (N_6776,N_4272,N_4962);
xor U6777 (N_6777,N_4175,N_5324);
nor U6778 (N_6778,N_5169,N_4403);
nand U6779 (N_6779,N_5678,N_4178);
and U6780 (N_6780,N_5631,N_5004);
nand U6781 (N_6781,N_4778,N_5340);
nand U6782 (N_6782,N_5381,N_4173);
nor U6783 (N_6783,N_5577,N_5759);
and U6784 (N_6784,N_5584,N_5221);
or U6785 (N_6785,N_4905,N_5524);
nand U6786 (N_6786,N_5196,N_5163);
nor U6787 (N_6787,N_4841,N_4921);
nor U6788 (N_6788,N_5153,N_4611);
nand U6789 (N_6789,N_5230,N_4628);
and U6790 (N_6790,N_4149,N_5411);
nor U6791 (N_6791,N_4957,N_5737);
and U6792 (N_6792,N_4102,N_4135);
nand U6793 (N_6793,N_4975,N_4303);
nand U6794 (N_6794,N_5874,N_5657);
nor U6795 (N_6795,N_4581,N_4386);
or U6796 (N_6796,N_4490,N_4799);
nand U6797 (N_6797,N_5234,N_4440);
nand U6798 (N_6798,N_5158,N_4784);
nand U6799 (N_6799,N_5903,N_5083);
nand U6800 (N_6800,N_5333,N_5345);
nor U6801 (N_6801,N_5076,N_4699);
or U6802 (N_6802,N_4544,N_5532);
and U6803 (N_6803,N_4239,N_5425);
nor U6804 (N_6804,N_4764,N_5761);
xor U6805 (N_6805,N_5430,N_5920);
nand U6806 (N_6806,N_4358,N_5780);
nand U6807 (N_6807,N_4010,N_5146);
and U6808 (N_6808,N_5558,N_4649);
nor U6809 (N_6809,N_5015,N_5367);
nor U6810 (N_6810,N_5961,N_4832);
and U6811 (N_6811,N_5962,N_5377);
or U6812 (N_6812,N_5307,N_5149);
and U6813 (N_6813,N_4790,N_5278);
nor U6814 (N_6814,N_4837,N_5758);
or U6815 (N_6815,N_4309,N_4729);
nor U6816 (N_6816,N_4402,N_4410);
nand U6817 (N_6817,N_4867,N_5028);
xor U6818 (N_6818,N_5932,N_5288);
or U6819 (N_6819,N_4089,N_5789);
nand U6820 (N_6820,N_4811,N_4892);
and U6821 (N_6821,N_4111,N_5614);
or U6822 (N_6822,N_4934,N_4168);
or U6823 (N_6823,N_5055,N_4037);
and U6824 (N_6824,N_5253,N_5827);
and U6825 (N_6825,N_4693,N_5646);
or U6826 (N_6826,N_5648,N_4755);
or U6827 (N_6827,N_4651,N_5974);
xor U6828 (N_6828,N_5310,N_4545);
or U6829 (N_6829,N_4633,N_5576);
nand U6830 (N_6830,N_4327,N_4608);
nand U6831 (N_6831,N_4737,N_5305);
xnor U6832 (N_6832,N_4232,N_4547);
or U6833 (N_6833,N_4567,N_5575);
nand U6834 (N_6834,N_5468,N_4333);
nand U6835 (N_6835,N_5794,N_4174);
or U6836 (N_6836,N_4552,N_5777);
nand U6837 (N_6837,N_4418,N_4573);
nor U6838 (N_6838,N_5900,N_5187);
nand U6839 (N_6839,N_5449,N_4179);
and U6840 (N_6840,N_4599,N_5346);
nor U6841 (N_6841,N_4226,N_5847);
nand U6842 (N_6842,N_5570,N_4108);
nand U6843 (N_6843,N_4055,N_4320);
nand U6844 (N_6844,N_5024,N_5923);
nor U6845 (N_6845,N_5736,N_5134);
or U6846 (N_6846,N_4119,N_5935);
and U6847 (N_6847,N_5870,N_4125);
and U6848 (N_6848,N_5972,N_4064);
nor U6849 (N_6849,N_4779,N_5297);
nor U6850 (N_6850,N_5093,N_5331);
nand U6851 (N_6851,N_5427,N_5611);
and U6852 (N_6852,N_4681,N_5218);
nand U6853 (N_6853,N_5070,N_4377);
and U6854 (N_6854,N_5978,N_5557);
or U6855 (N_6855,N_4147,N_5660);
nand U6856 (N_6856,N_5066,N_4941);
or U6857 (N_6857,N_4246,N_4211);
and U6858 (N_6858,N_4714,N_4244);
or U6859 (N_6859,N_5469,N_5429);
nor U6860 (N_6860,N_5826,N_4332);
and U6861 (N_6861,N_5124,N_4949);
nand U6862 (N_6862,N_4542,N_4710);
nand U6863 (N_6863,N_4093,N_4933);
or U6864 (N_6864,N_4392,N_4367);
and U6865 (N_6865,N_5672,N_4571);
nor U6866 (N_6866,N_5325,N_4369);
or U6867 (N_6867,N_5550,N_4450);
and U6868 (N_6868,N_5287,N_5131);
nand U6869 (N_6869,N_5866,N_4263);
nor U6870 (N_6870,N_5352,N_4442);
nand U6871 (N_6871,N_4073,N_5061);
or U6872 (N_6872,N_4106,N_5498);
nor U6873 (N_6873,N_5593,N_4053);
or U6874 (N_6874,N_5982,N_5222);
nand U6875 (N_6875,N_4688,N_5936);
xor U6876 (N_6876,N_4121,N_5798);
and U6877 (N_6877,N_5649,N_5823);
nand U6878 (N_6878,N_4766,N_5743);
or U6879 (N_6879,N_5082,N_4818);
or U6880 (N_6880,N_5699,N_5328);
and U6881 (N_6881,N_5078,N_4139);
or U6882 (N_6882,N_4536,N_4550);
nand U6883 (N_6883,N_4136,N_4654);
and U6884 (N_6884,N_4923,N_4759);
and U6885 (N_6885,N_4906,N_4181);
nor U6886 (N_6886,N_4577,N_4133);
and U6887 (N_6887,N_4313,N_5721);
nand U6888 (N_6888,N_5641,N_5011);
nand U6889 (N_6889,N_4794,N_4040);
or U6890 (N_6890,N_5828,N_4408);
or U6891 (N_6891,N_4304,N_4956);
nand U6892 (N_6892,N_5056,N_4137);
and U6893 (N_6893,N_5209,N_5819);
or U6894 (N_6894,N_4112,N_4110);
nand U6895 (N_6895,N_4634,N_5781);
or U6896 (N_6896,N_4088,N_5530);
or U6897 (N_6897,N_5988,N_5893);
nor U6898 (N_6898,N_5444,N_4939);
and U6899 (N_6899,N_5374,N_4708);
or U6900 (N_6900,N_4758,N_4115);
or U6901 (N_6901,N_4565,N_5534);
nand U6902 (N_6902,N_5125,N_4117);
nand U6903 (N_6903,N_5261,N_4362);
nand U6904 (N_6904,N_4815,N_5493);
nor U6905 (N_6905,N_5813,N_5100);
nor U6906 (N_6906,N_5300,N_5633);
and U6907 (N_6907,N_4590,N_4240);
or U6908 (N_6908,N_5627,N_5003);
or U6909 (N_6909,N_5994,N_5740);
nor U6910 (N_6910,N_5160,N_4411);
nor U6911 (N_6911,N_5846,N_4075);
and U6912 (N_6912,N_5606,N_4783);
nand U6913 (N_6913,N_4564,N_5705);
or U6914 (N_6914,N_4227,N_4159);
nor U6915 (N_6915,N_4551,N_5398);
or U6916 (N_6916,N_4270,N_5482);
nand U6917 (N_6917,N_4297,N_4493);
or U6918 (N_6918,N_4680,N_5709);
nand U6919 (N_6919,N_4292,N_4052);
or U6920 (N_6920,N_4868,N_5335);
or U6921 (N_6921,N_5652,N_5835);
or U6922 (N_6922,N_5526,N_4495);
or U6923 (N_6923,N_4492,N_5628);
and U6924 (N_6924,N_5871,N_4425);
and U6925 (N_6925,N_4998,N_4194);
xor U6926 (N_6926,N_4260,N_5053);
nor U6927 (N_6927,N_4787,N_4936);
and U6928 (N_6928,N_4019,N_4041);
nand U6929 (N_6929,N_5107,N_4039);
nor U6930 (N_6930,N_4430,N_4202);
nor U6931 (N_6931,N_4084,N_5993);
nand U6932 (N_6932,N_5453,N_5268);
nor U6933 (N_6933,N_5912,N_4529);
nor U6934 (N_6934,N_5095,N_5005);
or U6935 (N_6935,N_5792,N_4903);
or U6936 (N_6936,N_4926,N_4390);
nor U6937 (N_6937,N_4623,N_4576);
nor U6938 (N_6938,N_4154,N_5738);
or U6939 (N_6939,N_5054,N_4561);
nor U6940 (N_6940,N_4104,N_4141);
or U6941 (N_6941,N_5989,N_5560);
and U6942 (N_6942,N_4948,N_5914);
or U6943 (N_6943,N_5272,N_5727);
nand U6944 (N_6944,N_4880,N_4364);
and U6945 (N_6945,N_4444,N_4176);
and U6946 (N_6946,N_4724,N_4541);
or U6947 (N_6947,N_4095,N_4530);
nor U6948 (N_6948,N_4735,N_5966);
or U6949 (N_6949,N_5049,N_4578);
and U6950 (N_6950,N_5442,N_4875);
nand U6951 (N_6951,N_4234,N_4507);
or U6952 (N_6952,N_5714,N_4641);
nand U6953 (N_6953,N_5383,N_4991);
nand U6954 (N_6954,N_4511,N_4231);
or U6955 (N_6955,N_5072,N_5586);
or U6956 (N_6956,N_4157,N_4979);
or U6957 (N_6957,N_4470,N_4387);
or U6958 (N_6958,N_4438,N_5785);
and U6959 (N_6959,N_5080,N_4151);
xnor U6960 (N_6960,N_5476,N_4672);
nand U6961 (N_6961,N_4098,N_4209);
nor U6962 (N_6962,N_5313,N_5505);
nand U6963 (N_6963,N_4889,N_5320);
or U6964 (N_6964,N_4000,N_5868);
xnor U6965 (N_6965,N_5707,N_5022);
nor U6966 (N_6966,N_5902,N_5409);
nor U6967 (N_6967,N_5040,N_5795);
or U6968 (N_6968,N_5748,N_5441);
nor U6969 (N_6969,N_5552,N_4123);
nand U6970 (N_6970,N_4673,N_5126);
or U6971 (N_6971,N_5248,N_5654);
nor U6972 (N_6972,N_4825,N_5723);
and U6973 (N_6973,N_4230,N_5173);
or U6974 (N_6974,N_4678,N_4994);
and U6975 (N_6975,N_5765,N_5379);
or U6976 (N_6976,N_5448,N_5872);
nor U6977 (N_6977,N_4517,N_5851);
or U6978 (N_6978,N_5492,N_4268);
nand U6979 (N_6979,N_5888,N_5647);
and U6980 (N_6980,N_4250,N_4314);
and U6981 (N_6981,N_5204,N_4286);
nor U6982 (N_6982,N_5112,N_5266);
or U6983 (N_6983,N_4942,N_4574);
nor U6984 (N_6984,N_4038,N_4918);
nand U6985 (N_6985,N_4554,N_5984);
or U6986 (N_6986,N_4723,N_5579);
or U6987 (N_6987,N_5263,N_5536);
nand U6988 (N_6988,N_5856,N_4805);
and U6989 (N_6989,N_5949,N_5206);
nand U6990 (N_6990,N_4348,N_4518);
nor U6991 (N_6991,N_4985,N_5760);
and U6992 (N_6992,N_4166,N_5034);
xnor U6993 (N_6993,N_5845,N_4999);
or U6994 (N_6994,N_4996,N_5193);
and U6995 (N_6995,N_5317,N_5508);
nor U6996 (N_6996,N_5465,N_5318);
nor U6997 (N_6997,N_4195,N_5432);
nand U6998 (N_6998,N_5540,N_4214);
or U6999 (N_6999,N_4990,N_4993);
nand U7000 (N_7000,N_4690,N_5667);
nand U7001 (N_7001,N_4497,N_5395);
and U7002 (N_7002,N_4298,N_4320);
or U7003 (N_7003,N_5138,N_4318);
xnor U7004 (N_7004,N_5833,N_4749);
and U7005 (N_7005,N_5328,N_5643);
and U7006 (N_7006,N_5094,N_5882);
nand U7007 (N_7007,N_4059,N_5142);
and U7008 (N_7008,N_5495,N_4161);
and U7009 (N_7009,N_5292,N_5307);
or U7010 (N_7010,N_4842,N_4601);
and U7011 (N_7011,N_5606,N_5969);
nor U7012 (N_7012,N_5323,N_4045);
or U7013 (N_7013,N_5230,N_5847);
nand U7014 (N_7014,N_4804,N_4809);
or U7015 (N_7015,N_4629,N_5965);
nand U7016 (N_7016,N_5148,N_5064);
nor U7017 (N_7017,N_4997,N_5083);
or U7018 (N_7018,N_4843,N_5108);
nor U7019 (N_7019,N_4754,N_4433);
nand U7020 (N_7020,N_5306,N_4363);
or U7021 (N_7021,N_4625,N_5928);
nor U7022 (N_7022,N_4975,N_5888);
and U7023 (N_7023,N_5185,N_4151);
nor U7024 (N_7024,N_5757,N_4625);
nor U7025 (N_7025,N_4809,N_4697);
and U7026 (N_7026,N_5854,N_5054);
nand U7027 (N_7027,N_4974,N_4272);
and U7028 (N_7028,N_4753,N_5620);
nand U7029 (N_7029,N_4248,N_5742);
nand U7030 (N_7030,N_5529,N_4813);
or U7031 (N_7031,N_5163,N_4524);
nor U7032 (N_7032,N_4294,N_4685);
nor U7033 (N_7033,N_4299,N_4869);
nand U7034 (N_7034,N_4189,N_5554);
and U7035 (N_7035,N_4029,N_4972);
nand U7036 (N_7036,N_5651,N_4388);
or U7037 (N_7037,N_4237,N_5636);
nand U7038 (N_7038,N_4999,N_4767);
nor U7039 (N_7039,N_5031,N_4274);
nor U7040 (N_7040,N_5643,N_4634);
nand U7041 (N_7041,N_5617,N_4302);
and U7042 (N_7042,N_5341,N_5351);
nor U7043 (N_7043,N_4867,N_4353);
and U7044 (N_7044,N_5445,N_4557);
nor U7045 (N_7045,N_5911,N_5001);
nand U7046 (N_7046,N_4895,N_5859);
or U7047 (N_7047,N_5270,N_4481);
and U7048 (N_7048,N_4414,N_4594);
and U7049 (N_7049,N_5910,N_5188);
and U7050 (N_7050,N_4500,N_4959);
and U7051 (N_7051,N_5438,N_4761);
and U7052 (N_7052,N_5740,N_4839);
and U7053 (N_7053,N_5334,N_4104);
nor U7054 (N_7054,N_4213,N_4065);
or U7055 (N_7055,N_5226,N_5959);
or U7056 (N_7056,N_4174,N_5962);
nor U7057 (N_7057,N_4093,N_4027);
and U7058 (N_7058,N_5292,N_4175);
nand U7059 (N_7059,N_5127,N_5313);
nor U7060 (N_7060,N_5091,N_5052);
nand U7061 (N_7061,N_4874,N_4308);
or U7062 (N_7062,N_4112,N_4088);
and U7063 (N_7063,N_4505,N_5148);
xnor U7064 (N_7064,N_4917,N_4594);
or U7065 (N_7065,N_4109,N_5297);
nand U7066 (N_7066,N_5977,N_5978);
and U7067 (N_7067,N_5229,N_5503);
and U7068 (N_7068,N_4680,N_5767);
or U7069 (N_7069,N_4118,N_5891);
or U7070 (N_7070,N_5743,N_5304);
and U7071 (N_7071,N_4389,N_4320);
and U7072 (N_7072,N_5945,N_5864);
nand U7073 (N_7073,N_4607,N_5903);
nor U7074 (N_7074,N_5487,N_4274);
or U7075 (N_7075,N_5366,N_4950);
or U7076 (N_7076,N_4595,N_4524);
nor U7077 (N_7077,N_4615,N_5210);
and U7078 (N_7078,N_4937,N_5379);
nor U7079 (N_7079,N_5819,N_5752);
and U7080 (N_7080,N_5737,N_4796);
and U7081 (N_7081,N_4566,N_4128);
nor U7082 (N_7082,N_5329,N_5132);
nor U7083 (N_7083,N_5731,N_4205);
or U7084 (N_7084,N_5948,N_4959);
or U7085 (N_7085,N_4430,N_5437);
and U7086 (N_7086,N_4689,N_5697);
or U7087 (N_7087,N_5943,N_5124);
nand U7088 (N_7088,N_4625,N_4471);
and U7089 (N_7089,N_5481,N_5980);
nand U7090 (N_7090,N_5056,N_5388);
or U7091 (N_7091,N_4653,N_4939);
nand U7092 (N_7092,N_5061,N_5619);
or U7093 (N_7093,N_4626,N_5414);
xor U7094 (N_7094,N_4737,N_4773);
and U7095 (N_7095,N_4447,N_5946);
nand U7096 (N_7096,N_5870,N_5279);
nor U7097 (N_7097,N_5346,N_4650);
nor U7098 (N_7098,N_5484,N_5217);
or U7099 (N_7099,N_5484,N_4351);
nand U7100 (N_7100,N_4432,N_5201);
nand U7101 (N_7101,N_5745,N_5420);
or U7102 (N_7102,N_5793,N_4603);
and U7103 (N_7103,N_4448,N_4378);
nand U7104 (N_7104,N_4303,N_4967);
or U7105 (N_7105,N_4573,N_5491);
or U7106 (N_7106,N_4374,N_4711);
and U7107 (N_7107,N_5587,N_5496);
nand U7108 (N_7108,N_5781,N_4241);
and U7109 (N_7109,N_4729,N_5152);
and U7110 (N_7110,N_5761,N_4074);
and U7111 (N_7111,N_5606,N_5104);
and U7112 (N_7112,N_4768,N_4124);
and U7113 (N_7113,N_4308,N_5467);
and U7114 (N_7114,N_4138,N_5905);
and U7115 (N_7115,N_4590,N_4939);
nor U7116 (N_7116,N_5882,N_4731);
xor U7117 (N_7117,N_5464,N_5029);
or U7118 (N_7118,N_5668,N_4577);
nor U7119 (N_7119,N_4315,N_4593);
nor U7120 (N_7120,N_5045,N_5695);
nor U7121 (N_7121,N_4207,N_5304);
nand U7122 (N_7122,N_5582,N_4257);
nand U7123 (N_7123,N_5207,N_4725);
nor U7124 (N_7124,N_5946,N_5036);
nand U7125 (N_7125,N_4586,N_4683);
nor U7126 (N_7126,N_4776,N_4484);
or U7127 (N_7127,N_5253,N_4810);
or U7128 (N_7128,N_4463,N_5240);
and U7129 (N_7129,N_5898,N_5632);
and U7130 (N_7130,N_5348,N_5598);
and U7131 (N_7131,N_4435,N_4564);
nor U7132 (N_7132,N_5059,N_4414);
nor U7133 (N_7133,N_4457,N_5862);
or U7134 (N_7134,N_5893,N_5432);
nand U7135 (N_7135,N_4190,N_5998);
and U7136 (N_7136,N_5087,N_5370);
nand U7137 (N_7137,N_5800,N_4636);
nand U7138 (N_7138,N_5468,N_5849);
or U7139 (N_7139,N_5955,N_5499);
or U7140 (N_7140,N_5426,N_4433);
nor U7141 (N_7141,N_4227,N_4068);
nand U7142 (N_7142,N_4463,N_4029);
and U7143 (N_7143,N_4640,N_4742);
or U7144 (N_7144,N_5898,N_4607);
xnor U7145 (N_7145,N_4596,N_4604);
nand U7146 (N_7146,N_4739,N_5015);
and U7147 (N_7147,N_4231,N_5588);
xnor U7148 (N_7148,N_5243,N_4406);
nor U7149 (N_7149,N_5712,N_5470);
or U7150 (N_7150,N_5160,N_4290);
and U7151 (N_7151,N_5133,N_4886);
nand U7152 (N_7152,N_4676,N_4992);
xor U7153 (N_7153,N_5221,N_4268);
nor U7154 (N_7154,N_4511,N_5422);
xor U7155 (N_7155,N_5120,N_5949);
and U7156 (N_7156,N_4085,N_5531);
xor U7157 (N_7157,N_5591,N_5119);
or U7158 (N_7158,N_5519,N_4005);
nor U7159 (N_7159,N_4788,N_4696);
and U7160 (N_7160,N_5893,N_4993);
nand U7161 (N_7161,N_5047,N_5129);
or U7162 (N_7162,N_4160,N_5410);
nor U7163 (N_7163,N_5585,N_5211);
and U7164 (N_7164,N_4642,N_4817);
nor U7165 (N_7165,N_4557,N_4424);
or U7166 (N_7166,N_4855,N_4490);
nor U7167 (N_7167,N_4609,N_4299);
nand U7168 (N_7168,N_5262,N_4976);
nor U7169 (N_7169,N_5533,N_5585);
or U7170 (N_7170,N_5777,N_5422);
and U7171 (N_7171,N_4892,N_4943);
or U7172 (N_7172,N_5656,N_5462);
nand U7173 (N_7173,N_5396,N_4878);
nor U7174 (N_7174,N_4820,N_5424);
or U7175 (N_7175,N_4472,N_5222);
nand U7176 (N_7176,N_4038,N_4298);
nand U7177 (N_7177,N_5436,N_5964);
nand U7178 (N_7178,N_5715,N_5169);
and U7179 (N_7179,N_5498,N_4480);
nor U7180 (N_7180,N_4586,N_5751);
nor U7181 (N_7181,N_5406,N_5056);
nand U7182 (N_7182,N_4889,N_4615);
or U7183 (N_7183,N_4596,N_5077);
nand U7184 (N_7184,N_4003,N_4620);
nand U7185 (N_7185,N_4764,N_4201);
nand U7186 (N_7186,N_4003,N_5522);
nand U7187 (N_7187,N_4219,N_4074);
nand U7188 (N_7188,N_5609,N_5716);
and U7189 (N_7189,N_4430,N_5532);
nand U7190 (N_7190,N_4785,N_5290);
and U7191 (N_7191,N_4369,N_4544);
and U7192 (N_7192,N_5167,N_4723);
nand U7193 (N_7193,N_4796,N_4854);
or U7194 (N_7194,N_4263,N_4303);
and U7195 (N_7195,N_5592,N_5431);
xnor U7196 (N_7196,N_5453,N_4160);
or U7197 (N_7197,N_4622,N_4429);
nor U7198 (N_7198,N_5834,N_4028);
and U7199 (N_7199,N_4228,N_4888);
and U7200 (N_7200,N_5296,N_5728);
nor U7201 (N_7201,N_5842,N_4884);
and U7202 (N_7202,N_5785,N_5458);
or U7203 (N_7203,N_4663,N_4009);
and U7204 (N_7204,N_4376,N_5334);
nand U7205 (N_7205,N_4184,N_4170);
nand U7206 (N_7206,N_5646,N_5674);
nor U7207 (N_7207,N_4979,N_5155);
nand U7208 (N_7208,N_4346,N_5624);
nand U7209 (N_7209,N_4843,N_4776);
or U7210 (N_7210,N_5460,N_5666);
nand U7211 (N_7211,N_4025,N_5243);
and U7212 (N_7212,N_4312,N_4246);
and U7213 (N_7213,N_4570,N_4625);
nand U7214 (N_7214,N_4738,N_5036);
nand U7215 (N_7215,N_4686,N_5724);
and U7216 (N_7216,N_4711,N_5779);
or U7217 (N_7217,N_4958,N_4057);
and U7218 (N_7218,N_4691,N_4492);
and U7219 (N_7219,N_5986,N_4146);
xor U7220 (N_7220,N_5465,N_4848);
nor U7221 (N_7221,N_5755,N_5846);
and U7222 (N_7222,N_4500,N_4427);
nor U7223 (N_7223,N_5817,N_5422);
nand U7224 (N_7224,N_5489,N_4801);
nand U7225 (N_7225,N_5919,N_4843);
or U7226 (N_7226,N_4116,N_5657);
nand U7227 (N_7227,N_4815,N_4364);
nand U7228 (N_7228,N_4689,N_5534);
nor U7229 (N_7229,N_4542,N_5640);
nor U7230 (N_7230,N_5157,N_4057);
or U7231 (N_7231,N_5566,N_4695);
nand U7232 (N_7232,N_5898,N_5130);
nand U7233 (N_7233,N_4621,N_4093);
and U7234 (N_7234,N_5011,N_5206);
and U7235 (N_7235,N_4603,N_4702);
nor U7236 (N_7236,N_4779,N_4536);
nand U7237 (N_7237,N_4217,N_5376);
nor U7238 (N_7238,N_4751,N_5225);
nor U7239 (N_7239,N_4922,N_5353);
nand U7240 (N_7240,N_4648,N_5998);
and U7241 (N_7241,N_5632,N_4858);
nor U7242 (N_7242,N_4962,N_4738);
xnor U7243 (N_7243,N_5988,N_5062);
or U7244 (N_7244,N_5751,N_5264);
nand U7245 (N_7245,N_4424,N_4419);
and U7246 (N_7246,N_5431,N_4902);
nor U7247 (N_7247,N_4110,N_4594);
nor U7248 (N_7248,N_5102,N_5717);
or U7249 (N_7249,N_5537,N_5866);
or U7250 (N_7250,N_5806,N_4731);
xor U7251 (N_7251,N_5013,N_5359);
and U7252 (N_7252,N_4940,N_5076);
and U7253 (N_7253,N_4847,N_4383);
and U7254 (N_7254,N_5000,N_4339);
or U7255 (N_7255,N_5338,N_5989);
or U7256 (N_7256,N_4865,N_4417);
and U7257 (N_7257,N_5475,N_4185);
and U7258 (N_7258,N_4661,N_5730);
nand U7259 (N_7259,N_4257,N_4291);
and U7260 (N_7260,N_4591,N_5736);
nand U7261 (N_7261,N_4459,N_4927);
nand U7262 (N_7262,N_4914,N_5065);
nor U7263 (N_7263,N_5967,N_4816);
or U7264 (N_7264,N_4342,N_5151);
or U7265 (N_7265,N_5166,N_4082);
or U7266 (N_7266,N_5063,N_5773);
nand U7267 (N_7267,N_4173,N_4121);
and U7268 (N_7268,N_5093,N_4088);
nor U7269 (N_7269,N_4536,N_5531);
nor U7270 (N_7270,N_4493,N_4265);
nor U7271 (N_7271,N_4716,N_4726);
or U7272 (N_7272,N_4197,N_4185);
and U7273 (N_7273,N_4034,N_4080);
nor U7274 (N_7274,N_5868,N_4726);
and U7275 (N_7275,N_5516,N_5616);
xor U7276 (N_7276,N_5489,N_5037);
or U7277 (N_7277,N_5212,N_4784);
or U7278 (N_7278,N_4215,N_5502);
and U7279 (N_7279,N_5260,N_5181);
nand U7280 (N_7280,N_5486,N_5688);
nand U7281 (N_7281,N_4791,N_4371);
nor U7282 (N_7282,N_4101,N_5926);
nor U7283 (N_7283,N_5696,N_4246);
nand U7284 (N_7284,N_4338,N_4251);
or U7285 (N_7285,N_4796,N_4936);
and U7286 (N_7286,N_4404,N_4110);
or U7287 (N_7287,N_4312,N_5404);
nor U7288 (N_7288,N_5954,N_4478);
nor U7289 (N_7289,N_4056,N_4344);
or U7290 (N_7290,N_4684,N_4665);
or U7291 (N_7291,N_5860,N_4236);
or U7292 (N_7292,N_4897,N_5779);
or U7293 (N_7293,N_5722,N_5840);
nor U7294 (N_7294,N_5117,N_5724);
and U7295 (N_7295,N_4229,N_5385);
and U7296 (N_7296,N_5216,N_5887);
nand U7297 (N_7297,N_4211,N_4829);
and U7298 (N_7298,N_5941,N_5509);
nor U7299 (N_7299,N_4762,N_5478);
and U7300 (N_7300,N_4978,N_5260);
nor U7301 (N_7301,N_5217,N_4276);
or U7302 (N_7302,N_5529,N_5019);
nor U7303 (N_7303,N_4242,N_4617);
nand U7304 (N_7304,N_4581,N_5451);
nand U7305 (N_7305,N_5981,N_5523);
nand U7306 (N_7306,N_5749,N_4986);
nand U7307 (N_7307,N_5527,N_4486);
nor U7308 (N_7308,N_5430,N_5521);
nor U7309 (N_7309,N_5119,N_5497);
nor U7310 (N_7310,N_5544,N_5853);
nor U7311 (N_7311,N_4563,N_4255);
nor U7312 (N_7312,N_5496,N_5744);
or U7313 (N_7313,N_4882,N_4238);
nand U7314 (N_7314,N_4053,N_4288);
and U7315 (N_7315,N_4099,N_5335);
or U7316 (N_7316,N_4754,N_4888);
nor U7317 (N_7317,N_4696,N_5230);
nor U7318 (N_7318,N_4901,N_4709);
nor U7319 (N_7319,N_5717,N_5896);
or U7320 (N_7320,N_4607,N_5563);
or U7321 (N_7321,N_5627,N_4060);
nor U7322 (N_7322,N_4447,N_5233);
nand U7323 (N_7323,N_5547,N_4157);
nor U7324 (N_7324,N_5053,N_4824);
nand U7325 (N_7325,N_5679,N_5466);
nand U7326 (N_7326,N_5315,N_4317);
or U7327 (N_7327,N_4032,N_4715);
or U7328 (N_7328,N_4950,N_5471);
nor U7329 (N_7329,N_4236,N_5388);
nor U7330 (N_7330,N_5513,N_5136);
or U7331 (N_7331,N_4624,N_5801);
or U7332 (N_7332,N_4911,N_5688);
or U7333 (N_7333,N_5269,N_5923);
and U7334 (N_7334,N_4577,N_5178);
and U7335 (N_7335,N_4745,N_5228);
nand U7336 (N_7336,N_5857,N_5565);
nor U7337 (N_7337,N_5739,N_4008);
nand U7338 (N_7338,N_4509,N_4275);
and U7339 (N_7339,N_5360,N_5903);
and U7340 (N_7340,N_5560,N_4718);
nand U7341 (N_7341,N_4997,N_4540);
or U7342 (N_7342,N_5726,N_4825);
or U7343 (N_7343,N_4489,N_4120);
nand U7344 (N_7344,N_5990,N_5050);
and U7345 (N_7345,N_5754,N_5020);
and U7346 (N_7346,N_5937,N_5985);
nand U7347 (N_7347,N_4865,N_5904);
or U7348 (N_7348,N_4477,N_4613);
nor U7349 (N_7349,N_4320,N_4453);
nor U7350 (N_7350,N_4062,N_5888);
and U7351 (N_7351,N_4634,N_5937);
nor U7352 (N_7352,N_4092,N_5148);
nand U7353 (N_7353,N_4327,N_5510);
and U7354 (N_7354,N_5154,N_5119);
nand U7355 (N_7355,N_5761,N_4958);
nand U7356 (N_7356,N_4236,N_4201);
or U7357 (N_7357,N_5184,N_4559);
or U7358 (N_7358,N_4620,N_4358);
and U7359 (N_7359,N_4758,N_4351);
nor U7360 (N_7360,N_5647,N_5965);
nor U7361 (N_7361,N_5373,N_5119);
nand U7362 (N_7362,N_4306,N_4469);
and U7363 (N_7363,N_4004,N_5285);
nor U7364 (N_7364,N_4047,N_5488);
nand U7365 (N_7365,N_4963,N_5002);
or U7366 (N_7366,N_4124,N_5246);
nor U7367 (N_7367,N_4724,N_5021);
nor U7368 (N_7368,N_5654,N_4832);
or U7369 (N_7369,N_4185,N_4160);
nor U7370 (N_7370,N_5555,N_4623);
nor U7371 (N_7371,N_5711,N_4204);
nand U7372 (N_7372,N_5955,N_5652);
and U7373 (N_7373,N_4084,N_4872);
and U7374 (N_7374,N_5093,N_4831);
and U7375 (N_7375,N_5088,N_4706);
and U7376 (N_7376,N_5719,N_4629);
nand U7377 (N_7377,N_5102,N_5666);
nand U7378 (N_7378,N_4824,N_5002);
or U7379 (N_7379,N_4538,N_5066);
nand U7380 (N_7380,N_4154,N_4182);
nor U7381 (N_7381,N_4422,N_5991);
and U7382 (N_7382,N_5619,N_4897);
and U7383 (N_7383,N_4927,N_4142);
or U7384 (N_7384,N_5186,N_4371);
or U7385 (N_7385,N_4704,N_4726);
nand U7386 (N_7386,N_4985,N_5661);
xor U7387 (N_7387,N_5745,N_5266);
and U7388 (N_7388,N_4899,N_5806);
or U7389 (N_7389,N_4359,N_5691);
xor U7390 (N_7390,N_5626,N_4924);
or U7391 (N_7391,N_4017,N_4941);
nand U7392 (N_7392,N_4705,N_4736);
and U7393 (N_7393,N_5132,N_5307);
nor U7394 (N_7394,N_4842,N_5935);
or U7395 (N_7395,N_4839,N_5465);
nor U7396 (N_7396,N_5878,N_5238);
nand U7397 (N_7397,N_4873,N_4620);
or U7398 (N_7398,N_5338,N_5452);
nor U7399 (N_7399,N_4565,N_5040);
nor U7400 (N_7400,N_4269,N_5148);
or U7401 (N_7401,N_5049,N_4895);
nand U7402 (N_7402,N_5581,N_5347);
nor U7403 (N_7403,N_5490,N_4935);
or U7404 (N_7404,N_4455,N_4016);
or U7405 (N_7405,N_4633,N_5384);
and U7406 (N_7406,N_4037,N_5175);
or U7407 (N_7407,N_4385,N_4902);
or U7408 (N_7408,N_4115,N_4941);
nand U7409 (N_7409,N_5745,N_5552);
nor U7410 (N_7410,N_5486,N_5662);
nor U7411 (N_7411,N_4861,N_4600);
and U7412 (N_7412,N_4042,N_5424);
and U7413 (N_7413,N_5588,N_5180);
nand U7414 (N_7414,N_4772,N_5580);
nor U7415 (N_7415,N_4361,N_4061);
and U7416 (N_7416,N_4567,N_5591);
or U7417 (N_7417,N_5228,N_4030);
and U7418 (N_7418,N_5657,N_5250);
and U7419 (N_7419,N_4917,N_4740);
nor U7420 (N_7420,N_4751,N_5866);
or U7421 (N_7421,N_4411,N_4657);
and U7422 (N_7422,N_4842,N_4792);
or U7423 (N_7423,N_5142,N_5910);
nor U7424 (N_7424,N_5319,N_5754);
or U7425 (N_7425,N_4861,N_4944);
and U7426 (N_7426,N_5948,N_5706);
nand U7427 (N_7427,N_4851,N_4642);
nand U7428 (N_7428,N_4157,N_5031);
nor U7429 (N_7429,N_4663,N_5928);
and U7430 (N_7430,N_5063,N_4730);
nor U7431 (N_7431,N_4155,N_5351);
and U7432 (N_7432,N_4234,N_5890);
or U7433 (N_7433,N_5771,N_5474);
and U7434 (N_7434,N_4631,N_5853);
and U7435 (N_7435,N_5672,N_4398);
nand U7436 (N_7436,N_4739,N_4648);
or U7437 (N_7437,N_4829,N_4605);
nand U7438 (N_7438,N_5165,N_4190);
or U7439 (N_7439,N_5092,N_4369);
and U7440 (N_7440,N_5392,N_5143);
nor U7441 (N_7441,N_4189,N_4104);
nor U7442 (N_7442,N_5357,N_5740);
or U7443 (N_7443,N_5542,N_5478);
nor U7444 (N_7444,N_4450,N_5112);
and U7445 (N_7445,N_5807,N_4636);
or U7446 (N_7446,N_5431,N_5148);
nor U7447 (N_7447,N_5745,N_5729);
or U7448 (N_7448,N_5708,N_5056);
or U7449 (N_7449,N_5774,N_5160);
nor U7450 (N_7450,N_5612,N_5445);
or U7451 (N_7451,N_5806,N_4638);
nor U7452 (N_7452,N_5632,N_4632);
or U7453 (N_7453,N_4114,N_4607);
or U7454 (N_7454,N_5588,N_4182);
nand U7455 (N_7455,N_4828,N_4884);
and U7456 (N_7456,N_4072,N_4837);
nand U7457 (N_7457,N_5628,N_4356);
or U7458 (N_7458,N_4525,N_5853);
nand U7459 (N_7459,N_4095,N_5626);
nor U7460 (N_7460,N_5048,N_5545);
nor U7461 (N_7461,N_5820,N_4150);
and U7462 (N_7462,N_5880,N_5411);
or U7463 (N_7463,N_4130,N_5815);
nand U7464 (N_7464,N_4235,N_5403);
or U7465 (N_7465,N_4248,N_5876);
and U7466 (N_7466,N_4285,N_4529);
and U7467 (N_7467,N_4477,N_4325);
nor U7468 (N_7468,N_4747,N_4662);
and U7469 (N_7469,N_5505,N_5859);
or U7470 (N_7470,N_4113,N_5714);
and U7471 (N_7471,N_5999,N_5775);
and U7472 (N_7472,N_4971,N_5513);
and U7473 (N_7473,N_4528,N_5831);
nor U7474 (N_7474,N_5716,N_5590);
or U7475 (N_7475,N_5912,N_5199);
or U7476 (N_7476,N_4234,N_5779);
or U7477 (N_7477,N_5829,N_5053);
nor U7478 (N_7478,N_5492,N_4943);
nor U7479 (N_7479,N_5656,N_5400);
or U7480 (N_7480,N_5017,N_4824);
or U7481 (N_7481,N_4167,N_5796);
and U7482 (N_7482,N_5308,N_4039);
nor U7483 (N_7483,N_4736,N_4215);
nand U7484 (N_7484,N_5031,N_4666);
nand U7485 (N_7485,N_5223,N_4103);
nand U7486 (N_7486,N_4417,N_4510);
nor U7487 (N_7487,N_5933,N_5744);
and U7488 (N_7488,N_4516,N_4785);
nand U7489 (N_7489,N_4644,N_4160);
nor U7490 (N_7490,N_4192,N_4549);
and U7491 (N_7491,N_4816,N_4326);
nor U7492 (N_7492,N_5627,N_5712);
nand U7493 (N_7493,N_5263,N_5793);
nor U7494 (N_7494,N_4415,N_5493);
nor U7495 (N_7495,N_4327,N_5857);
nor U7496 (N_7496,N_5606,N_5426);
or U7497 (N_7497,N_4828,N_5004);
nand U7498 (N_7498,N_4441,N_4072);
xor U7499 (N_7499,N_4792,N_4286);
nor U7500 (N_7500,N_5242,N_4316);
and U7501 (N_7501,N_4396,N_4705);
nor U7502 (N_7502,N_4311,N_4073);
and U7503 (N_7503,N_4065,N_5199);
and U7504 (N_7504,N_5398,N_5416);
nand U7505 (N_7505,N_5603,N_4035);
nor U7506 (N_7506,N_5271,N_5721);
or U7507 (N_7507,N_5367,N_4475);
nor U7508 (N_7508,N_5505,N_4489);
nand U7509 (N_7509,N_4342,N_5967);
and U7510 (N_7510,N_4128,N_4805);
nand U7511 (N_7511,N_4254,N_5313);
nor U7512 (N_7512,N_5700,N_5401);
nor U7513 (N_7513,N_5283,N_5367);
and U7514 (N_7514,N_5947,N_4682);
nor U7515 (N_7515,N_5719,N_5340);
nand U7516 (N_7516,N_4674,N_4550);
nand U7517 (N_7517,N_5058,N_4578);
nor U7518 (N_7518,N_4175,N_5305);
nand U7519 (N_7519,N_5770,N_5324);
xor U7520 (N_7520,N_5254,N_4744);
and U7521 (N_7521,N_4678,N_4007);
nor U7522 (N_7522,N_4745,N_5293);
or U7523 (N_7523,N_4708,N_5569);
nand U7524 (N_7524,N_5438,N_5534);
nand U7525 (N_7525,N_4609,N_4175);
nor U7526 (N_7526,N_4419,N_4487);
nor U7527 (N_7527,N_5338,N_4921);
nand U7528 (N_7528,N_5097,N_4159);
nand U7529 (N_7529,N_5031,N_5741);
nand U7530 (N_7530,N_5636,N_5768);
nand U7531 (N_7531,N_5045,N_4868);
and U7532 (N_7532,N_5395,N_5925);
nor U7533 (N_7533,N_5572,N_4062);
nor U7534 (N_7534,N_5792,N_5174);
nor U7535 (N_7535,N_5127,N_5856);
and U7536 (N_7536,N_4805,N_4618);
nand U7537 (N_7537,N_5312,N_4664);
or U7538 (N_7538,N_4300,N_4760);
nor U7539 (N_7539,N_4227,N_4568);
or U7540 (N_7540,N_4913,N_5545);
xor U7541 (N_7541,N_5820,N_4936);
nand U7542 (N_7542,N_5275,N_5086);
and U7543 (N_7543,N_4195,N_4970);
and U7544 (N_7544,N_4646,N_4777);
and U7545 (N_7545,N_5266,N_4794);
or U7546 (N_7546,N_5501,N_5888);
nor U7547 (N_7547,N_4952,N_5610);
and U7548 (N_7548,N_4922,N_4674);
nand U7549 (N_7549,N_4519,N_5244);
nor U7550 (N_7550,N_4234,N_5295);
and U7551 (N_7551,N_4213,N_4759);
and U7552 (N_7552,N_5972,N_4092);
and U7553 (N_7553,N_5501,N_5664);
nor U7554 (N_7554,N_5162,N_4290);
nand U7555 (N_7555,N_4890,N_5037);
or U7556 (N_7556,N_4774,N_4117);
nand U7557 (N_7557,N_4412,N_5089);
nand U7558 (N_7558,N_4643,N_4488);
nand U7559 (N_7559,N_4625,N_5884);
xnor U7560 (N_7560,N_4320,N_5644);
nand U7561 (N_7561,N_4204,N_5640);
or U7562 (N_7562,N_4980,N_4608);
or U7563 (N_7563,N_4514,N_4947);
and U7564 (N_7564,N_5982,N_5681);
nand U7565 (N_7565,N_5335,N_5448);
nor U7566 (N_7566,N_4093,N_5886);
nand U7567 (N_7567,N_4436,N_5092);
nand U7568 (N_7568,N_4057,N_5049);
or U7569 (N_7569,N_4005,N_5087);
or U7570 (N_7570,N_5063,N_5561);
or U7571 (N_7571,N_5227,N_4360);
nor U7572 (N_7572,N_4027,N_5980);
or U7573 (N_7573,N_5425,N_4887);
or U7574 (N_7574,N_5098,N_4275);
nor U7575 (N_7575,N_5173,N_5487);
and U7576 (N_7576,N_4028,N_4569);
or U7577 (N_7577,N_5789,N_4250);
nand U7578 (N_7578,N_4764,N_5503);
nand U7579 (N_7579,N_5671,N_5080);
and U7580 (N_7580,N_4627,N_4252);
nand U7581 (N_7581,N_5655,N_5549);
and U7582 (N_7582,N_4529,N_4714);
nand U7583 (N_7583,N_4245,N_4876);
or U7584 (N_7584,N_5198,N_4475);
nand U7585 (N_7585,N_4650,N_4116);
or U7586 (N_7586,N_4743,N_5795);
or U7587 (N_7587,N_4212,N_4292);
and U7588 (N_7588,N_5495,N_4388);
or U7589 (N_7589,N_5145,N_5244);
or U7590 (N_7590,N_5652,N_5337);
or U7591 (N_7591,N_5430,N_4788);
nor U7592 (N_7592,N_5375,N_5767);
or U7593 (N_7593,N_4888,N_5815);
nor U7594 (N_7594,N_5917,N_5560);
and U7595 (N_7595,N_4919,N_4262);
nor U7596 (N_7596,N_5114,N_4441);
nand U7597 (N_7597,N_4168,N_4421);
nor U7598 (N_7598,N_5069,N_4879);
nor U7599 (N_7599,N_4000,N_5264);
and U7600 (N_7600,N_5411,N_5959);
nor U7601 (N_7601,N_4579,N_5426);
or U7602 (N_7602,N_5193,N_4795);
nand U7603 (N_7603,N_5733,N_4740);
nand U7604 (N_7604,N_5866,N_5396);
and U7605 (N_7605,N_4537,N_5273);
and U7606 (N_7606,N_5472,N_4290);
or U7607 (N_7607,N_5331,N_4990);
nand U7608 (N_7608,N_4255,N_5191);
nand U7609 (N_7609,N_4921,N_5689);
and U7610 (N_7610,N_4118,N_5727);
nand U7611 (N_7611,N_4680,N_5919);
or U7612 (N_7612,N_5325,N_4994);
nor U7613 (N_7613,N_5131,N_5546);
nand U7614 (N_7614,N_5282,N_5611);
nor U7615 (N_7615,N_5438,N_5055);
and U7616 (N_7616,N_4675,N_5585);
and U7617 (N_7617,N_5714,N_5890);
or U7618 (N_7618,N_4881,N_5739);
or U7619 (N_7619,N_4170,N_5354);
xor U7620 (N_7620,N_5878,N_5344);
nand U7621 (N_7621,N_4922,N_4086);
nor U7622 (N_7622,N_5428,N_4719);
or U7623 (N_7623,N_4643,N_4104);
and U7624 (N_7624,N_5719,N_4065);
nand U7625 (N_7625,N_4101,N_4342);
nor U7626 (N_7626,N_4014,N_5563);
or U7627 (N_7627,N_4068,N_4846);
nor U7628 (N_7628,N_4398,N_4815);
nor U7629 (N_7629,N_5635,N_5285);
or U7630 (N_7630,N_5510,N_5525);
and U7631 (N_7631,N_5970,N_5579);
or U7632 (N_7632,N_5455,N_4160);
or U7633 (N_7633,N_5088,N_5817);
or U7634 (N_7634,N_5289,N_4441);
nand U7635 (N_7635,N_4943,N_4476);
and U7636 (N_7636,N_5668,N_4126);
nor U7637 (N_7637,N_4517,N_5774);
nand U7638 (N_7638,N_5889,N_4814);
nand U7639 (N_7639,N_4361,N_4999);
nand U7640 (N_7640,N_4618,N_5802);
nor U7641 (N_7641,N_5418,N_4605);
xor U7642 (N_7642,N_5784,N_5714);
or U7643 (N_7643,N_5091,N_4582);
or U7644 (N_7644,N_4653,N_4620);
and U7645 (N_7645,N_4596,N_4019);
or U7646 (N_7646,N_4851,N_4436);
or U7647 (N_7647,N_4914,N_5669);
nand U7648 (N_7648,N_5321,N_4873);
nor U7649 (N_7649,N_5033,N_4417);
nand U7650 (N_7650,N_5308,N_4493);
nand U7651 (N_7651,N_4200,N_5221);
and U7652 (N_7652,N_4346,N_5644);
nor U7653 (N_7653,N_5857,N_5635);
nor U7654 (N_7654,N_4374,N_4128);
nor U7655 (N_7655,N_5810,N_5850);
and U7656 (N_7656,N_4743,N_5431);
and U7657 (N_7657,N_4190,N_5371);
nor U7658 (N_7658,N_5257,N_5952);
nand U7659 (N_7659,N_4813,N_5204);
nor U7660 (N_7660,N_4944,N_4733);
nand U7661 (N_7661,N_4890,N_5111);
or U7662 (N_7662,N_5363,N_4222);
and U7663 (N_7663,N_4867,N_4747);
nand U7664 (N_7664,N_5040,N_5149);
nor U7665 (N_7665,N_5866,N_5111);
and U7666 (N_7666,N_4332,N_4972);
nor U7667 (N_7667,N_5747,N_5461);
and U7668 (N_7668,N_4817,N_5551);
xor U7669 (N_7669,N_4791,N_5139);
nand U7670 (N_7670,N_5263,N_5865);
xnor U7671 (N_7671,N_5397,N_5631);
and U7672 (N_7672,N_4330,N_5451);
or U7673 (N_7673,N_5040,N_4816);
and U7674 (N_7674,N_4768,N_5805);
nand U7675 (N_7675,N_5519,N_4378);
and U7676 (N_7676,N_4986,N_4411);
and U7677 (N_7677,N_5817,N_4812);
nand U7678 (N_7678,N_5171,N_4136);
nor U7679 (N_7679,N_4544,N_4222);
and U7680 (N_7680,N_4691,N_5123);
and U7681 (N_7681,N_5210,N_5218);
or U7682 (N_7682,N_4116,N_5363);
nand U7683 (N_7683,N_4813,N_5178);
or U7684 (N_7684,N_4644,N_4946);
and U7685 (N_7685,N_4317,N_4781);
nor U7686 (N_7686,N_5953,N_4256);
or U7687 (N_7687,N_4070,N_5894);
or U7688 (N_7688,N_4683,N_4506);
and U7689 (N_7689,N_4815,N_5995);
and U7690 (N_7690,N_5795,N_5972);
nor U7691 (N_7691,N_5037,N_5709);
and U7692 (N_7692,N_4008,N_5620);
or U7693 (N_7693,N_4285,N_4392);
nor U7694 (N_7694,N_4726,N_5661);
or U7695 (N_7695,N_5115,N_5073);
and U7696 (N_7696,N_5866,N_5411);
nand U7697 (N_7697,N_4582,N_4546);
or U7698 (N_7698,N_5804,N_5483);
nand U7699 (N_7699,N_5544,N_5572);
nand U7700 (N_7700,N_5896,N_5495);
or U7701 (N_7701,N_4505,N_4193);
nand U7702 (N_7702,N_5225,N_5261);
and U7703 (N_7703,N_5957,N_5222);
nor U7704 (N_7704,N_4861,N_4055);
and U7705 (N_7705,N_4076,N_5521);
or U7706 (N_7706,N_5818,N_4743);
nor U7707 (N_7707,N_4555,N_4310);
nand U7708 (N_7708,N_4971,N_5133);
or U7709 (N_7709,N_4329,N_4007);
nor U7710 (N_7710,N_4132,N_5677);
nand U7711 (N_7711,N_5979,N_4459);
or U7712 (N_7712,N_5671,N_5789);
xnor U7713 (N_7713,N_4851,N_4090);
nand U7714 (N_7714,N_4164,N_5483);
nand U7715 (N_7715,N_5258,N_5873);
nor U7716 (N_7716,N_4061,N_5019);
nand U7717 (N_7717,N_5346,N_5468);
and U7718 (N_7718,N_5043,N_4286);
nor U7719 (N_7719,N_5774,N_4775);
nand U7720 (N_7720,N_5613,N_4270);
nor U7721 (N_7721,N_5998,N_5271);
and U7722 (N_7722,N_4210,N_4524);
nand U7723 (N_7723,N_4413,N_4722);
and U7724 (N_7724,N_4859,N_5381);
and U7725 (N_7725,N_4996,N_5829);
or U7726 (N_7726,N_5291,N_5039);
and U7727 (N_7727,N_5922,N_4871);
nor U7728 (N_7728,N_5315,N_4945);
nand U7729 (N_7729,N_4374,N_4199);
nand U7730 (N_7730,N_5190,N_4636);
and U7731 (N_7731,N_5600,N_5705);
nor U7732 (N_7732,N_4962,N_5574);
nor U7733 (N_7733,N_4470,N_4045);
or U7734 (N_7734,N_4723,N_5860);
nand U7735 (N_7735,N_5109,N_4661);
nand U7736 (N_7736,N_5923,N_4344);
and U7737 (N_7737,N_4053,N_4063);
and U7738 (N_7738,N_4260,N_5225);
nor U7739 (N_7739,N_4966,N_5804);
nor U7740 (N_7740,N_5466,N_5003);
or U7741 (N_7741,N_4804,N_5298);
nor U7742 (N_7742,N_4581,N_4693);
nand U7743 (N_7743,N_4366,N_4989);
or U7744 (N_7744,N_4634,N_4718);
nand U7745 (N_7745,N_4175,N_5997);
nand U7746 (N_7746,N_4667,N_5211);
and U7747 (N_7747,N_5565,N_4658);
and U7748 (N_7748,N_4265,N_4982);
or U7749 (N_7749,N_5779,N_4086);
or U7750 (N_7750,N_5832,N_4294);
nor U7751 (N_7751,N_4923,N_4395);
or U7752 (N_7752,N_5997,N_4911);
nand U7753 (N_7753,N_4399,N_5245);
nor U7754 (N_7754,N_5926,N_5325);
xnor U7755 (N_7755,N_5081,N_4400);
nand U7756 (N_7756,N_5982,N_5826);
and U7757 (N_7757,N_5559,N_5637);
or U7758 (N_7758,N_4207,N_5669);
nor U7759 (N_7759,N_4743,N_5956);
nand U7760 (N_7760,N_4234,N_5034);
nand U7761 (N_7761,N_4057,N_5473);
nand U7762 (N_7762,N_5259,N_5444);
or U7763 (N_7763,N_4708,N_5893);
or U7764 (N_7764,N_4209,N_4713);
and U7765 (N_7765,N_4023,N_4452);
and U7766 (N_7766,N_4998,N_4320);
nand U7767 (N_7767,N_5612,N_5203);
nor U7768 (N_7768,N_4055,N_5429);
and U7769 (N_7769,N_5859,N_5327);
or U7770 (N_7770,N_4739,N_4173);
xnor U7771 (N_7771,N_4888,N_4893);
or U7772 (N_7772,N_5482,N_4778);
nor U7773 (N_7773,N_4033,N_5687);
or U7774 (N_7774,N_5057,N_5237);
and U7775 (N_7775,N_4230,N_4704);
nand U7776 (N_7776,N_4618,N_4552);
nor U7777 (N_7777,N_5338,N_4038);
or U7778 (N_7778,N_5811,N_4949);
nor U7779 (N_7779,N_4775,N_5932);
or U7780 (N_7780,N_5460,N_4297);
xor U7781 (N_7781,N_5571,N_4047);
nor U7782 (N_7782,N_5287,N_4746);
and U7783 (N_7783,N_4053,N_5496);
or U7784 (N_7784,N_5845,N_5417);
xnor U7785 (N_7785,N_4096,N_5606);
and U7786 (N_7786,N_5439,N_4119);
nor U7787 (N_7787,N_4376,N_5920);
and U7788 (N_7788,N_5770,N_5480);
and U7789 (N_7789,N_5889,N_5090);
nor U7790 (N_7790,N_4624,N_5237);
xnor U7791 (N_7791,N_5342,N_5136);
and U7792 (N_7792,N_5583,N_4850);
nand U7793 (N_7793,N_4551,N_4899);
and U7794 (N_7794,N_5857,N_5880);
or U7795 (N_7795,N_5563,N_5198);
or U7796 (N_7796,N_5450,N_5287);
and U7797 (N_7797,N_5225,N_5772);
nand U7798 (N_7798,N_5383,N_5724);
nor U7799 (N_7799,N_4387,N_4968);
nor U7800 (N_7800,N_5054,N_4037);
or U7801 (N_7801,N_4144,N_4232);
or U7802 (N_7802,N_5598,N_5346);
and U7803 (N_7803,N_5673,N_5155);
nand U7804 (N_7804,N_4354,N_5370);
or U7805 (N_7805,N_5508,N_5861);
or U7806 (N_7806,N_5385,N_5508);
nor U7807 (N_7807,N_5405,N_4041);
nand U7808 (N_7808,N_5944,N_4866);
nor U7809 (N_7809,N_4515,N_5093);
nor U7810 (N_7810,N_4238,N_4530);
nand U7811 (N_7811,N_4431,N_5331);
or U7812 (N_7812,N_4692,N_4081);
nand U7813 (N_7813,N_4060,N_4972);
or U7814 (N_7814,N_5974,N_4081);
or U7815 (N_7815,N_4395,N_4319);
nor U7816 (N_7816,N_4949,N_5881);
or U7817 (N_7817,N_4922,N_5509);
nand U7818 (N_7818,N_5290,N_4418);
or U7819 (N_7819,N_5940,N_4826);
nand U7820 (N_7820,N_5680,N_4395);
nor U7821 (N_7821,N_4885,N_4822);
nand U7822 (N_7822,N_4576,N_4357);
nor U7823 (N_7823,N_4890,N_5463);
nand U7824 (N_7824,N_4354,N_4318);
nand U7825 (N_7825,N_4094,N_4421);
or U7826 (N_7826,N_4314,N_5999);
nand U7827 (N_7827,N_5250,N_5397);
or U7828 (N_7828,N_5789,N_5990);
nand U7829 (N_7829,N_5710,N_4282);
nor U7830 (N_7830,N_4376,N_5799);
nand U7831 (N_7831,N_4757,N_5490);
or U7832 (N_7832,N_5176,N_4247);
nor U7833 (N_7833,N_4633,N_5605);
and U7834 (N_7834,N_5196,N_4689);
or U7835 (N_7835,N_5766,N_5839);
or U7836 (N_7836,N_5358,N_4473);
or U7837 (N_7837,N_4868,N_5843);
or U7838 (N_7838,N_4158,N_4280);
nand U7839 (N_7839,N_5127,N_5411);
nand U7840 (N_7840,N_4636,N_4756);
and U7841 (N_7841,N_4782,N_4459);
nand U7842 (N_7842,N_4701,N_4036);
nand U7843 (N_7843,N_4081,N_4322);
nand U7844 (N_7844,N_5196,N_5503);
nor U7845 (N_7845,N_5004,N_4150);
and U7846 (N_7846,N_5245,N_5902);
nor U7847 (N_7847,N_4356,N_4060);
and U7848 (N_7848,N_4313,N_4014);
nand U7849 (N_7849,N_4718,N_4128);
and U7850 (N_7850,N_4246,N_4419);
or U7851 (N_7851,N_5940,N_5699);
nand U7852 (N_7852,N_4759,N_4362);
or U7853 (N_7853,N_5894,N_4820);
and U7854 (N_7854,N_5414,N_4371);
and U7855 (N_7855,N_4427,N_5244);
nand U7856 (N_7856,N_5003,N_5670);
nand U7857 (N_7857,N_5240,N_4840);
nor U7858 (N_7858,N_4566,N_5719);
or U7859 (N_7859,N_5727,N_5703);
nor U7860 (N_7860,N_4184,N_5974);
or U7861 (N_7861,N_4018,N_4425);
and U7862 (N_7862,N_5640,N_4313);
or U7863 (N_7863,N_5394,N_4959);
and U7864 (N_7864,N_5951,N_4088);
and U7865 (N_7865,N_5848,N_5506);
nand U7866 (N_7866,N_4774,N_5704);
nand U7867 (N_7867,N_4536,N_5260);
and U7868 (N_7868,N_4006,N_4576);
nor U7869 (N_7869,N_4357,N_4239);
or U7870 (N_7870,N_5699,N_5819);
nor U7871 (N_7871,N_5667,N_5530);
and U7872 (N_7872,N_4360,N_5249);
and U7873 (N_7873,N_5468,N_5705);
or U7874 (N_7874,N_5972,N_4875);
xnor U7875 (N_7875,N_5160,N_5798);
and U7876 (N_7876,N_4028,N_5320);
or U7877 (N_7877,N_5523,N_5896);
or U7878 (N_7878,N_5830,N_5326);
and U7879 (N_7879,N_4663,N_5407);
nand U7880 (N_7880,N_4261,N_4271);
nor U7881 (N_7881,N_5927,N_4913);
or U7882 (N_7882,N_5576,N_5920);
or U7883 (N_7883,N_5131,N_5260);
nor U7884 (N_7884,N_5147,N_4568);
nand U7885 (N_7885,N_5883,N_4540);
xor U7886 (N_7886,N_4361,N_4832);
and U7887 (N_7887,N_4305,N_5618);
nand U7888 (N_7888,N_4329,N_4934);
nand U7889 (N_7889,N_5144,N_5817);
or U7890 (N_7890,N_4049,N_5245);
and U7891 (N_7891,N_4414,N_4326);
and U7892 (N_7892,N_4293,N_5690);
or U7893 (N_7893,N_4480,N_5822);
or U7894 (N_7894,N_4520,N_4500);
nor U7895 (N_7895,N_5593,N_4350);
or U7896 (N_7896,N_4414,N_4787);
nor U7897 (N_7897,N_4505,N_4734);
and U7898 (N_7898,N_4601,N_5807);
and U7899 (N_7899,N_5266,N_4974);
or U7900 (N_7900,N_4298,N_5659);
and U7901 (N_7901,N_4462,N_4571);
nand U7902 (N_7902,N_5653,N_4420);
nor U7903 (N_7903,N_4702,N_5251);
nor U7904 (N_7904,N_4843,N_5111);
or U7905 (N_7905,N_4556,N_5385);
or U7906 (N_7906,N_5835,N_5944);
and U7907 (N_7907,N_4432,N_4693);
or U7908 (N_7908,N_5350,N_4496);
nand U7909 (N_7909,N_5049,N_5640);
and U7910 (N_7910,N_5846,N_5733);
nor U7911 (N_7911,N_4816,N_4689);
or U7912 (N_7912,N_4920,N_4662);
or U7913 (N_7913,N_4739,N_4804);
or U7914 (N_7914,N_5956,N_5273);
and U7915 (N_7915,N_5330,N_5842);
nor U7916 (N_7916,N_4718,N_5964);
or U7917 (N_7917,N_4812,N_5570);
and U7918 (N_7918,N_4915,N_5624);
and U7919 (N_7919,N_5140,N_5619);
and U7920 (N_7920,N_5675,N_4686);
xnor U7921 (N_7921,N_5435,N_5737);
or U7922 (N_7922,N_5425,N_5963);
nand U7923 (N_7923,N_5633,N_5981);
and U7924 (N_7924,N_4706,N_5502);
nor U7925 (N_7925,N_4404,N_5149);
xor U7926 (N_7926,N_4309,N_5795);
nand U7927 (N_7927,N_4689,N_4265);
nand U7928 (N_7928,N_4099,N_5291);
and U7929 (N_7929,N_4038,N_5530);
nand U7930 (N_7930,N_5770,N_5863);
nand U7931 (N_7931,N_4167,N_4154);
nor U7932 (N_7932,N_4267,N_4597);
and U7933 (N_7933,N_4749,N_4480);
or U7934 (N_7934,N_5535,N_4730);
nand U7935 (N_7935,N_4593,N_5879);
and U7936 (N_7936,N_4735,N_5062);
nor U7937 (N_7937,N_5665,N_4123);
or U7938 (N_7938,N_4398,N_5693);
or U7939 (N_7939,N_5575,N_5677);
and U7940 (N_7940,N_4039,N_5162);
or U7941 (N_7941,N_5546,N_5560);
or U7942 (N_7942,N_5609,N_4211);
nor U7943 (N_7943,N_5775,N_4279);
nand U7944 (N_7944,N_5829,N_4588);
xor U7945 (N_7945,N_4758,N_4569);
nor U7946 (N_7946,N_5664,N_5839);
or U7947 (N_7947,N_4672,N_4828);
or U7948 (N_7948,N_5753,N_4821);
nand U7949 (N_7949,N_4853,N_4925);
nor U7950 (N_7950,N_5741,N_4733);
or U7951 (N_7951,N_5968,N_5284);
nand U7952 (N_7952,N_5767,N_4010);
nor U7953 (N_7953,N_4584,N_4367);
and U7954 (N_7954,N_5025,N_4864);
or U7955 (N_7955,N_5869,N_5670);
or U7956 (N_7956,N_4237,N_5290);
and U7957 (N_7957,N_4798,N_5328);
nor U7958 (N_7958,N_5674,N_4686);
or U7959 (N_7959,N_4585,N_5814);
nor U7960 (N_7960,N_5436,N_5635);
nor U7961 (N_7961,N_5846,N_4649);
and U7962 (N_7962,N_5691,N_5959);
or U7963 (N_7963,N_5124,N_4051);
nor U7964 (N_7964,N_4674,N_5782);
nor U7965 (N_7965,N_4977,N_5217);
and U7966 (N_7966,N_5901,N_4490);
nor U7967 (N_7967,N_4251,N_5860);
or U7968 (N_7968,N_5693,N_4690);
and U7969 (N_7969,N_5974,N_4328);
nand U7970 (N_7970,N_4671,N_4267);
nor U7971 (N_7971,N_4566,N_4709);
and U7972 (N_7972,N_5849,N_4148);
or U7973 (N_7973,N_4261,N_4953);
nor U7974 (N_7974,N_4464,N_4778);
nor U7975 (N_7975,N_4744,N_5747);
nor U7976 (N_7976,N_5127,N_4157);
nand U7977 (N_7977,N_4879,N_5835);
nand U7978 (N_7978,N_4807,N_5985);
nand U7979 (N_7979,N_5970,N_5740);
nor U7980 (N_7980,N_4668,N_4899);
nand U7981 (N_7981,N_4979,N_5363);
or U7982 (N_7982,N_4418,N_4206);
or U7983 (N_7983,N_5686,N_4446);
or U7984 (N_7984,N_5016,N_4209);
nand U7985 (N_7985,N_4663,N_5725);
nand U7986 (N_7986,N_4876,N_4095);
nand U7987 (N_7987,N_5363,N_4527);
xnor U7988 (N_7988,N_4106,N_5914);
nand U7989 (N_7989,N_5192,N_4602);
nand U7990 (N_7990,N_5249,N_5270);
nor U7991 (N_7991,N_4412,N_5438);
nor U7992 (N_7992,N_5050,N_5838);
nor U7993 (N_7993,N_5860,N_4694);
or U7994 (N_7994,N_4964,N_5468);
nor U7995 (N_7995,N_4325,N_4711);
and U7996 (N_7996,N_4323,N_5287);
and U7997 (N_7997,N_4636,N_4511);
and U7998 (N_7998,N_4208,N_5008);
nor U7999 (N_7999,N_5164,N_4101);
nor U8000 (N_8000,N_6846,N_7493);
xnor U8001 (N_8001,N_7911,N_6082);
and U8002 (N_8002,N_6802,N_6137);
nand U8003 (N_8003,N_6539,N_7351);
and U8004 (N_8004,N_6132,N_7776);
nand U8005 (N_8005,N_7293,N_7314);
or U8006 (N_8006,N_6217,N_6519);
or U8007 (N_8007,N_7298,N_7604);
nand U8008 (N_8008,N_7942,N_7921);
nand U8009 (N_8009,N_7663,N_7023);
or U8010 (N_8010,N_7737,N_6793);
nor U8011 (N_8011,N_7723,N_6167);
nor U8012 (N_8012,N_7499,N_6529);
nor U8013 (N_8013,N_6530,N_6316);
nand U8014 (N_8014,N_7052,N_6238);
nand U8015 (N_8015,N_7046,N_6555);
nor U8016 (N_8016,N_6885,N_7098);
nand U8017 (N_8017,N_6170,N_7416);
and U8018 (N_8018,N_7773,N_6800);
nand U8019 (N_8019,N_7446,N_7277);
nor U8020 (N_8020,N_7067,N_7016);
nand U8021 (N_8021,N_7585,N_6647);
and U8022 (N_8022,N_6333,N_7848);
nor U8023 (N_8023,N_7906,N_7278);
or U8024 (N_8024,N_6856,N_7506);
or U8025 (N_8025,N_7496,N_6209);
or U8026 (N_8026,N_7486,N_6889);
or U8027 (N_8027,N_6141,N_7320);
nand U8028 (N_8028,N_7321,N_7841);
nand U8029 (N_8029,N_6135,N_6895);
nand U8030 (N_8030,N_7369,N_6504);
nor U8031 (N_8031,N_7478,N_7471);
nand U8032 (N_8032,N_7181,N_7629);
or U8033 (N_8033,N_7466,N_7104);
nand U8034 (N_8034,N_7691,N_7717);
or U8035 (N_8035,N_6868,N_7134);
nor U8036 (N_8036,N_6925,N_6041);
nand U8037 (N_8037,N_7642,N_6438);
and U8038 (N_8038,N_6280,N_7721);
nand U8039 (N_8039,N_6662,N_6129);
nor U8040 (N_8040,N_6317,N_6225);
and U8041 (N_8041,N_7299,N_6271);
nand U8042 (N_8042,N_6327,N_6680);
nand U8043 (N_8043,N_7275,N_6259);
or U8044 (N_8044,N_6377,N_7144);
or U8045 (N_8045,N_7910,N_7583);
nand U8046 (N_8046,N_7756,N_6951);
nor U8047 (N_8047,N_6894,N_7001);
nor U8048 (N_8048,N_7065,N_7334);
nand U8049 (N_8049,N_7532,N_7235);
or U8050 (N_8050,N_7337,N_6696);
and U8051 (N_8051,N_7402,N_6184);
or U8052 (N_8052,N_6248,N_6841);
or U8053 (N_8053,N_6291,N_7959);
or U8054 (N_8054,N_7544,N_7264);
nor U8055 (N_8055,N_7704,N_7409);
and U8056 (N_8056,N_6873,N_6983);
or U8057 (N_8057,N_6422,N_6096);
and U8058 (N_8058,N_7513,N_7839);
or U8059 (N_8059,N_7706,N_6848);
and U8060 (N_8060,N_7892,N_6034);
or U8061 (N_8061,N_6131,N_7648);
nor U8062 (N_8062,N_6151,N_6541);
nor U8063 (N_8063,N_7178,N_6969);
nand U8064 (N_8064,N_7058,N_6579);
nor U8065 (N_8065,N_6211,N_6515);
xor U8066 (N_8066,N_7433,N_7296);
nand U8067 (N_8067,N_6477,N_7873);
nor U8068 (N_8068,N_7442,N_7850);
nor U8069 (N_8069,N_7196,N_7907);
or U8070 (N_8070,N_6549,N_6581);
xor U8071 (N_8071,N_7972,N_6010);
and U8072 (N_8072,N_6126,N_7414);
nand U8073 (N_8073,N_7215,N_7820);
nor U8074 (N_8074,N_6007,N_7385);
nor U8075 (N_8075,N_7861,N_6352);
xnor U8076 (N_8076,N_6302,N_7659);
and U8077 (N_8077,N_6079,N_7517);
and U8078 (N_8078,N_7376,N_6116);
or U8079 (N_8079,N_7957,N_7990);
or U8080 (N_8080,N_7720,N_7832);
xnor U8081 (N_8081,N_7224,N_7488);
nor U8082 (N_8082,N_7452,N_6074);
or U8083 (N_8083,N_7699,N_6391);
nor U8084 (N_8084,N_6510,N_6786);
nand U8085 (N_8085,N_7947,N_7151);
and U8086 (N_8086,N_6021,N_7204);
nand U8087 (N_8087,N_6308,N_6744);
nor U8088 (N_8088,N_7010,N_6585);
nor U8089 (N_8089,N_6008,N_7961);
nor U8090 (N_8090,N_7944,N_6412);
nor U8091 (N_8091,N_7458,N_6626);
nand U8092 (N_8092,N_7743,N_7362);
nor U8093 (N_8093,N_6285,N_6914);
and U8094 (N_8094,N_6303,N_6649);
nand U8095 (N_8095,N_6845,N_7999);
and U8096 (N_8096,N_6413,N_7904);
or U8097 (N_8097,N_7905,N_7523);
nor U8098 (N_8098,N_6053,N_7881);
and U8099 (N_8099,N_7232,N_7213);
and U8100 (N_8100,N_7459,N_6849);
nor U8101 (N_8101,N_7986,N_7120);
xnor U8102 (N_8102,N_7390,N_6306);
and U8103 (N_8103,N_7135,N_7847);
nand U8104 (N_8104,N_6173,N_7794);
nor U8105 (N_8105,N_7610,N_6208);
nand U8106 (N_8106,N_7487,N_7138);
nor U8107 (N_8107,N_6994,N_7602);
or U8108 (N_8108,N_7419,N_7811);
and U8109 (N_8109,N_6268,N_7948);
nor U8110 (N_8110,N_7695,N_7034);
or U8111 (N_8111,N_6437,N_7669);
nand U8112 (N_8112,N_7083,N_7966);
nand U8113 (N_8113,N_6354,N_7650);
or U8114 (N_8114,N_6548,N_7474);
nor U8115 (N_8115,N_7318,N_7088);
nor U8116 (N_8116,N_7073,N_7370);
nand U8117 (N_8117,N_6617,N_7462);
nor U8118 (N_8118,N_7457,N_7760);
and U8119 (N_8119,N_6811,N_6472);
or U8120 (N_8120,N_6702,N_7189);
nor U8121 (N_8121,N_7516,N_7177);
or U8122 (N_8122,N_7327,N_7927);
and U8123 (N_8123,N_7603,N_7826);
and U8124 (N_8124,N_6334,N_7793);
nand U8125 (N_8125,N_6644,N_6659);
and U8126 (N_8126,N_6386,N_7226);
nor U8127 (N_8127,N_6060,N_7554);
and U8128 (N_8128,N_7778,N_7212);
nor U8129 (N_8129,N_7955,N_7359);
or U8130 (N_8130,N_7566,N_6410);
nand U8131 (N_8131,N_6538,N_6424);
nor U8132 (N_8132,N_6368,N_7038);
nor U8133 (N_8133,N_6573,N_7392);
nand U8134 (N_8134,N_7476,N_7284);
or U8135 (N_8135,N_6991,N_7356);
or U8136 (N_8136,N_7511,N_7230);
and U8137 (N_8137,N_7057,N_7797);
nor U8138 (N_8138,N_7423,N_7443);
nor U8139 (N_8139,N_7345,N_7260);
nor U8140 (N_8140,N_6342,N_7343);
or U8141 (N_8141,N_7619,N_7792);
and U8142 (N_8142,N_6785,N_7191);
nor U8143 (N_8143,N_7586,N_6557);
nor U8144 (N_8144,N_7757,N_7971);
nand U8145 (N_8145,N_7024,N_7882);
nand U8146 (N_8146,N_7441,N_6887);
nor U8147 (N_8147,N_6653,N_7363);
nand U8148 (N_8148,N_7465,N_6943);
and U8149 (N_8149,N_7075,N_7079);
or U8150 (N_8150,N_6293,N_6678);
nor U8151 (N_8151,N_6528,N_6789);
nand U8152 (N_8152,N_6743,N_6932);
nand U8153 (N_8153,N_6719,N_7835);
xor U8154 (N_8154,N_7862,N_7161);
or U8155 (N_8155,N_7871,N_6987);
nand U8156 (N_8156,N_6756,N_6803);
nor U8157 (N_8157,N_7365,N_6267);
or U8158 (N_8158,N_7606,N_6457);
nor U8159 (N_8159,N_7908,N_7111);
nand U8160 (N_8160,N_7520,N_7308);
or U8161 (N_8161,N_7245,N_7581);
nand U8162 (N_8162,N_6487,N_6736);
nor U8163 (N_8163,N_6329,N_7097);
nand U8164 (N_8164,N_7371,N_6262);
or U8165 (N_8165,N_7682,N_6415);
nor U8166 (N_8166,N_7157,N_6018);
nand U8167 (N_8167,N_7461,N_7349);
nand U8168 (N_8168,N_7087,N_7507);
nor U8169 (N_8169,N_6809,N_7313);
or U8170 (N_8170,N_7742,N_6922);
nand U8171 (N_8171,N_6174,N_7615);
nand U8172 (N_8172,N_6858,N_6652);
nand U8173 (N_8173,N_6506,N_7558);
or U8174 (N_8174,N_6956,N_7833);
nor U8175 (N_8175,N_7089,N_6503);
and U8176 (N_8176,N_6613,N_6307);
nand U8177 (N_8177,N_6661,N_6075);
or U8178 (N_8178,N_7049,N_6150);
nor U8179 (N_8179,N_7796,N_6192);
nor U8180 (N_8180,N_6533,N_6323);
nor U8181 (N_8181,N_6411,N_7738);
nand U8182 (N_8182,N_7933,N_7454);
or U8183 (N_8183,N_6855,N_6818);
and U8184 (N_8184,N_7130,N_7121);
and U8185 (N_8185,N_6171,N_6599);
and U8186 (N_8186,N_6568,N_7019);
or U8187 (N_8187,N_6988,N_7802);
nand U8188 (N_8188,N_6026,N_6179);
xor U8189 (N_8189,N_6219,N_7596);
or U8190 (N_8190,N_6820,N_7272);
and U8191 (N_8191,N_6304,N_6901);
nor U8192 (N_8192,N_7062,N_6029);
and U8193 (N_8193,N_7726,N_6928);
nor U8194 (N_8194,N_7160,N_6561);
or U8195 (N_8195,N_6518,N_7621);
or U8196 (N_8196,N_7338,N_7749);
or U8197 (N_8197,N_6364,N_6388);
or U8198 (N_8198,N_7562,N_7968);
or U8199 (N_8199,N_6582,N_7424);
or U8200 (N_8200,N_6972,N_6850);
or U8201 (N_8201,N_7624,N_6658);
nor U8202 (N_8202,N_6783,N_6758);
and U8203 (N_8203,N_6938,N_6038);
and U8204 (N_8204,N_6181,N_7434);
nand U8205 (N_8205,N_7611,N_7219);
xor U8206 (N_8206,N_6833,N_6872);
nor U8207 (N_8207,N_7578,N_7573);
nor U8208 (N_8208,N_6746,N_6862);
and U8209 (N_8209,N_6926,N_6616);
nand U8210 (N_8210,N_7113,N_6063);
or U8211 (N_8211,N_6861,N_6350);
and U8212 (N_8212,N_6940,N_6618);
nor U8213 (N_8213,N_6936,N_7779);
nand U8214 (N_8214,N_7956,N_7096);
nand U8215 (N_8215,N_7818,N_7309);
nand U8216 (N_8216,N_7608,N_6888);
or U8217 (N_8217,N_7675,N_7436);
or U8218 (N_8218,N_6752,N_7837);
nand U8219 (N_8219,N_7731,N_7868);
and U8220 (N_8220,N_6832,N_6000);
or U8221 (N_8221,N_6904,N_7439);
and U8222 (N_8222,N_7262,N_6546);
or U8223 (N_8223,N_7282,N_7694);
or U8224 (N_8224,N_7233,N_7970);
nor U8225 (N_8225,N_6570,N_6870);
nor U8226 (N_8226,N_6500,N_6356);
nor U8227 (N_8227,N_6997,N_7569);
and U8228 (N_8228,N_7590,N_6300);
and U8229 (N_8229,N_6036,N_7665);
and U8230 (N_8230,N_6019,N_6452);
nor U8231 (N_8231,N_7567,N_7598);
nor U8232 (N_8232,N_7547,N_6403);
nand U8233 (N_8233,N_7919,N_6269);
nand U8234 (N_8234,N_6565,N_7754);
nor U8235 (N_8235,N_7004,N_6360);
or U8236 (N_8236,N_6960,N_7382);
or U8237 (N_8237,N_7774,N_7216);
or U8238 (N_8238,N_7510,N_7077);
or U8239 (N_8239,N_7464,N_6012);
or U8240 (N_8240,N_6204,N_7982);
xnor U8241 (N_8241,N_6892,N_6989);
nor U8242 (N_8242,N_7662,N_6483);
or U8243 (N_8243,N_6276,N_6338);
nand U8244 (N_8244,N_6148,N_6876);
nor U8245 (N_8245,N_6602,N_6340);
nor U8246 (N_8246,N_7071,N_7386);
nor U8247 (N_8247,N_7391,N_7217);
nand U8248 (N_8248,N_7628,N_6020);
nor U8249 (N_8249,N_7543,N_7003);
or U8250 (N_8250,N_6138,N_6247);
and U8251 (N_8251,N_7552,N_6735);
nand U8252 (N_8252,N_6713,N_6840);
and U8253 (N_8253,N_7887,N_6183);
and U8254 (N_8254,N_6980,N_7722);
nor U8255 (N_8255,N_6374,N_6473);
and U8256 (N_8256,N_6062,N_7770);
or U8257 (N_8257,N_7225,N_7623);
nor U8258 (N_8258,N_6898,N_6884);
nor U8259 (N_8259,N_6981,N_7381);
nand U8260 (N_8260,N_7495,N_7925);
or U8261 (N_8261,N_6023,N_7500);
nor U8262 (N_8262,N_7588,N_7035);
or U8263 (N_8263,N_6953,N_6175);
or U8264 (N_8264,N_6115,N_7574);
or U8265 (N_8265,N_6331,N_6398);
nand U8266 (N_8266,N_6772,N_6596);
nand U8267 (N_8267,N_7239,N_7884);
or U8268 (N_8268,N_7983,N_6463);
and U8269 (N_8269,N_6679,N_6145);
or U8270 (N_8270,N_6512,N_6918);
or U8271 (N_8271,N_6777,N_7253);
nor U8272 (N_8272,N_6432,N_7045);
and U8273 (N_8273,N_7198,N_6740);
nand U8274 (N_8274,N_6113,N_7555);
or U8275 (N_8275,N_7660,N_7490);
nand U8276 (N_8276,N_7438,N_6475);
nand U8277 (N_8277,N_7310,N_6081);
or U8278 (N_8278,N_6249,N_6425);
nand U8279 (N_8279,N_7480,N_6706);
nor U8280 (N_8280,N_6650,N_7112);
nand U8281 (N_8281,N_6742,N_7145);
and U8282 (N_8282,N_6843,N_6134);
and U8283 (N_8283,N_6830,N_7549);
and U8284 (N_8284,N_6695,N_7806);
and U8285 (N_8285,N_6726,N_7782);
nand U8286 (N_8286,N_7859,N_7022);
or U8287 (N_8287,N_6770,N_6636);
or U8288 (N_8288,N_7952,N_7124);
nor U8289 (N_8289,N_7410,N_7689);
nor U8290 (N_8290,N_7658,N_6622);
and U8291 (N_8291,N_7162,N_6601);
and U8292 (N_8292,N_7333,N_6737);
or U8293 (N_8293,N_6235,N_6054);
nand U8294 (N_8294,N_6258,N_6088);
and U8295 (N_8295,N_7348,N_7341);
nor U8296 (N_8296,N_6687,N_7821);
or U8297 (N_8297,N_7938,N_7918);
or U8298 (N_8298,N_6385,N_7888);
or U8299 (N_8299,N_7194,N_7211);
nand U8300 (N_8300,N_6144,N_6284);
nand U8301 (N_8301,N_6003,N_6125);
or U8302 (N_8302,N_6031,N_7323);
nand U8303 (N_8303,N_6189,N_7234);
and U8304 (N_8304,N_6524,N_7188);
nor U8305 (N_8305,N_6837,N_6540);
and U8306 (N_8306,N_7877,N_7147);
or U8307 (N_8307,N_7231,N_6716);
and U8308 (N_8308,N_6731,N_6796);
or U8309 (N_8309,N_7290,N_7780);
and U8310 (N_8310,N_6996,N_6478);
nand U8311 (N_8311,N_6640,N_7316);
xnor U8312 (N_8312,N_6279,N_7240);
nand U8313 (N_8313,N_7631,N_6387);
nor U8314 (N_8314,N_6883,N_6362);
or U8315 (N_8315,N_6908,N_6239);
and U8316 (N_8316,N_7960,N_6660);
or U8317 (N_8317,N_6455,N_7561);
nand U8318 (N_8318,N_7958,N_7677);
nand U8319 (N_8319,N_6574,N_7548);
nand U8320 (N_8320,N_7741,N_7367);
and U8321 (N_8321,N_7784,N_6159);
or U8322 (N_8322,N_6314,N_7306);
nand U8323 (N_8323,N_6025,N_7613);
and U8324 (N_8324,N_7330,N_7479);
or U8325 (N_8325,N_6376,N_7238);
nand U8326 (N_8326,N_6343,N_6900);
or U8327 (N_8327,N_6619,N_6212);
and U8328 (N_8328,N_6289,N_6717);
or U8329 (N_8329,N_7664,N_7612);
and U8330 (N_8330,N_7814,N_6361);
and U8331 (N_8331,N_7002,N_6164);
and U8332 (N_8332,N_7775,N_6621);
and U8333 (N_8333,N_7257,N_7989);
nor U8334 (N_8334,N_6322,N_7118);
nor U8335 (N_8335,N_7954,N_6408);
nand U8336 (N_8336,N_6748,N_7626);
xor U8337 (N_8337,N_6022,N_7406);
and U8338 (N_8338,N_7830,N_7709);
and U8339 (N_8339,N_7336,N_6149);
nor U8340 (N_8340,N_6166,N_6807);
nand U8341 (N_8341,N_6474,N_6236);
and U8342 (N_8342,N_7127,N_7758);
and U8343 (N_8343,N_7750,N_6345);
nand U8344 (N_8344,N_7844,N_7788);
nor U8345 (N_8345,N_6064,N_6897);
nand U8346 (N_8346,N_7636,N_7048);
nand U8347 (N_8347,N_6851,N_7146);
or U8348 (N_8348,N_7752,N_7872);
nor U8349 (N_8349,N_7714,N_6798);
nand U8350 (N_8350,N_7672,N_6782);
xnor U8351 (N_8351,N_6152,N_6363);
nor U8352 (N_8352,N_7154,N_6979);
and U8353 (N_8353,N_6709,N_7354);
nor U8354 (N_8354,N_7223,N_7489);
nor U8355 (N_8355,N_7502,N_7378);
nor U8356 (N_8356,N_6040,N_6684);
nor U8357 (N_8357,N_6576,N_7683);
and U8358 (N_8358,N_7771,N_6383);
nor U8359 (N_8359,N_6418,N_7395);
nand U8360 (N_8360,N_7969,N_7831);
nor U8361 (N_8361,N_6977,N_7455);
and U8362 (N_8362,N_7915,N_7587);
and U8363 (N_8363,N_6930,N_6465);
nand U8364 (N_8364,N_7736,N_6015);
nor U8365 (N_8365,N_6569,N_7273);
nand U8366 (N_8366,N_6799,N_6421);
xnor U8367 (N_8367,N_7640,N_7870);
nand U8368 (N_8368,N_6227,N_6700);
nor U8369 (N_8369,N_6032,N_7319);
or U8370 (N_8370,N_7377,N_7759);
nor U8371 (N_8371,N_7114,N_6456);
nand U8372 (N_8372,N_6186,N_7360);
or U8373 (N_8373,N_6946,N_7165);
or U8374 (N_8374,N_7418,N_6093);
and U8375 (N_8375,N_6486,N_7182);
xor U8376 (N_8376,N_7117,N_7156);
nor U8377 (N_8377,N_6123,N_6630);
and U8378 (N_8378,N_6722,N_6016);
and U8379 (N_8379,N_7241,N_7804);
nor U8380 (N_8380,N_7595,N_7123);
and U8381 (N_8381,N_7498,N_7931);
or U8382 (N_8382,N_6825,N_7195);
or U8383 (N_8383,N_6241,N_6337);
nand U8384 (N_8384,N_6246,N_6112);
nor U8385 (N_8385,N_7705,N_7867);
nand U8386 (N_8386,N_7249,N_7857);
and U8387 (N_8387,N_7582,N_7874);
and U8388 (N_8388,N_7980,N_6532);
nand U8389 (N_8389,N_6627,N_7786);
and U8390 (N_8390,N_7374,N_7202);
nand U8391 (N_8391,N_6160,N_7258);
and U8392 (N_8392,N_6124,N_7148);
nor U8393 (N_8393,N_7460,N_6266);
nand U8394 (N_8394,N_6610,N_7158);
nand U8395 (N_8395,N_6780,N_7680);
nor U8396 (N_8396,N_7800,N_6543);
or U8397 (N_8397,N_6315,N_7505);
and U8398 (N_8398,N_6162,N_7846);
and U8399 (N_8399,N_7842,N_6683);
or U8400 (N_8400,N_6970,N_7690);
nand U8401 (N_8401,N_6583,N_6929);
nand U8402 (N_8402,N_7304,N_7641);
and U8403 (N_8403,N_7977,N_6729);
and U8404 (N_8404,N_6589,N_7651);
nand U8405 (N_8405,N_6194,N_6459);
nor U8406 (N_8406,N_7400,N_7655);
and U8407 (N_8407,N_7200,N_6982);
nor U8408 (N_8408,N_6451,N_7214);
and U8409 (N_8409,N_7589,N_6450);
or U8410 (N_8410,N_6600,N_7432);
nand U8411 (N_8411,N_7030,N_7951);
and U8412 (N_8412,N_7748,N_7286);
nand U8413 (N_8413,N_7404,N_6859);
nor U8414 (N_8414,N_6625,N_6829);
and U8415 (N_8415,N_7013,N_7509);
nor U8416 (N_8416,N_7428,N_6311);
nor U8417 (N_8417,N_7103,N_7407);
nand U8418 (N_8418,N_6947,N_7063);
and U8419 (N_8419,N_7576,N_7526);
nor U8420 (N_8420,N_6638,N_6339);
and U8421 (N_8421,N_7827,N_6142);
nor U8422 (N_8422,N_6407,N_6395);
or U8423 (N_8423,N_7484,N_7477);
nand U8424 (N_8424,N_6513,N_6933);
nor U8425 (N_8425,N_7838,N_6784);
or U8426 (N_8426,N_6215,N_7492);
and U8427 (N_8427,N_6349,N_6781);
nand U8428 (N_8428,N_6937,N_7700);
and U8429 (N_8429,N_6864,N_6494);
or U8430 (N_8430,N_7143,N_7777);
nand U8431 (N_8431,N_6787,N_6866);
or U8432 (N_8432,N_6577,N_7429);
nand U8433 (N_8433,N_7261,N_6757);
and U8434 (N_8434,N_6009,N_7551);
nand U8435 (N_8435,N_7537,N_6773);
nor U8436 (N_8436,N_7978,N_6401);
or U8437 (N_8437,N_6537,N_7183);
or U8438 (N_8438,N_7399,N_6373);
and U8439 (N_8439,N_6196,N_6252);
nand U8440 (N_8440,N_7252,N_7136);
nand U8441 (N_8441,N_7875,N_7497);
and U8442 (N_8442,N_7179,N_7854);
nand U8443 (N_8443,N_7236,N_7852);
or U8444 (N_8444,N_7383,N_6516);
nor U8445 (N_8445,N_6446,N_7607);
nand U8446 (N_8446,N_6823,N_6370);
or U8447 (N_8447,N_6955,N_7963);
nor U8448 (N_8448,N_7076,N_7991);
and U8449 (N_8449,N_7483,N_6492);
and U8450 (N_8450,N_6597,N_7995);
or U8451 (N_8451,N_6165,N_6119);
or U8452 (N_8452,N_6443,N_6428);
and U8453 (N_8453,N_7274,N_7373);
and U8454 (N_8454,N_6250,N_7294);
or U8455 (N_8455,N_6877,N_7855);
nand U8456 (N_8456,N_7066,N_7425);
nor U8457 (N_8457,N_7364,N_6718);
nand U8458 (N_8458,N_7440,N_6397);
nor U8459 (N_8459,N_6667,N_7845);
and U8460 (N_8460,N_6819,N_6052);
nor U8461 (N_8461,N_7012,N_7394);
or U8462 (N_8462,N_7453,N_6891);
or U8463 (N_8463,N_6995,N_6461);
and U8464 (N_8464,N_6962,N_6689);
nand U8465 (N_8465,N_6468,N_7992);
nor U8466 (N_8466,N_7131,N_7535);
or U8467 (N_8467,N_6035,N_7289);
nand U8468 (N_8468,N_7617,N_6091);
nand U8469 (N_8469,N_7643,N_7912);
and U8470 (N_8470,N_6067,N_7579);
nor U8471 (N_8471,N_6426,N_6263);
and U8472 (N_8472,N_7084,N_7227);
and U8473 (N_8473,N_6654,N_7803);
nand U8474 (N_8474,N_6882,N_6594);
nor U8475 (N_8475,N_7317,N_6312);
nand U8476 (N_8476,N_7637,N_7184);
or U8477 (N_8477,N_7017,N_6221);
and U8478 (N_8478,N_6328,N_6578);
and U8479 (N_8479,N_6086,N_6641);
or U8480 (N_8480,N_7889,N_6567);
and U8481 (N_8481,N_6704,N_6853);
nor U8482 (N_8482,N_7153,N_7295);
and U8483 (N_8483,N_6923,N_6673);
and U8484 (N_8484,N_7616,N_6471);
or U8485 (N_8485,N_7541,N_7530);
nand U8486 (N_8486,N_7920,N_6842);
and U8487 (N_8487,N_6121,N_7916);
nand U8488 (N_8488,N_6098,N_6815);
nor U8489 (N_8489,N_6732,N_7408);
nand U8490 (N_8490,N_6629,N_7974);
nor U8491 (N_8491,N_6677,N_7863);
nand U8492 (N_8492,N_6698,N_7524);
and U8493 (N_8493,N_7542,N_6598);
nor U8494 (N_8494,N_6986,N_6675);
or U8495 (N_8495,N_6156,N_7880);
and U8496 (N_8496,N_6643,N_6277);
xor U8497 (N_8497,N_7652,N_6645);
xnor U8498 (N_8498,N_6488,N_7203);
nand U8499 (N_8499,N_6335,N_7122);
nor U8500 (N_8500,N_7342,N_7550);
or U8501 (N_8501,N_7568,N_6489);
nand U8502 (N_8502,N_7755,N_7817);
nand U8503 (N_8503,N_6794,N_7531);
nor U8504 (N_8504,N_6027,N_6633);
nand U8505 (N_8505,N_6551,N_7246);
or U8506 (N_8506,N_6118,N_7767);
nand U8507 (N_8507,N_6595,N_6292);
and U8508 (N_8508,N_7649,N_6559);
or U8509 (N_8509,N_6915,N_7584);
nand U8510 (N_8510,N_6490,N_6298);
or U8511 (N_8511,N_7387,N_6222);
and U8512 (N_8512,N_6656,N_6493);
nor U8513 (N_8513,N_7059,N_7305);
nand U8514 (N_8514,N_6734,N_7597);
and U8515 (N_8515,N_6497,N_7557);
nor U8516 (N_8516,N_6393,N_6485);
and U8517 (N_8517,N_7287,N_7020);
nand U8518 (N_8518,N_7671,N_6801);
or U8519 (N_8519,N_7435,N_6371);
nand U8520 (N_8520,N_6632,N_7346);
or U8521 (N_8521,N_6536,N_6379);
nand U8522 (N_8522,N_6768,N_6542);
nand U8523 (N_8523,N_7288,N_6496);
nand U8524 (N_8524,N_6187,N_6664);
nand U8525 (N_8525,N_7785,N_7593);
nand U8526 (N_8526,N_7155,N_7924);
nand U8527 (N_8527,N_6685,N_7199);
and U8528 (N_8528,N_7600,N_7678);
or U8529 (N_8529,N_7929,N_7413);
or U8530 (N_8530,N_7251,N_7080);
or U8531 (N_8531,N_6320,N_7009);
and U8532 (N_8532,N_6727,N_7858);
and U8533 (N_8533,N_7941,N_6005);
and U8534 (N_8534,N_7292,N_7141);
nor U8535 (N_8535,N_7108,N_7673);
xor U8536 (N_8536,N_7315,N_6792);
or U8537 (N_8537,N_6006,N_6919);
nor U8538 (N_8538,N_7221,N_6094);
or U8539 (N_8539,N_6207,N_6101);
and U8540 (N_8540,N_6414,N_6836);
nor U8541 (N_8541,N_6526,N_6234);
nand U8542 (N_8542,N_7988,N_6624);
or U8543 (N_8543,N_7421,N_7475);
or U8544 (N_8544,N_6896,N_6871);
or U8545 (N_8545,N_6560,N_6048);
or U8546 (N_8546,N_6274,N_7248);
and U8547 (N_8547,N_6201,N_7824);
nand U8548 (N_8548,N_7622,N_6993);
or U8549 (N_8549,N_7033,N_6409);
nor U8550 (N_8550,N_6514,N_6233);
or U8551 (N_8551,N_6523,N_6476);
nor U8552 (N_8552,N_7119,N_6163);
nor U8553 (N_8553,N_6944,N_6984);
xor U8554 (N_8554,N_7086,N_7560);
nand U8555 (N_8555,N_6655,N_7815);
nand U8556 (N_8556,N_6612,N_6971);
or U8557 (N_8557,N_7405,N_6230);
and U8558 (N_8558,N_7379,N_6216);
and U8559 (N_8559,N_6253,N_6066);
or U8560 (N_8560,N_6287,N_7044);
nor U8561 (N_8561,N_6692,N_7069);
nor U8562 (N_8562,N_6672,N_6776);
and U8563 (N_8563,N_7891,N_7326);
nand U8564 (N_8564,N_7007,N_7668);
nand U8565 (N_8565,N_6033,N_6275);
or U8566 (N_8566,N_6921,N_6085);
and U8567 (N_8567,N_7322,N_6244);
and U8568 (N_8568,N_6665,N_6501);
nand U8569 (N_8569,N_7269,N_6348);
nand U8570 (N_8570,N_6703,N_6055);
nand U8571 (N_8571,N_6255,N_6902);
or U8572 (N_8572,N_6102,N_6071);
and U8573 (N_8573,N_6299,N_6347);
and U8574 (N_8574,N_7099,N_6080);
nor U8575 (N_8575,N_6069,N_7300);
and U8576 (N_8576,N_6440,N_6992);
nand U8577 (N_8577,N_7396,N_7040);
nand U8578 (N_8578,N_6566,N_7192);
or U8579 (N_8579,N_7808,N_6751);
and U8580 (N_8580,N_7485,N_7564);
or U8581 (N_8581,N_6562,N_6434);
nor U8582 (N_8582,N_6449,N_6813);
nand U8583 (N_8583,N_7350,N_6050);
nor U8584 (N_8584,N_6620,N_6205);
or U8585 (N_8585,N_6694,N_6998);
or U8586 (N_8586,N_6931,N_7430);
xnor U8587 (N_8587,N_6881,N_6464);
nor U8588 (N_8588,N_6389,N_7353);
or U8589 (N_8589,N_7368,N_7412);
and U8590 (N_8590,N_6606,N_7397);
and U8591 (N_8591,N_7437,N_6857);
nand U8592 (N_8592,N_7109,N_6445);
nand U8593 (N_8593,N_7897,N_6591);
and U8594 (N_8594,N_6935,N_6875);
nor U8595 (N_8595,N_7899,N_7137);
or U8596 (N_8596,N_7638,N_6554);
nand U8597 (N_8597,N_7152,N_7021);
and U8598 (N_8598,N_7692,N_7703);
nand U8599 (N_8599,N_6073,N_6745);
nor U8600 (N_8600,N_7572,N_6251);
nand U8601 (N_8601,N_6865,N_6976);
nand U8602 (N_8602,N_6531,N_7491);
and U8603 (N_8603,N_6436,N_6178);
nor U8604 (N_8604,N_7280,N_6905);
nand U8605 (N_8605,N_6957,N_7032);
nor U8606 (N_8606,N_7816,N_7653);
nor U8607 (N_8607,N_6002,N_6755);
or U8608 (N_8608,N_7008,N_6087);
and U8609 (N_8609,N_7591,N_6575);
nor U8610 (N_8610,N_7945,N_7472);
or U8611 (N_8611,N_7388,N_6635);
nor U8612 (N_8612,N_6648,N_7900);
or U8613 (N_8613,N_6140,N_6394);
nand U8614 (N_8614,N_6961,N_6828);
nand U8615 (N_8615,N_6273,N_7139);
nor U8616 (N_8616,N_6310,N_7501);
and U8617 (N_8617,N_6402,N_6963);
and U8618 (N_8618,N_7674,N_6242);
or U8619 (N_8619,N_7559,N_6834);
and U8620 (N_8620,N_6959,N_7061);
nand U8621 (N_8621,N_7834,N_6231);
nand U8622 (N_8622,N_6671,N_7250);
and U8623 (N_8623,N_7783,N_7060);
nor U8624 (N_8624,N_7923,N_7267);
xnor U8625 (N_8625,N_6747,N_6290);
nand U8626 (N_8626,N_7268,N_7594);
xor U8627 (N_8627,N_6707,N_6004);
nor U8628 (N_8628,N_7670,N_6824);
nor U8629 (N_8629,N_6441,N_6769);
or U8630 (N_8630,N_6103,N_6321);
and U8631 (N_8631,N_6774,N_6874);
xor U8632 (N_8632,N_7657,N_7027);
nand U8633 (N_8633,N_6642,N_7206);
nand U8634 (N_8634,N_6941,N_7344);
and U8635 (N_8635,N_7055,N_6344);
and U8636 (N_8636,N_7218,N_6161);
xor U8637 (N_8637,N_7840,N_6948);
nor U8638 (N_8638,N_7744,N_6739);
or U8639 (N_8639,N_7661,N_7647);
nor U8640 (N_8640,N_6454,N_6521);
nor U8641 (N_8641,N_7463,N_7876);
nor U8642 (N_8642,N_6065,N_6697);
or U8643 (N_8643,N_6762,N_6197);
or U8644 (N_8644,N_6564,N_6039);
nor U8645 (N_8645,N_6708,N_7256);
xnor U8646 (N_8646,N_7243,N_6479);
or U8647 (N_8647,N_7747,N_6975);
nor U8648 (N_8648,N_6967,N_6056);
nor U8649 (N_8649,N_7140,N_6157);
and U8650 (N_8650,N_7810,N_7903);
nand U8651 (N_8651,N_6199,N_6592);
or U8652 (N_8652,N_6517,N_6417);
or U8653 (N_8653,N_7276,N_7018);
and U8654 (N_8654,N_6688,N_6631);
and U8655 (N_8655,N_6917,N_6358);
or U8656 (N_8656,N_6505,N_7174);
and U8657 (N_8657,N_6804,N_7962);
nor U8658 (N_8658,N_6580,N_6324);
nand U8659 (N_8659,N_6553,N_6508);
nand U8660 (N_8660,N_7633,N_7599);
and U8661 (N_8661,N_6042,N_6111);
or U8662 (N_8662,N_6313,N_6095);
nand U8663 (N_8663,N_6447,N_7540);
nor U8664 (N_8664,N_6202,N_7693);
nor U8665 (N_8665,N_6608,N_6346);
or U8666 (N_8666,N_6525,N_6623);
nand U8667 (N_8667,N_6639,N_6381);
nand U8668 (N_8668,N_7822,N_7922);
nand U8669 (N_8669,N_6046,N_7210);
nand U8670 (N_8670,N_6044,N_7133);
or U8671 (N_8671,N_7102,N_6139);
nor U8672 (N_8672,N_6260,N_7666);
or U8673 (N_8673,N_7914,N_6330);
or U8674 (N_8674,N_6122,N_7166);
or U8675 (N_8675,N_6952,N_6001);
and U8676 (N_8676,N_6458,N_7570);
or U8677 (N_8677,N_7745,N_6097);
or U8678 (N_8678,N_7893,N_6110);
or U8679 (N_8679,N_6147,N_7790);
and U8680 (N_8680,N_6435,N_6507);
nand U8681 (N_8681,N_6106,N_7696);
or U8682 (N_8682,N_7533,N_6498);
nand U8683 (N_8683,N_6188,N_7514);
nand U8684 (N_8684,N_7515,N_6404);
or U8685 (N_8685,N_6068,N_6484);
nand U8686 (N_8686,N_7470,N_7823);
nor U8687 (N_8687,N_7358,N_7037);
and U8688 (N_8688,N_6699,N_7934);
nor U8689 (N_8689,N_6682,N_6826);
nor U8690 (N_8690,N_7522,N_7761);
and U8691 (N_8691,N_6844,N_7228);
or U8692 (N_8692,N_6558,N_7444);
nand U8693 (N_8693,N_7527,N_6305);
nand U8694 (N_8694,N_7482,N_7366);
and U8695 (N_8695,N_6927,N_6369);
or U8696 (N_8696,N_6462,N_6535);
or U8697 (N_8697,N_6604,N_6827);
nand U8698 (N_8698,N_6127,N_6228);
nor U8699 (N_8699,N_7639,N_6916);
nor U8700 (N_8700,N_6572,N_6332);
nor U8701 (N_8701,N_6058,N_6805);
nor U8702 (N_8702,N_7627,N_6808);
or U8703 (N_8703,N_7185,N_6420);
or U8704 (N_8704,N_6676,N_7635);
or U8705 (N_8705,N_7813,N_7041);
or U8706 (N_8706,N_6817,N_6037);
or U8707 (N_8707,N_7285,N_6117);
or U8708 (N_8708,N_6847,N_7329);
and U8709 (N_8709,N_7115,N_7930);
nand U8710 (N_8710,N_6177,N_6092);
nand U8711 (N_8711,N_6950,N_6198);
nand U8712 (N_8712,N_6527,N_7539);
nand U8713 (N_8713,N_7176,N_7718);
nor U8714 (N_8714,N_6763,N_7255);
nand U8715 (N_8715,N_7031,N_7725);
or U8716 (N_8716,N_7679,N_7291);
and U8717 (N_8717,N_6693,N_6705);
nand U8718 (N_8718,N_7528,N_6681);
nor U8719 (N_8719,N_6353,N_6014);
or U8720 (N_8720,N_7301,N_7791);
nor U8721 (N_8721,N_7091,N_7170);
or U8722 (N_8722,N_7688,N_7132);
xnor U8723 (N_8723,N_6759,N_7687);
or U8724 (N_8724,N_6835,N_7265);
or U8725 (N_8725,N_6378,N_7719);
nand U8726 (N_8726,N_6605,N_6480);
and U8727 (N_8727,N_6790,N_6136);
nor U8728 (N_8728,N_7716,N_6964);
nor U8729 (N_8729,N_7751,N_6544);
nor U8730 (N_8730,N_6511,N_7565);
and U8731 (N_8731,N_6089,N_6185);
and U8732 (N_8732,N_7996,N_7028);
nor U8733 (N_8733,N_7529,N_7577);
nor U8734 (N_8734,N_7283,N_7768);
or U8735 (N_8735,N_6448,N_7043);
nor U8736 (N_8736,N_7860,N_6224);
xor U8737 (N_8737,N_7545,N_7054);
nor U8738 (N_8738,N_6587,N_6728);
or U8739 (N_8739,N_7765,N_7676);
nor U8740 (N_8740,N_6965,N_6470);
nor U8741 (N_8741,N_7415,N_7347);
or U8742 (N_8742,N_7324,N_7064);
and U8743 (N_8743,N_6220,N_6545);
nand U8744 (N_8744,N_6090,N_7926);
and U8745 (N_8745,N_6366,N_7618);
and U8746 (N_8746,N_7445,N_6105);
or U8747 (N_8747,N_7812,N_7101);
nand U8748 (N_8748,N_7580,N_6686);
and U8749 (N_8749,N_7592,N_6154);
nor U8750 (N_8750,N_7710,N_7167);
and U8751 (N_8751,N_6024,N_6482);
nor U8752 (N_8752,N_7015,N_7186);
nand U8753 (N_8753,N_7074,N_6288);
or U8754 (N_8754,N_7312,N_7355);
nor U8755 (N_8755,N_6810,N_7701);
nor U8756 (N_8756,N_6714,N_6223);
or U8757 (N_8757,N_6282,N_6614);
nand U8758 (N_8758,N_7518,N_7172);
or U8759 (N_8759,N_7422,N_6431);
and U8760 (N_8760,N_7403,N_7384);
and U8761 (N_8761,N_7646,N_6439);
nand U8762 (N_8762,N_6384,N_6168);
nand U8763 (N_8763,N_6852,N_6104);
or U8764 (N_8764,N_6509,N_6615);
and U8765 (N_8765,N_7856,N_7935);
nor U8766 (N_8766,N_7732,N_7050);
nor U8767 (N_8767,N_7081,N_6084);
and U8768 (N_8768,N_7467,N_7973);
xnor U8769 (N_8769,N_7244,N_6100);
and U8770 (N_8770,N_7764,N_7036);
or U8771 (N_8771,N_7070,N_6771);
nand U8772 (N_8772,N_7625,N_6272);
nand U8773 (N_8773,N_6990,N_7473);
or U8774 (N_8774,N_7895,N_7828);
nor U8775 (N_8775,N_7508,N_6611);
nand U8776 (N_8776,N_6467,N_7481);
nand U8777 (N_8777,N_7896,N_6556);
or U8778 (N_8778,N_6586,N_6720);
or U8779 (N_8779,N_6571,N_7142);
nand U8780 (N_8780,N_7042,N_6715);
and U8781 (N_8781,N_6051,N_6270);
nand U8782 (N_8782,N_7005,N_6359);
and U8783 (N_8783,N_6670,N_6382);
nand U8784 (N_8784,N_7546,N_6083);
nor U8785 (N_8785,N_7000,N_6120);
and U8786 (N_8786,N_6711,N_6172);
nand U8787 (N_8787,N_6107,N_7068);
nor U8788 (N_8788,N_6047,N_7209);
and U8789 (N_8789,N_6942,N_7266);
or U8790 (N_8790,N_6724,N_7993);
nand U8791 (N_8791,N_7708,N_7994);
nand U8792 (N_8792,N_6767,N_6301);
or U8793 (N_8793,N_7259,N_7866);
or U8794 (N_8794,N_7078,N_6043);
nand U8795 (N_8795,N_7735,N_7781);
nor U8796 (N_8796,N_6761,N_6663);
or U8797 (N_8797,N_6797,N_6460);
nand U8798 (N_8798,N_6669,N_6416);
nor U8799 (N_8799,N_6760,N_7702);
nor U8800 (N_8800,N_7512,N_7953);
nand U8801 (N_8801,N_6791,N_7987);
and U8802 (N_8802,N_7698,N_7825);
and U8803 (N_8803,N_7150,N_7684);
nor U8804 (N_8804,N_6355,N_6218);
nor U8805 (N_8805,N_7898,N_7632);
or U8806 (N_8806,N_7431,N_6869);
nor U8807 (N_8807,N_6939,N_7085);
and U8808 (N_8808,N_7985,N_6741);
nand U8809 (N_8809,N_7686,N_6070);
nor U8810 (N_8810,N_7116,N_7917);
and U8811 (N_8811,N_7082,N_7197);
nand U8812 (N_8812,N_6351,N_7801);
nor U8813 (N_8813,N_6466,N_6380);
and U8814 (N_8814,N_6788,N_6750);
or U8815 (N_8815,N_7795,N_7601);
nor U8816 (N_8816,N_6213,N_7449);
nor U8817 (N_8817,N_6076,N_6195);
nand U8818 (N_8818,N_7222,N_6427);
or U8819 (N_8819,N_6229,N_6133);
and U8820 (N_8820,N_7536,N_7964);
nor U8821 (N_8821,N_7940,N_6057);
nor U8822 (N_8822,N_7372,N_6232);
nand U8823 (N_8823,N_6550,N_6723);
and U8824 (N_8824,N_6297,N_7967);
nand U8825 (N_8825,N_6365,N_7939);
nor U8826 (N_8826,N_7879,N_6590);
nand U8827 (N_8827,N_7878,N_6628);
or U8828 (N_8828,N_7168,N_6237);
or U8829 (N_8829,N_7411,N_6795);
nor U8830 (N_8830,N_7339,N_6754);
nand U8831 (N_8831,N_6880,N_6710);
and U8832 (N_8832,N_7494,N_7129);
nand U8833 (N_8833,N_7728,N_6128);
nand U8834 (N_8834,N_7712,N_6913);
and U8835 (N_8835,N_7946,N_6072);
nand U8836 (N_8836,N_6153,N_6108);
and U8837 (N_8837,N_6907,N_7913);
and U8838 (N_8838,N_6028,N_7053);
or U8839 (N_8839,N_6375,N_6372);
xor U8840 (N_8840,N_7724,N_6911);
and U8841 (N_8841,N_6593,N_6190);
nor U8842 (N_8842,N_7890,N_7740);
or U8843 (N_8843,N_6563,N_6910);
or U8844 (N_8844,N_7984,N_6924);
nor U8845 (N_8845,N_7380,N_6584);
nor U8846 (N_8846,N_7375,N_7468);
or U8847 (N_8847,N_7159,N_7789);
and U8848 (N_8848,N_7681,N_7864);
and U8849 (N_8849,N_7047,N_7807);
nor U8850 (N_8850,N_6030,N_7092);
or U8851 (N_8851,N_6469,N_7328);
and U8852 (N_8852,N_7630,N_6281);
or U8853 (N_8853,N_7039,N_6668);
or U8854 (N_8854,N_7427,N_6733);
nand U8855 (N_8855,N_7451,N_6721);
or U8856 (N_8856,N_6011,N_7901);
nand U8857 (N_8857,N_7729,N_6390);
and U8858 (N_8858,N_7763,N_6265);
nand U8859 (N_8859,N_6812,N_7331);
and U8860 (N_8860,N_6906,N_6099);
nor U8861 (N_8861,N_6400,N_6433);
nor U8862 (N_8862,N_6779,N_7340);
and U8863 (N_8863,N_7849,N_7503);
or U8864 (N_8864,N_6903,N_6945);
or U8865 (N_8865,N_6130,N_6890);
nor U8866 (N_8866,N_6143,N_6912);
and U8867 (N_8867,N_7656,N_7398);
nor U8868 (N_8868,N_7220,N_7389);
nand U8869 (N_8869,N_6609,N_6886);
and U8870 (N_8870,N_7169,N_6367);
and U8871 (N_8871,N_7357,N_6077);
or U8872 (N_8872,N_7667,N_7107);
or U8873 (N_8873,N_6176,N_7620);
nor U8874 (N_8874,N_6206,N_7352);
or U8875 (N_8875,N_6978,N_7932);
or U8876 (N_8876,N_6822,N_6766);
or U8877 (N_8877,N_7909,N_7819);
nor U8878 (N_8878,N_6283,N_6657);
or U8879 (N_8879,N_6491,N_7762);
or U8880 (N_8880,N_6603,N_7943);
nor U8881 (N_8881,N_7271,N_7707);
and U8882 (N_8882,N_7311,N_6934);
nor U8883 (N_8883,N_7869,N_6806);
and U8884 (N_8884,N_7208,N_6245);
nand U8885 (N_8885,N_6712,N_6278);
and U8886 (N_8886,N_7975,N_7685);
and U8887 (N_8887,N_7270,N_6481);
nor U8888 (N_8888,N_6442,N_6816);
nor U8889 (N_8889,N_7851,N_6839);
or U8890 (N_8890,N_7979,N_7727);
nand U8891 (N_8891,N_6419,N_6200);
or U8892 (N_8892,N_6256,N_7229);
and U8893 (N_8893,N_7538,N_6854);
and U8894 (N_8894,N_7242,N_6775);
nor U8895 (N_8895,N_6899,N_7769);
and U8896 (N_8896,N_6749,N_6257);
and U8897 (N_8897,N_6909,N_7556);
or U8898 (N_8898,N_7998,N_6180);
nor U8899 (N_8899,N_6863,N_7949);
and U8900 (N_8900,N_7734,N_7281);
nand U8901 (N_8901,N_6879,N_7809);
nand U8902 (N_8902,N_7072,N_7634);
nor U8903 (N_8903,N_6588,N_7936);
or U8904 (N_8904,N_7805,N_7605);
or U8905 (N_8905,N_6968,N_7885);
nor U8906 (N_8906,N_7644,N_7163);
or U8907 (N_8907,N_7697,N_7715);
nor U8908 (N_8908,N_7297,N_7095);
or U8909 (N_8909,N_7125,N_7447);
and U8910 (N_8910,N_6146,N_7469);
or U8911 (N_8911,N_7937,N_7902);
nor U8912 (N_8912,N_6878,N_6607);
nor U8913 (N_8913,N_7521,N_6499);
nor U8914 (N_8914,N_7175,N_6325);
nand U8915 (N_8915,N_7279,N_6954);
nor U8916 (N_8916,N_6974,N_6309);
and U8917 (N_8917,N_6357,N_6753);
nand U8918 (N_8918,N_6264,N_6958);
and U8919 (N_8919,N_7886,N_7325);
and U8920 (N_8920,N_6392,N_6765);
or U8921 (N_8921,N_7393,N_6701);
nand U8922 (N_8922,N_6240,N_7190);
nor U8923 (N_8923,N_6730,N_7563);
and U8924 (N_8924,N_7056,N_6158);
nand U8925 (N_8925,N_7051,N_7553);
or U8926 (N_8926,N_6831,N_6651);
nor U8927 (N_8927,N_7187,N_7237);
or U8928 (N_8928,N_7928,N_7504);
nor U8929 (N_8929,N_6182,N_7614);
and U8930 (N_8930,N_7609,N_6226);
or U8931 (N_8931,N_7417,N_7787);
and U8932 (N_8932,N_7025,N_6406);
nor U8933 (N_8933,N_6017,N_6547);
and U8934 (N_8934,N_7110,N_7128);
nor U8935 (N_8935,N_7094,N_7853);
xnor U8936 (N_8936,N_7207,N_6049);
and U8937 (N_8937,N_6495,N_7843);
nor U8938 (N_8938,N_7420,N_7263);
nand U8939 (N_8939,N_7307,N_6821);
or U8940 (N_8940,N_6341,N_7894);
and U8941 (N_8941,N_7534,N_7426);
and U8942 (N_8942,N_6243,N_7753);
or U8943 (N_8943,N_7733,N_7799);
nor U8944 (N_8944,N_6637,N_7335);
nand U8945 (N_8945,N_7997,N_7332);
xor U8946 (N_8946,N_7519,N_7798);
nor U8947 (N_8947,N_6646,N_6552);
or U8948 (N_8948,N_6502,N_6920);
nand U8949 (N_8949,N_6405,N_6893);
or U8950 (N_8950,N_7772,N_7201);
or U8951 (N_8951,N_7106,N_7173);
and U8952 (N_8952,N_6294,N_6814);
nand U8953 (N_8953,N_7093,N_7401);
nor U8954 (N_8954,N_6059,N_7836);
nor U8955 (N_8955,N_7645,N_7950);
and U8956 (N_8956,N_7180,N_6453);
nor U8957 (N_8957,N_7865,N_7654);
or U8958 (N_8958,N_6261,N_7575);
nand U8959 (N_8959,N_7361,N_6210);
or U8960 (N_8960,N_7193,N_6013);
nand U8961 (N_8961,N_7171,N_7739);
nor U8962 (N_8962,N_6520,N_6860);
or U8963 (N_8963,N_7571,N_6674);
nor U8964 (N_8964,N_6691,N_6423);
nor U8965 (N_8965,N_6522,N_6114);
and U8966 (N_8966,N_6966,N_6061);
or U8967 (N_8967,N_6973,N_7164);
nand U8968 (N_8968,N_7254,N_7981);
or U8969 (N_8969,N_6336,N_7247);
nand U8970 (N_8970,N_6319,N_7746);
nand U8971 (N_8971,N_7711,N_7029);
and U8972 (N_8972,N_6326,N_7448);
and U8973 (N_8973,N_7829,N_6109);
nor U8974 (N_8974,N_6725,N_6838);
and U8975 (N_8975,N_6295,N_7014);
nand U8976 (N_8976,N_6191,N_6634);
nor U8977 (N_8977,N_7026,N_6738);
nor U8978 (N_8978,N_7303,N_6296);
nand U8979 (N_8979,N_7525,N_7965);
or U8980 (N_8980,N_7100,N_7883);
nor U8981 (N_8981,N_6078,N_7302);
nor U8982 (N_8982,N_7450,N_6999);
nor U8983 (N_8983,N_7205,N_6690);
and U8984 (N_8984,N_7713,N_7105);
xnor U8985 (N_8985,N_6155,N_7456);
or U8986 (N_8986,N_6429,N_6399);
nor U8987 (N_8987,N_6534,N_7006);
nor U8988 (N_8988,N_6867,N_7730);
nand U8989 (N_8989,N_6193,N_7126);
nor U8990 (N_8990,N_6778,N_6254);
nor U8991 (N_8991,N_7090,N_6396);
and U8992 (N_8992,N_6203,N_6444);
nand U8993 (N_8993,N_6764,N_6214);
nor U8994 (N_8994,N_7149,N_6286);
or U8995 (N_8995,N_6169,N_7976);
nand U8996 (N_8996,N_6666,N_6045);
nor U8997 (N_8997,N_6430,N_7766);
and U8998 (N_8998,N_6318,N_6949);
nand U8999 (N_8999,N_7011,N_6985);
nor U9000 (N_9000,N_6018,N_7604);
or U9001 (N_9001,N_7120,N_7225);
nand U9002 (N_9002,N_7054,N_7812);
nand U9003 (N_9003,N_6045,N_6143);
nand U9004 (N_9004,N_7032,N_7931);
nand U9005 (N_9005,N_7339,N_7864);
nand U9006 (N_9006,N_6609,N_7013);
or U9007 (N_9007,N_6680,N_6948);
nor U9008 (N_9008,N_6909,N_6457);
nor U9009 (N_9009,N_6480,N_7663);
nand U9010 (N_9010,N_7224,N_7034);
nor U9011 (N_9011,N_6963,N_7525);
nand U9012 (N_9012,N_7806,N_7690);
or U9013 (N_9013,N_6561,N_6871);
nor U9014 (N_9014,N_7561,N_6437);
nor U9015 (N_9015,N_7820,N_6117);
and U9016 (N_9016,N_6762,N_7660);
or U9017 (N_9017,N_6007,N_7277);
or U9018 (N_9018,N_7224,N_7768);
nand U9019 (N_9019,N_6333,N_6407);
and U9020 (N_9020,N_6721,N_6323);
or U9021 (N_9021,N_6370,N_6442);
nand U9022 (N_9022,N_6690,N_6553);
or U9023 (N_9023,N_6313,N_7269);
nor U9024 (N_9024,N_6428,N_6708);
xnor U9025 (N_9025,N_7910,N_7942);
or U9026 (N_9026,N_7956,N_6005);
xor U9027 (N_9027,N_6348,N_7593);
nand U9028 (N_9028,N_6270,N_6866);
nand U9029 (N_9029,N_7813,N_7546);
and U9030 (N_9030,N_6368,N_6830);
or U9031 (N_9031,N_7302,N_6483);
or U9032 (N_9032,N_7203,N_7171);
nand U9033 (N_9033,N_6864,N_7077);
nand U9034 (N_9034,N_7705,N_7039);
and U9035 (N_9035,N_7225,N_6909);
and U9036 (N_9036,N_6951,N_7844);
or U9037 (N_9037,N_7003,N_6600);
or U9038 (N_9038,N_7670,N_7268);
or U9039 (N_9039,N_6105,N_6791);
and U9040 (N_9040,N_7439,N_6754);
and U9041 (N_9041,N_6120,N_6854);
nor U9042 (N_9042,N_7253,N_7376);
and U9043 (N_9043,N_6055,N_7535);
nand U9044 (N_9044,N_6266,N_7138);
nor U9045 (N_9045,N_6609,N_6037);
and U9046 (N_9046,N_6171,N_7444);
and U9047 (N_9047,N_6521,N_6958);
nand U9048 (N_9048,N_6042,N_6092);
nand U9049 (N_9049,N_7097,N_6277);
and U9050 (N_9050,N_7664,N_6319);
and U9051 (N_9051,N_7741,N_6249);
and U9052 (N_9052,N_7953,N_6047);
nor U9053 (N_9053,N_6205,N_6616);
or U9054 (N_9054,N_7563,N_7254);
and U9055 (N_9055,N_7363,N_7844);
xor U9056 (N_9056,N_6127,N_7442);
and U9057 (N_9057,N_7483,N_6645);
and U9058 (N_9058,N_6894,N_7628);
nor U9059 (N_9059,N_7747,N_6267);
or U9060 (N_9060,N_7099,N_6996);
nand U9061 (N_9061,N_7184,N_7388);
and U9062 (N_9062,N_6724,N_7540);
nor U9063 (N_9063,N_7331,N_6472);
nor U9064 (N_9064,N_7302,N_6972);
and U9065 (N_9065,N_6697,N_7760);
or U9066 (N_9066,N_6206,N_6808);
or U9067 (N_9067,N_6886,N_6020);
or U9068 (N_9068,N_7707,N_7585);
nor U9069 (N_9069,N_7171,N_7720);
nor U9070 (N_9070,N_6049,N_6429);
nand U9071 (N_9071,N_7552,N_7309);
nand U9072 (N_9072,N_6415,N_6740);
or U9073 (N_9073,N_7164,N_6504);
nand U9074 (N_9074,N_7184,N_6913);
or U9075 (N_9075,N_6321,N_7449);
or U9076 (N_9076,N_6704,N_6385);
nor U9077 (N_9077,N_7790,N_7760);
or U9078 (N_9078,N_6865,N_6130);
and U9079 (N_9079,N_6459,N_7072);
nor U9080 (N_9080,N_7453,N_7119);
and U9081 (N_9081,N_7832,N_7366);
or U9082 (N_9082,N_6057,N_6468);
nor U9083 (N_9083,N_7857,N_7331);
nor U9084 (N_9084,N_6199,N_7578);
nor U9085 (N_9085,N_7175,N_7344);
nand U9086 (N_9086,N_7560,N_7655);
xor U9087 (N_9087,N_6409,N_6636);
or U9088 (N_9088,N_6441,N_6179);
nand U9089 (N_9089,N_6157,N_6160);
nand U9090 (N_9090,N_7820,N_7190);
or U9091 (N_9091,N_6943,N_6914);
and U9092 (N_9092,N_6773,N_6565);
nand U9093 (N_9093,N_6764,N_7786);
nor U9094 (N_9094,N_6771,N_7542);
or U9095 (N_9095,N_6994,N_7589);
nor U9096 (N_9096,N_7519,N_6032);
or U9097 (N_9097,N_6899,N_7952);
or U9098 (N_9098,N_7989,N_6248);
nand U9099 (N_9099,N_7800,N_6928);
or U9100 (N_9100,N_6588,N_7342);
nor U9101 (N_9101,N_6000,N_6211);
and U9102 (N_9102,N_7067,N_7282);
or U9103 (N_9103,N_7443,N_6358);
or U9104 (N_9104,N_6505,N_7022);
nand U9105 (N_9105,N_6430,N_7198);
and U9106 (N_9106,N_7179,N_6899);
or U9107 (N_9107,N_7350,N_6155);
and U9108 (N_9108,N_7702,N_6046);
nor U9109 (N_9109,N_6457,N_6491);
nor U9110 (N_9110,N_7256,N_6789);
or U9111 (N_9111,N_7326,N_7195);
or U9112 (N_9112,N_7374,N_7134);
and U9113 (N_9113,N_6004,N_7610);
or U9114 (N_9114,N_6025,N_7811);
and U9115 (N_9115,N_7374,N_7949);
nor U9116 (N_9116,N_6441,N_7078);
nand U9117 (N_9117,N_6883,N_6931);
nor U9118 (N_9118,N_6341,N_6071);
xnor U9119 (N_9119,N_6685,N_7972);
and U9120 (N_9120,N_6702,N_6472);
nand U9121 (N_9121,N_6160,N_7542);
and U9122 (N_9122,N_7653,N_6670);
and U9123 (N_9123,N_6734,N_6512);
nand U9124 (N_9124,N_6805,N_7969);
or U9125 (N_9125,N_6780,N_6291);
and U9126 (N_9126,N_7310,N_6855);
or U9127 (N_9127,N_7865,N_7800);
or U9128 (N_9128,N_7351,N_7746);
and U9129 (N_9129,N_6381,N_7209);
and U9130 (N_9130,N_6503,N_7942);
nand U9131 (N_9131,N_6195,N_6185);
and U9132 (N_9132,N_6825,N_7250);
and U9133 (N_9133,N_7669,N_7363);
xor U9134 (N_9134,N_7167,N_6898);
nand U9135 (N_9135,N_6748,N_7139);
nor U9136 (N_9136,N_7298,N_7265);
or U9137 (N_9137,N_6454,N_7831);
or U9138 (N_9138,N_7414,N_7159);
and U9139 (N_9139,N_6426,N_7982);
or U9140 (N_9140,N_7412,N_7433);
nor U9141 (N_9141,N_7515,N_6940);
and U9142 (N_9142,N_7714,N_6727);
and U9143 (N_9143,N_6462,N_6765);
nand U9144 (N_9144,N_7561,N_7695);
and U9145 (N_9145,N_7953,N_7381);
or U9146 (N_9146,N_6410,N_6426);
nor U9147 (N_9147,N_6674,N_6911);
and U9148 (N_9148,N_7791,N_6364);
nor U9149 (N_9149,N_7556,N_6686);
nand U9150 (N_9150,N_6343,N_7734);
nor U9151 (N_9151,N_7465,N_6541);
nand U9152 (N_9152,N_6705,N_6681);
nor U9153 (N_9153,N_6733,N_6974);
and U9154 (N_9154,N_6024,N_7299);
and U9155 (N_9155,N_6721,N_6812);
or U9156 (N_9156,N_6244,N_6610);
or U9157 (N_9157,N_6136,N_6382);
or U9158 (N_9158,N_7570,N_6807);
and U9159 (N_9159,N_7535,N_7692);
or U9160 (N_9160,N_6606,N_7338);
nor U9161 (N_9161,N_6525,N_7758);
and U9162 (N_9162,N_6654,N_6378);
xnor U9163 (N_9163,N_7118,N_6991);
nand U9164 (N_9164,N_6885,N_6514);
nand U9165 (N_9165,N_7501,N_6159);
nand U9166 (N_9166,N_6735,N_7011);
and U9167 (N_9167,N_7982,N_6501);
nor U9168 (N_9168,N_7283,N_6919);
and U9169 (N_9169,N_6655,N_6895);
nand U9170 (N_9170,N_6332,N_6507);
nor U9171 (N_9171,N_6828,N_6366);
or U9172 (N_9172,N_7268,N_6386);
nand U9173 (N_9173,N_7995,N_6610);
or U9174 (N_9174,N_7739,N_6150);
nor U9175 (N_9175,N_7072,N_7888);
nand U9176 (N_9176,N_7594,N_7181);
and U9177 (N_9177,N_7858,N_7622);
xor U9178 (N_9178,N_6605,N_7049);
nand U9179 (N_9179,N_7247,N_7579);
and U9180 (N_9180,N_7000,N_6837);
or U9181 (N_9181,N_7835,N_6565);
and U9182 (N_9182,N_6421,N_6778);
or U9183 (N_9183,N_6713,N_7602);
nand U9184 (N_9184,N_7556,N_6606);
and U9185 (N_9185,N_6506,N_6016);
nor U9186 (N_9186,N_7165,N_6610);
nand U9187 (N_9187,N_6148,N_6149);
nor U9188 (N_9188,N_6233,N_6745);
and U9189 (N_9189,N_6309,N_6541);
and U9190 (N_9190,N_7978,N_7346);
or U9191 (N_9191,N_7190,N_7787);
nand U9192 (N_9192,N_7647,N_6278);
nand U9193 (N_9193,N_7171,N_6277);
nand U9194 (N_9194,N_7052,N_6254);
xor U9195 (N_9195,N_7698,N_7376);
nand U9196 (N_9196,N_6596,N_7583);
nor U9197 (N_9197,N_6376,N_6076);
nand U9198 (N_9198,N_7711,N_7704);
xnor U9199 (N_9199,N_7716,N_7242);
nor U9200 (N_9200,N_7057,N_6656);
and U9201 (N_9201,N_7432,N_6923);
and U9202 (N_9202,N_7007,N_7388);
and U9203 (N_9203,N_6089,N_7250);
nor U9204 (N_9204,N_7903,N_7259);
nor U9205 (N_9205,N_6548,N_7832);
nand U9206 (N_9206,N_7585,N_7287);
xor U9207 (N_9207,N_7373,N_6845);
nor U9208 (N_9208,N_7927,N_6471);
nor U9209 (N_9209,N_6786,N_7535);
nor U9210 (N_9210,N_7390,N_6971);
nor U9211 (N_9211,N_6907,N_7812);
nand U9212 (N_9212,N_7687,N_7361);
nor U9213 (N_9213,N_6075,N_7189);
nor U9214 (N_9214,N_6806,N_6563);
and U9215 (N_9215,N_6360,N_6777);
nand U9216 (N_9216,N_7352,N_6188);
nand U9217 (N_9217,N_7423,N_6343);
and U9218 (N_9218,N_7075,N_6980);
or U9219 (N_9219,N_6779,N_7585);
or U9220 (N_9220,N_6806,N_7239);
nor U9221 (N_9221,N_6721,N_7641);
or U9222 (N_9222,N_6519,N_7698);
nor U9223 (N_9223,N_6907,N_6120);
and U9224 (N_9224,N_6408,N_6458);
nor U9225 (N_9225,N_7538,N_6730);
xor U9226 (N_9226,N_6432,N_7176);
xnor U9227 (N_9227,N_6059,N_6529);
nor U9228 (N_9228,N_6678,N_7669);
and U9229 (N_9229,N_6979,N_7225);
or U9230 (N_9230,N_7742,N_7718);
and U9231 (N_9231,N_6564,N_7402);
nor U9232 (N_9232,N_6895,N_6225);
nand U9233 (N_9233,N_7998,N_6521);
and U9234 (N_9234,N_7186,N_7867);
nor U9235 (N_9235,N_7293,N_7321);
nand U9236 (N_9236,N_7073,N_6684);
nor U9237 (N_9237,N_6149,N_6703);
and U9238 (N_9238,N_7383,N_7642);
and U9239 (N_9239,N_6920,N_7613);
and U9240 (N_9240,N_6229,N_6803);
or U9241 (N_9241,N_7085,N_6997);
nor U9242 (N_9242,N_6254,N_6675);
nor U9243 (N_9243,N_6531,N_6192);
and U9244 (N_9244,N_6662,N_7386);
and U9245 (N_9245,N_7418,N_7466);
nand U9246 (N_9246,N_6217,N_6436);
or U9247 (N_9247,N_7044,N_6375);
or U9248 (N_9248,N_7660,N_7342);
or U9249 (N_9249,N_7335,N_7214);
nand U9250 (N_9250,N_6034,N_7310);
nand U9251 (N_9251,N_7434,N_6874);
xor U9252 (N_9252,N_7585,N_6631);
nand U9253 (N_9253,N_7626,N_6058);
nand U9254 (N_9254,N_7215,N_6093);
or U9255 (N_9255,N_7576,N_7897);
and U9256 (N_9256,N_6318,N_7556);
or U9257 (N_9257,N_7707,N_7645);
and U9258 (N_9258,N_6977,N_7590);
nand U9259 (N_9259,N_6506,N_6702);
nand U9260 (N_9260,N_6684,N_7741);
or U9261 (N_9261,N_6534,N_6245);
nor U9262 (N_9262,N_7006,N_7129);
nor U9263 (N_9263,N_6823,N_6953);
nor U9264 (N_9264,N_6298,N_6661);
or U9265 (N_9265,N_7586,N_6488);
or U9266 (N_9266,N_6885,N_6137);
nor U9267 (N_9267,N_7043,N_7637);
or U9268 (N_9268,N_7318,N_6890);
nand U9269 (N_9269,N_7052,N_6116);
nor U9270 (N_9270,N_6748,N_6102);
or U9271 (N_9271,N_6781,N_6426);
nor U9272 (N_9272,N_7525,N_7292);
or U9273 (N_9273,N_7679,N_6358);
or U9274 (N_9274,N_6496,N_7180);
or U9275 (N_9275,N_6557,N_7005);
or U9276 (N_9276,N_7162,N_7746);
nor U9277 (N_9277,N_7349,N_6326);
nand U9278 (N_9278,N_7853,N_6573);
nor U9279 (N_9279,N_7531,N_7254);
nand U9280 (N_9280,N_7356,N_6460);
and U9281 (N_9281,N_7204,N_7784);
nor U9282 (N_9282,N_7911,N_6301);
nand U9283 (N_9283,N_6353,N_6912);
nand U9284 (N_9284,N_6084,N_7896);
xor U9285 (N_9285,N_6953,N_7317);
nor U9286 (N_9286,N_7579,N_6916);
nor U9287 (N_9287,N_7226,N_7949);
and U9288 (N_9288,N_7445,N_7424);
or U9289 (N_9289,N_6326,N_7502);
xor U9290 (N_9290,N_7179,N_6298);
nor U9291 (N_9291,N_6697,N_6481);
and U9292 (N_9292,N_6326,N_6305);
nor U9293 (N_9293,N_6298,N_7290);
and U9294 (N_9294,N_7640,N_7413);
nor U9295 (N_9295,N_6091,N_6362);
nand U9296 (N_9296,N_7015,N_6423);
nand U9297 (N_9297,N_7183,N_6387);
nand U9298 (N_9298,N_6440,N_6486);
nor U9299 (N_9299,N_7872,N_7941);
nand U9300 (N_9300,N_7707,N_7323);
or U9301 (N_9301,N_6474,N_7399);
or U9302 (N_9302,N_6316,N_7909);
nor U9303 (N_9303,N_6785,N_7703);
nand U9304 (N_9304,N_7488,N_6881);
nand U9305 (N_9305,N_7039,N_6865);
nor U9306 (N_9306,N_6803,N_7379);
or U9307 (N_9307,N_6000,N_6035);
nor U9308 (N_9308,N_6239,N_6886);
nand U9309 (N_9309,N_7272,N_7717);
xor U9310 (N_9310,N_6865,N_6385);
nor U9311 (N_9311,N_6994,N_6933);
or U9312 (N_9312,N_6583,N_6432);
and U9313 (N_9313,N_7380,N_7382);
and U9314 (N_9314,N_7437,N_6196);
and U9315 (N_9315,N_7425,N_7703);
nand U9316 (N_9316,N_7219,N_6603);
nand U9317 (N_9317,N_6403,N_6110);
and U9318 (N_9318,N_7652,N_7756);
nand U9319 (N_9319,N_6685,N_7448);
and U9320 (N_9320,N_6255,N_6242);
and U9321 (N_9321,N_6508,N_6576);
or U9322 (N_9322,N_7538,N_7088);
nand U9323 (N_9323,N_6773,N_7260);
nand U9324 (N_9324,N_6571,N_6889);
or U9325 (N_9325,N_6682,N_7569);
nor U9326 (N_9326,N_6539,N_6629);
and U9327 (N_9327,N_6043,N_7883);
nor U9328 (N_9328,N_6206,N_6549);
and U9329 (N_9329,N_6624,N_7452);
nand U9330 (N_9330,N_7970,N_7038);
and U9331 (N_9331,N_7410,N_7580);
or U9332 (N_9332,N_7220,N_6217);
nor U9333 (N_9333,N_7190,N_6834);
or U9334 (N_9334,N_6630,N_6598);
nor U9335 (N_9335,N_7929,N_6614);
nand U9336 (N_9336,N_7354,N_7848);
xnor U9337 (N_9337,N_7893,N_7334);
or U9338 (N_9338,N_6737,N_7775);
nand U9339 (N_9339,N_6739,N_7050);
or U9340 (N_9340,N_7716,N_6519);
and U9341 (N_9341,N_7301,N_6321);
nand U9342 (N_9342,N_7756,N_6593);
and U9343 (N_9343,N_7982,N_7286);
or U9344 (N_9344,N_7104,N_7049);
or U9345 (N_9345,N_7619,N_6342);
nor U9346 (N_9346,N_6397,N_6686);
or U9347 (N_9347,N_7356,N_6105);
nor U9348 (N_9348,N_6637,N_6117);
nor U9349 (N_9349,N_7862,N_7883);
nand U9350 (N_9350,N_6560,N_6756);
nor U9351 (N_9351,N_7465,N_7478);
nand U9352 (N_9352,N_7340,N_6438);
or U9353 (N_9353,N_6330,N_6765);
nand U9354 (N_9354,N_7152,N_6121);
and U9355 (N_9355,N_7018,N_6246);
or U9356 (N_9356,N_7562,N_6329);
nor U9357 (N_9357,N_6545,N_6267);
nor U9358 (N_9358,N_7386,N_6081);
or U9359 (N_9359,N_7290,N_7455);
and U9360 (N_9360,N_6587,N_6190);
nor U9361 (N_9361,N_7857,N_7481);
nand U9362 (N_9362,N_7369,N_7646);
or U9363 (N_9363,N_7942,N_7687);
and U9364 (N_9364,N_7365,N_7904);
nand U9365 (N_9365,N_6437,N_7417);
nor U9366 (N_9366,N_7222,N_6160);
nand U9367 (N_9367,N_7319,N_7726);
nor U9368 (N_9368,N_6544,N_7161);
or U9369 (N_9369,N_6950,N_6617);
nor U9370 (N_9370,N_7902,N_7504);
or U9371 (N_9371,N_7394,N_7698);
and U9372 (N_9372,N_7492,N_6216);
nand U9373 (N_9373,N_6599,N_7785);
nor U9374 (N_9374,N_7447,N_6760);
and U9375 (N_9375,N_6343,N_7000);
nand U9376 (N_9376,N_6713,N_6421);
xnor U9377 (N_9377,N_6659,N_7818);
nand U9378 (N_9378,N_7594,N_6638);
nand U9379 (N_9379,N_7392,N_6682);
nor U9380 (N_9380,N_6051,N_7312);
and U9381 (N_9381,N_7073,N_6470);
nand U9382 (N_9382,N_6060,N_7060);
nor U9383 (N_9383,N_6384,N_7938);
and U9384 (N_9384,N_7398,N_7144);
and U9385 (N_9385,N_7041,N_6054);
nand U9386 (N_9386,N_7761,N_6526);
nand U9387 (N_9387,N_6472,N_6042);
or U9388 (N_9388,N_7581,N_6623);
nand U9389 (N_9389,N_7293,N_6064);
or U9390 (N_9390,N_7964,N_6424);
and U9391 (N_9391,N_7198,N_7085);
and U9392 (N_9392,N_7810,N_7313);
nor U9393 (N_9393,N_7810,N_7948);
and U9394 (N_9394,N_7231,N_7341);
and U9395 (N_9395,N_7824,N_6628);
nand U9396 (N_9396,N_6086,N_7292);
and U9397 (N_9397,N_7678,N_6490);
and U9398 (N_9398,N_6423,N_7245);
and U9399 (N_9399,N_7542,N_7247);
or U9400 (N_9400,N_7365,N_6398);
and U9401 (N_9401,N_6831,N_7439);
or U9402 (N_9402,N_7137,N_7661);
or U9403 (N_9403,N_7595,N_6251);
or U9404 (N_9404,N_7393,N_6897);
and U9405 (N_9405,N_6743,N_6836);
or U9406 (N_9406,N_6165,N_7737);
and U9407 (N_9407,N_6734,N_7686);
nand U9408 (N_9408,N_7533,N_7811);
nor U9409 (N_9409,N_6078,N_6308);
or U9410 (N_9410,N_6603,N_6567);
or U9411 (N_9411,N_7690,N_7799);
nor U9412 (N_9412,N_7809,N_6935);
or U9413 (N_9413,N_6353,N_7644);
nand U9414 (N_9414,N_7244,N_7057);
xnor U9415 (N_9415,N_7053,N_6353);
nand U9416 (N_9416,N_7891,N_7687);
and U9417 (N_9417,N_7951,N_6311);
nand U9418 (N_9418,N_7471,N_7948);
nor U9419 (N_9419,N_7836,N_6268);
and U9420 (N_9420,N_6666,N_7751);
nor U9421 (N_9421,N_6939,N_6600);
or U9422 (N_9422,N_6167,N_6657);
nor U9423 (N_9423,N_6159,N_6513);
xor U9424 (N_9424,N_6981,N_6720);
nand U9425 (N_9425,N_7806,N_7447);
or U9426 (N_9426,N_7339,N_6833);
nand U9427 (N_9427,N_6108,N_6551);
nor U9428 (N_9428,N_6891,N_7451);
and U9429 (N_9429,N_7324,N_6039);
nor U9430 (N_9430,N_7287,N_7351);
nand U9431 (N_9431,N_6046,N_7762);
nor U9432 (N_9432,N_6870,N_7794);
nand U9433 (N_9433,N_6635,N_7974);
nor U9434 (N_9434,N_7170,N_7112);
xor U9435 (N_9435,N_7883,N_7658);
nor U9436 (N_9436,N_6477,N_6535);
or U9437 (N_9437,N_6493,N_7827);
nor U9438 (N_9438,N_6273,N_6047);
nand U9439 (N_9439,N_7856,N_7865);
and U9440 (N_9440,N_6621,N_6928);
nor U9441 (N_9441,N_7281,N_6946);
or U9442 (N_9442,N_6337,N_6106);
and U9443 (N_9443,N_6817,N_6333);
nor U9444 (N_9444,N_6328,N_6201);
nand U9445 (N_9445,N_6762,N_6379);
nor U9446 (N_9446,N_7891,N_6177);
nor U9447 (N_9447,N_7668,N_6882);
or U9448 (N_9448,N_7116,N_6188);
xnor U9449 (N_9449,N_7795,N_6181);
and U9450 (N_9450,N_7095,N_6143);
or U9451 (N_9451,N_7120,N_7256);
nor U9452 (N_9452,N_6799,N_6765);
and U9453 (N_9453,N_6663,N_6647);
and U9454 (N_9454,N_6602,N_6815);
or U9455 (N_9455,N_6351,N_7777);
xor U9456 (N_9456,N_6360,N_6648);
or U9457 (N_9457,N_7625,N_6401);
xnor U9458 (N_9458,N_6490,N_6339);
or U9459 (N_9459,N_6636,N_7333);
nand U9460 (N_9460,N_6523,N_7867);
or U9461 (N_9461,N_7690,N_6750);
and U9462 (N_9462,N_7766,N_7257);
or U9463 (N_9463,N_7365,N_6231);
nand U9464 (N_9464,N_7436,N_6710);
or U9465 (N_9465,N_7072,N_7258);
nand U9466 (N_9466,N_6989,N_6721);
and U9467 (N_9467,N_7984,N_7285);
nand U9468 (N_9468,N_7528,N_6212);
or U9469 (N_9469,N_6950,N_6930);
nor U9470 (N_9470,N_6673,N_7174);
nor U9471 (N_9471,N_7918,N_6719);
and U9472 (N_9472,N_6224,N_6170);
nor U9473 (N_9473,N_6275,N_7684);
nor U9474 (N_9474,N_6151,N_6427);
nor U9475 (N_9475,N_7293,N_7438);
nor U9476 (N_9476,N_7697,N_7083);
and U9477 (N_9477,N_7431,N_7083);
or U9478 (N_9478,N_7136,N_6502);
or U9479 (N_9479,N_6321,N_6033);
nand U9480 (N_9480,N_7911,N_6843);
or U9481 (N_9481,N_7228,N_7676);
nor U9482 (N_9482,N_6127,N_6847);
xnor U9483 (N_9483,N_6885,N_7280);
or U9484 (N_9484,N_6460,N_6488);
and U9485 (N_9485,N_7282,N_7571);
xor U9486 (N_9486,N_7042,N_7760);
or U9487 (N_9487,N_6290,N_6406);
nand U9488 (N_9488,N_6763,N_7461);
and U9489 (N_9489,N_7834,N_7338);
or U9490 (N_9490,N_6463,N_7603);
or U9491 (N_9491,N_6936,N_6421);
or U9492 (N_9492,N_7271,N_7909);
or U9493 (N_9493,N_6813,N_6127);
nor U9494 (N_9494,N_6079,N_6294);
nor U9495 (N_9495,N_6577,N_6085);
and U9496 (N_9496,N_6178,N_7768);
or U9497 (N_9497,N_6075,N_6057);
or U9498 (N_9498,N_7071,N_7286);
nor U9499 (N_9499,N_7815,N_6982);
and U9500 (N_9500,N_7227,N_7872);
or U9501 (N_9501,N_6622,N_6619);
nand U9502 (N_9502,N_6246,N_6028);
or U9503 (N_9503,N_6357,N_7009);
and U9504 (N_9504,N_6190,N_7699);
nand U9505 (N_9505,N_7231,N_7270);
nand U9506 (N_9506,N_6122,N_7506);
nand U9507 (N_9507,N_7220,N_7734);
or U9508 (N_9508,N_7642,N_6082);
nand U9509 (N_9509,N_6409,N_7178);
or U9510 (N_9510,N_7411,N_6306);
nor U9511 (N_9511,N_6043,N_6441);
nor U9512 (N_9512,N_6996,N_6830);
and U9513 (N_9513,N_7037,N_6883);
and U9514 (N_9514,N_6542,N_6500);
or U9515 (N_9515,N_6950,N_7601);
nand U9516 (N_9516,N_6666,N_7256);
or U9517 (N_9517,N_6556,N_6525);
and U9518 (N_9518,N_6714,N_6487);
nand U9519 (N_9519,N_7485,N_7848);
nand U9520 (N_9520,N_6958,N_7425);
nor U9521 (N_9521,N_6373,N_6621);
and U9522 (N_9522,N_7698,N_7993);
nand U9523 (N_9523,N_7890,N_7201);
and U9524 (N_9524,N_6921,N_6150);
and U9525 (N_9525,N_6279,N_6182);
and U9526 (N_9526,N_7725,N_7529);
nor U9527 (N_9527,N_7888,N_6720);
and U9528 (N_9528,N_7175,N_6834);
or U9529 (N_9529,N_6800,N_6531);
nor U9530 (N_9530,N_6736,N_7155);
nand U9531 (N_9531,N_7847,N_7961);
or U9532 (N_9532,N_6401,N_7686);
nor U9533 (N_9533,N_7202,N_7586);
nand U9534 (N_9534,N_6846,N_6294);
nand U9535 (N_9535,N_7991,N_6879);
nor U9536 (N_9536,N_6493,N_6489);
and U9537 (N_9537,N_6492,N_7226);
and U9538 (N_9538,N_6643,N_6497);
nand U9539 (N_9539,N_7010,N_6495);
or U9540 (N_9540,N_6014,N_6996);
or U9541 (N_9541,N_6580,N_6204);
nor U9542 (N_9542,N_6659,N_6614);
or U9543 (N_9543,N_7827,N_7836);
nand U9544 (N_9544,N_7641,N_6070);
nand U9545 (N_9545,N_6230,N_6517);
nand U9546 (N_9546,N_6251,N_7955);
nor U9547 (N_9547,N_7589,N_6177);
or U9548 (N_9548,N_7864,N_7593);
and U9549 (N_9549,N_6027,N_7486);
or U9550 (N_9550,N_7624,N_7248);
xnor U9551 (N_9551,N_7933,N_7566);
or U9552 (N_9552,N_6063,N_7152);
and U9553 (N_9553,N_7132,N_6188);
nand U9554 (N_9554,N_6040,N_6163);
and U9555 (N_9555,N_6018,N_7778);
and U9556 (N_9556,N_6860,N_6803);
nand U9557 (N_9557,N_6318,N_7675);
nand U9558 (N_9558,N_7948,N_7453);
and U9559 (N_9559,N_6670,N_6339);
nor U9560 (N_9560,N_6389,N_6793);
or U9561 (N_9561,N_6712,N_6539);
nor U9562 (N_9562,N_6576,N_6449);
or U9563 (N_9563,N_6991,N_7944);
nand U9564 (N_9564,N_6742,N_7392);
nand U9565 (N_9565,N_6297,N_7807);
or U9566 (N_9566,N_7286,N_6400);
nand U9567 (N_9567,N_6380,N_6553);
nand U9568 (N_9568,N_7075,N_6488);
and U9569 (N_9569,N_6484,N_7131);
or U9570 (N_9570,N_7454,N_7183);
and U9571 (N_9571,N_6631,N_7155);
xnor U9572 (N_9572,N_7721,N_6680);
nand U9573 (N_9573,N_7345,N_7292);
nor U9574 (N_9574,N_7607,N_6987);
and U9575 (N_9575,N_6154,N_7435);
and U9576 (N_9576,N_7054,N_7454);
or U9577 (N_9577,N_7579,N_7925);
and U9578 (N_9578,N_7688,N_6044);
nand U9579 (N_9579,N_7637,N_6563);
nand U9580 (N_9580,N_7891,N_6569);
nand U9581 (N_9581,N_6724,N_7758);
and U9582 (N_9582,N_7544,N_6834);
nor U9583 (N_9583,N_7339,N_6769);
and U9584 (N_9584,N_6835,N_7773);
nand U9585 (N_9585,N_7527,N_6151);
nand U9586 (N_9586,N_6033,N_7178);
nand U9587 (N_9587,N_6115,N_6940);
or U9588 (N_9588,N_7943,N_7400);
nor U9589 (N_9589,N_7018,N_7215);
nand U9590 (N_9590,N_7806,N_7665);
nor U9591 (N_9591,N_7444,N_7275);
or U9592 (N_9592,N_7791,N_6738);
and U9593 (N_9593,N_6896,N_7494);
or U9594 (N_9594,N_6583,N_7259);
or U9595 (N_9595,N_6352,N_7103);
and U9596 (N_9596,N_7148,N_6951);
nand U9597 (N_9597,N_6726,N_6741);
nand U9598 (N_9598,N_7333,N_6765);
and U9599 (N_9599,N_6223,N_7695);
and U9600 (N_9600,N_7534,N_7505);
nor U9601 (N_9601,N_6556,N_6209);
nand U9602 (N_9602,N_6948,N_6535);
nor U9603 (N_9603,N_6195,N_6786);
nor U9604 (N_9604,N_7527,N_6907);
and U9605 (N_9605,N_7722,N_7620);
nand U9606 (N_9606,N_7525,N_6937);
or U9607 (N_9607,N_7173,N_7054);
and U9608 (N_9608,N_6547,N_7367);
or U9609 (N_9609,N_6801,N_7605);
and U9610 (N_9610,N_6337,N_7506);
nor U9611 (N_9611,N_6862,N_6139);
or U9612 (N_9612,N_6712,N_6976);
or U9613 (N_9613,N_7475,N_6219);
or U9614 (N_9614,N_7778,N_6208);
nor U9615 (N_9615,N_6356,N_6734);
or U9616 (N_9616,N_6945,N_6823);
nor U9617 (N_9617,N_6276,N_6645);
or U9618 (N_9618,N_7950,N_7383);
nand U9619 (N_9619,N_7877,N_6260);
xor U9620 (N_9620,N_6757,N_7617);
or U9621 (N_9621,N_7748,N_7674);
and U9622 (N_9622,N_6590,N_7283);
nand U9623 (N_9623,N_7571,N_7704);
xnor U9624 (N_9624,N_7550,N_7906);
or U9625 (N_9625,N_6623,N_6713);
or U9626 (N_9626,N_7509,N_7645);
and U9627 (N_9627,N_6821,N_6750);
nor U9628 (N_9628,N_6948,N_7740);
and U9629 (N_9629,N_6432,N_6303);
nor U9630 (N_9630,N_6380,N_7144);
or U9631 (N_9631,N_7462,N_6653);
nor U9632 (N_9632,N_7969,N_6738);
xor U9633 (N_9633,N_6638,N_6517);
xor U9634 (N_9634,N_7957,N_6269);
nand U9635 (N_9635,N_7283,N_7730);
nor U9636 (N_9636,N_6104,N_6298);
or U9637 (N_9637,N_6864,N_7134);
and U9638 (N_9638,N_7198,N_7418);
xnor U9639 (N_9639,N_7747,N_7259);
nor U9640 (N_9640,N_7928,N_6442);
and U9641 (N_9641,N_7731,N_6410);
nor U9642 (N_9642,N_6682,N_6504);
nand U9643 (N_9643,N_7599,N_6836);
nor U9644 (N_9644,N_6314,N_6488);
or U9645 (N_9645,N_7650,N_7576);
or U9646 (N_9646,N_7339,N_7360);
and U9647 (N_9647,N_6534,N_6557);
nor U9648 (N_9648,N_7656,N_7937);
xnor U9649 (N_9649,N_6640,N_6784);
nand U9650 (N_9650,N_7043,N_7396);
and U9651 (N_9651,N_7360,N_7202);
and U9652 (N_9652,N_6863,N_7859);
nor U9653 (N_9653,N_6010,N_7684);
nand U9654 (N_9654,N_6823,N_6855);
nor U9655 (N_9655,N_7108,N_6361);
and U9656 (N_9656,N_6737,N_6996);
xnor U9657 (N_9657,N_7139,N_7912);
nand U9658 (N_9658,N_7284,N_6776);
nor U9659 (N_9659,N_6085,N_6319);
nand U9660 (N_9660,N_6448,N_6474);
nor U9661 (N_9661,N_7305,N_7526);
xnor U9662 (N_9662,N_7060,N_6328);
or U9663 (N_9663,N_6625,N_7874);
and U9664 (N_9664,N_6145,N_6361);
or U9665 (N_9665,N_6429,N_6708);
nor U9666 (N_9666,N_6141,N_6989);
nor U9667 (N_9667,N_6675,N_7011);
nand U9668 (N_9668,N_6378,N_7605);
nand U9669 (N_9669,N_7840,N_6628);
nor U9670 (N_9670,N_6950,N_7541);
nor U9671 (N_9671,N_7082,N_6390);
or U9672 (N_9672,N_7859,N_7175);
and U9673 (N_9673,N_7739,N_6767);
or U9674 (N_9674,N_7016,N_6797);
nor U9675 (N_9675,N_6895,N_7007);
nor U9676 (N_9676,N_6106,N_7689);
nor U9677 (N_9677,N_6035,N_6158);
and U9678 (N_9678,N_7613,N_7096);
and U9679 (N_9679,N_7130,N_7122);
or U9680 (N_9680,N_6560,N_7979);
nor U9681 (N_9681,N_7766,N_7566);
or U9682 (N_9682,N_6860,N_6939);
nor U9683 (N_9683,N_6204,N_6094);
and U9684 (N_9684,N_7775,N_6003);
nand U9685 (N_9685,N_7386,N_6600);
nand U9686 (N_9686,N_7843,N_7006);
or U9687 (N_9687,N_7715,N_7446);
nand U9688 (N_9688,N_7790,N_6902);
nand U9689 (N_9689,N_7023,N_6707);
nor U9690 (N_9690,N_6813,N_6040);
nand U9691 (N_9691,N_7759,N_7757);
and U9692 (N_9692,N_7447,N_6300);
nand U9693 (N_9693,N_6365,N_7770);
nor U9694 (N_9694,N_6415,N_7946);
nor U9695 (N_9695,N_7339,N_6828);
nand U9696 (N_9696,N_6704,N_6109);
nor U9697 (N_9697,N_7319,N_6912);
and U9698 (N_9698,N_6373,N_7241);
nor U9699 (N_9699,N_7780,N_7925);
or U9700 (N_9700,N_7764,N_7182);
and U9701 (N_9701,N_7403,N_6244);
nor U9702 (N_9702,N_6975,N_6582);
nor U9703 (N_9703,N_7781,N_7369);
nor U9704 (N_9704,N_7440,N_6382);
and U9705 (N_9705,N_7905,N_6537);
nor U9706 (N_9706,N_7423,N_6272);
nor U9707 (N_9707,N_6528,N_7658);
nor U9708 (N_9708,N_6627,N_6882);
or U9709 (N_9709,N_7320,N_6273);
and U9710 (N_9710,N_7734,N_7038);
or U9711 (N_9711,N_7706,N_7505);
nand U9712 (N_9712,N_7843,N_6663);
nor U9713 (N_9713,N_6158,N_6349);
or U9714 (N_9714,N_7638,N_7684);
or U9715 (N_9715,N_7391,N_7394);
nor U9716 (N_9716,N_7544,N_6312);
or U9717 (N_9717,N_6598,N_6492);
and U9718 (N_9718,N_6897,N_7810);
nand U9719 (N_9719,N_7445,N_6992);
nor U9720 (N_9720,N_7146,N_7892);
nand U9721 (N_9721,N_6370,N_7641);
and U9722 (N_9722,N_6725,N_7615);
or U9723 (N_9723,N_6833,N_6641);
and U9724 (N_9724,N_7682,N_7273);
nand U9725 (N_9725,N_6824,N_6445);
or U9726 (N_9726,N_6893,N_6292);
and U9727 (N_9727,N_6302,N_7768);
nand U9728 (N_9728,N_6816,N_6567);
and U9729 (N_9729,N_6962,N_7741);
nand U9730 (N_9730,N_7783,N_6451);
and U9731 (N_9731,N_6364,N_6917);
nand U9732 (N_9732,N_7871,N_6538);
nor U9733 (N_9733,N_7795,N_7593);
and U9734 (N_9734,N_7691,N_6400);
nand U9735 (N_9735,N_6047,N_7629);
xnor U9736 (N_9736,N_6039,N_6044);
and U9737 (N_9737,N_7015,N_6844);
nand U9738 (N_9738,N_6249,N_7329);
nand U9739 (N_9739,N_7338,N_7069);
nand U9740 (N_9740,N_6431,N_6250);
nor U9741 (N_9741,N_6663,N_6075);
nand U9742 (N_9742,N_7209,N_6580);
nand U9743 (N_9743,N_7835,N_7193);
and U9744 (N_9744,N_6896,N_6195);
and U9745 (N_9745,N_7872,N_6007);
nand U9746 (N_9746,N_6026,N_7514);
nand U9747 (N_9747,N_7750,N_7114);
and U9748 (N_9748,N_7616,N_6421);
and U9749 (N_9749,N_7019,N_7291);
and U9750 (N_9750,N_7168,N_7928);
and U9751 (N_9751,N_6821,N_7827);
nor U9752 (N_9752,N_7749,N_6074);
nand U9753 (N_9753,N_7382,N_6486);
nor U9754 (N_9754,N_7240,N_7958);
or U9755 (N_9755,N_6390,N_6333);
nor U9756 (N_9756,N_7321,N_6365);
nand U9757 (N_9757,N_7890,N_7678);
or U9758 (N_9758,N_7664,N_7649);
nor U9759 (N_9759,N_6300,N_7053);
or U9760 (N_9760,N_7675,N_7504);
or U9761 (N_9761,N_6422,N_7120);
or U9762 (N_9762,N_6927,N_6637);
nand U9763 (N_9763,N_7846,N_6419);
nor U9764 (N_9764,N_7750,N_6690);
xor U9765 (N_9765,N_7941,N_7521);
xor U9766 (N_9766,N_6699,N_6957);
nor U9767 (N_9767,N_7069,N_7183);
nor U9768 (N_9768,N_6935,N_6972);
or U9769 (N_9769,N_7225,N_6819);
and U9770 (N_9770,N_7303,N_7365);
nor U9771 (N_9771,N_7299,N_6717);
or U9772 (N_9772,N_6460,N_6615);
nor U9773 (N_9773,N_6092,N_7191);
nand U9774 (N_9774,N_6220,N_7040);
and U9775 (N_9775,N_7583,N_7008);
or U9776 (N_9776,N_6226,N_6962);
and U9777 (N_9777,N_7630,N_7017);
nand U9778 (N_9778,N_6051,N_6608);
nand U9779 (N_9779,N_6019,N_7103);
nor U9780 (N_9780,N_7485,N_6976);
and U9781 (N_9781,N_6658,N_7536);
or U9782 (N_9782,N_7885,N_6721);
nand U9783 (N_9783,N_6680,N_6182);
nand U9784 (N_9784,N_7225,N_6122);
or U9785 (N_9785,N_6376,N_6762);
nor U9786 (N_9786,N_7602,N_6534);
and U9787 (N_9787,N_6286,N_7483);
nand U9788 (N_9788,N_7419,N_7253);
and U9789 (N_9789,N_6429,N_6890);
and U9790 (N_9790,N_6275,N_6763);
or U9791 (N_9791,N_7639,N_6182);
and U9792 (N_9792,N_7149,N_6165);
or U9793 (N_9793,N_6359,N_7191);
xnor U9794 (N_9794,N_6526,N_6859);
or U9795 (N_9795,N_7779,N_6156);
and U9796 (N_9796,N_6716,N_7461);
nand U9797 (N_9797,N_7560,N_6625);
nor U9798 (N_9798,N_7884,N_6299);
nand U9799 (N_9799,N_6492,N_6234);
nor U9800 (N_9800,N_6137,N_6866);
and U9801 (N_9801,N_6695,N_6015);
nand U9802 (N_9802,N_7434,N_6889);
nor U9803 (N_9803,N_7505,N_7952);
or U9804 (N_9804,N_7868,N_6549);
nand U9805 (N_9805,N_7385,N_7873);
and U9806 (N_9806,N_7737,N_6476);
or U9807 (N_9807,N_6249,N_7826);
or U9808 (N_9808,N_6104,N_7542);
and U9809 (N_9809,N_6679,N_7627);
or U9810 (N_9810,N_6765,N_7837);
or U9811 (N_9811,N_7321,N_6959);
nor U9812 (N_9812,N_7465,N_6580);
nor U9813 (N_9813,N_7636,N_6621);
nor U9814 (N_9814,N_7152,N_6729);
or U9815 (N_9815,N_7189,N_7320);
nand U9816 (N_9816,N_7866,N_6327);
nand U9817 (N_9817,N_6521,N_6190);
and U9818 (N_9818,N_7920,N_6735);
and U9819 (N_9819,N_7603,N_6028);
nand U9820 (N_9820,N_7838,N_7127);
nand U9821 (N_9821,N_6300,N_6013);
nand U9822 (N_9822,N_7104,N_6536);
nor U9823 (N_9823,N_6735,N_7070);
or U9824 (N_9824,N_7200,N_7812);
nand U9825 (N_9825,N_7561,N_7066);
nand U9826 (N_9826,N_7044,N_6355);
xor U9827 (N_9827,N_7421,N_6328);
nor U9828 (N_9828,N_7899,N_6579);
and U9829 (N_9829,N_6551,N_6172);
and U9830 (N_9830,N_7248,N_6943);
and U9831 (N_9831,N_6643,N_6227);
nand U9832 (N_9832,N_7636,N_6677);
or U9833 (N_9833,N_7137,N_6682);
nor U9834 (N_9834,N_7965,N_7286);
or U9835 (N_9835,N_7829,N_6010);
or U9836 (N_9836,N_7998,N_6478);
nand U9837 (N_9837,N_6237,N_6856);
or U9838 (N_9838,N_6038,N_7203);
and U9839 (N_9839,N_7834,N_7919);
nand U9840 (N_9840,N_7434,N_6708);
nor U9841 (N_9841,N_6802,N_6614);
and U9842 (N_9842,N_6091,N_6088);
nand U9843 (N_9843,N_7857,N_7126);
nor U9844 (N_9844,N_7726,N_7968);
or U9845 (N_9845,N_7388,N_7696);
and U9846 (N_9846,N_7285,N_7686);
and U9847 (N_9847,N_6373,N_7101);
nand U9848 (N_9848,N_7630,N_7192);
nor U9849 (N_9849,N_6966,N_6128);
nor U9850 (N_9850,N_6919,N_7909);
and U9851 (N_9851,N_7855,N_7246);
nor U9852 (N_9852,N_6579,N_7347);
xor U9853 (N_9853,N_6206,N_6703);
or U9854 (N_9854,N_7543,N_6144);
nand U9855 (N_9855,N_6627,N_6587);
and U9856 (N_9856,N_7202,N_6819);
nand U9857 (N_9857,N_7637,N_7439);
nand U9858 (N_9858,N_6341,N_7984);
and U9859 (N_9859,N_6104,N_7837);
nor U9860 (N_9860,N_6184,N_6930);
nor U9861 (N_9861,N_7364,N_7008);
and U9862 (N_9862,N_7484,N_7541);
or U9863 (N_9863,N_7601,N_6988);
or U9864 (N_9864,N_6824,N_6191);
nor U9865 (N_9865,N_6435,N_6654);
or U9866 (N_9866,N_7909,N_6288);
or U9867 (N_9867,N_6423,N_7669);
or U9868 (N_9868,N_7461,N_7311);
or U9869 (N_9869,N_6546,N_7679);
nor U9870 (N_9870,N_6624,N_6325);
xnor U9871 (N_9871,N_6851,N_6688);
or U9872 (N_9872,N_6007,N_6067);
and U9873 (N_9873,N_7966,N_7135);
nand U9874 (N_9874,N_7418,N_7773);
nand U9875 (N_9875,N_7112,N_6896);
nor U9876 (N_9876,N_7952,N_7621);
or U9877 (N_9877,N_7735,N_6653);
or U9878 (N_9878,N_6574,N_7500);
nand U9879 (N_9879,N_7033,N_7440);
nor U9880 (N_9880,N_6510,N_6893);
nand U9881 (N_9881,N_6392,N_6120);
and U9882 (N_9882,N_7864,N_7847);
and U9883 (N_9883,N_7552,N_6139);
and U9884 (N_9884,N_7863,N_6320);
and U9885 (N_9885,N_7475,N_7788);
nand U9886 (N_9886,N_6683,N_7345);
or U9887 (N_9887,N_7869,N_7820);
nand U9888 (N_9888,N_6464,N_6279);
nor U9889 (N_9889,N_6928,N_7527);
nand U9890 (N_9890,N_6405,N_7139);
or U9891 (N_9891,N_7868,N_6164);
nand U9892 (N_9892,N_6093,N_6116);
and U9893 (N_9893,N_7071,N_7898);
or U9894 (N_9894,N_7325,N_7355);
and U9895 (N_9895,N_6434,N_6087);
or U9896 (N_9896,N_6011,N_7499);
nor U9897 (N_9897,N_6623,N_7039);
or U9898 (N_9898,N_6221,N_7423);
nor U9899 (N_9899,N_7173,N_6970);
nand U9900 (N_9900,N_7536,N_7150);
nor U9901 (N_9901,N_7926,N_6852);
or U9902 (N_9902,N_6559,N_7212);
or U9903 (N_9903,N_6674,N_6113);
nand U9904 (N_9904,N_7339,N_6332);
or U9905 (N_9905,N_6422,N_7651);
or U9906 (N_9906,N_7435,N_7444);
or U9907 (N_9907,N_6951,N_7709);
nor U9908 (N_9908,N_7804,N_7038);
nand U9909 (N_9909,N_6473,N_6553);
and U9910 (N_9910,N_7434,N_7259);
nor U9911 (N_9911,N_7074,N_6992);
nor U9912 (N_9912,N_6981,N_6430);
and U9913 (N_9913,N_6016,N_7863);
nor U9914 (N_9914,N_6991,N_6577);
nand U9915 (N_9915,N_7813,N_6703);
nor U9916 (N_9916,N_6178,N_7009);
nor U9917 (N_9917,N_7397,N_6572);
or U9918 (N_9918,N_7169,N_7699);
nor U9919 (N_9919,N_7987,N_7633);
xnor U9920 (N_9920,N_6045,N_7249);
nor U9921 (N_9921,N_6789,N_6136);
nand U9922 (N_9922,N_7046,N_6814);
nand U9923 (N_9923,N_6636,N_6653);
xor U9924 (N_9924,N_6266,N_7189);
nand U9925 (N_9925,N_6006,N_7183);
and U9926 (N_9926,N_6489,N_6836);
or U9927 (N_9927,N_6806,N_6494);
and U9928 (N_9928,N_7467,N_6523);
or U9929 (N_9929,N_6164,N_6056);
nand U9930 (N_9930,N_6951,N_6621);
and U9931 (N_9931,N_7969,N_6942);
nand U9932 (N_9932,N_6174,N_6063);
or U9933 (N_9933,N_6487,N_6927);
xnor U9934 (N_9934,N_7753,N_6663);
nand U9935 (N_9935,N_6646,N_7162);
and U9936 (N_9936,N_7311,N_6039);
xor U9937 (N_9937,N_7950,N_6322);
nand U9938 (N_9938,N_7603,N_7681);
and U9939 (N_9939,N_6540,N_7640);
and U9940 (N_9940,N_7955,N_7655);
and U9941 (N_9941,N_6151,N_6599);
and U9942 (N_9942,N_7300,N_6748);
or U9943 (N_9943,N_7645,N_6882);
or U9944 (N_9944,N_6081,N_7652);
nand U9945 (N_9945,N_7996,N_7195);
or U9946 (N_9946,N_7479,N_6593);
xor U9947 (N_9947,N_6439,N_6529);
nand U9948 (N_9948,N_7220,N_6135);
nor U9949 (N_9949,N_6650,N_6025);
or U9950 (N_9950,N_7240,N_7738);
or U9951 (N_9951,N_6639,N_7760);
nand U9952 (N_9952,N_6382,N_7898);
nand U9953 (N_9953,N_6773,N_6877);
nor U9954 (N_9954,N_6310,N_7112);
nor U9955 (N_9955,N_7538,N_6040);
nor U9956 (N_9956,N_6426,N_7758);
and U9957 (N_9957,N_7706,N_7117);
or U9958 (N_9958,N_6122,N_6080);
and U9959 (N_9959,N_6149,N_6123);
nor U9960 (N_9960,N_7451,N_7016);
and U9961 (N_9961,N_7746,N_6790);
and U9962 (N_9962,N_7688,N_6258);
nor U9963 (N_9963,N_6947,N_7764);
nor U9964 (N_9964,N_7097,N_7607);
or U9965 (N_9965,N_7401,N_6864);
nand U9966 (N_9966,N_7127,N_7657);
and U9967 (N_9967,N_6383,N_6278);
and U9968 (N_9968,N_6874,N_6007);
nand U9969 (N_9969,N_6933,N_7100);
or U9970 (N_9970,N_6670,N_7185);
or U9971 (N_9971,N_6978,N_7214);
and U9972 (N_9972,N_6241,N_6778);
and U9973 (N_9973,N_6891,N_7050);
nand U9974 (N_9974,N_7664,N_7432);
or U9975 (N_9975,N_7618,N_7879);
nand U9976 (N_9976,N_6145,N_6728);
nand U9977 (N_9977,N_6143,N_7027);
nor U9978 (N_9978,N_7699,N_6564);
nand U9979 (N_9979,N_7535,N_7083);
or U9980 (N_9980,N_7883,N_6245);
and U9981 (N_9981,N_7882,N_6904);
or U9982 (N_9982,N_6456,N_6701);
nand U9983 (N_9983,N_6843,N_6444);
nand U9984 (N_9984,N_6815,N_7019);
nor U9985 (N_9985,N_7520,N_6362);
or U9986 (N_9986,N_7166,N_6472);
and U9987 (N_9987,N_6262,N_7958);
nor U9988 (N_9988,N_7433,N_7872);
nand U9989 (N_9989,N_7226,N_7833);
nor U9990 (N_9990,N_6896,N_7898);
and U9991 (N_9991,N_7561,N_6702);
and U9992 (N_9992,N_6807,N_7464);
nor U9993 (N_9993,N_6194,N_6662);
nand U9994 (N_9994,N_6669,N_7931);
and U9995 (N_9995,N_7764,N_6179);
or U9996 (N_9996,N_7968,N_6817);
and U9997 (N_9997,N_6792,N_6005);
and U9998 (N_9998,N_7500,N_7284);
nor U9999 (N_9999,N_6251,N_7640);
nand UO_0 (O_0,N_9795,N_9215);
and UO_1 (O_1,N_8053,N_8403);
nand UO_2 (O_2,N_9762,N_9454);
and UO_3 (O_3,N_9477,N_8899);
or UO_4 (O_4,N_8726,N_8978);
xor UO_5 (O_5,N_8027,N_9276);
xor UO_6 (O_6,N_8633,N_9257);
or UO_7 (O_7,N_9888,N_8811);
nor UO_8 (O_8,N_9841,N_8764);
xor UO_9 (O_9,N_9283,N_9529);
or UO_10 (O_10,N_9719,N_9449);
and UO_11 (O_11,N_9740,N_8971);
or UO_12 (O_12,N_9839,N_9993);
nor UO_13 (O_13,N_9510,N_9297);
and UO_14 (O_14,N_9524,N_8320);
nor UO_15 (O_15,N_8526,N_9899);
nand UO_16 (O_16,N_9934,N_9351);
nand UO_17 (O_17,N_9229,N_8779);
nand UO_18 (O_18,N_9178,N_9633);
nor UO_19 (O_19,N_8574,N_9213);
or UO_20 (O_20,N_9159,N_8326);
or UO_21 (O_21,N_9954,N_9600);
and UO_22 (O_22,N_8641,N_8891);
and UO_23 (O_23,N_8478,N_9165);
nor UO_24 (O_24,N_9258,N_8557);
and UO_25 (O_25,N_9079,N_9402);
xnor UO_26 (O_26,N_9866,N_8244);
nor UO_27 (O_27,N_9830,N_8289);
nor UO_28 (O_28,N_9743,N_8437);
or UO_29 (O_29,N_9950,N_8904);
nand UO_30 (O_30,N_8803,N_8112);
nand UO_31 (O_31,N_9733,N_8008);
nand UO_32 (O_32,N_8973,N_8265);
and UO_33 (O_33,N_8476,N_8900);
and UO_34 (O_34,N_9472,N_9628);
nand UO_35 (O_35,N_8506,N_9667);
or UO_36 (O_36,N_8657,N_9296);
and UO_37 (O_37,N_9167,N_8037);
and UO_38 (O_38,N_8511,N_8042);
xnor UO_39 (O_39,N_9038,N_9148);
nand UO_40 (O_40,N_8233,N_9071);
or UO_41 (O_41,N_9797,N_8603);
nor UO_42 (O_42,N_8194,N_8737);
nor UO_43 (O_43,N_8531,N_9826);
and UO_44 (O_44,N_8733,N_9659);
nand UO_45 (O_45,N_9509,N_8102);
xor UO_46 (O_46,N_8043,N_9308);
nand UO_47 (O_47,N_9483,N_8386);
and UO_48 (O_48,N_8409,N_9371);
or UO_49 (O_49,N_8601,N_8154);
nand UO_50 (O_50,N_8463,N_8308);
nand UO_51 (O_51,N_9379,N_8746);
and UO_52 (O_52,N_9244,N_8932);
and UO_53 (O_53,N_8290,N_8253);
or UO_54 (O_54,N_9340,N_8843);
nor UO_55 (O_55,N_9066,N_9879);
nand UO_56 (O_56,N_8470,N_9890);
or UO_57 (O_57,N_8549,N_8399);
and UO_58 (O_58,N_8938,N_9043);
nand UO_59 (O_59,N_9317,N_8946);
or UO_60 (O_60,N_9228,N_9173);
nor UO_61 (O_61,N_9818,N_8040);
nor UO_62 (O_62,N_9282,N_8237);
nand UO_63 (O_63,N_8931,N_9534);
or UO_64 (O_64,N_9774,N_9551);
or UO_65 (O_65,N_9288,N_9220);
or UO_66 (O_66,N_9344,N_8546);
and UO_67 (O_67,N_8278,N_8353);
or UO_68 (O_68,N_9267,N_8302);
and UO_69 (O_69,N_8280,N_9124);
nor UO_70 (O_70,N_8520,N_8689);
and UO_71 (O_71,N_9722,N_8207);
nand UO_72 (O_72,N_9717,N_8268);
or UO_73 (O_73,N_9552,N_9238);
nand UO_74 (O_74,N_9876,N_8175);
and UO_75 (O_75,N_9655,N_8436);
nand UO_76 (O_76,N_9753,N_9977);
and UO_77 (O_77,N_9156,N_9983);
nor UO_78 (O_78,N_8365,N_9496);
and UO_79 (O_79,N_9251,N_9764);
nor UO_80 (O_80,N_8793,N_8415);
nand UO_81 (O_81,N_8044,N_8515);
nor UO_82 (O_82,N_8917,N_9759);
nand UO_83 (O_83,N_9959,N_8431);
nand UO_84 (O_84,N_8611,N_8024);
and UO_85 (O_85,N_9834,N_8056);
and UO_86 (O_86,N_9180,N_9651);
or UO_87 (O_87,N_9923,N_9532);
nand UO_88 (O_88,N_8490,N_8495);
or UO_89 (O_89,N_8128,N_8393);
nand UO_90 (O_90,N_9768,N_9381);
nand UO_91 (O_91,N_8615,N_9395);
or UO_92 (O_92,N_8923,N_9003);
nor UO_93 (O_93,N_9973,N_8929);
nor UO_94 (O_94,N_9627,N_9137);
and UO_95 (O_95,N_9144,N_9788);
or UO_96 (O_96,N_8139,N_8903);
and UO_97 (O_97,N_9987,N_8573);
and UO_98 (O_98,N_8665,N_9745);
nand UO_99 (O_99,N_8853,N_9514);
or UO_100 (O_100,N_8823,N_9341);
and UO_101 (O_101,N_9186,N_9166);
and UO_102 (O_102,N_9550,N_8831);
nor UO_103 (O_103,N_9869,N_8387);
and UO_104 (O_104,N_8739,N_8980);
and UO_105 (O_105,N_8182,N_8167);
or UO_106 (O_106,N_8335,N_9274);
and UO_107 (O_107,N_8632,N_9965);
nand UO_108 (O_108,N_9938,N_9980);
and UO_109 (O_109,N_9356,N_9836);
nor UO_110 (O_110,N_8169,N_9968);
and UO_111 (O_111,N_9578,N_8304);
and UO_112 (O_112,N_8795,N_8006);
nand UO_113 (O_113,N_8510,N_9737);
or UO_114 (O_114,N_9445,N_8584);
nor UO_115 (O_115,N_8448,N_9117);
nor UO_116 (O_116,N_9320,N_9061);
and UO_117 (O_117,N_9666,N_8004);
nand UO_118 (O_118,N_9595,N_8566);
or UO_119 (O_119,N_9948,N_8597);
nand UO_120 (O_120,N_8508,N_8651);
and UO_121 (O_121,N_8408,N_9937);
or UO_122 (O_122,N_9140,N_9732);
and UO_123 (O_123,N_9766,N_8872);
and UO_124 (O_124,N_9527,N_9261);
or UO_125 (O_125,N_9077,N_9598);
and UO_126 (O_126,N_9898,N_8367);
and UO_127 (O_127,N_9746,N_9988);
or UO_128 (O_128,N_9011,N_9444);
or UO_129 (O_129,N_8672,N_8878);
or UO_130 (O_130,N_8455,N_8196);
nor UO_131 (O_131,N_8125,N_9157);
and UO_132 (O_132,N_9918,N_8228);
or UO_133 (O_133,N_8886,N_9252);
nor UO_134 (O_134,N_8357,N_8921);
or UO_135 (O_135,N_8071,N_9591);
nor UO_136 (O_136,N_8781,N_9913);
and UO_137 (O_137,N_9045,N_9548);
nand UO_138 (O_138,N_9602,N_9645);
nor UO_139 (O_139,N_9592,N_8569);
nand UO_140 (O_140,N_9129,N_9330);
nand UO_141 (O_141,N_8579,N_9603);
xor UO_142 (O_142,N_8619,N_8673);
and UO_143 (O_143,N_8636,N_8119);
nor UO_144 (O_144,N_8306,N_8682);
nand UO_145 (O_145,N_8930,N_8854);
and UO_146 (O_146,N_9136,N_8589);
nand UO_147 (O_147,N_8558,N_8956);
nor UO_148 (O_148,N_8951,N_8765);
nor UO_149 (O_149,N_8761,N_8411);
xor UO_150 (O_150,N_8227,N_8539);
or UO_151 (O_151,N_9217,N_9275);
nand UO_152 (O_152,N_9232,N_9845);
nand UO_153 (O_153,N_8688,N_9366);
and UO_154 (O_154,N_8457,N_9599);
nor UO_155 (O_155,N_8235,N_8276);
or UO_156 (O_156,N_9690,N_9616);
and UO_157 (O_157,N_9110,N_8679);
or UO_158 (O_158,N_9424,N_8991);
nor UO_159 (O_159,N_9631,N_8492);
nor UO_160 (O_160,N_8618,N_9706);
nor UO_161 (O_161,N_8552,N_8631);
and UO_162 (O_162,N_8816,N_9100);
and UO_163 (O_163,N_9469,N_8936);
or UO_164 (O_164,N_8583,N_8146);
nor UO_165 (O_165,N_9513,N_9546);
and UO_166 (O_166,N_9498,N_8525);
nor UO_167 (O_167,N_9787,N_9557);
and UO_168 (O_168,N_9701,N_9189);
nor UO_169 (O_169,N_9908,N_8430);
nand UO_170 (O_170,N_9139,N_8143);
nand UO_171 (O_171,N_8887,N_8116);
or UO_172 (O_172,N_8544,N_9052);
and UO_173 (O_173,N_8255,N_9847);
or UO_174 (O_174,N_9790,N_9319);
xor UO_175 (O_175,N_8216,N_8987);
nand UO_176 (O_176,N_8469,N_9596);
nor UO_177 (O_177,N_8787,N_8523);
or UO_178 (O_178,N_8693,N_8661);
or UO_179 (O_179,N_8424,N_9235);
xor UO_180 (O_180,N_9280,N_8806);
nand UO_181 (O_181,N_9375,N_9806);
nor UO_182 (O_182,N_9799,N_9700);
xnor UO_183 (O_183,N_9254,N_8848);
and UO_184 (O_184,N_8874,N_8261);
and UO_185 (O_185,N_8701,N_9050);
and UO_186 (O_186,N_9922,N_9128);
nand UO_187 (O_187,N_9930,N_8660);
or UO_188 (O_188,N_8824,N_9972);
or UO_189 (O_189,N_9624,N_8485);
or UO_190 (O_190,N_9162,N_9486);
nor UO_191 (O_191,N_8076,N_9284);
or UO_192 (O_192,N_9369,N_9864);
nand UO_193 (O_193,N_8217,N_9104);
nand UO_194 (O_194,N_9540,N_9115);
and UO_195 (O_195,N_8988,N_9002);
nor UO_196 (O_196,N_8427,N_9131);
nor UO_197 (O_197,N_8942,N_9149);
or UO_198 (O_198,N_8590,N_8814);
nor UO_199 (O_199,N_9095,N_8807);
or UO_200 (O_200,N_9141,N_9756);
and UO_201 (O_201,N_9322,N_8364);
or UO_202 (O_202,N_8949,N_9384);
nand UO_203 (O_203,N_8108,N_9412);
or UO_204 (O_204,N_9125,N_9408);
and UO_205 (O_205,N_9023,N_8029);
and UO_206 (O_206,N_8686,N_8471);
or UO_207 (O_207,N_8655,N_9849);
or UO_208 (O_208,N_9088,N_8148);
and UO_209 (O_209,N_9091,N_9353);
and UO_210 (O_210,N_8059,N_9786);
nand UO_211 (O_211,N_8294,N_8384);
nor UO_212 (O_212,N_9017,N_9164);
nand UO_213 (O_213,N_9517,N_8763);
nor UO_214 (O_214,N_8998,N_9286);
or UO_215 (O_215,N_8567,N_9448);
nor UO_216 (O_216,N_9172,N_9670);
or UO_217 (O_217,N_9501,N_8120);
nand UO_218 (O_218,N_9004,N_8620);
nand UO_219 (O_219,N_8434,N_8513);
or UO_220 (O_220,N_8363,N_8674);
nor UO_221 (O_221,N_8911,N_9863);
and UO_222 (O_222,N_9176,N_9843);
or UO_223 (O_223,N_8400,N_8465);
or UO_224 (O_224,N_9446,N_9685);
and UO_225 (O_225,N_8133,N_9179);
nor UO_226 (O_226,N_8089,N_9113);
nor UO_227 (O_227,N_8473,N_8069);
nand UO_228 (O_228,N_8284,N_9470);
nand UO_229 (O_229,N_9521,N_9474);
and UO_230 (O_230,N_8010,N_9678);
or UO_231 (O_231,N_9230,N_8340);
or UO_232 (O_232,N_8016,N_9279);
or UO_233 (O_233,N_8106,N_8487);
nand UO_234 (O_234,N_9635,N_9236);
nand UO_235 (O_235,N_8318,N_9777);
nor UO_236 (O_236,N_9407,N_9370);
nor UO_237 (O_237,N_8161,N_8272);
or UO_238 (O_238,N_9323,N_8309);
nand UO_239 (O_239,N_9058,N_8132);
or UO_240 (O_240,N_8080,N_9941);
and UO_241 (O_241,N_9741,N_8729);
and UO_242 (O_242,N_8716,N_8860);
and UO_243 (O_243,N_8014,N_8524);
nand UO_244 (O_244,N_8234,N_9982);
and UO_245 (O_245,N_9570,N_8757);
nand UO_246 (O_246,N_9415,N_9300);
nand UO_247 (O_247,N_9856,N_9302);
nand UO_248 (O_248,N_8861,N_9770);
xor UO_249 (O_249,N_9464,N_8639);
nor UO_250 (O_250,N_8038,N_9458);
nor UO_251 (O_251,N_9343,N_9331);
or UO_252 (O_252,N_8591,N_8162);
or UO_253 (O_253,N_9332,N_8799);
nor UO_254 (O_254,N_8736,N_9417);
and UO_255 (O_255,N_8989,N_8755);
nor UO_256 (O_256,N_9372,N_9969);
or UO_257 (O_257,N_8052,N_8221);
nand UO_258 (O_258,N_9271,N_8545);
and UO_259 (O_259,N_9074,N_8993);
or UO_260 (O_260,N_9198,N_8606);
and UO_261 (O_261,N_9175,N_9944);
nand UO_262 (O_262,N_9897,N_8559);
or UO_263 (O_263,N_9580,N_8575);
nor UO_264 (O_264,N_9422,N_9465);
or UO_265 (O_265,N_9942,N_8624);
nor UO_266 (O_266,N_9022,N_8751);
nand UO_267 (O_267,N_8652,N_9976);
or UO_268 (O_268,N_8060,N_9833);
nor UO_269 (O_269,N_9224,N_9646);
and UO_270 (O_270,N_9698,N_9975);
nor UO_271 (O_271,N_9304,N_8068);
nand UO_272 (O_272,N_8165,N_9535);
nand UO_273 (O_273,N_9001,N_8241);
or UO_274 (O_274,N_9577,N_8982);
nor UO_275 (O_275,N_8756,N_8486);
or UO_276 (O_276,N_8433,N_9842);
nor UO_277 (O_277,N_9119,N_9250);
and UO_278 (O_278,N_9339,N_8159);
or UO_279 (O_279,N_8168,N_9710);
xnor UO_280 (O_280,N_8481,N_8179);
nand UO_281 (O_281,N_9055,N_9953);
nand UO_282 (O_282,N_8031,N_9605);
or UO_283 (O_283,N_8542,N_9730);
or UO_284 (O_284,N_9014,N_8875);
nor UO_285 (O_285,N_9769,N_9837);
nor UO_286 (O_286,N_9440,N_8499);
or UO_287 (O_287,N_9970,N_8181);
nand UO_288 (O_288,N_8201,N_8890);
nand UO_289 (O_289,N_9193,N_8858);
or UO_290 (O_290,N_9122,N_8087);
xnor UO_291 (O_291,N_9335,N_9964);
or UO_292 (O_292,N_8883,N_9028);
nand UO_293 (O_293,N_9971,N_8644);
nor UO_294 (O_294,N_9721,N_8171);
nor UO_295 (O_295,N_8215,N_9857);
nand UO_296 (O_296,N_9493,N_8681);
and UO_297 (O_297,N_8459,N_8637);
nor UO_298 (O_298,N_9924,N_9200);
nor UO_299 (O_299,N_9438,N_8186);
or UO_300 (O_300,N_8416,N_8372);
xor UO_301 (O_301,N_9728,N_9309);
or UO_302 (O_302,N_8849,N_8464);
and UO_303 (O_303,N_8738,N_8088);
nor UO_304 (O_304,N_8915,N_9135);
or UO_305 (O_305,N_9084,N_9273);
and UO_306 (O_306,N_8759,N_9738);
nor UO_307 (O_307,N_9348,N_9029);
and UO_308 (O_308,N_8402,N_8896);
or UO_309 (O_309,N_8985,N_8236);
or UO_310 (O_310,N_8645,N_8809);
nand UO_311 (O_311,N_9219,N_9822);
or UO_312 (O_312,N_9755,N_8676);
nor UO_313 (O_313,N_8174,N_9855);
and UO_314 (O_314,N_8784,N_9488);
or UO_315 (O_315,N_8086,N_8009);
and UO_316 (O_316,N_8718,N_9827);
or UO_317 (O_317,N_9447,N_9831);
and UO_318 (O_318,N_8914,N_9221);
or UO_319 (O_319,N_8741,N_9383);
nor UO_320 (O_320,N_8802,N_8417);
or UO_321 (O_321,N_9560,N_9939);
nor UO_322 (O_322,N_8205,N_8333);
or UO_323 (O_323,N_9943,N_8684);
nand UO_324 (O_324,N_8663,N_8766);
nor UO_325 (O_325,N_9979,N_8964);
or UO_326 (O_326,N_9542,N_8392);
nand UO_327 (O_327,N_9709,N_8817);
and UO_328 (O_328,N_9249,N_8908);
xor UO_329 (O_329,N_8062,N_9880);
and UO_330 (O_330,N_9579,N_9634);
or UO_331 (O_331,N_9437,N_8594);
nand UO_332 (O_332,N_9227,N_8220);
or UO_333 (O_333,N_9889,N_9497);
nor UO_334 (O_334,N_9647,N_8397);
or UO_335 (O_335,N_9760,N_9278);
or UO_336 (O_336,N_8163,N_9325);
nor UO_337 (O_337,N_9195,N_8852);
and UO_338 (O_338,N_9558,N_9997);
and UO_339 (O_339,N_9809,N_9457);
nor UO_340 (O_340,N_9643,N_9089);
or UO_341 (O_341,N_8141,N_8300);
nand UO_342 (O_342,N_9355,N_9967);
or UO_343 (O_343,N_8343,N_9114);
or UO_344 (O_344,N_9290,N_9033);
nor UO_345 (O_345,N_8156,N_8669);
nand UO_346 (O_346,N_9027,N_9805);
and UO_347 (O_347,N_9848,N_9099);
or UO_348 (O_348,N_8534,N_8983);
or UO_349 (O_349,N_8258,N_8940);
or UO_350 (O_350,N_8580,N_9608);
or UO_351 (O_351,N_9365,N_9823);
nand UO_352 (O_352,N_8360,N_8836);
nand UO_353 (O_353,N_8398,N_9295);
and UO_354 (O_354,N_9758,N_9485);
xnor UO_355 (O_355,N_9385,N_9702);
nand UO_356 (O_356,N_8346,N_9868);
nor UO_357 (O_357,N_9169,N_9773);
and UO_358 (O_358,N_9453,N_8152);
or UO_359 (O_359,N_8239,N_8414);
nor UO_360 (O_360,N_9452,N_9692);
or UO_361 (O_361,N_8871,N_9928);
nor UO_362 (O_362,N_9204,N_8722);
nand UO_363 (O_363,N_8475,N_9450);
or UO_364 (O_364,N_8178,N_8097);
nor UO_365 (O_365,N_9508,N_8453);
or UO_366 (O_366,N_9482,N_8491);
nor UO_367 (O_367,N_9281,N_9377);
nor UO_368 (O_368,N_9660,N_9075);
nor UO_369 (O_369,N_8747,N_8254);
and UO_370 (O_370,N_8913,N_9468);
and UO_371 (O_371,N_8893,N_8137);
or UO_372 (O_372,N_8648,N_8283);
nand UO_373 (O_373,N_8924,N_8981);
nor UO_374 (O_374,N_8692,N_9399);
and UO_375 (O_375,N_9202,N_9932);
nand UO_376 (O_376,N_9555,N_8586);
nor UO_377 (O_377,N_9413,N_8190);
nor UO_378 (O_378,N_8996,N_9649);
nor UO_379 (O_379,N_8151,N_9504);
xnor UO_380 (O_380,N_8328,N_9704);
nor UO_381 (O_381,N_9199,N_8571);
nor UO_382 (O_382,N_9259,N_9336);
nor UO_383 (O_383,N_8719,N_8562);
and UO_384 (O_384,N_8945,N_8138);
and UO_385 (O_385,N_8131,N_8734);
or UO_386 (O_386,N_9442,N_9143);
or UO_387 (O_387,N_8551,N_8404);
xor UO_388 (O_388,N_8440,N_9750);
nor UO_389 (O_389,N_9053,N_8588);
nand UO_390 (O_390,N_8378,N_8394);
nor UO_391 (O_391,N_9851,N_8028);
nor UO_392 (O_392,N_9187,N_9487);
or UO_393 (O_393,N_9991,N_9321);
nor UO_394 (O_394,N_8844,N_9588);
nand UO_395 (O_395,N_9190,N_8117);
nor UO_396 (O_396,N_8093,N_8257);
xnor UO_397 (O_397,N_8828,N_8472);
and UO_398 (O_398,N_9907,N_9373);
or UO_399 (O_399,N_8967,N_8785);
nor UO_400 (O_400,N_8685,N_9334);
nand UO_401 (O_401,N_9623,N_8846);
nand UO_402 (O_402,N_8348,N_8715);
or UO_403 (O_403,N_9796,N_8339);
nand UO_404 (O_404,N_8390,N_8720);
nor UO_405 (O_405,N_8647,N_8356);
and UO_406 (O_406,N_8422,N_8005);
and UO_407 (O_407,N_9461,N_9726);
nand UO_408 (O_408,N_9478,N_9500);
or UO_409 (O_409,N_8382,N_9963);
and UO_410 (O_410,N_8565,N_9039);
and UO_411 (O_411,N_9009,N_8202);
or UO_412 (O_412,N_8177,N_9671);
nor UO_413 (O_413,N_9751,N_8856);
nor UO_414 (O_414,N_9048,N_8301);
and UO_415 (O_415,N_9059,N_9467);
and UO_416 (O_416,N_9723,N_9617);
nor UO_417 (O_417,N_8548,N_8296);
or UO_418 (O_418,N_9311,N_8332);
nand UO_419 (O_419,N_9632,N_9664);
nor UO_420 (O_420,N_9060,N_9123);
nand UO_421 (O_421,N_9626,N_8002);
nor UO_422 (O_422,N_8845,N_9929);
nor UO_423 (O_423,N_8493,N_8347);
or UO_424 (O_424,N_8798,N_9846);
nand UO_425 (O_425,N_9567,N_9511);
and UO_426 (O_426,N_9024,N_9451);
nand UO_427 (O_427,N_9265,N_8745);
and UO_428 (O_428,N_9638,N_9231);
and UO_429 (O_429,N_8825,N_8773);
and UO_430 (O_430,N_8266,N_9518);
or UO_431 (O_431,N_8659,N_8721);
nand UO_432 (O_432,N_8048,N_9393);
nand UO_433 (O_433,N_9080,N_8047);
or UO_434 (O_434,N_8728,N_9118);
and UO_435 (O_435,N_9688,N_9037);
and UO_436 (O_436,N_8725,N_8259);
nand UO_437 (O_437,N_9881,N_8780);
and UO_438 (O_438,N_9593,N_8772);
nand UO_439 (O_439,N_8480,N_8577);
nor UO_440 (O_440,N_9829,N_9032);
nor UO_441 (O_441,N_9432,N_8144);
or UO_442 (O_442,N_8600,N_9589);
nor UO_443 (O_443,N_9962,N_9584);
or UO_444 (O_444,N_9705,N_9502);
or UO_445 (O_445,N_8851,N_8643);
nor UO_446 (O_446,N_8555,N_9919);
nand UO_447 (O_447,N_9463,N_8813);
and UO_448 (O_448,N_9367,N_9046);
or UO_449 (O_449,N_8876,N_8275);
nand UO_450 (O_450,N_8602,N_9661);
and UO_451 (O_451,N_8023,N_8095);
or UO_452 (O_452,N_8768,N_9269);
and UO_453 (O_453,N_9072,N_8812);
or UO_454 (O_454,N_8810,N_8041);
nand UO_455 (O_455,N_8727,N_9403);
nor UO_456 (O_456,N_8295,N_8198);
and UO_457 (O_457,N_9877,N_9120);
or UO_458 (O_458,N_9107,N_9966);
nor UO_459 (O_459,N_9804,N_9289);
or UO_460 (O_460,N_8176,N_8704);
nor UO_461 (O_461,N_9318,N_9132);
or UO_462 (O_462,N_8322,N_9677);
or UO_463 (O_463,N_9063,N_9819);
or UO_464 (O_464,N_8185,N_9170);
nand UO_465 (O_465,N_9350,N_9731);
or UO_466 (O_466,N_9266,N_8240);
or UO_467 (O_467,N_8281,N_8114);
and UO_468 (O_468,N_8359,N_8344);
nand UO_469 (O_469,N_8839,N_8820);
nand UO_470 (O_470,N_8456,N_9225);
nand UO_471 (O_471,N_9392,N_8211);
nand UO_472 (O_472,N_8642,N_8935);
nor UO_473 (O_473,N_9142,N_8351);
xnor UO_474 (O_474,N_8064,N_9689);
nor UO_475 (O_475,N_9040,N_9310);
xor UO_476 (O_476,N_8975,N_8032);
or UO_477 (O_477,N_9946,N_9042);
and UO_478 (O_478,N_9708,N_8497);
or UO_479 (O_479,N_9947,N_8918);
or UO_480 (O_480,N_8694,N_9716);
or UO_481 (O_481,N_9785,N_9216);
nor UO_482 (O_482,N_8695,N_8075);
and UO_483 (O_483,N_8092,N_8107);
nand UO_484 (O_484,N_9637,N_8966);
nand UO_485 (O_485,N_9499,N_9338);
or UO_486 (O_486,N_9382,N_8135);
and UO_487 (O_487,N_9581,N_9808);
nor UO_488 (O_488,N_8420,N_8355);
or UO_489 (O_489,N_8498,N_8249);
nand UO_490 (O_490,N_9630,N_9106);
or UO_491 (O_491,N_9414,N_9902);
and UO_492 (O_492,N_9476,N_8553);
and UO_493 (O_493,N_9360,N_8428);
nor UO_494 (O_494,N_9391,N_8595);
and UO_495 (O_495,N_8614,N_9358);
nand UO_496 (O_496,N_8572,N_9354);
or UO_497 (O_497,N_8105,N_9427);
and UO_498 (O_498,N_8748,N_9812);
or UO_499 (O_499,N_8954,N_9208);
and UO_500 (O_500,N_8833,N_8556);
and UO_501 (O_501,N_8790,N_9696);
or UO_502 (O_502,N_9679,N_8955);
nor UO_503 (O_503,N_9171,N_9620);
nand UO_504 (O_504,N_8977,N_9247);
nand UO_505 (O_505,N_8279,N_9357);
nand UO_506 (O_506,N_8214,N_8880);
nor UO_507 (O_507,N_9754,N_8317);
and UO_508 (O_508,N_9174,N_9861);
nor UO_509 (O_509,N_9421,N_9815);
nor UO_510 (O_510,N_9530,N_9906);
or UO_511 (O_511,N_8262,N_9161);
nor UO_512 (O_512,N_8671,N_8101);
and UO_513 (O_513,N_9772,N_9801);
nand UO_514 (O_514,N_9329,N_9085);
or UO_515 (O_515,N_9270,N_8519);
nand UO_516 (O_516,N_8192,N_8910);
nor UO_517 (O_517,N_9388,N_9840);
and UO_518 (O_518,N_8050,N_9695);
and UO_519 (O_519,N_9019,N_9347);
nor UO_520 (O_520,N_9878,N_9747);
nor UO_521 (O_521,N_8576,N_8113);
or UO_522 (O_522,N_9194,N_9425);
and UO_523 (O_523,N_9374,N_9663);
or UO_524 (O_524,N_9999,N_8145);
nor UO_525 (O_525,N_8484,N_8570);
or UO_526 (O_526,N_8501,N_8026);
or UO_527 (O_527,N_9241,N_9489);
nand UO_528 (O_528,N_9800,N_8342);
nor UO_529 (O_529,N_8869,N_9867);
nand UO_530 (O_530,N_9952,N_8587);
xnor UO_531 (O_531,N_8898,N_8953);
or UO_532 (O_532,N_8449,N_8460);
and UO_533 (O_533,N_9327,N_9955);
and UO_534 (O_534,N_9995,N_8122);
and UO_535 (O_535,N_9301,N_8371);
nand UO_536 (O_536,N_8219,N_9763);
nor UO_537 (O_537,N_8706,N_8925);
nand UO_538 (O_538,N_8646,N_8022);
nand UO_539 (O_539,N_9883,N_9859);
nand UO_540 (O_540,N_8818,N_9587);
and UO_541 (O_541,N_8316,N_8270);
or UO_542 (O_542,N_9697,N_8293);
nor UO_543 (O_543,N_8329,N_9361);
and UO_544 (O_544,N_9070,N_8528);
nand UO_545 (O_545,N_9562,N_9539);
or UO_546 (O_546,N_8832,N_8677);
nor UO_547 (O_547,N_8466,N_9031);
and UO_548 (O_548,N_9739,N_9386);
nor UO_549 (O_549,N_9583,N_9126);
and UO_550 (O_550,N_9835,N_9349);
or UO_551 (O_551,N_8121,N_9669);
nor UO_552 (O_552,N_8083,N_8709);
and UO_553 (O_553,N_9000,N_9192);
or UO_554 (O_554,N_8054,N_9087);
nor UO_555 (O_555,N_8321,N_8445);
nand UO_556 (O_556,N_8617,N_9744);
nor UO_557 (O_557,N_8410,N_9672);
nand UO_558 (O_558,N_8888,N_8479);
or UO_559 (O_559,N_9475,N_9506);
and UO_560 (O_560,N_8968,N_9543);
and UO_561 (O_561,N_8909,N_9949);
nand UO_562 (O_562,N_9083,N_9418);
nor UO_563 (O_563,N_9155,N_8130);
and UO_564 (O_564,N_8438,N_9484);
nor UO_565 (O_565,N_9572,N_8700);
nand UO_566 (O_566,N_9563,N_9860);
or UO_567 (O_567,N_9749,N_8605);
xnor UO_568 (O_568,N_8783,N_8862);
or UO_569 (O_569,N_8905,N_9152);
nand UO_570 (O_570,N_8838,N_9134);
nand UO_571 (O_571,N_8061,N_9056);
and UO_572 (O_572,N_9793,N_9268);
and UO_573 (O_573,N_8452,N_8338);
nor UO_574 (O_574,N_9853,N_9915);
and UO_575 (O_575,N_8961,N_8919);
nand UO_576 (O_576,N_8815,N_8389);
and UO_577 (O_577,N_8530,N_9291);
and UO_578 (O_578,N_9168,N_8774);
nor UO_579 (O_579,N_9736,N_8859);
xnor UO_580 (O_580,N_8821,N_8902);
and UO_581 (O_581,N_9435,N_9612);
nand UO_582 (O_582,N_9294,N_8243);
nor UO_583 (O_583,N_8391,N_9707);
and UO_584 (O_584,N_9871,N_8482);
and UO_585 (O_585,N_8786,N_8286);
nor UO_586 (O_586,N_8269,N_8502);
and UO_587 (O_587,N_8863,N_9020);
and UO_588 (O_588,N_9036,N_8675);
nand UO_589 (O_589,N_9197,N_8752);
and UO_590 (O_590,N_9111,N_8376);
and UO_591 (O_591,N_9609,N_9996);
or UO_592 (O_592,N_8885,N_9886);
nor UO_593 (O_593,N_9255,N_9057);
nor UO_594 (O_594,N_9650,N_9503);
or UO_595 (O_595,N_8303,N_9345);
or UO_596 (O_596,N_9742,N_8634);
or UO_597 (O_597,N_9601,N_8533);
nor UO_598 (O_598,N_8366,N_9406);
nand UO_599 (O_599,N_8462,N_8442);
or UO_600 (O_600,N_8653,N_9858);
nor UO_601 (O_601,N_9621,N_9462);
nor UO_602 (O_602,N_8494,N_8826);
nor UO_603 (O_603,N_8717,N_9012);
nand UO_604 (O_604,N_9526,N_9802);
or UO_605 (O_605,N_9892,N_9090);
nand UO_606 (O_606,N_9233,N_9916);
and UO_607 (O_607,N_9434,N_8808);
nor UO_608 (O_608,N_9622,N_8699);
nand UO_609 (O_609,N_8067,N_8496);
nand UO_610 (O_610,N_9376,N_9363);
and UO_611 (O_611,N_8662,N_8230);
nor UO_612 (O_612,N_9430,N_8331);
nor UO_613 (O_613,N_8251,N_9724);
nor UO_614 (O_614,N_8879,N_9875);
or UO_615 (O_615,N_9337,N_9912);
nor UO_616 (O_616,N_8248,N_8001);
or UO_617 (O_617,N_8568,N_8769);
and UO_618 (O_618,N_9459,N_8585);
or UO_619 (O_619,N_8090,N_9315);
nand UO_620 (O_620,N_8703,N_9874);
nor UO_621 (O_621,N_8760,N_8724);
nor UO_622 (O_622,N_9479,N_9703);
or UO_623 (O_623,N_8226,N_8708);
or UO_624 (O_624,N_8247,N_9223);
nor UO_625 (O_625,N_9911,N_9185);
nor UO_626 (O_626,N_9429,N_8952);
nand UO_627 (O_627,N_8654,N_8477);
and UO_628 (O_628,N_8109,N_8084);
or UO_629 (O_629,N_9956,N_9794);
or UO_630 (O_630,N_8173,N_8950);
and UO_631 (O_631,N_8238,N_8776);
and UO_632 (O_632,N_8668,N_9680);
and UO_633 (O_633,N_9507,N_9673);
or UO_634 (O_634,N_9234,N_8974);
or UO_635 (O_635,N_8444,N_8960);
or UO_636 (O_636,N_9067,N_8801);
xnor UO_637 (O_637,N_8610,N_9516);
nor UO_638 (O_638,N_8383,N_8274);
nor UO_639 (O_639,N_9207,N_9984);
or UO_640 (O_640,N_9597,N_8933);
and UO_641 (O_641,N_8413,N_8829);
xnor UO_642 (O_642,N_9765,N_8742);
or UO_643 (O_643,N_9030,N_8907);
nand UO_644 (O_644,N_8285,N_9151);
and UO_645 (O_645,N_9652,N_9784);
or UO_646 (O_646,N_8629,N_8635);
and UO_647 (O_647,N_9333,N_9307);
nor UO_648 (O_648,N_9158,N_9277);
and UO_649 (O_649,N_9803,N_8670);
nor UO_650 (O_650,N_9094,N_9729);
nand UO_651 (O_651,N_8690,N_9910);
and UO_652 (O_652,N_9662,N_9287);
nor UO_653 (O_653,N_8012,N_8311);
and UO_654 (O_654,N_8129,N_9814);
nand UO_655 (O_655,N_8051,N_8319);
or UO_656 (O_656,N_9687,N_9314);
nor UO_657 (O_657,N_8944,N_8560);
nand UO_658 (O_658,N_9798,N_9364);
nand UO_659 (O_659,N_9069,N_8927);
nand UO_660 (O_660,N_8621,N_9935);
and UO_661 (O_661,N_9328,N_8521);
and UO_662 (O_662,N_9885,N_9205);
nor UO_663 (O_663,N_9016,N_8103);
nand UO_664 (O_664,N_9163,N_8782);
nand UO_665 (O_665,N_8959,N_9614);
or UO_666 (O_666,N_9191,N_8827);
nor UO_667 (O_667,N_9904,N_8426);
nor UO_668 (O_668,N_9433,N_9748);
and UO_669 (O_669,N_9817,N_8325);
nand UO_670 (O_670,N_8246,N_9285);
xnor UO_671 (O_671,N_8696,N_8423);
and UO_672 (O_672,N_9054,N_9778);
and UO_673 (O_673,N_8252,N_8349);
or UO_674 (O_674,N_9436,N_8870);
or UO_675 (O_675,N_8379,N_9303);
nand UO_676 (O_676,N_9398,N_9576);
nand UO_677 (O_677,N_8310,N_9590);
or UO_678 (O_678,N_8374,N_9900);
nor UO_679 (O_679,N_9242,N_9389);
and UO_680 (O_680,N_8789,N_8550);
nand UO_681 (O_681,N_9574,N_8740);
nand UO_682 (O_682,N_8538,N_9010);
or UO_683 (O_683,N_8264,N_8866);
nor UO_684 (O_684,N_9378,N_9184);
nor UO_685 (O_685,N_9693,N_9699);
or UO_686 (O_686,N_8350,N_8749);
nor UO_687 (O_687,N_9466,N_9894);
and UO_688 (O_688,N_8094,N_9346);
and UO_689 (O_689,N_9718,N_8507);
nand UO_690 (O_690,N_8723,N_8223);
nor UO_691 (O_691,N_8771,N_9264);
nor UO_692 (O_692,N_9177,N_8997);
nor UO_693 (O_693,N_8313,N_8203);
and UO_694 (O_694,N_8157,N_8271);
nor UO_695 (O_695,N_8758,N_8081);
xnor UO_696 (O_696,N_8912,N_9553);
or UO_697 (O_697,N_8540,N_9810);
nor UO_698 (O_698,N_8446,N_8419);
and UO_699 (O_699,N_9896,N_8666);
nor UO_700 (O_700,N_9961,N_8948);
nand UO_701 (O_701,N_8123,N_9537);
and UO_702 (O_702,N_9713,N_8381);
nand UO_703 (O_703,N_9791,N_9419);
nand UO_704 (O_704,N_9619,N_8451);
nand UO_705 (O_705,N_9901,N_9735);
nor UO_706 (O_706,N_9905,N_9657);
nand UO_707 (O_707,N_8034,N_9544);
xor UO_708 (O_708,N_9974,N_8352);
nor UO_709 (O_709,N_8292,N_8797);
or UO_710 (O_710,N_8916,N_8536);
nor UO_711 (O_711,N_9933,N_8057);
and UO_712 (O_712,N_8976,N_8065);
nand UO_713 (O_713,N_8489,N_9986);
and UO_714 (O_714,N_9051,N_8714);
or UO_715 (O_715,N_9262,N_8775);
and UO_716 (O_716,N_9734,N_8124);
nor UO_717 (O_717,N_8504,N_8018);
and UO_718 (O_718,N_8712,N_9887);
and UO_719 (O_719,N_9305,N_8204);
nand UO_720 (O_720,N_9884,N_8791);
nor UO_721 (O_721,N_8070,N_8767);
or UO_722 (O_722,N_9439,N_9564);
nand UO_723 (O_723,N_9480,N_9260);
or UO_724 (O_724,N_8375,N_8013);
nand UO_725 (O_725,N_9201,N_9081);
nor UO_726 (O_726,N_8011,N_9639);
and UO_727 (O_727,N_9752,N_9681);
nor UO_728 (O_728,N_9642,N_9850);
or UO_729 (O_729,N_8256,N_9989);
and UO_730 (O_730,N_9653,N_9715);
and UO_731 (O_731,N_8395,N_9927);
nor UO_732 (O_732,N_9536,N_9410);
or UO_733 (O_733,N_9957,N_8578);
and UO_734 (O_734,N_8922,N_8187);
nor UO_735 (O_735,N_8835,N_8612);
and UO_736 (O_736,N_9239,N_8972);
or UO_737 (O_737,N_8926,N_9554);
or UO_738 (O_738,N_8777,N_9188);
nor UO_739 (O_739,N_9675,N_8315);
nor UO_740 (O_740,N_9068,N_8541);
and UO_741 (O_741,N_9342,N_8564);
or UO_742 (O_742,N_8638,N_8664);
or UO_743 (O_743,N_8140,N_8458);
nor UO_744 (O_744,N_9781,N_8889);
and UO_745 (O_745,N_8206,N_9604);
nor UO_746 (O_746,N_8345,N_8461);
nand UO_747 (O_747,N_8796,N_9561);
nand UO_748 (O_748,N_9390,N_8225);
or UO_749 (O_749,N_8505,N_9914);
nand UO_750 (O_750,N_8881,N_8969);
and UO_751 (O_751,N_8920,N_9293);
nor UO_752 (O_752,N_9362,N_8134);
and UO_753 (O_753,N_9101,N_8503);
nand UO_754 (O_754,N_9396,N_8208);
nor UO_755 (O_755,N_9844,N_9138);
or UO_756 (O_756,N_8743,N_8195);
and UO_757 (O_757,N_9783,N_9676);
nor UO_758 (O_758,N_9683,N_9312);
and UO_759 (O_759,N_9183,N_8649);
and UO_760 (O_760,N_9041,N_8324);
nand UO_761 (O_761,N_9431,N_8850);
nand UO_762 (O_762,N_9549,N_8036);
and UO_763 (O_763,N_9565,N_8019);
and UO_764 (O_764,N_9387,N_9585);
and UO_765 (O_765,N_9541,N_9725);
and UO_766 (O_766,N_8855,N_8099);
or UO_767 (O_767,N_8085,N_9523);
and UO_768 (O_768,N_9062,N_9891);
nand UO_769 (O_769,N_8153,N_8142);
nor UO_770 (O_770,N_9610,N_8155);
nand UO_771 (O_771,N_9441,N_9127);
or UO_772 (O_772,N_8864,N_8500);
and UO_773 (O_773,N_8962,N_9153);
nand UO_774 (O_774,N_9926,N_8224);
and UO_775 (O_775,N_8963,N_9575);
nor UO_776 (O_776,N_8762,N_9005);
nor UO_777 (O_777,N_8115,N_9211);
and UO_778 (O_778,N_9636,N_8609);
nand UO_779 (O_779,N_9245,N_8711);
nor UO_780 (O_780,N_9668,N_9160);
or UO_781 (O_781,N_9073,N_9568);
and UO_782 (O_782,N_8713,N_8242);
nand UO_783 (O_783,N_9682,N_8608);
and UO_784 (O_784,N_9559,N_8432);
nor UO_785 (O_785,N_9694,N_8388);
and UO_786 (O_786,N_8096,N_8868);
and UO_787 (O_787,N_9298,N_9981);
nand UO_788 (O_788,N_8598,N_9103);
and UO_789 (O_789,N_8937,N_9512);
and UO_790 (O_790,N_8822,N_9248);
or UO_791 (O_791,N_8327,N_9044);
or UO_792 (O_792,N_8025,N_9780);
nor UO_793 (O_793,N_9326,N_8622);
or UO_794 (O_794,N_8164,N_9226);
or UO_795 (O_795,N_8197,N_9078);
nand UO_796 (O_796,N_9108,N_8058);
nor UO_797 (O_797,N_8222,N_9299);
nand UO_798 (O_798,N_8707,N_9093);
nor UO_799 (O_799,N_9105,N_8792);
nand UO_800 (O_800,N_8210,N_9359);
and UO_801 (O_801,N_9792,N_8939);
and UO_802 (O_802,N_9313,N_8158);
nand UO_803 (O_803,N_8509,N_8616);
nor UO_804 (O_804,N_8593,N_8063);
nor UO_805 (O_805,N_8750,N_8406);
nand UO_806 (O_806,N_9013,N_9116);
or UO_807 (O_807,N_9428,N_9775);
nand UO_808 (O_808,N_8468,N_8867);
xor UO_809 (O_809,N_9007,N_8607);
and UO_810 (O_810,N_9455,N_9243);
or UO_811 (O_811,N_9951,N_8518);
and UO_812 (O_812,N_8021,N_9994);
nand UO_813 (O_813,N_8017,N_9648);
xnor UO_814 (O_814,N_9538,N_8999);
nand UO_815 (O_815,N_8079,N_9893);
nand UO_816 (O_816,N_8020,N_9545);
nand UO_817 (O_817,N_8710,N_9405);
nor UO_818 (O_818,N_9895,N_8517);
nor UO_819 (O_819,N_9519,N_9034);
nand UO_820 (O_820,N_8547,N_8035);
and UO_821 (O_821,N_8447,N_8299);
or UO_822 (O_822,N_8901,N_8986);
nand UO_823 (O_823,N_8369,N_8184);
and UO_824 (O_824,N_9873,N_9025);
nor UO_825 (O_825,N_9181,N_9714);
nor UO_826 (O_826,N_9882,N_9613);
or UO_827 (O_827,N_9352,N_8819);
or UO_828 (O_828,N_8516,N_8628);
or UO_829 (O_829,N_8857,N_8554);
or UO_830 (O_830,N_8697,N_8894);
nor UO_831 (O_831,N_8735,N_8613);
or UO_832 (O_832,N_8263,N_9210);
and UO_833 (O_833,N_8837,N_8421);
nand UO_834 (O_834,N_8842,N_8847);
nor UO_835 (O_835,N_8744,N_9909);
and UO_836 (O_836,N_9237,N_9443);
nor UO_837 (O_837,N_9026,N_8623);
or UO_838 (O_838,N_8015,N_8160);
and UO_839 (O_839,N_8277,N_9018);
or UO_840 (O_840,N_9035,N_9811);
or UO_841 (O_841,N_9615,N_9571);
or UO_842 (O_842,N_8098,N_8582);
nor UO_843 (O_843,N_8705,N_9086);
nor UO_844 (O_844,N_9214,N_8055);
nand UO_845 (O_845,N_9920,N_8561);
or UO_846 (O_846,N_8199,N_8698);
or UO_847 (O_847,N_8003,N_9958);
xnor UO_848 (O_848,N_9522,N_9771);
nand UO_849 (O_849,N_9240,N_9145);
and UO_850 (O_850,N_8287,N_9368);
nor UO_851 (O_851,N_9761,N_8188);
xnor UO_852 (O_852,N_9821,N_9582);
xor UO_853 (O_853,N_9606,N_8794);
and UO_854 (O_854,N_8625,N_9782);
nand UO_855 (O_855,N_8604,N_8934);
nand UO_856 (O_856,N_9640,N_8091);
nand UO_857 (O_857,N_9625,N_9256);
nor UO_858 (O_858,N_8877,N_9547);
or UO_859 (O_859,N_8947,N_9978);
nor UO_860 (O_860,N_8995,N_8592);
or UO_861 (O_861,N_9686,N_9047);
nand UO_862 (O_862,N_8965,N_8368);
nand UO_863 (O_863,N_9656,N_8110);
or UO_864 (O_864,N_9505,N_8800);
and UO_865 (O_865,N_8298,N_8683);
or UO_866 (O_866,N_8957,N_8341);
nand UO_867 (O_867,N_8189,N_8370);
nor UO_868 (O_868,N_9109,N_8958);
or UO_869 (O_869,N_9490,N_9065);
nor UO_870 (O_870,N_9492,N_8841);
nand UO_871 (O_871,N_8073,N_9146);
nor UO_872 (O_872,N_8834,N_8046);
nor UO_873 (O_873,N_9654,N_8830);
nor UO_874 (O_874,N_9990,N_9306);
or UO_875 (O_875,N_9566,N_9411);
and UO_876 (O_876,N_8401,N_9263);
nand UO_877 (O_877,N_9691,N_8512);
nand UO_878 (O_878,N_9102,N_8441);
or UO_879 (O_879,N_8291,N_8897);
nand UO_880 (O_880,N_8250,N_9420);
nor UO_881 (O_881,N_8147,N_8314);
and UO_882 (O_882,N_9015,N_9931);
xnor UO_883 (O_883,N_9573,N_9154);
nand UO_884 (O_884,N_8354,N_8778);
and UO_885 (O_885,N_9776,N_9816);
or UO_886 (O_886,N_9985,N_9021);
nor UO_887 (O_887,N_9528,N_9925);
nand UO_888 (O_888,N_9586,N_8439);
or UO_889 (O_889,N_9789,N_8687);
and UO_890 (O_890,N_8873,N_8640);
nor UO_891 (O_891,N_8865,N_8149);
or UO_892 (O_892,N_8150,N_8529);
or UO_893 (O_893,N_9206,N_9711);
nor UO_894 (O_894,N_9292,N_9272);
or UO_895 (O_895,N_9854,N_9767);
and UO_896 (O_896,N_9471,N_8074);
nor UO_897 (O_897,N_8474,N_9594);
nor UO_898 (O_898,N_8407,N_8100);
or UO_899 (O_899,N_9397,N_9820);
nor UO_900 (O_900,N_8405,N_8072);
and UO_901 (O_901,N_9253,N_8172);
nand UO_902 (O_902,N_9209,N_9727);
nor UO_903 (O_903,N_8537,N_8362);
nand UO_904 (O_904,N_9076,N_8127);
nor UO_905 (O_905,N_9569,N_9096);
nor UO_906 (O_906,N_9473,N_9380);
nand UO_907 (O_907,N_8111,N_9665);
nor UO_908 (O_908,N_8535,N_8532);
nand UO_909 (O_909,N_8418,N_8488);
nand UO_910 (O_910,N_8581,N_8218);
and UO_911 (O_911,N_8066,N_9460);
and UO_912 (O_912,N_9992,N_9316);
nand UO_913 (O_913,N_9049,N_8941);
nand UO_914 (O_914,N_9862,N_8702);
nor UO_915 (O_915,N_8377,N_9684);
and UO_916 (O_916,N_8658,N_8882);
or UO_917 (O_917,N_9611,N_9658);
and UO_918 (O_918,N_9618,N_8312);
nor UO_919 (O_919,N_9828,N_8180);
and UO_920 (O_920,N_8104,N_8928);
nor UO_921 (O_921,N_9838,N_8288);
nand UO_922 (O_922,N_9960,N_9945);
and UO_923 (O_923,N_8788,N_8193);
nor UO_924 (O_924,N_8334,N_8191);
or UO_925 (O_925,N_9423,N_8323);
nand UO_926 (O_926,N_9133,N_9416);
nor UO_927 (O_927,N_9196,N_8118);
xnor UO_928 (O_928,N_9757,N_9525);
and UO_929 (O_929,N_8231,N_9940);
nand UO_930 (O_930,N_8307,N_9674);
nand UO_931 (O_931,N_8906,N_8126);
or UO_932 (O_932,N_8425,N_8626);
or UO_933 (O_933,N_8454,N_8082);
nor UO_934 (O_934,N_9409,N_8979);
nor UO_935 (O_935,N_8731,N_8730);
nand UO_936 (O_936,N_8984,N_8754);
or UO_937 (O_937,N_8596,N_9813);
and UO_938 (O_938,N_8077,N_9064);
and UO_939 (O_939,N_8136,N_8078);
or UO_940 (O_940,N_8267,N_9533);
nor UO_941 (O_941,N_9629,N_9531);
nand UO_942 (O_942,N_9121,N_8361);
xor UO_943 (O_943,N_9097,N_9130);
nor UO_944 (O_944,N_8770,N_9807);
nand UO_945 (O_945,N_9456,N_9400);
nor UO_946 (O_946,N_8273,N_9556);
or UO_947 (O_947,N_8412,N_9998);
and UO_948 (O_948,N_9218,N_9852);
nor UO_949 (O_949,N_9720,N_9222);
nand UO_950 (O_950,N_8045,N_8429);
nor UO_951 (O_951,N_8650,N_8033);
and UO_952 (O_952,N_8170,N_8840);
xor UO_953 (O_953,N_8380,N_8229);
and UO_954 (O_954,N_9515,N_9491);
xnor UO_955 (O_955,N_9921,N_9481);
or UO_956 (O_956,N_8970,N_9607);
or UO_957 (O_957,N_8514,N_9008);
or UO_958 (O_958,N_8443,N_8892);
nor UO_959 (O_959,N_8039,N_8305);
and UO_960 (O_960,N_8994,N_9644);
or UO_961 (O_961,N_9832,N_9150);
nor UO_962 (O_962,N_8450,N_8691);
nor UO_963 (O_963,N_8200,N_8884);
or UO_964 (O_964,N_8183,N_8990);
and UO_965 (O_965,N_9495,N_9712);
and UO_966 (O_966,N_8753,N_9872);
or UO_967 (O_967,N_8007,N_8260);
nor UO_968 (O_968,N_9246,N_8358);
nor UO_969 (O_969,N_8000,N_9147);
or UO_970 (O_970,N_8543,N_8667);
nand UO_971 (O_971,N_8732,N_9917);
and UO_972 (O_972,N_9098,N_9494);
or UO_973 (O_973,N_9092,N_8049);
nor UO_974 (O_974,N_9936,N_9865);
nor UO_975 (O_975,N_9824,N_8467);
nor UO_976 (O_976,N_8435,N_8336);
and UO_977 (O_977,N_8680,N_9426);
nand UO_978 (O_978,N_8483,N_9212);
nand UO_979 (O_979,N_8337,N_8563);
nor UO_980 (O_980,N_8656,N_8030);
nor UO_981 (O_981,N_9825,N_9779);
nor UO_982 (O_982,N_8212,N_8627);
nor UO_983 (O_983,N_9870,N_8805);
nor UO_984 (O_984,N_8992,N_8599);
nor UO_985 (O_985,N_8232,N_8804);
nand UO_986 (O_986,N_9404,N_9401);
nor UO_987 (O_987,N_8330,N_9520);
or UO_988 (O_988,N_8678,N_8385);
nor UO_989 (O_989,N_8373,N_9182);
or UO_990 (O_990,N_8282,N_9641);
nor UO_991 (O_991,N_9203,N_9082);
nor UO_992 (O_992,N_8297,N_9006);
or UO_993 (O_993,N_8522,N_8527);
nor UO_994 (O_994,N_8209,N_9903);
nor UO_995 (O_995,N_8943,N_9324);
or UO_996 (O_996,N_8245,N_8895);
and UO_997 (O_997,N_8166,N_9112);
nand UO_998 (O_998,N_8396,N_8213);
nand UO_999 (O_999,N_9394,N_8630);
nand UO_1000 (O_1000,N_8208,N_9657);
nor UO_1001 (O_1001,N_8794,N_8623);
nor UO_1002 (O_1002,N_8477,N_8531);
and UO_1003 (O_1003,N_9262,N_9197);
and UO_1004 (O_1004,N_8005,N_9255);
and UO_1005 (O_1005,N_8539,N_9919);
and UO_1006 (O_1006,N_9106,N_9906);
nand UO_1007 (O_1007,N_9608,N_8230);
nor UO_1008 (O_1008,N_9760,N_9106);
or UO_1009 (O_1009,N_8887,N_9594);
or UO_1010 (O_1010,N_9435,N_8970);
nand UO_1011 (O_1011,N_9718,N_8240);
and UO_1012 (O_1012,N_8793,N_9177);
nand UO_1013 (O_1013,N_9605,N_8163);
or UO_1014 (O_1014,N_9520,N_9779);
and UO_1015 (O_1015,N_8525,N_9460);
or UO_1016 (O_1016,N_9617,N_8261);
nand UO_1017 (O_1017,N_9085,N_9587);
nand UO_1018 (O_1018,N_8386,N_9520);
or UO_1019 (O_1019,N_9297,N_9968);
nor UO_1020 (O_1020,N_8201,N_9216);
nand UO_1021 (O_1021,N_8340,N_8406);
nor UO_1022 (O_1022,N_9559,N_8163);
nand UO_1023 (O_1023,N_8888,N_9068);
or UO_1024 (O_1024,N_8765,N_9034);
or UO_1025 (O_1025,N_9533,N_9446);
nor UO_1026 (O_1026,N_8039,N_9295);
or UO_1027 (O_1027,N_9684,N_8064);
and UO_1028 (O_1028,N_8441,N_9176);
nand UO_1029 (O_1029,N_8561,N_8601);
nor UO_1030 (O_1030,N_8922,N_9749);
or UO_1031 (O_1031,N_9336,N_9389);
and UO_1032 (O_1032,N_8271,N_9187);
or UO_1033 (O_1033,N_9854,N_8324);
or UO_1034 (O_1034,N_8460,N_9213);
nand UO_1035 (O_1035,N_8348,N_9311);
nor UO_1036 (O_1036,N_8711,N_9036);
or UO_1037 (O_1037,N_9380,N_9004);
nor UO_1038 (O_1038,N_9449,N_8287);
and UO_1039 (O_1039,N_8019,N_8807);
and UO_1040 (O_1040,N_9025,N_8019);
and UO_1041 (O_1041,N_8626,N_9078);
and UO_1042 (O_1042,N_9709,N_8666);
and UO_1043 (O_1043,N_8033,N_9199);
nand UO_1044 (O_1044,N_9283,N_8455);
xor UO_1045 (O_1045,N_9162,N_9481);
or UO_1046 (O_1046,N_9584,N_9256);
nand UO_1047 (O_1047,N_8888,N_8317);
or UO_1048 (O_1048,N_9613,N_9329);
or UO_1049 (O_1049,N_8286,N_8209);
nor UO_1050 (O_1050,N_9203,N_8294);
and UO_1051 (O_1051,N_8788,N_8359);
nor UO_1052 (O_1052,N_9116,N_9242);
nand UO_1053 (O_1053,N_9620,N_9574);
nor UO_1054 (O_1054,N_9805,N_8601);
xnor UO_1055 (O_1055,N_9427,N_9310);
nor UO_1056 (O_1056,N_9795,N_9641);
and UO_1057 (O_1057,N_8921,N_9889);
and UO_1058 (O_1058,N_9513,N_8012);
and UO_1059 (O_1059,N_8926,N_8169);
or UO_1060 (O_1060,N_8698,N_8003);
or UO_1061 (O_1061,N_8876,N_8015);
nand UO_1062 (O_1062,N_8405,N_9294);
and UO_1063 (O_1063,N_8571,N_8415);
xor UO_1064 (O_1064,N_8406,N_8615);
nor UO_1065 (O_1065,N_8870,N_9254);
nand UO_1066 (O_1066,N_8678,N_8240);
nor UO_1067 (O_1067,N_8005,N_9418);
nand UO_1068 (O_1068,N_8219,N_9072);
nand UO_1069 (O_1069,N_9048,N_9098);
nand UO_1070 (O_1070,N_9386,N_8060);
nand UO_1071 (O_1071,N_8669,N_8673);
and UO_1072 (O_1072,N_9972,N_8031);
nor UO_1073 (O_1073,N_9463,N_9981);
nand UO_1074 (O_1074,N_8265,N_8101);
or UO_1075 (O_1075,N_9362,N_9054);
nor UO_1076 (O_1076,N_9260,N_8292);
nand UO_1077 (O_1077,N_8019,N_8287);
nor UO_1078 (O_1078,N_8038,N_9589);
and UO_1079 (O_1079,N_9009,N_8646);
nor UO_1080 (O_1080,N_9543,N_8956);
or UO_1081 (O_1081,N_8919,N_8689);
or UO_1082 (O_1082,N_8257,N_8375);
and UO_1083 (O_1083,N_8484,N_8149);
or UO_1084 (O_1084,N_9554,N_9237);
or UO_1085 (O_1085,N_9689,N_8571);
nand UO_1086 (O_1086,N_8172,N_8194);
and UO_1087 (O_1087,N_8581,N_8107);
and UO_1088 (O_1088,N_9618,N_8820);
and UO_1089 (O_1089,N_9525,N_8252);
nand UO_1090 (O_1090,N_8128,N_8469);
or UO_1091 (O_1091,N_8194,N_9982);
nor UO_1092 (O_1092,N_8466,N_9081);
and UO_1093 (O_1093,N_8321,N_9302);
nor UO_1094 (O_1094,N_8240,N_8044);
nand UO_1095 (O_1095,N_9347,N_8280);
xor UO_1096 (O_1096,N_8561,N_8991);
nand UO_1097 (O_1097,N_8367,N_9053);
nor UO_1098 (O_1098,N_8599,N_8654);
xnor UO_1099 (O_1099,N_8032,N_9481);
or UO_1100 (O_1100,N_9049,N_8245);
and UO_1101 (O_1101,N_8120,N_9462);
and UO_1102 (O_1102,N_9940,N_8603);
nor UO_1103 (O_1103,N_8908,N_9438);
nor UO_1104 (O_1104,N_8605,N_9962);
nand UO_1105 (O_1105,N_9121,N_9405);
nand UO_1106 (O_1106,N_9457,N_8540);
nor UO_1107 (O_1107,N_8395,N_8856);
or UO_1108 (O_1108,N_8588,N_9884);
nor UO_1109 (O_1109,N_8357,N_8286);
nor UO_1110 (O_1110,N_8660,N_8959);
nand UO_1111 (O_1111,N_9860,N_8567);
or UO_1112 (O_1112,N_9626,N_8694);
nor UO_1113 (O_1113,N_8130,N_8060);
nor UO_1114 (O_1114,N_8020,N_8984);
and UO_1115 (O_1115,N_8100,N_8565);
and UO_1116 (O_1116,N_9375,N_8305);
nor UO_1117 (O_1117,N_9547,N_9885);
nor UO_1118 (O_1118,N_9763,N_9603);
and UO_1119 (O_1119,N_9446,N_9191);
nor UO_1120 (O_1120,N_9188,N_8944);
or UO_1121 (O_1121,N_8091,N_8176);
and UO_1122 (O_1122,N_8497,N_9622);
and UO_1123 (O_1123,N_8900,N_9783);
and UO_1124 (O_1124,N_9061,N_9481);
or UO_1125 (O_1125,N_8316,N_8740);
and UO_1126 (O_1126,N_8606,N_9293);
nand UO_1127 (O_1127,N_8348,N_8853);
and UO_1128 (O_1128,N_8741,N_9734);
nor UO_1129 (O_1129,N_8643,N_8890);
and UO_1130 (O_1130,N_8066,N_8544);
nor UO_1131 (O_1131,N_8456,N_9004);
nor UO_1132 (O_1132,N_8950,N_9912);
or UO_1133 (O_1133,N_9568,N_8104);
and UO_1134 (O_1134,N_8405,N_8647);
or UO_1135 (O_1135,N_9678,N_8839);
nor UO_1136 (O_1136,N_9983,N_9858);
or UO_1137 (O_1137,N_8741,N_9024);
or UO_1138 (O_1138,N_9987,N_9724);
nand UO_1139 (O_1139,N_9743,N_9028);
nor UO_1140 (O_1140,N_9001,N_8112);
nor UO_1141 (O_1141,N_8642,N_9988);
or UO_1142 (O_1142,N_9671,N_9589);
nor UO_1143 (O_1143,N_8450,N_8309);
xor UO_1144 (O_1144,N_9652,N_9697);
or UO_1145 (O_1145,N_8271,N_8878);
nand UO_1146 (O_1146,N_8600,N_9721);
xor UO_1147 (O_1147,N_8029,N_9027);
nand UO_1148 (O_1148,N_9242,N_8913);
nand UO_1149 (O_1149,N_9899,N_8859);
nand UO_1150 (O_1150,N_8541,N_8230);
and UO_1151 (O_1151,N_9118,N_9488);
nor UO_1152 (O_1152,N_9549,N_8909);
and UO_1153 (O_1153,N_8074,N_8925);
or UO_1154 (O_1154,N_8200,N_8056);
and UO_1155 (O_1155,N_8948,N_8553);
or UO_1156 (O_1156,N_8555,N_9079);
nor UO_1157 (O_1157,N_9533,N_9411);
xnor UO_1158 (O_1158,N_9248,N_9872);
nand UO_1159 (O_1159,N_8816,N_9633);
nor UO_1160 (O_1160,N_9159,N_9182);
and UO_1161 (O_1161,N_8698,N_9369);
and UO_1162 (O_1162,N_8866,N_9936);
and UO_1163 (O_1163,N_8650,N_9644);
nor UO_1164 (O_1164,N_9341,N_8215);
nor UO_1165 (O_1165,N_8678,N_9393);
and UO_1166 (O_1166,N_8687,N_8748);
and UO_1167 (O_1167,N_9563,N_8888);
or UO_1168 (O_1168,N_8224,N_9276);
and UO_1169 (O_1169,N_9431,N_8102);
nor UO_1170 (O_1170,N_9294,N_9804);
or UO_1171 (O_1171,N_9029,N_8037);
nor UO_1172 (O_1172,N_9473,N_9331);
nor UO_1173 (O_1173,N_8294,N_9995);
nand UO_1174 (O_1174,N_9539,N_9555);
and UO_1175 (O_1175,N_9572,N_8024);
or UO_1176 (O_1176,N_8656,N_8905);
nand UO_1177 (O_1177,N_8800,N_9783);
nand UO_1178 (O_1178,N_9578,N_8457);
nor UO_1179 (O_1179,N_8808,N_9740);
nor UO_1180 (O_1180,N_9486,N_9093);
or UO_1181 (O_1181,N_9016,N_9371);
or UO_1182 (O_1182,N_8453,N_8378);
nor UO_1183 (O_1183,N_8089,N_9700);
and UO_1184 (O_1184,N_8804,N_9886);
nor UO_1185 (O_1185,N_9816,N_9772);
nor UO_1186 (O_1186,N_8785,N_8492);
or UO_1187 (O_1187,N_8547,N_9091);
nor UO_1188 (O_1188,N_9830,N_8019);
or UO_1189 (O_1189,N_8213,N_9185);
nor UO_1190 (O_1190,N_8662,N_9024);
nor UO_1191 (O_1191,N_8666,N_9442);
nand UO_1192 (O_1192,N_8855,N_9378);
and UO_1193 (O_1193,N_9466,N_9905);
nand UO_1194 (O_1194,N_9169,N_8421);
nand UO_1195 (O_1195,N_8845,N_8790);
and UO_1196 (O_1196,N_8863,N_9012);
or UO_1197 (O_1197,N_9272,N_8635);
nand UO_1198 (O_1198,N_8234,N_9419);
nor UO_1199 (O_1199,N_9753,N_9671);
and UO_1200 (O_1200,N_9481,N_9419);
nor UO_1201 (O_1201,N_8268,N_8043);
nand UO_1202 (O_1202,N_8790,N_8152);
or UO_1203 (O_1203,N_8957,N_9485);
or UO_1204 (O_1204,N_8008,N_9628);
nor UO_1205 (O_1205,N_9778,N_8986);
nand UO_1206 (O_1206,N_9006,N_9342);
nor UO_1207 (O_1207,N_8160,N_9230);
nor UO_1208 (O_1208,N_9403,N_9656);
or UO_1209 (O_1209,N_8962,N_9998);
nand UO_1210 (O_1210,N_9348,N_8989);
nand UO_1211 (O_1211,N_8765,N_8553);
nor UO_1212 (O_1212,N_8031,N_8244);
or UO_1213 (O_1213,N_8894,N_8066);
nand UO_1214 (O_1214,N_8914,N_9475);
or UO_1215 (O_1215,N_8797,N_9209);
and UO_1216 (O_1216,N_8534,N_8523);
and UO_1217 (O_1217,N_9424,N_8401);
or UO_1218 (O_1218,N_9010,N_9466);
and UO_1219 (O_1219,N_8245,N_9203);
or UO_1220 (O_1220,N_8091,N_8487);
or UO_1221 (O_1221,N_8169,N_8422);
nor UO_1222 (O_1222,N_9957,N_9383);
nor UO_1223 (O_1223,N_8960,N_8670);
or UO_1224 (O_1224,N_8155,N_9701);
or UO_1225 (O_1225,N_9725,N_8970);
and UO_1226 (O_1226,N_8744,N_9579);
nand UO_1227 (O_1227,N_9262,N_9583);
or UO_1228 (O_1228,N_9174,N_9743);
nor UO_1229 (O_1229,N_8425,N_8558);
or UO_1230 (O_1230,N_9975,N_9189);
nor UO_1231 (O_1231,N_8097,N_9220);
and UO_1232 (O_1232,N_8076,N_9730);
nand UO_1233 (O_1233,N_9992,N_8006);
and UO_1234 (O_1234,N_9764,N_8521);
nor UO_1235 (O_1235,N_9263,N_8210);
nor UO_1236 (O_1236,N_9385,N_9851);
nand UO_1237 (O_1237,N_8043,N_8281);
or UO_1238 (O_1238,N_8213,N_9288);
nor UO_1239 (O_1239,N_9249,N_9011);
nor UO_1240 (O_1240,N_8050,N_9448);
or UO_1241 (O_1241,N_9976,N_8898);
and UO_1242 (O_1242,N_9073,N_8682);
nand UO_1243 (O_1243,N_9579,N_9077);
and UO_1244 (O_1244,N_9839,N_8994);
or UO_1245 (O_1245,N_9837,N_8222);
nor UO_1246 (O_1246,N_9224,N_8140);
or UO_1247 (O_1247,N_8230,N_9594);
nand UO_1248 (O_1248,N_8824,N_9995);
and UO_1249 (O_1249,N_8352,N_9190);
or UO_1250 (O_1250,N_8703,N_8721);
or UO_1251 (O_1251,N_9701,N_9145);
and UO_1252 (O_1252,N_8070,N_9854);
or UO_1253 (O_1253,N_8742,N_9096);
nand UO_1254 (O_1254,N_9977,N_9167);
nand UO_1255 (O_1255,N_9447,N_8045);
xnor UO_1256 (O_1256,N_8777,N_9206);
nand UO_1257 (O_1257,N_8712,N_9156);
nor UO_1258 (O_1258,N_8424,N_8606);
or UO_1259 (O_1259,N_8762,N_9848);
and UO_1260 (O_1260,N_9185,N_9189);
and UO_1261 (O_1261,N_8845,N_8552);
or UO_1262 (O_1262,N_9307,N_8333);
nand UO_1263 (O_1263,N_9495,N_8503);
or UO_1264 (O_1264,N_9272,N_8939);
or UO_1265 (O_1265,N_9142,N_9170);
nand UO_1266 (O_1266,N_8376,N_9686);
or UO_1267 (O_1267,N_8125,N_8581);
or UO_1268 (O_1268,N_8835,N_8009);
and UO_1269 (O_1269,N_8257,N_9627);
nor UO_1270 (O_1270,N_9805,N_8084);
nand UO_1271 (O_1271,N_8253,N_8642);
and UO_1272 (O_1272,N_9266,N_9409);
nand UO_1273 (O_1273,N_8655,N_9620);
nor UO_1274 (O_1274,N_8610,N_9820);
or UO_1275 (O_1275,N_9520,N_9282);
or UO_1276 (O_1276,N_9704,N_8493);
nand UO_1277 (O_1277,N_9770,N_8348);
nand UO_1278 (O_1278,N_9256,N_8442);
nor UO_1279 (O_1279,N_9026,N_9303);
or UO_1280 (O_1280,N_8606,N_8931);
and UO_1281 (O_1281,N_9315,N_9357);
or UO_1282 (O_1282,N_8351,N_8811);
and UO_1283 (O_1283,N_9858,N_8770);
and UO_1284 (O_1284,N_8470,N_8855);
or UO_1285 (O_1285,N_8763,N_8979);
and UO_1286 (O_1286,N_8010,N_9953);
nor UO_1287 (O_1287,N_8549,N_8211);
nor UO_1288 (O_1288,N_8129,N_8616);
nor UO_1289 (O_1289,N_9259,N_8021);
and UO_1290 (O_1290,N_9472,N_8661);
and UO_1291 (O_1291,N_9709,N_9894);
and UO_1292 (O_1292,N_8728,N_9255);
nor UO_1293 (O_1293,N_8125,N_8960);
and UO_1294 (O_1294,N_9684,N_9266);
nand UO_1295 (O_1295,N_9752,N_8060);
nor UO_1296 (O_1296,N_8286,N_9559);
xor UO_1297 (O_1297,N_9219,N_9802);
and UO_1298 (O_1298,N_8857,N_9163);
and UO_1299 (O_1299,N_9758,N_8615);
nor UO_1300 (O_1300,N_9706,N_9906);
nand UO_1301 (O_1301,N_9987,N_8232);
or UO_1302 (O_1302,N_9406,N_8076);
xnor UO_1303 (O_1303,N_9036,N_8137);
nor UO_1304 (O_1304,N_8927,N_9809);
nor UO_1305 (O_1305,N_9503,N_9266);
and UO_1306 (O_1306,N_9433,N_9072);
and UO_1307 (O_1307,N_8575,N_9014);
nand UO_1308 (O_1308,N_8533,N_9111);
nor UO_1309 (O_1309,N_8250,N_8632);
nand UO_1310 (O_1310,N_8056,N_9548);
and UO_1311 (O_1311,N_9625,N_8899);
nand UO_1312 (O_1312,N_9218,N_8876);
nor UO_1313 (O_1313,N_9971,N_8214);
nand UO_1314 (O_1314,N_8368,N_9006);
and UO_1315 (O_1315,N_9327,N_9534);
nor UO_1316 (O_1316,N_8101,N_9232);
and UO_1317 (O_1317,N_8752,N_8578);
nand UO_1318 (O_1318,N_9751,N_8415);
nor UO_1319 (O_1319,N_8226,N_8374);
or UO_1320 (O_1320,N_9155,N_9100);
or UO_1321 (O_1321,N_8427,N_8235);
and UO_1322 (O_1322,N_9698,N_9120);
or UO_1323 (O_1323,N_8856,N_8526);
and UO_1324 (O_1324,N_8453,N_9967);
nor UO_1325 (O_1325,N_8238,N_9755);
nand UO_1326 (O_1326,N_9867,N_8616);
nand UO_1327 (O_1327,N_9027,N_8969);
or UO_1328 (O_1328,N_8027,N_8548);
and UO_1329 (O_1329,N_8853,N_8825);
nand UO_1330 (O_1330,N_9382,N_9534);
nor UO_1331 (O_1331,N_8667,N_8966);
nor UO_1332 (O_1332,N_9512,N_9345);
xnor UO_1333 (O_1333,N_8765,N_8980);
xnor UO_1334 (O_1334,N_8316,N_9467);
or UO_1335 (O_1335,N_8904,N_9955);
xor UO_1336 (O_1336,N_8534,N_9532);
nand UO_1337 (O_1337,N_9496,N_8922);
nand UO_1338 (O_1338,N_8469,N_9402);
or UO_1339 (O_1339,N_8209,N_8100);
nor UO_1340 (O_1340,N_8886,N_8480);
nor UO_1341 (O_1341,N_8571,N_8318);
and UO_1342 (O_1342,N_8256,N_9324);
nor UO_1343 (O_1343,N_8247,N_8646);
nor UO_1344 (O_1344,N_8962,N_9607);
nor UO_1345 (O_1345,N_8566,N_9759);
nor UO_1346 (O_1346,N_8931,N_8969);
or UO_1347 (O_1347,N_9183,N_8915);
and UO_1348 (O_1348,N_9323,N_9285);
nor UO_1349 (O_1349,N_9658,N_9471);
and UO_1350 (O_1350,N_9749,N_8867);
or UO_1351 (O_1351,N_9576,N_8159);
nor UO_1352 (O_1352,N_8330,N_8885);
nor UO_1353 (O_1353,N_8586,N_9836);
and UO_1354 (O_1354,N_9077,N_9130);
nand UO_1355 (O_1355,N_8733,N_8516);
nor UO_1356 (O_1356,N_8846,N_9153);
and UO_1357 (O_1357,N_8916,N_9154);
nor UO_1358 (O_1358,N_8569,N_9816);
and UO_1359 (O_1359,N_9336,N_8983);
or UO_1360 (O_1360,N_9327,N_9148);
nand UO_1361 (O_1361,N_9628,N_9871);
nor UO_1362 (O_1362,N_9322,N_9239);
and UO_1363 (O_1363,N_9522,N_8437);
nand UO_1364 (O_1364,N_8190,N_8000);
nand UO_1365 (O_1365,N_8489,N_8592);
nand UO_1366 (O_1366,N_9586,N_9306);
nor UO_1367 (O_1367,N_8493,N_9718);
nand UO_1368 (O_1368,N_8842,N_9665);
nand UO_1369 (O_1369,N_9185,N_9740);
and UO_1370 (O_1370,N_8918,N_8379);
or UO_1371 (O_1371,N_8911,N_8491);
and UO_1372 (O_1372,N_9230,N_8263);
nor UO_1373 (O_1373,N_9068,N_8297);
and UO_1374 (O_1374,N_9916,N_8465);
nor UO_1375 (O_1375,N_9590,N_8621);
and UO_1376 (O_1376,N_8907,N_9624);
or UO_1377 (O_1377,N_9161,N_8364);
nor UO_1378 (O_1378,N_8344,N_9148);
and UO_1379 (O_1379,N_9975,N_9115);
and UO_1380 (O_1380,N_9233,N_8337);
nand UO_1381 (O_1381,N_8840,N_9003);
nor UO_1382 (O_1382,N_8854,N_9221);
or UO_1383 (O_1383,N_8168,N_9556);
nor UO_1384 (O_1384,N_9590,N_8636);
or UO_1385 (O_1385,N_9747,N_9505);
nor UO_1386 (O_1386,N_8213,N_9824);
or UO_1387 (O_1387,N_9502,N_9536);
nand UO_1388 (O_1388,N_8415,N_8707);
nand UO_1389 (O_1389,N_8185,N_9017);
and UO_1390 (O_1390,N_9572,N_8506);
nor UO_1391 (O_1391,N_9824,N_8203);
and UO_1392 (O_1392,N_9697,N_9168);
or UO_1393 (O_1393,N_8020,N_9509);
and UO_1394 (O_1394,N_8370,N_8916);
nor UO_1395 (O_1395,N_9172,N_8256);
nand UO_1396 (O_1396,N_9173,N_8657);
and UO_1397 (O_1397,N_9318,N_9843);
nand UO_1398 (O_1398,N_9864,N_9329);
xor UO_1399 (O_1399,N_8385,N_9317);
nor UO_1400 (O_1400,N_9800,N_8947);
nor UO_1401 (O_1401,N_9824,N_8967);
nand UO_1402 (O_1402,N_8508,N_9250);
and UO_1403 (O_1403,N_8050,N_9229);
and UO_1404 (O_1404,N_9679,N_9286);
nor UO_1405 (O_1405,N_9627,N_9384);
or UO_1406 (O_1406,N_9713,N_9962);
or UO_1407 (O_1407,N_9898,N_8285);
nor UO_1408 (O_1408,N_9565,N_8163);
or UO_1409 (O_1409,N_8158,N_9830);
nand UO_1410 (O_1410,N_8224,N_8302);
nor UO_1411 (O_1411,N_8181,N_8847);
nand UO_1412 (O_1412,N_9131,N_9561);
nor UO_1413 (O_1413,N_9719,N_8046);
nor UO_1414 (O_1414,N_8066,N_9560);
nor UO_1415 (O_1415,N_8288,N_9036);
or UO_1416 (O_1416,N_9030,N_8168);
or UO_1417 (O_1417,N_8257,N_8437);
nor UO_1418 (O_1418,N_9080,N_9141);
nor UO_1419 (O_1419,N_8487,N_9255);
and UO_1420 (O_1420,N_8740,N_9024);
nand UO_1421 (O_1421,N_8994,N_8881);
and UO_1422 (O_1422,N_8235,N_8359);
or UO_1423 (O_1423,N_9760,N_9835);
or UO_1424 (O_1424,N_8957,N_9880);
nor UO_1425 (O_1425,N_9844,N_8020);
and UO_1426 (O_1426,N_8577,N_8201);
xnor UO_1427 (O_1427,N_8186,N_8901);
or UO_1428 (O_1428,N_8209,N_8019);
or UO_1429 (O_1429,N_9010,N_8489);
or UO_1430 (O_1430,N_9278,N_8510);
or UO_1431 (O_1431,N_9448,N_9801);
nor UO_1432 (O_1432,N_9016,N_9439);
nand UO_1433 (O_1433,N_8601,N_9306);
and UO_1434 (O_1434,N_8225,N_9629);
or UO_1435 (O_1435,N_8047,N_8778);
and UO_1436 (O_1436,N_9965,N_9326);
or UO_1437 (O_1437,N_8012,N_8052);
nor UO_1438 (O_1438,N_8991,N_8548);
and UO_1439 (O_1439,N_8664,N_9463);
or UO_1440 (O_1440,N_9169,N_9623);
or UO_1441 (O_1441,N_8395,N_8657);
or UO_1442 (O_1442,N_8084,N_9979);
or UO_1443 (O_1443,N_9129,N_9140);
and UO_1444 (O_1444,N_8980,N_8903);
nand UO_1445 (O_1445,N_8326,N_9499);
nand UO_1446 (O_1446,N_8566,N_8173);
nand UO_1447 (O_1447,N_9184,N_8516);
nor UO_1448 (O_1448,N_9533,N_9706);
and UO_1449 (O_1449,N_8393,N_8103);
or UO_1450 (O_1450,N_9499,N_8863);
nor UO_1451 (O_1451,N_9927,N_9530);
xor UO_1452 (O_1452,N_8836,N_8680);
and UO_1453 (O_1453,N_9307,N_9118);
nor UO_1454 (O_1454,N_9049,N_8926);
or UO_1455 (O_1455,N_8223,N_8497);
or UO_1456 (O_1456,N_8314,N_9578);
and UO_1457 (O_1457,N_9943,N_9206);
and UO_1458 (O_1458,N_8843,N_8663);
or UO_1459 (O_1459,N_8565,N_9451);
and UO_1460 (O_1460,N_8016,N_9817);
and UO_1461 (O_1461,N_9263,N_8986);
nor UO_1462 (O_1462,N_8096,N_9812);
and UO_1463 (O_1463,N_9821,N_9197);
or UO_1464 (O_1464,N_8828,N_9106);
xnor UO_1465 (O_1465,N_8081,N_9705);
and UO_1466 (O_1466,N_8247,N_9424);
and UO_1467 (O_1467,N_9745,N_9564);
or UO_1468 (O_1468,N_9839,N_9080);
nand UO_1469 (O_1469,N_9445,N_9440);
nand UO_1470 (O_1470,N_9294,N_9543);
nand UO_1471 (O_1471,N_9270,N_8644);
nand UO_1472 (O_1472,N_9264,N_8768);
nand UO_1473 (O_1473,N_8154,N_9759);
and UO_1474 (O_1474,N_9890,N_8135);
nor UO_1475 (O_1475,N_9970,N_9813);
and UO_1476 (O_1476,N_8977,N_8822);
or UO_1477 (O_1477,N_8197,N_9458);
and UO_1478 (O_1478,N_8422,N_8875);
and UO_1479 (O_1479,N_9453,N_9962);
and UO_1480 (O_1480,N_8346,N_8029);
nor UO_1481 (O_1481,N_9376,N_9920);
nor UO_1482 (O_1482,N_8155,N_9321);
nor UO_1483 (O_1483,N_9909,N_8373);
and UO_1484 (O_1484,N_9222,N_8379);
nor UO_1485 (O_1485,N_9172,N_8626);
xnor UO_1486 (O_1486,N_8616,N_9618);
nand UO_1487 (O_1487,N_9869,N_8879);
nand UO_1488 (O_1488,N_8570,N_8652);
nand UO_1489 (O_1489,N_8235,N_8504);
nor UO_1490 (O_1490,N_8980,N_9092);
xnor UO_1491 (O_1491,N_9970,N_8967);
nand UO_1492 (O_1492,N_9138,N_9419);
and UO_1493 (O_1493,N_8010,N_8481);
or UO_1494 (O_1494,N_8975,N_8442);
and UO_1495 (O_1495,N_8174,N_8354);
nand UO_1496 (O_1496,N_9483,N_8058);
nor UO_1497 (O_1497,N_8496,N_8569);
nand UO_1498 (O_1498,N_9729,N_8028);
or UO_1499 (O_1499,N_8822,N_8090);
endmodule