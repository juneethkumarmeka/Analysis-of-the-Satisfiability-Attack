module basic_500_3000_500_4_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_118,In_329);
nand U1 (N_1,In_222,In_301);
nor U2 (N_2,In_185,In_424);
nor U3 (N_3,In_278,In_60);
nand U4 (N_4,In_23,In_227);
nor U5 (N_5,In_228,In_247);
and U6 (N_6,In_498,In_359);
nor U7 (N_7,In_331,In_203);
or U8 (N_8,In_148,In_313);
nand U9 (N_9,In_262,In_320);
nor U10 (N_10,In_443,In_92);
and U11 (N_11,In_449,In_404);
or U12 (N_12,In_490,In_171);
nor U13 (N_13,In_215,In_459);
nand U14 (N_14,In_4,In_131);
and U15 (N_15,In_432,In_62);
or U16 (N_16,In_241,In_291);
xor U17 (N_17,In_16,In_188);
xor U18 (N_18,In_415,In_343);
nor U19 (N_19,In_173,In_18);
xor U20 (N_20,In_293,In_63);
nor U21 (N_21,In_493,In_226);
nor U22 (N_22,In_39,In_183);
or U23 (N_23,In_192,In_378);
nor U24 (N_24,In_371,In_104);
nand U25 (N_25,In_152,In_91);
or U26 (N_26,In_204,In_54);
nand U27 (N_27,In_272,In_349);
and U28 (N_28,In_164,In_207);
or U29 (N_29,In_335,In_474);
xor U30 (N_30,In_158,In_242);
nand U31 (N_31,In_24,In_315);
or U32 (N_32,In_191,In_6);
nor U33 (N_33,In_360,In_64);
or U34 (N_34,In_20,In_362);
nand U35 (N_35,In_211,In_441);
and U36 (N_36,In_466,In_197);
nand U37 (N_37,In_477,In_352);
and U38 (N_38,In_412,In_193);
nor U39 (N_39,In_475,In_346);
nand U40 (N_40,In_271,In_409);
or U41 (N_41,In_422,In_107);
or U42 (N_42,In_196,In_316);
nand U43 (N_43,In_119,In_435);
and U44 (N_44,In_369,In_174);
xnor U45 (N_45,In_172,In_431);
and U46 (N_46,In_7,In_296);
xor U47 (N_47,In_421,In_200);
or U48 (N_48,In_51,In_299);
and U49 (N_49,In_396,In_476);
nand U50 (N_50,In_465,In_334);
or U51 (N_51,In_286,In_22);
or U52 (N_52,In_43,In_231);
nand U53 (N_53,In_442,In_143);
nand U54 (N_54,In_394,In_95);
nand U55 (N_55,In_217,In_52);
and U56 (N_56,In_125,In_235);
or U57 (N_57,In_406,In_232);
nand U58 (N_58,In_113,In_120);
and U59 (N_59,In_298,In_85);
nor U60 (N_60,In_489,In_124);
nor U61 (N_61,In_492,In_347);
nand U62 (N_62,In_336,In_309);
or U63 (N_63,In_410,In_59);
and U64 (N_64,In_450,In_479);
nand U65 (N_65,In_234,In_401);
nand U66 (N_66,In_209,In_236);
or U67 (N_67,In_245,In_267);
or U68 (N_68,In_13,In_295);
or U69 (N_69,In_283,In_150);
and U70 (N_70,In_5,In_244);
or U71 (N_71,In_494,In_99);
or U72 (N_72,In_134,In_314);
or U73 (N_73,In_463,In_32);
and U74 (N_74,In_468,In_121);
nor U75 (N_75,In_408,In_73);
or U76 (N_76,In_497,In_74);
nand U77 (N_77,In_201,In_42);
nor U78 (N_78,In_169,In_116);
and U79 (N_79,In_65,In_472);
and U80 (N_80,In_260,In_444);
and U81 (N_81,In_275,In_71);
nor U82 (N_82,In_327,In_375);
xnor U83 (N_83,In_487,In_344);
xor U84 (N_84,In_36,In_302);
xnor U85 (N_85,In_438,In_189);
or U86 (N_86,In_257,In_46);
nor U87 (N_87,In_282,In_304);
and U88 (N_88,In_256,In_470);
and U89 (N_89,In_445,In_87);
nand U90 (N_90,In_212,In_11);
nor U91 (N_91,In_276,In_128);
or U92 (N_92,In_457,In_354);
nand U93 (N_93,In_337,In_14);
and U94 (N_94,In_420,In_138);
or U95 (N_95,In_265,In_345);
and U96 (N_96,In_248,In_102);
or U97 (N_97,In_111,In_467);
and U98 (N_98,In_130,In_103);
and U99 (N_99,In_80,In_368);
nand U100 (N_100,In_142,In_448);
or U101 (N_101,In_68,In_277);
nand U102 (N_102,In_194,In_2);
nand U103 (N_103,In_122,In_210);
and U104 (N_104,In_440,In_198);
nand U105 (N_105,In_446,In_168);
or U106 (N_106,In_53,In_289);
or U107 (N_107,In_384,In_31);
or U108 (N_108,In_478,In_153);
nor U109 (N_109,In_108,In_139);
or U110 (N_110,In_340,In_380);
and U111 (N_111,In_429,In_311);
nand U112 (N_112,In_184,In_392);
nand U113 (N_113,In_310,In_141);
and U114 (N_114,In_307,In_373);
xnor U115 (N_115,In_269,In_281);
nor U116 (N_116,In_3,In_97);
and U117 (N_117,In_284,In_195);
nand U118 (N_118,In_253,In_25);
nand U119 (N_119,In_0,In_90);
nand U120 (N_120,In_55,In_83);
or U121 (N_121,In_485,In_224);
and U122 (N_122,In_67,In_140);
nand U123 (N_123,In_136,In_40);
nand U124 (N_124,In_179,In_387);
and U125 (N_125,In_82,In_353);
or U126 (N_126,In_213,In_145);
and U127 (N_127,In_250,In_325);
or U128 (N_128,In_177,In_280);
xor U129 (N_129,In_482,In_333);
or U130 (N_130,In_259,In_312);
nand U131 (N_131,In_88,In_418);
nand U132 (N_132,In_416,In_390);
nor U133 (N_133,In_132,In_484);
or U134 (N_134,In_330,In_464);
and U135 (N_135,In_423,In_214);
nor U136 (N_136,In_338,In_402);
nand U137 (N_137,In_37,In_400);
and U138 (N_138,In_377,In_414);
nor U139 (N_139,In_285,In_341);
nor U140 (N_140,In_1,In_181);
and U141 (N_141,In_462,In_255);
and U142 (N_142,In_399,In_49);
nand U143 (N_143,In_9,In_61);
nand U144 (N_144,In_389,In_274);
nand U145 (N_145,In_86,In_317);
and U146 (N_146,In_160,In_461);
nand U147 (N_147,In_486,In_318);
nor U148 (N_148,In_50,In_33);
nor U149 (N_149,In_163,In_100);
nor U150 (N_150,In_319,In_385);
nor U151 (N_151,In_10,In_225);
xor U152 (N_152,In_292,In_456);
xnor U153 (N_153,In_306,In_56);
nand U154 (N_154,In_84,In_187);
or U155 (N_155,In_21,In_287);
or U156 (N_156,In_175,In_167);
and U157 (N_157,In_428,In_382);
nor U158 (N_158,In_202,In_28);
or U159 (N_159,In_279,In_126);
nand U160 (N_160,In_154,In_366);
and U161 (N_161,In_17,In_324);
and U162 (N_162,In_115,In_238);
nor U163 (N_163,In_72,In_166);
nor U164 (N_164,In_452,In_146);
nand U165 (N_165,In_199,In_129);
nor U166 (N_166,In_391,In_495);
and U167 (N_167,In_162,In_41);
xnor U168 (N_168,In_161,In_155);
or U169 (N_169,In_35,In_261);
or U170 (N_170,In_254,In_270);
or U171 (N_171,In_332,In_297);
nor U172 (N_172,In_433,In_308);
and U173 (N_173,In_182,In_427);
and U174 (N_174,In_117,In_112);
nor U175 (N_175,In_263,In_388);
xnor U176 (N_176,In_451,In_469);
nor U177 (N_177,In_403,In_361);
or U178 (N_178,In_426,In_106);
nor U179 (N_179,In_439,In_45);
nor U180 (N_180,In_101,In_34);
or U181 (N_181,In_290,In_437);
or U182 (N_182,In_157,In_96);
nor U183 (N_183,In_499,In_237);
and U184 (N_184,In_326,In_246);
and U185 (N_185,In_149,In_358);
and U186 (N_186,In_381,In_363);
xor U187 (N_187,In_481,In_109);
and U188 (N_188,In_454,In_205);
nor U189 (N_189,In_342,In_348);
and U190 (N_190,In_480,In_81);
or U191 (N_191,In_133,In_70);
nor U192 (N_192,In_218,In_239);
or U193 (N_193,In_434,In_137);
nor U194 (N_194,In_127,In_57);
nor U195 (N_195,In_288,In_75);
or U196 (N_196,In_110,In_294);
and U197 (N_197,In_27,In_233);
xor U198 (N_198,In_273,In_219);
nor U199 (N_199,In_252,In_58);
nand U200 (N_200,In_144,In_156);
and U201 (N_201,In_176,In_407);
nor U202 (N_202,In_93,In_78);
or U203 (N_203,In_483,In_393);
or U204 (N_204,In_223,In_165);
nand U205 (N_205,In_47,In_147);
or U206 (N_206,In_398,In_491);
or U207 (N_207,In_488,In_220);
or U208 (N_208,In_370,In_365);
nand U209 (N_209,In_395,In_471);
nor U210 (N_210,In_240,In_372);
xor U211 (N_211,In_496,In_114);
nand U212 (N_212,In_30,In_98);
nor U213 (N_213,In_397,In_15);
nand U214 (N_214,In_453,In_249);
or U215 (N_215,In_123,In_44);
nor U216 (N_216,In_351,In_221);
nand U217 (N_217,In_321,In_460);
or U218 (N_218,In_208,In_425);
xnor U219 (N_219,In_386,In_300);
or U220 (N_220,In_350,In_376);
or U221 (N_221,In_251,In_48);
nor U222 (N_222,In_186,In_19);
nand U223 (N_223,In_229,In_328);
nor U224 (N_224,In_89,In_264);
xor U225 (N_225,In_411,In_364);
and U226 (N_226,In_473,In_374);
nand U227 (N_227,In_405,In_206);
and U228 (N_228,In_458,In_8);
and U229 (N_229,In_367,In_180);
nand U230 (N_230,In_26,In_12);
or U231 (N_231,In_419,In_305);
and U232 (N_232,In_436,In_178);
and U233 (N_233,In_135,In_323);
nor U234 (N_234,In_76,In_105);
nor U235 (N_235,In_170,In_383);
and U236 (N_236,In_151,In_66);
nor U237 (N_237,In_266,In_230);
and U238 (N_238,In_357,In_455);
or U239 (N_239,In_243,In_339);
xnor U240 (N_240,In_79,In_29);
nand U241 (N_241,In_69,In_190);
xnor U242 (N_242,In_303,In_94);
nor U243 (N_243,In_430,In_413);
nand U244 (N_244,In_379,In_356);
and U245 (N_245,In_77,In_258);
xnor U246 (N_246,In_268,In_322);
and U247 (N_247,In_447,In_38);
and U248 (N_248,In_417,In_216);
nand U249 (N_249,In_159,In_355);
or U250 (N_250,In_165,In_252);
xnor U251 (N_251,In_351,In_20);
nand U252 (N_252,In_364,In_213);
nand U253 (N_253,In_95,In_57);
and U254 (N_254,In_468,In_95);
nor U255 (N_255,In_439,In_265);
and U256 (N_256,In_136,In_174);
and U257 (N_257,In_73,In_244);
nand U258 (N_258,In_414,In_6);
or U259 (N_259,In_384,In_276);
or U260 (N_260,In_424,In_365);
and U261 (N_261,In_423,In_8);
or U262 (N_262,In_432,In_205);
nor U263 (N_263,In_326,In_172);
and U264 (N_264,In_296,In_352);
nand U265 (N_265,In_340,In_304);
nor U266 (N_266,In_397,In_87);
and U267 (N_267,In_58,In_447);
nor U268 (N_268,In_30,In_118);
nor U269 (N_269,In_221,In_332);
and U270 (N_270,In_153,In_347);
and U271 (N_271,In_313,In_183);
xnor U272 (N_272,In_371,In_125);
nor U273 (N_273,In_291,In_58);
or U274 (N_274,In_278,In_420);
nor U275 (N_275,In_187,In_5);
xnor U276 (N_276,In_379,In_344);
or U277 (N_277,In_62,In_255);
nand U278 (N_278,In_252,In_478);
and U279 (N_279,In_289,In_496);
xnor U280 (N_280,In_130,In_473);
and U281 (N_281,In_260,In_224);
xnor U282 (N_282,In_83,In_468);
and U283 (N_283,In_189,In_190);
nand U284 (N_284,In_444,In_263);
xor U285 (N_285,In_199,In_289);
and U286 (N_286,In_475,In_155);
nor U287 (N_287,In_333,In_0);
and U288 (N_288,In_123,In_432);
nor U289 (N_289,In_406,In_285);
nand U290 (N_290,In_65,In_146);
nand U291 (N_291,In_467,In_275);
xor U292 (N_292,In_207,In_320);
and U293 (N_293,In_139,In_52);
or U294 (N_294,In_76,In_60);
nor U295 (N_295,In_93,In_284);
nand U296 (N_296,In_340,In_206);
or U297 (N_297,In_437,In_78);
nor U298 (N_298,In_267,In_280);
and U299 (N_299,In_238,In_256);
nor U300 (N_300,In_186,In_461);
xnor U301 (N_301,In_357,In_106);
nor U302 (N_302,In_419,In_19);
nor U303 (N_303,In_387,In_432);
and U304 (N_304,In_159,In_368);
or U305 (N_305,In_149,In_375);
and U306 (N_306,In_207,In_168);
nor U307 (N_307,In_88,In_332);
or U308 (N_308,In_286,In_319);
or U309 (N_309,In_21,In_330);
or U310 (N_310,In_336,In_250);
and U311 (N_311,In_112,In_102);
or U312 (N_312,In_289,In_58);
or U313 (N_313,In_190,In_427);
xnor U314 (N_314,In_33,In_150);
nand U315 (N_315,In_401,In_407);
nand U316 (N_316,In_426,In_459);
or U317 (N_317,In_157,In_143);
nor U318 (N_318,In_176,In_174);
nand U319 (N_319,In_50,In_196);
and U320 (N_320,In_408,In_107);
or U321 (N_321,In_369,In_431);
nand U322 (N_322,In_242,In_485);
xor U323 (N_323,In_382,In_133);
nor U324 (N_324,In_9,In_348);
or U325 (N_325,In_157,In_12);
or U326 (N_326,In_150,In_375);
and U327 (N_327,In_84,In_192);
and U328 (N_328,In_116,In_279);
and U329 (N_329,In_12,In_213);
nor U330 (N_330,In_242,In_257);
and U331 (N_331,In_403,In_458);
and U332 (N_332,In_24,In_22);
nand U333 (N_333,In_411,In_357);
and U334 (N_334,In_79,In_410);
nor U335 (N_335,In_242,In_166);
nor U336 (N_336,In_30,In_160);
nand U337 (N_337,In_119,In_102);
and U338 (N_338,In_239,In_400);
nor U339 (N_339,In_344,In_52);
nor U340 (N_340,In_97,In_206);
nor U341 (N_341,In_403,In_303);
or U342 (N_342,In_166,In_73);
and U343 (N_343,In_78,In_82);
and U344 (N_344,In_143,In_493);
nand U345 (N_345,In_254,In_288);
or U346 (N_346,In_309,In_377);
nand U347 (N_347,In_370,In_216);
nand U348 (N_348,In_337,In_307);
and U349 (N_349,In_62,In_182);
or U350 (N_350,In_143,In_288);
or U351 (N_351,In_354,In_315);
nor U352 (N_352,In_143,In_244);
nor U353 (N_353,In_193,In_272);
nor U354 (N_354,In_479,In_4);
nand U355 (N_355,In_444,In_408);
nand U356 (N_356,In_205,In_293);
nor U357 (N_357,In_189,In_371);
nand U358 (N_358,In_169,In_233);
nor U359 (N_359,In_495,In_326);
or U360 (N_360,In_151,In_83);
or U361 (N_361,In_353,In_63);
and U362 (N_362,In_331,In_106);
or U363 (N_363,In_61,In_333);
nor U364 (N_364,In_180,In_61);
xnor U365 (N_365,In_257,In_111);
nand U366 (N_366,In_126,In_197);
or U367 (N_367,In_37,In_94);
nand U368 (N_368,In_201,In_325);
or U369 (N_369,In_412,In_402);
nand U370 (N_370,In_266,In_322);
nand U371 (N_371,In_171,In_394);
nor U372 (N_372,In_72,In_106);
and U373 (N_373,In_471,In_492);
or U374 (N_374,In_347,In_6);
and U375 (N_375,In_34,In_225);
nor U376 (N_376,In_411,In_166);
nor U377 (N_377,In_80,In_397);
nor U378 (N_378,In_471,In_212);
and U379 (N_379,In_370,In_250);
nor U380 (N_380,In_260,In_194);
and U381 (N_381,In_113,In_187);
xor U382 (N_382,In_144,In_90);
or U383 (N_383,In_143,In_55);
nand U384 (N_384,In_418,In_389);
and U385 (N_385,In_55,In_261);
or U386 (N_386,In_445,In_35);
and U387 (N_387,In_290,In_346);
or U388 (N_388,In_279,In_299);
nand U389 (N_389,In_230,In_350);
nand U390 (N_390,In_116,In_406);
and U391 (N_391,In_64,In_252);
nor U392 (N_392,In_40,In_383);
nand U393 (N_393,In_52,In_407);
nand U394 (N_394,In_325,In_100);
or U395 (N_395,In_92,In_383);
and U396 (N_396,In_99,In_407);
nor U397 (N_397,In_41,In_389);
and U398 (N_398,In_445,In_232);
or U399 (N_399,In_265,In_355);
and U400 (N_400,In_63,In_81);
nor U401 (N_401,In_267,In_194);
nor U402 (N_402,In_145,In_94);
xnor U403 (N_403,In_170,In_339);
nor U404 (N_404,In_285,In_326);
nand U405 (N_405,In_306,In_162);
or U406 (N_406,In_485,In_244);
or U407 (N_407,In_378,In_430);
or U408 (N_408,In_237,In_22);
nor U409 (N_409,In_238,In_106);
or U410 (N_410,In_299,In_458);
xor U411 (N_411,In_422,In_93);
nand U412 (N_412,In_127,In_346);
nand U413 (N_413,In_103,In_144);
nor U414 (N_414,In_4,In_1);
or U415 (N_415,In_114,In_146);
nand U416 (N_416,In_58,In_445);
xnor U417 (N_417,In_137,In_113);
nor U418 (N_418,In_193,In_431);
nor U419 (N_419,In_303,In_72);
xnor U420 (N_420,In_79,In_437);
nand U421 (N_421,In_182,In_261);
and U422 (N_422,In_406,In_31);
nand U423 (N_423,In_191,In_331);
or U424 (N_424,In_134,In_272);
or U425 (N_425,In_213,In_233);
or U426 (N_426,In_297,In_474);
nand U427 (N_427,In_258,In_366);
nand U428 (N_428,In_364,In_195);
and U429 (N_429,In_187,In_413);
and U430 (N_430,In_155,In_454);
nand U431 (N_431,In_292,In_132);
nand U432 (N_432,In_366,In_422);
nor U433 (N_433,In_283,In_250);
or U434 (N_434,In_352,In_343);
and U435 (N_435,In_194,In_72);
nand U436 (N_436,In_119,In_219);
or U437 (N_437,In_69,In_173);
or U438 (N_438,In_188,In_440);
nand U439 (N_439,In_483,In_238);
and U440 (N_440,In_309,In_166);
or U441 (N_441,In_226,In_411);
nor U442 (N_442,In_213,In_466);
and U443 (N_443,In_33,In_325);
or U444 (N_444,In_213,In_48);
nand U445 (N_445,In_151,In_120);
nor U446 (N_446,In_305,In_116);
and U447 (N_447,In_491,In_112);
and U448 (N_448,In_417,In_197);
nand U449 (N_449,In_0,In_161);
nand U450 (N_450,In_35,In_337);
nor U451 (N_451,In_368,In_148);
or U452 (N_452,In_197,In_410);
nor U453 (N_453,In_296,In_231);
nand U454 (N_454,In_286,In_453);
nand U455 (N_455,In_300,In_167);
or U456 (N_456,In_179,In_389);
nor U457 (N_457,In_468,In_283);
or U458 (N_458,In_146,In_1);
xor U459 (N_459,In_467,In_333);
and U460 (N_460,In_494,In_32);
or U461 (N_461,In_290,In_236);
or U462 (N_462,In_20,In_158);
xor U463 (N_463,In_40,In_170);
nor U464 (N_464,In_21,In_6);
or U465 (N_465,In_457,In_132);
xnor U466 (N_466,In_59,In_62);
nand U467 (N_467,In_244,In_412);
nand U468 (N_468,In_314,In_472);
xor U469 (N_469,In_390,In_2);
or U470 (N_470,In_354,In_16);
nand U471 (N_471,In_487,In_201);
nand U472 (N_472,In_394,In_409);
nor U473 (N_473,In_77,In_46);
and U474 (N_474,In_6,In_59);
or U475 (N_475,In_476,In_162);
nor U476 (N_476,In_130,In_400);
xnor U477 (N_477,In_286,In_192);
or U478 (N_478,In_353,In_300);
and U479 (N_479,In_116,In_201);
or U480 (N_480,In_187,In_10);
nor U481 (N_481,In_285,In_200);
or U482 (N_482,In_26,In_53);
nor U483 (N_483,In_439,In_398);
and U484 (N_484,In_375,In_282);
nor U485 (N_485,In_20,In_85);
nor U486 (N_486,In_147,In_241);
nor U487 (N_487,In_467,In_233);
and U488 (N_488,In_381,In_70);
and U489 (N_489,In_429,In_84);
nor U490 (N_490,In_130,In_490);
and U491 (N_491,In_274,In_356);
and U492 (N_492,In_188,In_406);
and U493 (N_493,In_144,In_411);
or U494 (N_494,In_253,In_474);
or U495 (N_495,In_444,In_15);
nor U496 (N_496,In_101,In_210);
nor U497 (N_497,In_23,In_158);
nand U498 (N_498,In_1,In_161);
or U499 (N_499,In_92,In_428);
xnor U500 (N_500,In_252,In_387);
nor U501 (N_501,In_402,In_455);
nand U502 (N_502,In_177,In_100);
nor U503 (N_503,In_270,In_445);
and U504 (N_504,In_197,In_492);
nand U505 (N_505,In_235,In_154);
nand U506 (N_506,In_373,In_462);
and U507 (N_507,In_6,In_92);
and U508 (N_508,In_269,In_340);
xor U509 (N_509,In_431,In_25);
or U510 (N_510,In_123,In_364);
and U511 (N_511,In_448,In_56);
nor U512 (N_512,In_38,In_139);
or U513 (N_513,In_281,In_13);
nand U514 (N_514,In_440,In_190);
or U515 (N_515,In_94,In_479);
nand U516 (N_516,In_121,In_444);
nor U517 (N_517,In_49,In_372);
nand U518 (N_518,In_488,In_161);
and U519 (N_519,In_2,In_492);
nor U520 (N_520,In_170,In_465);
nand U521 (N_521,In_184,In_52);
nand U522 (N_522,In_107,In_294);
nor U523 (N_523,In_478,In_322);
and U524 (N_524,In_100,In_200);
and U525 (N_525,In_193,In_263);
and U526 (N_526,In_215,In_124);
nor U527 (N_527,In_296,In_248);
nand U528 (N_528,In_49,In_214);
nor U529 (N_529,In_397,In_398);
xnor U530 (N_530,In_407,In_452);
nor U531 (N_531,In_275,In_208);
nand U532 (N_532,In_214,In_154);
and U533 (N_533,In_195,In_137);
xnor U534 (N_534,In_292,In_370);
xnor U535 (N_535,In_146,In_240);
nor U536 (N_536,In_117,In_377);
or U537 (N_537,In_240,In_407);
and U538 (N_538,In_355,In_264);
and U539 (N_539,In_83,In_144);
xor U540 (N_540,In_380,In_403);
or U541 (N_541,In_178,In_50);
nor U542 (N_542,In_465,In_137);
or U543 (N_543,In_53,In_370);
nand U544 (N_544,In_12,In_391);
and U545 (N_545,In_115,In_134);
and U546 (N_546,In_308,In_290);
nand U547 (N_547,In_308,In_180);
or U548 (N_548,In_406,In_24);
or U549 (N_549,In_64,In_109);
nor U550 (N_550,In_234,In_51);
nand U551 (N_551,In_39,In_126);
and U552 (N_552,In_343,In_106);
and U553 (N_553,In_84,In_147);
xnor U554 (N_554,In_304,In_494);
or U555 (N_555,In_133,In_373);
and U556 (N_556,In_261,In_452);
xor U557 (N_557,In_341,In_63);
or U558 (N_558,In_302,In_339);
nand U559 (N_559,In_255,In_5);
or U560 (N_560,In_461,In_441);
and U561 (N_561,In_403,In_297);
and U562 (N_562,In_117,In_91);
or U563 (N_563,In_112,In_27);
nand U564 (N_564,In_252,In_300);
or U565 (N_565,In_155,In_18);
nand U566 (N_566,In_29,In_86);
or U567 (N_567,In_99,In_161);
or U568 (N_568,In_336,In_486);
nand U569 (N_569,In_429,In_55);
or U570 (N_570,In_474,In_325);
or U571 (N_571,In_352,In_480);
and U572 (N_572,In_2,In_79);
and U573 (N_573,In_333,In_93);
nor U574 (N_574,In_243,In_196);
or U575 (N_575,In_298,In_91);
nand U576 (N_576,In_360,In_17);
nand U577 (N_577,In_163,In_313);
xor U578 (N_578,In_259,In_93);
and U579 (N_579,In_241,In_483);
nor U580 (N_580,In_162,In_404);
and U581 (N_581,In_379,In_423);
nand U582 (N_582,In_216,In_359);
nor U583 (N_583,In_409,In_71);
nor U584 (N_584,In_214,In_403);
or U585 (N_585,In_253,In_43);
nand U586 (N_586,In_134,In_269);
nor U587 (N_587,In_14,In_7);
nor U588 (N_588,In_205,In_167);
and U589 (N_589,In_440,In_240);
and U590 (N_590,In_145,In_379);
nand U591 (N_591,In_328,In_350);
nand U592 (N_592,In_136,In_213);
nor U593 (N_593,In_324,In_130);
nor U594 (N_594,In_465,In_293);
xor U595 (N_595,In_16,In_161);
nand U596 (N_596,In_371,In_240);
and U597 (N_597,In_408,In_96);
nor U598 (N_598,In_372,In_327);
and U599 (N_599,In_344,In_390);
and U600 (N_600,In_14,In_247);
and U601 (N_601,In_364,In_3);
and U602 (N_602,In_244,In_219);
nand U603 (N_603,In_360,In_458);
nand U604 (N_604,In_485,In_359);
xnor U605 (N_605,In_168,In_136);
or U606 (N_606,In_416,In_201);
nand U607 (N_607,In_196,In_386);
or U608 (N_608,In_37,In_179);
xnor U609 (N_609,In_143,In_128);
nor U610 (N_610,In_331,In_35);
or U611 (N_611,In_330,In_388);
and U612 (N_612,In_147,In_126);
xor U613 (N_613,In_457,In_312);
nor U614 (N_614,In_331,In_117);
or U615 (N_615,In_229,In_243);
and U616 (N_616,In_44,In_52);
xnor U617 (N_617,In_299,In_389);
nand U618 (N_618,In_463,In_79);
nor U619 (N_619,In_43,In_36);
and U620 (N_620,In_17,In_490);
and U621 (N_621,In_402,In_173);
and U622 (N_622,In_35,In_471);
and U623 (N_623,In_88,In_240);
or U624 (N_624,In_383,In_419);
nor U625 (N_625,In_21,In_411);
or U626 (N_626,In_79,In_377);
xnor U627 (N_627,In_203,In_426);
or U628 (N_628,In_239,In_356);
and U629 (N_629,In_158,In_187);
nand U630 (N_630,In_167,In_362);
nand U631 (N_631,In_125,In_31);
nand U632 (N_632,In_49,In_263);
and U633 (N_633,In_61,In_259);
or U634 (N_634,In_376,In_143);
nor U635 (N_635,In_50,In_254);
xnor U636 (N_636,In_248,In_128);
and U637 (N_637,In_230,In_295);
and U638 (N_638,In_365,In_171);
nand U639 (N_639,In_433,In_157);
or U640 (N_640,In_112,In_106);
and U641 (N_641,In_66,In_218);
nand U642 (N_642,In_223,In_145);
and U643 (N_643,In_425,In_366);
nor U644 (N_644,In_439,In_24);
nor U645 (N_645,In_98,In_471);
nor U646 (N_646,In_65,In_417);
nand U647 (N_647,In_81,In_87);
nor U648 (N_648,In_342,In_315);
or U649 (N_649,In_51,In_139);
nor U650 (N_650,In_493,In_38);
nand U651 (N_651,In_130,In_445);
and U652 (N_652,In_267,In_158);
xor U653 (N_653,In_496,In_279);
and U654 (N_654,In_271,In_365);
and U655 (N_655,In_128,In_206);
and U656 (N_656,In_272,In_384);
nand U657 (N_657,In_426,In_387);
nand U658 (N_658,In_94,In_293);
nand U659 (N_659,In_204,In_431);
nand U660 (N_660,In_84,In_491);
and U661 (N_661,In_262,In_410);
nor U662 (N_662,In_303,In_107);
xor U663 (N_663,In_63,In_163);
xnor U664 (N_664,In_20,In_292);
and U665 (N_665,In_400,In_129);
and U666 (N_666,In_179,In_129);
xnor U667 (N_667,In_222,In_413);
nor U668 (N_668,In_396,In_189);
nor U669 (N_669,In_251,In_19);
nand U670 (N_670,In_223,In_324);
or U671 (N_671,In_119,In_5);
and U672 (N_672,In_80,In_458);
nor U673 (N_673,In_291,In_300);
nor U674 (N_674,In_200,In_126);
nor U675 (N_675,In_396,In_37);
nor U676 (N_676,In_237,In_27);
nand U677 (N_677,In_231,In_8);
and U678 (N_678,In_337,In_11);
nor U679 (N_679,In_414,In_193);
nor U680 (N_680,In_107,In_167);
nand U681 (N_681,In_96,In_196);
and U682 (N_682,In_413,In_480);
or U683 (N_683,In_175,In_384);
nor U684 (N_684,In_431,In_332);
or U685 (N_685,In_249,In_419);
or U686 (N_686,In_413,In_411);
nand U687 (N_687,In_380,In_454);
nor U688 (N_688,In_219,In_447);
or U689 (N_689,In_203,In_421);
nor U690 (N_690,In_381,In_353);
nand U691 (N_691,In_395,In_13);
nand U692 (N_692,In_199,In_132);
nand U693 (N_693,In_437,In_119);
nor U694 (N_694,In_158,In_69);
nor U695 (N_695,In_16,In_48);
or U696 (N_696,In_367,In_172);
nand U697 (N_697,In_138,In_299);
nor U698 (N_698,In_322,In_148);
or U699 (N_699,In_242,In_404);
nand U700 (N_700,In_325,In_249);
or U701 (N_701,In_131,In_477);
or U702 (N_702,In_139,In_320);
and U703 (N_703,In_231,In_381);
or U704 (N_704,In_330,In_359);
nand U705 (N_705,In_123,In_368);
nand U706 (N_706,In_431,In_304);
or U707 (N_707,In_288,In_491);
and U708 (N_708,In_132,In_230);
nand U709 (N_709,In_304,In_337);
or U710 (N_710,In_193,In_310);
nor U711 (N_711,In_211,In_74);
or U712 (N_712,In_394,In_15);
and U713 (N_713,In_116,In_435);
nand U714 (N_714,In_376,In_13);
and U715 (N_715,In_470,In_275);
or U716 (N_716,In_33,In_345);
nand U717 (N_717,In_227,In_445);
and U718 (N_718,In_58,In_385);
nor U719 (N_719,In_113,In_89);
and U720 (N_720,In_57,In_401);
and U721 (N_721,In_319,In_243);
nor U722 (N_722,In_2,In_284);
nand U723 (N_723,In_334,In_484);
nor U724 (N_724,In_277,In_357);
nand U725 (N_725,In_120,In_345);
nor U726 (N_726,In_193,In_336);
or U727 (N_727,In_370,In_84);
nor U728 (N_728,In_309,In_170);
or U729 (N_729,In_379,In_422);
xor U730 (N_730,In_50,In_117);
nor U731 (N_731,In_48,In_401);
nand U732 (N_732,In_409,In_3);
or U733 (N_733,In_241,In_101);
and U734 (N_734,In_482,In_436);
nor U735 (N_735,In_232,In_299);
xor U736 (N_736,In_398,In_261);
or U737 (N_737,In_305,In_295);
or U738 (N_738,In_408,In_295);
nor U739 (N_739,In_132,In_109);
and U740 (N_740,In_219,In_387);
or U741 (N_741,In_292,In_22);
nand U742 (N_742,In_129,In_430);
nand U743 (N_743,In_307,In_121);
nand U744 (N_744,In_294,In_397);
xnor U745 (N_745,In_52,In_19);
or U746 (N_746,In_8,In_410);
and U747 (N_747,In_229,In_219);
nor U748 (N_748,In_45,In_28);
xor U749 (N_749,In_243,In_388);
nor U750 (N_750,N_541,N_248);
and U751 (N_751,N_285,N_196);
nor U752 (N_752,N_145,N_165);
and U753 (N_753,N_202,N_233);
or U754 (N_754,N_289,N_504);
nand U755 (N_755,N_444,N_224);
xor U756 (N_756,N_727,N_589);
xnor U757 (N_757,N_572,N_602);
nand U758 (N_758,N_477,N_743);
or U759 (N_759,N_489,N_84);
and U760 (N_760,N_734,N_671);
and U761 (N_761,N_140,N_95);
and U762 (N_762,N_211,N_388);
and U763 (N_763,N_736,N_520);
or U764 (N_764,N_551,N_240);
nor U765 (N_765,N_10,N_218);
or U766 (N_766,N_630,N_176);
or U767 (N_767,N_302,N_507);
or U768 (N_768,N_369,N_535);
xor U769 (N_769,N_310,N_144);
or U770 (N_770,N_215,N_604);
nand U771 (N_771,N_665,N_637);
or U772 (N_772,N_282,N_299);
nand U773 (N_773,N_22,N_413);
nor U774 (N_774,N_314,N_415);
or U775 (N_775,N_169,N_78);
or U776 (N_776,N_168,N_505);
nand U777 (N_777,N_385,N_228);
or U778 (N_778,N_308,N_737);
nand U779 (N_779,N_153,N_182);
or U780 (N_780,N_405,N_493);
and U781 (N_781,N_105,N_148);
nand U782 (N_782,N_594,N_568);
and U783 (N_783,N_300,N_36);
and U784 (N_784,N_728,N_287);
and U785 (N_785,N_690,N_217);
xnor U786 (N_786,N_673,N_348);
xor U787 (N_787,N_487,N_279);
and U788 (N_788,N_375,N_509);
xor U789 (N_789,N_591,N_376);
and U790 (N_790,N_7,N_267);
or U791 (N_791,N_398,N_523);
nand U792 (N_792,N_648,N_281);
nand U793 (N_793,N_212,N_409);
nor U794 (N_794,N_1,N_570);
and U795 (N_795,N_117,N_81);
nor U796 (N_796,N_463,N_599);
nor U797 (N_797,N_465,N_296);
or U798 (N_798,N_94,N_685);
nand U799 (N_799,N_596,N_155);
or U800 (N_800,N_692,N_198);
and U801 (N_801,N_163,N_587);
or U802 (N_802,N_634,N_435);
nor U803 (N_803,N_738,N_357);
xor U804 (N_804,N_120,N_46);
nand U805 (N_805,N_735,N_622);
nand U806 (N_806,N_683,N_749);
or U807 (N_807,N_266,N_733);
and U808 (N_808,N_386,N_460);
nor U809 (N_809,N_380,N_701);
or U810 (N_810,N_66,N_558);
nor U811 (N_811,N_331,N_152);
nor U812 (N_812,N_70,N_53);
nand U813 (N_813,N_724,N_542);
nor U814 (N_814,N_134,N_639);
nor U815 (N_815,N_329,N_499);
xnor U816 (N_816,N_87,N_355);
nand U817 (N_817,N_723,N_434);
and U818 (N_818,N_108,N_421);
or U819 (N_819,N_617,N_312);
xnor U820 (N_820,N_40,N_318);
xnor U821 (N_821,N_137,N_748);
and U822 (N_822,N_691,N_132);
and U823 (N_823,N_255,N_26);
nor U824 (N_824,N_631,N_326);
nand U825 (N_825,N_472,N_112);
xor U826 (N_826,N_585,N_107);
nor U827 (N_827,N_88,N_82);
or U828 (N_828,N_554,N_346);
nand U829 (N_829,N_330,N_401);
or U830 (N_830,N_470,N_223);
or U831 (N_831,N_426,N_588);
or U832 (N_832,N_616,N_33);
nand U833 (N_833,N_361,N_216);
or U834 (N_834,N_263,N_127);
nand U835 (N_835,N_44,N_500);
nor U836 (N_836,N_49,N_313);
nand U837 (N_837,N_320,N_553);
nand U838 (N_838,N_130,N_632);
nand U839 (N_839,N_442,N_580);
nor U840 (N_840,N_670,N_52);
nand U841 (N_841,N_277,N_220);
and U842 (N_842,N_422,N_75);
nor U843 (N_843,N_534,N_412);
nand U844 (N_844,N_204,N_529);
or U845 (N_845,N_337,N_304);
xor U846 (N_846,N_328,N_322);
nand U847 (N_847,N_103,N_272);
nor U848 (N_848,N_62,N_582);
xor U849 (N_849,N_124,N_700);
nor U850 (N_850,N_403,N_370);
nand U851 (N_851,N_703,N_48);
and U852 (N_852,N_364,N_129);
and U853 (N_853,N_239,N_14);
xor U854 (N_854,N_192,N_543);
and U855 (N_855,N_180,N_41);
and U856 (N_856,N_595,N_419);
nor U857 (N_857,N_525,N_186);
and U858 (N_858,N_25,N_447);
nor U859 (N_859,N_90,N_571);
or U860 (N_860,N_390,N_86);
or U861 (N_861,N_417,N_485);
and U862 (N_862,N_92,N_63);
and U863 (N_863,N_338,N_37);
nand U864 (N_864,N_236,N_677);
or U865 (N_865,N_600,N_423);
xnor U866 (N_866,N_546,N_650);
nor U867 (N_867,N_544,N_77);
and U868 (N_868,N_657,N_626);
or U869 (N_869,N_190,N_275);
or U870 (N_870,N_540,N_245);
nor U871 (N_871,N_478,N_147);
nor U872 (N_872,N_290,N_379);
xnor U873 (N_873,N_327,N_511);
and U874 (N_874,N_150,N_432);
nor U875 (N_875,N_722,N_424);
and U876 (N_876,N_642,N_383);
and U877 (N_877,N_252,N_425);
nand U878 (N_878,N_476,N_698);
xnor U879 (N_879,N_658,N_539);
or U880 (N_880,N_619,N_11);
or U881 (N_881,N_611,N_199);
and U882 (N_882,N_537,N_552);
or U883 (N_883,N_297,N_638);
or U884 (N_884,N_454,N_60);
nor U885 (N_885,N_271,N_237);
nand U886 (N_886,N_747,N_406);
nor U887 (N_887,N_185,N_740);
nand U888 (N_888,N_362,N_16);
nor U889 (N_889,N_446,N_621);
and U890 (N_890,N_342,N_100);
and U891 (N_891,N_394,N_227);
and U892 (N_892,N_651,N_73);
and U893 (N_893,N_433,N_118);
and U894 (N_894,N_506,N_166);
nor U895 (N_895,N_503,N_704);
or U896 (N_896,N_324,N_254);
nor U897 (N_897,N_384,N_280);
nand U898 (N_898,N_54,N_106);
nand U899 (N_899,N_162,N_353);
nand U900 (N_900,N_56,N_354);
or U901 (N_901,N_514,N_85);
nor U902 (N_902,N_668,N_494);
nand U903 (N_903,N_205,N_68);
nand U904 (N_904,N_65,N_456);
or U905 (N_905,N_177,N_656);
nand U906 (N_906,N_556,N_193);
nand U907 (N_907,N_512,N_625);
nor U908 (N_908,N_241,N_74);
nor U909 (N_909,N_0,N_713);
and U910 (N_910,N_586,N_437);
nand U911 (N_911,N_675,N_4);
nand U912 (N_912,N_45,N_203);
nand U913 (N_913,N_680,N_262);
nor U914 (N_914,N_726,N_57);
nor U915 (N_915,N_699,N_19);
or U916 (N_916,N_530,N_410);
or U917 (N_917,N_209,N_400);
and U918 (N_918,N_416,N_455);
and U919 (N_919,N_628,N_559);
nand U920 (N_920,N_560,N_715);
or U921 (N_921,N_532,N_238);
xnor U922 (N_922,N_366,N_207);
nor U923 (N_923,N_496,N_573);
nand U924 (N_924,N_574,N_678);
and U925 (N_925,N_276,N_578);
nor U926 (N_926,N_261,N_428);
and U927 (N_927,N_119,N_109);
or U928 (N_928,N_623,N_381);
or U929 (N_929,N_194,N_491);
xnor U930 (N_930,N_206,N_635);
nand U931 (N_931,N_646,N_319);
nand U932 (N_932,N_468,N_116);
and U933 (N_933,N_718,N_32);
or U934 (N_934,N_295,N_633);
and U935 (N_935,N_647,N_521);
nand U936 (N_936,N_110,N_563);
or U937 (N_937,N_59,N_242);
nand U938 (N_938,N_243,N_244);
nor U939 (N_939,N_641,N_609);
nor U940 (N_940,N_79,N_681);
nand U941 (N_941,N_502,N_482);
nand U942 (N_942,N_663,N_284);
or U943 (N_943,N_114,N_99);
nor U944 (N_944,N_122,N_689);
xnor U945 (N_945,N_184,N_745);
and U946 (N_946,N_89,N_712);
nand U947 (N_947,N_93,N_246);
nor U948 (N_948,N_360,N_195);
or U949 (N_949,N_576,N_21);
and U950 (N_950,N_50,N_682);
nand U951 (N_951,N_363,N_181);
xnor U952 (N_952,N_259,N_501);
nor U953 (N_953,N_159,N_654);
nor U954 (N_954,N_707,N_598);
nor U955 (N_955,N_717,N_133);
nand U956 (N_956,N_368,N_336);
xnor U957 (N_957,N_377,N_136);
nor U958 (N_958,N_160,N_76);
or U959 (N_959,N_288,N_229);
nor U960 (N_960,N_28,N_549);
nor U961 (N_961,N_349,N_567);
or U962 (N_962,N_666,N_323);
and U963 (N_963,N_102,N_725);
and U964 (N_964,N_438,N_164);
nor U965 (N_965,N_614,N_339);
nor U966 (N_966,N_58,N_581);
nand U967 (N_967,N_524,N_694);
or U968 (N_968,N_676,N_513);
xnor U969 (N_969,N_325,N_200);
or U970 (N_970,N_382,N_12);
nor U971 (N_971,N_387,N_292);
and U972 (N_972,N_457,N_464);
and U973 (N_973,N_389,N_96);
and U974 (N_974,N_146,N_575);
nor U975 (N_975,N_706,N_605);
xnor U976 (N_976,N_13,N_729);
nand U977 (N_977,N_309,N_606);
nand U978 (N_978,N_555,N_175);
or U979 (N_979,N_693,N_347);
xnor U980 (N_980,N_142,N_436);
and U981 (N_981,N_561,N_115);
nor U982 (N_982,N_174,N_125);
nor U983 (N_983,N_445,N_643);
nand U984 (N_984,N_18,N_67);
and U985 (N_985,N_101,N_51);
nor U986 (N_986,N_492,N_564);
nor U987 (N_987,N_592,N_474);
xor U988 (N_988,N_538,N_340);
nand U989 (N_989,N_188,N_332);
nand U990 (N_990,N_257,N_526);
nand U991 (N_991,N_480,N_247);
and U992 (N_992,N_143,N_427);
and U993 (N_993,N_311,N_629);
or U994 (N_994,N_20,N_550);
or U995 (N_995,N_226,N_395);
nor U996 (N_996,N_321,N_178);
or U997 (N_997,N_141,N_61);
nand U998 (N_998,N_627,N_443);
or U999 (N_999,N_30,N_131);
and U1000 (N_1000,N_579,N_516);
nor U1001 (N_1001,N_431,N_655);
or U1002 (N_1002,N_372,N_291);
nor U1003 (N_1003,N_149,N_352);
nor U1004 (N_1004,N_15,N_171);
or U1005 (N_1005,N_545,N_221);
or U1006 (N_1006,N_730,N_705);
nor U1007 (N_1007,N_157,N_31);
nand U1008 (N_1008,N_222,N_613);
nor U1009 (N_1009,N_333,N_98);
nand U1010 (N_1010,N_104,N_123);
or U1011 (N_1011,N_6,N_294);
nand U1012 (N_1012,N_138,N_404);
or U1013 (N_1013,N_742,N_660);
xor U1014 (N_1014,N_91,N_721);
or U1015 (N_1015,N_548,N_172);
nand U1016 (N_1016,N_43,N_620);
or U1017 (N_1017,N_597,N_695);
and U1018 (N_1018,N_231,N_430);
nand U1019 (N_1019,N_283,N_429);
or U1020 (N_1020,N_47,N_508);
xor U1021 (N_1021,N_306,N_462);
or U1022 (N_1022,N_459,N_714);
or U1023 (N_1023,N_270,N_659);
nand U1024 (N_1024,N_744,N_527);
nand U1025 (N_1025,N_256,N_481);
nand U1026 (N_1026,N_497,N_316);
and U1027 (N_1027,N_38,N_391);
nand U1028 (N_1028,N_378,N_732);
and U1029 (N_1029,N_286,N_536);
or U1030 (N_1030,N_479,N_187);
and U1031 (N_1031,N_615,N_402);
and U1032 (N_1032,N_518,N_746);
or U1033 (N_1033,N_709,N_126);
and U1034 (N_1034,N_315,N_225);
nand U1035 (N_1035,N_197,N_664);
or U1036 (N_1036,N_461,N_121);
and U1037 (N_1037,N_640,N_161);
nand U1038 (N_1038,N_686,N_250);
or U1039 (N_1039,N_618,N_399);
and U1040 (N_1040,N_2,N_716);
or U1041 (N_1041,N_469,N_533);
nand U1042 (N_1042,N_167,N_359);
and U1043 (N_1043,N_343,N_158);
xor U1044 (N_1044,N_374,N_358);
nand U1045 (N_1045,N_213,N_498);
nand U1046 (N_1046,N_420,N_293);
xor U1047 (N_1047,N_557,N_9);
nand U1048 (N_1048,N_230,N_335);
or U1049 (N_1049,N_269,N_475);
or U1050 (N_1050,N_562,N_232);
and U1051 (N_1051,N_264,N_128);
or U1052 (N_1052,N_607,N_189);
nand U1053 (N_1053,N_590,N_34);
xor U1054 (N_1054,N_486,N_8);
nand U1055 (N_1055,N_179,N_397);
or U1056 (N_1056,N_111,N_392);
and U1057 (N_1057,N_139,N_356);
or U1058 (N_1058,N_69,N_24);
xnor U1059 (N_1059,N_303,N_42);
or U1060 (N_1060,N_739,N_97);
nand U1061 (N_1061,N_696,N_334);
nand U1062 (N_1062,N_408,N_510);
nor U1063 (N_1063,N_577,N_83);
or U1064 (N_1064,N_55,N_684);
xor U1065 (N_1065,N_731,N_64);
nor U1066 (N_1066,N_448,N_667);
or U1067 (N_1067,N_365,N_547);
and U1068 (N_1068,N_584,N_407);
nand U1069 (N_1069,N_608,N_583);
and U1070 (N_1070,N_495,N_687);
or U1071 (N_1071,N_636,N_260);
xor U1072 (N_1072,N_234,N_273);
and U1073 (N_1073,N_235,N_531);
nand U1074 (N_1074,N_569,N_317);
or U1075 (N_1075,N_307,N_17);
nand U1076 (N_1076,N_305,N_515);
or U1077 (N_1077,N_344,N_483);
and U1078 (N_1078,N_214,N_458);
or U1079 (N_1079,N_719,N_345);
xor U1080 (N_1080,N_27,N_414);
nand U1081 (N_1081,N_441,N_249);
nand U1082 (N_1082,N_439,N_528);
nand U1083 (N_1083,N_624,N_210);
or U1084 (N_1084,N_490,N_173);
nor U1085 (N_1085,N_373,N_672);
and U1086 (N_1086,N_29,N_350);
or U1087 (N_1087,N_697,N_80);
or U1088 (N_1088,N_201,N_471);
xor U1089 (N_1089,N_522,N_156);
nand U1090 (N_1090,N_467,N_3);
or U1091 (N_1091,N_612,N_151);
or U1092 (N_1092,N_488,N_278);
nor U1093 (N_1093,N_5,N_39);
and U1094 (N_1094,N_661,N_451);
and U1095 (N_1095,N_452,N_720);
and U1096 (N_1096,N_440,N_711);
nor U1097 (N_1097,N_265,N_274);
and U1098 (N_1098,N_593,N_708);
nand U1099 (N_1099,N_396,N_453);
and U1100 (N_1100,N_35,N_418);
xor U1101 (N_1101,N_298,N_484);
nand U1102 (N_1102,N_258,N_351);
nand U1103 (N_1103,N_702,N_517);
or U1104 (N_1104,N_610,N_411);
nand U1105 (N_1105,N_450,N_741);
nand U1106 (N_1106,N_649,N_253);
nand U1107 (N_1107,N_183,N_393);
or U1108 (N_1108,N_72,N_449);
xor U1109 (N_1109,N_644,N_601);
nor U1110 (N_1110,N_653,N_688);
or U1111 (N_1111,N_135,N_23);
nor U1112 (N_1112,N_566,N_662);
xor U1113 (N_1113,N_669,N_191);
and U1114 (N_1114,N_466,N_652);
xnor U1115 (N_1115,N_341,N_268);
or U1116 (N_1116,N_603,N_674);
xor U1117 (N_1117,N_170,N_645);
or U1118 (N_1118,N_71,N_473);
or U1119 (N_1119,N_371,N_519);
or U1120 (N_1120,N_113,N_251);
nand U1121 (N_1121,N_367,N_565);
nor U1122 (N_1122,N_208,N_710);
nand U1123 (N_1123,N_301,N_154);
nor U1124 (N_1124,N_219,N_679);
nand U1125 (N_1125,N_291,N_287);
nand U1126 (N_1126,N_469,N_311);
or U1127 (N_1127,N_226,N_16);
nand U1128 (N_1128,N_390,N_645);
and U1129 (N_1129,N_482,N_422);
or U1130 (N_1130,N_567,N_641);
xnor U1131 (N_1131,N_279,N_703);
xnor U1132 (N_1132,N_306,N_394);
nand U1133 (N_1133,N_175,N_171);
nand U1134 (N_1134,N_420,N_257);
nor U1135 (N_1135,N_278,N_612);
xor U1136 (N_1136,N_643,N_76);
and U1137 (N_1137,N_197,N_534);
nor U1138 (N_1138,N_29,N_554);
nor U1139 (N_1139,N_146,N_112);
or U1140 (N_1140,N_318,N_500);
and U1141 (N_1141,N_349,N_697);
nor U1142 (N_1142,N_558,N_414);
xor U1143 (N_1143,N_232,N_25);
or U1144 (N_1144,N_699,N_257);
and U1145 (N_1145,N_40,N_593);
xnor U1146 (N_1146,N_112,N_292);
nor U1147 (N_1147,N_470,N_221);
nor U1148 (N_1148,N_352,N_287);
and U1149 (N_1149,N_450,N_388);
nor U1150 (N_1150,N_270,N_80);
or U1151 (N_1151,N_409,N_139);
or U1152 (N_1152,N_280,N_737);
xnor U1153 (N_1153,N_572,N_427);
or U1154 (N_1154,N_469,N_15);
and U1155 (N_1155,N_33,N_412);
nand U1156 (N_1156,N_91,N_79);
or U1157 (N_1157,N_256,N_603);
nand U1158 (N_1158,N_71,N_70);
nand U1159 (N_1159,N_405,N_105);
xor U1160 (N_1160,N_81,N_652);
nor U1161 (N_1161,N_446,N_366);
and U1162 (N_1162,N_661,N_479);
nand U1163 (N_1163,N_155,N_180);
or U1164 (N_1164,N_606,N_55);
or U1165 (N_1165,N_560,N_439);
or U1166 (N_1166,N_628,N_748);
nand U1167 (N_1167,N_66,N_267);
nand U1168 (N_1168,N_180,N_578);
and U1169 (N_1169,N_725,N_650);
or U1170 (N_1170,N_425,N_396);
xnor U1171 (N_1171,N_42,N_424);
and U1172 (N_1172,N_39,N_37);
nand U1173 (N_1173,N_338,N_564);
or U1174 (N_1174,N_710,N_131);
and U1175 (N_1175,N_153,N_126);
and U1176 (N_1176,N_552,N_299);
xnor U1177 (N_1177,N_506,N_690);
or U1178 (N_1178,N_140,N_214);
and U1179 (N_1179,N_748,N_348);
nor U1180 (N_1180,N_307,N_637);
and U1181 (N_1181,N_705,N_184);
xor U1182 (N_1182,N_564,N_667);
and U1183 (N_1183,N_502,N_519);
or U1184 (N_1184,N_661,N_318);
nand U1185 (N_1185,N_359,N_360);
nor U1186 (N_1186,N_419,N_59);
nand U1187 (N_1187,N_307,N_240);
nand U1188 (N_1188,N_467,N_690);
and U1189 (N_1189,N_361,N_230);
nor U1190 (N_1190,N_403,N_0);
and U1191 (N_1191,N_109,N_619);
nand U1192 (N_1192,N_162,N_315);
nor U1193 (N_1193,N_722,N_158);
nand U1194 (N_1194,N_381,N_436);
nand U1195 (N_1195,N_447,N_339);
nor U1196 (N_1196,N_711,N_689);
and U1197 (N_1197,N_237,N_161);
xor U1198 (N_1198,N_551,N_108);
or U1199 (N_1199,N_584,N_528);
nand U1200 (N_1200,N_387,N_618);
nand U1201 (N_1201,N_481,N_98);
nor U1202 (N_1202,N_26,N_212);
or U1203 (N_1203,N_26,N_492);
and U1204 (N_1204,N_320,N_440);
nor U1205 (N_1205,N_702,N_474);
and U1206 (N_1206,N_532,N_386);
or U1207 (N_1207,N_376,N_319);
and U1208 (N_1208,N_373,N_589);
nor U1209 (N_1209,N_636,N_313);
or U1210 (N_1210,N_349,N_690);
or U1211 (N_1211,N_432,N_54);
and U1212 (N_1212,N_254,N_522);
or U1213 (N_1213,N_448,N_259);
nand U1214 (N_1214,N_248,N_282);
nor U1215 (N_1215,N_11,N_673);
nor U1216 (N_1216,N_81,N_722);
or U1217 (N_1217,N_100,N_285);
and U1218 (N_1218,N_209,N_377);
nor U1219 (N_1219,N_59,N_738);
xor U1220 (N_1220,N_206,N_554);
and U1221 (N_1221,N_226,N_348);
nand U1222 (N_1222,N_711,N_695);
xnor U1223 (N_1223,N_649,N_687);
xor U1224 (N_1224,N_286,N_248);
nor U1225 (N_1225,N_99,N_27);
xor U1226 (N_1226,N_445,N_380);
nor U1227 (N_1227,N_547,N_664);
xnor U1228 (N_1228,N_138,N_214);
nor U1229 (N_1229,N_619,N_282);
nand U1230 (N_1230,N_245,N_382);
and U1231 (N_1231,N_680,N_626);
nor U1232 (N_1232,N_583,N_547);
nand U1233 (N_1233,N_242,N_724);
nor U1234 (N_1234,N_358,N_146);
xor U1235 (N_1235,N_501,N_499);
and U1236 (N_1236,N_274,N_355);
or U1237 (N_1237,N_0,N_92);
and U1238 (N_1238,N_303,N_154);
nand U1239 (N_1239,N_493,N_445);
nor U1240 (N_1240,N_711,N_155);
nand U1241 (N_1241,N_455,N_747);
nor U1242 (N_1242,N_86,N_197);
nor U1243 (N_1243,N_13,N_638);
xor U1244 (N_1244,N_517,N_28);
xnor U1245 (N_1245,N_56,N_155);
or U1246 (N_1246,N_662,N_28);
nor U1247 (N_1247,N_674,N_72);
or U1248 (N_1248,N_439,N_237);
xnor U1249 (N_1249,N_210,N_543);
and U1250 (N_1250,N_141,N_551);
nand U1251 (N_1251,N_710,N_577);
and U1252 (N_1252,N_221,N_21);
or U1253 (N_1253,N_287,N_492);
nor U1254 (N_1254,N_598,N_461);
nand U1255 (N_1255,N_586,N_594);
nand U1256 (N_1256,N_445,N_451);
nor U1257 (N_1257,N_46,N_257);
or U1258 (N_1258,N_344,N_337);
or U1259 (N_1259,N_686,N_690);
nor U1260 (N_1260,N_334,N_454);
or U1261 (N_1261,N_118,N_141);
or U1262 (N_1262,N_297,N_197);
and U1263 (N_1263,N_569,N_5);
and U1264 (N_1264,N_148,N_677);
xor U1265 (N_1265,N_390,N_356);
or U1266 (N_1266,N_58,N_376);
nand U1267 (N_1267,N_180,N_716);
and U1268 (N_1268,N_380,N_21);
or U1269 (N_1269,N_486,N_552);
and U1270 (N_1270,N_512,N_384);
xor U1271 (N_1271,N_553,N_706);
nand U1272 (N_1272,N_703,N_14);
nand U1273 (N_1273,N_330,N_638);
and U1274 (N_1274,N_744,N_359);
nand U1275 (N_1275,N_57,N_16);
nand U1276 (N_1276,N_264,N_17);
or U1277 (N_1277,N_469,N_126);
nand U1278 (N_1278,N_400,N_61);
nor U1279 (N_1279,N_631,N_692);
nand U1280 (N_1280,N_701,N_733);
or U1281 (N_1281,N_1,N_613);
nand U1282 (N_1282,N_173,N_273);
and U1283 (N_1283,N_257,N_693);
nor U1284 (N_1284,N_331,N_268);
nand U1285 (N_1285,N_81,N_417);
or U1286 (N_1286,N_120,N_282);
nor U1287 (N_1287,N_77,N_64);
or U1288 (N_1288,N_15,N_706);
nor U1289 (N_1289,N_414,N_464);
or U1290 (N_1290,N_617,N_339);
nor U1291 (N_1291,N_71,N_525);
or U1292 (N_1292,N_481,N_261);
or U1293 (N_1293,N_623,N_17);
xor U1294 (N_1294,N_266,N_157);
or U1295 (N_1295,N_531,N_713);
nand U1296 (N_1296,N_282,N_374);
or U1297 (N_1297,N_146,N_443);
nor U1298 (N_1298,N_90,N_685);
and U1299 (N_1299,N_29,N_411);
or U1300 (N_1300,N_189,N_630);
or U1301 (N_1301,N_318,N_389);
nand U1302 (N_1302,N_238,N_680);
nand U1303 (N_1303,N_344,N_350);
nor U1304 (N_1304,N_533,N_667);
nand U1305 (N_1305,N_107,N_455);
nand U1306 (N_1306,N_418,N_269);
nand U1307 (N_1307,N_363,N_208);
and U1308 (N_1308,N_597,N_550);
and U1309 (N_1309,N_94,N_607);
or U1310 (N_1310,N_185,N_411);
nand U1311 (N_1311,N_717,N_151);
xor U1312 (N_1312,N_282,N_155);
nor U1313 (N_1313,N_622,N_744);
and U1314 (N_1314,N_41,N_635);
xor U1315 (N_1315,N_126,N_5);
xnor U1316 (N_1316,N_86,N_438);
and U1317 (N_1317,N_681,N_356);
or U1318 (N_1318,N_34,N_532);
and U1319 (N_1319,N_170,N_440);
and U1320 (N_1320,N_232,N_417);
or U1321 (N_1321,N_319,N_256);
nor U1322 (N_1322,N_86,N_623);
nand U1323 (N_1323,N_275,N_141);
nand U1324 (N_1324,N_189,N_423);
nor U1325 (N_1325,N_727,N_717);
xor U1326 (N_1326,N_422,N_653);
nand U1327 (N_1327,N_466,N_676);
or U1328 (N_1328,N_261,N_449);
and U1329 (N_1329,N_746,N_193);
and U1330 (N_1330,N_283,N_30);
nor U1331 (N_1331,N_725,N_122);
and U1332 (N_1332,N_671,N_632);
and U1333 (N_1333,N_132,N_146);
and U1334 (N_1334,N_134,N_346);
or U1335 (N_1335,N_42,N_146);
nor U1336 (N_1336,N_122,N_314);
nor U1337 (N_1337,N_549,N_579);
or U1338 (N_1338,N_298,N_478);
or U1339 (N_1339,N_663,N_165);
or U1340 (N_1340,N_695,N_11);
nor U1341 (N_1341,N_305,N_28);
nor U1342 (N_1342,N_494,N_593);
or U1343 (N_1343,N_530,N_363);
nor U1344 (N_1344,N_456,N_149);
nand U1345 (N_1345,N_184,N_241);
nor U1346 (N_1346,N_468,N_150);
or U1347 (N_1347,N_663,N_259);
xnor U1348 (N_1348,N_745,N_596);
or U1349 (N_1349,N_746,N_679);
nand U1350 (N_1350,N_659,N_247);
nor U1351 (N_1351,N_77,N_190);
nor U1352 (N_1352,N_66,N_696);
or U1353 (N_1353,N_5,N_288);
nand U1354 (N_1354,N_497,N_135);
and U1355 (N_1355,N_380,N_275);
or U1356 (N_1356,N_256,N_360);
nand U1357 (N_1357,N_284,N_344);
or U1358 (N_1358,N_748,N_653);
or U1359 (N_1359,N_148,N_8);
nand U1360 (N_1360,N_431,N_518);
or U1361 (N_1361,N_108,N_238);
and U1362 (N_1362,N_23,N_632);
and U1363 (N_1363,N_646,N_297);
xnor U1364 (N_1364,N_498,N_620);
nor U1365 (N_1365,N_489,N_608);
nand U1366 (N_1366,N_480,N_606);
and U1367 (N_1367,N_525,N_160);
nand U1368 (N_1368,N_707,N_682);
and U1369 (N_1369,N_368,N_395);
and U1370 (N_1370,N_447,N_434);
xor U1371 (N_1371,N_130,N_9);
nand U1372 (N_1372,N_509,N_707);
nand U1373 (N_1373,N_249,N_69);
and U1374 (N_1374,N_425,N_187);
and U1375 (N_1375,N_316,N_326);
nand U1376 (N_1376,N_515,N_270);
or U1377 (N_1377,N_638,N_462);
or U1378 (N_1378,N_262,N_640);
nand U1379 (N_1379,N_23,N_299);
xor U1380 (N_1380,N_749,N_338);
nand U1381 (N_1381,N_396,N_229);
nand U1382 (N_1382,N_418,N_21);
nand U1383 (N_1383,N_181,N_285);
and U1384 (N_1384,N_417,N_716);
or U1385 (N_1385,N_197,N_132);
nand U1386 (N_1386,N_211,N_265);
xnor U1387 (N_1387,N_202,N_341);
and U1388 (N_1388,N_471,N_273);
and U1389 (N_1389,N_121,N_445);
nand U1390 (N_1390,N_530,N_229);
nor U1391 (N_1391,N_58,N_658);
nand U1392 (N_1392,N_31,N_625);
and U1393 (N_1393,N_346,N_383);
nor U1394 (N_1394,N_310,N_615);
and U1395 (N_1395,N_399,N_9);
xnor U1396 (N_1396,N_36,N_313);
nand U1397 (N_1397,N_486,N_305);
and U1398 (N_1398,N_681,N_611);
nand U1399 (N_1399,N_539,N_650);
xor U1400 (N_1400,N_562,N_24);
nor U1401 (N_1401,N_613,N_587);
nor U1402 (N_1402,N_603,N_529);
nand U1403 (N_1403,N_580,N_550);
and U1404 (N_1404,N_102,N_121);
or U1405 (N_1405,N_36,N_295);
nand U1406 (N_1406,N_740,N_159);
nand U1407 (N_1407,N_497,N_403);
nand U1408 (N_1408,N_252,N_729);
nor U1409 (N_1409,N_114,N_196);
xor U1410 (N_1410,N_550,N_326);
nor U1411 (N_1411,N_171,N_44);
or U1412 (N_1412,N_69,N_576);
nor U1413 (N_1413,N_734,N_302);
and U1414 (N_1414,N_344,N_482);
or U1415 (N_1415,N_415,N_296);
or U1416 (N_1416,N_628,N_636);
nand U1417 (N_1417,N_365,N_716);
or U1418 (N_1418,N_119,N_419);
nand U1419 (N_1419,N_327,N_364);
or U1420 (N_1420,N_54,N_245);
and U1421 (N_1421,N_252,N_236);
nand U1422 (N_1422,N_179,N_224);
or U1423 (N_1423,N_302,N_270);
nor U1424 (N_1424,N_435,N_368);
and U1425 (N_1425,N_396,N_0);
xnor U1426 (N_1426,N_738,N_217);
xor U1427 (N_1427,N_586,N_564);
or U1428 (N_1428,N_712,N_688);
xnor U1429 (N_1429,N_259,N_186);
xor U1430 (N_1430,N_417,N_225);
nor U1431 (N_1431,N_336,N_115);
and U1432 (N_1432,N_249,N_160);
or U1433 (N_1433,N_299,N_682);
xor U1434 (N_1434,N_123,N_175);
or U1435 (N_1435,N_700,N_480);
xor U1436 (N_1436,N_178,N_165);
nand U1437 (N_1437,N_60,N_656);
or U1438 (N_1438,N_46,N_16);
xor U1439 (N_1439,N_436,N_97);
or U1440 (N_1440,N_214,N_747);
and U1441 (N_1441,N_107,N_688);
xor U1442 (N_1442,N_110,N_730);
nand U1443 (N_1443,N_144,N_617);
nand U1444 (N_1444,N_203,N_138);
nor U1445 (N_1445,N_557,N_14);
nor U1446 (N_1446,N_111,N_668);
nand U1447 (N_1447,N_669,N_464);
and U1448 (N_1448,N_271,N_259);
and U1449 (N_1449,N_624,N_639);
nand U1450 (N_1450,N_676,N_558);
or U1451 (N_1451,N_304,N_339);
and U1452 (N_1452,N_460,N_78);
and U1453 (N_1453,N_241,N_630);
nor U1454 (N_1454,N_685,N_574);
nand U1455 (N_1455,N_129,N_182);
nand U1456 (N_1456,N_119,N_695);
nand U1457 (N_1457,N_711,N_167);
and U1458 (N_1458,N_692,N_439);
and U1459 (N_1459,N_208,N_35);
nor U1460 (N_1460,N_542,N_30);
nor U1461 (N_1461,N_168,N_637);
and U1462 (N_1462,N_209,N_734);
nor U1463 (N_1463,N_663,N_267);
and U1464 (N_1464,N_568,N_72);
nor U1465 (N_1465,N_703,N_47);
nor U1466 (N_1466,N_252,N_387);
or U1467 (N_1467,N_25,N_102);
and U1468 (N_1468,N_729,N_659);
or U1469 (N_1469,N_10,N_274);
xor U1470 (N_1470,N_466,N_430);
nor U1471 (N_1471,N_120,N_630);
nor U1472 (N_1472,N_259,N_442);
or U1473 (N_1473,N_39,N_396);
or U1474 (N_1474,N_489,N_194);
or U1475 (N_1475,N_727,N_441);
xor U1476 (N_1476,N_603,N_68);
nand U1477 (N_1477,N_589,N_397);
xor U1478 (N_1478,N_34,N_605);
nand U1479 (N_1479,N_128,N_559);
or U1480 (N_1480,N_425,N_374);
nand U1481 (N_1481,N_237,N_542);
nor U1482 (N_1482,N_366,N_113);
nor U1483 (N_1483,N_603,N_677);
and U1484 (N_1484,N_639,N_244);
nand U1485 (N_1485,N_1,N_54);
or U1486 (N_1486,N_68,N_219);
or U1487 (N_1487,N_384,N_327);
nand U1488 (N_1488,N_459,N_435);
nor U1489 (N_1489,N_704,N_57);
nor U1490 (N_1490,N_384,N_689);
xnor U1491 (N_1491,N_503,N_398);
nor U1492 (N_1492,N_236,N_110);
or U1493 (N_1493,N_399,N_577);
or U1494 (N_1494,N_146,N_212);
nor U1495 (N_1495,N_143,N_199);
xnor U1496 (N_1496,N_70,N_737);
nor U1497 (N_1497,N_244,N_728);
nand U1498 (N_1498,N_313,N_409);
nor U1499 (N_1499,N_353,N_497);
or U1500 (N_1500,N_1108,N_1376);
nand U1501 (N_1501,N_1161,N_1462);
nor U1502 (N_1502,N_1229,N_1134);
nand U1503 (N_1503,N_816,N_1252);
nor U1504 (N_1504,N_1042,N_1228);
nor U1505 (N_1505,N_974,N_1341);
nor U1506 (N_1506,N_951,N_903);
nand U1507 (N_1507,N_995,N_1198);
or U1508 (N_1508,N_1118,N_1374);
and U1509 (N_1509,N_1052,N_895);
and U1510 (N_1510,N_1081,N_893);
or U1511 (N_1511,N_1095,N_1420);
and U1512 (N_1512,N_971,N_1343);
nand U1513 (N_1513,N_1226,N_1127);
nor U1514 (N_1514,N_1295,N_1002);
or U1515 (N_1515,N_1274,N_976);
nand U1516 (N_1516,N_1003,N_1211);
nand U1517 (N_1517,N_1050,N_1218);
or U1518 (N_1518,N_763,N_1415);
nor U1519 (N_1519,N_755,N_1357);
nor U1520 (N_1520,N_937,N_868);
or U1521 (N_1521,N_1079,N_1253);
nand U1522 (N_1522,N_1383,N_1309);
nand U1523 (N_1523,N_1496,N_1280);
nand U1524 (N_1524,N_1275,N_1167);
nor U1525 (N_1525,N_1290,N_1470);
nor U1526 (N_1526,N_784,N_943);
nor U1527 (N_1527,N_1099,N_1163);
and U1528 (N_1528,N_1306,N_1122);
and U1529 (N_1529,N_1273,N_878);
nand U1530 (N_1530,N_1331,N_1460);
xor U1531 (N_1531,N_914,N_1175);
or U1532 (N_1532,N_1251,N_1245);
nor U1533 (N_1533,N_1027,N_1112);
nor U1534 (N_1534,N_1440,N_970);
nand U1535 (N_1535,N_1354,N_945);
nand U1536 (N_1536,N_1443,N_1316);
nand U1537 (N_1537,N_1086,N_942);
nand U1538 (N_1538,N_1008,N_894);
nand U1539 (N_1539,N_1171,N_876);
or U1540 (N_1540,N_1344,N_1259);
or U1541 (N_1541,N_1399,N_1381);
nand U1542 (N_1542,N_1054,N_1428);
xor U1543 (N_1543,N_1311,N_1370);
or U1544 (N_1544,N_1166,N_1117);
or U1545 (N_1545,N_778,N_800);
nor U1546 (N_1546,N_1413,N_1024);
or U1547 (N_1547,N_1059,N_925);
nor U1548 (N_1548,N_1410,N_799);
nor U1549 (N_1549,N_991,N_968);
xor U1550 (N_1550,N_766,N_1098);
and U1551 (N_1551,N_1206,N_1084);
or U1552 (N_1552,N_1037,N_1405);
nand U1553 (N_1553,N_1009,N_883);
or U1554 (N_1554,N_1264,N_963);
or U1555 (N_1555,N_1493,N_1185);
nor U1556 (N_1556,N_844,N_1326);
and U1557 (N_1557,N_1312,N_1479);
or U1558 (N_1558,N_757,N_1269);
nand U1559 (N_1559,N_777,N_1395);
xnor U1560 (N_1560,N_1313,N_1058);
and U1561 (N_1561,N_1102,N_1246);
nand U1562 (N_1562,N_1499,N_1115);
nand U1563 (N_1563,N_980,N_1157);
nor U1564 (N_1564,N_1183,N_865);
nor U1565 (N_1565,N_1406,N_1408);
or U1566 (N_1566,N_1116,N_789);
and U1567 (N_1567,N_1466,N_1071);
nand U1568 (N_1568,N_1421,N_1109);
nor U1569 (N_1569,N_803,N_1392);
nand U1570 (N_1570,N_1317,N_1184);
nand U1571 (N_1571,N_910,N_1203);
nand U1572 (N_1572,N_785,N_1485);
or U1573 (N_1573,N_1459,N_1138);
and U1574 (N_1574,N_847,N_1400);
or U1575 (N_1575,N_798,N_1451);
and U1576 (N_1576,N_1414,N_1104);
nand U1577 (N_1577,N_1186,N_1474);
nand U1578 (N_1578,N_1256,N_939);
or U1579 (N_1579,N_1366,N_1445);
xor U1580 (N_1580,N_1461,N_1358);
nand U1581 (N_1581,N_1178,N_790);
or U1582 (N_1582,N_905,N_1193);
nand U1583 (N_1583,N_1465,N_1267);
or U1584 (N_1584,N_1236,N_959);
nand U1585 (N_1585,N_1080,N_1154);
nand U1586 (N_1586,N_975,N_1205);
and U1587 (N_1587,N_912,N_1452);
nor U1588 (N_1588,N_954,N_1135);
and U1589 (N_1589,N_1006,N_852);
or U1590 (N_1590,N_873,N_1097);
nor U1591 (N_1591,N_885,N_1279);
nand U1592 (N_1592,N_882,N_1302);
nand U1593 (N_1593,N_787,N_794);
or U1594 (N_1594,N_1417,N_1332);
or U1595 (N_1595,N_916,N_753);
nor U1596 (N_1596,N_1215,N_855);
nor U1597 (N_1597,N_819,N_1057);
or U1598 (N_1598,N_839,N_1026);
nand U1599 (N_1599,N_1077,N_1022);
or U1600 (N_1600,N_1068,N_1450);
nor U1601 (N_1601,N_933,N_960);
and U1602 (N_1602,N_1333,N_831);
nor U1603 (N_1603,N_890,N_775);
nand U1604 (N_1604,N_1238,N_1260);
nand U1605 (N_1605,N_1004,N_926);
and U1606 (N_1606,N_824,N_1321);
nand U1607 (N_1607,N_817,N_1268);
nor U1608 (N_1608,N_1085,N_1149);
nor U1609 (N_1609,N_1000,N_1001);
nor U1610 (N_1610,N_961,N_1403);
or U1611 (N_1611,N_825,N_857);
xor U1612 (N_1612,N_1363,N_1033);
and U1613 (N_1613,N_1012,N_1423);
and U1614 (N_1614,N_1367,N_1432);
nor U1615 (N_1615,N_1481,N_1338);
or U1616 (N_1616,N_1488,N_1457);
xor U1617 (N_1617,N_812,N_1244);
nor U1618 (N_1618,N_1285,N_1032);
and U1619 (N_1619,N_1204,N_1362);
nand U1620 (N_1620,N_1239,N_1340);
or U1621 (N_1621,N_1296,N_1231);
nor U1622 (N_1622,N_1299,N_1463);
nand U1623 (N_1623,N_1441,N_1349);
and U1624 (N_1624,N_1491,N_1062);
nor U1625 (N_1625,N_1293,N_966);
nand U1626 (N_1626,N_849,N_1212);
nand U1627 (N_1627,N_801,N_1105);
and U1628 (N_1628,N_1276,N_1156);
nor U1629 (N_1629,N_987,N_1137);
nor U1630 (N_1630,N_1436,N_1458);
nand U1631 (N_1631,N_913,N_1390);
and U1632 (N_1632,N_1036,N_1411);
nor U1633 (N_1633,N_811,N_1132);
and U1634 (N_1634,N_908,N_906);
or U1635 (N_1635,N_899,N_887);
or U1636 (N_1636,N_822,N_1017);
nor U1637 (N_1637,N_1224,N_953);
nand U1638 (N_1638,N_1483,N_1325);
nor U1639 (N_1639,N_802,N_1110);
nor U1640 (N_1640,N_1075,N_917);
nor U1641 (N_1641,N_1195,N_769);
or U1642 (N_1642,N_1010,N_1375);
or U1643 (N_1643,N_1409,N_752);
or U1644 (N_1644,N_1160,N_1039);
nor U1645 (N_1645,N_998,N_901);
nor U1646 (N_1646,N_1048,N_1418);
nor U1647 (N_1647,N_754,N_1490);
and U1648 (N_1648,N_1216,N_1043);
nand U1649 (N_1649,N_1119,N_1208);
and U1650 (N_1650,N_1250,N_1072);
and U1651 (N_1651,N_1223,N_1412);
and U1652 (N_1652,N_1194,N_973);
or U1653 (N_1653,N_772,N_1155);
and U1654 (N_1654,N_1067,N_1255);
or U1655 (N_1655,N_904,N_1243);
nand U1656 (N_1656,N_947,N_1439);
and U1657 (N_1657,N_1069,N_1126);
or U1658 (N_1658,N_877,N_1368);
nor U1659 (N_1659,N_773,N_1284);
nand U1660 (N_1660,N_919,N_1046);
and U1661 (N_1661,N_923,N_1301);
xor U1662 (N_1662,N_1448,N_1217);
nand U1663 (N_1663,N_1304,N_1329);
nor U1664 (N_1664,N_1242,N_1143);
nor U1665 (N_1665,N_964,N_1360);
nand U1666 (N_1666,N_1416,N_1453);
or U1667 (N_1667,N_1222,N_1371);
nand U1668 (N_1668,N_1484,N_1425);
nor U1669 (N_1669,N_1107,N_922);
and U1670 (N_1670,N_1189,N_1020);
or U1671 (N_1671,N_1289,N_1153);
nand U1672 (N_1672,N_1078,N_997);
and U1673 (N_1673,N_1021,N_863);
or U1674 (N_1674,N_1292,N_1121);
or U1675 (N_1675,N_815,N_1031);
and U1676 (N_1676,N_1064,N_999);
or U1677 (N_1677,N_1364,N_1431);
nand U1678 (N_1678,N_793,N_1356);
and U1679 (N_1679,N_1232,N_765);
nand U1680 (N_1680,N_1045,N_946);
nor U1681 (N_1681,N_1380,N_1144);
nor U1682 (N_1682,N_1388,N_1477);
or U1683 (N_1683,N_1398,N_1319);
xnor U1684 (N_1684,N_1318,N_761);
or U1685 (N_1685,N_1190,N_940);
nor U1686 (N_1686,N_762,N_1047);
and U1687 (N_1687,N_1365,N_1327);
nand U1688 (N_1688,N_1261,N_1014);
or U1689 (N_1689,N_1051,N_1262);
nor U1690 (N_1690,N_860,N_1391);
nand U1691 (N_1691,N_1307,N_1019);
nor U1692 (N_1692,N_1191,N_1225);
nor U1693 (N_1693,N_1049,N_1114);
or U1694 (N_1694,N_788,N_1288);
nor U1695 (N_1695,N_935,N_758);
nand U1696 (N_1696,N_1435,N_770);
or U1697 (N_1697,N_1430,N_1145);
or U1698 (N_1698,N_934,N_1029);
xor U1699 (N_1699,N_921,N_1422);
xnor U1700 (N_1700,N_1053,N_1397);
and U1701 (N_1701,N_1424,N_1091);
nor U1702 (N_1702,N_928,N_1182);
nand U1703 (N_1703,N_1188,N_1350);
and U1704 (N_1704,N_909,N_1221);
or U1705 (N_1705,N_1489,N_1196);
and U1706 (N_1706,N_833,N_1162);
or U1707 (N_1707,N_1164,N_1283);
or U1708 (N_1708,N_892,N_814);
or U1709 (N_1709,N_1214,N_1455);
nand U1710 (N_1710,N_1468,N_1101);
nand U1711 (N_1711,N_1096,N_861);
nand U1712 (N_1712,N_1007,N_977);
nand U1713 (N_1713,N_1035,N_1240);
nand U1714 (N_1714,N_897,N_872);
and U1715 (N_1715,N_1330,N_1070);
or U1716 (N_1716,N_1347,N_911);
and U1717 (N_1717,N_1192,N_1136);
or U1718 (N_1718,N_1265,N_829);
or U1719 (N_1719,N_1278,N_841);
nand U1720 (N_1720,N_1492,N_1005);
nand U1721 (N_1721,N_1056,N_1148);
nand U1722 (N_1722,N_992,N_1300);
nor U1723 (N_1723,N_949,N_1237);
nand U1724 (N_1724,N_907,N_988);
nand U1725 (N_1725,N_871,N_936);
xnor U1726 (N_1726,N_1170,N_948);
xnor U1727 (N_1727,N_938,N_950);
nand U1728 (N_1728,N_821,N_981);
nand U1729 (N_1729,N_1444,N_955);
nand U1730 (N_1730,N_1201,N_1103);
and U1731 (N_1731,N_1241,N_1387);
and U1732 (N_1732,N_902,N_978);
nor U1733 (N_1733,N_1011,N_1210);
and U1734 (N_1734,N_1315,N_989);
and U1735 (N_1735,N_780,N_809);
xnor U1736 (N_1736,N_1066,N_1179);
and U1737 (N_1737,N_856,N_1257);
nand U1738 (N_1738,N_1025,N_1339);
nor U1739 (N_1739,N_1176,N_1073);
xnor U1740 (N_1740,N_826,N_783);
nand U1741 (N_1741,N_1482,N_1016);
and U1742 (N_1742,N_804,N_1034);
or U1743 (N_1743,N_1040,N_1041);
nand U1744 (N_1744,N_1291,N_867);
nor U1745 (N_1745,N_1270,N_786);
nor U1746 (N_1746,N_1351,N_1158);
nand U1747 (N_1747,N_1092,N_1335);
and U1748 (N_1748,N_1233,N_781);
nand U1749 (N_1749,N_862,N_1087);
or U1750 (N_1750,N_927,N_898);
or U1751 (N_1751,N_1133,N_1038);
nor U1752 (N_1752,N_779,N_1235);
nor U1753 (N_1753,N_854,N_1028);
xor U1754 (N_1754,N_1456,N_1227);
nand U1755 (N_1755,N_1230,N_836);
nor U1756 (N_1756,N_797,N_1180);
xnor U1757 (N_1757,N_1013,N_792);
or U1758 (N_1758,N_1181,N_1476);
or U1759 (N_1759,N_1100,N_1248);
nor U1760 (N_1760,N_1487,N_1345);
nor U1761 (N_1761,N_1386,N_1464);
or U1762 (N_1762,N_929,N_1055);
nor U1763 (N_1763,N_1174,N_918);
or U1764 (N_1764,N_1199,N_1384);
and U1765 (N_1765,N_1207,N_1377);
nor U1766 (N_1766,N_1478,N_986);
nor U1767 (N_1767,N_1297,N_984);
nor U1768 (N_1768,N_771,N_866);
and U1769 (N_1769,N_838,N_1131);
nand U1770 (N_1770,N_967,N_807);
xnor U1771 (N_1771,N_834,N_1219);
xnor U1772 (N_1772,N_979,N_1310);
nand U1773 (N_1773,N_759,N_810);
and U1774 (N_1774,N_805,N_1385);
and U1775 (N_1775,N_1060,N_1082);
or U1776 (N_1776,N_1369,N_827);
nor U1777 (N_1777,N_1177,N_782);
and U1778 (N_1778,N_931,N_1447);
nand U1779 (N_1779,N_851,N_1169);
nor U1780 (N_1780,N_982,N_1434);
or U1781 (N_1781,N_1497,N_1352);
nand U1782 (N_1782,N_1187,N_972);
nand U1783 (N_1783,N_858,N_1437);
or U1784 (N_1784,N_1378,N_845);
or U1785 (N_1785,N_1475,N_1328);
nor U1786 (N_1786,N_1258,N_1234);
or U1787 (N_1787,N_1030,N_1125);
and U1788 (N_1788,N_1427,N_1090);
or U1789 (N_1789,N_796,N_1438);
nor U1790 (N_1790,N_843,N_1140);
nor U1791 (N_1791,N_1308,N_1172);
and U1792 (N_1792,N_932,N_1382);
and U1793 (N_1793,N_1372,N_944);
and U1794 (N_1794,N_837,N_806);
nand U1795 (N_1795,N_888,N_830);
nand U1796 (N_1796,N_1220,N_1141);
nor U1797 (N_1797,N_985,N_1094);
nand U1798 (N_1798,N_1498,N_1023);
nor U1799 (N_1799,N_1173,N_768);
or U1800 (N_1800,N_1305,N_1197);
nand U1801 (N_1801,N_1467,N_1083);
and U1802 (N_1802,N_1247,N_1353);
nand U1803 (N_1803,N_1433,N_1480);
nand U1804 (N_1804,N_1159,N_869);
xnor U1805 (N_1805,N_983,N_1394);
nand U1806 (N_1806,N_1142,N_1129);
nand U1807 (N_1807,N_1359,N_1337);
xor U1808 (N_1808,N_1200,N_1287);
or U1809 (N_1809,N_930,N_832);
nor U1810 (N_1810,N_828,N_884);
and U1811 (N_1811,N_1015,N_1389);
nand U1812 (N_1812,N_840,N_850);
or U1813 (N_1813,N_750,N_859);
nor U1814 (N_1814,N_1471,N_924);
nand U1815 (N_1815,N_958,N_1130);
and U1816 (N_1816,N_1379,N_1202);
nor U1817 (N_1817,N_1303,N_891);
or U1818 (N_1818,N_1076,N_760);
nand U1819 (N_1819,N_823,N_874);
or U1820 (N_1820,N_1402,N_915);
nand U1821 (N_1821,N_756,N_1147);
or U1822 (N_1822,N_1113,N_957);
and U1823 (N_1823,N_1286,N_751);
xor U1824 (N_1824,N_1263,N_791);
nor U1825 (N_1825,N_1088,N_1213);
or U1826 (N_1826,N_864,N_1150);
nand U1827 (N_1827,N_1146,N_875);
or U1828 (N_1828,N_1419,N_962);
xnor U1829 (N_1829,N_1209,N_1314);
or U1830 (N_1830,N_941,N_969);
or U1831 (N_1831,N_1320,N_1089);
and U1832 (N_1832,N_965,N_886);
or U1833 (N_1833,N_1271,N_1336);
xor U1834 (N_1834,N_1124,N_764);
xnor U1835 (N_1835,N_1323,N_1429);
and U1836 (N_1836,N_1106,N_774);
xnor U1837 (N_1837,N_1044,N_1342);
or U1838 (N_1838,N_993,N_1074);
nor U1839 (N_1839,N_1401,N_1281);
or U1840 (N_1840,N_1346,N_808);
nor U1841 (N_1841,N_1249,N_1018);
or U1842 (N_1842,N_1348,N_1324);
xor U1843 (N_1843,N_870,N_881);
nand U1844 (N_1844,N_1373,N_842);
xnor U1845 (N_1845,N_900,N_1266);
and U1846 (N_1846,N_1355,N_1128);
or U1847 (N_1847,N_1152,N_920);
nand U1848 (N_1848,N_1426,N_1151);
nand U1849 (N_1849,N_1407,N_853);
nor U1850 (N_1850,N_1282,N_1472);
or U1851 (N_1851,N_1065,N_1093);
nor U1852 (N_1852,N_956,N_1396);
nor U1853 (N_1853,N_1111,N_896);
nor U1854 (N_1854,N_820,N_1165);
nor U1855 (N_1855,N_990,N_994);
or U1856 (N_1856,N_1322,N_846);
nor U1857 (N_1857,N_1449,N_776);
and U1858 (N_1858,N_1123,N_1277);
or U1859 (N_1859,N_1294,N_1494);
or U1860 (N_1860,N_1061,N_1404);
nor U1861 (N_1861,N_1063,N_1254);
nand U1862 (N_1862,N_1495,N_1469);
or U1863 (N_1863,N_1454,N_889);
nand U1864 (N_1864,N_835,N_1168);
or U1865 (N_1865,N_1486,N_1446);
xnor U1866 (N_1866,N_818,N_848);
or U1867 (N_1867,N_880,N_1272);
nand U1868 (N_1868,N_1442,N_1361);
xnor U1869 (N_1869,N_767,N_1473);
or U1870 (N_1870,N_813,N_795);
or U1871 (N_1871,N_952,N_1393);
or U1872 (N_1872,N_1334,N_1120);
and U1873 (N_1873,N_1298,N_996);
xor U1874 (N_1874,N_1139,N_879);
nor U1875 (N_1875,N_918,N_1039);
nand U1876 (N_1876,N_765,N_1031);
and U1877 (N_1877,N_1093,N_886);
nand U1878 (N_1878,N_1149,N_1310);
nand U1879 (N_1879,N_893,N_1009);
or U1880 (N_1880,N_1216,N_752);
xnor U1881 (N_1881,N_1075,N_1069);
or U1882 (N_1882,N_1079,N_1046);
nand U1883 (N_1883,N_914,N_1168);
nand U1884 (N_1884,N_873,N_901);
and U1885 (N_1885,N_1310,N_1263);
nor U1886 (N_1886,N_1391,N_1234);
nand U1887 (N_1887,N_964,N_949);
and U1888 (N_1888,N_1047,N_1142);
nor U1889 (N_1889,N_1353,N_1328);
and U1890 (N_1890,N_1225,N_826);
or U1891 (N_1891,N_1412,N_984);
nor U1892 (N_1892,N_1275,N_896);
and U1893 (N_1893,N_1453,N_1117);
and U1894 (N_1894,N_808,N_814);
nor U1895 (N_1895,N_885,N_1023);
or U1896 (N_1896,N_1286,N_1042);
nor U1897 (N_1897,N_1227,N_761);
and U1898 (N_1898,N_1018,N_1407);
nand U1899 (N_1899,N_1176,N_1431);
and U1900 (N_1900,N_980,N_1038);
nor U1901 (N_1901,N_1411,N_1197);
and U1902 (N_1902,N_1419,N_946);
nand U1903 (N_1903,N_1163,N_1313);
and U1904 (N_1904,N_1285,N_944);
and U1905 (N_1905,N_1488,N_775);
or U1906 (N_1906,N_1198,N_1002);
nand U1907 (N_1907,N_1129,N_765);
nand U1908 (N_1908,N_1097,N_1278);
and U1909 (N_1909,N_1468,N_772);
nor U1910 (N_1910,N_1064,N_1319);
nand U1911 (N_1911,N_766,N_805);
or U1912 (N_1912,N_859,N_1211);
nand U1913 (N_1913,N_819,N_1063);
and U1914 (N_1914,N_1127,N_1430);
nand U1915 (N_1915,N_862,N_1461);
nand U1916 (N_1916,N_914,N_1357);
nor U1917 (N_1917,N_1026,N_796);
nand U1918 (N_1918,N_1460,N_941);
or U1919 (N_1919,N_960,N_1242);
nand U1920 (N_1920,N_852,N_901);
nand U1921 (N_1921,N_976,N_1194);
and U1922 (N_1922,N_1158,N_1424);
and U1923 (N_1923,N_1361,N_1068);
and U1924 (N_1924,N_963,N_763);
nor U1925 (N_1925,N_943,N_1351);
nand U1926 (N_1926,N_1377,N_1399);
xnor U1927 (N_1927,N_821,N_1036);
xnor U1928 (N_1928,N_770,N_787);
and U1929 (N_1929,N_1422,N_980);
nand U1930 (N_1930,N_1233,N_861);
and U1931 (N_1931,N_1189,N_1062);
nand U1932 (N_1932,N_769,N_1387);
nand U1933 (N_1933,N_1384,N_956);
nor U1934 (N_1934,N_1287,N_1465);
or U1935 (N_1935,N_1244,N_1490);
or U1936 (N_1936,N_1374,N_1249);
or U1937 (N_1937,N_1157,N_1317);
nand U1938 (N_1938,N_1377,N_856);
nor U1939 (N_1939,N_782,N_941);
or U1940 (N_1940,N_1437,N_803);
or U1941 (N_1941,N_1083,N_820);
and U1942 (N_1942,N_1398,N_1330);
and U1943 (N_1943,N_1339,N_1056);
and U1944 (N_1944,N_757,N_1233);
nor U1945 (N_1945,N_757,N_1438);
nor U1946 (N_1946,N_1110,N_1180);
nor U1947 (N_1947,N_895,N_1019);
nand U1948 (N_1948,N_1333,N_1487);
nand U1949 (N_1949,N_789,N_851);
xnor U1950 (N_1950,N_925,N_1201);
and U1951 (N_1951,N_828,N_1469);
and U1952 (N_1952,N_770,N_1007);
or U1953 (N_1953,N_1202,N_1168);
nor U1954 (N_1954,N_875,N_1214);
or U1955 (N_1955,N_963,N_865);
and U1956 (N_1956,N_1267,N_1284);
or U1957 (N_1957,N_1399,N_1076);
nand U1958 (N_1958,N_817,N_1048);
nand U1959 (N_1959,N_1150,N_894);
or U1960 (N_1960,N_1161,N_957);
and U1961 (N_1961,N_1340,N_1168);
nor U1962 (N_1962,N_1352,N_997);
or U1963 (N_1963,N_1306,N_854);
and U1964 (N_1964,N_1204,N_1304);
or U1965 (N_1965,N_969,N_1181);
nand U1966 (N_1966,N_1304,N_1060);
nor U1967 (N_1967,N_1473,N_1043);
or U1968 (N_1968,N_1030,N_983);
xor U1969 (N_1969,N_955,N_1034);
nor U1970 (N_1970,N_840,N_789);
or U1971 (N_1971,N_1207,N_1315);
nand U1972 (N_1972,N_944,N_1392);
nor U1973 (N_1973,N_780,N_1300);
or U1974 (N_1974,N_1031,N_1390);
and U1975 (N_1975,N_1115,N_1070);
and U1976 (N_1976,N_1196,N_1309);
xor U1977 (N_1977,N_1499,N_996);
xor U1978 (N_1978,N_1039,N_1314);
nand U1979 (N_1979,N_1293,N_1394);
nand U1980 (N_1980,N_1338,N_1428);
and U1981 (N_1981,N_1489,N_1076);
xor U1982 (N_1982,N_924,N_1107);
and U1983 (N_1983,N_849,N_1066);
nor U1984 (N_1984,N_1225,N_1248);
nor U1985 (N_1985,N_1104,N_1074);
nor U1986 (N_1986,N_1467,N_949);
and U1987 (N_1987,N_843,N_1438);
or U1988 (N_1988,N_1233,N_810);
and U1989 (N_1989,N_882,N_789);
nor U1990 (N_1990,N_821,N_813);
nor U1991 (N_1991,N_1332,N_1114);
nand U1992 (N_1992,N_1432,N_979);
and U1993 (N_1993,N_1141,N_1058);
nand U1994 (N_1994,N_968,N_855);
nand U1995 (N_1995,N_1453,N_761);
nor U1996 (N_1996,N_1120,N_1155);
or U1997 (N_1997,N_1104,N_1218);
nand U1998 (N_1998,N_1485,N_1426);
nor U1999 (N_1999,N_880,N_871);
xnor U2000 (N_2000,N_1462,N_917);
and U2001 (N_2001,N_996,N_817);
nor U2002 (N_2002,N_904,N_932);
nor U2003 (N_2003,N_1261,N_1086);
nor U2004 (N_2004,N_1043,N_1484);
or U2005 (N_2005,N_845,N_1221);
and U2006 (N_2006,N_1096,N_1384);
nand U2007 (N_2007,N_1045,N_1046);
nor U2008 (N_2008,N_1350,N_1132);
or U2009 (N_2009,N_1222,N_1032);
nor U2010 (N_2010,N_1036,N_823);
xnor U2011 (N_2011,N_998,N_954);
and U2012 (N_2012,N_840,N_1112);
nand U2013 (N_2013,N_1283,N_1093);
nor U2014 (N_2014,N_929,N_852);
xor U2015 (N_2015,N_767,N_751);
or U2016 (N_2016,N_1196,N_1441);
nor U2017 (N_2017,N_811,N_1481);
and U2018 (N_2018,N_1449,N_981);
nor U2019 (N_2019,N_853,N_1319);
and U2020 (N_2020,N_875,N_1143);
and U2021 (N_2021,N_1378,N_790);
and U2022 (N_2022,N_1393,N_1171);
nand U2023 (N_2023,N_883,N_1304);
nor U2024 (N_2024,N_1321,N_1005);
and U2025 (N_2025,N_924,N_1139);
and U2026 (N_2026,N_1250,N_1042);
and U2027 (N_2027,N_1440,N_1259);
or U2028 (N_2028,N_1469,N_1464);
xor U2029 (N_2029,N_1133,N_1132);
nand U2030 (N_2030,N_1084,N_1350);
or U2031 (N_2031,N_959,N_1342);
or U2032 (N_2032,N_1005,N_858);
or U2033 (N_2033,N_1320,N_1134);
or U2034 (N_2034,N_788,N_1146);
nor U2035 (N_2035,N_902,N_880);
nand U2036 (N_2036,N_822,N_1355);
nand U2037 (N_2037,N_1496,N_1055);
nand U2038 (N_2038,N_815,N_1207);
or U2039 (N_2039,N_1317,N_842);
nand U2040 (N_2040,N_932,N_1185);
or U2041 (N_2041,N_819,N_766);
nand U2042 (N_2042,N_981,N_1137);
nor U2043 (N_2043,N_1056,N_1197);
or U2044 (N_2044,N_1264,N_1094);
nand U2045 (N_2045,N_921,N_1177);
nand U2046 (N_2046,N_1007,N_1419);
nand U2047 (N_2047,N_777,N_1055);
nor U2048 (N_2048,N_922,N_1256);
or U2049 (N_2049,N_1071,N_1328);
xor U2050 (N_2050,N_1140,N_1326);
or U2051 (N_2051,N_1231,N_841);
and U2052 (N_2052,N_1158,N_1272);
and U2053 (N_2053,N_1436,N_879);
xnor U2054 (N_2054,N_914,N_937);
or U2055 (N_2055,N_1163,N_1392);
nand U2056 (N_2056,N_992,N_999);
or U2057 (N_2057,N_1252,N_959);
and U2058 (N_2058,N_1020,N_1169);
nor U2059 (N_2059,N_871,N_1294);
nand U2060 (N_2060,N_1210,N_858);
and U2061 (N_2061,N_1405,N_1417);
nand U2062 (N_2062,N_1299,N_1333);
and U2063 (N_2063,N_1301,N_1091);
or U2064 (N_2064,N_1139,N_1408);
nor U2065 (N_2065,N_1383,N_1045);
or U2066 (N_2066,N_869,N_1065);
nand U2067 (N_2067,N_1297,N_1305);
or U2068 (N_2068,N_949,N_943);
nand U2069 (N_2069,N_1050,N_920);
and U2070 (N_2070,N_1132,N_1393);
nor U2071 (N_2071,N_893,N_1128);
nor U2072 (N_2072,N_1108,N_1269);
nor U2073 (N_2073,N_1078,N_774);
nand U2074 (N_2074,N_1246,N_1453);
xor U2075 (N_2075,N_1458,N_944);
or U2076 (N_2076,N_1364,N_791);
nand U2077 (N_2077,N_1028,N_1371);
or U2078 (N_2078,N_1497,N_1275);
xnor U2079 (N_2079,N_963,N_1099);
and U2080 (N_2080,N_1032,N_1001);
xor U2081 (N_2081,N_810,N_931);
or U2082 (N_2082,N_1035,N_1145);
nand U2083 (N_2083,N_897,N_870);
nand U2084 (N_2084,N_1362,N_1000);
xnor U2085 (N_2085,N_1334,N_911);
xnor U2086 (N_2086,N_757,N_1495);
and U2087 (N_2087,N_1052,N_1469);
and U2088 (N_2088,N_789,N_1319);
and U2089 (N_2089,N_1126,N_1016);
nor U2090 (N_2090,N_1100,N_1251);
nor U2091 (N_2091,N_1283,N_1073);
or U2092 (N_2092,N_832,N_1497);
nand U2093 (N_2093,N_751,N_1430);
or U2094 (N_2094,N_973,N_1017);
nor U2095 (N_2095,N_766,N_1389);
nor U2096 (N_2096,N_856,N_1263);
nand U2097 (N_2097,N_1031,N_1266);
nor U2098 (N_2098,N_1232,N_1002);
nand U2099 (N_2099,N_940,N_1273);
and U2100 (N_2100,N_979,N_828);
nand U2101 (N_2101,N_835,N_941);
or U2102 (N_2102,N_800,N_927);
nand U2103 (N_2103,N_805,N_1397);
and U2104 (N_2104,N_884,N_883);
and U2105 (N_2105,N_1025,N_1187);
and U2106 (N_2106,N_921,N_888);
or U2107 (N_2107,N_1035,N_1010);
nor U2108 (N_2108,N_1343,N_1210);
xnor U2109 (N_2109,N_1369,N_1034);
and U2110 (N_2110,N_1275,N_1399);
nand U2111 (N_2111,N_979,N_1115);
and U2112 (N_2112,N_815,N_925);
or U2113 (N_2113,N_1215,N_870);
xor U2114 (N_2114,N_1440,N_916);
nand U2115 (N_2115,N_1431,N_1343);
nor U2116 (N_2116,N_1035,N_1327);
nand U2117 (N_2117,N_756,N_811);
or U2118 (N_2118,N_949,N_1255);
nand U2119 (N_2119,N_1096,N_758);
nand U2120 (N_2120,N_814,N_974);
and U2121 (N_2121,N_996,N_994);
nand U2122 (N_2122,N_960,N_997);
or U2123 (N_2123,N_1323,N_803);
nor U2124 (N_2124,N_1337,N_1421);
and U2125 (N_2125,N_1201,N_908);
nor U2126 (N_2126,N_1247,N_1429);
xnor U2127 (N_2127,N_1030,N_1000);
or U2128 (N_2128,N_1373,N_1299);
nor U2129 (N_2129,N_1202,N_1425);
nand U2130 (N_2130,N_865,N_1056);
xnor U2131 (N_2131,N_1203,N_1007);
or U2132 (N_2132,N_1387,N_1204);
or U2133 (N_2133,N_945,N_1014);
and U2134 (N_2134,N_1327,N_1072);
and U2135 (N_2135,N_931,N_1120);
nor U2136 (N_2136,N_1143,N_1412);
nand U2137 (N_2137,N_1088,N_1205);
and U2138 (N_2138,N_784,N_1034);
nand U2139 (N_2139,N_1428,N_1224);
and U2140 (N_2140,N_1333,N_1356);
nand U2141 (N_2141,N_946,N_1222);
nand U2142 (N_2142,N_1109,N_958);
and U2143 (N_2143,N_959,N_1288);
or U2144 (N_2144,N_1348,N_1107);
nor U2145 (N_2145,N_1448,N_842);
and U2146 (N_2146,N_1309,N_760);
or U2147 (N_2147,N_1164,N_1208);
or U2148 (N_2148,N_1463,N_1228);
xnor U2149 (N_2149,N_1172,N_750);
nor U2150 (N_2150,N_1312,N_888);
and U2151 (N_2151,N_752,N_1381);
xor U2152 (N_2152,N_1486,N_1077);
and U2153 (N_2153,N_1146,N_1456);
and U2154 (N_2154,N_801,N_1075);
xor U2155 (N_2155,N_1276,N_962);
or U2156 (N_2156,N_1244,N_787);
or U2157 (N_2157,N_763,N_1232);
and U2158 (N_2158,N_1289,N_1495);
nand U2159 (N_2159,N_838,N_797);
or U2160 (N_2160,N_794,N_1106);
and U2161 (N_2161,N_762,N_1324);
and U2162 (N_2162,N_811,N_986);
and U2163 (N_2163,N_1116,N_784);
and U2164 (N_2164,N_835,N_940);
or U2165 (N_2165,N_1487,N_1309);
nand U2166 (N_2166,N_819,N_1142);
xnor U2167 (N_2167,N_1121,N_1499);
or U2168 (N_2168,N_938,N_1131);
and U2169 (N_2169,N_1227,N_1463);
or U2170 (N_2170,N_792,N_873);
or U2171 (N_2171,N_1231,N_1155);
xor U2172 (N_2172,N_786,N_1229);
nand U2173 (N_2173,N_967,N_1156);
nor U2174 (N_2174,N_1025,N_1299);
or U2175 (N_2175,N_1488,N_1036);
and U2176 (N_2176,N_854,N_834);
and U2177 (N_2177,N_1147,N_957);
and U2178 (N_2178,N_1146,N_1110);
nand U2179 (N_2179,N_1028,N_828);
and U2180 (N_2180,N_1007,N_1259);
and U2181 (N_2181,N_1447,N_1226);
nand U2182 (N_2182,N_1452,N_1018);
or U2183 (N_2183,N_940,N_990);
and U2184 (N_2184,N_1207,N_830);
or U2185 (N_2185,N_1382,N_1231);
and U2186 (N_2186,N_1247,N_784);
and U2187 (N_2187,N_1334,N_1092);
and U2188 (N_2188,N_771,N_952);
nor U2189 (N_2189,N_1320,N_880);
nor U2190 (N_2190,N_1357,N_1365);
nand U2191 (N_2191,N_1187,N_1195);
or U2192 (N_2192,N_829,N_1122);
nor U2193 (N_2193,N_1255,N_1470);
xnor U2194 (N_2194,N_1034,N_1434);
nand U2195 (N_2195,N_1494,N_786);
xnor U2196 (N_2196,N_758,N_1000);
and U2197 (N_2197,N_1138,N_812);
and U2198 (N_2198,N_1377,N_1091);
or U2199 (N_2199,N_991,N_1468);
or U2200 (N_2200,N_826,N_1485);
xnor U2201 (N_2201,N_971,N_1256);
nor U2202 (N_2202,N_1048,N_775);
nor U2203 (N_2203,N_1340,N_1390);
and U2204 (N_2204,N_1434,N_1011);
or U2205 (N_2205,N_1319,N_1385);
or U2206 (N_2206,N_913,N_1370);
xor U2207 (N_2207,N_1262,N_846);
nor U2208 (N_2208,N_987,N_1074);
nor U2209 (N_2209,N_857,N_1408);
nor U2210 (N_2210,N_1279,N_1375);
nand U2211 (N_2211,N_831,N_1122);
or U2212 (N_2212,N_1465,N_864);
or U2213 (N_2213,N_1197,N_1496);
nor U2214 (N_2214,N_1314,N_924);
nand U2215 (N_2215,N_853,N_1216);
or U2216 (N_2216,N_814,N_1390);
and U2217 (N_2217,N_887,N_1016);
nor U2218 (N_2218,N_1336,N_1101);
or U2219 (N_2219,N_1271,N_954);
xor U2220 (N_2220,N_952,N_1117);
and U2221 (N_2221,N_1356,N_1250);
xor U2222 (N_2222,N_1162,N_800);
or U2223 (N_2223,N_1195,N_750);
or U2224 (N_2224,N_1134,N_1257);
xnor U2225 (N_2225,N_1315,N_1452);
nand U2226 (N_2226,N_1019,N_1140);
nor U2227 (N_2227,N_1058,N_772);
nand U2228 (N_2228,N_950,N_760);
or U2229 (N_2229,N_1245,N_1216);
xor U2230 (N_2230,N_1352,N_1247);
and U2231 (N_2231,N_1448,N_857);
and U2232 (N_2232,N_1073,N_1033);
or U2233 (N_2233,N_1117,N_1263);
or U2234 (N_2234,N_1229,N_864);
and U2235 (N_2235,N_1463,N_1114);
nor U2236 (N_2236,N_1277,N_1399);
nor U2237 (N_2237,N_1363,N_1292);
and U2238 (N_2238,N_778,N_1327);
nor U2239 (N_2239,N_1047,N_895);
or U2240 (N_2240,N_1246,N_1291);
nand U2241 (N_2241,N_844,N_1090);
and U2242 (N_2242,N_1438,N_1494);
or U2243 (N_2243,N_1480,N_1421);
nand U2244 (N_2244,N_990,N_936);
and U2245 (N_2245,N_1276,N_852);
or U2246 (N_2246,N_1410,N_1097);
and U2247 (N_2247,N_1140,N_1325);
xnor U2248 (N_2248,N_828,N_1480);
xor U2249 (N_2249,N_1020,N_934);
nand U2250 (N_2250,N_1826,N_1818);
or U2251 (N_2251,N_1979,N_1726);
or U2252 (N_2252,N_2137,N_1529);
or U2253 (N_2253,N_2227,N_1583);
or U2254 (N_2254,N_1517,N_1674);
or U2255 (N_2255,N_1736,N_2125);
nor U2256 (N_2256,N_1947,N_1924);
nand U2257 (N_2257,N_2210,N_2169);
nand U2258 (N_2258,N_2195,N_2171);
or U2259 (N_2259,N_1989,N_2203);
xor U2260 (N_2260,N_1602,N_1768);
nand U2261 (N_2261,N_1506,N_1860);
nor U2262 (N_2262,N_1510,N_1977);
nand U2263 (N_2263,N_1591,N_1821);
and U2264 (N_2264,N_1878,N_2035);
xnor U2265 (N_2265,N_1548,N_1737);
and U2266 (N_2266,N_1767,N_1573);
xnor U2267 (N_2267,N_1787,N_1663);
nor U2268 (N_2268,N_1556,N_1544);
nand U2269 (N_2269,N_2181,N_1961);
or U2270 (N_2270,N_2016,N_1533);
nand U2271 (N_2271,N_2060,N_1960);
or U2272 (N_2272,N_1953,N_1992);
nand U2273 (N_2273,N_1935,N_1746);
and U2274 (N_2274,N_1791,N_1797);
nor U2275 (N_2275,N_1714,N_1862);
nor U2276 (N_2276,N_1687,N_1630);
xor U2277 (N_2277,N_1608,N_1908);
or U2278 (N_2278,N_2116,N_1955);
nor U2279 (N_2279,N_2164,N_1537);
and U2280 (N_2280,N_1691,N_1643);
and U2281 (N_2281,N_1902,N_2220);
or U2282 (N_2282,N_1595,N_1628);
or U2283 (N_2283,N_1684,N_1887);
and U2284 (N_2284,N_1637,N_1766);
nand U2285 (N_2285,N_2108,N_2192);
xor U2286 (N_2286,N_1672,N_1567);
nor U2287 (N_2287,N_1799,N_2160);
nand U2288 (N_2288,N_1692,N_2003);
and U2289 (N_2289,N_1964,N_2061);
nor U2290 (N_2290,N_1871,N_2008);
and U2291 (N_2291,N_2162,N_1699);
and U2292 (N_2292,N_2165,N_1842);
and U2293 (N_2293,N_1632,N_1621);
xor U2294 (N_2294,N_1521,N_1718);
and U2295 (N_2295,N_2004,N_1694);
and U2296 (N_2296,N_2123,N_1706);
xnor U2297 (N_2297,N_2119,N_2026);
nand U2298 (N_2298,N_2244,N_1679);
nor U2299 (N_2299,N_2041,N_1807);
and U2300 (N_2300,N_1942,N_1557);
or U2301 (N_2301,N_1934,N_2063);
or U2302 (N_2302,N_2083,N_1614);
and U2303 (N_2303,N_2094,N_2110);
nand U2304 (N_2304,N_1783,N_1975);
nand U2305 (N_2305,N_1834,N_2229);
nor U2306 (N_2306,N_1764,N_2222);
or U2307 (N_2307,N_1893,N_1505);
nand U2308 (N_2308,N_2045,N_1816);
nor U2309 (N_2309,N_1833,N_1645);
and U2310 (N_2310,N_1617,N_2246);
nand U2311 (N_2311,N_2068,N_1541);
or U2312 (N_2312,N_1585,N_2019);
and U2313 (N_2313,N_1873,N_1864);
xor U2314 (N_2314,N_1748,N_2018);
and U2315 (N_2315,N_2212,N_1693);
and U2316 (N_2316,N_1732,N_1677);
and U2317 (N_2317,N_1530,N_1671);
nor U2318 (N_2318,N_1929,N_1911);
and U2319 (N_2319,N_2052,N_2226);
nor U2320 (N_2320,N_1644,N_1782);
nor U2321 (N_2321,N_1755,N_1571);
nand U2322 (N_2322,N_1555,N_1713);
xor U2323 (N_2323,N_2039,N_1523);
or U2324 (N_2324,N_1622,N_1612);
xor U2325 (N_2325,N_1963,N_1788);
xnor U2326 (N_2326,N_1669,N_1804);
nor U2327 (N_2327,N_1638,N_1972);
xnor U2328 (N_2328,N_1962,N_1828);
nand U2329 (N_2329,N_1519,N_1627);
and U2330 (N_2330,N_2077,N_1577);
or U2331 (N_2331,N_1906,N_1957);
or U2332 (N_2332,N_1666,N_1550);
and U2333 (N_2333,N_2175,N_1905);
nand U2334 (N_2334,N_1656,N_2059);
and U2335 (N_2335,N_2170,N_1681);
and U2336 (N_2336,N_1938,N_2231);
or U2337 (N_2337,N_1922,N_1763);
nand U2338 (N_2338,N_1704,N_2032);
or U2339 (N_2339,N_1970,N_1985);
or U2340 (N_2340,N_1697,N_1610);
nor U2341 (N_2341,N_2146,N_1940);
and U2342 (N_2342,N_1615,N_1852);
nor U2343 (N_2343,N_2188,N_2058);
or U2344 (N_2344,N_2000,N_2030);
or U2345 (N_2345,N_1786,N_1832);
or U2346 (N_2346,N_1877,N_1798);
and U2347 (N_2347,N_1855,N_1857);
nand U2348 (N_2348,N_2109,N_1631);
nor U2349 (N_2349,N_1731,N_2036);
and U2350 (N_2350,N_1520,N_2071);
nand U2351 (N_2351,N_2033,N_2102);
or U2352 (N_2352,N_2107,N_1849);
and U2353 (N_2353,N_1626,N_2152);
and U2354 (N_2354,N_2114,N_1965);
nand U2355 (N_2355,N_2075,N_1512);
nand U2356 (N_2356,N_1946,N_2135);
nand U2357 (N_2357,N_2213,N_1507);
nor U2358 (N_2358,N_2242,N_1664);
or U2359 (N_2359,N_2245,N_1894);
nor U2360 (N_2360,N_1662,N_1721);
and U2361 (N_2361,N_1995,N_1760);
and U2362 (N_2362,N_2104,N_1884);
nand U2363 (N_2363,N_1647,N_1733);
nand U2364 (N_2364,N_2073,N_1657);
or U2365 (N_2365,N_2219,N_1723);
nor U2366 (N_2366,N_2120,N_2134);
or U2367 (N_2367,N_1619,N_2141);
nand U2368 (N_2368,N_2122,N_1785);
nand U2369 (N_2369,N_1700,N_1812);
and U2370 (N_2370,N_1969,N_1921);
nor U2371 (N_2371,N_1903,N_1604);
nand U2372 (N_2372,N_2022,N_1527);
and U2373 (N_2373,N_1729,N_1870);
nand U2374 (N_2374,N_2067,N_2236);
and U2375 (N_2375,N_1954,N_1897);
or U2376 (N_2376,N_2084,N_1830);
xor U2377 (N_2377,N_1711,N_1735);
and U2378 (N_2378,N_2194,N_1745);
nor U2379 (N_2379,N_1620,N_2124);
or U2380 (N_2380,N_1844,N_2157);
or U2381 (N_2381,N_2012,N_1971);
or U2382 (N_2382,N_1837,N_1931);
nand U2383 (N_2383,N_1850,N_1918);
nand U2384 (N_2384,N_1728,N_1588);
nor U2385 (N_2385,N_1686,N_1930);
or U2386 (N_2386,N_1705,N_1784);
nor U2387 (N_2387,N_2193,N_1559);
nand U2388 (N_2388,N_2190,N_1915);
or U2389 (N_2389,N_1659,N_1951);
nand U2390 (N_2390,N_2156,N_1890);
nor U2391 (N_2391,N_2002,N_1720);
nand U2392 (N_2392,N_2034,N_1685);
nand U2393 (N_2393,N_1606,N_1593);
nand U2394 (N_2394,N_2099,N_1762);
and U2395 (N_2395,N_1866,N_1993);
nor U2396 (N_2396,N_1561,N_1682);
nand U2397 (N_2397,N_1534,N_1562);
nor U2398 (N_2398,N_2015,N_1531);
and U2399 (N_2399,N_1936,N_1625);
nand U2400 (N_2400,N_1611,N_2158);
and U2401 (N_2401,N_1725,N_1769);
nand U2402 (N_2402,N_1802,N_1859);
and U2403 (N_2403,N_1563,N_1817);
nor U2404 (N_2404,N_2209,N_1670);
and U2405 (N_2405,N_2100,N_1978);
nor U2406 (N_2406,N_1564,N_1819);
nand U2407 (N_2407,N_1886,N_2147);
nand U2408 (N_2408,N_2153,N_1539);
xnor U2409 (N_2409,N_1543,N_2074);
and U2410 (N_2410,N_2148,N_2183);
or U2411 (N_2411,N_1803,N_1920);
nor U2412 (N_2412,N_1795,N_1554);
and U2413 (N_2413,N_1917,N_1503);
nor U2414 (N_2414,N_1854,N_1904);
or U2415 (N_2415,N_2054,N_2239);
nand U2416 (N_2416,N_1820,N_1513);
xor U2417 (N_2417,N_1914,N_1727);
nor U2418 (N_2418,N_1761,N_1605);
and U2419 (N_2419,N_2009,N_1973);
and U2420 (N_2420,N_1771,N_1586);
or U2421 (N_2421,N_2224,N_1990);
nor U2422 (N_2422,N_2031,N_1765);
nor U2423 (N_2423,N_1508,N_1629);
or U2424 (N_2424,N_2096,N_1640);
nor U2425 (N_2425,N_1966,N_1623);
nor U2426 (N_2426,N_1509,N_2218);
nand U2427 (N_2427,N_1590,N_1758);
nand U2428 (N_2428,N_2053,N_2180);
and U2429 (N_2429,N_1879,N_2248);
nor U2430 (N_2430,N_1825,N_1809);
nor U2431 (N_2431,N_1635,N_2066);
nor U2432 (N_2432,N_1851,N_1853);
or U2433 (N_2433,N_1861,N_2230);
nor U2434 (N_2434,N_1649,N_2021);
and U2435 (N_2435,N_1982,N_1780);
and U2436 (N_2436,N_1532,N_2235);
nand U2437 (N_2437,N_2121,N_2082);
and U2438 (N_2438,N_1909,N_1945);
nand U2439 (N_2439,N_1724,N_1941);
xor U2440 (N_2440,N_1998,N_1575);
nand U2441 (N_2441,N_1542,N_1739);
and U2442 (N_2442,N_1757,N_1813);
nand U2443 (N_2443,N_2225,N_1968);
xnor U2444 (N_2444,N_2070,N_1883);
and U2445 (N_2445,N_1545,N_1944);
and U2446 (N_2446,N_2241,N_1937);
nand U2447 (N_2447,N_2144,N_1843);
nand U2448 (N_2448,N_2161,N_2072);
and U2449 (N_2449,N_1863,N_1948);
nand U2450 (N_2450,N_2106,N_1753);
or U2451 (N_2451,N_2143,N_1584);
nor U2452 (N_2452,N_2081,N_2043);
and U2453 (N_2453,N_2129,N_1715);
or U2454 (N_2454,N_1609,N_2025);
or U2455 (N_2455,N_1880,N_1540);
nand U2456 (N_2456,N_2178,N_1808);
and U2457 (N_2457,N_1774,N_1933);
nor U2458 (N_2458,N_1695,N_2208);
or U2459 (N_2459,N_1829,N_2095);
nor U2460 (N_2460,N_2130,N_2127);
and U2461 (N_2461,N_1996,N_1698);
nand U2462 (N_2462,N_1578,N_2056);
nand U2463 (N_2463,N_1815,N_1675);
xor U2464 (N_2464,N_1689,N_1574);
or U2465 (N_2465,N_1589,N_1927);
or U2466 (N_2466,N_2133,N_1999);
nand U2467 (N_2467,N_1709,N_2184);
or U2468 (N_2468,N_2204,N_1892);
xnor U2469 (N_2469,N_1781,N_1553);
or U2470 (N_2470,N_1881,N_1889);
nand U2471 (N_2471,N_1566,N_1839);
or U2472 (N_2472,N_1653,N_1516);
nand U2473 (N_2473,N_2040,N_1949);
nand U2474 (N_2474,N_1518,N_1702);
nor U2475 (N_2475,N_1717,N_1738);
nor U2476 (N_2476,N_1901,N_1565);
nor U2477 (N_2477,N_1525,N_1551);
and U2478 (N_2478,N_1734,N_1740);
nand U2479 (N_2479,N_1668,N_2199);
xnor U2480 (N_2480,N_2051,N_2089);
and U2481 (N_2481,N_1896,N_2044);
or U2482 (N_2482,N_2017,N_2042);
nand U2483 (N_2483,N_2149,N_2233);
nor U2484 (N_2484,N_1576,N_1607);
and U2485 (N_2485,N_1660,N_1919);
or U2486 (N_2486,N_1501,N_2014);
nand U2487 (N_2487,N_1618,N_1750);
nand U2488 (N_2488,N_1703,N_1823);
nor U2489 (N_2489,N_2189,N_1504);
and U2490 (N_2490,N_1912,N_1810);
xor U2491 (N_2491,N_1654,N_1558);
nor U2492 (N_2492,N_2069,N_1974);
nand U2493 (N_2493,N_1658,N_2001);
or U2494 (N_2494,N_2028,N_1596);
or U2495 (N_2495,N_1747,N_1744);
or U2496 (N_2496,N_2215,N_1676);
or U2497 (N_2497,N_2132,N_1742);
nand U2498 (N_2498,N_1549,N_1950);
nor U2499 (N_2499,N_1661,N_2047);
nor U2500 (N_2500,N_1641,N_2177);
nor U2501 (N_2501,N_1624,N_1932);
nor U2502 (N_2502,N_2191,N_2176);
or U2503 (N_2503,N_1526,N_2216);
and U2504 (N_2504,N_1546,N_1582);
nor U2505 (N_2505,N_1984,N_1865);
nor U2506 (N_2506,N_2023,N_2007);
nor U2507 (N_2507,N_1789,N_1800);
nand U2508 (N_2508,N_1848,N_2247);
and U2509 (N_2509,N_1683,N_1592);
nand U2510 (N_2510,N_1888,N_2145);
or U2511 (N_2511,N_1722,N_1958);
nor U2512 (N_2512,N_1667,N_2185);
nor U2513 (N_2513,N_2234,N_2038);
and U2514 (N_2514,N_1775,N_2172);
or U2515 (N_2515,N_1570,N_2159);
xor U2516 (N_2516,N_2238,N_1603);
and U2517 (N_2517,N_2010,N_1708);
xnor U2518 (N_2518,N_1655,N_2037);
nor U2519 (N_2519,N_1794,N_1868);
or U2520 (N_2520,N_1874,N_2186);
nor U2521 (N_2521,N_1840,N_1569);
and U2522 (N_2522,N_1613,N_1600);
xnor U2523 (N_2523,N_1847,N_1594);
or U2524 (N_2524,N_2112,N_1925);
nor U2525 (N_2525,N_2049,N_2011);
and U2526 (N_2526,N_1811,N_2166);
or U2527 (N_2527,N_1778,N_1956);
nand U2528 (N_2528,N_1712,N_1882);
nand U2529 (N_2529,N_1943,N_1898);
or U2530 (N_2530,N_1678,N_1997);
xnor U2531 (N_2531,N_2221,N_1579);
nor U2532 (N_2532,N_1749,N_1772);
or U2533 (N_2533,N_2173,N_1568);
nand U2534 (N_2534,N_2128,N_1680);
and U2535 (N_2535,N_2200,N_1587);
or U2536 (N_2536,N_1856,N_1967);
or U2537 (N_2537,N_1822,N_1976);
nand U2538 (N_2538,N_1899,N_1926);
nand U2539 (N_2539,N_2101,N_2240);
nor U2540 (N_2540,N_1988,N_2167);
or U2541 (N_2541,N_2005,N_2064);
nor U2542 (N_2542,N_1779,N_2086);
and U2543 (N_2543,N_1547,N_1876);
nand U2544 (N_2544,N_1845,N_1831);
or U2545 (N_2545,N_1636,N_2105);
nor U2546 (N_2546,N_2154,N_1777);
and U2547 (N_2547,N_1846,N_2020);
and U2548 (N_2548,N_2006,N_2080);
nor U2549 (N_2549,N_2237,N_1756);
or U2550 (N_2550,N_2151,N_1601);
nand U2551 (N_2551,N_1616,N_1502);
and U2552 (N_2552,N_1528,N_2078);
and U2553 (N_2553,N_1959,N_1875);
xor U2554 (N_2554,N_2113,N_2046);
nand U2555 (N_2555,N_1633,N_1754);
nand U2556 (N_2556,N_2050,N_1923);
or U2557 (N_2557,N_1867,N_2088);
or U2558 (N_2558,N_1980,N_1952);
nand U2559 (N_2559,N_1690,N_1648);
and U2560 (N_2560,N_1524,N_1719);
nand U2561 (N_2561,N_1752,N_1814);
or U2562 (N_2562,N_2249,N_2048);
nor U2563 (N_2563,N_2163,N_2087);
or U2564 (N_2564,N_1696,N_1646);
nand U2565 (N_2565,N_1872,N_2228);
and U2566 (N_2566,N_1827,N_2055);
nor U2567 (N_2567,N_1560,N_1916);
nand U2568 (N_2568,N_2065,N_1891);
nor U2569 (N_2569,N_1599,N_1716);
xnor U2570 (N_2570,N_2142,N_1522);
nand U2571 (N_2571,N_1650,N_2027);
and U2572 (N_2572,N_1652,N_2196);
or U2573 (N_2573,N_2155,N_1580);
and U2574 (N_2574,N_1869,N_2205);
xnor U2575 (N_2575,N_1536,N_2217);
and U2576 (N_2576,N_2062,N_1981);
and U2577 (N_2577,N_1598,N_2126);
nor U2578 (N_2578,N_2057,N_1515);
nor U2579 (N_2579,N_2140,N_2111);
nor U2580 (N_2580,N_2201,N_1838);
nand U2581 (N_2581,N_1751,N_1900);
and U2582 (N_2582,N_1792,N_1581);
nand U2583 (N_2583,N_1651,N_2197);
nor U2584 (N_2584,N_2090,N_1986);
and U2585 (N_2585,N_1885,N_1836);
and U2586 (N_2586,N_1913,N_2232);
nor U2587 (N_2587,N_2117,N_2206);
nor U2588 (N_2588,N_2202,N_1790);
or U2589 (N_2589,N_1910,N_1673);
or U2590 (N_2590,N_1597,N_2168);
nand U2591 (N_2591,N_2187,N_1987);
and U2592 (N_2592,N_2243,N_1538);
nor U2593 (N_2593,N_1514,N_1824);
or U2594 (N_2594,N_2076,N_2211);
xnor U2595 (N_2595,N_2097,N_1773);
nor U2596 (N_2596,N_2138,N_2198);
and U2597 (N_2597,N_2174,N_1806);
and U2598 (N_2598,N_1776,N_2139);
nand U2599 (N_2599,N_1907,N_2013);
xor U2600 (N_2600,N_1805,N_1793);
nand U2601 (N_2601,N_2091,N_1743);
nor U2602 (N_2602,N_1759,N_2092);
nor U2603 (N_2603,N_1730,N_1535);
nand U2604 (N_2604,N_1642,N_2150);
nor U2605 (N_2605,N_2024,N_2098);
or U2606 (N_2606,N_1710,N_1983);
or U2607 (N_2607,N_1707,N_1639);
or U2608 (N_2608,N_1665,N_2131);
or U2609 (N_2609,N_1634,N_2115);
and U2610 (N_2610,N_1796,N_2093);
xnor U2611 (N_2611,N_2029,N_1572);
nor U2612 (N_2612,N_1500,N_2079);
and U2613 (N_2613,N_1741,N_2207);
or U2614 (N_2614,N_1994,N_1552);
xnor U2615 (N_2615,N_1841,N_1770);
and U2616 (N_2616,N_1895,N_1801);
or U2617 (N_2617,N_1858,N_2136);
nor U2618 (N_2618,N_2182,N_1835);
and U2619 (N_2619,N_2223,N_1511);
and U2620 (N_2620,N_2179,N_1688);
xnor U2621 (N_2621,N_1701,N_1939);
xnor U2622 (N_2622,N_1928,N_1991);
nor U2623 (N_2623,N_2214,N_2103);
or U2624 (N_2624,N_2085,N_2118);
and U2625 (N_2625,N_1992,N_1947);
or U2626 (N_2626,N_2148,N_1888);
nor U2627 (N_2627,N_1889,N_1526);
nor U2628 (N_2628,N_1830,N_1930);
xor U2629 (N_2629,N_1888,N_2220);
or U2630 (N_2630,N_1880,N_2207);
or U2631 (N_2631,N_1844,N_1848);
and U2632 (N_2632,N_2071,N_2113);
nand U2633 (N_2633,N_1566,N_2182);
or U2634 (N_2634,N_1969,N_2042);
nor U2635 (N_2635,N_1886,N_1780);
nor U2636 (N_2636,N_1913,N_1631);
and U2637 (N_2637,N_1753,N_2018);
nand U2638 (N_2638,N_1637,N_1944);
xnor U2639 (N_2639,N_1666,N_1549);
xor U2640 (N_2640,N_2053,N_1573);
or U2641 (N_2641,N_1515,N_1661);
and U2642 (N_2642,N_2131,N_1500);
xnor U2643 (N_2643,N_2144,N_1994);
and U2644 (N_2644,N_1582,N_1911);
or U2645 (N_2645,N_2193,N_2134);
xnor U2646 (N_2646,N_1803,N_1515);
or U2647 (N_2647,N_1698,N_1788);
nand U2648 (N_2648,N_2207,N_2200);
nor U2649 (N_2649,N_1958,N_2091);
nand U2650 (N_2650,N_1520,N_1890);
nand U2651 (N_2651,N_2144,N_1931);
nand U2652 (N_2652,N_1633,N_1904);
nand U2653 (N_2653,N_2215,N_1519);
nand U2654 (N_2654,N_1991,N_2190);
or U2655 (N_2655,N_1533,N_2060);
nand U2656 (N_2656,N_2103,N_1892);
nor U2657 (N_2657,N_1696,N_1590);
nor U2658 (N_2658,N_2230,N_1672);
or U2659 (N_2659,N_1624,N_2236);
and U2660 (N_2660,N_1893,N_1738);
xnor U2661 (N_2661,N_1650,N_1647);
nand U2662 (N_2662,N_1634,N_1922);
and U2663 (N_2663,N_1720,N_2182);
nor U2664 (N_2664,N_1546,N_1866);
and U2665 (N_2665,N_2219,N_2017);
or U2666 (N_2666,N_2142,N_1707);
xor U2667 (N_2667,N_1758,N_2117);
xnor U2668 (N_2668,N_2024,N_1868);
xnor U2669 (N_2669,N_1772,N_1966);
xor U2670 (N_2670,N_1571,N_1509);
nand U2671 (N_2671,N_1509,N_1799);
or U2672 (N_2672,N_1942,N_2130);
and U2673 (N_2673,N_2203,N_2178);
nand U2674 (N_2674,N_1736,N_2209);
nor U2675 (N_2675,N_1852,N_1609);
xnor U2676 (N_2676,N_1763,N_2223);
or U2677 (N_2677,N_1759,N_1569);
nand U2678 (N_2678,N_2083,N_2126);
nand U2679 (N_2679,N_1900,N_2147);
nand U2680 (N_2680,N_1586,N_1823);
nor U2681 (N_2681,N_1784,N_1956);
nor U2682 (N_2682,N_1505,N_1822);
nor U2683 (N_2683,N_1619,N_1905);
nor U2684 (N_2684,N_1630,N_1541);
nand U2685 (N_2685,N_1580,N_1900);
nor U2686 (N_2686,N_2131,N_2015);
nand U2687 (N_2687,N_1968,N_1784);
and U2688 (N_2688,N_1794,N_1748);
nor U2689 (N_2689,N_1949,N_2205);
nand U2690 (N_2690,N_2195,N_1869);
and U2691 (N_2691,N_1824,N_1582);
nand U2692 (N_2692,N_1665,N_1600);
and U2693 (N_2693,N_1628,N_1569);
nand U2694 (N_2694,N_1992,N_1771);
and U2695 (N_2695,N_2078,N_1994);
xnor U2696 (N_2696,N_2150,N_2130);
and U2697 (N_2697,N_1677,N_2175);
nand U2698 (N_2698,N_1701,N_2089);
and U2699 (N_2699,N_1923,N_1813);
nor U2700 (N_2700,N_2117,N_1932);
xnor U2701 (N_2701,N_1933,N_2027);
and U2702 (N_2702,N_2080,N_1919);
or U2703 (N_2703,N_1608,N_1975);
or U2704 (N_2704,N_2096,N_1822);
or U2705 (N_2705,N_1719,N_1506);
nor U2706 (N_2706,N_1597,N_2206);
or U2707 (N_2707,N_1648,N_1910);
nor U2708 (N_2708,N_2249,N_1682);
nand U2709 (N_2709,N_1755,N_1814);
or U2710 (N_2710,N_1958,N_1897);
or U2711 (N_2711,N_2240,N_1591);
nor U2712 (N_2712,N_1972,N_2092);
nand U2713 (N_2713,N_1764,N_1570);
or U2714 (N_2714,N_1690,N_1618);
and U2715 (N_2715,N_2185,N_2133);
nand U2716 (N_2716,N_1585,N_2087);
nor U2717 (N_2717,N_1744,N_1937);
and U2718 (N_2718,N_2131,N_1616);
and U2719 (N_2719,N_1674,N_2060);
or U2720 (N_2720,N_1582,N_2113);
nor U2721 (N_2721,N_1879,N_2063);
and U2722 (N_2722,N_1898,N_2169);
nand U2723 (N_2723,N_1612,N_2205);
and U2724 (N_2724,N_1865,N_2129);
and U2725 (N_2725,N_2142,N_2057);
nand U2726 (N_2726,N_1746,N_1812);
and U2727 (N_2727,N_1751,N_2128);
nor U2728 (N_2728,N_1951,N_1750);
xnor U2729 (N_2729,N_1966,N_1590);
nor U2730 (N_2730,N_1928,N_1569);
nor U2731 (N_2731,N_1755,N_1779);
and U2732 (N_2732,N_1784,N_1688);
and U2733 (N_2733,N_1720,N_1550);
or U2734 (N_2734,N_1547,N_1679);
nor U2735 (N_2735,N_1772,N_1874);
nand U2736 (N_2736,N_1618,N_1663);
nand U2737 (N_2737,N_1945,N_1530);
nor U2738 (N_2738,N_1858,N_1882);
xnor U2739 (N_2739,N_1980,N_1614);
nor U2740 (N_2740,N_1759,N_1823);
nand U2741 (N_2741,N_2106,N_2005);
nor U2742 (N_2742,N_1847,N_2098);
and U2743 (N_2743,N_1973,N_1943);
or U2744 (N_2744,N_2238,N_2105);
nand U2745 (N_2745,N_1884,N_1675);
or U2746 (N_2746,N_2105,N_1740);
nor U2747 (N_2747,N_2127,N_1618);
nand U2748 (N_2748,N_2001,N_1741);
nand U2749 (N_2749,N_1665,N_2054);
and U2750 (N_2750,N_1999,N_1946);
nor U2751 (N_2751,N_2168,N_2161);
and U2752 (N_2752,N_1746,N_1771);
or U2753 (N_2753,N_1884,N_1666);
nor U2754 (N_2754,N_1509,N_1988);
and U2755 (N_2755,N_1791,N_1545);
and U2756 (N_2756,N_2145,N_2111);
nor U2757 (N_2757,N_2004,N_2080);
or U2758 (N_2758,N_1541,N_1659);
or U2759 (N_2759,N_2102,N_1991);
nand U2760 (N_2760,N_1661,N_1765);
and U2761 (N_2761,N_1887,N_2108);
nand U2762 (N_2762,N_2037,N_1529);
and U2763 (N_2763,N_1840,N_1953);
and U2764 (N_2764,N_2228,N_1879);
or U2765 (N_2765,N_1594,N_1860);
or U2766 (N_2766,N_1777,N_2074);
nor U2767 (N_2767,N_1564,N_1985);
nand U2768 (N_2768,N_1903,N_2075);
and U2769 (N_2769,N_1937,N_2150);
nand U2770 (N_2770,N_2042,N_1648);
nor U2771 (N_2771,N_1918,N_1756);
nor U2772 (N_2772,N_1901,N_1644);
xnor U2773 (N_2773,N_1734,N_1889);
or U2774 (N_2774,N_1792,N_1579);
or U2775 (N_2775,N_2009,N_1527);
nor U2776 (N_2776,N_1747,N_2026);
and U2777 (N_2777,N_1932,N_2062);
xnor U2778 (N_2778,N_2165,N_1662);
nor U2779 (N_2779,N_2119,N_1726);
or U2780 (N_2780,N_1778,N_2125);
nand U2781 (N_2781,N_1526,N_1613);
or U2782 (N_2782,N_1554,N_2244);
nor U2783 (N_2783,N_1648,N_1602);
nand U2784 (N_2784,N_2102,N_2050);
nor U2785 (N_2785,N_2072,N_1852);
and U2786 (N_2786,N_1998,N_1538);
or U2787 (N_2787,N_1557,N_2178);
nor U2788 (N_2788,N_2023,N_1997);
nand U2789 (N_2789,N_2171,N_1597);
nor U2790 (N_2790,N_2017,N_1971);
and U2791 (N_2791,N_2247,N_1659);
and U2792 (N_2792,N_1891,N_1631);
xnor U2793 (N_2793,N_1671,N_1852);
nand U2794 (N_2794,N_2207,N_2136);
nand U2795 (N_2795,N_1920,N_1851);
or U2796 (N_2796,N_1909,N_1803);
and U2797 (N_2797,N_1681,N_1784);
xor U2798 (N_2798,N_1822,N_1609);
and U2799 (N_2799,N_2123,N_1844);
or U2800 (N_2800,N_1950,N_1572);
nand U2801 (N_2801,N_1588,N_1623);
nand U2802 (N_2802,N_1973,N_2241);
nand U2803 (N_2803,N_1507,N_1807);
and U2804 (N_2804,N_1814,N_1507);
xnor U2805 (N_2805,N_1900,N_1654);
nor U2806 (N_2806,N_2020,N_1634);
or U2807 (N_2807,N_1999,N_1858);
xnor U2808 (N_2808,N_2231,N_2062);
nor U2809 (N_2809,N_1992,N_1784);
and U2810 (N_2810,N_1642,N_2243);
and U2811 (N_2811,N_1701,N_2244);
or U2812 (N_2812,N_2024,N_1943);
and U2813 (N_2813,N_1586,N_2141);
and U2814 (N_2814,N_1669,N_1817);
nor U2815 (N_2815,N_1546,N_1755);
or U2816 (N_2816,N_1523,N_1990);
nor U2817 (N_2817,N_2136,N_2003);
and U2818 (N_2818,N_2047,N_2223);
and U2819 (N_2819,N_1706,N_2026);
xnor U2820 (N_2820,N_1798,N_1879);
nand U2821 (N_2821,N_1601,N_2091);
nand U2822 (N_2822,N_1555,N_2237);
and U2823 (N_2823,N_1638,N_1886);
nor U2824 (N_2824,N_1817,N_2160);
or U2825 (N_2825,N_2065,N_2222);
or U2826 (N_2826,N_1566,N_1778);
nor U2827 (N_2827,N_2067,N_1663);
and U2828 (N_2828,N_2167,N_1821);
nand U2829 (N_2829,N_1526,N_2089);
or U2830 (N_2830,N_1790,N_1553);
nand U2831 (N_2831,N_1506,N_2046);
nor U2832 (N_2832,N_2023,N_1819);
and U2833 (N_2833,N_1708,N_1796);
and U2834 (N_2834,N_2169,N_1970);
and U2835 (N_2835,N_1514,N_1522);
nand U2836 (N_2836,N_1522,N_1534);
nand U2837 (N_2837,N_1739,N_1554);
and U2838 (N_2838,N_2101,N_2001);
or U2839 (N_2839,N_2039,N_1615);
nor U2840 (N_2840,N_1631,N_2235);
and U2841 (N_2841,N_2221,N_1614);
nand U2842 (N_2842,N_1576,N_1778);
xnor U2843 (N_2843,N_1838,N_2066);
nand U2844 (N_2844,N_1833,N_1767);
or U2845 (N_2845,N_1709,N_2140);
and U2846 (N_2846,N_1623,N_1568);
nand U2847 (N_2847,N_2043,N_1600);
or U2848 (N_2848,N_1574,N_1972);
nand U2849 (N_2849,N_1823,N_1903);
nand U2850 (N_2850,N_1650,N_2033);
and U2851 (N_2851,N_2046,N_1752);
nor U2852 (N_2852,N_2027,N_2243);
or U2853 (N_2853,N_1562,N_1665);
and U2854 (N_2854,N_1812,N_2030);
and U2855 (N_2855,N_1685,N_1895);
nand U2856 (N_2856,N_1969,N_1652);
and U2857 (N_2857,N_2064,N_1621);
xor U2858 (N_2858,N_1685,N_1818);
or U2859 (N_2859,N_2027,N_1999);
nand U2860 (N_2860,N_2035,N_1898);
xnor U2861 (N_2861,N_1530,N_1641);
xnor U2862 (N_2862,N_1565,N_1860);
and U2863 (N_2863,N_1501,N_1728);
nor U2864 (N_2864,N_1944,N_2239);
or U2865 (N_2865,N_2109,N_2045);
nor U2866 (N_2866,N_1722,N_2193);
or U2867 (N_2867,N_1731,N_2045);
and U2868 (N_2868,N_2036,N_2032);
and U2869 (N_2869,N_1817,N_1765);
and U2870 (N_2870,N_1983,N_1987);
nor U2871 (N_2871,N_1698,N_2028);
nor U2872 (N_2872,N_1604,N_1533);
or U2873 (N_2873,N_1547,N_1783);
or U2874 (N_2874,N_1548,N_1617);
xor U2875 (N_2875,N_1654,N_1503);
nand U2876 (N_2876,N_1576,N_2079);
or U2877 (N_2877,N_1560,N_1653);
and U2878 (N_2878,N_1603,N_1553);
or U2879 (N_2879,N_1864,N_1734);
nor U2880 (N_2880,N_1607,N_1929);
or U2881 (N_2881,N_1597,N_2140);
nand U2882 (N_2882,N_1543,N_1929);
or U2883 (N_2883,N_1541,N_1519);
or U2884 (N_2884,N_1796,N_1731);
or U2885 (N_2885,N_1839,N_1856);
nor U2886 (N_2886,N_1924,N_1604);
or U2887 (N_2887,N_1653,N_1583);
or U2888 (N_2888,N_1686,N_2161);
nand U2889 (N_2889,N_2044,N_1744);
xnor U2890 (N_2890,N_1842,N_1936);
or U2891 (N_2891,N_1827,N_1742);
nand U2892 (N_2892,N_1701,N_1957);
xnor U2893 (N_2893,N_1879,N_1571);
xor U2894 (N_2894,N_2167,N_1782);
nand U2895 (N_2895,N_1883,N_1632);
nand U2896 (N_2896,N_2045,N_1862);
or U2897 (N_2897,N_1991,N_1964);
nand U2898 (N_2898,N_1536,N_1612);
nor U2899 (N_2899,N_1652,N_1673);
nor U2900 (N_2900,N_1634,N_1670);
nor U2901 (N_2901,N_2041,N_2165);
nor U2902 (N_2902,N_2141,N_1615);
nand U2903 (N_2903,N_1819,N_2058);
nand U2904 (N_2904,N_2035,N_2091);
nand U2905 (N_2905,N_1805,N_2054);
or U2906 (N_2906,N_1870,N_2053);
nor U2907 (N_2907,N_1769,N_1610);
xor U2908 (N_2908,N_1560,N_1771);
and U2909 (N_2909,N_1943,N_2058);
nor U2910 (N_2910,N_1910,N_2091);
and U2911 (N_2911,N_2188,N_2144);
xor U2912 (N_2912,N_2241,N_1594);
nor U2913 (N_2913,N_2072,N_2017);
nand U2914 (N_2914,N_2064,N_2047);
and U2915 (N_2915,N_1855,N_1591);
or U2916 (N_2916,N_1778,N_2247);
nand U2917 (N_2917,N_2238,N_1767);
and U2918 (N_2918,N_1711,N_1627);
nand U2919 (N_2919,N_1631,N_2140);
and U2920 (N_2920,N_1943,N_2086);
or U2921 (N_2921,N_2161,N_1863);
or U2922 (N_2922,N_2183,N_2110);
and U2923 (N_2923,N_1745,N_2037);
nand U2924 (N_2924,N_1503,N_2045);
xnor U2925 (N_2925,N_1956,N_1510);
xnor U2926 (N_2926,N_1974,N_1989);
nor U2927 (N_2927,N_1745,N_1743);
and U2928 (N_2928,N_2134,N_2080);
or U2929 (N_2929,N_2026,N_2128);
nor U2930 (N_2930,N_1794,N_2068);
or U2931 (N_2931,N_1963,N_2082);
nand U2932 (N_2932,N_1658,N_1547);
nor U2933 (N_2933,N_1839,N_1726);
nand U2934 (N_2934,N_1817,N_1557);
or U2935 (N_2935,N_1607,N_1617);
and U2936 (N_2936,N_1556,N_1789);
nor U2937 (N_2937,N_1870,N_1912);
nor U2938 (N_2938,N_1718,N_1794);
nand U2939 (N_2939,N_1964,N_1583);
and U2940 (N_2940,N_1620,N_1546);
nand U2941 (N_2941,N_2202,N_2155);
and U2942 (N_2942,N_1522,N_2170);
nand U2943 (N_2943,N_1631,N_1790);
and U2944 (N_2944,N_1751,N_1668);
nor U2945 (N_2945,N_2023,N_1589);
and U2946 (N_2946,N_1677,N_1537);
nor U2947 (N_2947,N_1559,N_1615);
or U2948 (N_2948,N_1821,N_1951);
nor U2949 (N_2949,N_2207,N_1876);
nand U2950 (N_2950,N_1702,N_1619);
nand U2951 (N_2951,N_2154,N_2100);
or U2952 (N_2952,N_1762,N_1947);
nand U2953 (N_2953,N_1893,N_1974);
and U2954 (N_2954,N_1703,N_1757);
nand U2955 (N_2955,N_1687,N_1775);
nor U2956 (N_2956,N_1566,N_2141);
nand U2957 (N_2957,N_2199,N_1553);
and U2958 (N_2958,N_2019,N_1659);
and U2959 (N_2959,N_1766,N_1660);
nor U2960 (N_2960,N_2068,N_1945);
or U2961 (N_2961,N_1899,N_1728);
or U2962 (N_2962,N_2033,N_1698);
and U2963 (N_2963,N_2102,N_2060);
and U2964 (N_2964,N_2242,N_1950);
xnor U2965 (N_2965,N_2083,N_2235);
nor U2966 (N_2966,N_2085,N_1703);
xor U2967 (N_2967,N_2202,N_2179);
xor U2968 (N_2968,N_2061,N_1674);
nand U2969 (N_2969,N_2075,N_1660);
and U2970 (N_2970,N_2038,N_2240);
xnor U2971 (N_2971,N_2236,N_2235);
nand U2972 (N_2972,N_2007,N_1564);
or U2973 (N_2973,N_1977,N_2238);
or U2974 (N_2974,N_1815,N_1693);
or U2975 (N_2975,N_1886,N_2012);
or U2976 (N_2976,N_2085,N_1647);
or U2977 (N_2977,N_2249,N_1507);
or U2978 (N_2978,N_1506,N_1503);
nor U2979 (N_2979,N_1841,N_2139);
nand U2980 (N_2980,N_1992,N_1521);
nand U2981 (N_2981,N_1554,N_2177);
nor U2982 (N_2982,N_1818,N_2027);
xor U2983 (N_2983,N_2057,N_2024);
nand U2984 (N_2984,N_1935,N_1986);
or U2985 (N_2985,N_1888,N_1932);
xor U2986 (N_2986,N_2016,N_2137);
nand U2987 (N_2987,N_1828,N_1569);
xnor U2988 (N_2988,N_1691,N_2129);
nand U2989 (N_2989,N_2053,N_1534);
nand U2990 (N_2990,N_1528,N_1883);
nor U2991 (N_2991,N_1932,N_1806);
nor U2992 (N_2992,N_1558,N_1800);
xnor U2993 (N_2993,N_1817,N_2121);
and U2994 (N_2994,N_1676,N_2221);
nand U2995 (N_2995,N_1526,N_1798);
nand U2996 (N_2996,N_1904,N_1829);
nand U2997 (N_2997,N_1693,N_1618);
or U2998 (N_2998,N_1634,N_1682);
and U2999 (N_2999,N_2009,N_1792);
and UO_0 (O_0,N_2489,N_2673);
nor UO_1 (O_1,N_2805,N_2779);
and UO_2 (O_2,N_2338,N_2789);
nor UO_3 (O_3,N_2927,N_2409);
xor UO_4 (O_4,N_2833,N_2456);
or UO_5 (O_5,N_2413,N_2497);
and UO_6 (O_6,N_2374,N_2990);
nand UO_7 (O_7,N_2555,N_2324);
xor UO_8 (O_8,N_2457,N_2751);
nor UO_9 (O_9,N_2542,N_2634);
and UO_10 (O_10,N_2523,N_2276);
nor UO_11 (O_11,N_2577,N_2871);
nand UO_12 (O_12,N_2788,N_2704);
and UO_13 (O_13,N_2652,N_2628);
nor UO_14 (O_14,N_2358,N_2316);
nor UO_15 (O_15,N_2705,N_2425);
xnor UO_16 (O_16,N_2662,N_2718);
and UO_17 (O_17,N_2441,N_2916);
nand UO_18 (O_18,N_2414,N_2514);
and UO_19 (O_19,N_2430,N_2627);
nand UO_20 (O_20,N_2560,N_2888);
xnor UO_21 (O_21,N_2884,N_2415);
and UO_22 (O_22,N_2664,N_2680);
or UO_23 (O_23,N_2807,N_2418);
or UO_24 (O_24,N_2391,N_2856);
nand UO_25 (O_25,N_2530,N_2925);
or UO_26 (O_26,N_2632,N_2329);
nor UO_27 (O_27,N_2361,N_2912);
nor UO_28 (O_28,N_2808,N_2516);
or UO_29 (O_29,N_2707,N_2904);
xor UO_30 (O_30,N_2345,N_2446);
and UO_31 (O_31,N_2283,N_2802);
or UO_32 (O_32,N_2622,N_2593);
nand UO_33 (O_33,N_2625,N_2943);
or UO_34 (O_34,N_2398,N_2701);
nand UO_35 (O_35,N_2852,N_2638);
and UO_36 (O_36,N_2545,N_2534);
nor UO_37 (O_37,N_2824,N_2510);
or UO_38 (O_38,N_2928,N_2365);
xnor UO_39 (O_39,N_2408,N_2983);
nor UO_40 (O_40,N_2333,N_2343);
nor UO_41 (O_41,N_2954,N_2655);
nor UO_42 (O_42,N_2863,N_2416);
and UO_43 (O_43,N_2988,N_2533);
xnor UO_44 (O_44,N_2695,N_2763);
or UO_45 (O_45,N_2535,N_2868);
or UO_46 (O_46,N_2476,N_2780);
nand UO_47 (O_47,N_2406,N_2266);
or UO_48 (O_48,N_2500,N_2359);
xor UO_49 (O_49,N_2287,N_2919);
nand UO_50 (O_50,N_2811,N_2909);
xnor UO_51 (O_51,N_2384,N_2606);
or UO_52 (O_52,N_2568,N_2468);
nand UO_53 (O_53,N_2923,N_2496);
or UO_54 (O_54,N_2796,N_2736);
and UO_55 (O_55,N_2537,N_2561);
nor UO_56 (O_56,N_2926,N_2719);
and UO_57 (O_57,N_2573,N_2387);
or UO_58 (O_58,N_2825,N_2827);
and UO_59 (O_59,N_2386,N_2536);
or UO_60 (O_60,N_2251,N_2956);
nand UO_61 (O_61,N_2716,N_2587);
nand UO_62 (O_62,N_2921,N_2422);
xnor UO_63 (O_63,N_2583,N_2752);
and UO_64 (O_64,N_2485,N_2371);
nor UO_65 (O_65,N_2840,N_2549);
or UO_66 (O_66,N_2502,N_2375);
and UO_67 (O_67,N_2299,N_2838);
nor UO_68 (O_68,N_2259,N_2854);
nand UO_69 (O_69,N_2797,N_2920);
and UO_70 (O_70,N_2651,N_2557);
or UO_71 (O_71,N_2309,N_2645);
and UO_72 (O_72,N_2311,N_2624);
nor UO_73 (O_73,N_2582,N_2750);
nor UO_74 (O_74,N_2396,N_2698);
xor UO_75 (O_75,N_2597,N_2334);
or UO_76 (O_76,N_2350,N_2964);
or UO_77 (O_77,N_2541,N_2263);
nand UO_78 (O_78,N_2279,N_2454);
or UO_79 (O_79,N_2323,N_2335);
nor UO_80 (O_80,N_2442,N_2347);
nor UO_81 (O_81,N_2623,N_2635);
and UO_82 (O_82,N_2370,N_2894);
xor UO_83 (O_83,N_2431,N_2615);
xor UO_84 (O_84,N_2977,N_2971);
xor UO_85 (O_85,N_2783,N_2314);
xor UO_86 (O_86,N_2574,N_2326);
and UO_87 (O_87,N_2972,N_2467);
and UO_88 (O_88,N_2548,N_2458);
and UO_89 (O_89,N_2969,N_2547);
and UO_90 (O_90,N_2281,N_2941);
and UO_91 (O_91,N_2506,N_2295);
or UO_92 (O_92,N_2958,N_2613);
and UO_93 (O_93,N_2887,N_2460);
nor UO_94 (O_94,N_2286,N_2804);
nand UO_95 (O_95,N_2434,N_2368);
nor UO_96 (O_96,N_2531,N_2945);
or UO_97 (O_97,N_2449,N_2924);
or UO_98 (O_98,N_2621,N_2626);
nor UO_99 (O_99,N_2839,N_2886);
nand UO_100 (O_100,N_2274,N_2951);
nand UO_101 (O_101,N_2936,N_2666);
xnor UO_102 (O_102,N_2566,N_2672);
nand UO_103 (O_103,N_2596,N_2284);
nand UO_104 (O_104,N_2772,N_2985);
xnor UO_105 (O_105,N_2417,N_2721);
and UO_106 (O_106,N_2993,N_2520);
nor UO_107 (O_107,N_2289,N_2429);
nor UO_108 (O_108,N_2602,N_2942);
xor UO_109 (O_109,N_2690,N_2499);
or UO_110 (O_110,N_2676,N_2405);
nand UO_111 (O_111,N_2300,N_2355);
and UO_112 (O_112,N_2841,N_2823);
and UO_113 (O_113,N_2726,N_2671);
nor UO_114 (O_114,N_2614,N_2801);
nor UO_115 (O_115,N_2660,N_2722);
nand UO_116 (O_116,N_2539,N_2362);
or UO_117 (O_117,N_2490,N_2509);
and UO_118 (O_118,N_2952,N_2911);
or UO_119 (O_119,N_2585,N_2619);
nand UO_120 (O_120,N_2296,N_2766);
and UO_121 (O_121,N_2525,N_2455);
nor UO_122 (O_122,N_2865,N_2790);
or UO_123 (O_123,N_2426,N_2641);
xor UO_124 (O_124,N_2661,N_2843);
nor UO_125 (O_125,N_2328,N_2949);
nand UO_126 (O_126,N_2570,N_2255);
and UO_127 (O_127,N_2795,N_2914);
and UO_128 (O_128,N_2553,N_2592);
or UO_129 (O_129,N_2663,N_2778);
nand UO_130 (O_130,N_2647,N_2744);
and UO_131 (O_131,N_2538,N_2702);
nand UO_132 (O_132,N_2770,N_2963);
xor UO_133 (O_133,N_2607,N_2654);
or UO_134 (O_134,N_2569,N_2742);
nor UO_135 (O_135,N_2421,N_2720);
or UO_136 (O_136,N_2901,N_2853);
or UO_137 (O_137,N_2906,N_2946);
and UO_138 (O_138,N_2617,N_2379);
nor UO_139 (O_139,N_2761,N_2493);
nor UO_140 (O_140,N_2918,N_2540);
nand UO_141 (O_141,N_2862,N_2610);
or UO_142 (O_142,N_2675,N_2732);
nand UO_143 (O_143,N_2965,N_2630);
nor UO_144 (O_144,N_2526,N_2315);
or UO_145 (O_145,N_2997,N_2771);
and UO_146 (O_146,N_2837,N_2341);
or UO_147 (O_147,N_2558,N_2544);
nand UO_148 (O_148,N_2354,N_2412);
or UO_149 (O_149,N_2799,N_2685);
xor UO_150 (O_150,N_2774,N_2492);
or UO_151 (O_151,N_2339,N_2659);
nand UO_152 (O_152,N_2301,N_2764);
xnor UO_153 (O_153,N_2452,N_2260);
or UO_154 (O_154,N_2723,N_2961);
nor UO_155 (O_155,N_2803,N_2447);
and UO_156 (O_156,N_2684,N_2294);
or UO_157 (O_157,N_2435,N_2929);
nand UO_158 (O_158,N_2995,N_2465);
and UO_159 (O_159,N_2340,N_2765);
xor UO_160 (O_160,N_2581,N_2401);
nand UO_161 (O_161,N_2745,N_2327);
or UO_162 (O_162,N_2267,N_2832);
or UO_163 (O_163,N_2905,N_2356);
nand UO_164 (O_164,N_2775,N_2688);
or UO_165 (O_165,N_2512,N_2992);
nand UO_166 (O_166,N_2879,N_2953);
or UO_167 (O_167,N_2846,N_2631);
or UO_168 (O_168,N_2528,N_2453);
or UO_169 (O_169,N_2353,N_2423);
and UO_170 (O_170,N_2419,N_2565);
and UO_171 (O_171,N_2609,N_2830);
nand UO_172 (O_172,N_2973,N_2519);
and UO_173 (O_173,N_2572,N_2470);
nor UO_174 (O_174,N_2855,N_2527);
nand UO_175 (O_175,N_2895,N_2649);
nor UO_176 (O_176,N_2336,N_2265);
xor UO_177 (O_177,N_2381,N_2709);
and UO_178 (O_178,N_2962,N_2658);
nor UO_179 (O_179,N_2792,N_2728);
xnor UO_180 (O_180,N_2346,N_2305);
and UO_181 (O_181,N_2567,N_2877);
xor UO_182 (O_182,N_2984,N_2910);
or UO_183 (O_183,N_2682,N_2575);
nor UO_184 (O_184,N_2922,N_2440);
nand UO_185 (O_185,N_2507,N_2829);
nand UO_186 (O_186,N_2819,N_2578);
nand UO_187 (O_187,N_2321,N_2989);
or UO_188 (O_188,N_2849,N_2648);
and UO_189 (O_189,N_2696,N_2411);
nand UO_190 (O_190,N_2437,N_2633);
and UO_191 (O_191,N_2693,N_2932);
nor UO_192 (O_192,N_2950,N_2428);
nand UO_193 (O_193,N_2897,N_2691);
and UO_194 (O_194,N_2616,N_2938);
nor UO_195 (O_195,N_2757,N_2970);
nor UO_196 (O_196,N_2306,N_2407);
nand UO_197 (O_197,N_2687,N_2640);
nor UO_198 (O_198,N_2944,N_2318);
xor UO_199 (O_199,N_2699,N_2834);
or UO_200 (O_200,N_2273,N_2337);
nor UO_201 (O_201,N_2292,N_2781);
and UO_202 (O_202,N_2466,N_2308);
or UO_203 (O_203,N_2382,N_2257);
and UO_204 (O_204,N_2629,N_2955);
and UO_205 (O_205,N_2317,N_2364);
nor UO_206 (O_206,N_2873,N_2822);
nand UO_207 (O_207,N_2798,N_2586);
and UO_208 (O_208,N_2933,N_2270);
nand UO_209 (O_209,N_2250,N_2665);
nand UO_210 (O_210,N_2599,N_2360);
nand UO_211 (O_211,N_2598,N_2793);
or UO_212 (O_212,N_2275,N_2399);
nand UO_213 (O_213,N_2828,N_2760);
nor UO_214 (O_214,N_2390,N_2471);
nor UO_215 (O_215,N_2312,N_2727);
or UO_216 (O_216,N_2982,N_2870);
and UO_217 (O_217,N_2473,N_2319);
and UO_218 (O_218,N_2258,N_2352);
nand UO_219 (O_219,N_2380,N_2650);
or UO_220 (O_220,N_2282,N_2515);
or UO_221 (O_221,N_2791,N_2373);
nor UO_222 (O_222,N_2987,N_2410);
nor UO_223 (O_223,N_2522,N_2703);
or UO_224 (O_224,N_2351,N_2809);
nand UO_225 (O_225,N_2730,N_2959);
nor UO_226 (O_226,N_2461,N_2821);
nand UO_227 (O_227,N_2505,N_2331);
and UO_228 (O_228,N_2253,N_2363);
and UO_229 (O_229,N_2681,N_2494);
xnor UO_230 (O_230,N_2511,N_2885);
nand UO_231 (O_231,N_2483,N_2860);
and UO_232 (O_232,N_2898,N_2372);
and UO_233 (O_233,N_2291,N_2302);
nor UO_234 (O_234,N_2636,N_2739);
nand UO_235 (O_235,N_2858,N_2589);
and UO_236 (O_236,N_2782,N_2268);
or UO_237 (O_237,N_2448,N_2402);
or UO_238 (O_238,N_2290,N_2298);
and UO_239 (O_239,N_2342,N_2403);
nand UO_240 (O_240,N_2710,N_2262);
xnor UO_241 (O_241,N_2563,N_2521);
and UO_242 (O_242,N_2420,N_2388);
nand UO_243 (O_243,N_2734,N_2395);
and UO_244 (O_244,N_2835,N_2786);
xnor UO_245 (O_245,N_2404,N_2677);
and UO_246 (O_246,N_2310,N_2325);
nor UO_247 (O_247,N_2469,N_2875);
nor UO_248 (O_248,N_2818,N_2715);
nand UO_249 (O_249,N_2344,N_2293);
nor UO_250 (O_250,N_2759,N_2900);
xor UO_251 (O_251,N_2551,N_2491);
and UO_252 (O_252,N_2889,N_2307);
nand UO_253 (O_253,N_2639,N_2367);
or UO_254 (O_254,N_2882,N_2608);
xnor UO_255 (O_255,N_2271,N_2785);
or UO_256 (O_256,N_2842,N_2472);
xor UO_257 (O_257,N_2773,N_2644);
or UO_258 (O_258,N_2717,N_2817);
xor UO_259 (O_259,N_2850,N_2836);
or UO_260 (O_260,N_2656,N_2612);
and UO_261 (O_261,N_2686,N_2432);
nand UO_262 (O_262,N_2503,N_2867);
nor UO_263 (O_263,N_2482,N_2980);
and UO_264 (O_264,N_2588,N_2501);
nor UO_265 (O_265,N_2504,N_2712);
or UO_266 (O_266,N_2595,N_2394);
nor UO_267 (O_267,N_2477,N_2800);
or UO_268 (O_268,N_2976,N_2729);
and UO_269 (O_269,N_2436,N_2591);
and UO_270 (O_270,N_2366,N_2646);
nor UO_271 (O_271,N_2564,N_2261);
xnor UO_272 (O_272,N_2451,N_2668);
or UO_273 (O_273,N_2847,N_2810);
nand UO_274 (O_274,N_2899,N_2277);
nor UO_275 (O_275,N_2313,N_2883);
and UO_276 (O_276,N_2474,N_2383);
nand UO_277 (O_277,N_2931,N_2741);
nor UO_278 (O_278,N_2749,N_2708);
nor UO_279 (O_279,N_2994,N_2815);
nand UO_280 (O_280,N_2939,N_2896);
or UO_281 (O_281,N_2445,N_2433);
nand UO_282 (O_282,N_2618,N_2576);
nand UO_283 (O_283,N_2532,N_2304);
or UO_284 (O_284,N_2320,N_2462);
or UO_285 (O_285,N_2488,N_2256);
or UO_286 (O_286,N_2733,N_2913);
nor UO_287 (O_287,N_2484,N_2459);
nor UO_288 (O_288,N_2288,N_2679);
or UO_289 (O_289,N_2444,N_2940);
and UO_290 (O_290,N_2322,N_2252);
and UO_291 (O_291,N_2713,N_2642);
or UO_292 (O_292,N_2479,N_2937);
nor UO_293 (O_293,N_2330,N_2278);
xor UO_294 (O_294,N_2667,N_2747);
or UO_295 (O_295,N_2683,N_2580);
nand UO_296 (O_296,N_2397,N_2814);
nand UO_297 (O_297,N_2820,N_2603);
xor UO_298 (O_298,N_2670,N_2857);
nand UO_299 (O_299,N_2643,N_2753);
and UO_300 (O_300,N_2864,N_2996);
or UO_301 (O_301,N_2816,N_2981);
and UO_302 (O_302,N_2376,N_2392);
xnor UO_303 (O_303,N_2915,N_2264);
nor UO_304 (O_304,N_2784,N_2439);
nand UO_305 (O_305,N_2787,N_2611);
or UO_306 (O_306,N_2812,N_2393);
nand UO_307 (O_307,N_2806,N_2604);
xor UO_308 (O_308,N_2513,N_2400);
nor UO_309 (O_309,N_2594,N_2562);
and UO_310 (O_310,N_2762,N_2859);
or UO_311 (O_311,N_2697,N_2826);
or UO_312 (O_312,N_2848,N_2552);
or UO_313 (O_313,N_2902,N_2349);
nand UO_314 (O_314,N_2450,N_2427);
nand UO_315 (O_315,N_2890,N_2743);
nor UO_316 (O_316,N_2878,N_2463);
and UO_317 (O_317,N_2754,N_2880);
nor UO_318 (O_318,N_2487,N_2700);
and UO_319 (O_319,N_2908,N_2481);
nor UO_320 (O_320,N_2748,N_2711);
and UO_321 (O_321,N_2556,N_2794);
and UO_322 (O_322,N_2498,N_2694);
nor UO_323 (O_323,N_2991,N_2657);
and UO_324 (O_324,N_2480,N_2424);
or UO_325 (O_325,N_2979,N_2872);
or UO_326 (O_326,N_2620,N_2524);
nor UO_327 (O_327,N_2269,N_2601);
nand UO_328 (O_328,N_2935,N_2332);
nor UO_329 (O_329,N_2948,N_2517);
nor UO_330 (O_330,N_2637,N_2590);
nand UO_331 (O_331,N_2605,N_2735);
and UO_332 (O_332,N_2738,N_2844);
or UO_333 (O_333,N_2669,N_2689);
nand UO_334 (O_334,N_2907,N_2600);
nand UO_335 (O_335,N_2866,N_2280);
nand UO_336 (O_336,N_2947,N_2724);
and UO_337 (O_337,N_2579,N_2776);
nand UO_338 (O_338,N_2861,N_2554);
nor UO_339 (O_339,N_2377,N_2740);
and UO_340 (O_340,N_2348,N_2706);
and UO_341 (O_341,N_2584,N_2303);
xnor UO_342 (O_342,N_2385,N_2475);
and UO_343 (O_343,N_2874,N_2881);
nor UO_344 (O_344,N_2653,N_2930);
and UO_345 (O_345,N_2998,N_2903);
nand UO_346 (O_346,N_2678,N_2546);
and UO_347 (O_347,N_2746,N_2767);
or UO_348 (O_348,N_2755,N_2986);
nand UO_349 (O_349,N_2692,N_2957);
and UO_350 (O_350,N_2571,N_2974);
nor UO_351 (O_351,N_2731,N_2518);
or UO_352 (O_352,N_2272,N_2550);
nor UO_353 (O_353,N_2725,N_2917);
nand UO_354 (O_354,N_2758,N_2369);
nand UO_355 (O_355,N_2674,N_2968);
nand UO_356 (O_356,N_2254,N_2508);
or UO_357 (O_357,N_2876,N_2999);
or UO_358 (O_358,N_2378,N_2966);
and UO_359 (O_359,N_2529,N_2869);
nand UO_360 (O_360,N_2813,N_2893);
and UO_361 (O_361,N_2495,N_2934);
nor UO_362 (O_362,N_2967,N_2478);
or UO_363 (O_363,N_2891,N_2357);
xnor UO_364 (O_364,N_2756,N_2559);
nand UO_365 (O_365,N_2769,N_2978);
nor UO_366 (O_366,N_2768,N_2443);
or UO_367 (O_367,N_2975,N_2543);
nor UO_368 (O_368,N_2892,N_2438);
or UO_369 (O_369,N_2389,N_2831);
nor UO_370 (O_370,N_2714,N_2486);
or UO_371 (O_371,N_2737,N_2960);
nand UO_372 (O_372,N_2845,N_2297);
nor UO_373 (O_373,N_2464,N_2851);
or UO_374 (O_374,N_2285,N_2777);
and UO_375 (O_375,N_2497,N_2498);
and UO_376 (O_376,N_2437,N_2641);
nor UO_377 (O_377,N_2969,N_2253);
nand UO_378 (O_378,N_2501,N_2962);
nor UO_379 (O_379,N_2976,N_2843);
nand UO_380 (O_380,N_2484,N_2898);
nand UO_381 (O_381,N_2626,N_2557);
or UO_382 (O_382,N_2281,N_2970);
or UO_383 (O_383,N_2649,N_2604);
nand UO_384 (O_384,N_2306,N_2821);
or UO_385 (O_385,N_2375,N_2955);
nand UO_386 (O_386,N_2865,N_2576);
or UO_387 (O_387,N_2831,N_2712);
nor UO_388 (O_388,N_2528,N_2524);
or UO_389 (O_389,N_2430,N_2426);
xnor UO_390 (O_390,N_2904,N_2368);
or UO_391 (O_391,N_2661,N_2625);
nor UO_392 (O_392,N_2564,N_2413);
or UO_393 (O_393,N_2909,N_2313);
and UO_394 (O_394,N_2711,N_2905);
nor UO_395 (O_395,N_2938,N_2403);
nor UO_396 (O_396,N_2401,N_2675);
nand UO_397 (O_397,N_2407,N_2816);
and UO_398 (O_398,N_2354,N_2440);
nand UO_399 (O_399,N_2858,N_2563);
nor UO_400 (O_400,N_2526,N_2979);
nand UO_401 (O_401,N_2853,N_2899);
and UO_402 (O_402,N_2806,N_2701);
and UO_403 (O_403,N_2573,N_2506);
and UO_404 (O_404,N_2921,N_2281);
xor UO_405 (O_405,N_2823,N_2814);
xnor UO_406 (O_406,N_2663,N_2544);
nand UO_407 (O_407,N_2472,N_2926);
nand UO_408 (O_408,N_2533,N_2962);
nand UO_409 (O_409,N_2977,N_2416);
and UO_410 (O_410,N_2776,N_2353);
and UO_411 (O_411,N_2849,N_2507);
or UO_412 (O_412,N_2684,N_2314);
or UO_413 (O_413,N_2634,N_2893);
nor UO_414 (O_414,N_2621,N_2985);
xor UO_415 (O_415,N_2495,N_2772);
or UO_416 (O_416,N_2366,N_2421);
and UO_417 (O_417,N_2682,N_2568);
nor UO_418 (O_418,N_2654,N_2339);
nor UO_419 (O_419,N_2314,N_2560);
or UO_420 (O_420,N_2356,N_2304);
nand UO_421 (O_421,N_2661,N_2955);
and UO_422 (O_422,N_2311,N_2627);
nor UO_423 (O_423,N_2262,N_2866);
and UO_424 (O_424,N_2791,N_2850);
nor UO_425 (O_425,N_2423,N_2994);
or UO_426 (O_426,N_2900,N_2607);
xnor UO_427 (O_427,N_2905,N_2825);
nor UO_428 (O_428,N_2711,N_2818);
or UO_429 (O_429,N_2905,N_2774);
nor UO_430 (O_430,N_2366,N_2349);
nor UO_431 (O_431,N_2920,N_2997);
or UO_432 (O_432,N_2453,N_2747);
or UO_433 (O_433,N_2957,N_2601);
nor UO_434 (O_434,N_2760,N_2282);
and UO_435 (O_435,N_2774,N_2716);
xnor UO_436 (O_436,N_2786,N_2985);
xnor UO_437 (O_437,N_2453,N_2825);
and UO_438 (O_438,N_2528,N_2478);
nor UO_439 (O_439,N_2647,N_2846);
nand UO_440 (O_440,N_2606,N_2911);
and UO_441 (O_441,N_2611,N_2753);
xor UO_442 (O_442,N_2345,N_2604);
nor UO_443 (O_443,N_2704,N_2782);
xor UO_444 (O_444,N_2596,N_2738);
and UO_445 (O_445,N_2643,N_2311);
nor UO_446 (O_446,N_2265,N_2691);
nor UO_447 (O_447,N_2613,N_2910);
or UO_448 (O_448,N_2274,N_2869);
and UO_449 (O_449,N_2456,N_2882);
or UO_450 (O_450,N_2398,N_2531);
nor UO_451 (O_451,N_2962,N_2817);
nand UO_452 (O_452,N_2786,N_2673);
nor UO_453 (O_453,N_2720,N_2812);
xnor UO_454 (O_454,N_2849,N_2537);
nand UO_455 (O_455,N_2730,N_2879);
xor UO_456 (O_456,N_2637,N_2680);
nand UO_457 (O_457,N_2778,N_2559);
and UO_458 (O_458,N_2612,N_2584);
nand UO_459 (O_459,N_2783,N_2624);
nor UO_460 (O_460,N_2833,N_2426);
nor UO_461 (O_461,N_2908,N_2425);
nand UO_462 (O_462,N_2499,N_2389);
or UO_463 (O_463,N_2747,N_2709);
or UO_464 (O_464,N_2885,N_2402);
nand UO_465 (O_465,N_2394,N_2588);
nor UO_466 (O_466,N_2987,N_2890);
or UO_467 (O_467,N_2559,N_2642);
or UO_468 (O_468,N_2759,N_2336);
nor UO_469 (O_469,N_2561,N_2456);
nor UO_470 (O_470,N_2567,N_2966);
xor UO_471 (O_471,N_2904,N_2353);
nor UO_472 (O_472,N_2283,N_2763);
xnor UO_473 (O_473,N_2343,N_2295);
and UO_474 (O_474,N_2618,N_2566);
nor UO_475 (O_475,N_2467,N_2984);
nand UO_476 (O_476,N_2413,N_2867);
and UO_477 (O_477,N_2261,N_2316);
nor UO_478 (O_478,N_2827,N_2716);
nand UO_479 (O_479,N_2382,N_2994);
and UO_480 (O_480,N_2806,N_2915);
or UO_481 (O_481,N_2418,N_2599);
and UO_482 (O_482,N_2995,N_2770);
nand UO_483 (O_483,N_2990,N_2622);
xor UO_484 (O_484,N_2377,N_2718);
or UO_485 (O_485,N_2397,N_2467);
or UO_486 (O_486,N_2843,N_2842);
nor UO_487 (O_487,N_2662,N_2905);
xnor UO_488 (O_488,N_2677,N_2767);
nand UO_489 (O_489,N_2432,N_2632);
xnor UO_490 (O_490,N_2630,N_2531);
or UO_491 (O_491,N_2690,N_2941);
and UO_492 (O_492,N_2414,N_2617);
or UO_493 (O_493,N_2719,N_2394);
xor UO_494 (O_494,N_2919,N_2976);
nor UO_495 (O_495,N_2605,N_2801);
nor UO_496 (O_496,N_2732,N_2761);
xnor UO_497 (O_497,N_2967,N_2437);
nand UO_498 (O_498,N_2873,N_2519);
and UO_499 (O_499,N_2850,N_2529);
endmodule