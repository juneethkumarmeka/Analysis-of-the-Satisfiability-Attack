module basic_2000_20000_2500_100_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1358,In_86);
or U1 (N_1,In_245,In_346);
and U2 (N_2,In_1630,In_1506);
and U3 (N_3,In_840,In_1297);
nand U4 (N_4,In_607,In_790);
or U5 (N_5,In_1375,In_110);
nand U6 (N_6,In_1330,In_890);
nor U7 (N_7,In_1899,In_1897);
xnor U8 (N_8,In_1214,In_829);
nand U9 (N_9,In_1977,In_658);
and U10 (N_10,In_311,In_217);
or U11 (N_11,In_1288,In_1107);
or U12 (N_12,In_165,In_33);
nand U13 (N_13,In_308,In_1846);
and U14 (N_14,In_1440,In_1929);
nand U15 (N_15,In_1124,In_998);
nand U16 (N_16,In_1989,In_1179);
xor U17 (N_17,In_1346,In_661);
or U18 (N_18,In_1064,In_1021);
and U19 (N_19,In_690,In_995);
nand U20 (N_20,In_147,In_940);
nand U21 (N_21,In_946,In_1725);
and U22 (N_22,In_1101,In_1232);
xor U23 (N_23,In_27,In_764);
nor U24 (N_24,In_836,In_935);
and U25 (N_25,In_618,In_934);
nor U26 (N_26,In_1295,In_51);
nor U27 (N_27,In_1813,In_1408);
xnor U28 (N_28,In_1642,In_1025);
nand U29 (N_29,In_140,In_803);
xnor U30 (N_30,In_1139,In_1456);
and U31 (N_31,In_653,In_208);
nor U32 (N_32,In_1721,In_1906);
nor U33 (N_33,In_593,In_1320);
nand U34 (N_34,In_1728,In_69);
nor U35 (N_35,In_1390,In_533);
nor U36 (N_36,In_1678,In_169);
xnor U37 (N_37,In_1606,In_1473);
nor U38 (N_38,In_539,In_1381);
or U39 (N_39,In_315,In_1837);
nor U40 (N_40,In_1955,In_977);
nor U41 (N_41,In_1959,In_131);
nor U42 (N_42,In_104,In_993);
and U43 (N_43,In_1791,In_1026);
nand U44 (N_44,In_302,In_1760);
and U45 (N_45,In_473,In_806);
nand U46 (N_46,In_19,In_1009);
and U47 (N_47,In_886,In_303);
and U48 (N_48,In_163,In_791);
and U49 (N_49,In_895,In_421);
xnor U50 (N_50,In_15,In_422);
xnor U51 (N_51,In_1947,In_952);
or U52 (N_52,In_1076,In_854);
and U53 (N_53,In_894,In_1963);
and U54 (N_54,In_1762,In_1414);
or U55 (N_55,In_943,In_1600);
nor U56 (N_56,In_601,In_1127);
and U57 (N_57,In_435,In_1255);
nor U58 (N_58,In_1044,In_1551);
and U59 (N_59,In_730,In_160);
or U60 (N_60,In_1635,In_1941);
and U61 (N_61,In_613,In_1409);
and U62 (N_62,In_556,In_1495);
xnor U63 (N_63,In_1294,In_387);
xnor U64 (N_64,In_915,In_476);
and U65 (N_65,In_974,In_1772);
xor U66 (N_66,In_1264,In_445);
nand U67 (N_67,In_340,In_324);
xor U68 (N_68,In_591,In_862);
nor U69 (N_69,In_198,In_1571);
xnor U70 (N_70,In_1450,In_1911);
nand U71 (N_71,In_1313,In_1786);
nor U72 (N_72,In_1849,In_1377);
nor U73 (N_73,In_1140,In_1596);
and U74 (N_74,In_1823,In_863);
nor U75 (N_75,In_1744,In_23);
and U76 (N_76,In_1084,In_10);
nand U77 (N_77,In_686,In_1158);
or U78 (N_78,In_382,In_24);
and U79 (N_79,In_639,In_454);
or U80 (N_80,In_1833,In_1287);
nand U81 (N_81,In_606,In_641);
and U82 (N_82,In_930,In_920);
nor U83 (N_83,In_1080,In_747);
nand U84 (N_84,In_1467,In_365);
or U85 (N_85,In_910,In_1558);
nor U86 (N_86,In_620,In_203);
nand U87 (N_87,In_158,In_156);
or U88 (N_88,In_1661,In_558);
or U89 (N_89,In_299,In_1144);
or U90 (N_90,In_631,In_972);
nor U91 (N_91,In_1610,In_710);
nor U92 (N_92,In_646,In_1844);
xor U93 (N_93,In_278,In_336);
and U94 (N_94,In_1822,In_1985);
nand U95 (N_95,In_1994,In_1563);
xor U96 (N_96,In_314,In_553);
nor U97 (N_97,In_922,In_638);
nor U98 (N_98,In_1307,In_580);
or U99 (N_99,In_162,In_1736);
xor U100 (N_100,In_680,In_616);
nor U101 (N_101,In_1676,In_1904);
nand U102 (N_102,In_583,In_1914);
xor U103 (N_103,In_1344,In_841);
xor U104 (N_104,In_1516,In_538);
and U105 (N_105,In_50,In_726);
and U106 (N_106,In_1509,In_979);
or U107 (N_107,In_1182,In_1188);
nor U108 (N_108,In_885,In_1260);
nand U109 (N_109,In_1479,In_413);
nor U110 (N_110,In_735,In_1494);
or U111 (N_111,In_967,In_545);
nor U112 (N_112,In_508,In_1712);
and U113 (N_113,In_360,In_1001);
nor U114 (N_114,In_526,In_490);
or U115 (N_115,In_17,In_92);
nor U116 (N_116,In_1618,In_236);
nor U117 (N_117,In_1037,In_701);
nor U118 (N_118,In_1011,In_677);
and U119 (N_119,In_1389,In_222);
xor U120 (N_120,In_1034,In_1089);
nor U121 (N_121,In_1131,In_1388);
nand U122 (N_122,In_91,In_745);
and U123 (N_123,In_1687,In_1866);
and U124 (N_124,In_1591,In_849);
nor U125 (N_125,In_213,In_1343);
or U126 (N_126,In_118,In_414);
or U127 (N_127,In_150,In_1159);
or U128 (N_128,In_1907,In_1428);
or U129 (N_129,In_858,In_740);
and U130 (N_130,In_1898,In_1226);
and U131 (N_131,In_1711,In_1134);
xor U132 (N_132,In_1922,In_1587);
nand U133 (N_133,In_1379,In_1054);
or U134 (N_134,In_1119,In_544);
xor U135 (N_135,In_507,In_497);
nand U136 (N_136,In_725,In_781);
or U137 (N_137,In_1246,In_1468);
or U138 (N_138,In_189,In_1231);
and U139 (N_139,In_1259,In_325);
nor U140 (N_140,In_1268,In_1302);
or U141 (N_141,In_808,In_1520);
nand U142 (N_142,In_479,In_471);
xor U143 (N_143,In_1718,In_1812);
xnor U144 (N_144,In_1719,In_1930);
and U145 (N_145,In_557,In_866);
xnor U146 (N_146,In_1632,In_997);
xnor U147 (N_147,In_1471,In_477);
and U148 (N_148,In_1197,In_855);
xor U149 (N_149,In_579,In_185);
and U150 (N_150,In_876,In_1);
xnor U151 (N_151,In_736,In_1239);
nand U152 (N_152,In_959,In_154);
xor U153 (N_153,In_1281,In_218);
xor U154 (N_154,In_941,In_295);
nand U155 (N_155,In_342,In_563);
and U156 (N_156,In_180,In_955);
or U157 (N_157,In_1589,In_1583);
nand U158 (N_158,In_1656,In_1171);
nand U159 (N_159,In_715,In_501);
xnor U160 (N_160,In_722,In_1802);
and U161 (N_161,In_1191,In_847);
nand U162 (N_162,In_1835,In_1794);
or U163 (N_163,In_1187,In_403);
or U164 (N_164,In_1938,In_333);
nand U165 (N_165,In_1174,In_1219);
and U166 (N_166,In_1086,In_491);
nor U167 (N_167,In_173,In_559);
xor U168 (N_168,In_456,In_1000);
and U169 (N_169,In_186,In_1910);
and U170 (N_170,In_817,In_892);
nand U171 (N_171,In_1433,In_1141);
or U172 (N_172,In_681,In_1106);
and U173 (N_173,In_1045,In_1057);
nand U174 (N_174,In_531,In_1636);
nand U175 (N_175,In_472,In_1517);
or U176 (N_176,In_1586,In_1236);
or U177 (N_177,In_448,In_9);
or U178 (N_178,In_564,In_1122);
xor U179 (N_179,In_835,In_289);
nor U180 (N_180,In_1138,In_505);
xnor U181 (N_181,In_64,In_684);
and U182 (N_182,In_767,In_1406);
and U183 (N_183,In_1043,In_447);
or U184 (N_184,In_351,In_1785);
nor U185 (N_185,In_1204,In_1085);
xnor U186 (N_186,In_624,In_1942);
xor U187 (N_187,In_1623,In_90);
nand U188 (N_188,In_1900,In_199);
and U189 (N_189,In_1499,In_1709);
nand U190 (N_190,In_54,In_1177);
nor U191 (N_191,In_306,In_947);
or U192 (N_192,In_1919,In_1758);
xor U193 (N_193,In_1189,In_376);
and U194 (N_194,In_980,In_1284);
and U195 (N_195,In_845,In_994);
and U196 (N_196,In_436,In_673);
nand U197 (N_197,In_515,In_1658);
or U198 (N_198,In_8,In_101);
or U199 (N_199,In_1990,In_1493);
or U200 (N_200,In_1901,N_71);
nor U201 (N_201,In_1402,In_1308);
or U202 (N_202,In_280,In_773);
and U203 (N_203,In_1427,In_400);
and U204 (N_204,In_1625,In_540);
and U205 (N_205,In_588,In_1407);
nor U206 (N_206,N_19,In_1372);
nand U207 (N_207,In_1361,In_1761);
nor U208 (N_208,In_38,In_685);
nor U209 (N_209,In_1706,In_1114);
and U210 (N_210,In_1505,N_94);
xor U211 (N_211,In_427,In_753);
nand U212 (N_212,In_159,In_1273);
xor U213 (N_213,In_1518,In_1053);
nand U214 (N_214,In_29,In_1422);
or U215 (N_215,In_1326,N_168);
nor U216 (N_216,In_1002,In_720);
nor U217 (N_217,In_1503,In_1796);
or U218 (N_218,In_590,In_1477);
and U219 (N_219,In_519,In_1199);
nor U220 (N_220,In_1240,In_1363);
and U221 (N_221,In_1838,In_39);
or U222 (N_222,In_1031,In_903);
nor U223 (N_223,In_1885,In_1827);
xnor U224 (N_224,In_431,In_1731);
xor U225 (N_225,In_269,In_493);
nand U226 (N_226,In_1175,In_465);
nor U227 (N_227,In_549,In_1155);
and U228 (N_228,In_951,In_450);
and U229 (N_229,In_528,In_1017);
or U230 (N_230,In_697,In_1385);
nor U231 (N_231,In_461,In_834);
nor U232 (N_232,In_734,In_1418);
xnor U233 (N_233,In_1865,In_1047);
nand U234 (N_234,In_1194,In_396);
nor U235 (N_235,N_130,In_1764);
nor U236 (N_236,In_1617,In_389);
nor U237 (N_237,In_41,In_1225);
nor U238 (N_238,In_296,In_35);
xor U239 (N_239,In_711,N_40);
and U240 (N_240,In_323,In_1576);
xnor U241 (N_241,In_1980,In_148);
or U242 (N_242,In_1429,In_81);
and U243 (N_243,In_717,In_1525);
nand U244 (N_244,In_819,In_356);
nor U245 (N_245,In_1527,In_1223);
xor U246 (N_246,In_879,In_309);
xor U247 (N_247,In_569,In_1546);
nand U248 (N_248,In_1829,In_1986);
or U249 (N_249,In_712,In_1071);
or U250 (N_250,N_86,N_153);
nor U251 (N_251,In_1847,In_455);
nor U252 (N_252,In_566,In_1027);
and U253 (N_253,In_1018,N_174);
or U254 (N_254,In_322,N_62);
and U255 (N_255,In_1894,In_1501);
and U256 (N_256,In_729,In_965);
or U257 (N_257,In_152,In_242);
and U258 (N_258,N_133,In_667);
or U259 (N_259,In_1956,N_163);
xor U260 (N_260,In_1354,In_107);
nand U261 (N_261,In_1347,In_1208);
nand U262 (N_262,In_1153,In_831);
and U263 (N_263,In_1335,In_687);
and U264 (N_264,In_870,N_132);
nor U265 (N_265,In_1277,In_1637);
xor U266 (N_266,In_1275,In_1150);
and U267 (N_267,In_1304,In_543);
and U268 (N_268,In_758,In_73);
nand U269 (N_269,In_509,In_1063);
nand U270 (N_270,N_53,N_21);
or U271 (N_271,In_184,In_728);
xnor U272 (N_272,In_1593,In_1650);
nor U273 (N_273,In_292,In_1133);
xnor U274 (N_274,N_1,N_106);
nand U275 (N_275,In_562,In_457);
or U276 (N_276,In_757,In_1857);
nand U277 (N_277,In_122,In_989);
nand U278 (N_278,In_688,In_1060);
nor U279 (N_279,In_766,In_142);
nor U280 (N_280,In_931,In_1909);
nor U281 (N_281,In_742,In_708);
and U282 (N_282,In_317,In_443);
nand U283 (N_283,In_1003,N_5);
nor U284 (N_284,In_1818,In_77);
and U285 (N_285,In_640,In_370);
nor U286 (N_286,In_1222,In_1881);
or U287 (N_287,In_1944,In_1769);
and U288 (N_288,In_584,In_11);
xor U289 (N_289,In_1006,In_1365);
or U290 (N_290,In_1807,In_1181);
and U291 (N_291,In_1452,In_626);
nand U292 (N_292,In_1918,In_644);
xnor U293 (N_293,In_338,In_1903);
and U294 (N_294,In_1373,In_1569);
or U295 (N_295,In_1781,In_1183);
xor U296 (N_296,N_102,In_304);
nand U297 (N_297,In_825,N_198);
and U298 (N_298,In_214,N_43);
xnor U299 (N_299,In_749,In_348);
or U300 (N_300,In_1982,In_671);
or U301 (N_301,In_1988,N_85);
and U302 (N_302,In_1668,N_88);
xnor U303 (N_303,In_1950,In_1537);
nor U304 (N_304,N_98,In_1359);
or U305 (N_305,In_1640,In_398);
nor U306 (N_306,In_1341,In_578);
or U307 (N_307,In_1476,In_762);
xor U308 (N_308,In_875,In_1714);
or U309 (N_309,In_1300,In_1701);
nor U310 (N_310,In_62,In_380);
or U311 (N_311,In_1775,In_1212);
and U312 (N_312,In_1698,In_797);
and U313 (N_313,In_694,In_359);
or U314 (N_314,In_43,In_1530);
xnor U315 (N_315,N_107,In_1108);
and U316 (N_316,In_210,In_1132);
or U317 (N_317,In_1931,In_530);
xor U318 (N_318,In_489,In_355);
and U319 (N_319,N_52,N_48);
xor U320 (N_320,In_1889,In_779);
and U321 (N_321,In_621,N_78);
xor U322 (N_322,N_135,In_369);
nand U323 (N_323,In_756,In_224);
nand U324 (N_324,In_78,In_1555);
or U325 (N_325,In_1624,N_118);
or U326 (N_326,In_138,In_1686);
xnor U327 (N_327,In_957,In_1371);
nand U328 (N_328,In_1608,In_1483);
xnor U329 (N_329,In_743,In_1038);
nand U330 (N_330,In_813,In_871);
and U331 (N_331,In_1464,In_1792);
or U332 (N_332,In_1562,In_5);
or U333 (N_333,In_884,N_89);
xor U334 (N_334,In_1351,In_239);
or U335 (N_335,In_1425,N_191);
nor U336 (N_336,In_1875,In_1755);
nor U337 (N_337,In_1474,In_964);
xor U338 (N_338,In_1532,N_172);
nand U339 (N_339,In_896,N_199);
or U340 (N_340,In_195,In_1748);
nand U341 (N_341,In_1660,In_985);
nand U342 (N_342,In_1804,In_469);
nor U343 (N_343,In_1960,In_1543);
or U344 (N_344,In_882,In_284);
xor U345 (N_345,In_880,In_171);
or U346 (N_346,N_15,In_1083);
nand U347 (N_347,In_1568,In_911);
and U348 (N_348,In_1766,In_6);
and U349 (N_349,In_512,N_195);
or U350 (N_350,In_281,In_1780);
nand U351 (N_351,N_141,In_452);
xor U352 (N_352,N_196,In_1392);
and U353 (N_353,In_551,In_263);
or U354 (N_354,In_1578,In_552);
or U355 (N_355,In_1949,In_776);
nor U356 (N_356,In_1074,In_785);
nand U357 (N_357,N_38,In_377);
and U358 (N_358,In_226,N_128);
xnor U359 (N_359,In_1717,In_230);
nand U360 (N_360,In_738,In_602);
xnor U361 (N_361,In_14,In_1357);
xnor U362 (N_362,N_54,In_1504);
nor U363 (N_363,N_184,N_57);
nor U364 (N_364,In_1536,N_123);
or U365 (N_365,In_554,In_268);
xor U366 (N_366,In_1258,In_912);
nand U367 (N_367,In_1752,In_570);
and U368 (N_368,In_1803,In_332);
and U369 (N_369,In_1957,In_1943);
nor U370 (N_370,In_1056,In_625);
nor U371 (N_371,N_105,In_1102);
xor U372 (N_372,In_1227,In_1852);
or U373 (N_373,In_1328,In_488);
nand U374 (N_374,In_1376,In_1249);
or U375 (N_375,In_378,In_1314);
nand U376 (N_376,In_1272,In_1020);
or U377 (N_377,In_1285,In_1380);
nor U378 (N_378,In_1306,In_1192);
and U379 (N_379,In_649,In_192);
nor U380 (N_380,In_804,In_1121);
or U381 (N_381,In_1475,In_1271);
nand U382 (N_382,In_859,N_33);
and U383 (N_383,In_164,In_264);
and U384 (N_384,N_187,In_1662);
xnor U385 (N_385,In_642,In_698);
nand U386 (N_386,In_968,In_1560);
nor U387 (N_387,In_670,In_132);
nor U388 (N_388,In_1008,In_251);
nor U389 (N_389,In_1173,In_1213);
nor U390 (N_390,In_1200,In_1767);
or U391 (N_391,N_145,In_99);
nor U392 (N_392,In_1247,In_1861);
xor U393 (N_393,In_739,In_1378);
nor U394 (N_394,In_1682,In_265);
or U395 (N_395,In_1633,In_1186);
or U396 (N_396,N_164,In_391);
or U397 (N_397,N_157,In_20);
xor U398 (N_398,In_683,N_192);
nor U399 (N_399,In_1828,In_1859);
xnor U400 (N_400,N_116,In_547);
or U401 (N_401,In_659,In_1577);
and U402 (N_402,In_761,In_1496);
nand U403 (N_403,In_1394,In_520);
nor U404 (N_404,In_233,In_1350);
nand U405 (N_405,N_285,In_1399);
and U406 (N_406,In_1393,In_320);
nor U407 (N_407,In_1729,In_1099);
xor U408 (N_408,In_460,In_1292);
and U409 (N_409,N_356,In_674);
xor U410 (N_410,N_49,In_1110);
or U411 (N_411,In_798,In_1515);
and U412 (N_412,In_828,In_318);
or U413 (N_413,In_1870,In_1436);
or U414 (N_414,In_966,N_272);
xnor U415 (N_415,In_1443,In_917);
and U416 (N_416,In_741,In_630);
xnor U417 (N_417,In_1411,In_206);
xor U418 (N_418,In_115,In_1492);
or U419 (N_419,In_286,In_1739);
nand U420 (N_420,In_668,N_287);
or U421 (N_421,In_787,In_1417);
nand U422 (N_422,In_1973,In_521);
and U423 (N_423,In_794,In_1848);
nand U424 (N_424,In_976,In_282);
xor U425 (N_425,N_255,In_1839);
or U426 (N_426,N_129,In_45);
and U427 (N_427,In_1644,In_120);
xnor U428 (N_428,N_311,In_243);
or U429 (N_429,N_306,In_1749);
xnor U430 (N_430,In_1740,N_304);
nor U431 (N_431,In_430,N_109);
and U432 (N_432,In_883,In_1075);
xnor U433 (N_433,In_1735,In_449);
or U434 (N_434,In_1896,In_1081);
and U435 (N_435,In_769,In_1565);
nand U436 (N_436,In_1799,N_253);
nor U437 (N_437,In_1311,In_648);
and U438 (N_438,In_793,N_335);
nand U439 (N_439,In_978,In_1773);
and U440 (N_440,In_58,N_16);
nor U441 (N_441,N_271,N_66);
xor U442 (N_442,N_370,In_235);
and U443 (N_443,In_1680,In_498);
or U444 (N_444,In_874,In_72);
xor U445 (N_445,In_1220,In_1010);
nand U446 (N_446,In_604,N_312);
nor U447 (N_447,In_774,N_250);
xnor U448 (N_448,In_316,In_1190);
or U449 (N_449,In_353,N_270);
nand U450 (N_450,In_1730,In_177);
nor U451 (N_451,In_1609,In_1603);
or U452 (N_452,In_215,In_1743);
and U453 (N_453,In_902,In_384);
nand U454 (N_454,N_140,N_32);
or U455 (N_455,In_1856,N_59);
and U456 (N_456,N_277,In_1090);
nand U457 (N_457,In_536,In_1825);
xor U458 (N_458,In_357,In_1882);
nand U459 (N_459,In_1125,N_210);
nand U460 (N_460,In_1531,In_1522);
nor U461 (N_461,In_1424,In_113);
or U462 (N_462,In_1757,In_1946);
or U463 (N_463,In_1235,In_439);
or U464 (N_464,In_522,N_146);
or U465 (N_465,N_228,In_628);
nor U466 (N_466,In_1871,N_342);
nor U467 (N_467,In_1607,In_1404);
nor U468 (N_468,In_1572,In_1510);
or U469 (N_469,In_386,In_1978);
and U470 (N_470,N_127,In_1035);
xnor U471 (N_471,In_1327,In_788);
and U472 (N_472,In_300,In_1832);
nor U473 (N_473,In_853,In_1103);
xor U474 (N_474,In_991,In_223);
nor U475 (N_475,In_1078,In_1670);
and U476 (N_476,In_1004,N_61);
xor U477 (N_477,In_617,N_267);
nand U478 (N_478,In_1178,In_1143);
and U479 (N_479,In_1854,In_1843);
or U480 (N_480,In_1550,In_79);
or U481 (N_481,In_466,In_1283);
and U482 (N_482,In_1933,In_900);
nand U483 (N_483,In_405,In_1545);
nand U484 (N_484,In_128,In_703);
or U485 (N_485,In_83,N_131);
and U486 (N_486,N_395,In_1912);
nor U487 (N_487,In_330,In_799);
nor U488 (N_488,In_248,In_1783);
nand U489 (N_489,In_394,In_714);
and U490 (N_490,N_39,In_692);
nor U491 (N_491,In_1401,N_266);
xor U492 (N_492,In_1750,In_938);
xor U493 (N_493,N_314,In_59);
xnor U494 (N_494,In_25,In_1584);
nand U495 (N_495,N_67,In_1917);
and U496 (N_496,In_963,In_1689);
and U497 (N_497,N_238,In_253);
xor U498 (N_498,In_1597,In_746);
xnor U499 (N_499,In_153,In_1163);
nand U500 (N_500,In_600,In_1325);
and U501 (N_501,In_1789,In_272);
nand U502 (N_502,N_317,In_1458);
and U503 (N_503,In_155,In_878);
nor U504 (N_504,N_331,In_1423);
and U505 (N_505,In_1629,In_1442);
nor U506 (N_506,In_635,In_502);
nand U507 (N_507,N_215,In_1999);
nor U508 (N_508,In_301,N_189);
nand U509 (N_509,N_47,N_261);
nor U510 (N_510,In_1831,In_220);
and U511 (N_511,In_662,N_41);
xor U512 (N_512,N_136,In_125);
nor U513 (N_513,In_1157,In_1318);
nor U514 (N_514,In_1156,In_1673);
or U515 (N_515,In_983,In_129);
nor U516 (N_516,In_1615,In_1397);
and U517 (N_517,In_1485,In_1290);
xnor U518 (N_518,In_1254,In_1855);
nor U519 (N_519,In_1396,N_97);
and U520 (N_520,N_366,In_1671);
or U521 (N_521,In_1552,In_197);
or U522 (N_522,N_364,In_948);
or U523 (N_523,In_75,In_221);
xnor U524 (N_524,In_546,In_1118);
xnor U525 (N_525,In_893,In_1966);
and U526 (N_526,N_9,In_307);
nor U527 (N_527,In_723,In_1449);
or U528 (N_528,N_328,In_1954);
xnor U529 (N_529,In_76,N_319);
and U530 (N_530,N_384,In_108);
and U531 (N_531,In_942,In_247);
or U532 (N_532,N_185,In_1599);
nor U533 (N_533,In_257,In_1659);
or U534 (N_534,N_180,N_382);
nor U535 (N_535,In_1228,In_1142);
and U536 (N_536,In_1455,In_1962);
or U537 (N_537,In_909,In_1095);
or U538 (N_538,In_1841,In_792);
or U539 (N_539,In_402,In_1274);
nor U540 (N_540,In_191,In_1908);
and U541 (N_541,In_468,In_1621);
xor U542 (N_542,In_704,N_288);
nand U543 (N_543,In_1322,In_1461);
and U544 (N_544,In_1146,In_1776);
or U545 (N_545,In_1309,In_106);
or U546 (N_546,In_1958,N_313);
nor U547 (N_547,In_1602,In_1256);
or U548 (N_548,In_754,In_971);
xor U549 (N_549,In_1788,In_926);
or U550 (N_550,In_1710,In_7);
xnor U551 (N_551,N_171,In_329);
or U552 (N_552,N_29,In_1867);
and U553 (N_553,In_605,N_231);
xnor U554 (N_554,In_707,In_1257);
xnor U555 (N_555,In_1457,In_61);
nand U556 (N_556,In_1312,In_1446);
nand U557 (N_557,In_470,In_1708);
or U558 (N_558,In_227,In_172);
xor U559 (N_559,In_312,N_18);
and U560 (N_560,N_92,In_1688);
nor U561 (N_561,In_428,N_346);
nand U562 (N_562,In_1170,In_1400);
nor U563 (N_563,In_2,In_1800);
or U564 (N_564,In_1195,In_1556);
nand U565 (N_565,In_1421,N_193);
and U566 (N_566,In_1250,In_1905);
or U567 (N_567,In_1123,In_897);
xnor U568 (N_568,N_302,In_945);
and U569 (N_569,In_833,In_144);
nor U570 (N_570,In_1595,In_1759);
nor U571 (N_571,In_1815,In_241);
nand U572 (N_572,In_82,In_1147);
xor U573 (N_573,In_867,In_367);
nand U574 (N_574,In_811,In_1104);
nor U575 (N_575,N_147,In_1713);
nand U576 (N_576,In_499,N_63);
nand U577 (N_577,In_1362,In_527);
and U578 (N_578,In_999,In_1939);
nor U579 (N_579,N_14,N_121);
xor U580 (N_580,N_308,N_173);
nor U581 (N_581,In_1310,In_13);
nor U582 (N_582,In_1419,In_1851);
and U583 (N_583,In_31,In_181);
nand U584 (N_584,In_187,In_973);
and U585 (N_585,In_1996,In_201);
and U586 (N_586,N_298,In_992);
nor U587 (N_587,In_541,In_293);
xor U588 (N_588,In_1111,In_55);
or U589 (N_589,In_283,In_1547);
xor U590 (N_590,In_582,In_1180);
xnor U591 (N_591,In_313,In_1432);
nand U592 (N_592,In_1211,In_581);
and U593 (N_593,In_778,In_1160);
xnor U594 (N_594,In_1117,In_225);
nor U595 (N_595,In_1333,In_1243);
or U596 (N_596,In_383,In_1810);
and U597 (N_597,In_1932,In_1533);
or U598 (N_598,In_111,In_373);
xnor U599 (N_599,In_908,In_1667);
and U600 (N_600,In_1066,N_523);
xnor U601 (N_601,In_1198,In_399);
nor U602 (N_602,In_1319,In_869);
or U603 (N_603,In_1620,N_451);
nor U604 (N_604,In_366,N_516);
and U605 (N_605,In_1681,N_264);
and U606 (N_606,N_353,In_525);
and U607 (N_607,N_8,In_1166);
nand U608 (N_608,In_202,N_183);
xnor U609 (N_609,In_901,In_1965);
nor U610 (N_610,In_877,N_511);
nor U611 (N_611,N_46,N_589);
nand U612 (N_612,N_422,In_1028);
xor U613 (N_613,In_1233,In_1924);
nor U614 (N_614,N_540,In_1926);
xnor U615 (N_615,N_229,In_30);
nor U616 (N_616,In_207,In_1185);
nor U617 (N_617,In_462,N_249);
nand U618 (N_618,N_352,In_1937);
or U619 (N_619,In_1573,In_1774);
and U620 (N_620,N_430,In_1073);
nand U621 (N_621,In_1466,In_1218);
and U622 (N_622,N_404,In_275);
nor U623 (N_623,In_262,In_1613);
nand U624 (N_624,N_158,N_112);
and U625 (N_625,In_1022,In_1270);
and U626 (N_626,N_20,In_364);
nand U627 (N_627,In_397,In_343);
or U628 (N_628,In_151,N_380);
nand U629 (N_629,N_561,In_1679);
and U630 (N_630,In_744,In_807);
and U631 (N_631,In_949,N_381);
or U632 (N_632,In_1094,In_274);
xor U633 (N_633,N_432,In_1113);
and U634 (N_634,N_398,In_702);
nor U635 (N_635,N_426,In_109);
or U636 (N_636,In_1567,In_1278);
nand U637 (N_637,N_201,In_1727);
xor U638 (N_638,In_37,In_1012);
and U639 (N_639,In_881,In_629);
and U640 (N_640,In_1451,N_592);
nor U641 (N_641,N_558,In_550);
nand U642 (N_642,In_1983,In_228);
nand U643 (N_643,In_1923,In_127);
and U644 (N_644,In_1176,In_1093);
nor U645 (N_645,In_1934,N_148);
and U646 (N_646,In_843,In_1165);
or U647 (N_647,In_487,In_1940);
nor U648 (N_648,N_110,In_1145);
nor U649 (N_649,In_112,In_962);
xor U650 (N_650,In_1777,N_60);
nand U651 (N_651,In_1674,N_418);
xnor U652 (N_652,In_1005,In_786);
nor U653 (N_653,In_1805,N_421);
nand U654 (N_654,In_1540,N_336);
or U655 (N_655,In_246,In_368);
nor U656 (N_656,In_627,N_491);
and U657 (N_657,In_529,N_125);
xor U658 (N_658,N_486,In_1070);
nand U659 (N_659,In_1077,N_456);
nor U660 (N_660,N_549,In_1353);
and U661 (N_661,N_521,In_1383);
nand U662 (N_662,N_76,In_857);
and U663 (N_663,In_103,In_1694);
nor U664 (N_664,N_474,In_211);
nor U665 (N_665,In_417,N_509);
and U666 (N_666,In_1203,N_417);
or U667 (N_667,In_928,In_285);
nor U668 (N_668,In_1486,In_1779);
or U669 (N_669,In_575,N_396);
or U670 (N_670,In_1765,N_472);
nand U671 (N_671,N_160,In_1069);
and U672 (N_672,In_1067,In_1747);
xor U673 (N_673,In_1611,In_1519);
nand U674 (N_674,In_1352,In_732);
nand U675 (N_675,In_1500,N_351);
nor U676 (N_676,In_157,In_665);
nand U677 (N_677,N_10,N_350);
nand U678 (N_678,In_655,In_1315);
and U679 (N_679,In_1570,In_1329);
xnor U680 (N_680,In_1763,In_433);
xnor U681 (N_681,In_705,In_1628);
and U682 (N_682,In_1991,In_1580);
nand U683 (N_683,N_246,N_532);
and U684 (N_684,In_319,N_150);
and U685 (N_685,In_1193,In_205);
or U686 (N_686,In_956,N_575);
and U687 (N_687,N_460,In_1685);
or U688 (N_688,In_1130,N_137);
nand U689 (N_689,In_810,N_468);
nor U690 (N_690,N_56,In_724);
nand U691 (N_691,In_846,In_1403);
xor U692 (N_692,N_194,In_1265);
xnor U693 (N_693,In_1888,In_496);
nand U694 (N_694,In_200,In_193);
nand U695 (N_695,In_1690,N_295);
nor U696 (N_696,In_699,In_1324);
nor U697 (N_697,N_262,In_234);
xor U698 (N_698,N_594,In_1478);
nor U699 (N_699,In_800,In_212);
nand U700 (N_700,N_392,N_347);
nand U701 (N_701,In_100,N_409);
or U702 (N_702,In_1715,In_68);
nor U703 (N_703,In_1059,N_386);
nand U704 (N_704,In_393,N_179);
or U705 (N_705,In_654,In_689);
nor U706 (N_706,In_258,In_1024);
xor U707 (N_707,In_1826,In_1023);
xnor U708 (N_708,N_119,N_282);
xnor U709 (N_709,N_383,N_591);
and U710 (N_710,In_1033,N_571);
xor U711 (N_711,In_350,In_1431);
xnor U712 (N_712,In_237,In_1454);
nor U713 (N_713,In_102,In_49);
nand U714 (N_714,In_1512,N_537);
nor U715 (N_715,In_982,In_117);
or U716 (N_716,In_1819,In_812);
or U717 (N_717,In_1554,In_1019);
and U718 (N_718,N_560,N_457);
and U719 (N_719,N_96,In_988);
xnor U720 (N_720,In_669,N_506);
nor U721 (N_721,In_1205,N_507);
nor U722 (N_722,N_235,In_595);
nor U723 (N_723,In_768,In_484);
or U724 (N_724,N_565,N_520);
or U725 (N_725,In_503,In_16);
or U726 (N_726,In_1669,In_1282);
or U727 (N_727,In_1162,In_252);
nor U728 (N_728,In_44,In_1705);
xor U729 (N_729,In_271,In_1091);
xor U730 (N_730,In_105,In_927);
xnor U731 (N_731,In_832,In_1581);
xnor U732 (N_732,N_212,In_255);
or U733 (N_733,In_149,N_385);
nand U734 (N_734,N_569,In_190);
nand U735 (N_735,In_1677,In_805);
xnor U736 (N_736,In_143,In_1697);
nand U737 (N_737,In_1834,In_1969);
and U738 (N_738,N_553,N_543);
and U739 (N_739,In_1797,In_1135);
nor U740 (N_740,N_80,In_1387);
xnor U741 (N_741,In_634,N_4);
nor U742 (N_742,N_497,In_1215);
nand U743 (N_743,In_1097,In_1538);
or U744 (N_744,N_379,In_254);
xor U745 (N_745,In_48,In_1601);
or U746 (N_746,N_226,N_538);
or U747 (N_747,In_1703,In_672);
or U748 (N_748,In_36,In_1751);
nand U749 (N_749,In_1754,In_410);
nand U750 (N_750,N_139,In_209);
or U751 (N_751,N_22,In_1920);
nand U752 (N_752,N_590,In_916);
nor U753 (N_753,In_572,In_1915);
nor U754 (N_754,In_1741,In_1210);
and U755 (N_755,In_987,In_94);
or U756 (N_756,In_1109,In_1230);
nand U757 (N_757,In_1790,N_36);
nor U758 (N_758,In_864,In_1087);
xnor U759 (N_759,N_586,N_577);
and U760 (N_760,N_263,In_1972);
or U761 (N_761,N_340,N_545);
or U762 (N_762,N_449,In_1869);
xor U763 (N_763,N_394,In_1887);
nor U764 (N_764,In_1331,In_1997);
nand U765 (N_765,In_84,In_71);
or U766 (N_766,In_1840,In_887);
or U767 (N_767,In_1202,In_1614);
or U768 (N_768,N_300,In_1663);
xnor U769 (N_769,N_429,In_1575);
nor U770 (N_770,In_1267,In_438);
xor U771 (N_771,N_256,In_1641);
and U772 (N_772,In_1465,In_1566);
nand U773 (N_773,In_1695,In_560);
xnor U774 (N_774,N_581,N_478);
and U775 (N_775,In_594,N_464);
xor U776 (N_776,In_182,N_232);
and U777 (N_777,In_589,N_550);
nand U778 (N_778,In_1605,In_1415);
xnor U779 (N_779,N_480,In_1391);
nand U780 (N_780,N_359,N_416);
or U781 (N_781,In_598,In_534);
or U782 (N_782,In_1814,In_1793);
nor U783 (N_783,In_760,In_70);
nor U784 (N_784,In_1987,N_223);
and U785 (N_785,N_224,In_1420);
nand U786 (N_786,N_548,In_249);
and U787 (N_787,In_905,N_439);
or U788 (N_788,N_260,In_119);
nor U789 (N_789,In_1726,In_411);
nand U790 (N_790,N_167,In_771);
nor U791 (N_791,In_341,In_1691);
nand U792 (N_792,N_170,In_1784);
and U793 (N_793,In_63,N_316);
and U794 (N_794,In_1746,In_250);
nor U795 (N_795,In_537,In_1348);
and U796 (N_796,In_816,In_657);
xor U797 (N_797,In_1405,N_269);
nand U798 (N_798,N_70,N_403);
nor U799 (N_799,In_1692,N_64);
nor U800 (N_800,N_764,In_1303);
or U801 (N_801,N_789,In_483);
nand U802 (N_802,N_257,In_1666);
or U803 (N_803,In_1514,In_1463);
or U804 (N_804,N_241,In_1638);
and U805 (N_805,In_375,N_108);
nor U806 (N_806,In_1342,In_1136);
nor U807 (N_807,In_1459,N_220);
xnor U808 (N_808,In_907,In_1808);
or U809 (N_809,N_390,In_1448);
and U810 (N_810,In_609,N_332);
or U811 (N_811,In_1345,In_385);
nand U812 (N_812,N_329,N_562);
xor U813 (N_813,In_969,In_97);
nor U814 (N_814,In_610,N_406);
and U815 (N_815,In_1092,In_1830);
or U816 (N_816,In_1877,N_126);
or U817 (N_817,N_496,N_159);
nor U818 (N_818,N_355,In_1370);
xnor U819 (N_819,In_660,N_309);
and U820 (N_820,N_17,In_524);
nand U821 (N_821,N_205,N_602);
xnor U822 (N_822,N_774,N_616);
and U823 (N_823,N_371,In_1672);
xor U824 (N_824,In_358,In_1862);
nand U825 (N_825,N_415,In_1161);
xor U826 (N_826,N_402,In_66);
nor U827 (N_827,N_682,N_761);
nor U828 (N_828,In_650,In_1116);
xnor U829 (N_829,N_685,In_85);
xnor U830 (N_830,In_1340,N_552);
nor U831 (N_831,N_554,N_149);
nor U832 (N_832,In_1732,N_481);
or U833 (N_833,N_613,In_232);
nor U834 (N_834,In_1564,In_1129);
nor U835 (N_835,N_671,In_1058);
and U836 (N_836,N_697,N_276);
xnor U837 (N_837,N_652,In_795);
or U838 (N_838,N_597,In_133);
nor U839 (N_839,In_1209,In_716);
and U840 (N_840,N_599,N_13);
xor U841 (N_841,In_1384,In_1262);
and U842 (N_842,In_441,In_56);
xnor U843 (N_843,N_709,N_547);
xor U844 (N_844,N_700,N_469);
xnor U845 (N_845,In_838,In_814);
nand U846 (N_846,In_924,In_1511);
and U847 (N_847,In_1652,N_624);
or U848 (N_848,In_1206,In_1716);
nand U849 (N_849,In_748,In_1439);
nor U850 (N_850,N_372,N_369);
nor U851 (N_851,In_1482,N_462);
nor U852 (N_852,N_563,N_413);
xnor U853 (N_853,N_445,In_651);
and U854 (N_854,N_93,In_801);
xnor U855 (N_855,In_1626,In_585);
nand U856 (N_856,In_1657,In_780);
nor U857 (N_857,N_791,In_229);
and U858 (N_858,In_830,In_1269);
nand U859 (N_859,N_544,N_693);
or U860 (N_860,In_40,N_588);
or U861 (N_861,N_206,In_852);
xnor U862 (N_862,In_1876,N_144);
nor U863 (N_863,In_424,N_176);
xnor U864 (N_864,N_604,N_598);
nand U865 (N_865,N_368,N_11);
xnor U866 (N_866,In_1544,In_1072);
or U867 (N_867,N_117,In_1253);
nor U868 (N_868,In_899,N_557);
nand U869 (N_869,In_865,N_120);
nor U870 (N_870,In_1040,N_407);
or U871 (N_871,In_1498,N_758);
or U872 (N_872,In_238,N_444);
nand U873 (N_873,N_733,N_211);
nand U874 (N_874,In_666,N_735);
or U875 (N_875,N_362,In_820);
and U876 (N_876,N_784,N_465);
or U877 (N_877,In_827,N_691);
nor U878 (N_878,In_1039,In_328);
nor U879 (N_879,N_473,N_412);
and U880 (N_880,In_577,N_679);
nand U881 (N_881,In_176,In_1487);
and U882 (N_882,In_1367,In_1820);
xor U883 (N_883,N_749,N_753);
and U884 (N_884,In_1594,N_684);
nand U885 (N_885,N_639,N_542);
and U886 (N_886,In_1878,N_217);
nand U887 (N_887,N_82,N_712);
or U888 (N_888,N_305,In_1782);
or U889 (N_889,N_441,In_1699);
or U890 (N_890,In_1707,In_1296);
and U891 (N_891,N_799,In_446);
nor U892 (N_892,In_1654,In_1874);
and U893 (N_893,In_759,In_467);
xnor U894 (N_894,N_593,In_244);
and U895 (N_895,N_87,N_408);
nor U896 (N_896,In_932,In_406);
or U897 (N_897,N_640,In_576);
or U898 (N_898,N_6,In_868);
and U899 (N_899,N_436,In_1237);
xor U900 (N_900,N_746,N_695);
nand U901 (N_901,N_650,N_719);
nand U902 (N_902,In_939,N_155);
and U903 (N_903,N_258,In_1971);
nor U904 (N_904,In_1864,In_1298);
xnor U905 (N_905,N_546,N_143);
xor U906 (N_906,N_254,In_510);
nand U907 (N_907,In_1369,In_1998);
and U908 (N_908,In_451,N_587);
and U909 (N_909,In_1007,In_464);
nor U910 (N_910,N_103,In_872);
xnor U911 (N_911,In_463,In_1497);
nand U912 (N_912,In_898,N_605);
or U913 (N_913,In_850,In_1460);
nand U914 (N_914,N_467,N_727);
nor U915 (N_915,In_22,In_1062);
and U916 (N_916,N_522,In_1032);
or U917 (N_917,N_579,In_121);
xnor U918 (N_918,In_1964,N_788);
nor U919 (N_919,N_202,N_517);
nor U920 (N_920,N_777,N_420);
or U921 (N_921,N_663,In_1491);
or U922 (N_922,N_459,In_240);
and U923 (N_923,In_1928,N_559);
xnor U924 (N_924,In_1148,N_233);
or U925 (N_925,N_572,N_752);
nor U926 (N_926,In_344,N_721);
or U927 (N_927,In_1883,N_625);
and U928 (N_928,In_231,In_481);
and U929 (N_929,In_713,N_675);
nand U930 (N_930,In_603,In_1088);
nor U931 (N_931,N_787,In_1700);
nor U932 (N_932,N_483,N_530);
xnor U933 (N_933,In_1280,N_237);
and U934 (N_934,In_1356,In_419);
or U935 (N_935,N_177,N_2);
nand U936 (N_936,N_162,N_601);
xnor U937 (N_937,N_7,N_297);
nor U938 (N_938,In_700,N_293);
nor U939 (N_939,In_954,In_475);
or U940 (N_940,N_248,N_512);
or U941 (N_941,In_1836,N_186);
xor U942 (N_942,In_1816,In_98);
xor U943 (N_943,In_1355,In_861);
nand U944 (N_944,In_440,N_503);
nor U945 (N_945,N_704,N_674);
and U946 (N_946,N_711,N_99);
xnor U947 (N_947,N_450,In_1016);
nor U948 (N_948,N_619,In_379);
nor U949 (N_949,N_500,In_194);
and U950 (N_950,N_515,In_1470);
or U951 (N_951,N_536,In_1806);
xnor U952 (N_952,In_371,N_534);
or U953 (N_953,In_52,N_609);
or U954 (N_954,N_477,N_216);
or U955 (N_955,In_936,N_595);
or U956 (N_956,N_633,In_1438);
nor U957 (N_957,In_1434,N_279);
nor U958 (N_958,N_337,N_169);
nor U959 (N_959,In_1588,N_730);
or U960 (N_960,N_771,In_1733);
or U961 (N_961,N_247,In_297);
and U962 (N_962,N_664,In_950);
or U963 (N_963,In_216,N_769);
nand U964 (N_964,N_573,In_442);
and U965 (N_965,In_1995,N_213);
and U966 (N_966,In_335,In_1238);
nand U967 (N_967,In_1042,In_480);
xor U968 (N_968,N_615,N_284);
or U969 (N_969,In_18,N_699);
nand U970 (N_970,N_45,N_626);
xor U971 (N_971,N_737,N_447);
nand U972 (N_972,N_794,N_236);
or U973 (N_973,In_1902,N_576);
xor U974 (N_974,N_708,In_3);
nor U975 (N_975,In_1722,In_587);
nor U976 (N_976,N_68,N_244);
and U977 (N_977,In_1734,N_683);
nor U978 (N_978,N_427,N_618);
or U979 (N_979,In_392,In_718);
nand U980 (N_980,In_1604,N_12);
nand U981 (N_981,In_719,In_1305);
and U982 (N_982,In_1234,In_134);
and U983 (N_983,In_919,In_1105);
nand U984 (N_984,N_606,In_1649);
and U985 (N_985,N_762,In_913);
xor U986 (N_986,N_175,N_101);
nand U987 (N_987,In_1374,In_511);
nor U988 (N_988,N_533,In_390);
and U989 (N_989,N_122,N_214);
nand U990 (N_990,N_376,N_360);
or U991 (N_991,In_733,In_1778);
nor U992 (N_992,In_1612,N_275);
and U993 (N_993,In_782,N_600);
and U994 (N_994,In_633,In_777);
and U995 (N_995,N_499,N_528);
or U996 (N_996,N_320,N_703);
nor U997 (N_997,In_1579,In_1100);
nand U998 (N_998,N_722,N_283);
xor U999 (N_999,In_1742,In_1893);
nor U1000 (N_1000,In_418,N_632);
or U1001 (N_1001,N_668,N_178);
xnor U1002 (N_1002,In_622,N_808);
nor U1003 (N_1003,In_273,N_330);
or U1004 (N_1004,N_800,N_608);
or U1005 (N_1005,N_658,N_959);
xor U1006 (N_1006,In_1513,In_770);
nand U1007 (N_1007,N_113,In_261);
nor U1008 (N_1008,N_960,In_1229);
nand U1009 (N_1009,N_286,In_664);
or U1010 (N_1010,In_426,N_919);
xnor U1011 (N_1011,N_996,N_713);
nor U1012 (N_1012,N_424,N_908);
or U1013 (N_1013,In_663,In_288);
and U1014 (N_1014,N_348,In_137);
nand U1015 (N_1015,N_823,In_259);
nand U1016 (N_1016,In_1872,N_798);
nand U1017 (N_1017,N_647,N_51);
nor U1018 (N_1018,In_395,In_1167);
nand U1019 (N_1019,N_903,In_1252);
xnor U1020 (N_1020,In_459,In_826);
and U1021 (N_1021,N_763,N_539);
nor U1022 (N_1022,N_811,N_221);
or U1023 (N_1023,N_373,N_829);
and U1024 (N_1024,N_966,In_474);
nor U1025 (N_1025,N_865,In_986);
and U1026 (N_1026,N_251,In_823);
and U1027 (N_1027,In_1619,In_1981);
and U1028 (N_1028,In_573,N_470);
xor U1029 (N_1029,N_803,N_914);
nand U1030 (N_1030,In_775,N_884);
or U1031 (N_1031,N_879,N_448);
xnor U1032 (N_1032,N_868,In_1079);
nor U1033 (N_1033,In_260,In_1745);
nand U1034 (N_1034,N_689,N_649);
nor U1035 (N_1035,In_458,N_74);
and U1036 (N_1036,In_1753,N_124);
nor U1037 (N_1037,In_1925,In_944);
and U1038 (N_1038,In_1154,In_1631);
and U1039 (N_1039,N_268,In_1951);
nor U1040 (N_1040,N_690,In_1128);
nand U1041 (N_1041,N_446,In_535);
or U1042 (N_1042,N_25,N_728);
and U1043 (N_1043,N_344,In_506);
nor U1044 (N_1044,N_785,N_861);
or U1045 (N_1045,In_842,N_898);
or U1046 (N_1046,N_956,N_743);
xnor U1047 (N_1047,N_992,In_1015);
or U1048 (N_1048,N_281,N_461);
or U1049 (N_1049,N_611,N_827);
or U1050 (N_1050,In_1337,In_1221);
xnor U1051 (N_1051,N_873,N_111);
or U1052 (N_1052,N_943,N_698);
or U1053 (N_1053,N_475,N_154);
or U1054 (N_1054,N_333,In_1366);
xor U1055 (N_1055,In_923,N_732);
xnor U1056 (N_1056,In_1065,In_555);
nor U1057 (N_1057,N_874,In_486);
and U1058 (N_1058,N_200,In_1051);
and U1059 (N_1059,N_965,N_463);
or U1060 (N_1060,N_886,In_1014);
or U1061 (N_1061,N_939,In_4);
and U1062 (N_1062,In_331,In_571);
nand U1063 (N_1063,N_654,N_391);
and U1064 (N_1064,N_717,In_1216);
xor U1065 (N_1065,In_46,N_906);
and U1066 (N_1066,In_596,In_1480);
nand U1067 (N_1067,In_478,N_259);
xor U1068 (N_1068,N_651,In_1041);
nor U1069 (N_1069,In_1890,N_678);
or U1070 (N_1070,In_1992,In_65);
or U1071 (N_1071,In_141,N_585);
xor U1072 (N_1072,In_818,N_744);
nor U1073 (N_1073,In_1655,In_1821);
or U1074 (N_1074,N_883,In_361);
or U1075 (N_1075,In_1447,N_455);
nor U1076 (N_1076,N_222,In_1364);
and U1077 (N_1077,In_1481,N_104);
nor U1078 (N_1078,N_648,N_58);
nor U1079 (N_1079,In_1643,N_555);
and U1080 (N_1080,N_818,In_1768);
and U1081 (N_1081,In_518,N_849);
or U1082 (N_1082,N_243,In_87);
and U1083 (N_1083,N_902,N_240);
xnor U1084 (N_1084,N_397,In_513);
nor U1085 (N_1085,In_1245,N_878);
nor U1086 (N_1086,N_28,N_638);
xor U1087 (N_1087,In_279,N_138);
and U1088 (N_1088,In_1653,N_947);
or U1089 (N_1089,N_388,N_414);
nor U1090 (N_1090,In_305,In_975);
or U1091 (N_1091,In_656,In_1845);
and U1092 (N_1092,N_855,In_696);
or U1093 (N_1093,In_1115,N_296);
xnor U1094 (N_1094,N_688,In_1720);
nand U1095 (N_1095,N_801,In_429);
xor U1096 (N_1096,N_705,In_136);
nand U1097 (N_1097,N_508,N_858);
and U1098 (N_1098,In_1046,N_950);
xor U1099 (N_1099,N_526,In_1323);
and U1100 (N_1100,In_615,N_326);
nor U1101 (N_1101,N_245,In_1557);
nand U1102 (N_1102,In_1413,In_93);
nand U1103 (N_1103,N_754,N_844);
or U1104 (N_1104,In_1913,In_67);
nand U1105 (N_1105,N_617,In_1534);
nor U1106 (N_1106,N_476,In_1970);
nand U1107 (N_1107,N_623,N_837);
or U1108 (N_1108,N_760,N_807);
nand U1109 (N_1109,In_388,N_814);
nand U1110 (N_1110,In_1338,N_510);
xor U1111 (N_1111,N_782,In_783);
or U1112 (N_1112,In_1850,N_864);
or U1113 (N_1113,N_780,N_853);
or U1114 (N_1114,In_960,N_954);
nand U1115 (N_1115,N_751,N_363);
and U1116 (N_1116,In_219,In_765);
nand U1117 (N_1117,N_979,In_1266);
nand U1118 (N_1118,N_920,N_318);
nor U1119 (N_1119,In_1916,N_389);
or U1120 (N_1120,N_114,N_568);
nor U1121 (N_1121,In_1030,N_928);
nand U1122 (N_1122,N_970,In_652);
xor U1123 (N_1123,In_420,N_826);
nor U1124 (N_1124,In_860,N_891);
xor U1125 (N_1125,In_1801,N_893);
or U1126 (N_1126,N_857,N_993);
nand U1127 (N_1127,N_790,N_871);
nand U1128 (N_1128,In_401,N_745);
nor U1129 (N_1129,In_412,N_911);
nand U1130 (N_1130,In_1445,In_196);
nor U1131 (N_1131,In_1858,N_620);
nand U1132 (N_1132,In_695,In_408);
nand U1133 (N_1133,N_151,N_303);
nand U1134 (N_1134,N_786,N_775);
or U1135 (N_1135,In_1541,N_915);
xnor U1136 (N_1136,N_834,In_482);
or U1137 (N_1137,In_1184,N_440);
xor U1138 (N_1138,In_851,N_912);
nand U1139 (N_1139,In_891,N_603);
nand U1140 (N_1140,In_958,In_592);
xnor U1141 (N_1141,In_1242,N_905);
nand U1142 (N_1142,N_929,In_751);
nand U1143 (N_1143,N_492,In_1539);
nand U1144 (N_1144,In_179,N_289);
and U1145 (N_1145,In_116,N_997);
nor U1146 (N_1146,In_492,N_378);
nor U1147 (N_1147,In_981,N_866);
and U1148 (N_1148,In_647,N_292);
or U1149 (N_1149,N_951,N_981);
xor U1150 (N_1150,N_636,N_341);
and U1151 (N_1151,N_846,In_1286);
and U1152 (N_1152,In_1201,N_845);
nor U1153 (N_1153,N_81,N_948);
nor U1154 (N_1154,N_957,In_574);
nor U1155 (N_1155,N_926,In_611);
or U1156 (N_1156,N_955,N_203);
or U1157 (N_1157,N_900,N_802);
xnor U1158 (N_1158,In_809,N_875);
nand U1159 (N_1159,In_1704,In_755);
and U1160 (N_1160,In_1149,N_838);
and U1161 (N_1161,In_374,In_12);
nand U1162 (N_1162,N_901,N_755);
or U1163 (N_1163,In_914,In_1948);
nand U1164 (N_1164,In_95,N_681);
and U1165 (N_1165,In_1895,N_338);
nor U1166 (N_1166,N_934,N_665);
or U1167 (N_1167,N_770,N_442);
nand U1168 (N_1168,In_1860,In_354);
and U1169 (N_1169,N_768,In_166);
and U1170 (N_1170,N_643,In_337);
nor U1171 (N_1171,In_1386,N_963);
and U1172 (N_1172,In_32,N_927);
or U1173 (N_1173,N_634,N_466);
nor U1174 (N_1174,In_1935,In_345);
and U1175 (N_1175,N_797,In_568);
nand U1176 (N_1176,N_922,In_1489);
xor U1177 (N_1177,In_1993,N_750);
or U1178 (N_1178,N_687,N_888);
nand U1179 (N_1179,N_998,In_404);
nor U1180 (N_1180,N_227,N_265);
and U1181 (N_1181,In_856,N_976);
and U1182 (N_1182,N_301,N_962);
xnor U1183 (N_1183,In_984,N_504);
xor U1184 (N_1184,N_635,In_1316);
nor U1185 (N_1185,In_532,N_584);
nor U1186 (N_1186,N_453,N_909);
and U1187 (N_1187,In_1968,In_267);
xnor U1188 (N_1188,N_280,N_673);
nand U1189 (N_1189,In_675,In_1811);
and U1190 (N_1190,N_583,In_1756);
nor U1191 (N_1191,N_847,N_612);
and U1192 (N_1192,N_531,In_1590);
nand U1193 (N_1193,In_352,In_1217);
or U1194 (N_1194,N_747,In_1412);
or U1195 (N_1195,N_930,N_374);
nand U1196 (N_1196,In_1952,In_1349);
xor U1197 (N_1197,N_984,N_686);
and U1198 (N_1198,In_1639,In_1975);
and U1199 (N_1199,In_1508,N_323);
xor U1200 (N_1200,N_859,In_1112);
nand U1201 (N_1201,N_1092,In_1724);
nand U1202 (N_1202,N_1070,In_124);
nand U1203 (N_1203,In_1842,N_824);
and U1204 (N_1204,In_565,N_830);
and U1205 (N_1205,N_165,N_1065);
nand U1206 (N_1206,N_1185,N_958);
and U1207 (N_1207,N_405,N_1090);
and U1208 (N_1208,N_1168,In_1961);
nand U1209 (N_1209,N_239,N_860);
or U1210 (N_1210,N_290,N_1162);
nor U1211 (N_1211,In_60,N_1071);
and U1212 (N_1212,N_765,In_1817);
or U1213 (N_1213,N_629,In_1120);
xnor U1214 (N_1214,In_918,N_501);
xor U1215 (N_1215,N_1196,N_1189);
xnor U1216 (N_1216,In_1207,In_276);
xnor U1217 (N_1217,In_423,In_953);
xor U1218 (N_1218,N_428,N_870);
and U1219 (N_1219,N_741,N_819);
nor U1220 (N_1220,N_156,In_1592);
or U1221 (N_1221,N_291,N_1088);
xnor U1222 (N_1222,N_899,N_513);
or U1223 (N_1223,N_614,In_839);
or U1224 (N_1224,N_1097,N_1055);
nand U1225 (N_1225,In_1395,N_739);
and U1226 (N_1226,N_1126,N_1042);
nor U1227 (N_1227,N_566,N_1130);
or U1228 (N_1228,N_1155,In_1574);
or U1229 (N_1229,N_622,N_435);
or U1230 (N_1230,N_1190,In_74);
nor U1231 (N_1231,N_1188,N_1001);
xnor U1232 (N_1232,In_1336,In_1824);
nor U1233 (N_1233,N_971,N_204);
or U1234 (N_1234,N_181,In_727);
xor U1235 (N_1235,N_969,In_636);
xnor U1236 (N_1236,N_1122,N_1083);
or U1237 (N_1237,In_1646,N_77);
or U1238 (N_1238,N_896,In_821);
and U1239 (N_1239,N_24,N_672);
or U1240 (N_1240,N_1067,In_57);
nor U1241 (N_1241,In_409,N_207);
xor U1242 (N_1242,N_925,N_645);
nor U1243 (N_1243,N_471,N_1016);
nand U1244 (N_1244,In_1279,N_1087);
or U1245 (N_1245,N_1095,In_1049);
nand U1246 (N_1246,N_835,In_1523);
xor U1247 (N_1247,In_523,N_1192);
or U1248 (N_1248,N_225,In_632);
or U1249 (N_1249,N_1187,N_1044);
nand U1250 (N_1250,N_423,In_1055);
nor U1251 (N_1251,In_763,In_1029);
or U1252 (N_1252,N_339,N_377);
xor U1253 (N_1253,In_1339,N_1150);
xnor U1254 (N_1254,In_434,N_1161);
nand U1255 (N_1255,N_27,N_1186);
and U1256 (N_1256,N_1159,N_1111);
and U1257 (N_1257,In_425,In_822);
and U1258 (N_1258,In_1261,N_100);
nand U1259 (N_1259,N_574,N_1170);
nand U1260 (N_1260,N_630,N_715);
xor U1261 (N_1261,N_1056,N_989);
and U1262 (N_1262,In_996,N_367);
nor U1263 (N_1263,In_339,N_1048);
or U1264 (N_1264,N_452,N_759);
nor U1265 (N_1265,N_458,N_1107);
and U1266 (N_1266,In_1927,In_327);
nand U1267 (N_1267,In_1665,N_766);
and U1268 (N_1268,N_278,N_964);
and U1269 (N_1269,In_1332,N_990);
nand U1270 (N_1270,N_724,N_399);
xnor U1271 (N_1271,N_987,In_28);
or U1272 (N_1272,In_437,N_694);
nor U1273 (N_1273,N_1081,In_291);
and U1274 (N_1274,N_1163,In_1936);
and U1275 (N_1275,In_1368,N_1195);
nor U1276 (N_1276,N_95,In_608);
xor U1277 (N_1277,In_737,N_387);
nand U1278 (N_1278,N_1074,N_637);
nand U1279 (N_1279,N_357,N_1180);
or U1280 (N_1280,N_852,N_748);
and U1281 (N_1281,N_518,N_1129);
nand U1282 (N_1282,N_1064,N_676);
and U1283 (N_1283,N_1157,In_266);
or U1284 (N_1284,N_1057,N_502);
xnor U1285 (N_1285,In_1437,N_1102);
and U1286 (N_1286,In_1559,N_1183);
xor U1287 (N_1287,N_1002,N_655);
xor U1288 (N_1288,N_209,N_646);
xnor U1289 (N_1289,N_941,N_1193);
nand U1290 (N_1290,In_1096,N_1005);
xor U1291 (N_1291,In_287,N_35);
xnor U1292 (N_1292,N_918,N_778);
xnor U1293 (N_1293,N_1032,N_299);
or U1294 (N_1294,In_334,In_145);
nor U1295 (N_1295,N_134,N_779);
xnor U1296 (N_1296,In_21,In_789);
nor U1297 (N_1297,In_645,In_561);
and U1298 (N_1298,N_494,N_69);
nand U1299 (N_1299,In_1126,N_1082);
and U1300 (N_1300,In_256,N_1121);
nor U1301 (N_1301,In_599,N_1103);
or U1302 (N_1302,In_990,N_1060);
and U1303 (N_1303,In_873,N_680);
nor U1304 (N_1304,In_679,N_1054);
and U1305 (N_1305,N_1007,N_968);
or U1306 (N_1306,In_1795,N_570);
nor U1307 (N_1307,N_1051,N_393);
and U1308 (N_1308,In_1648,In_1868);
xnor U1309 (N_1309,In_321,In_1528);
xnor U1310 (N_1310,In_1416,In_904);
nand U1311 (N_1311,In_1627,N_944);
nand U1312 (N_1312,N_1084,N_813);
nand U1313 (N_1313,N_1047,N_274);
nand U1314 (N_1314,N_524,N_1052);
or U1315 (N_1315,N_1026,N_988);
and U1316 (N_1316,N_1166,In_1472);
xor U1317 (N_1317,In_1891,N_1011);
nor U1318 (N_1318,N_991,In_444);
or U1319 (N_1319,In_889,N_188);
or U1320 (N_1320,N_1023,N_454);
nor U1321 (N_1321,N_832,In_42);
nand U1322 (N_1322,In_270,N_932);
nand U1323 (N_1323,N_894,N_438);
or U1324 (N_1324,N_1117,N_696);
xnor U1325 (N_1325,N_1176,In_721);
and U1326 (N_1326,N_1094,In_542);
nand U1327 (N_1327,In_1048,N_627);
or U1328 (N_1328,In_1549,N_843);
or U1329 (N_1329,In_139,N_657);
or U1330 (N_1330,N_707,In_678);
nor U1331 (N_1331,N_425,N_978);
or U1332 (N_1332,N_1105,N_667);
nand U1333 (N_1333,N_734,N_793);
nor U1334 (N_1334,N_1118,N_479);
xor U1335 (N_1335,N_1146,In_188);
or U1336 (N_1336,In_1524,N_809);
or U1337 (N_1337,N_653,N_1108);
nor U1338 (N_1338,N_815,In_1299);
nand U1339 (N_1339,N_1006,N_1080);
and U1340 (N_1340,N_692,N_938);
nand U1341 (N_1341,N_792,In_1622);
or U1342 (N_1342,In_1548,N_1139);
and U1343 (N_1343,N_720,N_541);
or U1344 (N_1344,In_123,N_1147);
xnor U1345 (N_1345,In_1974,N_1131);
nand U1346 (N_1346,In_1224,N_973);
nand U1347 (N_1347,N_1012,N_1091);
nand U1348 (N_1348,N_876,In_848);
nand U1349 (N_1349,N_400,N_1173);
and U1350 (N_1350,N_1149,N_949);
or U1351 (N_1351,In_504,N_1079);
xor U1352 (N_1352,N_897,In_1137);
nor U1353 (N_1353,N_580,N_1154);
nor U1354 (N_1354,N_723,N_1142);
and U1355 (N_1355,N_1182,N_726);
xnor U1356 (N_1356,N_931,In_1444);
or U1357 (N_1357,N_877,N_607);
and U1358 (N_1358,In_1169,N_490);
or U1359 (N_1359,In_1892,In_1723);
and U1360 (N_1360,N_659,N_889);
or U1361 (N_1361,N_1123,N_365);
nor U1362 (N_1362,In_204,In_1598);
and U1363 (N_1363,N_1061,N_1171);
nand U1364 (N_1364,N_1073,In_170);
nand U1365 (N_1365,In_691,N_701);
and U1366 (N_1366,In_1787,In_1068);
or U1367 (N_1367,N_1028,N_1015);
nand U1368 (N_1368,In_1098,N_882);
nor U1369 (N_1369,N_273,N_50);
nand U1370 (N_1370,N_325,N_890);
nand U1371 (N_1371,In_1241,In_407);
and U1372 (N_1372,N_1109,N_1013);
or U1373 (N_1373,In_1953,N_434);
xnor U1374 (N_1374,N_152,In_961);
nand U1375 (N_1375,N_1038,In_175);
and U1376 (N_1376,N_710,In_1263);
xor U1377 (N_1377,In_146,N_1020);
and U1378 (N_1378,N_869,N_885);
and U1379 (N_1379,In_1526,N_482);
or U1380 (N_1380,In_1984,N_840);
and U1381 (N_1381,N_851,N_961);
or U1382 (N_1382,N_1096,In_1036);
or U1383 (N_1383,N_315,N_1169);
nand U1384 (N_1384,N_1136,In_548);
xnor U1385 (N_1385,In_1426,In_1507);
xnor U1386 (N_1386,In_1469,N_872);
xnor U1387 (N_1387,In_0,N_493);
and U1388 (N_1388,N_529,In_34);
nand U1389 (N_1389,In_26,N_1033);
and U1390 (N_1390,N_995,In_1244);
nor U1391 (N_1391,N_334,In_1453);
or U1392 (N_1392,N_933,In_1647);
nand U1393 (N_1393,In_1886,In_135);
and U1394 (N_1394,N_1125,In_906);
nand U1395 (N_1395,N_661,N_756);
nand U1396 (N_1396,In_130,N_327);
or U1397 (N_1397,N_1089,N_806);
nand U1398 (N_1398,In_1921,N_73);
nand U1399 (N_1399,In_89,N_1116);
nor U1400 (N_1400,N_1115,N_1258);
and U1401 (N_1401,N_1148,N_1027);
and U1402 (N_1402,N_1304,In_614);
or U1403 (N_1403,N_1320,N_1383);
or U1404 (N_1404,In_752,In_1382);
xnor U1405 (N_1405,N_1198,N_1245);
nor U1406 (N_1406,N_1308,N_1210);
nand U1407 (N_1407,In_362,In_96);
nor U1408 (N_1408,N_83,N_1368);
and U1409 (N_1409,N_1272,N_945);
nand U1410 (N_1410,N_1324,N_773);
or U1411 (N_1411,N_1069,N_1128);
xor U1412 (N_1412,N_1252,N_642);
or U1413 (N_1413,N_1230,N_551);
or U1414 (N_1414,N_1254,N_1339);
nand U1415 (N_1415,N_1326,N_917);
and U1416 (N_1416,N_1200,In_676);
nand U1417 (N_1417,N_443,N_610);
nand U1418 (N_1418,N_974,In_183);
and U1419 (N_1419,In_1702,N_1341);
xnor U1420 (N_1420,N_1266,N_1325);
or U1421 (N_1421,In_1490,N_375);
nor U1422 (N_1422,N_489,N_1276);
nand U1423 (N_1423,N_527,N_1381);
and U1424 (N_1424,In_1675,N_1305);
and U1425 (N_1425,N_1158,N_1268);
or U1426 (N_1426,N_1376,N_1177);
and U1427 (N_1427,N_862,N_936);
nor U1428 (N_1428,In_1976,N_1025);
nand U1429 (N_1429,N_1068,N_1141);
and U1430 (N_1430,N_1045,In_1561);
nand U1431 (N_1431,N_1024,N_1086);
xor U1432 (N_1432,N_1172,N_1350);
nor U1433 (N_1433,N_84,N_1249);
xnor U1434 (N_1434,N_1374,N_1264);
or U1435 (N_1435,N_1019,N_488);
or U1436 (N_1436,N_812,N_1352);
nand U1437 (N_1437,N_1330,N_1004);
and U1438 (N_1438,N_1058,N_817);
nand U1439 (N_1439,In_495,In_114);
xor U1440 (N_1440,N_208,N_1314);
xor U1441 (N_1441,N_660,N_1263);
or U1442 (N_1442,N_1299,N_349);
xor U1443 (N_1443,N_1250,N_1093);
or U1444 (N_1444,N_952,N_1390);
xnor U1445 (N_1445,N_1357,N_1235);
nand U1446 (N_1446,In_168,N_1346);
nor U1447 (N_1447,N_182,In_294);
nand U1448 (N_1448,In_1863,N_1321);
or U1449 (N_1449,N_842,In_784);
nand U1450 (N_1450,In_750,N_1078);
nor U1451 (N_1451,In_643,N_1184);
nor U1452 (N_1452,N_776,N_1000);
and U1453 (N_1453,In_970,N_1290);
or U1454 (N_1454,In_517,In_1542);
nand U1455 (N_1455,N_1298,N_1377);
and U1456 (N_1456,N_535,In_921);
nor U1457 (N_1457,N_42,N_1137);
nand U1458 (N_1458,N_1132,N_1355);
and U1459 (N_1459,N_913,N_1336);
or U1460 (N_1460,N_358,In_167);
nand U1461 (N_1461,N_1380,N_1309);
or U1462 (N_1462,N_1285,N_1217);
or U1463 (N_1463,N_714,N_1291);
and U1464 (N_1464,N_1251,N_310);
and U1465 (N_1465,N_190,N_977);
nor U1466 (N_1466,N_1215,N_1396);
nand U1467 (N_1467,In_637,N_1269);
nand U1468 (N_1468,N_1367,N_161);
nor U1469 (N_1469,N_1144,N_564);
nand U1470 (N_1470,N_505,N_1009);
nor U1471 (N_1471,In_1276,N_578);
or U1472 (N_1472,In_290,N_1363);
xor U1473 (N_1473,N_1289,N_942);
and U1474 (N_1474,N_967,N_1369);
nor U1475 (N_1475,N_1119,N_1329);
xnor U1476 (N_1476,N_431,In_1441);
and U1477 (N_1477,N_1295,N_91);
xnor U1478 (N_1478,N_783,N_1322);
nor U1479 (N_1479,N_1342,N_1359);
nor U1480 (N_1480,N_904,N_1294);
nand U1481 (N_1481,N_1385,N_1348);
xor U1482 (N_1482,In_326,N_841);
nand U1483 (N_1483,N_1153,In_1967);
xnor U1484 (N_1484,In_1809,N_1394);
and U1485 (N_1485,N_1029,In_1050);
nand U1486 (N_1486,N_662,N_1283);
or U1487 (N_1487,N_37,In_80);
xor U1488 (N_1488,In_706,In_485);
xnor U1489 (N_1489,N_767,In_432);
and U1490 (N_1490,N_1260,N_115);
nand U1491 (N_1491,N_1391,In_53);
nand U1492 (N_1492,N_1328,N_1278);
and U1493 (N_1493,N_514,In_1521);
nor U1494 (N_1494,In_349,N_485);
xor U1495 (N_1495,N_1306,N_1035);
nor U1496 (N_1496,In_1634,N_1398);
and U1497 (N_1497,N_1041,N_1275);
and U1498 (N_1498,N_1372,In_1317);
or U1499 (N_1499,N_1114,N_1030);
or U1500 (N_1500,N_656,N_916);
nand U1501 (N_1501,N_411,N_1059);
or U1502 (N_1502,N_1053,N_1008);
nand U1503 (N_1503,N_1104,N_1244);
nand U1504 (N_1504,N_1282,N_935);
or U1505 (N_1505,In_174,N_1072);
nand U1506 (N_1506,N_731,N_1307);
nor U1507 (N_1507,N_1344,N_1099);
nand U1508 (N_1508,N_3,In_802);
nand U1509 (N_1509,N_1296,N_940);
and U1510 (N_1510,N_946,N_1207);
nor U1511 (N_1511,In_693,N_1243);
and U1512 (N_1512,In_1164,N_1127);
nand U1513 (N_1513,N_1362,N_1361);
and U1514 (N_1514,N_487,N_1262);
or U1515 (N_1515,N_321,N_1257);
nand U1516 (N_1516,N_1338,In_1684);
nand U1517 (N_1517,N_1286,N_498);
nand U1518 (N_1518,N_1206,N_831);
nand U1519 (N_1519,In_453,In_796);
and U1520 (N_1520,N_1145,In_567);
xnor U1521 (N_1521,N_242,N_1395);
nand U1522 (N_1522,In_347,N_666);
nor U1523 (N_1523,In_310,N_628);
and U1524 (N_1524,In_1301,N_1393);
xnor U1525 (N_1525,In_1884,N_1311);
and U1526 (N_1526,N_1036,N_556);
and U1527 (N_1527,N_166,N_1265);
xnor U1528 (N_1528,N_354,N_621);
xor U1529 (N_1529,N_1201,In_1398);
xnor U1530 (N_1530,N_796,N_26);
or U1531 (N_1531,N_1270,In_88);
nor U1532 (N_1532,N_1277,In_1585);
and U1533 (N_1533,In_1334,In_1738);
or U1534 (N_1534,N_1208,In_1289);
or U1535 (N_1535,N_1347,N_1333);
nor U1536 (N_1536,N_1046,N_1140);
nand U1537 (N_1537,N_795,N_1287);
xor U1538 (N_1538,N_1373,N_1101);
nor U1539 (N_1539,In_1535,In_1798);
xor U1540 (N_1540,N_1098,N_836);
xnor U1541 (N_1541,In_1616,N_1018);
nor U1542 (N_1542,N_1351,In_1291);
nand U1543 (N_1543,In_888,N_230);
and U1544 (N_1544,N_1040,In_1651);
or U1545 (N_1545,N_1358,N_1366);
nand U1546 (N_1546,N_1345,In_47);
and U1547 (N_1547,In_731,In_1462);
and U1548 (N_1548,N_1043,N_596);
xor U1549 (N_1549,In_1664,N_863);
and U1550 (N_1550,N_1310,N_839);
or U1551 (N_1551,N_1022,N_822);
and U1552 (N_1552,N_1194,In_619);
or U1553 (N_1553,N_1174,In_815);
or U1554 (N_1554,N_1151,N_1143);
nand U1555 (N_1555,In_298,N_825);
or U1556 (N_1556,N_345,In_1488);
and U1557 (N_1557,N_1343,N_982);
nand U1558 (N_1558,N_1219,N_410);
nor U1559 (N_1559,N_1317,In_1151);
or U1560 (N_1560,N_1222,N_1164);
nand U1561 (N_1561,In_1853,N_994);
nor U1562 (N_1562,N_1156,N_90);
or U1563 (N_1563,N_1247,N_892);
nor U1564 (N_1564,N_1216,In_1082);
and U1565 (N_1565,N_1349,In_1152);
and U1566 (N_1566,N_1334,N_31);
or U1567 (N_1567,N_781,N_401);
nand U1568 (N_1568,N_670,In_1693);
xor U1569 (N_1569,N_1273,N_75);
or U1570 (N_1570,N_1062,N_985);
nand U1571 (N_1571,N_142,In_516);
nand U1572 (N_1572,In_416,N_1316);
xnor U1573 (N_1573,N_816,In_1321);
nand U1574 (N_1574,N_820,N_234);
or U1575 (N_1575,N_1375,N_1234);
xor U1576 (N_1576,N_1167,N_525);
and U1577 (N_1577,N_1138,N_1292);
xor U1578 (N_1578,N_1233,N_1039);
or U1579 (N_1579,N_433,N_1165);
xnor U1580 (N_1580,N_1297,In_1435);
xnor U1581 (N_1581,In_161,N_1392);
or U1582 (N_1582,N_1152,N_923);
xor U1583 (N_1583,N_1077,In_1770);
nand U1584 (N_1584,N_1370,N_1232);
or U1585 (N_1585,N_1382,N_1100);
or U1586 (N_1586,In_1645,N_1255);
and U1587 (N_1587,N_1335,N_983);
or U1588 (N_1588,N_1204,N_1340);
xor U1589 (N_1589,N_1191,N_1010);
nor U1590 (N_1590,N_631,N_706);
nor U1591 (N_1591,N_924,N_23);
and U1592 (N_1592,N_218,N_1227);
xor U1593 (N_1593,In_1248,N_1327);
or U1594 (N_1594,N_1226,N_986);
nand U1595 (N_1595,N_1160,N_644);
xnor U1596 (N_1596,N_1246,N_343);
nand U1597 (N_1597,In_1251,N_1066);
nor U1598 (N_1598,N_716,In_372);
nor U1599 (N_1599,N_729,In_1771);
and U1600 (N_1600,N_1561,N_1438);
xnor U1601 (N_1601,N_1448,N_1534);
xnor U1602 (N_1602,N_1315,N_1420);
nor U1603 (N_1603,N_1259,N_810);
xor U1604 (N_1604,N_1211,N_219);
and U1605 (N_1605,N_1545,N_1505);
and U1606 (N_1606,N_1544,In_1502);
or U1607 (N_1607,N_1503,N_1223);
and U1608 (N_1608,In_929,In_1880);
or U1609 (N_1609,N_1037,In_597);
or U1610 (N_1610,N_1228,In_363);
nand U1611 (N_1611,N_1569,N_1549);
nor U1612 (N_1612,N_718,N_0);
xnor U1613 (N_1613,N_1496,N_1491);
nor U1614 (N_1614,In_1683,N_880);
or U1615 (N_1615,N_72,N_1591);
and U1616 (N_1616,In_178,N_34);
xnor U1617 (N_1617,N_1124,In_1052);
or U1618 (N_1618,N_1580,N_1267);
nor U1619 (N_1619,N_1540,N_1354);
xnor U1620 (N_1620,In_500,N_1432);
nor U1621 (N_1621,N_1423,N_1241);
and U1622 (N_1622,N_1487,N_1454);
and U1623 (N_1623,N_1318,N_1274);
or U1624 (N_1624,N_1364,N_1451);
nor U1625 (N_1625,N_1389,N_1181);
and U1626 (N_1626,In_1696,N_1465);
nor U1627 (N_1627,N_1431,N_322);
and U1628 (N_1628,N_1488,N_1134);
or U1629 (N_1629,N_1213,N_1525);
nor U1630 (N_1630,N_1527,N_1595);
and U1631 (N_1631,N_1224,N_1419);
nor U1632 (N_1632,N_1592,N_669);
and U1633 (N_1633,N_1236,N_1479);
and U1634 (N_1634,N_1478,N_1430);
and U1635 (N_1635,N_1501,N_1112);
nand U1636 (N_1636,N_1332,N_1494);
nand U1637 (N_1637,N_1412,N_1511);
or U1638 (N_1638,In_1061,N_1356);
and U1639 (N_1639,N_1353,In_824);
or U1640 (N_1640,N_1416,N_641);
or U1641 (N_1641,N_1429,N_1085);
xor U1642 (N_1642,N_1212,N_1179);
nor U1643 (N_1643,N_1466,N_1360);
xor U1644 (N_1644,In_1582,N_1453);
or U1645 (N_1645,N_1576,N_1439);
nor U1646 (N_1646,N_1288,N_1424);
or U1647 (N_1647,N_1445,N_1197);
and U1648 (N_1648,N_1464,N_1508);
xor U1649 (N_1649,N_1568,N_1458);
xor U1650 (N_1650,N_1567,N_1408);
xor U1651 (N_1651,N_1587,N_1021);
xor U1652 (N_1652,N_1063,N_1486);
xnor U1653 (N_1653,N_1583,N_1452);
nor U1654 (N_1654,N_1474,N_419);
and U1655 (N_1655,In_1410,N_1566);
nor U1656 (N_1656,N_1106,N_65);
nand U1657 (N_1657,N_740,N_937);
nor U1658 (N_1658,N_1548,N_1521);
nor U1659 (N_1659,N_1437,N_1386);
xnor U1660 (N_1660,N_1584,N_1578);
nand U1661 (N_1661,N_1536,N_1572);
nand U1662 (N_1662,N_1203,N_1242);
nor U1663 (N_1663,N_999,N_1441);
nand U1664 (N_1664,N_1303,N_1014);
nor U1665 (N_1665,N_1365,N_252);
xor U1666 (N_1666,N_1518,N_1443);
or U1667 (N_1667,N_1414,N_1279);
nor U1668 (N_1668,In_1293,N_828);
nor U1669 (N_1669,N_1240,N_582);
and U1670 (N_1670,N_1444,N_1399);
nor U1671 (N_1671,N_1564,N_757);
or U1672 (N_1672,N_821,N_1457);
xnor U1673 (N_1673,N_1574,N_1434);
and U1674 (N_1674,N_1471,N_55);
or U1675 (N_1675,N_1514,N_1220);
nand U1676 (N_1676,N_324,N_1462);
nand U1677 (N_1677,N_1426,N_1199);
or U1678 (N_1678,In_514,N_1323);
xnor U1679 (N_1679,N_1524,N_1594);
xor U1680 (N_1680,N_1522,N_1502);
nand U1681 (N_1681,N_856,N_1485);
nor U1682 (N_1682,In_612,In_1013);
or U1683 (N_1683,N_850,N_1588);
nor U1684 (N_1684,N_1379,N_1049);
nor U1685 (N_1685,In_925,N_307);
and U1686 (N_1686,N_1520,N_1415);
and U1687 (N_1687,N_1401,N_1472);
and U1688 (N_1688,N_1178,N_804);
or U1689 (N_1689,N_1550,N_975);
nor U1690 (N_1690,N_1559,N_736);
or U1691 (N_1691,In_1879,N_1532);
nand U1692 (N_1692,N_921,N_1535);
and U1693 (N_1693,N_1205,N_567);
nand U1694 (N_1694,N_1542,N_1593);
nor U1695 (N_1695,In_933,N_1442);
nand U1696 (N_1696,N_1475,N_1565);
and U1697 (N_1697,N_1516,N_1489);
xor U1698 (N_1698,N_1293,N_1400);
or U1699 (N_1699,N_1513,N_1214);
xnor U1700 (N_1700,N_1492,N_953);
nor U1701 (N_1701,In_844,N_1425);
and U1702 (N_1702,N_1468,In_1196);
nor U1703 (N_1703,N_1499,N_907);
and U1704 (N_1704,N_1579,N_1031);
or U1705 (N_1705,N_1538,In_1360);
xnor U1706 (N_1706,N_1530,N_1543);
and U1707 (N_1707,N_1417,N_1413);
nand U1708 (N_1708,N_772,N_895);
or U1709 (N_1709,N_1281,N_1337);
and U1710 (N_1710,N_1388,In_1979);
nand U1711 (N_1711,N_1509,N_1312);
and U1712 (N_1712,N_848,N_1371);
nor U1713 (N_1713,In_415,In_1172);
nor U1714 (N_1714,N_1421,N_1470);
and U1715 (N_1715,N_1581,N_30);
nor U1716 (N_1716,N_1135,N_1555);
or U1717 (N_1717,N_1557,N_1484);
xor U1718 (N_1718,N_738,N_1407);
xor U1719 (N_1719,N_1433,N_1599);
nor U1720 (N_1720,N_361,In_1553);
and U1721 (N_1721,N_1570,In_937);
and U1722 (N_1722,N_1387,N_980);
and U1723 (N_1723,N_1221,N_1428);
xor U1724 (N_1724,N_1110,In_837);
nor U1725 (N_1725,N_1422,In_277);
and U1726 (N_1726,N_1515,In_1945);
or U1727 (N_1727,N_854,N_1504);
and U1728 (N_1728,N_1510,N_1531);
and U1729 (N_1729,N_1483,In_586);
nor U1730 (N_1730,N_1003,N_1500);
nand U1731 (N_1731,N_1113,N_1397);
nor U1732 (N_1732,N_44,N_1229);
nand U1733 (N_1733,N_1410,In_772);
xnor U1734 (N_1734,N_1586,N_1467);
or U1735 (N_1735,N_495,N_1427);
xnor U1736 (N_1736,N_1517,N_1556);
nor U1737 (N_1737,N_1480,N_1378);
nor U1738 (N_1738,In_1430,N_805);
nand U1739 (N_1739,N_1571,N_1597);
and U1740 (N_1740,In_1484,N_1238);
or U1741 (N_1741,N_1523,N_1519);
nor U1742 (N_1742,N_1495,N_1017);
and U1743 (N_1743,N_1533,In_682);
or U1744 (N_1744,N_1120,N_1476);
nor U1745 (N_1745,N_1575,N_1237);
nor U1746 (N_1746,N_79,N_1418);
or U1747 (N_1747,N_1598,N_1034);
nor U1748 (N_1748,N_519,N_702);
and U1749 (N_1749,N_1302,N_1300);
or U1750 (N_1750,N_1446,N_1440);
nor U1751 (N_1751,N_1248,N_1526);
and U1752 (N_1752,N_677,N_1577);
nor U1753 (N_1753,N_1589,N_1582);
and U1754 (N_1754,In_1737,N_1551);
nand U1755 (N_1755,N_1498,N_1506);
nand U1756 (N_1756,N_1469,N_742);
or U1757 (N_1757,N_1497,N_1301);
xor U1758 (N_1758,N_1405,In_1168);
nor U1759 (N_1759,N_1133,N_1596);
nand U1760 (N_1760,N_1563,N_1404);
xor U1761 (N_1761,N_1490,In_623);
nand U1762 (N_1762,N_1481,N_725);
and U1763 (N_1763,N_1507,N_1539);
nand U1764 (N_1764,N_1075,N_1313);
nand U1765 (N_1765,N_1271,N_1406);
nand U1766 (N_1766,N_1456,N_294);
xnor U1767 (N_1767,N_1512,N_1225);
and U1768 (N_1768,N_1560,N_1553);
xor U1769 (N_1769,N_1482,N_1541);
or U1770 (N_1770,N_1461,N_484);
nor U1771 (N_1771,N_1590,N_1175);
nand U1772 (N_1772,N_1076,N_1554);
nor U1773 (N_1773,N_1256,N_1209);
or U1774 (N_1774,N_972,N_197);
nand U1775 (N_1775,N_437,In_1873);
nand U1776 (N_1776,N_1455,N_1537);
xor U1777 (N_1777,N_887,N_1546);
nand U1778 (N_1778,N_1261,N_1463);
and U1779 (N_1779,N_1409,N_1435);
nand U1780 (N_1780,N_1239,N_1447);
or U1781 (N_1781,N_1218,In_126);
or U1782 (N_1782,N_1477,N_1231);
nor U1783 (N_1783,In_381,N_1562);
nor U1784 (N_1784,N_1280,N_1253);
xnor U1785 (N_1785,N_1558,N_1411);
nor U1786 (N_1786,N_1529,N_1547);
and U1787 (N_1787,N_1384,N_1459);
nor U1788 (N_1788,N_1319,N_1493);
nor U1789 (N_1789,N_1050,N_1450);
and U1790 (N_1790,N_867,N_1402);
nor U1791 (N_1791,N_881,N_1552);
or U1792 (N_1792,N_1449,N_1585);
and U1793 (N_1793,N_910,In_709);
xor U1794 (N_1794,N_1202,In_1529);
nand U1795 (N_1795,N_1460,N_833);
and U1796 (N_1796,In_494,N_1473);
nor U1797 (N_1797,N_1284,N_1528);
xor U1798 (N_1798,N_1331,N_1436);
and U1799 (N_1799,N_1403,N_1573);
nand U1800 (N_1800,N_1643,N_1731);
nand U1801 (N_1801,N_1695,N_1628);
xor U1802 (N_1802,N_1799,N_1627);
and U1803 (N_1803,N_1642,N_1703);
and U1804 (N_1804,N_1654,N_1748);
or U1805 (N_1805,N_1659,N_1791);
and U1806 (N_1806,N_1644,N_1651);
or U1807 (N_1807,N_1749,N_1713);
nor U1808 (N_1808,N_1770,N_1754);
xnor U1809 (N_1809,N_1685,N_1697);
nor U1810 (N_1810,N_1601,N_1751);
xor U1811 (N_1811,N_1636,N_1797);
and U1812 (N_1812,N_1710,N_1687);
nor U1813 (N_1813,N_1728,N_1622);
xor U1814 (N_1814,N_1649,N_1777);
or U1815 (N_1815,N_1656,N_1702);
xor U1816 (N_1816,N_1773,N_1690);
and U1817 (N_1817,N_1670,N_1787);
and U1818 (N_1818,N_1609,N_1708);
nand U1819 (N_1819,N_1701,N_1733);
nand U1820 (N_1820,N_1620,N_1735);
nand U1821 (N_1821,N_1704,N_1646);
xor U1822 (N_1822,N_1789,N_1779);
nand U1823 (N_1823,N_1674,N_1657);
and U1824 (N_1824,N_1612,N_1738);
nand U1825 (N_1825,N_1758,N_1747);
or U1826 (N_1826,N_1744,N_1768);
xor U1827 (N_1827,N_1658,N_1798);
or U1828 (N_1828,N_1705,N_1729);
xor U1829 (N_1829,N_1741,N_1737);
nand U1830 (N_1830,N_1684,N_1720);
xor U1831 (N_1831,N_1630,N_1785);
or U1832 (N_1832,N_1756,N_1727);
and U1833 (N_1833,N_1689,N_1761);
or U1834 (N_1834,N_1638,N_1730);
nand U1835 (N_1835,N_1764,N_1717);
or U1836 (N_1836,N_1795,N_1641);
or U1837 (N_1837,N_1614,N_1712);
nor U1838 (N_1838,N_1631,N_1757);
nor U1839 (N_1839,N_1769,N_1693);
and U1840 (N_1840,N_1718,N_1726);
nand U1841 (N_1841,N_1615,N_1650);
nand U1842 (N_1842,N_1743,N_1663);
nor U1843 (N_1843,N_1602,N_1767);
nand U1844 (N_1844,N_1632,N_1714);
xnor U1845 (N_1845,N_1745,N_1673);
nand U1846 (N_1846,N_1784,N_1725);
nand U1847 (N_1847,N_1780,N_1700);
nor U1848 (N_1848,N_1774,N_1635);
or U1849 (N_1849,N_1623,N_1639);
and U1850 (N_1850,N_1652,N_1610);
or U1851 (N_1851,N_1640,N_1679);
and U1852 (N_1852,N_1665,N_1606);
or U1853 (N_1853,N_1607,N_1686);
or U1854 (N_1854,N_1788,N_1611);
or U1855 (N_1855,N_1624,N_1699);
xnor U1856 (N_1856,N_1711,N_1691);
nand U1857 (N_1857,N_1739,N_1740);
nand U1858 (N_1858,N_1671,N_1750);
and U1859 (N_1859,N_1715,N_1600);
and U1860 (N_1860,N_1736,N_1648);
nand U1861 (N_1861,N_1698,N_1696);
or U1862 (N_1862,N_1682,N_1629);
and U1863 (N_1863,N_1792,N_1677);
nand U1864 (N_1864,N_1608,N_1625);
or U1865 (N_1865,N_1668,N_1794);
or U1866 (N_1866,N_1746,N_1734);
nand U1867 (N_1867,N_1662,N_1653);
and U1868 (N_1868,N_1634,N_1755);
or U1869 (N_1869,N_1721,N_1752);
nand U1870 (N_1870,N_1680,N_1763);
or U1871 (N_1871,N_1722,N_1647);
and U1872 (N_1872,N_1616,N_1766);
and U1873 (N_1873,N_1753,N_1790);
and U1874 (N_1874,N_1655,N_1633);
or U1875 (N_1875,N_1683,N_1742);
or U1876 (N_1876,N_1765,N_1676);
nor U1877 (N_1877,N_1603,N_1664);
nand U1878 (N_1878,N_1666,N_1618);
or U1879 (N_1879,N_1776,N_1661);
xor U1880 (N_1880,N_1716,N_1724);
and U1881 (N_1881,N_1617,N_1783);
xnor U1882 (N_1882,N_1681,N_1771);
xor U1883 (N_1883,N_1759,N_1672);
and U1884 (N_1884,N_1719,N_1772);
nor U1885 (N_1885,N_1775,N_1723);
nor U1886 (N_1886,N_1688,N_1637);
or U1887 (N_1887,N_1707,N_1667);
nor U1888 (N_1888,N_1782,N_1692);
or U1889 (N_1889,N_1706,N_1732);
or U1890 (N_1890,N_1605,N_1619);
or U1891 (N_1891,N_1762,N_1709);
and U1892 (N_1892,N_1760,N_1781);
nand U1893 (N_1893,N_1621,N_1613);
nand U1894 (N_1894,N_1778,N_1660);
or U1895 (N_1895,N_1604,N_1796);
and U1896 (N_1896,N_1793,N_1678);
and U1897 (N_1897,N_1694,N_1675);
or U1898 (N_1898,N_1645,N_1786);
nor U1899 (N_1899,N_1669,N_1626);
or U1900 (N_1900,N_1637,N_1750);
xor U1901 (N_1901,N_1607,N_1617);
and U1902 (N_1902,N_1784,N_1664);
nand U1903 (N_1903,N_1603,N_1691);
nand U1904 (N_1904,N_1624,N_1658);
nor U1905 (N_1905,N_1692,N_1652);
xor U1906 (N_1906,N_1791,N_1792);
or U1907 (N_1907,N_1716,N_1635);
or U1908 (N_1908,N_1702,N_1641);
and U1909 (N_1909,N_1762,N_1711);
and U1910 (N_1910,N_1606,N_1732);
nor U1911 (N_1911,N_1676,N_1769);
xor U1912 (N_1912,N_1617,N_1635);
and U1913 (N_1913,N_1636,N_1704);
xnor U1914 (N_1914,N_1688,N_1716);
or U1915 (N_1915,N_1664,N_1732);
or U1916 (N_1916,N_1725,N_1711);
nor U1917 (N_1917,N_1693,N_1763);
nand U1918 (N_1918,N_1629,N_1637);
xnor U1919 (N_1919,N_1794,N_1631);
nand U1920 (N_1920,N_1798,N_1713);
nand U1921 (N_1921,N_1749,N_1623);
nor U1922 (N_1922,N_1650,N_1716);
nand U1923 (N_1923,N_1747,N_1746);
and U1924 (N_1924,N_1635,N_1770);
xor U1925 (N_1925,N_1600,N_1676);
or U1926 (N_1926,N_1647,N_1643);
xnor U1927 (N_1927,N_1753,N_1698);
xnor U1928 (N_1928,N_1720,N_1644);
xnor U1929 (N_1929,N_1748,N_1716);
nor U1930 (N_1930,N_1779,N_1621);
nand U1931 (N_1931,N_1709,N_1727);
and U1932 (N_1932,N_1736,N_1705);
nand U1933 (N_1933,N_1675,N_1605);
or U1934 (N_1934,N_1741,N_1743);
xor U1935 (N_1935,N_1699,N_1762);
nand U1936 (N_1936,N_1752,N_1731);
or U1937 (N_1937,N_1655,N_1607);
and U1938 (N_1938,N_1617,N_1672);
nor U1939 (N_1939,N_1700,N_1672);
and U1940 (N_1940,N_1643,N_1754);
and U1941 (N_1941,N_1712,N_1737);
or U1942 (N_1942,N_1665,N_1786);
nor U1943 (N_1943,N_1707,N_1620);
and U1944 (N_1944,N_1621,N_1608);
xor U1945 (N_1945,N_1728,N_1643);
xor U1946 (N_1946,N_1755,N_1750);
and U1947 (N_1947,N_1663,N_1609);
nand U1948 (N_1948,N_1613,N_1738);
nand U1949 (N_1949,N_1759,N_1698);
xnor U1950 (N_1950,N_1693,N_1721);
or U1951 (N_1951,N_1798,N_1760);
and U1952 (N_1952,N_1740,N_1681);
or U1953 (N_1953,N_1644,N_1755);
or U1954 (N_1954,N_1683,N_1719);
and U1955 (N_1955,N_1649,N_1721);
nor U1956 (N_1956,N_1748,N_1734);
nor U1957 (N_1957,N_1610,N_1798);
nand U1958 (N_1958,N_1627,N_1784);
or U1959 (N_1959,N_1726,N_1623);
and U1960 (N_1960,N_1733,N_1762);
xor U1961 (N_1961,N_1743,N_1779);
and U1962 (N_1962,N_1609,N_1745);
or U1963 (N_1963,N_1602,N_1645);
or U1964 (N_1964,N_1613,N_1620);
nor U1965 (N_1965,N_1656,N_1645);
or U1966 (N_1966,N_1693,N_1617);
or U1967 (N_1967,N_1624,N_1629);
nor U1968 (N_1968,N_1627,N_1636);
and U1969 (N_1969,N_1714,N_1728);
and U1970 (N_1970,N_1624,N_1651);
nand U1971 (N_1971,N_1724,N_1646);
and U1972 (N_1972,N_1755,N_1636);
nand U1973 (N_1973,N_1656,N_1676);
and U1974 (N_1974,N_1759,N_1775);
nor U1975 (N_1975,N_1715,N_1636);
nor U1976 (N_1976,N_1736,N_1645);
nor U1977 (N_1977,N_1704,N_1652);
or U1978 (N_1978,N_1789,N_1774);
xnor U1979 (N_1979,N_1638,N_1698);
nand U1980 (N_1980,N_1752,N_1643);
or U1981 (N_1981,N_1661,N_1658);
or U1982 (N_1982,N_1799,N_1645);
nand U1983 (N_1983,N_1747,N_1616);
or U1984 (N_1984,N_1787,N_1721);
nor U1985 (N_1985,N_1757,N_1736);
or U1986 (N_1986,N_1619,N_1664);
nand U1987 (N_1987,N_1753,N_1735);
and U1988 (N_1988,N_1630,N_1757);
nor U1989 (N_1989,N_1663,N_1729);
or U1990 (N_1990,N_1628,N_1765);
or U1991 (N_1991,N_1649,N_1740);
nand U1992 (N_1992,N_1762,N_1627);
nand U1993 (N_1993,N_1647,N_1672);
or U1994 (N_1994,N_1682,N_1701);
or U1995 (N_1995,N_1616,N_1686);
nand U1996 (N_1996,N_1759,N_1716);
xnor U1997 (N_1997,N_1645,N_1664);
or U1998 (N_1998,N_1625,N_1675);
xnor U1999 (N_1999,N_1730,N_1739);
or U2000 (N_2000,N_1909,N_1875);
nor U2001 (N_2001,N_1859,N_1926);
xor U2002 (N_2002,N_1980,N_1810);
nand U2003 (N_2003,N_1869,N_1800);
nand U2004 (N_2004,N_1802,N_1920);
nor U2005 (N_2005,N_1831,N_1836);
nand U2006 (N_2006,N_1937,N_1812);
nand U2007 (N_2007,N_1919,N_1960);
nor U2008 (N_2008,N_1917,N_1955);
nand U2009 (N_2009,N_1826,N_1941);
xnor U2010 (N_2010,N_1858,N_1945);
or U2011 (N_2011,N_1978,N_1856);
nor U2012 (N_2012,N_1981,N_1938);
or U2013 (N_2013,N_1877,N_1809);
nor U2014 (N_2014,N_1896,N_1923);
nand U2015 (N_2015,N_1889,N_1934);
nor U2016 (N_2016,N_1973,N_1846);
nor U2017 (N_2017,N_1946,N_1864);
nand U2018 (N_2018,N_1962,N_1924);
xor U2019 (N_2019,N_1882,N_1940);
nand U2020 (N_2020,N_1985,N_1997);
xor U2021 (N_2021,N_1983,N_1850);
nand U2022 (N_2022,N_1820,N_1825);
or U2023 (N_2023,N_1977,N_1839);
or U2024 (N_2024,N_1976,N_1930);
nor U2025 (N_2025,N_1815,N_1880);
and U2026 (N_2026,N_1990,N_1901);
nand U2027 (N_2027,N_1890,N_1971);
xor U2028 (N_2028,N_1958,N_1833);
or U2029 (N_2029,N_1979,N_1936);
or U2030 (N_2030,N_1984,N_1866);
xor U2031 (N_2031,N_1835,N_1855);
xnor U2032 (N_2032,N_1989,N_1892);
xnor U2033 (N_2033,N_1849,N_1986);
and U2034 (N_2034,N_1963,N_1821);
nand U2035 (N_2035,N_1834,N_1817);
and U2036 (N_2036,N_1908,N_1927);
xnor U2037 (N_2037,N_1957,N_1914);
xnor U2038 (N_2038,N_1886,N_1944);
and U2039 (N_2039,N_1847,N_1993);
or U2040 (N_2040,N_1942,N_1956);
and U2041 (N_2041,N_1883,N_1925);
nand U2042 (N_2042,N_1863,N_1972);
nor U2043 (N_2043,N_1933,N_1819);
and U2044 (N_2044,N_1871,N_1975);
and U2045 (N_2045,N_1885,N_1903);
and U2046 (N_2046,N_1922,N_1954);
xnor U2047 (N_2047,N_1952,N_1998);
or U2048 (N_2048,N_1822,N_1891);
xnor U2049 (N_2049,N_1921,N_1827);
and U2050 (N_2050,N_1854,N_1844);
nor U2051 (N_2051,N_1840,N_1974);
or U2052 (N_2052,N_1876,N_1801);
or U2053 (N_2053,N_1929,N_1910);
and U2054 (N_2054,N_1906,N_1965);
and U2055 (N_2055,N_1884,N_1939);
or U2056 (N_2056,N_1803,N_1982);
and U2057 (N_2057,N_1828,N_1904);
or U2058 (N_2058,N_1959,N_1931);
and U2059 (N_2059,N_1838,N_1870);
nand U2060 (N_2060,N_1900,N_1852);
or U2061 (N_2061,N_1879,N_1966);
nand U2062 (N_2062,N_1807,N_1824);
nor U2063 (N_2063,N_1907,N_1913);
nand U2064 (N_2064,N_1806,N_1848);
or U2065 (N_2065,N_1935,N_1893);
nor U2066 (N_2066,N_1823,N_1968);
nand U2067 (N_2067,N_1967,N_1949);
nor U2068 (N_2068,N_1898,N_1996);
nor U2069 (N_2069,N_1932,N_1878);
and U2070 (N_2070,N_1867,N_1873);
and U2071 (N_2071,N_1964,N_1961);
or U2072 (N_2072,N_1912,N_1808);
nand U2073 (N_2073,N_1947,N_1951);
or U2074 (N_2074,N_1902,N_1987);
and U2075 (N_2075,N_1804,N_1853);
nand U2076 (N_2076,N_1992,N_1948);
or U2077 (N_2077,N_1953,N_1999);
xor U2078 (N_2078,N_1829,N_1991);
nor U2079 (N_2079,N_1832,N_1816);
nand U2080 (N_2080,N_1857,N_1905);
or U2081 (N_2081,N_1813,N_1970);
nor U2082 (N_2082,N_1837,N_1895);
xor U2083 (N_2083,N_1814,N_1860);
xnor U2084 (N_2084,N_1899,N_1995);
and U2085 (N_2085,N_1868,N_1950);
and U2086 (N_2086,N_1862,N_1874);
xor U2087 (N_2087,N_1818,N_1916);
xnor U2088 (N_2088,N_1928,N_1830);
or U2089 (N_2089,N_1915,N_1894);
nor U2090 (N_2090,N_1881,N_1851);
nand U2091 (N_2091,N_1994,N_1805);
nor U2092 (N_2092,N_1897,N_1842);
xnor U2093 (N_2093,N_1843,N_1888);
and U2094 (N_2094,N_1845,N_1811);
and U2095 (N_2095,N_1872,N_1988);
or U2096 (N_2096,N_1943,N_1841);
nor U2097 (N_2097,N_1887,N_1911);
nor U2098 (N_2098,N_1865,N_1918);
nor U2099 (N_2099,N_1969,N_1861);
and U2100 (N_2100,N_1970,N_1919);
nand U2101 (N_2101,N_1949,N_1813);
nor U2102 (N_2102,N_1884,N_1904);
nand U2103 (N_2103,N_1864,N_1989);
and U2104 (N_2104,N_1849,N_1919);
and U2105 (N_2105,N_1938,N_1964);
nand U2106 (N_2106,N_1853,N_1945);
nand U2107 (N_2107,N_1852,N_1973);
nor U2108 (N_2108,N_1911,N_1932);
xor U2109 (N_2109,N_1959,N_1849);
xnor U2110 (N_2110,N_1854,N_1918);
nor U2111 (N_2111,N_1974,N_1828);
or U2112 (N_2112,N_1953,N_1908);
nand U2113 (N_2113,N_1812,N_1839);
or U2114 (N_2114,N_1873,N_1856);
and U2115 (N_2115,N_1971,N_1888);
nor U2116 (N_2116,N_1957,N_1977);
xor U2117 (N_2117,N_1842,N_1855);
nor U2118 (N_2118,N_1845,N_1918);
or U2119 (N_2119,N_1998,N_1935);
nand U2120 (N_2120,N_1871,N_1878);
and U2121 (N_2121,N_1919,N_1823);
or U2122 (N_2122,N_1919,N_1917);
nand U2123 (N_2123,N_1934,N_1888);
and U2124 (N_2124,N_1800,N_1901);
or U2125 (N_2125,N_1936,N_1984);
and U2126 (N_2126,N_1955,N_1965);
or U2127 (N_2127,N_1916,N_1950);
or U2128 (N_2128,N_1835,N_1824);
or U2129 (N_2129,N_1920,N_1927);
or U2130 (N_2130,N_1956,N_1814);
nor U2131 (N_2131,N_1975,N_1959);
nand U2132 (N_2132,N_1883,N_1820);
nor U2133 (N_2133,N_1876,N_1815);
xnor U2134 (N_2134,N_1895,N_1887);
or U2135 (N_2135,N_1962,N_1944);
nand U2136 (N_2136,N_1846,N_1877);
nand U2137 (N_2137,N_1879,N_1997);
nand U2138 (N_2138,N_1977,N_1813);
xnor U2139 (N_2139,N_1938,N_1844);
xnor U2140 (N_2140,N_1910,N_1912);
nand U2141 (N_2141,N_1928,N_1871);
nor U2142 (N_2142,N_1848,N_1976);
or U2143 (N_2143,N_1991,N_1834);
nand U2144 (N_2144,N_1988,N_1919);
nand U2145 (N_2145,N_1995,N_1953);
or U2146 (N_2146,N_1823,N_1994);
nor U2147 (N_2147,N_1853,N_1877);
xnor U2148 (N_2148,N_1867,N_1977);
nor U2149 (N_2149,N_1956,N_1828);
xor U2150 (N_2150,N_1836,N_1854);
xnor U2151 (N_2151,N_1912,N_1888);
nand U2152 (N_2152,N_1863,N_1989);
nand U2153 (N_2153,N_1916,N_1867);
and U2154 (N_2154,N_1882,N_1941);
nor U2155 (N_2155,N_1916,N_1932);
or U2156 (N_2156,N_1938,N_1806);
nand U2157 (N_2157,N_1885,N_1827);
and U2158 (N_2158,N_1817,N_1800);
nor U2159 (N_2159,N_1924,N_1827);
nand U2160 (N_2160,N_1985,N_1906);
and U2161 (N_2161,N_1941,N_1839);
xnor U2162 (N_2162,N_1970,N_1890);
nor U2163 (N_2163,N_1986,N_1818);
xnor U2164 (N_2164,N_1918,N_1908);
nand U2165 (N_2165,N_1977,N_1884);
nand U2166 (N_2166,N_1912,N_1992);
nor U2167 (N_2167,N_1869,N_1930);
xor U2168 (N_2168,N_1848,N_1961);
xor U2169 (N_2169,N_1878,N_1859);
and U2170 (N_2170,N_1907,N_1943);
nand U2171 (N_2171,N_1961,N_1916);
or U2172 (N_2172,N_1969,N_1927);
nor U2173 (N_2173,N_1817,N_1807);
and U2174 (N_2174,N_1950,N_1843);
or U2175 (N_2175,N_1803,N_1879);
and U2176 (N_2176,N_1996,N_1936);
nor U2177 (N_2177,N_1869,N_1913);
nand U2178 (N_2178,N_1854,N_1812);
xnor U2179 (N_2179,N_1891,N_1804);
xor U2180 (N_2180,N_1864,N_1919);
or U2181 (N_2181,N_1859,N_1925);
and U2182 (N_2182,N_1816,N_1847);
and U2183 (N_2183,N_1965,N_1966);
and U2184 (N_2184,N_1826,N_1912);
nand U2185 (N_2185,N_1995,N_1965);
nand U2186 (N_2186,N_1993,N_1926);
xor U2187 (N_2187,N_1847,N_1959);
nand U2188 (N_2188,N_1902,N_1993);
and U2189 (N_2189,N_1882,N_1966);
xor U2190 (N_2190,N_1885,N_1969);
xnor U2191 (N_2191,N_1919,N_1996);
nor U2192 (N_2192,N_1899,N_1927);
and U2193 (N_2193,N_1951,N_1939);
and U2194 (N_2194,N_1851,N_1898);
nor U2195 (N_2195,N_1940,N_1961);
xor U2196 (N_2196,N_1880,N_1924);
nand U2197 (N_2197,N_1842,N_1827);
or U2198 (N_2198,N_1834,N_1826);
and U2199 (N_2199,N_1882,N_1977);
nand U2200 (N_2200,N_2158,N_2121);
and U2201 (N_2201,N_2083,N_2153);
nor U2202 (N_2202,N_2003,N_2031);
xnor U2203 (N_2203,N_2102,N_2006);
or U2204 (N_2204,N_2014,N_2117);
nand U2205 (N_2205,N_2135,N_2103);
or U2206 (N_2206,N_2110,N_2059);
nor U2207 (N_2207,N_2020,N_2148);
nor U2208 (N_2208,N_2111,N_2071);
nand U2209 (N_2209,N_2193,N_2104);
and U2210 (N_2210,N_2189,N_2073);
and U2211 (N_2211,N_2173,N_2064);
nand U2212 (N_2212,N_2051,N_2079);
xnor U2213 (N_2213,N_2048,N_2122);
nand U2214 (N_2214,N_2015,N_2030);
and U2215 (N_2215,N_2176,N_2047);
or U2216 (N_2216,N_2082,N_2085);
xnor U2217 (N_2217,N_2062,N_2128);
nor U2218 (N_2218,N_2115,N_2130);
and U2219 (N_2219,N_2178,N_2197);
nor U2220 (N_2220,N_2098,N_2044);
xnor U2221 (N_2221,N_2192,N_2074);
or U2222 (N_2222,N_2040,N_2077);
xor U2223 (N_2223,N_2187,N_2140);
nor U2224 (N_2224,N_2177,N_2039);
xor U2225 (N_2225,N_2155,N_2114);
xnor U2226 (N_2226,N_2163,N_2068);
nor U2227 (N_2227,N_2133,N_2021);
nand U2228 (N_2228,N_2033,N_2028);
or U2229 (N_2229,N_2183,N_2069);
nor U2230 (N_2230,N_2007,N_2019);
and U2231 (N_2231,N_2011,N_2113);
or U2232 (N_2232,N_2129,N_2185);
nand U2233 (N_2233,N_2032,N_2066);
nor U2234 (N_2234,N_2164,N_2027);
xnor U2235 (N_2235,N_2149,N_2131);
nor U2236 (N_2236,N_2005,N_2095);
or U2237 (N_2237,N_2023,N_2038);
xor U2238 (N_2238,N_2001,N_2154);
and U2239 (N_2239,N_2167,N_2170);
nor U2240 (N_2240,N_2088,N_2137);
xor U2241 (N_2241,N_2058,N_2134);
nor U2242 (N_2242,N_2159,N_2078);
nor U2243 (N_2243,N_2054,N_2081);
nand U2244 (N_2244,N_2060,N_2161);
or U2245 (N_2245,N_2004,N_2136);
nand U2246 (N_2246,N_2087,N_2141);
or U2247 (N_2247,N_2182,N_2156);
nand U2248 (N_2248,N_2127,N_2125);
and U2249 (N_2249,N_2094,N_2181);
nor U2250 (N_2250,N_2000,N_2165);
and U2251 (N_2251,N_2029,N_2057);
nor U2252 (N_2252,N_2090,N_2037);
xor U2253 (N_2253,N_2056,N_2179);
nand U2254 (N_2254,N_2067,N_2180);
nand U2255 (N_2255,N_2018,N_2184);
nor U2256 (N_2256,N_2106,N_2147);
nor U2257 (N_2257,N_2138,N_2045);
or U2258 (N_2258,N_2084,N_2145);
nor U2259 (N_2259,N_2035,N_2061);
nor U2260 (N_2260,N_2120,N_2162);
xor U2261 (N_2261,N_2052,N_2016);
nor U2262 (N_2262,N_2008,N_2175);
xnor U2263 (N_2263,N_2191,N_2118);
or U2264 (N_2264,N_2144,N_2072);
and U2265 (N_2265,N_2126,N_2050);
xnor U2266 (N_2266,N_2026,N_2076);
nand U2267 (N_2267,N_2013,N_2142);
nor U2268 (N_2268,N_2091,N_2157);
or U2269 (N_2269,N_2150,N_2107);
or U2270 (N_2270,N_2063,N_2041);
nor U2271 (N_2271,N_2196,N_2009);
and U2272 (N_2272,N_2188,N_2168);
and U2273 (N_2273,N_2124,N_2100);
nor U2274 (N_2274,N_2199,N_2112);
and U2275 (N_2275,N_2024,N_2171);
nor U2276 (N_2276,N_2092,N_2099);
nor U2277 (N_2277,N_2043,N_2132);
nand U2278 (N_2278,N_2116,N_2146);
and U2279 (N_2279,N_2096,N_2055);
nor U2280 (N_2280,N_2123,N_2151);
xnor U2281 (N_2281,N_2194,N_2101);
xnor U2282 (N_2282,N_2139,N_2097);
or U2283 (N_2283,N_2010,N_2172);
xor U2284 (N_2284,N_2049,N_2070);
or U2285 (N_2285,N_2169,N_2034);
nand U2286 (N_2286,N_2022,N_2089);
and U2287 (N_2287,N_2109,N_2025);
and U2288 (N_2288,N_2119,N_2012);
nor U2289 (N_2289,N_2065,N_2093);
nand U2290 (N_2290,N_2174,N_2160);
xnor U2291 (N_2291,N_2086,N_2042);
xor U2292 (N_2292,N_2143,N_2108);
xor U2293 (N_2293,N_2075,N_2036);
and U2294 (N_2294,N_2046,N_2186);
and U2295 (N_2295,N_2002,N_2195);
or U2296 (N_2296,N_2198,N_2080);
or U2297 (N_2297,N_2190,N_2166);
nor U2298 (N_2298,N_2105,N_2017);
and U2299 (N_2299,N_2152,N_2053);
xor U2300 (N_2300,N_2126,N_2188);
nand U2301 (N_2301,N_2091,N_2121);
and U2302 (N_2302,N_2046,N_2195);
xor U2303 (N_2303,N_2110,N_2025);
or U2304 (N_2304,N_2188,N_2037);
xnor U2305 (N_2305,N_2038,N_2095);
nand U2306 (N_2306,N_2037,N_2055);
and U2307 (N_2307,N_2128,N_2016);
nor U2308 (N_2308,N_2093,N_2073);
or U2309 (N_2309,N_2049,N_2112);
nor U2310 (N_2310,N_2025,N_2166);
xor U2311 (N_2311,N_2099,N_2056);
nand U2312 (N_2312,N_2090,N_2185);
nor U2313 (N_2313,N_2119,N_2054);
xor U2314 (N_2314,N_2014,N_2066);
nor U2315 (N_2315,N_2050,N_2197);
and U2316 (N_2316,N_2013,N_2021);
nand U2317 (N_2317,N_2170,N_2004);
or U2318 (N_2318,N_2137,N_2028);
and U2319 (N_2319,N_2127,N_2133);
xnor U2320 (N_2320,N_2103,N_2059);
or U2321 (N_2321,N_2007,N_2045);
nand U2322 (N_2322,N_2041,N_2187);
nand U2323 (N_2323,N_2066,N_2199);
nand U2324 (N_2324,N_2087,N_2155);
nor U2325 (N_2325,N_2192,N_2036);
nand U2326 (N_2326,N_2104,N_2094);
nand U2327 (N_2327,N_2074,N_2090);
and U2328 (N_2328,N_2041,N_2085);
nand U2329 (N_2329,N_2174,N_2180);
nor U2330 (N_2330,N_2054,N_2127);
and U2331 (N_2331,N_2199,N_2104);
or U2332 (N_2332,N_2053,N_2024);
nand U2333 (N_2333,N_2039,N_2181);
xor U2334 (N_2334,N_2177,N_2116);
and U2335 (N_2335,N_2096,N_2008);
or U2336 (N_2336,N_2098,N_2188);
and U2337 (N_2337,N_2004,N_2135);
and U2338 (N_2338,N_2027,N_2162);
or U2339 (N_2339,N_2056,N_2139);
xnor U2340 (N_2340,N_2189,N_2044);
or U2341 (N_2341,N_2194,N_2066);
or U2342 (N_2342,N_2066,N_2078);
or U2343 (N_2343,N_2168,N_2158);
nand U2344 (N_2344,N_2154,N_2151);
and U2345 (N_2345,N_2164,N_2198);
nor U2346 (N_2346,N_2140,N_2185);
xnor U2347 (N_2347,N_2175,N_2030);
xnor U2348 (N_2348,N_2104,N_2181);
xor U2349 (N_2349,N_2115,N_2119);
nor U2350 (N_2350,N_2013,N_2188);
or U2351 (N_2351,N_2152,N_2101);
nand U2352 (N_2352,N_2035,N_2163);
nand U2353 (N_2353,N_2120,N_2099);
and U2354 (N_2354,N_2006,N_2190);
xnor U2355 (N_2355,N_2105,N_2062);
nand U2356 (N_2356,N_2062,N_2029);
nor U2357 (N_2357,N_2089,N_2125);
nor U2358 (N_2358,N_2012,N_2111);
nand U2359 (N_2359,N_2044,N_2119);
xor U2360 (N_2360,N_2034,N_2047);
nand U2361 (N_2361,N_2182,N_2075);
nor U2362 (N_2362,N_2175,N_2137);
or U2363 (N_2363,N_2027,N_2144);
xnor U2364 (N_2364,N_2121,N_2097);
and U2365 (N_2365,N_2055,N_2143);
and U2366 (N_2366,N_2018,N_2062);
xnor U2367 (N_2367,N_2170,N_2049);
xnor U2368 (N_2368,N_2055,N_2015);
xnor U2369 (N_2369,N_2147,N_2163);
nor U2370 (N_2370,N_2041,N_2137);
or U2371 (N_2371,N_2093,N_2145);
xnor U2372 (N_2372,N_2110,N_2183);
nor U2373 (N_2373,N_2138,N_2037);
nand U2374 (N_2374,N_2019,N_2116);
xor U2375 (N_2375,N_2187,N_2051);
or U2376 (N_2376,N_2189,N_2127);
xor U2377 (N_2377,N_2036,N_2048);
or U2378 (N_2378,N_2149,N_2130);
nor U2379 (N_2379,N_2090,N_2083);
nand U2380 (N_2380,N_2076,N_2100);
nor U2381 (N_2381,N_2142,N_2026);
and U2382 (N_2382,N_2075,N_2029);
and U2383 (N_2383,N_2039,N_2032);
xnor U2384 (N_2384,N_2116,N_2131);
and U2385 (N_2385,N_2017,N_2071);
and U2386 (N_2386,N_2153,N_2150);
xor U2387 (N_2387,N_2191,N_2132);
nand U2388 (N_2388,N_2190,N_2161);
xor U2389 (N_2389,N_2014,N_2160);
xnor U2390 (N_2390,N_2183,N_2059);
or U2391 (N_2391,N_2171,N_2166);
nand U2392 (N_2392,N_2075,N_2068);
or U2393 (N_2393,N_2174,N_2045);
or U2394 (N_2394,N_2091,N_2033);
xor U2395 (N_2395,N_2074,N_2097);
nand U2396 (N_2396,N_2188,N_2085);
nor U2397 (N_2397,N_2020,N_2160);
xnor U2398 (N_2398,N_2049,N_2071);
or U2399 (N_2399,N_2008,N_2158);
or U2400 (N_2400,N_2354,N_2312);
nor U2401 (N_2401,N_2352,N_2249);
or U2402 (N_2402,N_2381,N_2275);
or U2403 (N_2403,N_2327,N_2245);
and U2404 (N_2404,N_2330,N_2271);
xnor U2405 (N_2405,N_2278,N_2235);
nand U2406 (N_2406,N_2389,N_2355);
and U2407 (N_2407,N_2399,N_2290);
nor U2408 (N_2408,N_2370,N_2234);
xor U2409 (N_2409,N_2241,N_2270);
or U2410 (N_2410,N_2340,N_2344);
or U2411 (N_2411,N_2374,N_2291);
nand U2412 (N_2412,N_2246,N_2227);
xnor U2413 (N_2413,N_2223,N_2318);
xor U2414 (N_2414,N_2390,N_2393);
nand U2415 (N_2415,N_2277,N_2365);
nand U2416 (N_2416,N_2301,N_2283);
nor U2417 (N_2417,N_2204,N_2305);
nand U2418 (N_2418,N_2345,N_2348);
and U2419 (N_2419,N_2296,N_2308);
or U2420 (N_2420,N_2297,N_2351);
or U2421 (N_2421,N_2218,N_2242);
nand U2422 (N_2422,N_2266,N_2203);
or U2423 (N_2423,N_2337,N_2251);
nor U2424 (N_2424,N_2237,N_2284);
nand U2425 (N_2425,N_2201,N_2346);
nand U2426 (N_2426,N_2213,N_2230);
and U2427 (N_2427,N_2379,N_2261);
nand U2428 (N_2428,N_2252,N_2395);
xor U2429 (N_2429,N_2356,N_2363);
nand U2430 (N_2430,N_2384,N_2216);
nor U2431 (N_2431,N_2286,N_2396);
nand U2432 (N_2432,N_2322,N_2397);
nand U2433 (N_2433,N_2229,N_2289);
and U2434 (N_2434,N_2281,N_2273);
and U2435 (N_2435,N_2364,N_2336);
nand U2436 (N_2436,N_2300,N_2255);
xnor U2437 (N_2437,N_2220,N_2309);
nand U2438 (N_2438,N_2238,N_2367);
or U2439 (N_2439,N_2285,N_2315);
or U2440 (N_2440,N_2302,N_2372);
or U2441 (N_2441,N_2321,N_2332);
nand U2442 (N_2442,N_2293,N_2298);
xnor U2443 (N_2443,N_2398,N_2225);
nor U2444 (N_2444,N_2392,N_2299);
nand U2445 (N_2445,N_2314,N_2265);
and U2446 (N_2446,N_2208,N_2373);
and U2447 (N_2447,N_2279,N_2377);
and U2448 (N_2448,N_2232,N_2259);
and U2449 (N_2449,N_2347,N_2219);
or U2450 (N_2450,N_2385,N_2316);
nor U2451 (N_2451,N_2335,N_2207);
xor U2452 (N_2452,N_2268,N_2215);
or U2453 (N_2453,N_2280,N_2254);
and U2454 (N_2454,N_2211,N_2228);
xnor U2455 (N_2455,N_2256,N_2383);
xnor U2456 (N_2456,N_2292,N_2317);
and U2457 (N_2457,N_2349,N_2366);
or U2458 (N_2458,N_2307,N_2224);
or U2459 (N_2459,N_2386,N_2391);
nor U2460 (N_2460,N_2304,N_2325);
nor U2461 (N_2461,N_2288,N_2212);
nand U2462 (N_2462,N_2388,N_2310);
or U2463 (N_2463,N_2360,N_2357);
or U2464 (N_2464,N_2264,N_2324);
xor U2465 (N_2465,N_2331,N_2358);
nor U2466 (N_2466,N_2319,N_2303);
nand U2467 (N_2467,N_2353,N_2250);
nor U2468 (N_2468,N_2338,N_2295);
nand U2469 (N_2469,N_2326,N_2329);
nand U2470 (N_2470,N_2267,N_2244);
xnor U2471 (N_2471,N_2239,N_2282);
nand U2472 (N_2472,N_2368,N_2214);
nand U2473 (N_2473,N_2362,N_2306);
and U2474 (N_2474,N_2236,N_2378);
or U2475 (N_2475,N_2287,N_2339);
nor U2476 (N_2476,N_2313,N_2311);
nand U2477 (N_2477,N_2272,N_2342);
nand U2478 (N_2478,N_2217,N_2320);
and U2479 (N_2479,N_2200,N_2269);
xor U2480 (N_2480,N_2240,N_2253);
or U2481 (N_2481,N_2209,N_2359);
xor U2482 (N_2482,N_2323,N_2233);
or U2483 (N_2483,N_2262,N_2263);
nor U2484 (N_2484,N_2202,N_2247);
nor U2485 (N_2485,N_2371,N_2206);
and U2486 (N_2486,N_2380,N_2334);
nor U2487 (N_2487,N_2382,N_2222);
nand U2488 (N_2488,N_2210,N_2369);
nand U2489 (N_2489,N_2260,N_2394);
nor U2490 (N_2490,N_2376,N_2231);
xnor U2491 (N_2491,N_2333,N_2375);
nor U2492 (N_2492,N_2258,N_2341);
or U2493 (N_2493,N_2221,N_2361);
nor U2494 (N_2494,N_2205,N_2226);
or U2495 (N_2495,N_2294,N_2343);
and U2496 (N_2496,N_2243,N_2328);
and U2497 (N_2497,N_2350,N_2387);
xnor U2498 (N_2498,N_2276,N_2248);
nor U2499 (N_2499,N_2274,N_2257);
and U2500 (N_2500,N_2266,N_2208);
nand U2501 (N_2501,N_2273,N_2373);
nand U2502 (N_2502,N_2235,N_2206);
xnor U2503 (N_2503,N_2212,N_2275);
or U2504 (N_2504,N_2380,N_2238);
and U2505 (N_2505,N_2304,N_2294);
nand U2506 (N_2506,N_2218,N_2203);
and U2507 (N_2507,N_2349,N_2312);
or U2508 (N_2508,N_2200,N_2292);
nand U2509 (N_2509,N_2368,N_2359);
or U2510 (N_2510,N_2376,N_2230);
nand U2511 (N_2511,N_2300,N_2211);
or U2512 (N_2512,N_2317,N_2275);
xnor U2513 (N_2513,N_2366,N_2238);
nor U2514 (N_2514,N_2319,N_2285);
nor U2515 (N_2515,N_2329,N_2317);
and U2516 (N_2516,N_2296,N_2325);
nor U2517 (N_2517,N_2334,N_2234);
or U2518 (N_2518,N_2304,N_2244);
xnor U2519 (N_2519,N_2317,N_2346);
and U2520 (N_2520,N_2223,N_2301);
or U2521 (N_2521,N_2327,N_2313);
nand U2522 (N_2522,N_2365,N_2305);
nor U2523 (N_2523,N_2335,N_2323);
nor U2524 (N_2524,N_2283,N_2316);
or U2525 (N_2525,N_2228,N_2210);
nor U2526 (N_2526,N_2337,N_2330);
nand U2527 (N_2527,N_2288,N_2277);
xor U2528 (N_2528,N_2299,N_2382);
nor U2529 (N_2529,N_2319,N_2207);
nor U2530 (N_2530,N_2277,N_2259);
nand U2531 (N_2531,N_2397,N_2396);
nor U2532 (N_2532,N_2320,N_2356);
nor U2533 (N_2533,N_2292,N_2222);
xnor U2534 (N_2534,N_2392,N_2221);
nand U2535 (N_2535,N_2282,N_2396);
nand U2536 (N_2536,N_2278,N_2329);
xor U2537 (N_2537,N_2373,N_2335);
and U2538 (N_2538,N_2268,N_2255);
and U2539 (N_2539,N_2204,N_2310);
nand U2540 (N_2540,N_2201,N_2282);
and U2541 (N_2541,N_2298,N_2271);
and U2542 (N_2542,N_2327,N_2332);
and U2543 (N_2543,N_2275,N_2220);
nand U2544 (N_2544,N_2230,N_2361);
xnor U2545 (N_2545,N_2380,N_2384);
xor U2546 (N_2546,N_2268,N_2305);
nor U2547 (N_2547,N_2312,N_2229);
or U2548 (N_2548,N_2246,N_2376);
xor U2549 (N_2549,N_2205,N_2206);
nor U2550 (N_2550,N_2295,N_2382);
nand U2551 (N_2551,N_2328,N_2377);
nor U2552 (N_2552,N_2355,N_2279);
and U2553 (N_2553,N_2395,N_2202);
xnor U2554 (N_2554,N_2294,N_2369);
nor U2555 (N_2555,N_2226,N_2370);
or U2556 (N_2556,N_2342,N_2220);
and U2557 (N_2557,N_2233,N_2368);
nand U2558 (N_2558,N_2282,N_2389);
or U2559 (N_2559,N_2311,N_2336);
xnor U2560 (N_2560,N_2282,N_2309);
nand U2561 (N_2561,N_2310,N_2214);
or U2562 (N_2562,N_2309,N_2235);
xnor U2563 (N_2563,N_2381,N_2291);
xnor U2564 (N_2564,N_2290,N_2267);
nand U2565 (N_2565,N_2223,N_2283);
and U2566 (N_2566,N_2374,N_2372);
xnor U2567 (N_2567,N_2216,N_2211);
xor U2568 (N_2568,N_2390,N_2212);
nor U2569 (N_2569,N_2347,N_2339);
nand U2570 (N_2570,N_2314,N_2390);
xnor U2571 (N_2571,N_2224,N_2242);
and U2572 (N_2572,N_2300,N_2360);
nand U2573 (N_2573,N_2378,N_2314);
xnor U2574 (N_2574,N_2231,N_2200);
and U2575 (N_2575,N_2238,N_2397);
xnor U2576 (N_2576,N_2219,N_2350);
nor U2577 (N_2577,N_2216,N_2298);
and U2578 (N_2578,N_2202,N_2337);
nand U2579 (N_2579,N_2352,N_2208);
and U2580 (N_2580,N_2296,N_2278);
and U2581 (N_2581,N_2303,N_2307);
and U2582 (N_2582,N_2227,N_2232);
nand U2583 (N_2583,N_2236,N_2391);
xnor U2584 (N_2584,N_2293,N_2303);
or U2585 (N_2585,N_2309,N_2332);
xor U2586 (N_2586,N_2301,N_2210);
xor U2587 (N_2587,N_2261,N_2269);
nand U2588 (N_2588,N_2278,N_2219);
or U2589 (N_2589,N_2394,N_2247);
or U2590 (N_2590,N_2238,N_2336);
and U2591 (N_2591,N_2351,N_2264);
nor U2592 (N_2592,N_2229,N_2369);
nand U2593 (N_2593,N_2252,N_2277);
and U2594 (N_2594,N_2367,N_2225);
and U2595 (N_2595,N_2351,N_2298);
or U2596 (N_2596,N_2283,N_2306);
nor U2597 (N_2597,N_2200,N_2301);
or U2598 (N_2598,N_2386,N_2286);
xor U2599 (N_2599,N_2282,N_2208);
or U2600 (N_2600,N_2415,N_2472);
nor U2601 (N_2601,N_2450,N_2526);
nor U2602 (N_2602,N_2439,N_2483);
nor U2603 (N_2603,N_2507,N_2473);
nor U2604 (N_2604,N_2531,N_2422);
or U2605 (N_2605,N_2591,N_2594);
nor U2606 (N_2606,N_2486,N_2465);
nor U2607 (N_2607,N_2420,N_2452);
and U2608 (N_2608,N_2555,N_2470);
xor U2609 (N_2609,N_2424,N_2409);
xor U2610 (N_2610,N_2417,N_2532);
and U2611 (N_2611,N_2568,N_2413);
nor U2612 (N_2612,N_2525,N_2504);
or U2613 (N_2613,N_2448,N_2400);
nand U2614 (N_2614,N_2442,N_2463);
nand U2615 (N_2615,N_2449,N_2534);
xnor U2616 (N_2616,N_2597,N_2547);
nor U2617 (N_2617,N_2469,N_2427);
xor U2618 (N_2618,N_2493,N_2587);
and U2619 (N_2619,N_2476,N_2481);
and U2620 (N_2620,N_2518,N_2574);
xnor U2621 (N_2621,N_2474,N_2535);
and U2622 (N_2622,N_2460,N_2468);
and U2623 (N_2623,N_2593,N_2499);
or U2624 (N_2624,N_2519,N_2479);
or U2625 (N_2625,N_2540,N_2436);
nor U2626 (N_2626,N_2488,N_2599);
nor U2627 (N_2627,N_2515,N_2596);
xor U2628 (N_2628,N_2494,N_2572);
or U2629 (N_2629,N_2554,N_2458);
xor U2630 (N_2630,N_2423,N_2576);
nor U2631 (N_2631,N_2431,N_2502);
xnor U2632 (N_2632,N_2434,N_2524);
xnor U2633 (N_2633,N_2557,N_2529);
nand U2634 (N_2634,N_2471,N_2567);
nand U2635 (N_2635,N_2435,N_2545);
nand U2636 (N_2636,N_2402,N_2560);
nand U2637 (N_2637,N_2577,N_2404);
or U2638 (N_2638,N_2497,N_2491);
or U2639 (N_2639,N_2520,N_2513);
or U2640 (N_2640,N_2405,N_2583);
and U2641 (N_2641,N_2533,N_2563);
xnor U2642 (N_2642,N_2457,N_2541);
xor U2643 (N_2643,N_2501,N_2408);
nand U2644 (N_2644,N_2522,N_2406);
nand U2645 (N_2645,N_2482,N_2584);
nor U2646 (N_2646,N_2517,N_2553);
nor U2647 (N_2647,N_2503,N_2546);
or U2648 (N_2648,N_2445,N_2419);
or U2649 (N_2649,N_2489,N_2530);
nand U2650 (N_2650,N_2425,N_2536);
nand U2651 (N_2651,N_2411,N_2559);
or U2652 (N_2652,N_2464,N_2564);
or U2653 (N_2653,N_2573,N_2492);
and U2654 (N_2654,N_2508,N_2510);
xnor U2655 (N_2655,N_2490,N_2509);
xnor U2656 (N_2656,N_2432,N_2523);
xor U2657 (N_2657,N_2443,N_2556);
nor U2658 (N_2658,N_2585,N_2410);
nor U2659 (N_2659,N_2544,N_2480);
nand U2660 (N_2660,N_2542,N_2444);
nand U2661 (N_2661,N_2462,N_2551);
xor U2662 (N_2662,N_2412,N_2438);
xnor U2663 (N_2663,N_2552,N_2477);
xnor U2664 (N_2664,N_2571,N_2485);
or U2665 (N_2665,N_2569,N_2511);
and U2666 (N_2666,N_2516,N_2418);
nor U2667 (N_2667,N_2421,N_2550);
or U2668 (N_2668,N_2426,N_2433);
nor U2669 (N_2669,N_2447,N_2401);
and U2670 (N_2670,N_2498,N_2500);
or U2671 (N_2671,N_2437,N_2527);
nor U2672 (N_2672,N_2588,N_2538);
nor U2673 (N_2673,N_2566,N_2440);
nand U2674 (N_2674,N_2496,N_2451);
or U2675 (N_2675,N_2561,N_2595);
xor U2676 (N_2676,N_2586,N_2407);
xnor U2677 (N_2677,N_2580,N_2429);
xnor U2678 (N_2678,N_2598,N_2570);
nor U2679 (N_2679,N_2543,N_2428);
nand U2680 (N_2680,N_2506,N_2505);
nand U2681 (N_2681,N_2467,N_2549);
nor U2682 (N_2682,N_2446,N_2558);
nand U2683 (N_2683,N_2466,N_2456);
nand U2684 (N_2684,N_2487,N_2453);
nand U2685 (N_2685,N_2459,N_2539);
nand U2686 (N_2686,N_2416,N_2562);
nor U2687 (N_2687,N_2537,N_2575);
nand U2688 (N_2688,N_2454,N_2578);
nor U2689 (N_2689,N_2592,N_2582);
and U2690 (N_2690,N_2495,N_2528);
or U2691 (N_2691,N_2441,N_2521);
nor U2692 (N_2692,N_2590,N_2565);
nand U2693 (N_2693,N_2589,N_2484);
or U2694 (N_2694,N_2512,N_2478);
or U2695 (N_2695,N_2403,N_2579);
or U2696 (N_2696,N_2514,N_2455);
or U2697 (N_2697,N_2414,N_2430);
nand U2698 (N_2698,N_2548,N_2461);
and U2699 (N_2699,N_2475,N_2581);
xnor U2700 (N_2700,N_2443,N_2425);
and U2701 (N_2701,N_2495,N_2445);
and U2702 (N_2702,N_2564,N_2473);
nand U2703 (N_2703,N_2473,N_2556);
or U2704 (N_2704,N_2415,N_2466);
nor U2705 (N_2705,N_2450,N_2524);
nor U2706 (N_2706,N_2502,N_2541);
or U2707 (N_2707,N_2514,N_2577);
nand U2708 (N_2708,N_2465,N_2435);
and U2709 (N_2709,N_2507,N_2461);
nor U2710 (N_2710,N_2524,N_2462);
nand U2711 (N_2711,N_2564,N_2509);
or U2712 (N_2712,N_2406,N_2552);
and U2713 (N_2713,N_2414,N_2438);
or U2714 (N_2714,N_2515,N_2514);
nor U2715 (N_2715,N_2463,N_2546);
nand U2716 (N_2716,N_2411,N_2505);
nand U2717 (N_2717,N_2525,N_2471);
or U2718 (N_2718,N_2595,N_2495);
xor U2719 (N_2719,N_2469,N_2428);
or U2720 (N_2720,N_2401,N_2514);
and U2721 (N_2721,N_2530,N_2557);
nor U2722 (N_2722,N_2463,N_2518);
and U2723 (N_2723,N_2408,N_2524);
nor U2724 (N_2724,N_2406,N_2593);
nor U2725 (N_2725,N_2575,N_2546);
nor U2726 (N_2726,N_2428,N_2479);
nor U2727 (N_2727,N_2460,N_2502);
nor U2728 (N_2728,N_2505,N_2540);
nand U2729 (N_2729,N_2483,N_2505);
or U2730 (N_2730,N_2430,N_2499);
nor U2731 (N_2731,N_2491,N_2478);
and U2732 (N_2732,N_2561,N_2530);
nand U2733 (N_2733,N_2427,N_2416);
or U2734 (N_2734,N_2472,N_2436);
nor U2735 (N_2735,N_2493,N_2442);
xor U2736 (N_2736,N_2477,N_2402);
or U2737 (N_2737,N_2533,N_2488);
nor U2738 (N_2738,N_2531,N_2552);
nand U2739 (N_2739,N_2571,N_2517);
or U2740 (N_2740,N_2599,N_2462);
nand U2741 (N_2741,N_2552,N_2422);
nor U2742 (N_2742,N_2404,N_2456);
xor U2743 (N_2743,N_2416,N_2524);
or U2744 (N_2744,N_2417,N_2582);
xnor U2745 (N_2745,N_2547,N_2592);
xor U2746 (N_2746,N_2566,N_2537);
nand U2747 (N_2747,N_2541,N_2555);
and U2748 (N_2748,N_2537,N_2420);
nor U2749 (N_2749,N_2559,N_2498);
nor U2750 (N_2750,N_2540,N_2536);
or U2751 (N_2751,N_2441,N_2540);
nor U2752 (N_2752,N_2522,N_2495);
and U2753 (N_2753,N_2430,N_2512);
xor U2754 (N_2754,N_2479,N_2440);
xor U2755 (N_2755,N_2574,N_2490);
nand U2756 (N_2756,N_2557,N_2540);
nor U2757 (N_2757,N_2547,N_2447);
nor U2758 (N_2758,N_2526,N_2441);
or U2759 (N_2759,N_2553,N_2455);
nor U2760 (N_2760,N_2465,N_2436);
or U2761 (N_2761,N_2404,N_2563);
nand U2762 (N_2762,N_2546,N_2587);
nor U2763 (N_2763,N_2526,N_2496);
or U2764 (N_2764,N_2494,N_2599);
nand U2765 (N_2765,N_2506,N_2507);
nand U2766 (N_2766,N_2473,N_2429);
xor U2767 (N_2767,N_2576,N_2556);
and U2768 (N_2768,N_2489,N_2579);
nor U2769 (N_2769,N_2434,N_2596);
and U2770 (N_2770,N_2439,N_2432);
xnor U2771 (N_2771,N_2498,N_2459);
and U2772 (N_2772,N_2487,N_2445);
nor U2773 (N_2773,N_2486,N_2566);
nand U2774 (N_2774,N_2512,N_2558);
nor U2775 (N_2775,N_2559,N_2533);
or U2776 (N_2776,N_2515,N_2412);
and U2777 (N_2777,N_2481,N_2418);
xor U2778 (N_2778,N_2437,N_2530);
and U2779 (N_2779,N_2598,N_2400);
xnor U2780 (N_2780,N_2536,N_2434);
or U2781 (N_2781,N_2599,N_2445);
and U2782 (N_2782,N_2402,N_2414);
or U2783 (N_2783,N_2436,N_2493);
and U2784 (N_2784,N_2488,N_2494);
or U2785 (N_2785,N_2403,N_2417);
nand U2786 (N_2786,N_2477,N_2413);
or U2787 (N_2787,N_2557,N_2438);
nand U2788 (N_2788,N_2473,N_2516);
xnor U2789 (N_2789,N_2497,N_2566);
xor U2790 (N_2790,N_2580,N_2401);
xnor U2791 (N_2791,N_2460,N_2466);
nor U2792 (N_2792,N_2538,N_2412);
nand U2793 (N_2793,N_2515,N_2523);
or U2794 (N_2794,N_2472,N_2507);
and U2795 (N_2795,N_2503,N_2490);
and U2796 (N_2796,N_2528,N_2413);
and U2797 (N_2797,N_2428,N_2558);
xor U2798 (N_2798,N_2538,N_2586);
or U2799 (N_2799,N_2451,N_2423);
xnor U2800 (N_2800,N_2760,N_2645);
nand U2801 (N_2801,N_2690,N_2679);
nor U2802 (N_2802,N_2661,N_2719);
and U2803 (N_2803,N_2635,N_2754);
or U2804 (N_2804,N_2771,N_2723);
or U2805 (N_2805,N_2693,N_2604);
xor U2806 (N_2806,N_2713,N_2736);
or U2807 (N_2807,N_2660,N_2772);
nor U2808 (N_2808,N_2765,N_2640);
xnor U2809 (N_2809,N_2721,N_2764);
and U2810 (N_2810,N_2676,N_2618);
and U2811 (N_2811,N_2731,N_2658);
nor U2812 (N_2812,N_2681,N_2694);
or U2813 (N_2813,N_2727,N_2770);
and U2814 (N_2814,N_2610,N_2733);
nand U2815 (N_2815,N_2725,N_2662);
xnor U2816 (N_2816,N_2687,N_2631);
or U2817 (N_2817,N_2684,N_2778);
nand U2818 (N_2818,N_2705,N_2626);
nor U2819 (N_2819,N_2619,N_2709);
nand U2820 (N_2820,N_2683,N_2794);
xnor U2821 (N_2821,N_2691,N_2606);
nand U2822 (N_2822,N_2643,N_2649);
nand U2823 (N_2823,N_2628,N_2665);
xor U2824 (N_2824,N_2629,N_2769);
and U2825 (N_2825,N_2624,N_2701);
xnor U2826 (N_2826,N_2680,N_2663);
xnor U2827 (N_2827,N_2755,N_2668);
xnor U2828 (N_2828,N_2766,N_2703);
and U2829 (N_2829,N_2729,N_2603);
and U2830 (N_2830,N_2792,N_2720);
or U2831 (N_2831,N_2704,N_2734);
xnor U2832 (N_2832,N_2717,N_2666);
or U2833 (N_2833,N_2762,N_2667);
nand U2834 (N_2834,N_2656,N_2797);
xnor U2835 (N_2835,N_2614,N_2671);
or U2836 (N_2836,N_2632,N_2622);
nand U2837 (N_2837,N_2742,N_2669);
nand U2838 (N_2838,N_2642,N_2695);
nand U2839 (N_2839,N_2747,N_2777);
nor U2840 (N_2840,N_2633,N_2746);
and U2841 (N_2841,N_2767,N_2616);
xnor U2842 (N_2842,N_2753,N_2637);
or U2843 (N_2843,N_2735,N_2763);
and U2844 (N_2844,N_2796,N_2609);
nor U2845 (N_2845,N_2788,N_2607);
nand U2846 (N_2846,N_2795,N_2710);
and U2847 (N_2847,N_2784,N_2670);
xnor U2848 (N_2848,N_2786,N_2749);
nand U2849 (N_2849,N_2756,N_2608);
nor U2850 (N_2850,N_2636,N_2790);
and U2851 (N_2851,N_2780,N_2634);
and U2852 (N_2852,N_2706,N_2648);
or U2853 (N_2853,N_2711,N_2715);
or U2854 (N_2854,N_2673,N_2782);
nand U2855 (N_2855,N_2600,N_2601);
or U2856 (N_2856,N_2689,N_2657);
or U2857 (N_2857,N_2625,N_2617);
xor U2858 (N_2858,N_2730,N_2664);
and U2859 (N_2859,N_2718,N_2650);
xor U2860 (N_2860,N_2744,N_2773);
and U2861 (N_2861,N_2728,N_2696);
or U2862 (N_2862,N_2682,N_2743);
nand U2863 (N_2863,N_2612,N_2737);
and U2864 (N_2864,N_2761,N_2707);
and U2865 (N_2865,N_2674,N_2787);
nand U2866 (N_2866,N_2639,N_2686);
and U2867 (N_2867,N_2702,N_2685);
and U2868 (N_2868,N_2672,N_2698);
and U2869 (N_2869,N_2783,N_2654);
nor U2870 (N_2870,N_2739,N_2789);
and U2871 (N_2871,N_2740,N_2651);
xnor U2872 (N_2872,N_2623,N_2613);
and U2873 (N_2873,N_2630,N_2653);
or U2874 (N_2874,N_2647,N_2757);
nor U2875 (N_2875,N_2605,N_2659);
nor U2876 (N_2876,N_2716,N_2644);
xor U2877 (N_2877,N_2700,N_2714);
nor U2878 (N_2878,N_2750,N_2745);
nand U2879 (N_2879,N_2779,N_2697);
and U2880 (N_2880,N_2675,N_2712);
and U2881 (N_2881,N_2655,N_2620);
nor U2882 (N_2882,N_2621,N_2768);
nand U2883 (N_2883,N_2738,N_2652);
nor U2884 (N_2884,N_2775,N_2726);
nor U2885 (N_2885,N_2692,N_2793);
xnor U2886 (N_2886,N_2646,N_2615);
nand U2887 (N_2887,N_2732,N_2791);
or U2888 (N_2888,N_2722,N_2638);
and U2889 (N_2889,N_2708,N_2781);
nand U2890 (N_2890,N_2799,N_2678);
nand U2891 (N_2891,N_2741,N_2677);
xnor U2892 (N_2892,N_2699,N_2602);
nor U2893 (N_2893,N_2688,N_2627);
xor U2894 (N_2894,N_2758,N_2751);
or U2895 (N_2895,N_2724,N_2785);
nor U2896 (N_2896,N_2611,N_2752);
nor U2897 (N_2897,N_2641,N_2759);
or U2898 (N_2898,N_2774,N_2776);
or U2899 (N_2899,N_2798,N_2748);
xor U2900 (N_2900,N_2742,N_2776);
and U2901 (N_2901,N_2656,N_2717);
nor U2902 (N_2902,N_2709,N_2720);
and U2903 (N_2903,N_2603,N_2635);
and U2904 (N_2904,N_2612,N_2704);
and U2905 (N_2905,N_2721,N_2681);
and U2906 (N_2906,N_2768,N_2620);
nor U2907 (N_2907,N_2720,N_2718);
nand U2908 (N_2908,N_2631,N_2761);
and U2909 (N_2909,N_2659,N_2742);
or U2910 (N_2910,N_2676,N_2651);
or U2911 (N_2911,N_2709,N_2603);
nor U2912 (N_2912,N_2701,N_2712);
nand U2913 (N_2913,N_2745,N_2785);
xnor U2914 (N_2914,N_2772,N_2779);
nand U2915 (N_2915,N_2767,N_2627);
and U2916 (N_2916,N_2745,N_2757);
or U2917 (N_2917,N_2775,N_2734);
nor U2918 (N_2918,N_2771,N_2649);
and U2919 (N_2919,N_2783,N_2795);
or U2920 (N_2920,N_2763,N_2789);
or U2921 (N_2921,N_2609,N_2747);
xor U2922 (N_2922,N_2750,N_2696);
or U2923 (N_2923,N_2786,N_2700);
and U2924 (N_2924,N_2619,N_2787);
xnor U2925 (N_2925,N_2774,N_2689);
nor U2926 (N_2926,N_2666,N_2602);
or U2927 (N_2927,N_2697,N_2795);
nand U2928 (N_2928,N_2645,N_2628);
and U2929 (N_2929,N_2703,N_2633);
and U2930 (N_2930,N_2679,N_2655);
nand U2931 (N_2931,N_2700,N_2701);
or U2932 (N_2932,N_2782,N_2771);
or U2933 (N_2933,N_2607,N_2772);
or U2934 (N_2934,N_2764,N_2760);
and U2935 (N_2935,N_2655,N_2795);
nand U2936 (N_2936,N_2630,N_2716);
nand U2937 (N_2937,N_2773,N_2776);
xor U2938 (N_2938,N_2721,N_2751);
nor U2939 (N_2939,N_2704,N_2710);
xor U2940 (N_2940,N_2710,N_2793);
xor U2941 (N_2941,N_2772,N_2671);
nand U2942 (N_2942,N_2712,N_2700);
or U2943 (N_2943,N_2767,N_2610);
xnor U2944 (N_2944,N_2627,N_2630);
nor U2945 (N_2945,N_2655,N_2721);
nand U2946 (N_2946,N_2603,N_2765);
nand U2947 (N_2947,N_2649,N_2775);
nor U2948 (N_2948,N_2721,N_2762);
nor U2949 (N_2949,N_2799,N_2746);
xor U2950 (N_2950,N_2692,N_2618);
xnor U2951 (N_2951,N_2777,N_2741);
and U2952 (N_2952,N_2723,N_2748);
nand U2953 (N_2953,N_2722,N_2618);
and U2954 (N_2954,N_2703,N_2721);
nand U2955 (N_2955,N_2641,N_2717);
nor U2956 (N_2956,N_2756,N_2625);
xor U2957 (N_2957,N_2653,N_2781);
and U2958 (N_2958,N_2712,N_2648);
nor U2959 (N_2959,N_2758,N_2749);
and U2960 (N_2960,N_2701,N_2633);
or U2961 (N_2961,N_2769,N_2757);
nand U2962 (N_2962,N_2698,N_2777);
and U2963 (N_2963,N_2797,N_2705);
nor U2964 (N_2964,N_2649,N_2689);
nand U2965 (N_2965,N_2653,N_2748);
nor U2966 (N_2966,N_2729,N_2659);
nor U2967 (N_2967,N_2673,N_2624);
xnor U2968 (N_2968,N_2634,N_2716);
nor U2969 (N_2969,N_2711,N_2641);
or U2970 (N_2970,N_2618,N_2627);
and U2971 (N_2971,N_2745,N_2665);
xor U2972 (N_2972,N_2615,N_2798);
or U2973 (N_2973,N_2750,N_2715);
xor U2974 (N_2974,N_2696,N_2706);
nor U2975 (N_2975,N_2637,N_2607);
xor U2976 (N_2976,N_2770,N_2783);
nand U2977 (N_2977,N_2767,N_2746);
nand U2978 (N_2978,N_2675,N_2798);
nor U2979 (N_2979,N_2737,N_2683);
xnor U2980 (N_2980,N_2643,N_2787);
xor U2981 (N_2981,N_2639,N_2652);
or U2982 (N_2982,N_2653,N_2613);
and U2983 (N_2983,N_2636,N_2630);
nor U2984 (N_2984,N_2684,N_2600);
or U2985 (N_2985,N_2690,N_2774);
nor U2986 (N_2986,N_2653,N_2792);
xnor U2987 (N_2987,N_2601,N_2783);
nor U2988 (N_2988,N_2675,N_2613);
nand U2989 (N_2989,N_2649,N_2784);
or U2990 (N_2990,N_2734,N_2752);
xor U2991 (N_2991,N_2653,N_2614);
nand U2992 (N_2992,N_2632,N_2647);
xor U2993 (N_2993,N_2688,N_2632);
xor U2994 (N_2994,N_2621,N_2753);
xnor U2995 (N_2995,N_2748,N_2703);
nand U2996 (N_2996,N_2667,N_2632);
xnor U2997 (N_2997,N_2703,N_2713);
nor U2998 (N_2998,N_2667,N_2781);
and U2999 (N_2999,N_2678,N_2718);
and U3000 (N_3000,N_2920,N_2880);
or U3001 (N_3001,N_2849,N_2881);
xor U3002 (N_3002,N_2898,N_2935);
nor U3003 (N_3003,N_2932,N_2865);
and U3004 (N_3004,N_2887,N_2851);
or U3005 (N_3005,N_2802,N_2815);
nor U3006 (N_3006,N_2919,N_2964);
and U3007 (N_3007,N_2924,N_2936);
nand U3008 (N_3008,N_2985,N_2906);
and U3009 (N_3009,N_2885,N_2943);
nor U3010 (N_3010,N_2941,N_2805);
or U3011 (N_3011,N_2835,N_2808);
and U3012 (N_3012,N_2972,N_2874);
and U3013 (N_3013,N_2965,N_2832);
nor U3014 (N_3014,N_2995,N_2809);
nor U3015 (N_3015,N_2925,N_2939);
or U3016 (N_3016,N_2961,N_2843);
or U3017 (N_3017,N_2928,N_2946);
nand U3018 (N_3018,N_2952,N_2971);
or U3019 (N_3019,N_2822,N_2868);
xor U3020 (N_3020,N_2857,N_2944);
or U3021 (N_3021,N_2947,N_2953);
or U3022 (N_3022,N_2914,N_2876);
or U3023 (N_3023,N_2813,N_2927);
and U3024 (N_3024,N_2890,N_2973);
nand U3025 (N_3025,N_2962,N_2847);
nand U3026 (N_3026,N_2866,N_2888);
or U3027 (N_3027,N_2839,N_2994);
and U3028 (N_3028,N_2875,N_2960);
nand U3029 (N_3029,N_2991,N_2967);
nand U3030 (N_3030,N_2986,N_2903);
or U3031 (N_3031,N_2836,N_2841);
and U3032 (N_3032,N_2891,N_2814);
nor U3033 (N_3033,N_2883,N_2894);
nand U3034 (N_3034,N_2882,N_2979);
nor U3035 (N_3035,N_2864,N_2934);
xnor U3036 (N_3036,N_2917,N_2933);
and U3037 (N_3037,N_2820,N_2913);
and U3038 (N_3038,N_2812,N_2884);
nor U3039 (N_3039,N_2938,N_2869);
xnor U3040 (N_3040,N_2845,N_2833);
xnor U3041 (N_3041,N_2983,N_2918);
nand U3042 (N_3042,N_2873,N_2957);
nor U3043 (N_3043,N_2800,N_2989);
or U3044 (N_3044,N_2877,N_2968);
xor U3045 (N_3045,N_2937,N_2801);
nor U3046 (N_3046,N_2998,N_2823);
xnor U3047 (N_3047,N_2963,N_2811);
or U3048 (N_3048,N_2804,N_2860);
xnor U3049 (N_3049,N_2966,N_2807);
xnor U3050 (N_3050,N_2976,N_2909);
and U3051 (N_3051,N_2827,N_2830);
or U3052 (N_3052,N_2893,N_2879);
nand U3053 (N_3053,N_2980,N_2831);
xnor U3054 (N_3054,N_2855,N_2867);
nand U3055 (N_3055,N_2988,N_2871);
nor U3056 (N_3056,N_2828,N_2949);
and U3057 (N_3057,N_2907,N_2999);
or U3058 (N_3058,N_2886,N_2862);
nor U3059 (N_3059,N_2850,N_2878);
or U3060 (N_3060,N_2911,N_2837);
nand U3061 (N_3061,N_2958,N_2806);
or U3062 (N_3062,N_2978,N_2895);
nand U3063 (N_3063,N_2993,N_2816);
nor U3064 (N_3064,N_2990,N_2940);
nand U3065 (N_3065,N_2861,N_2842);
nor U3066 (N_3066,N_2824,N_2910);
and U3067 (N_3067,N_2840,N_2969);
and U3068 (N_3068,N_2904,N_2955);
nand U3069 (N_3069,N_2977,N_2956);
xnor U3070 (N_3070,N_2829,N_2929);
nand U3071 (N_3071,N_2915,N_2922);
and U3072 (N_3072,N_2970,N_2858);
xor U3073 (N_3073,N_2926,N_2810);
nor U3074 (N_3074,N_2854,N_2902);
and U3075 (N_3075,N_2825,N_2900);
nand U3076 (N_3076,N_2916,N_2846);
xnor U3077 (N_3077,N_2889,N_2859);
xor U3078 (N_3078,N_2844,N_2945);
xnor U3079 (N_3079,N_2872,N_2954);
nor U3080 (N_3080,N_2981,N_2838);
or U3081 (N_3081,N_2848,N_2959);
xor U3082 (N_3082,N_2899,N_2996);
nand U3083 (N_3083,N_2931,N_2817);
nor U3084 (N_3084,N_2897,N_2982);
nand U3085 (N_3085,N_2853,N_2942);
or U3086 (N_3086,N_2975,N_2896);
xor U3087 (N_3087,N_2997,N_2863);
or U3088 (N_3088,N_2923,N_2821);
nor U3089 (N_3089,N_2818,N_2921);
or U3090 (N_3090,N_2901,N_2870);
or U3091 (N_3091,N_2826,N_2856);
nor U3092 (N_3092,N_2803,N_2950);
nor U3093 (N_3093,N_2892,N_2908);
nor U3094 (N_3094,N_2992,N_2912);
and U3095 (N_3095,N_2974,N_2852);
nor U3096 (N_3096,N_2984,N_2905);
or U3097 (N_3097,N_2987,N_2930);
and U3098 (N_3098,N_2951,N_2819);
nand U3099 (N_3099,N_2948,N_2834);
and U3100 (N_3100,N_2813,N_2871);
nand U3101 (N_3101,N_2927,N_2992);
nor U3102 (N_3102,N_2977,N_2911);
and U3103 (N_3103,N_2851,N_2854);
xnor U3104 (N_3104,N_2992,N_2961);
nand U3105 (N_3105,N_2827,N_2919);
and U3106 (N_3106,N_2810,N_2856);
or U3107 (N_3107,N_2868,N_2826);
nor U3108 (N_3108,N_2848,N_2865);
or U3109 (N_3109,N_2951,N_2870);
or U3110 (N_3110,N_2990,N_2804);
or U3111 (N_3111,N_2943,N_2963);
xnor U3112 (N_3112,N_2821,N_2848);
or U3113 (N_3113,N_2974,N_2823);
and U3114 (N_3114,N_2854,N_2908);
or U3115 (N_3115,N_2866,N_2946);
nor U3116 (N_3116,N_2950,N_2808);
nor U3117 (N_3117,N_2802,N_2873);
xor U3118 (N_3118,N_2926,N_2919);
or U3119 (N_3119,N_2824,N_2837);
nand U3120 (N_3120,N_2867,N_2892);
nand U3121 (N_3121,N_2976,N_2865);
or U3122 (N_3122,N_2898,N_2978);
or U3123 (N_3123,N_2871,N_2910);
xnor U3124 (N_3124,N_2969,N_2948);
nor U3125 (N_3125,N_2819,N_2980);
nor U3126 (N_3126,N_2878,N_2968);
and U3127 (N_3127,N_2965,N_2809);
xor U3128 (N_3128,N_2891,N_2903);
nand U3129 (N_3129,N_2972,N_2898);
nand U3130 (N_3130,N_2894,N_2945);
or U3131 (N_3131,N_2975,N_2919);
nor U3132 (N_3132,N_2807,N_2929);
or U3133 (N_3133,N_2937,N_2847);
xor U3134 (N_3134,N_2995,N_2806);
nand U3135 (N_3135,N_2885,N_2894);
nand U3136 (N_3136,N_2976,N_2987);
nor U3137 (N_3137,N_2802,N_2982);
nand U3138 (N_3138,N_2869,N_2898);
nor U3139 (N_3139,N_2935,N_2909);
or U3140 (N_3140,N_2925,N_2951);
nand U3141 (N_3141,N_2941,N_2822);
nand U3142 (N_3142,N_2868,N_2952);
nor U3143 (N_3143,N_2893,N_2823);
and U3144 (N_3144,N_2882,N_2843);
nand U3145 (N_3145,N_2868,N_2861);
or U3146 (N_3146,N_2816,N_2999);
xor U3147 (N_3147,N_2994,N_2945);
xnor U3148 (N_3148,N_2852,N_2927);
xor U3149 (N_3149,N_2816,N_2985);
nor U3150 (N_3150,N_2849,N_2804);
xnor U3151 (N_3151,N_2997,N_2818);
nor U3152 (N_3152,N_2947,N_2820);
nor U3153 (N_3153,N_2813,N_2860);
and U3154 (N_3154,N_2970,N_2977);
and U3155 (N_3155,N_2877,N_2982);
or U3156 (N_3156,N_2889,N_2904);
nand U3157 (N_3157,N_2916,N_2816);
xnor U3158 (N_3158,N_2846,N_2974);
nor U3159 (N_3159,N_2950,N_2924);
xnor U3160 (N_3160,N_2976,N_2910);
xnor U3161 (N_3161,N_2944,N_2988);
nand U3162 (N_3162,N_2852,N_2892);
nand U3163 (N_3163,N_2864,N_2933);
and U3164 (N_3164,N_2881,N_2887);
xnor U3165 (N_3165,N_2839,N_2888);
xor U3166 (N_3166,N_2843,N_2810);
nand U3167 (N_3167,N_2922,N_2956);
or U3168 (N_3168,N_2861,N_2901);
nand U3169 (N_3169,N_2979,N_2850);
or U3170 (N_3170,N_2838,N_2911);
xor U3171 (N_3171,N_2942,N_2802);
nand U3172 (N_3172,N_2910,N_2829);
nor U3173 (N_3173,N_2935,N_2828);
nand U3174 (N_3174,N_2812,N_2931);
or U3175 (N_3175,N_2831,N_2964);
or U3176 (N_3176,N_2926,N_2953);
xor U3177 (N_3177,N_2987,N_2838);
xor U3178 (N_3178,N_2963,N_2860);
and U3179 (N_3179,N_2932,N_2895);
or U3180 (N_3180,N_2884,N_2969);
and U3181 (N_3181,N_2897,N_2881);
nor U3182 (N_3182,N_2890,N_2938);
nor U3183 (N_3183,N_2987,N_2889);
and U3184 (N_3184,N_2907,N_2919);
nand U3185 (N_3185,N_2874,N_2955);
nor U3186 (N_3186,N_2821,N_2887);
xor U3187 (N_3187,N_2936,N_2882);
nor U3188 (N_3188,N_2962,N_2845);
and U3189 (N_3189,N_2965,N_2856);
and U3190 (N_3190,N_2932,N_2909);
xnor U3191 (N_3191,N_2937,N_2835);
nand U3192 (N_3192,N_2896,N_2800);
and U3193 (N_3193,N_2962,N_2834);
nor U3194 (N_3194,N_2992,N_2832);
nor U3195 (N_3195,N_2819,N_2968);
or U3196 (N_3196,N_2911,N_2874);
xor U3197 (N_3197,N_2947,N_2930);
nand U3198 (N_3198,N_2952,N_2866);
nand U3199 (N_3199,N_2925,N_2954);
nand U3200 (N_3200,N_3094,N_3192);
nand U3201 (N_3201,N_3175,N_3055);
nand U3202 (N_3202,N_3091,N_3116);
nor U3203 (N_3203,N_3155,N_3095);
xor U3204 (N_3204,N_3005,N_3132);
or U3205 (N_3205,N_3195,N_3032);
nor U3206 (N_3206,N_3072,N_3003);
xnor U3207 (N_3207,N_3104,N_3172);
or U3208 (N_3208,N_3142,N_3141);
nand U3209 (N_3209,N_3148,N_3147);
and U3210 (N_3210,N_3149,N_3133);
or U3211 (N_3211,N_3051,N_3182);
or U3212 (N_3212,N_3135,N_3043);
nor U3213 (N_3213,N_3040,N_3009);
xnor U3214 (N_3214,N_3093,N_3159);
xnor U3215 (N_3215,N_3008,N_3052);
xor U3216 (N_3216,N_3160,N_3112);
and U3217 (N_3217,N_3037,N_3111);
nor U3218 (N_3218,N_3083,N_3146);
xnor U3219 (N_3219,N_3176,N_3174);
nand U3220 (N_3220,N_3013,N_3106);
or U3221 (N_3221,N_3026,N_3157);
nand U3222 (N_3222,N_3066,N_3161);
xor U3223 (N_3223,N_3049,N_3011);
xnor U3224 (N_3224,N_3022,N_3084);
nand U3225 (N_3225,N_3124,N_3001);
nor U3226 (N_3226,N_3020,N_3016);
or U3227 (N_3227,N_3163,N_3186);
nor U3228 (N_3228,N_3087,N_3136);
xor U3229 (N_3229,N_3024,N_3030);
or U3230 (N_3230,N_3127,N_3078);
and U3231 (N_3231,N_3027,N_3038);
or U3232 (N_3232,N_3102,N_3025);
nor U3233 (N_3233,N_3173,N_3140);
nor U3234 (N_3234,N_3113,N_3057);
nand U3235 (N_3235,N_3041,N_3123);
nor U3236 (N_3236,N_3070,N_3126);
nor U3237 (N_3237,N_3031,N_3180);
nand U3238 (N_3238,N_3118,N_3082);
nand U3239 (N_3239,N_3048,N_3061);
and U3240 (N_3240,N_3117,N_3007);
nor U3241 (N_3241,N_3198,N_3179);
nor U3242 (N_3242,N_3134,N_3000);
nor U3243 (N_3243,N_3045,N_3191);
xnor U3244 (N_3244,N_3099,N_3079);
or U3245 (N_3245,N_3137,N_3101);
or U3246 (N_3246,N_3164,N_3128);
and U3247 (N_3247,N_3125,N_3019);
nand U3248 (N_3248,N_3119,N_3139);
nand U3249 (N_3249,N_3196,N_3089);
or U3250 (N_3250,N_3122,N_3108);
xnor U3251 (N_3251,N_3050,N_3171);
nand U3252 (N_3252,N_3075,N_3188);
xor U3253 (N_3253,N_3184,N_3002);
xnor U3254 (N_3254,N_3120,N_3042);
nand U3255 (N_3255,N_3017,N_3081);
or U3256 (N_3256,N_3073,N_3097);
nand U3257 (N_3257,N_3138,N_3162);
xnor U3258 (N_3258,N_3158,N_3100);
nand U3259 (N_3259,N_3088,N_3018);
xnor U3260 (N_3260,N_3069,N_3064);
nand U3261 (N_3261,N_3199,N_3105);
and U3262 (N_3262,N_3154,N_3194);
xnor U3263 (N_3263,N_3044,N_3065);
or U3264 (N_3264,N_3153,N_3189);
nor U3265 (N_3265,N_3115,N_3036);
nand U3266 (N_3266,N_3165,N_3028);
nand U3267 (N_3267,N_3086,N_3144);
and U3268 (N_3268,N_3058,N_3068);
or U3269 (N_3269,N_3033,N_3197);
or U3270 (N_3270,N_3054,N_3143);
and U3271 (N_3271,N_3167,N_3076);
and U3272 (N_3272,N_3130,N_3056);
nand U3273 (N_3273,N_3010,N_3177);
or U3274 (N_3274,N_3023,N_3169);
nand U3275 (N_3275,N_3085,N_3151);
nor U3276 (N_3276,N_3029,N_3187);
xnor U3277 (N_3277,N_3063,N_3014);
or U3278 (N_3278,N_3090,N_3178);
or U3279 (N_3279,N_3152,N_3156);
or U3280 (N_3280,N_3107,N_3166);
or U3281 (N_3281,N_3053,N_3183);
or U3282 (N_3282,N_3067,N_3181);
nand U3283 (N_3283,N_3004,N_3074);
and U3284 (N_3284,N_3190,N_3059);
or U3285 (N_3285,N_3170,N_3109);
nand U3286 (N_3286,N_3098,N_3015);
and U3287 (N_3287,N_3129,N_3092);
nand U3288 (N_3288,N_3021,N_3039);
and U3289 (N_3289,N_3185,N_3103);
xnor U3290 (N_3290,N_3006,N_3034);
xor U3291 (N_3291,N_3193,N_3071);
nor U3292 (N_3292,N_3046,N_3077);
and U3293 (N_3293,N_3110,N_3047);
nor U3294 (N_3294,N_3168,N_3096);
xor U3295 (N_3295,N_3012,N_3150);
or U3296 (N_3296,N_3062,N_3114);
and U3297 (N_3297,N_3145,N_3121);
nand U3298 (N_3298,N_3080,N_3035);
nand U3299 (N_3299,N_3060,N_3131);
nor U3300 (N_3300,N_3013,N_3056);
nor U3301 (N_3301,N_3195,N_3095);
and U3302 (N_3302,N_3030,N_3097);
nand U3303 (N_3303,N_3115,N_3024);
nand U3304 (N_3304,N_3165,N_3181);
or U3305 (N_3305,N_3001,N_3092);
xnor U3306 (N_3306,N_3156,N_3186);
or U3307 (N_3307,N_3133,N_3106);
xnor U3308 (N_3308,N_3089,N_3038);
nor U3309 (N_3309,N_3011,N_3062);
nand U3310 (N_3310,N_3189,N_3157);
and U3311 (N_3311,N_3152,N_3046);
nand U3312 (N_3312,N_3137,N_3039);
xnor U3313 (N_3313,N_3167,N_3013);
nor U3314 (N_3314,N_3072,N_3139);
nor U3315 (N_3315,N_3102,N_3111);
xor U3316 (N_3316,N_3147,N_3152);
or U3317 (N_3317,N_3139,N_3193);
xnor U3318 (N_3318,N_3086,N_3100);
xor U3319 (N_3319,N_3004,N_3077);
nand U3320 (N_3320,N_3172,N_3053);
or U3321 (N_3321,N_3011,N_3052);
or U3322 (N_3322,N_3050,N_3165);
or U3323 (N_3323,N_3176,N_3043);
and U3324 (N_3324,N_3077,N_3038);
and U3325 (N_3325,N_3147,N_3196);
nand U3326 (N_3326,N_3095,N_3028);
or U3327 (N_3327,N_3008,N_3071);
xor U3328 (N_3328,N_3082,N_3030);
and U3329 (N_3329,N_3124,N_3144);
nor U3330 (N_3330,N_3133,N_3175);
or U3331 (N_3331,N_3127,N_3196);
nand U3332 (N_3332,N_3042,N_3160);
or U3333 (N_3333,N_3167,N_3017);
nand U3334 (N_3334,N_3136,N_3182);
nor U3335 (N_3335,N_3036,N_3128);
and U3336 (N_3336,N_3199,N_3100);
or U3337 (N_3337,N_3081,N_3160);
nand U3338 (N_3338,N_3097,N_3078);
nor U3339 (N_3339,N_3108,N_3197);
nor U3340 (N_3340,N_3016,N_3130);
or U3341 (N_3341,N_3073,N_3142);
and U3342 (N_3342,N_3047,N_3096);
nand U3343 (N_3343,N_3192,N_3154);
or U3344 (N_3344,N_3055,N_3100);
xor U3345 (N_3345,N_3015,N_3025);
xor U3346 (N_3346,N_3105,N_3144);
xnor U3347 (N_3347,N_3169,N_3153);
or U3348 (N_3348,N_3157,N_3128);
and U3349 (N_3349,N_3082,N_3096);
or U3350 (N_3350,N_3109,N_3016);
nor U3351 (N_3351,N_3138,N_3117);
and U3352 (N_3352,N_3179,N_3173);
nand U3353 (N_3353,N_3180,N_3195);
nand U3354 (N_3354,N_3111,N_3012);
xnor U3355 (N_3355,N_3182,N_3134);
xor U3356 (N_3356,N_3148,N_3172);
xor U3357 (N_3357,N_3149,N_3136);
nor U3358 (N_3358,N_3005,N_3013);
or U3359 (N_3359,N_3100,N_3040);
nor U3360 (N_3360,N_3014,N_3195);
xnor U3361 (N_3361,N_3196,N_3195);
and U3362 (N_3362,N_3035,N_3143);
nor U3363 (N_3363,N_3100,N_3169);
or U3364 (N_3364,N_3015,N_3036);
nand U3365 (N_3365,N_3031,N_3054);
xor U3366 (N_3366,N_3178,N_3028);
or U3367 (N_3367,N_3165,N_3177);
nor U3368 (N_3368,N_3167,N_3094);
and U3369 (N_3369,N_3071,N_3054);
nand U3370 (N_3370,N_3132,N_3122);
nand U3371 (N_3371,N_3081,N_3063);
nand U3372 (N_3372,N_3091,N_3101);
nand U3373 (N_3373,N_3165,N_3191);
or U3374 (N_3374,N_3047,N_3184);
or U3375 (N_3375,N_3082,N_3164);
xnor U3376 (N_3376,N_3111,N_3062);
nand U3377 (N_3377,N_3070,N_3080);
xnor U3378 (N_3378,N_3101,N_3044);
or U3379 (N_3379,N_3024,N_3125);
and U3380 (N_3380,N_3115,N_3062);
nand U3381 (N_3381,N_3069,N_3180);
nor U3382 (N_3382,N_3111,N_3088);
nor U3383 (N_3383,N_3151,N_3121);
xor U3384 (N_3384,N_3010,N_3075);
nand U3385 (N_3385,N_3068,N_3112);
nand U3386 (N_3386,N_3068,N_3177);
nand U3387 (N_3387,N_3113,N_3179);
or U3388 (N_3388,N_3122,N_3104);
nor U3389 (N_3389,N_3062,N_3172);
or U3390 (N_3390,N_3140,N_3024);
xnor U3391 (N_3391,N_3050,N_3123);
nor U3392 (N_3392,N_3136,N_3191);
nand U3393 (N_3393,N_3090,N_3174);
nand U3394 (N_3394,N_3038,N_3117);
xor U3395 (N_3395,N_3094,N_3015);
or U3396 (N_3396,N_3164,N_3076);
nor U3397 (N_3397,N_3172,N_3011);
nand U3398 (N_3398,N_3125,N_3140);
xor U3399 (N_3399,N_3158,N_3064);
nor U3400 (N_3400,N_3361,N_3359);
nand U3401 (N_3401,N_3207,N_3298);
nor U3402 (N_3402,N_3340,N_3210);
or U3403 (N_3403,N_3391,N_3259);
or U3404 (N_3404,N_3203,N_3239);
nor U3405 (N_3405,N_3341,N_3290);
or U3406 (N_3406,N_3240,N_3328);
xor U3407 (N_3407,N_3204,N_3333);
or U3408 (N_3408,N_3354,N_3363);
xor U3409 (N_3409,N_3294,N_3241);
xnor U3410 (N_3410,N_3323,N_3389);
xnor U3411 (N_3411,N_3338,N_3344);
nor U3412 (N_3412,N_3273,N_3233);
nor U3413 (N_3413,N_3309,N_3395);
and U3414 (N_3414,N_3254,N_3276);
nand U3415 (N_3415,N_3398,N_3322);
and U3416 (N_3416,N_3225,N_3329);
or U3417 (N_3417,N_3200,N_3311);
or U3418 (N_3418,N_3201,N_3305);
or U3419 (N_3419,N_3252,N_3383);
nor U3420 (N_3420,N_3263,N_3301);
and U3421 (N_3421,N_3205,N_3351);
nor U3422 (N_3422,N_3295,N_3373);
nor U3423 (N_3423,N_3218,N_3347);
xor U3424 (N_3424,N_3397,N_3399);
xor U3425 (N_3425,N_3260,N_3337);
xnor U3426 (N_3426,N_3326,N_3221);
or U3427 (N_3427,N_3206,N_3320);
nor U3428 (N_3428,N_3316,N_3242);
and U3429 (N_3429,N_3300,N_3375);
nor U3430 (N_3430,N_3331,N_3350);
nand U3431 (N_3431,N_3312,N_3307);
xor U3432 (N_3432,N_3289,N_3283);
nor U3433 (N_3433,N_3216,N_3377);
xor U3434 (N_3434,N_3271,N_3379);
nor U3435 (N_3435,N_3334,N_3346);
nand U3436 (N_3436,N_3388,N_3237);
nand U3437 (N_3437,N_3268,N_3266);
nor U3438 (N_3438,N_3274,N_3292);
nor U3439 (N_3439,N_3356,N_3386);
nor U3440 (N_3440,N_3297,N_3360);
nor U3441 (N_3441,N_3234,N_3372);
or U3442 (N_3442,N_3214,N_3330);
and U3443 (N_3443,N_3258,N_3327);
and U3444 (N_3444,N_3228,N_3317);
nor U3445 (N_3445,N_3264,N_3394);
or U3446 (N_3446,N_3279,N_3376);
nand U3447 (N_3447,N_3364,N_3308);
or U3448 (N_3448,N_3250,N_3267);
or U3449 (N_3449,N_3227,N_3282);
nand U3450 (N_3450,N_3261,N_3371);
and U3451 (N_3451,N_3212,N_3335);
nor U3452 (N_3452,N_3357,N_3362);
nand U3453 (N_3453,N_3224,N_3269);
xor U3454 (N_3454,N_3304,N_3285);
nor U3455 (N_3455,N_3382,N_3396);
xnor U3456 (N_3456,N_3253,N_3255);
or U3457 (N_3457,N_3265,N_3336);
nand U3458 (N_3458,N_3310,N_3229);
or U3459 (N_3459,N_3286,N_3348);
nor U3460 (N_3460,N_3215,N_3277);
nand U3461 (N_3461,N_3370,N_3293);
nand U3462 (N_3462,N_3246,N_3202);
and U3463 (N_3463,N_3366,N_3226);
and U3464 (N_3464,N_3219,N_3302);
or U3465 (N_3465,N_3324,N_3378);
nor U3466 (N_3466,N_3387,N_3236);
or U3467 (N_3467,N_3367,N_3392);
xnor U3468 (N_3468,N_3209,N_3358);
and U3469 (N_3469,N_3381,N_3345);
and U3470 (N_3470,N_3374,N_3270);
nor U3471 (N_3471,N_3208,N_3249);
xor U3472 (N_3472,N_3314,N_3256);
nand U3473 (N_3473,N_3245,N_3235);
xor U3474 (N_3474,N_3287,N_3291);
and U3475 (N_3475,N_3251,N_3281);
nor U3476 (N_3476,N_3393,N_3220);
nor U3477 (N_3477,N_3390,N_3262);
or U3478 (N_3478,N_3352,N_3243);
and U3479 (N_3479,N_3232,N_3222);
nand U3480 (N_3480,N_3248,N_3342);
or U3481 (N_3481,N_3321,N_3318);
and U3482 (N_3482,N_3280,N_3230);
xnor U3483 (N_3483,N_3339,N_3355);
and U3484 (N_3484,N_3325,N_3247);
and U3485 (N_3485,N_3257,N_3278);
or U3486 (N_3486,N_3272,N_3288);
or U3487 (N_3487,N_3319,N_3384);
nand U3488 (N_3488,N_3385,N_3343);
nand U3489 (N_3489,N_3349,N_3332);
xnor U3490 (N_3490,N_3238,N_3368);
or U3491 (N_3491,N_3217,N_3299);
nor U3492 (N_3492,N_3303,N_3296);
or U3493 (N_3493,N_3315,N_3380);
or U3494 (N_3494,N_3365,N_3211);
and U3495 (N_3495,N_3213,N_3313);
nand U3496 (N_3496,N_3306,N_3231);
or U3497 (N_3497,N_3275,N_3244);
xnor U3498 (N_3498,N_3369,N_3223);
and U3499 (N_3499,N_3353,N_3284);
nand U3500 (N_3500,N_3391,N_3365);
xnor U3501 (N_3501,N_3253,N_3355);
or U3502 (N_3502,N_3376,N_3360);
nand U3503 (N_3503,N_3270,N_3255);
nor U3504 (N_3504,N_3364,N_3349);
xnor U3505 (N_3505,N_3265,N_3213);
nor U3506 (N_3506,N_3369,N_3397);
or U3507 (N_3507,N_3293,N_3360);
or U3508 (N_3508,N_3319,N_3246);
and U3509 (N_3509,N_3232,N_3269);
xor U3510 (N_3510,N_3354,N_3219);
nand U3511 (N_3511,N_3217,N_3394);
xor U3512 (N_3512,N_3304,N_3214);
xnor U3513 (N_3513,N_3250,N_3207);
nor U3514 (N_3514,N_3356,N_3310);
or U3515 (N_3515,N_3334,N_3242);
nand U3516 (N_3516,N_3290,N_3239);
nand U3517 (N_3517,N_3248,N_3290);
nor U3518 (N_3518,N_3345,N_3272);
or U3519 (N_3519,N_3322,N_3200);
nand U3520 (N_3520,N_3246,N_3249);
and U3521 (N_3521,N_3284,N_3352);
nor U3522 (N_3522,N_3395,N_3396);
nand U3523 (N_3523,N_3279,N_3394);
nand U3524 (N_3524,N_3335,N_3239);
nand U3525 (N_3525,N_3365,N_3299);
xor U3526 (N_3526,N_3267,N_3215);
nor U3527 (N_3527,N_3219,N_3235);
xnor U3528 (N_3528,N_3372,N_3368);
and U3529 (N_3529,N_3277,N_3326);
and U3530 (N_3530,N_3368,N_3328);
nand U3531 (N_3531,N_3277,N_3271);
nand U3532 (N_3532,N_3217,N_3202);
xnor U3533 (N_3533,N_3364,N_3297);
or U3534 (N_3534,N_3349,N_3297);
nand U3535 (N_3535,N_3265,N_3326);
xnor U3536 (N_3536,N_3352,N_3316);
nand U3537 (N_3537,N_3281,N_3311);
xor U3538 (N_3538,N_3389,N_3355);
or U3539 (N_3539,N_3245,N_3225);
and U3540 (N_3540,N_3255,N_3306);
xnor U3541 (N_3541,N_3271,N_3321);
and U3542 (N_3542,N_3338,N_3361);
or U3543 (N_3543,N_3322,N_3363);
nor U3544 (N_3544,N_3233,N_3385);
nand U3545 (N_3545,N_3243,N_3321);
and U3546 (N_3546,N_3396,N_3227);
nor U3547 (N_3547,N_3223,N_3219);
nor U3548 (N_3548,N_3287,N_3380);
or U3549 (N_3549,N_3310,N_3218);
xnor U3550 (N_3550,N_3312,N_3360);
nand U3551 (N_3551,N_3345,N_3391);
nor U3552 (N_3552,N_3249,N_3367);
xnor U3553 (N_3553,N_3296,N_3387);
nand U3554 (N_3554,N_3206,N_3325);
nand U3555 (N_3555,N_3232,N_3352);
xnor U3556 (N_3556,N_3240,N_3302);
xor U3557 (N_3557,N_3257,N_3265);
or U3558 (N_3558,N_3248,N_3211);
or U3559 (N_3559,N_3230,N_3218);
and U3560 (N_3560,N_3227,N_3208);
xnor U3561 (N_3561,N_3357,N_3259);
nand U3562 (N_3562,N_3268,N_3386);
and U3563 (N_3563,N_3315,N_3276);
and U3564 (N_3564,N_3234,N_3255);
and U3565 (N_3565,N_3335,N_3331);
or U3566 (N_3566,N_3320,N_3213);
or U3567 (N_3567,N_3257,N_3366);
or U3568 (N_3568,N_3277,N_3384);
and U3569 (N_3569,N_3333,N_3390);
or U3570 (N_3570,N_3264,N_3325);
nor U3571 (N_3571,N_3354,N_3383);
nand U3572 (N_3572,N_3301,N_3368);
or U3573 (N_3573,N_3321,N_3315);
nor U3574 (N_3574,N_3283,N_3391);
and U3575 (N_3575,N_3366,N_3318);
and U3576 (N_3576,N_3323,N_3276);
or U3577 (N_3577,N_3247,N_3387);
and U3578 (N_3578,N_3260,N_3312);
xor U3579 (N_3579,N_3270,N_3370);
nor U3580 (N_3580,N_3362,N_3302);
and U3581 (N_3581,N_3268,N_3369);
or U3582 (N_3582,N_3376,N_3264);
nand U3583 (N_3583,N_3323,N_3291);
nor U3584 (N_3584,N_3204,N_3235);
nand U3585 (N_3585,N_3269,N_3206);
nand U3586 (N_3586,N_3399,N_3398);
nand U3587 (N_3587,N_3344,N_3221);
nor U3588 (N_3588,N_3229,N_3225);
xor U3589 (N_3589,N_3292,N_3278);
nor U3590 (N_3590,N_3359,N_3384);
nor U3591 (N_3591,N_3344,N_3386);
nor U3592 (N_3592,N_3368,N_3253);
nor U3593 (N_3593,N_3279,N_3392);
and U3594 (N_3594,N_3388,N_3291);
nor U3595 (N_3595,N_3255,N_3205);
nor U3596 (N_3596,N_3293,N_3237);
nor U3597 (N_3597,N_3369,N_3352);
nor U3598 (N_3598,N_3260,N_3394);
and U3599 (N_3599,N_3247,N_3350);
and U3600 (N_3600,N_3579,N_3495);
xor U3601 (N_3601,N_3438,N_3481);
xor U3602 (N_3602,N_3565,N_3427);
nand U3603 (N_3603,N_3412,N_3563);
nor U3604 (N_3604,N_3413,N_3526);
nand U3605 (N_3605,N_3516,N_3588);
and U3606 (N_3606,N_3483,N_3560);
nor U3607 (N_3607,N_3492,N_3587);
xor U3608 (N_3608,N_3514,N_3420);
or U3609 (N_3609,N_3536,N_3582);
and U3610 (N_3610,N_3559,N_3401);
nor U3611 (N_3611,N_3513,N_3480);
nand U3612 (N_3612,N_3425,N_3486);
and U3613 (N_3613,N_3593,N_3595);
nor U3614 (N_3614,N_3437,N_3494);
nand U3615 (N_3615,N_3447,N_3446);
nor U3616 (N_3616,N_3457,N_3550);
or U3617 (N_3617,N_3461,N_3555);
nor U3618 (N_3618,N_3432,N_3415);
nand U3619 (N_3619,N_3557,N_3539);
nor U3620 (N_3620,N_3535,N_3510);
nand U3621 (N_3621,N_3428,N_3414);
and U3622 (N_3622,N_3489,N_3574);
xor U3623 (N_3623,N_3479,N_3571);
nor U3624 (N_3624,N_3505,N_3577);
nand U3625 (N_3625,N_3470,N_3500);
and U3626 (N_3626,N_3402,N_3502);
and U3627 (N_3627,N_3512,N_3580);
or U3628 (N_3628,N_3429,N_3453);
nand U3629 (N_3629,N_3452,N_3544);
and U3630 (N_3630,N_3435,N_3581);
nand U3631 (N_3631,N_3454,N_3556);
nand U3632 (N_3632,N_3410,N_3542);
nand U3633 (N_3633,N_3467,N_3472);
or U3634 (N_3634,N_3543,N_3541);
nor U3635 (N_3635,N_3417,N_3578);
and U3636 (N_3636,N_3408,N_3553);
xor U3637 (N_3637,N_3545,N_3532);
or U3638 (N_3638,N_3418,N_3522);
nor U3639 (N_3639,N_3552,N_3473);
and U3640 (N_3640,N_3404,N_3439);
and U3641 (N_3641,N_3475,N_3496);
nand U3642 (N_3642,N_3490,N_3534);
or U3643 (N_3643,N_3478,N_3421);
nor U3644 (N_3644,N_3466,N_3476);
or U3645 (N_3645,N_3530,N_3455);
nand U3646 (N_3646,N_3589,N_3459);
or U3647 (N_3647,N_3409,N_3436);
or U3648 (N_3648,N_3527,N_3540);
and U3649 (N_3649,N_3568,N_3583);
nand U3650 (N_3650,N_3442,N_3596);
or U3651 (N_3651,N_3592,N_3594);
nand U3652 (N_3652,N_3597,N_3487);
xnor U3653 (N_3653,N_3562,N_3474);
nand U3654 (N_3654,N_3507,N_3493);
nand U3655 (N_3655,N_3573,N_3572);
nor U3656 (N_3656,N_3598,N_3508);
xor U3657 (N_3657,N_3570,N_3445);
nor U3658 (N_3658,N_3517,N_3504);
nor U3659 (N_3659,N_3525,N_3554);
nor U3660 (N_3660,N_3511,N_3558);
xor U3661 (N_3661,N_3529,N_3521);
and U3662 (N_3662,N_3569,N_3464);
and U3663 (N_3663,N_3419,N_3548);
or U3664 (N_3664,N_3518,N_3537);
xnor U3665 (N_3665,N_3422,N_3531);
nor U3666 (N_3666,N_3599,N_3460);
and U3667 (N_3667,N_3566,N_3591);
xor U3668 (N_3668,N_3440,N_3485);
and U3669 (N_3669,N_3528,N_3564);
or U3670 (N_3670,N_3411,N_3523);
xnor U3671 (N_3671,N_3405,N_3506);
and U3672 (N_3672,N_3444,N_3585);
xor U3673 (N_3673,N_3458,N_3456);
nand U3674 (N_3674,N_3590,N_3503);
nor U3675 (N_3675,N_3431,N_3482);
nor U3676 (N_3676,N_3491,N_3551);
nor U3677 (N_3677,N_3538,N_3451);
nand U3678 (N_3678,N_3499,N_3524);
nor U3679 (N_3679,N_3519,N_3484);
or U3680 (N_3680,N_3448,N_3498);
nor U3681 (N_3681,N_3434,N_3549);
xor U3682 (N_3682,N_3520,N_3416);
or U3683 (N_3683,N_3407,N_3477);
xor U3684 (N_3684,N_3509,N_3546);
nand U3685 (N_3685,N_3586,N_3400);
nor U3686 (N_3686,N_3441,N_3576);
xor U3687 (N_3687,N_3424,N_3468);
xnor U3688 (N_3688,N_3567,N_3465);
xnor U3689 (N_3689,N_3515,N_3406);
and U3690 (N_3690,N_3463,N_3433);
or U3691 (N_3691,N_3423,N_3497);
xnor U3692 (N_3692,N_3443,N_3547);
or U3693 (N_3693,N_3533,N_3471);
nand U3694 (N_3694,N_3584,N_3449);
or U3695 (N_3695,N_3430,N_3403);
nand U3696 (N_3696,N_3426,N_3469);
nor U3697 (N_3697,N_3501,N_3488);
and U3698 (N_3698,N_3561,N_3462);
or U3699 (N_3699,N_3450,N_3575);
nor U3700 (N_3700,N_3486,N_3499);
nor U3701 (N_3701,N_3561,N_3490);
or U3702 (N_3702,N_3442,N_3461);
and U3703 (N_3703,N_3595,N_3490);
xor U3704 (N_3704,N_3459,N_3465);
nor U3705 (N_3705,N_3411,N_3586);
xor U3706 (N_3706,N_3578,N_3451);
nand U3707 (N_3707,N_3449,N_3466);
and U3708 (N_3708,N_3579,N_3429);
nor U3709 (N_3709,N_3402,N_3556);
or U3710 (N_3710,N_3594,N_3568);
nor U3711 (N_3711,N_3477,N_3497);
and U3712 (N_3712,N_3483,N_3544);
xor U3713 (N_3713,N_3502,N_3482);
nand U3714 (N_3714,N_3474,N_3592);
nand U3715 (N_3715,N_3400,N_3595);
nor U3716 (N_3716,N_3505,N_3538);
xor U3717 (N_3717,N_3454,N_3567);
and U3718 (N_3718,N_3526,N_3501);
nor U3719 (N_3719,N_3406,N_3498);
nand U3720 (N_3720,N_3596,N_3487);
or U3721 (N_3721,N_3421,N_3504);
nor U3722 (N_3722,N_3492,N_3441);
xnor U3723 (N_3723,N_3470,N_3514);
or U3724 (N_3724,N_3513,N_3496);
and U3725 (N_3725,N_3542,N_3429);
xor U3726 (N_3726,N_3413,N_3580);
xor U3727 (N_3727,N_3552,N_3451);
xnor U3728 (N_3728,N_3456,N_3577);
nor U3729 (N_3729,N_3472,N_3500);
and U3730 (N_3730,N_3405,N_3568);
or U3731 (N_3731,N_3584,N_3523);
nor U3732 (N_3732,N_3426,N_3548);
nor U3733 (N_3733,N_3491,N_3592);
nand U3734 (N_3734,N_3448,N_3519);
nor U3735 (N_3735,N_3437,N_3429);
and U3736 (N_3736,N_3574,N_3509);
xnor U3737 (N_3737,N_3573,N_3531);
xor U3738 (N_3738,N_3518,N_3530);
or U3739 (N_3739,N_3514,N_3462);
xor U3740 (N_3740,N_3434,N_3475);
nand U3741 (N_3741,N_3460,N_3554);
xnor U3742 (N_3742,N_3578,N_3487);
nor U3743 (N_3743,N_3502,N_3550);
nand U3744 (N_3744,N_3595,N_3594);
nand U3745 (N_3745,N_3415,N_3527);
nand U3746 (N_3746,N_3494,N_3479);
and U3747 (N_3747,N_3565,N_3417);
nand U3748 (N_3748,N_3487,N_3570);
and U3749 (N_3749,N_3462,N_3589);
nand U3750 (N_3750,N_3542,N_3556);
nor U3751 (N_3751,N_3419,N_3562);
nor U3752 (N_3752,N_3438,N_3421);
and U3753 (N_3753,N_3530,N_3486);
nand U3754 (N_3754,N_3458,N_3487);
and U3755 (N_3755,N_3444,N_3519);
and U3756 (N_3756,N_3404,N_3525);
nand U3757 (N_3757,N_3466,N_3448);
xor U3758 (N_3758,N_3558,N_3523);
nor U3759 (N_3759,N_3526,N_3505);
and U3760 (N_3760,N_3542,N_3529);
nor U3761 (N_3761,N_3426,N_3574);
xor U3762 (N_3762,N_3559,N_3426);
nor U3763 (N_3763,N_3525,N_3578);
xnor U3764 (N_3764,N_3543,N_3560);
and U3765 (N_3765,N_3426,N_3576);
or U3766 (N_3766,N_3544,N_3560);
and U3767 (N_3767,N_3472,N_3411);
xnor U3768 (N_3768,N_3528,N_3541);
or U3769 (N_3769,N_3422,N_3541);
nor U3770 (N_3770,N_3551,N_3535);
nand U3771 (N_3771,N_3529,N_3493);
xor U3772 (N_3772,N_3414,N_3455);
or U3773 (N_3773,N_3401,N_3544);
xnor U3774 (N_3774,N_3533,N_3404);
nor U3775 (N_3775,N_3431,N_3532);
nand U3776 (N_3776,N_3457,N_3402);
and U3777 (N_3777,N_3545,N_3555);
nor U3778 (N_3778,N_3595,N_3508);
nand U3779 (N_3779,N_3518,N_3553);
xnor U3780 (N_3780,N_3584,N_3597);
or U3781 (N_3781,N_3506,N_3401);
nor U3782 (N_3782,N_3527,N_3472);
nand U3783 (N_3783,N_3559,N_3472);
nand U3784 (N_3784,N_3478,N_3476);
or U3785 (N_3785,N_3435,N_3501);
nor U3786 (N_3786,N_3583,N_3507);
nor U3787 (N_3787,N_3553,N_3452);
or U3788 (N_3788,N_3555,N_3490);
xor U3789 (N_3789,N_3550,N_3416);
xor U3790 (N_3790,N_3461,N_3436);
nor U3791 (N_3791,N_3406,N_3417);
and U3792 (N_3792,N_3535,N_3413);
or U3793 (N_3793,N_3423,N_3502);
and U3794 (N_3794,N_3535,N_3409);
xor U3795 (N_3795,N_3449,N_3594);
xnor U3796 (N_3796,N_3453,N_3448);
or U3797 (N_3797,N_3448,N_3445);
xor U3798 (N_3798,N_3545,N_3497);
nand U3799 (N_3799,N_3552,N_3488);
or U3800 (N_3800,N_3670,N_3786);
nand U3801 (N_3801,N_3698,N_3669);
or U3802 (N_3802,N_3650,N_3609);
and U3803 (N_3803,N_3715,N_3766);
or U3804 (N_3804,N_3796,N_3620);
nand U3805 (N_3805,N_3740,N_3684);
and U3806 (N_3806,N_3783,N_3743);
or U3807 (N_3807,N_3687,N_3606);
nor U3808 (N_3808,N_3746,N_3759);
or U3809 (N_3809,N_3763,N_3726);
and U3810 (N_3810,N_3700,N_3711);
and U3811 (N_3811,N_3721,N_3776);
or U3812 (N_3812,N_3718,N_3720);
nand U3813 (N_3813,N_3768,N_3713);
and U3814 (N_3814,N_3625,N_3661);
and U3815 (N_3815,N_3790,N_3771);
or U3816 (N_3816,N_3723,N_3691);
nor U3817 (N_3817,N_3660,N_3689);
xnor U3818 (N_3818,N_3634,N_3794);
or U3819 (N_3819,N_3742,N_3610);
nor U3820 (N_3820,N_3638,N_3685);
or U3821 (N_3821,N_3765,N_3712);
and U3822 (N_3822,N_3795,N_3734);
nor U3823 (N_3823,N_3633,N_3753);
nor U3824 (N_3824,N_3652,N_3654);
nor U3825 (N_3825,N_3719,N_3642);
xor U3826 (N_3826,N_3714,N_3631);
nand U3827 (N_3827,N_3655,N_3601);
nand U3828 (N_3828,N_3667,N_3764);
xnor U3829 (N_3829,N_3651,N_3605);
nand U3830 (N_3830,N_3716,N_3617);
or U3831 (N_3831,N_3751,N_3775);
and U3832 (N_3832,N_3664,N_3778);
or U3833 (N_3833,N_3671,N_3704);
xnor U3834 (N_3834,N_3643,N_3663);
nand U3835 (N_3835,N_3741,N_3695);
xnor U3836 (N_3836,N_3611,N_3692);
or U3837 (N_3837,N_3614,N_3729);
xnor U3838 (N_3838,N_3750,N_3662);
and U3839 (N_3839,N_3693,N_3708);
xnor U3840 (N_3840,N_3773,N_3717);
and U3841 (N_3841,N_3789,N_3780);
nand U3842 (N_3842,N_3735,N_3672);
xnor U3843 (N_3843,N_3736,N_3756);
and U3844 (N_3844,N_3649,N_3732);
nor U3845 (N_3845,N_3739,N_3688);
xor U3846 (N_3846,N_3637,N_3608);
and U3847 (N_3847,N_3730,N_3607);
and U3848 (N_3848,N_3710,N_3630);
xnor U3849 (N_3849,N_3793,N_3602);
or U3850 (N_3850,N_3624,N_3781);
or U3851 (N_3851,N_3666,N_3603);
xor U3852 (N_3852,N_3622,N_3762);
xnor U3853 (N_3853,N_3797,N_3699);
and U3854 (N_3854,N_3644,N_3757);
xor U3855 (N_3855,N_3658,N_3646);
and U3856 (N_3856,N_3745,N_3653);
and U3857 (N_3857,N_3784,N_3747);
nor U3858 (N_3858,N_3779,N_3774);
nor U3859 (N_3859,N_3792,N_3618);
xor U3860 (N_3860,N_3705,N_3744);
xnor U3861 (N_3861,N_3760,N_3683);
or U3862 (N_3862,N_3682,N_3767);
or U3863 (N_3863,N_3709,N_3727);
xnor U3864 (N_3864,N_3673,N_3738);
xnor U3865 (N_3865,N_3694,N_3659);
nor U3866 (N_3866,N_3640,N_3702);
and U3867 (N_3867,N_3675,N_3725);
nor U3868 (N_3868,N_3706,N_3621);
nor U3869 (N_3869,N_3724,N_3681);
xor U3870 (N_3870,N_3613,N_3798);
nand U3871 (N_3871,N_3761,N_3772);
nor U3872 (N_3872,N_3686,N_3641);
or U3873 (N_3873,N_3676,N_3600);
and U3874 (N_3874,N_3707,N_3616);
nand U3875 (N_3875,N_3748,N_3782);
xor U3876 (N_3876,N_3701,N_3680);
nand U3877 (N_3877,N_3769,N_3656);
nor U3878 (N_3878,N_3787,N_3612);
and U3879 (N_3879,N_3647,N_3677);
nand U3880 (N_3880,N_3785,N_3696);
and U3881 (N_3881,N_3752,N_3635);
nor U3882 (N_3882,N_3639,N_3628);
or U3883 (N_3883,N_3678,N_3788);
xnor U3884 (N_3884,N_3777,N_3636);
nor U3885 (N_3885,N_3754,N_3619);
and U3886 (N_3886,N_3648,N_3674);
xor U3887 (N_3887,N_3703,N_3679);
and U3888 (N_3888,N_3791,N_3627);
or U3889 (N_3889,N_3668,N_3755);
nand U3890 (N_3890,N_3731,N_3623);
or U3891 (N_3891,N_3657,N_3737);
and U3892 (N_3892,N_3604,N_3758);
and U3893 (N_3893,N_3722,N_3728);
nand U3894 (N_3894,N_3615,N_3799);
or U3895 (N_3895,N_3749,N_3690);
nor U3896 (N_3896,N_3632,N_3665);
or U3897 (N_3897,N_3645,N_3626);
and U3898 (N_3898,N_3697,N_3629);
nand U3899 (N_3899,N_3770,N_3733);
xnor U3900 (N_3900,N_3680,N_3638);
or U3901 (N_3901,N_3698,N_3649);
or U3902 (N_3902,N_3652,N_3680);
nand U3903 (N_3903,N_3612,N_3781);
xnor U3904 (N_3904,N_3673,N_3699);
nor U3905 (N_3905,N_3665,N_3605);
and U3906 (N_3906,N_3658,N_3731);
or U3907 (N_3907,N_3747,N_3759);
nand U3908 (N_3908,N_3616,N_3629);
nand U3909 (N_3909,N_3707,N_3761);
xnor U3910 (N_3910,N_3784,N_3764);
nor U3911 (N_3911,N_3689,N_3656);
nand U3912 (N_3912,N_3786,N_3605);
or U3913 (N_3913,N_3680,N_3670);
nor U3914 (N_3914,N_3709,N_3759);
nor U3915 (N_3915,N_3756,N_3776);
xnor U3916 (N_3916,N_3616,N_3665);
or U3917 (N_3917,N_3626,N_3660);
xnor U3918 (N_3918,N_3669,N_3770);
nor U3919 (N_3919,N_3763,N_3655);
xnor U3920 (N_3920,N_3773,N_3667);
nor U3921 (N_3921,N_3707,N_3711);
xor U3922 (N_3922,N_3619,N_3609);
xor U3923 (N_3923,N_3661,N_3763);
nor U3924 (N_3924,N_3618,N_3658);
and U3925 (N_3925,N_3706,N_3746);
nor U3926 (N_3926,N_3746,N_3654);
xnor U3927 (N_3927,N_3728,N_3662);
nand U3928 (N_3928,N_3628,N_3675);
and U3929 (N_3929,N_3697,N_3603);
or U3930 (N_3930,N_3758,N_3654);
and U3931 (N_3931,N_3785,N_3771);
and U3932 (N_3932,N_3734,N_3654);
and U3933 (N_3933,N_3697,N_3776);
and U3934 (N_3934,N_3774,N_3699);
and U3935 (N_3935,N_3757,N_3698);
or U3936 (N_3936,N_3610,N_3746);
or U3937 (N_3937,N_3625,N_3677);
and U3938 (N_3938,N_3649,N_3674);
nand U3939 (N_3939,N_3643,N_3604);
and U3940 (N_3940,N_3670,N_3649);
nor U3941 (N_3941,N_3664,N_3760);
and U3942 (N_3942,N_3605,N_3626);
nand U3943 (N_3943,N_3724,N_3713);
or U3944 (N_3944,N_3795,N_3768);
nor U3945 (N_3945,N_3638,N_3631);
xor U3946 (N_3946,N_3717,N_3676);
and U3947 (N_3947,N_3626,N_3602);
nand U3948 (N_3948,N_3789,N_3720);
nand U3949 (N_3949,N_3635,N_3670);
or U3950 (N_3950,N_3783,N_3780);
or U3951 (N_3951,N_3619,N_3677);
or U3952 (N_3952,N_3688,N_3641);
xor U3953 (N_3953,N_3669,N_3690);
xnor U3954 (N_3954,N_3628,N_3652);
xor U3955 (N_3955,N_3780,N_3608);
nand U3956 (N_3956,N_3749,N_3617);
and U3957 (N_3957,N_3765,N_3764);
nand U3958 (N_3958,N_3687,N_3679);
xnor U3959 (N_3959,N_3779,N_3764);
and U3960 (N_3960,N_3736,N_3676);
nor U3961 (N_3961,N_3741,N_3677);
nor U3962 (N_3962,N_3772,N_3634);
nor U3963 (N_3963,N_3723,N_3756);
or U3964 (N_3964,N_3638,N_3646);
and U3965 (N_3965,N_3758,N_3606);
and U3966 (N_3966,N_3783,N_3669);
nor U3967 (N_3967,N_3723,N_3683);
or U3968 (N_3968,N_3768,N_3764);
and U3969 (N_3969,N_3726,N_3752);
or U3970 (N_3970,N_3758,N_3714);
nor U3971 (N_3971,N_3643,N_3690);
and U3972 (N_3972,N_3625,N_3775);
and U3973 (N_3973,N_3743,N_3694);
nand U3974 (N_3974,N_3786,N_3613);
or U3975 (N_3975,N_3604,N_3616);
xnor U3976 (N_3976,N_3647,N_3651);
nor U3977 (N_3977,N_3604,N_3659);
nand U3978 (N_3978,N_3768,N_3659);
nor U3979 (N_3979,N_3728,N_3712);
and U3980 (N_3980,N_3630,N_3733);
nand U3981 (N_3981,N_3715,N_3797);
or U3982 (N_3982,N_3604,N_3783);
nor U3983 (N_3983,N_3681,N_3640);
nor U3984 (N_3984,N_3730,N_3681);
nor U3985 (N_3985,N_3716,N_3690);
nand U3986 (N_3986,N_3745,N_3694);
and U3987 (N_3987,N_3785,N_3687);
nand U3988 (N_3988,N_3666,N_3776);
and U3989 (N_3989,N_3782,N_3787);
xor U3990 (N_3990,N_3740,N_3607);
xnor U3991 (N_3991,N_3717,N_3685);
nand U3992 (N_3992,N_3601,N_3617);
nand U3993 (N_3993,N_3610,N_3716);
and U3994 (N_3994,N_3647,N_3654);
nand U3995 (N_3995,N_3642,N_3631);
xor U3996 (N_3996,N_3781,N_3695);
xor U3997 (N_3997,N_3674,N_3708);
or U3998 (N_3998,N_3652,N_3739);
nor U3999 (N_3999,N_3710,N_3680);
nand U4000 (N_4000,N_3828,N_3816);
nand U4001 (N_4001,N_3845,N_3973);
nor U4002 (N_4002,N_3966,N_3930);
nor U4003 (N_4003,N_3810,N_3921);
and U4004 (N_4004,N_3942,N_3827);
nor U4005 (N_4005,N_3913,N_3922);
nor U4006 (N_4006,N_3887,N_3898);
xor U4007 (N_4007,N_3931,N_3969);
or U4008 (N_4008,N_3976,N_3809);
nand U4009 (N_4009,N_3951,N_3961);
nand U4010 (N_4010,N_3822,N_3927);
nand U4011 (N_4011,N_3992,N_3874);
and U4012 (N_4012,N_3863,N_3853);
nor U4013 (N_4013,N_3889,N_3938);
nand U4014 (N_4014,N_3873,N_3933);
or U4015 (N_4015,N_3999,N_3955);
and U4016 (N_4016,N_3974,N_3944);
nand U4017 (N_4017,N_3843,N_3858);
xor U4018 (N_4018,N_3917,N_3841);
xor U4019 (N_4019,N_3980,N_3947);
or U4020 (N_4020,N_3881,N_3901);
xnor U4021 (N_4021,N_3914,N_3803);
or U4022 (N_4022,N_3814,N_3997);
and U4023 (N_4023,N_3893,N_3865);
and U4024 (N_4024,N_3846,N_3824);
and U4025 (N_4025,N_3840,N_3948);
nor U4026 (N_4026,N_3993,N_3868);
and U4027 (N_4027,N_3842,N_3872);
and U4028 (N_4028,N_3855,N_3869);
or U4029 (N_4029,N_3970,N_3954);
or U4030 (N_4030,N_3959,N_3856);
and U4031 (N_4031,N_3844,N_3852);
nor U4032 (N_4032,N_3821,N_3916);
or U4033 (N_4033,N_3936,N_3885);
and U4034 (N_4034,N_3964,N_3836);
nor U4035 (N_4035,N_3823,N_3994);
and U4036 (N_4036,N_3949,N_3886);
xnor U4037 (N_4037,N_3943,N_3820);
nand U4038 (N_4038,N_3866,N_3965);
or U4039 (N_4039,N_3903,N_3906);
or U4040 (N_4040,N_3802,N_3945);
nand U4041 (N_4041,N_3982,N_3819);
or U4042 (N_4042,N_3900,N_3875);
and U4043 (N_4043,N_3818,N_3847);
nand U4044 (N_4044,N_3864,N_3977);
nor U4045 (N_4045,N_3862,N_3888);
xor U4046 (N_4046,N_3963,N_3876);
or U4047 (N_4047,N_3939,N_3952);
xor U4048 (N_4048,N_3908,N_3984);
and U4049 (N_4049,N_3801,N_3915);
nand U4050 (N_4050,N_3928,N_3879);
nand U4051 (N_4051,N_3925,N_3812);
and U4052 (N_4052,N_3892,N_3849);
xor U4053 (N_4053,N_3910,N_3912);
and U4054 (N_4054,N_3920,N_3957);
nor U4055 (N_4055,N_3904,N_3870);
xnor U4056 (N_4056,N_3941,N_3923);
xnor U4057 (N_4057,N_3817,N_3986);
xor U4058 (N_4058,N_3815,N_3946);
or U4059 (N_4059,N_3839,N_3830);
xnor U4060 (N_4060,N_3907,N_3940);
xor U4061 (N_4061,N_3890,N_3831);
nand U4062 (N_4062,N_3990,N_3806);
xor U4063 (N_4063,N_3985,N_3891);
and U4064 (N_4064,N_3899,N_3978);
nor U4065 (N_4065,N_3835,N_3979);
or U4066 (N_4066,N_3884,N_3919);
and U4067 (N_4067,N_3850,N_3860);
or U4068 (N_4068,N_3861,N_3929);
nor U4069 (N_4069,N_3958,N_3804);
and U4070 (N_4070,N_3848,N_3924);
and U4071 (N_4071,N_3867,N_3934);
nand U4072 (N_4072,N_3897,N_3805);
xnor U4073 (N_4073,N_3857,N_3800);
nand U4074 (N_4074,N_3981,N_3877);
xor U4075 (N_4075,N_3972,N_3878);
nor U4076 (N_4076,N_3960,N_3975);
nor U4077 (N_4077,N_3995,N_3956);
nor U4078 (N_4078,N_3926,N_3950);
or U4079 (N_4079,N_3883,N_3988);
xnor U4080 (N_4080,N_3825,N_3896);
and U4081 (N_4081,N_3854,N_3987);
nor U4082 (N_4082,N_3971,N_3895);
nand U4083 (N_4083,N_3962,N_3834);
or U4084 (N_4084,N_3808,N_3813);
or U4085 (N_4085,N_3935,N_3880);
nand U4086 (N_4086,N_3932,N_3911);
or U4087 (N_4087,N_3851,N_3953);
or U4088 (N_4088,N_3937,N_3905);
and U4089 (N_4089,N_3859,N_3998);
xnor U4090 (N_4090,N_3833,N_3968);
or U4091 (N_4091,N_3837,N_3996);
xnor U4092 (N_4092,N_3807,N_3909);
and U4093 (N_4093,N_3871,N_3826);
and U4094 (N_4094,N_3838,N_3832);
xnor U4095 (N_4095,N_3882,N_3918);
or U4096 (N_4096,N_3894,N_3902);
and U4097 (N_4097,N_3811,N_3991);
and U4098 (N_4098,N_3989,N_3983);
nor U4099 (N_4099,N_3829,N_3967);
nor U4100 (N_4100,N_3831,N_3912);
and U4101 (N_4101,N_3832,N_3928);
or U4102 (N_4102,N_3982,N_3980);
nand U4103 (N_4103,N_3865,N_3889);
or U4104 (N_4104,N_3846,N_3902);
nor U4105 (N_4105,N_3888,N_3982);
xnor U4106 (N_4106,N_3802,N_3993);
xor U4107 (N_4107,N_3994,N_3920);
xor U4108 (N_4108,N_3905,N_3834);
nor U4109 (N_4109,N_3897,N_3824);
and U4110 (N_4110,N_3886,N_3831);
or U4111 (N_4111,N_3803,N_3995);
and U4112 (N_4112,N_3847,N_3887);
xnor U4113 (N_4113,N_3825,N_3997);
and U4114 (N_4114,N_3894,N_3881);
or U4115 (N_4115,N_3879,N_3837);
xnor U4116 (N_4116,N_3865,N_3998);
nor U4117 (N_4117,N_3941,N_3907);
xnor U4118 (N_4118,N_3852,N_3924);
nand U4119 (N_4119,N_3889,N_3894);
nor U4120 (N_4120,N_3877,N_3857);
nand U4121 (N_4121,N_3944,N_3843);
or U4122 (N_4122,N_3962,N_3803);
and U4123 (N_4123,N_3978,N_3828);
and U4124 (N_4124,N_3953,N_3875);
xnor U4125 (N_4125,N_3923,N_3993);
nand U4126 (N_4126,N_3996,N_3810);
xnor U4127 (N_4127,N_3969,N_3872);
and U4128 (N_4128,N_3904,N_3959);
xor U4129 (N_4129,N_3905,N_3970);
and U4130 (N_4130,N_3929,N_3850);
xnor U4131 (N_4131,N_3990,N_3837);
nand U4132 (N_4132,N_3827,N_3869);
nor U4133 (N_4133,N_3943,N_3870);
or U4134 (N_4134,N_3930,N_3929);
nor U4135 (N_4135,N_3908,N_3871);
or U4136 (N_4136,N_3944,N_3915);
or U4137 (N_4137,N_3985,N_3941);
and U4138 (N_4138,N_3800,N_3981);
or U4139 (N_4139,N_3946,N_3878);
or U4140 (N_4140,N_3954,N_3860);
nand U4141 (N_4141,N_3817,N_3941);
or U4142 (N_4142,N_3886,N_3944);
nor U4143 (N_4143,N_3852,N_3818);
xnor U4144 (N_4144,N_3978,N_3854);
xor U4145 (N_4145,N_3833,N_3895);
nor U4146 (N_4146,N_3957,N_3997);
nand U4147 (N_4147,N_3957,N_3876);
xor U4148 (N_4148,N_3877,N_3929);
nand U4149 (N_4149,N_3932,N_3829);
and U4150 (N_4150,N_3956,N_3917);
or U4151 (N_4151,N_3935,N_3903);
nor U4152 (N_4152,N_3837,N_3843);
nor U4153 (N_4153,N_3928,N_3986);
nand U4154 (N_4154,N_3968,N_3880);
nand U4155 (N_4155,N_3931,N_3995);
xnor U4156 (N_4156,N_3896,N_3921);
and U4157 (N_4157,N_3833,N_3969);
nor U4158 (N_4158,N_3819,N_3995);
or U4159 (N_4159,N_3901,N_3904);
nor U4160 (N_4160,N_3930,N_3811);
or U4161 (N_4161,N_3923,N_3956);
nand U4162 (N_4162,N_3839,N_3926);
nor U4163 (N_4163,N_3800,N_3975);
or U4164 (N_4164,N_3862,N_3986);
nand U4165 (N_4165,N_3853,N_3961);
nor U4166 (N_4166,N_3885,N_3932);
xnor U4167 (N_4167,N_3857,N_3811);
or U4168 (N_4168,N_3949,N_3806);
xor U4169 (N_4169,N_3801,N_3892);
nand U4170 (N_4170,N_3844,N_3887);
or U4171 (N_4171,N_3857,N_3981);
nor U4172 (N_4172,N_3975,N_3953);
nor U4173 (N_4173,N_3871,N_3802);
nand U4174 (N_4174,N_3870,N_3967);
xor U4175 (N_4175,N_3800,N_3863);
nor U4176 (N_4176,N_3850,N_3971);
and U4177 (N_4177,N_3832,N_3923);
nand U4178 (N_4178,N_3840,N_3832);
nand U4179 (N_4179,N_3816,N_3994);
and U4180 (N_4180,N_3964,N_3992);
xor U4181 (N_4181,N_3863,N_3807);
nor U4182 (N_4182,N_3850,N_3994);
nor U4183 (N_4183,N_3867,N_3869);
nor U4184 (N_4184,N_3873,N_3810);
or U4185 (N_4185,N_3938,N_3840);
and U4186 (N_4186,N_3883,N_3877);
nand U4187 (N_4187,N_3965,N_3952);
or U4188 (N_4188,N_3881,N_3884);
nand U4189 (N_4189,N_3976,N_3975);
and U4190 (N_4190,N_3818,N_3998);
or U4191 (N_4191,N_3826,N_3810);
nor U4192 (N_4192,N_3984,N_3996);
xnor U4193 (N_4193,N_3803,N_3838);
or U4194 (N_4194,N_3934,N_3857);
or U4195 (N_4195,N_3816,N_3969);
or U4196 (N_4196,N_3885,N_3870);
xnor U4197 (N_4197,N_3927,N_3902);
nor U4198 (N_4198,N_3989,N_3878);
or U4199 (N_4199,N_3942,N_3876);
xnor U4200 (N_4200,N_4020,N_4152);
and U4201 (N_4201,N_4057,N_4153);
nand U4202 (N_4202,N_4055,N_4188);
nand U4203 (N_4203,N_4131,N_4166);
nand U4204 (N_4204,N_4069,N_4134);
and U4205 (N_4205,N_4129,N_4087);
nand U4206 (N_4206,N_4024,N_4080);
and U4207 (N_4207,N_4076,N_4155);
nor U4208 (N_4208,N_4074,N_4127);
nor U4209 (N_4209,N_4092,N_4165);
nand U4210 (N_4210,N_4082,N_4084);
or U4211 (N_4211,N_4041,N_4039);
xnor U4212 (N_4212,N_4177,N_4193);
or U4213 (N_4213,N_4123,N_4164);
xor U4214 (N_4214,N_4098,N_4112);
xnor U4215 (N_4215,N_4006,N_4178);
or U4216 (N_4216,N_4173,N_4023);
nand U4217 (N_4217,N_4190,N_4064);
xnor U4218 (N_4218,N_4027,N_4086);
and U4219 (N_4219,N_4099,N_4137);
and U4220 (N_4220,N_4182,N_4135);
xnor U4221 (N_4221,N_4090,N_4119);
nor U4222 (N_4222,N_4097,N_4083);
nor U4223 (N_4223,N_4011,N_4056);
and U4224 (N_4224,N_4003,N_4026);
and U4225 (N_4225,N_4044,N_4031);
nor U4226 (N_4226,N_4174,N_4068);
nand U4227 (N_4227,N_4028,N_4051);
and U4228 (N_4228,N_4101,N_4015);
and U4229 (N_4229,N_4091,N_4185);
and U4230 (N_4230,N_4000,N_4199);
nand U4231 (N_4231,N_4106,N_4070);
or U4232 (N_4232,N_4150,N_4159);
or U4233 (N_4233,N_4008,N_4018);
and U4234 (N_4234,N_4021,N_4128);
nand U4235 (N_4235,N_4133,N_4078);
xor U4236 (N_4236,N_4001,N_4117);
or U4237 (N_4237,N_4160,N_4170);
nor U4238 (N_4238,N_4060,N_4025);
and U4239 (N_4239,N_4010,N_4172);
or U4240 (N_4240,N_4122,N_4197);
or U4241 (N_4241,N_4143,N_4047);
xor U4242 (N_4242,N_4118,N_4045);
nor U4243 (N_4243,N_4065,N_4141);
nand U4244 (N_4244,N_4120,N_4162);
or U4245 (N_4245,N_4085,N_4105);
nand U4246 (N_4246,N_4077,N_4154);
or U4247 (N_4247,N_4111,N_4062);
and U4248 (N_4248,N_4108,N_4121);
xnor U4249 (N_4249,N_4196,N_4093);
nand U4250 (N_4250,N_4139,N_4017);
xor U4251 (N_4251,N_4138,N_4046);
xnor U4252 (N_4252,N_4163,N_4102);
nor U4253 (N_4253,N_4184,N_4029);
or U4254 (N_4254,N_4148,N_4038);
or U4255 (N_4255,N_4096,N_4187);
nand U4256 (N_4256,N_4124,N_4050);
nor U4257 (N_4257,N_4169,N_4140);
nand U4258 (N_4258,N_4073,N_4095);
nor U4259 (N_4259,N_4114,N_4180);
and U4260 (N_4260,N_4194,N_4004);
and U4261 (N_4261,N_4103,N_4126);
or U4262 (N_4262,N_4022,N_4158);
xnor U4263 (N_4263,N_4116,N_4066);
nand U4264 (N_4264,N_4110,N_4081);
or U4265 (N_4265,N_4071,N_4067);
and U4266 (N_4266,N_4186,N_4002);
and U4267 (N_4267,N_4104,N_4013);
and U4268 (N_4268,N_4168,N_4100);
nor U4269 (N_4269,N_4144,N_4130);
nor U4270 (N_4270,N_4035,N_4037);
and U4271 (N_4271,N_4175,N_4113);
or U4272 (N_4272,N_4125,N_4075);
nor U4273 (N_4273,N_4192,N_4043);
xor U4274 (N_4274,N_4179,N_4072);
nand U4275 (N_4275,N_4171,N_4014);
and U4276 (N_4276,N_4048,N_4058);
xnor U4277 (N_4277,N_4115,N_4191);
nand U4278 (N_4278,N_4157,N_4107);
nand U4279 (N_4279,N_4052,N_4142);
or U4280 (N_4280,N_4009,N_4030);
or U4281 (N_4281,N_4167,N_4146);
or U4282 (N_4282,N_4181,N_4063);
and U4283 (N_4283,N_4049,N_4079);
and U4284 (N_4284,N_4033,N_4088);
nor U4285 (N_4285,N_4042,N_4094);
nand U4286 (N_4286,N_4147,N_4151);
or U4287 (N_4287,N_4195,N_4189);
nand U4288 (N_4288,N_4149,N_4034);
nand U4289 (N_4289,N_4183,N_4053);
nor U4290 (N_4290,N_4007,N_4089);
or U4291 (N_4291,N_4019,N_4156);
xnor U4292 (N_4292,N_4136,N_4145);
xor U4293 (N_4293,N_4198,N_4012);
or U4294 (N_4294,N_4161,N_4032);
and U4295 (N_4295,N_4040,N_4005);
or U4296 (N_4296,N_4054,N_4109);
nand U4297 (N_4297,N_4176,N_4059);
or U4298 (N_4298,N_4132,N_4036);
and U4299 (N_4299,N_4061,N_4016);
and U4300 (N_4300,N_4183,N_4125);
nor U4301 (N_4301,N_4150,N_4122);
nand U4302 (N_4302,N_4036,N_4068);
nor U4303 (N_4303,N_4163,N_4080);
xor U4304 (N_4304,N_4102,N_4061);
nand U4305 (N_4305,N_4155,N_4121);
xnor U4306 (N_4306,N_4004,N_4002);
nand U4307 (N_4307,N_4087,N_4067);
xnor U4308 (N_4308,N_4018,N_4119);
nand U4309 (N_4309,N_4149,N_4170);
nand U4310 (N_4310,N_4040,N_4105);
nand U4311 (N_4311,N_4123,N_4087);
nor U4312 (N_4312,N_4052,N_4169);
nand U4313 (N_4313,N_4147,N_4114);
nor U4314 (N_4314,N_4160,N_4059);
nor U4315 (N_4315,N_4017,N_4130);
nor U4316 (N_4316,N_4153,N_4005);
and U4317 (N_4317,N_4006,N_4091);
xnor U4318 (N_4318,N_4030,N_4059);
nand U4319 (N_4319,N_4112,N_4006);
nor U4320 (N_4320,N_4109,N_4198);
or U4321 (N_4321,N_4066,N_4150);
and U4322 (N_4322,N_4022,N_4128);
and U4323 (N_4323,N_4133,N_4064);
xor U4324 (N_4324,N_4123,N_4069);
xnor U4325 (N_4325,N_4009,N_4193);
nor U4326 (N_4326,N_4044,N_4133);
xor U4327 (N_4327,N_4130,N_4066);
and U4328 (N_4328,N_4138,N_4081);
xor U4329 (N_4329,N_4184,N_4196);
xor U4330 (N_4330,N_4147,N_4120);
nor U4331 (N_4331,N_4009,N_4047);
xnor U4332 (N_4332,N_4089,N_4173);
xor U4333 (N_4333,N_4088,N_4120);
xnor U4334 (N_4334,N_4081,N_4106);
and U4335 (N_4335,N_4144,N_4128);
nand U4336 (N_4336,N_4007,N_4144);
xor U4337 (N_4337,N_4020,N_4036);
nand U4338 (N_4338,N_4158,N_4082);
or U4339 (N_4339,N_4070,N_4085);
xnor U4340 (N_4340,N_4043,N_4094);
and U4341 (N_4341,N_4038,N_4000);
nor U4342 (N_4342,N_4134,N_4067);
or U4343 (N_4343,N_4105,N_4164);
nand U4344 (N_4344,N_4078,N_4003);
or U4345 (N_4345,N_4158,N_4145);
nand U4346 (N_4346,N_4110,N_4046);
and U4347 (N_4347,N_4093,N_4113);
and U4348 (N_4348,N_4194,N_4033);
nand U4349 (N_4349,N_4178,N_4025);
and U4350 (N_4350,N_4118,N_4144);
and U4351 (N_4351,N_4190,N_4027);
nand U4352 (N_4352,N_4163,N_4090);
xnor U4353 (N_4353,N_4154,N_4078);
and U4354 (N_4354,N_4038,N_4028);
nand U4355 (N_4355,N_4059,N_4072);
nor U4356 (N_4356,N_4158,N_4181);
xor U4357 (N_4357,N_4137,N_4019);
xnor U4358 (N_4358,N_4021,N_4001);
and U4359 (N_4359,N_4012,N_4017);
and U4360 (N_4360,N_4138,N_4135);
xor U4361 (N_4361,N_4060,N_4033);
nand U4362 (N_4362,N_4127,N_4004);
or U4363 (N_4363,N_4007,N_4039);
and U4364 (N_4364,N_4093,N_4111);
or U4365 (N_4365,N_4187,N_4191);
and U4366 (N_4366,N_4099,N_4051);
nor U4367 (N_4367,N_4005,N_4135);
or U4368 (N_4368,N_4056,N_4114);
or U4369 (N_4369,N_4199,N_4102);
nand U4370 (N_4370,N_4186,N_4151);
or U4371 (N_4371,N_4145,N_4152);
and U4372 (N_4372,N_4067,N_4016);
nand U4373 (N_4373,N_4124,N_4033);
and U4374 (N_4374,N_4010,N_4018);
or U4375 (N_4375,N_4156,N_4158);
nor U4376 (N_4376,N_4176,N_4040);
and U4377 (N_4377,N_4169,N_4110);
nor U4378 (N_4378,N_4058,N_4163);
nor U4379 (N_4379,N_4016,N_4000);
or U4380 (N_4380,N_4158,N_4183);
nor U4381 (N_4381,N_4186,N_4180);
and U4382 (N_4382,N_4069,N_4194);
nor U4383 (N_4383,N_4196,N_4074);
or U4384 (N_4384,N_4056,N_4058);
or U4385 (N_4385,N_4128,N_4059);
nor U4386 (N_4386,N_4070,N_4000);
nor U4387 (N_4387,N_4013,N_4134);
xnor U4388 (N_4388,N_4048,N_4037);
and U4389 (N_4389,N_4047,N_4105);
xnor U4390 (N_4390,N_4119,N_4020);
and U4391 (N_4391,N_4003,N_4182);
and U4392 (N_4392,N_4144,N_4064);
nor U4393 (N_4393,N_4155,N_4112);
or U4394 (N_4394,N_4173,N_4007);
and U4395 (N_4395,N_4069,N_4171);
nand U4396 (N_4396,N_4196,N_4044);
and U4397 (N_4397,N_4159,N_4005);
nor U4398 (N_4398,N_4164,N_4106);
and U4399 (N_4399,N_4109,N_4148);
xnor U4400 (N_4400,N_4246,N_4271);
nor U4401 (N_4401,N_4390,N_4351);
xor U4402 (N_4402,N_4309,N_4243);
xnor U4403 (N_4403,N_4328,N_4232);
nor U4404 (N_4404,N_4259,N_4288);
nand U4405 (N_4405,N_4329,N_4379);
xor U4406 (N_4406,N_4388,N_4222);
or U4407 (N_4407,N_4394,N_4307);
or U4408 (N_4408,N_4220,N_4302);
or U4409 (N_4409,N_4252,N_4343);
xnor U4410 (N_4410,N_4283,N_4339);
and U4411 (N_4411,N_4265,N_4399);
or U4412 (N_4412,N_4371,N_4317);
xor U4413 (N_4413,N_4321,N_4346);
xnor U4414 (N_4414,N_4396,N_4392);
nand U4415 (N_4415,N_4359,N_4268);
nand U4416 (N_4416,N_4256,N_4284);
nor U4417 (N_4417,N_4255,N_4237);
nand U4418 (N_4418,N_4245,N_4357);
nand U4419 (N_4419,N_4311,N_4253);
or U4420 (N_4420,N_4204,N_4214);
nand U4421 (N_4421,N_4327,N_4316);
xor U4422 (N_4422,N_4331,N_4369);
xor U4423 (N_4423,N_4342,N_4276);
xor U4424 (N_4424,N_4207,N_4282);
or U4425 (N_4425,N_4341,N_4247);
and U4426 (N_4426,N_4372,N_4293);
nand U4427 (N_4427,N_4242,N_4300);
and U4428 (N_4428,N_4257,N_4365);
and U4429 (N_4429,N_4345,N_4398);
xor U4430 (N_4430,N_4229,N_4385);
xnor U4431 (N_4431,N_4249,N_4298);
xnor U4432 (N_4432,N_4393,N_4285);
xnor U4433 (N_4433,N_4354,N_4362);
nand U4434 (N_4434,N_4294,N_4270);
nand U4435 (N_4435,N_4308,N_4320);
or U4436 (N_4436,N_4289,N_4366);
xnor U4437 (N_4437,N_4340,N_4292);
xnor U4438 (N_4438,N_4216,N_4315);
nor U4439 (N_4439,N_4387,N_4248);
nor U4440 (N_4440,N_4269,N_4212);
xor U4441 (N_4441,N_4350,N_4224);
or U4442 (N_4442,N_4376,N_4363);
and U4443 (N_4443,N_4240,N_4250);
nand U4444 (N_4444,N_4356,N_4344);
and U4445 (N_4445,N_4382,N_4295);
nand U4446 (N_4446,N_4262,N_4275);
nor U4447 (N_4447,N_4352,N_4335);
and U4448 (N_4448,N_4378,N_4215);
nor U4449 (N_4449,N_4213,N_4347);
nand U4450 (N_4450,N_4266,N_4274);
nand U4451 (N_4451,N_4312,N_4277);
nor U4452 (N_4452,N_4230,N_4313);
or U4453 (N_4453,N_4297,N_4200);
xor U4454 (N_4454,N_4304,N_4368);
or U4455 (N_4455,N_4210,N_4349);
xor U4456 (N_4456,N_4279,N_4384);
or U4457 (N_4457,N_4323,N_4367);
nor U4458 (N_4458,N_4226,N_4234);
xnor U4459 (N_4459,N_4201,N_4218);
nand U4460 (N_4460,N_4296,N_4391);
xor U4461 (N_4461,N_4395,N_4205);
xor U4462 (N_4462,N_4364,N_4383);
nor U4463 (N_4463,N_4272,N_4386);
and U4464 (N_4464,N_4374,N_4303);
or U4465 (N_4465,N_4290,N_4358);
or U4466 (N_4466,N_4299,N_4332);
nor U4467 (N_4467,N_4260,N_4219);
and U4468 (N_4468,N_4370,N_4330);
nand U4469 (N_4469,N_4231,N_4336);
and U4470 (N_4470,N_4221,N_4211);
nand U4471 (N_4471,N_4381,N_4326);
xor U4472 (N_4472,N_4324,N_4217);
xnor U4473 (N_4473,N_4263,N_4389);
or U4474 (N_4474,N_4267,N_4238);
and U4475 (N_4475,N_4235,N_4228);
nand U4476 (N_4476,N_4319,N_4338);
or U4477 (N_4477,N_4227,N_4334);
and U4478 (N_4478,N_4223,N_4203);
and U4479 (N_4479,N_4353,N_4258);
nor U4480 (N_4480,N_4273,N_4291);
and U4481 (N_4481,N_4202,N_4278);
and U4482 (N_4482,N_4286,N_4251);
nor U4483 (N_4483,N_4361,N_4355);
and U4484 (N_4484,N_4264,N_4261);
xnor U4485 (N_4485,N_4233,N_4280);
xor U4486 (N_4486,N_4239,N_4241);
nand U4487 (N_4487,N_4209,N_4281);
xnor U4488 (N_4488,N_4225,N_4373);
nor U4489 (N_4489,N_4301,N_4314);
xnor U4490 (N_4490,N_4287,N_4206);
xnor U4491 (N_4491,N_4325,N_4348);
nand U4492 (N_4492,N_4310,N_4318);
nor U4493 (N_4493,N_4244,N_4360);
or U4494 (N_4494,N_4236,N_4254);
nor U4495 (N_4495,N_4306,N_4377);
or U4496 (N_4496,N_4305,N_4208);
nand U4497 (N_4497,N_4397,N_4322);
and U4498 (N_4498,N_4333,N_4375);
and U4499 (N_4499,N_4337,N_4380);
or U4500 (N_4500,N_4388,N_4282);
nand U4501 (N_4501,N_4218,N_4253);
nor U4502 (N_4502,N_4306,N_4330);
nand U4503 (N_4503,N_4343,N_4263);
or U4504 (N_4504,N_4361,N_4308);
nor U4505 (N_4505,N_4364,N_4207);
nor U4506 (N_4506,N_4357,N_4238);
xor U4507 (N_4507,N_4394,N_4309);
and U4508 (N_4508,N_4238,N_4335);
and U4509 (N_4509,N_4252,N_4322);
nor U4510 (N_4510,N_4268,N_4212);
xnor U4511 (N_4511,N_4206,N_4357);
xnor U4512 (N_4512,N_4264,N_4233);
xnor U4513 (N_4513,N_4268,N_4255);
xor U4514 (N_4514,N_4233,N_4367);
nor U4515 (N_4515,N_4263,N_4208);
nor U4516 (N_4516,N_4388,N_4285);
xor U4517 (N_4517,N_4250,N_4224);
and U4518 (N_4518,N_4320,N_4319);
nor U4519 (N_4519,N_4373,N_4275);
and U4520 (N_4520,N_4234,N_4260);
and U4521 (N_4521,N_4254,N_4266);
and U4522 (N_4522,N_4295,N_4283);
or U4523 (N_4523,N_4201,N_4238);
or U4524 (N_4524,N_4334,N_4391);
nor U4525 (N_4525,N_4252,N_4316);
xor U4526 (N_4526,N_4319,N_4356);
or U4527 (N_4527,N_4392,N_4337);
nor U4528 (N_4528,N_4306,N_4300);
nand U4529 (N_4529,N_4339,N_4330);
and U4530 (N_4530,N_4276,N_4230);
or U4531 (N_4531,N_4360,N_4239);
nand U4532 (N_4532,N_4244,N_4286);
and U4533 (N_4533,N_4391,N_4255);
xnor U4534 (N_4534,N_4382,N_4205);
and U4535 (N_4535,N_4309,N_4260);
nor U4536 (N_4536,N_4308,N_4248);
and U4537 (N_4537,N_4320,N_4255);
nor U4538 (N_4538,N_4287,N_4332);
nand U4539 (N_4539,N_4259,N_4394);
and U4540 (N_4540,N_4344,N_4399);
nor U4541 (N_4541,N_4232,N_4376);
nor U4542 (N_4542,N_4254,N_4346);
nand U4543 (N_4543,N_4243,N_4302);
nand U4544 (N_4544,N_4354,N_4204);
nor U4545 (N_4545,N_4246,N_4332);
xor U4546 (N_4546,N_4249,N_4236);
xor U4547 (N_4547,N_4220,N_4228);
and U4548 (N_4548,N_4217,N_4399);
xnor U4549 (N_4549,N_4223,N_4207);
nor U4550 (N_4550,N_4317,N_4342);
or U4551 (N_4551,N_4388,N_4299);
xnor U4552 (N_4552,N_4289,N_4378);
or U4553 (N_4553,N_4205,N_4228);
xor U4554 (N_4554,N_4328,N_4217);
xor U4555 (N_4555,N_4225,N_4396);
nor U4556 (N_4556,N_4219,N_4384);
or U4557 (N_4557,N_4219,N_4282);
or U4558 (N_4558,N_4223,N_4384);
xor U4559 (N_4559,N_4272,N_4236);
and U4560 (N_4560,N_4369,N_4210);
nor U4561 (N_4561,N_4285,N_4234);
xor U4562 (N_4562,N_4391,N_4373);
xnor U4563 (N_4563,N_4294,N_4387);
nor U4564 (N_4564,N_4367,N_4334);
nand U4565 (N_4565,N_4345,N_4252);
nor U4566 (N_4566,N_4361,N_4236);
or U4567 (N_4567,N_4300,N_4207);
xnor U4568 (N_4568,N_4360,N_4248);
and U4569 (N_4569,N_4325,N_4262);
and U4570 (N_4570,N_4366,N_4213);
nor U4571 (N_4571,N_4255,N_4375);
xor U4572 (N_4572,N_4228,N_4246);
or U4573 (N_4573,N_4367,N_4356);
xnor U4574 (N_4574,N_4350,N_4397);
xnor U4575 (N_4575,N_4260,N_4385);
or U4576 (N_4576,N_4216,N_4390);
and U4577 (N_4577,N_4342,N_4275);
or U4578 (N_4578,N_4208,N_4238);
nand U4579 (N_4579,N_4220,N_4217);
xor U4580 (N_4580,N_4319,N_4310);
or U4581 (N_4581,N_4273,N_4307);
and U4582 (N_4582,N_4264,N_4226);
or U4583 (N_4583,N_4286,N_4369);
or U4584 (N_4584,N_4394,N_4311);
xnor U4585 (N_4585,N_4253,N_4308);
nand U4586 (N_4586,N_4267,N_4229);
nand U4587 (N_4587,N_4347,N_4360);
nor U4588 (N_4588,N_4241,N_4232);
or U4589 (N_4589,N_4228,N_4208);
and U4590 (N_4590,N_4295,N_4277);
nor U4591 (N_4591,N_4240,N_4299);
xnor U4592 (N_4592,N_4226,N_4386);
nor U4593 (N_4593,N_4256,N_4215);
xnor U4594 (N_4594,N_4223,N_4314);
nand U4595 (N_4595,N_4373,N_4240);
and U4596 (N_4596,N_4217,N_4375);
and U4597 (N_4597,N_4205,N_4203);
or U4598 (N_4598,N_4284,N_4288);
and U4599 (N_4599,N_4353,N_4357);
nand U4600 (N_4600,N_4517,N_4542);
nor U4601 (N_4601,N_4485,N_4503);
or U4602 (N_4602,N_4477,N_4529);
xnor U4603 (N_4603,N_4445,N_4426);
nor U4604 (N_4604,N_4502,N_4535);
and U4605 (N_4605,N_4488,N_4504);
nand U4606 (N_4606,N_4516,N_4554);
and U4607 (N_4607,N_4437,N_4547);
xor U4608 (N_4608,N_4549,N_4548);
and U4609 (N_4609,N_4439,N_4557);
and U4610 (N_4610,N_4544,N_4474);
nand U4611 (N_4611,N_4460,N_4508);
nor U4612 (N_4612,N_4462,N_4422);
nand U4613 (N_4613,N_4457,N_4561);
and U4614 (N_4614,N_4435,N_4467);
nand U4615 (N_4615,N_4563,N_4412);
nor U4616 (N_4616,N_4597,N_4434);
nor U4617 (N_4617,N_4414,N_4566);
nor U4618 (N_4618,N_4475,N_4491);
xor U4619 (N_4619,N_4428,N_4487);
or U4620 (N_4620,N_4486,N_4550);
xor U4621 (N_4621,N_4559,N_4472);
xor U4622 (N_4622,N_4525,N_4568);
or U4623 (N_4623,N_4518,N_4584);
and U4624 (N_4624,N_4429,N_4579);
or U4625 (N_4625,N_4416,N_4415);
nor U4626 (N_4626,N_4524,N_4587);
and U4627 (N_4627,N_4465,N_4501);
and U4628 (N_4628,N_4410,N_4484);
nor U4629 (N_4629,N_4471,N_4521);
and U4630 (N_4630,N_4569,N_4417);
xnor U4631 (N_4631,N_4585,N_4555);
or U4632 (N_4632,N_4522,N_4556);
nor U4633 (N_4633,N_4515,N_4523);
and U4634 (N_4634,N_4466,N_4514);
nor U4635 (N_4635,N_4532,N_4576);
and U4636 (N_4636,N_4469,N_4436);
nor U4637 (N_4637,N_4552,N_4551);
or U4638 (N_4638,N_4401,N_4404);
nor U4639 (N_4639,N_4574,N_4592);
nor U4640 (N_4640,N_4496,N_4406);
nor U4641 (N_4641,N_4407,N_4418);
xor U4642 (N_4642,N_4438,N_4571);
or U4643 (N_4643,N_4553,N_4573);
nand U4644 (N_4644,N_4423,N_4433);
nand U4645 (N_4645,N_4531,N_4468);
and U4646 (N_4646,N_4509,N_4409);
xor U4647 (N_4647,N_4432,N_4500);
and U4648 (N_4648,N_4538,N_4581);
xor U4649 (N_4649,N_4577,N_4490);
nand U4650 (N_4650,N_4447,N_4572);
xor U4651 (N_4651,N_4430,N_4530);
nand U4652 (N_4652,N_4441,N_4420);
or U4653 (N_4653,N_4408,N_4519);
xor U4654 (N_4654,N_4510,N_4583);
or U4655 (N_4655,N_4478,N_4575);
nor U4656 (N_4656,N_4456,N_4565);
or U4657 (N_4657,N_4564,N_4463);
and U4658 (N_4658,N_4578,N_4543);
and U4659 (N_4659,N_4580,N_4449);
xnor U4660 (N_4660,N_4541,N_4505);
or U4661 (N_4661,N_4567,N_4444);
and U4662 (N_4662,N_4537,N_4513);
nand U4663 (N_4663,N_4419,N_4470);
or U4664 (N_4664,N_4411,N_4479);
or U4665 (N_4665,N_4424,N_4450);
nor U4666 (N_4666,N_4452,N_4526);
or U4667 (N_4667,N_4480,N_4400);
and U4668 (N_4668,N_4442,N_4493);
xnor U4669 (N_4669,N_4499,N_4431);
xor U4670 (N_4670,N_4482,N_4582);
and U4671 (N_4671,N_4527,N_4598);
xor U4672 (N_4672,N_4594,N_4539);
nor U4673 (N_4673,N_4511,N_4520);
xor U4674 (N_4674,N_4459,N_4586);
and U4675 (N_4675,N_4589,N_4421);
and U4676 (N_4676,N_4533,N_4461);
or U4677 (N_4677,N_4536,N_4425);
and U4678 (N_4678,N_4453,N_4455);
or U4679 (N_4679,N_4596,N_4446);
nand U4680 (N_4680,N_4562,N_4476);
and U4681 (N_4681,N_4546,N_4534);
xnor U4682 (N_4682,N_4506,N_4591);
or U4683 (N_4683,N_4413,N_4560);
and U4684 (N_4684,N_4495,N_4528);
nand U4685 (N_4685,N_4440,N_4483);
or U4686 (N_4686,N_4595,N_4545);
xor U4687 (N_4687,N_4443,N_4492);
nor U4688 (N_4688,N_4599,N_4464);
or U4689 (N_4689,N_4405,N_4590);
and U4690 (N_4690,N_4402,N_4454);
or U4691 (N_4691,N_4448,N_4494);
nor U4692 (N_4692,N_4497,N_4473);
xnor U4693 (N_4693,N_4498,N_4570);
or U4694 (N_4694,N_4593,N_4481);
nor U4695 (N_4695,N_4403,N_4588);
and U4696 (N_4696,N_4489,N_4540);
and U4697 (N_4697,N_4507,N_4512);
nor U4698 (N_4698,N_4451,N_4427);
nor U4699 (N_4699,N_4558,N_4458);
xor U4700 (N_4700,N_4426,N_4478);
xor U4701 (N_4701,N_4454,N_4537);
or U4702 (N_4702,N_4549,N_4412);
and U4703 (N_4703,N_4489,N_4533);
nor U4704 (N_4704,N_4525,N_4557);
nand U4705 (N_4705,N_4420,N_4451);
or U4706 (N_4706,N_4414,N_4547);
xor U4707 (N_4707,N_4496,N_4450);
or U4708 (N_4708,N_4510,N_4553);
nor U4709 (N_4709,N_4472,N_4554);
and U4710 (N_4710,N_4404,N_4557);
nor U4711 (N_4711,N_4410,N_4587);
or U4712 (N_4712,N_4515,N_4401);
nand U4713 (N_4713,N_4529,N_4589);
nor U4714 (N_4714,N_4512,N_4435);
nor U4715 (N_4715,N_4425,N_4472);
or U4716 (N_4716,N_4489,N_4501);
and U4717 (N_4717,N_4545,N_4511);
nand U4718 (N_4718,N_4499,N_4574);
nand U4719 (N_4719,N_4473,N_4437);
xnor U4720 (N_4720,N_4477,N_4572);
nor U4721 (N_4721,N_4435,N_4579);
xnor U4722 (N_4722,N_4411,N_4496);
xor U4723 (N_4723,N_4501,N_4425);
nand U4724 (N_4724,N_4587,N_4419);
and U4725 (N_4725,N_4502,N_4579);
nand U4726 (N_4726,N_4420,N_4564);
xnor U4727 (N_4727,N_4521,N_4475);
nand U4728 (N_4728,N_4587,N_4400);
and U4729 (N_4729,N_4414,N_4518);
or U4730 (N_4730,N_4462,N_4540);
and U4731 (N_4731,N_4557,N_4567);
nor U4732 (N_4732,N_4591,N_4540);
and U4733 (N_4733,N_4547,N_4507);
nor U4734 (N_4734,N_4537,N_4536);
xor U4735 (N_4735,N_4436,N_4599);
nor U4736 (N_4736,N_4491,N_4496);
xnor U4737 (N_4737,N_4463,N_4524);
nor U4738 (N_4738,N_4406,N_4564);
and U4739 (N_4739,N_4475,N_4492);
and U4740 (N_4740,N_4540,N_4524);
and U4741 (N_4741,N_4495,N_4470);
or U4742 (N_4742,N_4580,N_4422);
nor U4743 (N_4743,N_4491,N_4472);
or U4744 (N_4744,N_4539,N_4551);
and U4745 (N_4745,N_4475,N_4409);
and U4746 (N_4746,N_4494,N_4495);
or U4747 (N_4747,N_4595,N_4587);
or U4748 (N_4748,N_4473,N_4581);
xor U4749 (N_4749,N_4410,N_4541);
nand U4750 (N_4750,N_4479,N_4498);
nor U4751 (N_4751,N_4599,N_4584);
nand U4752 (N_4752,N_4469,N_4402);
nand U4753 (N_4753,N_4431,N_4522);
nor U4754 (N_4754,N_4506,N_4558);
xnor U4755 (N_4755,N_4572,N_4444);
or U4756 (N_4756,N_4545,N_4431);
nand U4757 (N_4757,N_4472,N_4514);
nand U4758 (N_4758,N_4478,N_4412);
and U4759 (N_4759,N_4538,N_4552);
or U4760 (N_4760,N_4524,N_4498);
and U4761 (N_4761,N_4483,N_4549);
xnor U4762 (N_4762,N_4541,N_4437);
or U4763 (N_4763,N_4480,N_4500);
nand U4764 (N_4764,N_4471,N_4482);
or U4765 (N_4765,N_4495,N_4421);
xnor U4766 (N_4766,N_4439,N_4423);
xor U4767 (N_4767,N_4516,N_4526);
or U4768 (N_4768,N_4573,N_4447);
and U4769 (N_4769,N_4537,N_4530);
and U4770 (N_4770,N_4596,N_4539);
nor U4771 (N_4771,N_4438,N_4565);
and U4772 (N_4772,N_4402,N_4461);
xor U4773 (N_4773,N_4443,N_4597);
and U4774 (N_4774,N_4596,N_4492);
xor U4775 (N_4775,N_4570,N_4510);
or U4776 (N_4776,N_4562,N_4432);
xnor U4777 (N_4777,N_4556,N_4435);
nand U4778 (N_4778,N_4565,N_4498);
and U4779 (N_4779,N_4405,N_4573);
or U4780 (N_4780,N_4590,N_4544);
or U4781 (N_4781,N_4426,N_4488);
and U4782 (N_4782,N_4595,N_4441);
nor U4783 (N_4783,N_4572,N_4446);
xnor U4784 (N_4784,N_4587,N_4536);
nor U4785 (N_4785,N_4553,N_4583);
nand U4786 (N_4786,N_4583,N_4494);
nand U4787 (N_4787,N_4502,N_4464);
and U4788 (N_4788,N_4484,N_4448);
nor U4789 (N_4789,N_4534,N_4597);
nand U4790 (N_4790,N_4523,N_4498);
and U4791 (N_4791,N_4511,N_4566);
nor U4792 (N_4792,N_4436,N_4490);
nand U4793 (N_4793,N_4466,N_4488);
nand U4794 (N_4794,N_4490,N_4494);
nand U4795 (N_4795,N_4548,N_4589);
nor U4796 (N_4796,N_4520,N_4536);
and U4797 (N_4797,N_4453,N_4552);
xnor U4798 (N_4798,N_4455,N_4430);
and U4799 (N_4799,N_4527,N_4597);
nand U4800 (N_4800,N_4792,N_4793);
and U4801 (N_4801,N_4623,N_4710);
and U4802 (N_4802,N_4739,N_4683);
and U4803 (N_4803,N_4732,N_4772);
nand U4804 (N_4804,N_4620,N_4673);
and U4805 (N_4805,N_4604,N_4628);
nor U4806 (N_4806,N_4670,N_4656);
or U4807 (N_4807,N_4609,N_4615);
xnor U4808 (N_4808,N_4664,N_4635);
nand U4809 (N_4809,N_4744,N_4791);
nor U4810 (N_4810,N_4736,N_4611);
xnor U4811 (N_4811,N_4689,N_4750);
and U4812 (N_4812,N_4759,N_4799);
xnor U4813 (N_4813,N_4704,N_4684);
nor U4814 (N_4814,N_4754,N_4687);
xnor U4815 (N_4815,N_4662,N_4636);
nand U4816 (N_4816,N_4785,N_4703);
nor U4817 (N_4817,N_4752,N_4761);
nor U4818 (N_4818,N_4679,N_4601);
nand U4819 (N_4819,N_4630,N_4600);
xnor U4820 (N_4820,N_4671,N_4651);
xor U4821 (N_4821,N_4603,N_4779);
and U4822 (N_4822,N_4705,N_4728);
nor U4823 (N_4823,N_4777,N_4794);
nor U4824 (N_4824,N_4631,N_4738);
and U4825 (N_4825,N_4654,N_4789);
xnor U4826 (N_4826,N_4743,N_4780);
nand U4827 (N_4827,N_4709,N_4617);
and U4828 (N_4828,N_4667,N_4742);
or U4829 (N_4829,N_4757,N_4790);
and U4830 (N_4830,N_4714,N_4768);
nor U4831 (N_4831,N_4725,N_4658);
or U4832 (N_4832,N_4763,N_4678);
and U4833 (N_4833,N_4606,N_4756);
and U4834 (N_4834,N_4610,N_4717);
nor U4835 (N_4835,N_4698,N_4706);
and U4836 (N_4836,N_4663,N_4760);
and U4837 (N_4837,N_4638,N_4637);
xor U4838 (N_4838,N_4659,N_4781);
or U4839 (N_4839,N_4712,N_4769);
nor U4840 (N_4840,N_4682,N_4640);
or U4841 (N_4841,N_4716,N_4618);
nor U4842 (N_4842,N_4775,N_4696);
xor U4843 (N_4843,N_4741,N_4770);
xnor U4844 (N_4844,N_4612,N_4788);
nand U4845 (N_4845,N_4622,N_4608);
or U4846 (N_4846,N_4646,N_4633);
or U4847 (N_4847,N_4669,N_4748);
or U4848 (N_4848,N_4680,N_4639);
nor U4849 (N_4849,N_4730,N_4765);
or U4850 (N_4850,N_4735,N_4771);
and U4851 (N_4851,N_4647,N_4677);
nand U4852 (N_4852,N_4688,N_4681);
and U4853 (N_4853,N_4672,N_4711);
nand U4854 (N_4854,N_4634,N_4700);
and U4855 (N_4855,N_4650,N_4783);
and U4856 (N_4856,N_4675,N_4708);
or U4857 (N_4857,N_4727,N_4740);
and U4858 (N_4858,N_4702,N_4699);
nand U4859 (N_4859,N_4755,N_4686);
xnor U4860 (N_4860,N_4753,N_4632);
or U4861 (N_4861,N_4605,N_4643);
xor U4862 (N_4862,N_4690,N_4695);
nor U4863 (N_4863,N_4674,N_4713);
and U4864 (N_4864,N_4784,N_4767);
or U4865 (N_4865,N_4642,N_4697);
xnor U4866 (N_4866,N_4701,N_4661);
or U4867 (N_4867,N_4676,N_4707);
nand U4868 (N_4868,N_4758,N_4733);
xnor U4869 (N_4869,N_4719,N_4614);
and U4870 (N_4870,N_4715,N_4796);
xor U4871 (N_4871,N_4607,N_4720);
nand U4872 (N_4872,N_4657,N_4747);
xor U4873 (N_4873,N_4749,N_4778);
or U4874 (N_4874,N_4645,N_4774);
xnor U4875 (N_4875,N_4762,N_4624);
and U4876 (N_4876,N_4724,N_4648);
or U4877 (N_4877,N_4764,N_4782);
xor U4878 (N_4878,N_4629,N_4685);
xor U4879 (N_4879,N_4786,N_4766);
or U4880 (N_4880,N_4722,N_4729);
and U4881 (N_4881,N_4726,N_4795);
or U4882 (N_4882,N_4691,N_4692);
xnor U4883 (N_4883,N_4731,N_4602);
xnor U4884 (N_4884,N_4751,N_4776);
xor U4885 (N_4885,N_4668,N_4649);
xor U4886 (N_4886,N_4746,N_4625);
and U4887 (N_4887,N_4619,N_4693);
nor U4888 (N_4888,N_4627,N_4734);
nand U4889 (N_4889,N_4655,N_4626);
or U4890 (N_4890,N_4644,N_4797);
nand U4891 (N_4891,N_4737,N_4616);
nor U4892 (N_4892,N_4745,N_4798);
and U4893 (N_4893,N_4665,N_4694);
nand U4894 (N_4894,N_4718,N_4641);
nor U4895 (N_4895,N_4621,N_4723);
nand U4896 (N_4896,N_4653,N_4773);
nand U4897 (N_4897,N_4787,N_4666);
and U4898 (N_4898,N_4721,N_4613);
xor U4899 (N_4899,N_4660,N_4652);
or U4900 (N_4900,N_4676,N_4787);
and U4901 (N_4901,N_4631,N_4635);
or U4902 (N_4902,N_4667,N_4635);
xor U4903 (N_4903,N_4604,N_4790);
or U4904 (N_4904,N_4619,N_4761);
or U4905 (N_4905,N_4726,N_4638);
nand U4906 (N_4906,N_4662,N_4634);
nand U4907 (N_4907,N_4744,N_4783);
or U4908 (N_4908,N_4685,N_4698);
and U4909 (N_4909,N_4646,N_4743);
nor U4910 (N_4910,N_4647,N_4633);
xnor U4911 (N_4911,N_4713,N_4643);
or U4912 (N_4912,N_4689,N_4686);
or U4913 (N_4913,N_4791,N_4623);
nor U4914 (N_4914,N_4648,N_4600);
xnor U4915 (N_4915,N_4726,N_4648);
and U4916 (N_4916,N_4745,N_4628);
xnor U4917 (N_4917,N_4792,N_4783);
or U4918 (N_4918,N_4786,N_4744);
nand U4919 (N_4919,N_4769,N_4684);
and U4920 (N_4920,N_4757,N_4655);
nand U4921 (N_4921,N_4790,N_4649);
nor U4922 (N_4922,N_4730,N_4653);
and U4923 (N_4923,N_4609,N_4640);
nand U4924 (N_4924,N_4753,N_4778);
nor U4925 (N_4925,N_4795,N_4791);
nor U4926 (N_4926,N_4715,N_4711);
xnor U4927 (N_4927,N_4664,N_4628);
xnor U4928 (N_4928,N_4783,N_4717);
and U4929 (N_4929,N_4708,N_4640);
and U4930 (N_4930,N_4755,N_4772);
and U4931 (N_4931,N_4762,N_4750);
and U4932 (N_4932,N_4686,N_4600);
nand U4933 (N_4933,N_4689,N_4642);
xnor U4934 (N_4934,N_4709,N_4765);
or U4935 (N_4935,N_4761,N_4789);
or U4936 (N_4936,N_4743,N_4624);
and U4937 (N_4937,N_4684,N_4664);
nor U4938 (N_4938,N_4606,N_4761);
or U4939 (N_4939,N_4693,N_4705);
xnor U4940 (N_4940,N_4797,N_4632);
nor U4941 (N_4941,N_4785,N_4675);
nor U4942 (N_4942,N_4656,N_4716);
and U4943 (N_4943,N_4716,N_4768);
or U4944 (N_4944,N_4617,N_4683);
nand U4945 (N_4945,N_4779,N_4767);
or U4946 (N_4946,N_4655,N_4615);
or U4947 (N_4947,N_4748,N_4736);
or U4948 (N_4948,N_4768,N_4736);
or U4949 (N_4949,N_4775,N_4728);
nor U4950 (N_4950,N_4717,N_4657);
or U4951 (N_4951,N_4732,N_4651);
xnor U4952 (N_4952,N_4661,N_4783);
nand U4953 (N_4953,N_4681,N_4617);
or U4954 (N_4954,N_4641,N_4683);
nand U4955 (N_4955,N_4694,N_4747);
nand U4956 (N_4956,N_4670,N_4720);
xnor U4957 (N_4957,N_4660,N_4600);
nor U4958 (N_4958,N_4651,N_4750);
or U4959 (N_4959,N_4613,N_4621);
xor U4960 (N_4960,N_4600,N_4748);
or U4961 (N_4961,N_4658,N_4751);
nand U4962 (N_4962,N_4745,N_4759);
nand U4963 (N_4963,N_4699,N_4797);
nand U4964 (N_4964,N_4694,N_4640);
or U4965 (N_4965,N_4731,N_4736);
nand U4966 (N_4966,N_4697,N_4695);
nor U4967 (N_4967,N_4748,N_4771);
and U4968 (N_4968,N_4744,N_4674);
and U4969 (N_4969,N_4647,N_4757);
nor U4970 (N_4970,N_4732,N_4763);
and U4971 (N_4971,N_4742,N_4610);
nor U4972 (N_4972,N_4772,N_4631);
or U4973 (N_4973,N_4776,N_4660);
xnor U4974 (N_4974,N_4745,N_4755);
nand U4975 (N_4975,N_4679,N_4693);
nand U4976 (N_4976,N_4708,N_4721);
nand U4977 (N_4977,N_4684,N_4707);
and U4978 (N_4978,N_4643,N_4727);
or U4979 (N_4979,N_4799,N_4770);
or U4980 (N_4980,N_4651,N_4632);
and U4981 (N_4981,N_4736,N_4752);
nand U4982 (N_4982,N_4664,N_4668);
or U4983 (N_4983,N_4750,N_4770);
and U4984 (N_4984,N_4642,N_4622);
nor U4985 (N_4985,N_4610,N_4682);
nor U4986 (N_4986,N_4704,N_4649);
nand U4987 (N_4987,N_4755,N_4613);
xor U4988 (N_4988,N_4612,N_4682);
nand U4989 (N_4989,N_4677,N_4786);
nand U4990 (N_4990,N_4737,N_4733);
and U4991 (N_4991,N_4632,N_4775);
or U4992 (N_4992,N_4795,N_4708);
or U4993 (N_4993,N_4632,N_4615);
nand U4994 (N_4994,N_4732,N_4724);
and U4995 (N_4995,N_4615,N_4665);
or U4996 (N_4996,N_4636,N_4706);
xor U4997 (N_4997,N_4655,N_4648);
and U4998 (N_4998,N_4637,N_4673);
and U4999 (N_4999,N_4650,N_4620);
or U5000 (N_5000,N_4911,N_4916);
or U5001 (N_5001,N_4805,N_4848);
or U5002 (N_5002,N_4997,N_4946);
or U5003 (N_5003,N_4941,N_4937);
and U5004 (N_5004,N_4966,N_4964);
and U5005 (N_5005,N_4923,N_4986);
or U5006 (N_5006,N_4870,N_4882);
and U5007 (N_5007,N_4902,N_4801);
nor U5008 (N_5008,N_4921,N_4854);
nand U5009 (N_5009,N_4855,N_4829);
nand U5010 (N_5010,N_4813,N_4896);
or U5011 (N_5011,N_4908,N_4863);
and U5012 (N_5012,N_4980,N_4967);
and U5013 (N_5013,N_4977,N_4856);
nor U5014 (N_5014,N_4837,N_4850);
nor U5015 (N_5015,N_4942,N_4808);
and U5016 (N_5016,N_4958,N_4812);
nor U5017 (N_5017,N_4886,N_4959);
xnor U5018 (N_5018,N_4872,N_4979);
nor U5019 (N_5019,N_4931,N_4885);
nor U5020 (N_5020,N_4834,N_4995);
or U5021 (N_5021,N_4960,N_4840);
nor U5022 (N_5022,N_4918,N_4858);
nor U5023 (N_5023,N_4888,N_4982);
or U5024 (N_5024,N_4910,N_4853);
nand U5025 (N_5025,N_4810,N_4935);
nor U5026 (N_5026,N_4996,N_4922);
and U5027 (N_5027,N_4845,N_4957);
or U5028 (N_5028,N_4818,N_4831);
and U5029 (N_5029,N_4892,N_4968);
or U5030 (N_5030,N_4930,N_4807);
xor U5031 (N_5031,N_4815,N_4984);
or U5032 (N_5032,N_4838,N_4836);
or U5033 (N_5033,N_4976,N_4944);
xnor U5034 (N_5034,N_4919,N_4992);
and U5035 (N_5035,N_4945,N_4800);
or U5036 (N_5036,N_4867,N_4904);
nor U5037 (N_5037,N_4926,N_4938);
and U5038 (N_5038,N_4825,N_4933);
nand U5039 (N_5039,N_4993,N_4869);
nand U5040 (N_5040,N_4985,N_4887);
or U5041 (N_5041,N_4906,N_4828);
xor U5042 (N_5042,N_4894,N_4874);
and U5043 (N_5043,N_4927,N_4865);
and U5044 (N_5044,N_4806,N_4975);
and U5045 (N_5045,N_4903,N_4851);
nand U5046 (N_5046,N_4832,N_4974);
nor U5047 (N_5047,N_4844,N_4880);
xnor U5048 (N_5048,N_4897,N_4951);
nand U5049 (N_5049,N_4804,N_4820);
xnor U5050 (N_5050,N_4881,N_4816);
and U5051 (N_5051,N_4868,N_4924);
nand U5052 (N_5052,N_4988,N_4893);
and U5053 (N_5053,N_4972,N_4823);
xor U5054 (N_5054,N_4913,N_4849);
nand U5055 (N_5055,N_4981,N_4920);
nand U5056 (N_5056,N_4917,N_4879);
and U5057 (N_5057,N_4971,N_4999);
and U5058 (N_5058,N_4817,N_4847);
nor U5059 (N_5059,N_4803,N_4835);
xnor U5060 (N_5060,N_4833,N_4952);
xor U5061 (N_5061,N_4884,N_4873);
and U5062 (N_5062,N_4866,N_4895);
nor U5063 (N_5063,N_4954,N_4987);
nand U5064 (N_5064,N_4900,N_4991);
nand U5065 (N_5065,N_4905,N_4852);
nand U5066 (N_5066,N_4962,N_4841);
xor U5067 (N_5067,N_4862,N_4934);
xor U5068 (N_5068,N_4998,N_4929);
nand U5069 (N_5069,N_4963,N_4824);
xnor U5070 (N_5070,N_4898,N_4814);
or U5071 (N_5071,N_4990,N_4883);
and U5072 (N_5072,N_4943,N_4878);
xor U5073 (N_5073,N_4821,N_4912);
nand U5074 (N_5074,N_4901,N_4839);
nor U5075 (N_5075,N_4842,N_4915);
and U5076 (N_5076,N_4961,N_4861);
nor U5077 (N_5077,N_4953,N_4819);
xor U5078 (N_5078,N_4936,N_4955);
or U5079 (N_5079,N_4846,N_4932);
nor U5080 (N_5080,N_4890,N_4877);
and U5081 (N_5081,N_4970,N_4928);
nand U5082 (N_5082,N_4857,N_4973);
nor U5083 (N_5083,N_4940,N_4876);
or U5084 (N_5084,N_4830,N_4859);
and U5085 (N_5085,N_4860,N_4843);
nor U5086 (N_5086,N_4969,N_4899);
nand U5087 (N_5087,N_4827,N_4949);
nand U5088 (N_5088,N_4948,N_4864);
and U5089 (N_5089,N_4909,N_4978);
or U5090 (N_5090,N_4822,N_4950);
or U5091 (N_5091,N_4871,N_4907);
and U5092 (N_5092,N_4826,N_4914);
nor U5093 (N_5093,N_4965,N_4889);
nand U5094 (N_5094,N_4925,N_4989);
nand U5095 (N_5095,N_4809,N_4811);
nand U5096 (N_5096,N_4875,N_4939);
nand U5097 (N_5097,N_4956,N_4891);
or U5098 (N_5098,N_4994,N_4947);
nand U5099 (N_5099,N_4802,N_4983);
or U5100 (N_5100,N_4882,N_4893);
xnor U5101 (N_5101,N_4929,N_4835);
nand U5102 (N_5102,N_4813,N_4969);
nand U5103 (N_5103,N_4870,N_4876);
or U5104 (N_5104,N_4845,N_4977);
nor U5105 (N_5105,N_4883,N_4896);
xnor U5106 (N_5106,N_4886,N_4938);
nor U5107 (N_5107,N_4887,N_4822);
or U5108 (N_5108,N_4907,N_4950);
or U5109 (N_5109,N_4809,N_4929);
or U5110 (N_5110,N_4934,N_4828);
nand U5111 (N_5111,N_4815,N_4987);
nor U5112 (N_5112,N_4970,N_4838);
and U5113 (N_5113,N_4923,N_4946);
nand U5114 (N_5114,N_4987,N_4882);
or U5115 (N_5115,N_4810,N_4982);
nand U5116 (N_5116,N_4803,N_4842);
xor U5117 (N_5117,N_4804,N_4829);
xor U5118 (N_5118,N_4873,N_4857);
nand U5119 (N_5119,N_4988,N_4898);
and U5120 (N_5120,N_4980,N_4857);
and U5121 (N_5121,N_4972,N_4802);
nand U5122 (N_5122,N_4893,N_4821);
or U5123 (N_5123,N_4977,N_4897);
nand U5124 (N_5124,N_4929,N_4903);
and U5125 (N_5125,N_4996,N_4804);
nor U5126 (N_5126,N_4982,N_4944);
and U5127 (N_5127,N_4842,N_4898);
nand U5128 (N_5128,N_4831,N_4803);
xor U5129 (N_5129,N_4928,N_4968);
nor U5130 (N_5130,N_4888,N_4881);
nor U5131 (N_5131,N_4958,N_4855);
and U5132 (N_5132,N_4827,N_4881);
nor U5133 (N_5133,N_4874,N_4978);
nand U5134 (N_5134,N_4815,N_4913);
nand U5135 (N_5135,N_4897,N_4922);
or U5136 (N_5136,N_4950,N_4867);
and U5137 (N_5137,N_4989,N_4937);
nor U5138 (N_5138,N_4912,N_4819);
and U5139 (N_5139,N_4943,N_4837);
and U5140 (N_5140,N_4984,N_4839);
or U5141 (N_5141,N_4886,N_4990);
and U5142 (N_5142,N_4840,N_4922);
nor U5143 (N_5143,N_4849,N_4819);
or U5144 (N_5144,N_4984,N_4857);
and U5145 (N_5145,N_4814,N_4869);
and U5146 (N_5146,N_4949,N_4905);
nor U5147 (N_5147,N_4825,N_4921);
nand U5148 (N_5148,N_4973,N_4871);
xor U5149 (N_5149,N_4818,N_4983);
and U5150 (N_5150,N_4993,N_4945);
xor U5151 (N_5151,N_4895,N_4939);
nand U5152 (N_5152,N_4946,N_4950);
or U5153 (N_5153,N_4822,N_4936);
xnor U5154 (N_5154,N_4903,N_4972);
nand U5155 (N_5155,N_4969,N_4846);
xnor U5156 (N_5156,N_4954,N_4881);
and U5157 (N_5157,N_4878,N_4892);
and U5158 (N_5158,N_4863,N_4887);
or U5159 (N_5159,N_4963,N_4894);
and U5160 (N_5160,N_4918,N_4938);
or U5161 (N_5161,N_4859,N_4933);
xnor U5162 (N_5162,N_4946,N_4842);
or U5163 (N_5163,N_4969,N_4872);
or U5164 (N_5164,N_4944,N_4929);
or U5165 (N_5165,N_4848,N_4976);
nand U5166 (N_5166,N_4983,N_4838);
and U5167 (N_5167,N_4958,N_4878);
or U5168 (N_5168,N_4824,N_4868);
nand U5169 (N_5169,N_4942,N_4903);
nand U5170 (N_5170,N_4906,N_4967);
xor U5171 (N_5171,N_4815,N_4859);
nand U5172 (N_5172,N_4896,N_4939);
nor U5173 (N_5173,N_4914,N_4807);
nor U5174 (N_5174,N_4963,N_4915);
and U5175 (N_5175,N_4984,N_4950);
nand U5176 (N_5176,N_4842,N_4934);
nand U5177 (N_5177,N_4841,N_4979);
nor U5178 (N_5178,N_4970,N_4996);
nor U5179 (N_5179,N_4808,N_4944);
nand U5180 (N_5180,N_4800,N_4870);
and U5181 (N_5181,N_4941,N_4902);
nand U5182 (N_5182,N_4864,N_4917);
nand U5183 (N_5183,N_4835,N_4879);
or U5184 (N_5184,N_4997,N_4933);
nor U5185 (N_5185,N_4820,N_4806);
or U5186 (N_5186,N_4995,N_4905);
or U5187 (N_5187,N_4823,N_4900);
nand U5188 (N_5188,N_4884,N_4839);
and U5189 (N_5189,N_4843,N_4816);
and U5190 (N_5190,N_4833,N_4848);
nor U5191 (N_5191,N_4897,N_4995);
or U5192 (N_5192,N_4811,N_4844);
or U5193 (N_5193,N_4831,N_4861);
and U5194 (N_5194,N_4878,N_4954);
xor U5195 (N_5195,N_4932,N_4825);
and U5196 (N_5196,N_4866,N_4993);
and U5197 (N_5197,N_4967,N_4833);
nand U5198 (N_5198,N_4809,N_4858);
nand U5199 (N_5199,N_4809,N_4959);
xnor U5200 (N_5200,N_5048,N_5185);
or U5201 (N_5201,N_5096,N_5115);
nand U5202 (N_5202,N_5127,N_5182);
and U5203 (N_5203,N_5052,N_5084);
or U5204 (N_5204,N_5059,N_5179);
and U5205 (N_5205,N_5132,N_5167);
nand U5206 (N_5206,N_5144,N_5186);
nor U5207 (N_5207,N_5134,N_5033);
xor U5208 (N_5208,N_5024,N_5197);
xnor U5209 (N_5209,N_5086,N_5000);
nand U5210 (N_5210,N_5135,N_5133);
nand U5211 (N_5211,N_5142,N_5175);
and U5212 (N_5212,N_5071,N_5094);
xor U5213 (N_5213,N_5015,N_5166);
and U5214 (N_5214,N_5170,N_5128);
and U5215 (N_5215,N_5005,N_5063);
or U5216 (N_5216,N_5074,N_5168);
nor U5217 (N_5217,N_5020,N_5110);
and U5218 (N_5218,N_5145,N_5093);
nand U5219 (N_5219,N_5113,N_5049);
nand U5220 (N_5220,N_5191,N_5088);
xor U5221 (N_5221,N_5176,N_5046);
and U5222 (N_5222,N_5114,N_5019);
and U5223 (N_5223,N_5180,N_5097);
nor U5224 (N_5224,N_5045,N_5009);
and U5225 (N_5225,N_5111,N_5174);
and U5226 (N_5226,N_5154,N_5003);
and U5227 (N_5227,N_5139,N_5161);
and U5228 (N_5228,N_5010,N_5075);
nor U5229 (N_5229,N_5108,N_5006);
or U5230 (N_5230,N_5160,N_5196);
nand U5231 (N_5231,N_5137,N_5156);
or U5232 (N_5232,N_5173,N_5053);
nand U5233 (N_5233,N_5038,N_5195);
nor U5234 (N_5234,N_5150,N_5007);
and U5235 (N_5235,N_5055,N_5169);
nand U5236 (N_5236,N_5021,N_5014);
nor U5237 (N_5237,N_5162,N_5079);
and U5238 (N_5238,N_5172,N_5130);
xnor U5239 (N_5239,N_5190,N_5092);
and U5240 (N_5240,N_5061,N_5044);
xnor U5241 (N_5241,N_5032,N_5087);
or U5242 (N_5242,N_5037,N_5028);
or U5243 (N_5243,N_5068,N_5100);
and U5244 (N_5244,N_5159,N_5104);
or U5245 (N_5245,N_5077,N_5157);
and U5246 (N_5246,N_5085,N_5107);
nand U5247 (N_5247,N_5118,N_5163);
xor U5248 (N_5248,N_5123,N_5136);
nand U5249 (N_5249,N_5188,N_5004);
nand U5250 (N_5250,N_5031,N_5147);
and U5251 (N_5251,N_5112,N_5072);
xnor U5252 (N_5252,N_5057,N_5164);
or U5253 (N_5253,N_5051,N_5109);
nor U5254 (N_5254,N_5039,N_5105);
or U5255 (N_5255,N_5078,N_5125);
nand U5256 (N_5256,N_5148,N_5189);
or U5257 (N_5257,N_5198,N_5155);
and U5258 (N_5258,N_5001,N_5013);
xor U5259 (N_5259,N_5102,N_5029);
xnor U5260 (N_5260,N_5040,N_5023);
or U5261 (N_5261,N_5117,N_5025);
xor U5262 (N_5262,N_5121,N_5103);
and U5263 (N_5263,N_5042,N_5011);
nor U5264 (N_5264,N_5120,N_5143);
nand U5265 (N_5265,N_5140,N_5062);
nand U5266 (N_5266,N_5126,N_5089);
nand U5267 (N_5267,N_5095,N_5076);
xnor U5268 (N_5268,N_5119,N_5194);
nand U5269 (N_5269,N_5193,N_5199);
xnor U5270 (N_5270,N_5122,N_5091);
xor U5271 (N_5271,N_5016,N_5138);
and U5272 (N_5272,N_5030,N_5192);
or U5273 (N_5273,N_5043,N_5036);
nand U5274 (N_5274,N_5069,N_5083);
or U5275 (N_5275,N_5177,N_5050);
nand U5276 (N_5276,N_5008,N_5054);
or U5277 (N_5277,N_5129,N_5012);
and U5278 (N_5278,N_5152,N_5181);
nor U5279 (N_5279,N_5060,N_5131);
or U5280 (N_5280,N_5178,N_5165);
nor U5281 (N_5281,N_5073,N_5018);
nor U5282 (N_5282,N_5017,N_5070);
or U5283 (N_5283,N_5098,N_5082);
or U5284 (N_5284,N_5171,N_5187);
nor U5285 (N_5285,N_5067,N_5027);
or U5286 (N_5286,N_5026,N_5146);
nor U5287 (N_5287,N_5184,N_5034);
or U5288 (N_5288,N_5047,N_5080);
nand U5289 (N_5289,N_5022,N_5058);
xor U5290 (N_5290,N_5041,N_5149);
and U5291 (N_5291,N_5158,N_5056);
nand U5292 (N_5292,N_5141,N_5065);
nor U5293 (N_5293,N_5153,N_5064);
nand U5294 (N_5294,N_5081,N_5002);
and U5295 (N_5295,N_5106,N_5116);
nand U5296 (N_5296,N_5124,N_5066);
xor U5297 (N_5297,N_5183,N_5101);
xor U5298 (N_5298,N_5151,N_5090);
nand U5299 (N_5299,N_5035,N_5099);
nor U5300 (N_5300,N_5107,N_5073);
nor U5301 (N_5301,N_5182,N_5083);
xor U5302 (N_5302,N_5014,N_5139);
or U5303 (N_5303,N_5190,N_5104);
or U5304 (N_5304,N_5099,N_5027);
and U5305 (N_5305,N_5100,N_5168);
or U5306 (N_5306,N_5062,N_5051);
and U5307 (N_5307,N_5004,N_5048);
nor U5308 (N_5308,N_5175,N_5134);
xor U5309 (N_5309,N_5106,N_5138);
nand U5310 (N_5310,N_5156,N_5121);
nor U5311 (N_5311,N_5089,N_5086);
or U5312 (N_5312,N_5195,N_5058);
or U5313 (N_5313,N_5049,N_5081);
and U5314 (N_5314,N_5177,N_5071);
and U5315 (N_5315,N_5171,N_5197);
xor U5316 (N_5316,N_5178,N_5179);
or U5317 (N_5317,N_5131,N_5095);
nand U5318 (N_5318,N_5077,N_5171);
nand U5319 (N_5319,N_5051,N_5087);
and U5320 (N_5320,N_5061,N_5077);
nor U5321 (N_5321,N_5181,N_5094);
or U5322 (N_5322,N_5049,N_5124);
nor U5323 (N_5323,N_5028,N_5085);
xnor U5324 (N_5324,N_5183,N_5189);
xor U5325 (N_5325,N_5092,N_5059);
nor U5326 (N_5326,N_5039,N_5104);
or U5327 (N_5327,N_5198,N_5186);
xnor U5328 (N_5328,N_5041,N_5023);
nor U5329 (N_5329,N_5156,N_5177);
or U5330 (N_5330,N_5089,N_5021);
or U5331 (N_5331,N_5007,N_5183);
nor U5332 (N_5332,N_5057,N_5093);
nor U5333 (N_5333,N_5116,N_5144);
or U5334 (N_5334,N_5070,N_5119);
or U5335 (N_5335,N_5024,N_5100);
or U5336 (N_5336,N_5155,N_5179);
xor U5337 (N_5337,N_5193,N_5195);
nor U5338 (N_5338,N_5149,N_5139);
nor U5339 (N_5339,N_5096,N_5048);
nand U5340 (N_5340,N_5134,N_5160);
xor U5341 (N_5341,N_5184,N_5149);
nand U5342 (N_5342,N_5113,N_5057);
and U5343 (N_5343,N_5082,N_5035);
and U5344 (N_5344,N_5062,N_5190);
xor U5345 (N_5345,N_5041,N_5165);
or U5346 (N_5346,N_5179,N_5007);
nand U5347 (N_5347,N_5013,N_5105);
or U5348 (N_5348,N_5064,N_5089);
and U5349 (N_5349,N_5113,N_5186);
or U5350 (N_5350,N_5135,N_5058);
and U5351 (N_5351,N_5089,N_5199);
or U5352 (N_5352,N_5048,N_5014);
nand U5353 (N_5353,N_5035,N_5199);
xnor U5354 (N_5354,N_5134,N_5081);
or U5355 (N_5355,N_5110,N_5063);
nand U5356 (N_5356,N_5027,N_5072);
xor U5357 (N_5357,N_5157,N_5158);
nand U5358 (N_5358,N_5107,N_5032);
nor U5359 (N_5359,N_5154,N_5095);
nor U5360 (N_5360,N_5002,N_5086);
xor U5361 (N_5361,N_5010,N_5162);
nand U5362 (N_5362,N_5075,N_5104);
nor U5363 (N_5363,N_5044,N_5055);
or U5364 (N_5364,N_5129,N_5199);
nand U5365 (N_5365,N_5135,N_5067);
xnor U5366 (N_5366,N_5143,N_5174);
xnor U5367 (N_5367,N_5049,N_5154);
nand U5368 (N_5368,N_5075,N_5178);
nand U5369 (N_5369,N_5140,N_5028);
and U5370 (N_5370,N_5120,N_5025);
xor U5371 (N_5371,N_5023,N_5042);
xor U5372 (N_5372,N_5127,N_5103);
and U5373 (N_5373,N_5199,N_5151);
nand U5374 (N_5374,N_5067,N_5188);
or U5375 (N_5375,N_5122,N_5110);
xor U5376 (N_5376,N_5040,N_5035);
xnor U5377 (N_5377,N_5092,N_5013);
and U5378 (N_5378,N_5075,N_5043);
xnor U5379 (N_5379,N_5171,N_5099);
nand U5380 (N_5380,N_5169,N_5096);
xnor U5381 (N_5381,N_5122,N_5059);
nand U5382 (N_5382,N_5195,N_5159);
nor U5383 (N_5383,N_5126,N_5004);
nor U5384 (N_5384,N_5188,N_5010);
and U5385 (N_5385,N_5034,N_5102);
and U5386 (N_5386,N_5018,N_5135);
nand U5387 (N_5387,N_5067,N_5092);
nor U5388 (N_5388,N_5018,N_5060);
xnor U5389 (N_5389,N_5121,N_5148);
xor U5390 (N_5390,N_5155,N_5106);
and U5391 (N_5391,N_5141,N_5170);
nand U5392 (N_5392,N_5196,N_5143);
nand U5393 (N_5393,N_5098,N_5126);
xnor U5394 (N_5394,N_5041,N_5011);
and U5395 (N_5395,N_5173,N_5127);
or U5396 (N_5396,N_5173,N_5155);
nor U5397 (N_5397,N_5085,N_5176);
nand U5398 (N_5398,N_5049,N_5089);
nor U5399 (N_5399,N_5123,N_5165);
xor U5400 (N_5400,N_5202,N_5305);
nor U5401 (N_5401,N_5357,N_5206);
and U5402 (N_5402,N_5396,N_5289);
nand U5403 (N_5403,N_5285,N_5394);
xnor U5404 (N_5404,N_5388,N_5264);
nand U5405 (N_5405,N_5350,N_5251);
nor U5406 (N_5406,N_5235,N_5329);
nor U5407 (N_5407,N_5359,N_5252);
or U5408 (N_5408,N_5232,N_5324);
or U5409 (N_5409,N_5327,N_5383);
and U5410 (N_5410,N_5227,N_5243);
xor U5411 (N_5411,N_5293,N_5333);
xnor U5412 (N_5412,N_5209,N_5328);
nor U5413 (N_5413,N_5247,N_5210);
xnor U5414 (N_5414,N_5279,N_5381);
nand U5415 (N_5415,N_5355,N_5341);
nor U5416 (N_5416,N_5398,N_5220);
nand U5417 (N_5417,N_5391,N_5307);
xnor U5418 (N_5418,N_5317,N_5239);
or U5419 (N_5419,N_5248,N_5298);
and U5420 (N_5420,N_5306,N_5343);
xor U5421 (N_5421,N_5346,N_5218);
nor U5422 (N_5422,N_5253,N_5284);
and U5423 (N_5423,N_5219,N_5356);
or U5424 (N_5424,N_5214,N_5382);
nor U5425 (N_5425,N_5311,N_5376);
xor U5426 (N_5426,N_5315,N_5348);
xnor U5427 (N_5427,N_5352,N_5222);
or U5428 (N_5428,N_5387,N_5399);
xnor U5429 (N_5429,N_5349,N_5308);
nor U5430 (N_5430,N_5332,N_5303);
or U5431 (N_5431,N_5286,N_5313);
and U5432 (N_5432,N_5360,N_5300);
nand U5433 (N_5433,N_5246,N_5345);
nand U5434 (N_5434,N_5371,N_5347);
and U5435 (N_5435,N_5295,N_5330);
nor U5436 (N_5436,N_5296,N_5212);
xnor U5437 (N_5437,N_5336,N_5390);
nor U5438 (N_5438,N_5310,N_5258);
nand U5439 (N_5439,N_5326,N_5229);
nor U5440 (N_5440,N_5379,N_5364);
nor U5441 (N_5441,N_5255,N_5369);
nand U5442 (N_5442,N_5297,N_5301);
nand U5443 (N_5443,N_5380,N_5234);
nor U5444 (N_5444,N_5339,N_5254);
or U5445 (N_5445,N_5216,N_5265);
nand U5446 (N_5446,N_5373,N_5276);
nor U5447 (N_5447,N_5211,N_5244);
or U5448 (N_5448,N_5316,N_5319);
and U5449 (N_5449,N_5240,N_5268);
nor U5450 (N_5450,N_5290,N_5367);
or U5451 (N_5451,N_5325,N_5304);
or U5452 (N_5452,N_5385,N_5272);
xor U5453 (N_5453,N_5250,N_5392);
xnor U5454 (N_5454,N_5335,N_5217);
xnor U5455 (N_5455,N_5269,N_5374);
or U5456 (N_5456,N_5368,N_5283);
nand U5457 (N_5457,N_5291,N_5204);
or U5458 (N_5458,N_5249,N_5275);
and U5459 (N_5459,N_5351,N_5337);
or U5460 (N_5460,N_5208,N_5215);
or U5461 (N_5461,N_5256,N_5205);
nand U5462 (N_5462,N_5362,N_5245);
nand U5463 (N_5463,N_5231,N_5302);
or U5464 (N_5464,N_5213,N_5358);
nor U5465 (N_5465,N_5226,N_5271);
xor U5466 (N_5466,N_5267,N_5228);
nor U5467 (N_5467,N_5340,N_5318);
xor U5468 (N_5468,N_5323,N_5363);
and U5469 (N_5469,N_5224,N_5354);
or U5470 (N_5470,N_5378,N_5281);
nand U5471 (N_5471,N_5263,N_5370);
nand U5472 (N_5472,N_5242,N_5273);
or U5473 (N_5473,N_5207,N_5334);
or U5474 (N_5474,N_5280,N_5299);
nand U5475 (N_5475,N_5366,N_5266);
and U5476 (N_5476,N_5389,N_5377);
xor U5477 (N_5477,N_5375,N_5331);
xnor U5478 (N_5478,N_5260,N_5322);
and U5479 (N_5479,N_5236,N_5277);
nor U5480 (N_5480,N_5344,N_5274);
or U5481 (N_5481,N_5312,N_5261);
nor U5482 (N_5482,N_5230,N_5225);
nor U5483 (N_5483,N_5238,N_5314);
or U5484 (N_5484,N_5221,N_5233);
xor U5485 (N_5485,N_5361,N_5200);
nor U5486 (N_5486,N_5282,N_5223);
xnor U5487 (N_5487,N_5393,N_5353);
xnor U5488 (N_5488,N_5342,N_5321);
nor U5489 (N_5489,N_5384,N_5278);
and U5490 (N_5490,N_5386,N_5309);
nand U5491 (N_5491,N_5287,N_5259);
nand U5492 (N_5492,N_5294,N_5395);
and U5493 (N_5493,N_5372,N_5237);
and U5494 (N_5494,N_5270,N_5262);
nand U5495 (N_5495,N_5397,N_5365);
nand U5496 (N_5496,N_5292,N_5288);
nand U5497 (N_5497,N_5320,N_5257);
xor U5498 (N_5498,N_5201,N_5338);
and U5499 (N_5499,N_5241,N_5203);
nand U5500 (N_5500,N_5365,N_5265);
nor U5501 (N_5501,N_5312,N_5359);
or U5502 (N_5502,N_5245,N_5227);
or U5503 (N_5503,N_5256,N_5351);
nand U5504 (N_5504,N_5313,N_5243);
or U5505 (N_5505,N_5220,N_5247);
xnor U5506 (N_5506,N_5286,N_5282);
nor U5507 (N_5507,N_5209,N_5368);
nor U5508 (N_5508,N_5383,N_5279);
nand U5509 (N_5509,N_5275,N_5379);
and U5510 (N_5510,N_5306,N_5281);
nand U5511 (N_5511,N_5314,N_5288);
xnor U5512 (N_5512,N_5259,N_5333);
and U5513 (N_5513,N_5278,N_5395);
or U5514 (N_5514,N_5372,N_5208);
nand U5515 (N_5515,N_5345,N_5314);
or U5516 (N_5516,N_5246,N_5377);
xnor U5517 (N_5517,N_5222,N_5362);
nor U5518 (N_5518,N_5316,N_5294);
xor U5519 (N_5519,N_5255,N_5397);
xnor U5520 (N_5520,N_5384,N_5319);
nand U5521 (N_5521,N_5204,N_5310);
or U5522 (N_5522,N_5337,N_5364);
nor U5523 (N_5523,N_5228,N_5358);
or U5524 (N_5524,N_5388,N_5287);
xnor U5525 (N_5525,N_5309,N_5211);
or U5526 (N_5526,N_5239,N_5203);
or U5527 (N_5527,N_5306,N_5207);
xor U5528 (N_5528,N_5248,N_5397);
nor U5529 (N_5529,N_5226,N_5303);
or U5530 (N_5530,N_5256,N_5329);
nor U5531 (N_5531,N_5261,N_5331);
nor U5532 (N_5532,N_5280,N_5255);
or U5533 (N_5533,N_5334,N_5298);
and U5534 (N_5534,N_5294,N_5330);
xor U5535 (N_5535,N_5219,N_5388);
and U5536 (N_5536,N_5275,N_5386);
or U5537 (N_5537,N_5270,N_5258);
or U5538 (N_5538,N_5217,N_5276);
nand U5539 (N_5539,N_5247,N_5344);
or U5540 (N_5540,N_5266,N_5339);
and U5541 (N_5541,N_5339,N_5323);
and U5542 (N_5542,N_5288,N_5336);
xor U5543 (N_5543,N_5360,N_5271);
nor U5544 (N_5544,N_5349,N_5394);
xnor U5545 (N_5545,N_5242,N_5371);
xnor U5546 (N_5546,N_5327,N_5298);
or U5547 (N_5547,N_5269,N_5382);
nor U5548 (N_5548,N_5356,N_5351);
or U5549 (N_5549,N_5389,N_5362);
or U5550 (N_5550,N_5231,N_5395);
xnor U5551 (N_5551,N_5265,N_5245);
xor U5552 (N_5552,N_5208,N_5270);
nor U5553 (N_5553,N_5380,N_5296);
and U5554 (N_5554,N_5384,N_5225);
and U5555 (N_5555,N_5207,N_5393);
nand U5556 (N_5556,N_5239,N_5208);
nor U5557 (N_5557,N_5387,N_5220);
and U5558 (N_5558,N_5351,N_5344);
xnor U5559 (N_5559,N_5329,N_5288);
nor U5560 (N_5560,N_5350,N_5203);
nor U5561 (N_5561,N_5214,N_5224);
xnor U5562 (N_5562,N_5338,N_5391);
xor U5563 (N_5563,N_5355,N_5382);
and U5564 (N_5564,N_5344,N_5298);
or U5565 (N_5565,N_5259,N_5362);
or U5566 (N_5566,N_5228,N_5269);
or U5567 (N_5567,N_5271,N_5272);
xnor U5568 (N_5568,N_5364,N_5206);
nor U5569 (N_5569,N_5330,N_5371);
xnor U5570 (N_5570,N_5291,N_5284);
nand U5571 (N_5571,N_5307,N_5206);
or U5572 (N_5572,N_5234,N_5210);
xnor U5573 (N_5573,N_5223,N_5347);
nand U5574 (N_5574,N_5295,N_5261);
nor U5575 (N_5575,N_5327,N_5310);
nand U5576 (N_5576,N_5212,N_5322);
and U5577 (N_5577,N_5219,N_5394);
xor U5578 (N_5578,N_5276,N_5206);
nor U5579 (N_5579,N_5268,N_5343);
xnor U5580 (N_5580,N_5219,N_5384);
nand U5581 (N_5581,N_5381,N_5335);
or U5582 (N_5582,N_5306,N_5251);
or U5583 (N_5583,N_5332,N_5243);
nand U5584 (N_5584,N_5327,N_5243);
and U5585 (N_5585,N_5349,N_5297);
and U5586 (N_5586,N_5291,N_5395);
and U5587 (N_5587,N_5331,N_5222);
nor U5588 (N_5588,N_5219,N_5222);
nor U5589 (N_5589,N_5244,N_5209);
or U5590 (N_5590,N_5306,N_5257);
nor U5591 (N_5591,N_5349,N_5315);
xnor U5592 (N_5592,N_5266,N_5340);
and U5593 (N_5593,N_5296,N_5214);
nor U5594 (N_5594,N_5217,N_5225);
and U5595 (N_5595,N_5284,N_5308);
nand U5596 (N_5596,N_5231,N_5342);
nand U5597 (N_5597,N_5258,N_5317);
nand U5598 (N_5598,N_5301,N_5239);
nor U5599 (N_5599,N_5241,N_5263);
xor U5600 (N_5600,N_5590,N_5403);
or U5601 (N_5601,N_5547,N_5516);
nor U5602 (N_5602,N_5566,N_5543);
or U5603 (N_5603,N_5520,N_5593);
nand U5604 (N_5604,N_5468,N_5570);
nor U5605 (N_5605,N_5506,N_5545);
nor U5606 (N_5606,N_5582,N_5558);
and U5607 (N_5607,N_5578,N_5544);
and U5608 (N_5608,N_5562,N_5458);
and U5609 (N_5609,N_5503,N_5555);
and U5610 (N_5610,N_5575,N_5454);
or U5611 (N_5611,N_5510,N_5477);
and U5612 (N_5612,N_5494,N_5469);
nor U5613 (N_5613,N_5493,N_5482);
xor U5614 (N_5614,N_5412,N_5483);
xnor U5615 (N_5615,N_5489,N_5530);
nand U5616 (N_5616,N_5485,N_5492);
nor U5617 (N_5617,N_5596,N_5434);
or U5618 (N_5618,N_5527,N_5406);
nand U5619 (N_5619,N_5580,N_5572);
nand U5620 (N_5620,N_5420,N_5442);
nor U5621 (N_5621,N_5504,N_5505);
nand U5622 (N_5622,N_5560,N_5535);
and U5623 (N_5623,N_5522,N_5411);
nand U5624 (N_5624,N_5481,N_5509);
xnor U5625 (N_5625,N_5508,N_5511);
or U5626 (N_5626,N_5437,N_5488);
or U5627 (N_5627,N_5444,N_5588);
and U5628 (N_5628,N_5402,N_5445);
xor U5629 (N_5629,N_5490,N_5597);
and U5630 (N_5630,N_5410,N_5497);
xor U5631 (N_5631,N_5447,N_5529);
nor U5632 (N_5632,N_5595,N_5592);
or U5633 (N_5633,N_5408,N_5479);
nor U5634 (N_5634,N_5589,N_5400);
or U5635 (N_5635,N_5579,N_5586);
xor U5636 (N_5636,N_5553,N_5542);
and U5637 (N_5637,N_5443,N_5428);
and U5638 (N_5638,N_5591,N_5474);
nand U5639 (N_5639,N_5568,N_5460);
nor U5640 (N_5640,N_5416,N_5540);
or U5641 (N_5641,N_5463,N_5452);
or U5642 (N_5642,N_5432,N_5431);
or U5643 (N_5643,N_5405,N_5475);
and U5644 (N_5644,N_5495,N_5557);
xor U5645 (N_5645,N_5513,N_5409);
nor U5646 (N_5646,N_5532,N_5531);
nor U5647 (N_5647,N_5414,N_5491);
nor U5648 (N_5648,N_5476,N_5450);
xnor U5649 (N_5649,N_5541,N_5466);
or U5650 (N_5650,N_5563,N_5449);
nand U5651 (N_5651,N_5561,N_5523);
and U5652 (N_5652,N_5424,N_5467);
xnor U5653 (N_5653,N_5521,N_5430);
and U5654 (N_5654,N_5427,N_5528);
nand U5655 (N_5655,N_5581,N_5576);
or U5656 (N_5656,N_5587,N_5425);
or U5657 (N_5657,N_5515,N_5500);
xnor U5658 (N_5658,N_5585,N_5407);
and U5659 (N_5659,N_5517,N_5539);
nor U5660 (N_5660,N_5546,N_5423);
or U5661 (N_5661,N_5524,N_5459);
nor U5662 (N_5662,N_5413,N_5533);
xnor U5663 (N_5663,N_5565,N_5550);
and U5664 (N_5664,N_5456,N_5426);
nor U5665 (N_5665,N_5470,N_5417);
nand U5666 (N_5666,N_5429,N_5538);
and U5667 (N_5667,N_5583,N_5573);
or U5668 (N_5668,N_5419,N_5441);
or U5669 (N_5669,N_5438,N_5552);
nor U5670 (N_5670,N_5418,N_5451);
nand U5671 (N_5671,N_5422,N_5537);
or U5672 (N_5672,N_5501,N_5549);
and U5673 (N_5673,N_5512,N_5448);
and U5674 (N_5674,N_5401,N_5487);
nor U5675 (N_5675,N_5571,N_5433);
or U5676 (N_5676,N_5496,N_5478);
nand U5677 (N_5677,N_5594,N_5480);
and U5678 (N_5678,N_5554,N_5536);
or U5679 (N_5679,N_5471,N_5551);
nand U5680 (N_5680,N_5548,N_5584);
nand U5681 (N_5681,N_5502,N_5574);
and U5682 (N_5682,N_5404,N_5525);
or U5683 (N_5683,N_5564,N_5462);
xnor U5684 (N_5684,N_5464,N_5473);
nor U5685 (N_5685,N_5439,N_5567);
and U5686 (N_5686,N_5534,N_5486);
xor U5687 (N_5687,N_5599,N_5577);
and U5688 (N_5688,N_5465,N_5598);
xnor U5689 (N_5689,N_5484,N_5436);
xor U5690 (N_5690,N_5440,N_5446);
xor U5691 (N_5691,N_5518,N_5559);
or U5692 (N_5692,N_5453,N_5519);
xor U5693 (N_5693,N_5472,N_5499);
nand U5694 (N_5694,N_5556,N_5455);
or U5695 (N_5695,N_5461,N_5457);
or U5696 (N_5696,N_5415,N_5526);
nand U5697 (N_5697,N_5421,N_5514);
and U5698 (N_5698,N_5569,N_5507);
nand U5699 (N_5699,N_5498,N_5435);
and U5700 (N_5700,N_5550,N_5429);
or U5701 (N_5701,N_5468,N_5521);
or U5702 (N_5702,N_5426,N_5527);
nand U5703 (N_5703,N_5441,N_5527);
xnor U5704 (N_5704,N_5497,N_5443);
xor U5705 (N_5705,N_5491,N_5554);
or U5706 (N_5706,N_5513,N_5572);
xor U5707 (N_5707,N_5461,N_5594);
xnor U5708 (N_5708,N_5597,N_5563);
nand U5709 (N_5709,N_5573,N_5584);
xnor U5710 (N_5710,N_5468,N_5511);
nor U5711 (N_5711,N_5524,N_5485);
nand U5712 (N_5712,N_5549,N_5592);
or U5713 (N_5713,N_5541,N_5441);
xor U5714 (N_5714,N_5466,N_5584);
nor U5715 (N_5715,N_5502,N_5516);
nor U5716 (N_5716,N_5574,N_5499);
or U5717 (N_5717,N_5420,N_5413);
nand U5718 (N_5718,N_5400,N_5505);
or U5719 (N_5719,N_5589,N_5449);
xnor U5720 (N_5720,N_5448,N_5433);
xor U5721 (N_5721,N_5422,N_5481);
nor U5722 (N_5722,N_5472,N_5410);
nor U5723 (N_5723,N_5466,N_5411);
and U5724 (N_5724,N_5427,N_5485);
nor U5725 (N_5725,N_5440,N_5537);
or U5726 (N_5726,N_5441,N_5448);
or U5727 (N_5727,N_5442,N_5422);
or U5728 (N_5728,N_5485,N_5412);
nor U5729 (N_5729,N_5578,N_5565);
nand U5730 (N_5730,N_5537,N_5530);
nand U5731 (N_5731,N_5539,N_5520);
nor U5732 (N_5732,N_5409,N_5599);
and U5733 (N_5733,N_5408,N_5575);
nand U5734 (N_5734,N_5561,N_5515);
nand U5735 (N_5735,N_5468,N_5425);
or U5736 (N_5736,N_5559,N_5599);
or U5737 (N_5737,N_5555,N_5546);
nand U5738 (N_5738,N_5591,N_5404);
or U5739 (N_5739,N_5443,N_5597);
or U5740 (N_5740,N_5537,N_5404);
xnor U5741 (N_5741,N_5561,N_5599);
or U5742 (N_5742,N_5575,N_5588);
xnor U5743 (N_5743,N_5551,N_5418);
nor U5744 (N_5744,N_5423,N_5529);
or U5745 (N_5745,N_5450,N_5424);
nor U5746 (N_5746,N_5499,N_5550);
nand U5747 (N_5747,N_5570,N_5590);
and U5748 (N_5748,N_5523,N_5440);
xor U5749 (N_5749,N_5404,N_5550);
nand U5750 (N_5750,N_5539,N_5427);
xor U5751 (N_5751,N_5599,N_5501);
or U5752 (N_5752,N_5434,N_5575);
nand U5753 (N_5753,N_5525,N_5501);
nand U5754 (N_5754,N_5443,N_5473);
xor U5755 (N_5755,N_5583,N_5578);
and U5756 (N_5756,N_5461,N_5501);
nand U5757 (N_5757,N_5468,N_5497);
xor U5758 (N_5758,N_5439,N_5407);
xor U5759 (N_5759,N_5568,N_5558);
nand U5760 (N_5760,N_5450,N_5502);
nor U5761 (N_5761,N_5412,N_5530);
nor U5762 (N_5762,N_5460,N_5587);
and U5763 (N_5763,N_5469,N_5465);
xnor U5764 (N_5764,N_5576,N_5552);
nor U5765 (N_5765,N_5406,N_5487);
or U5766 (N_5766,N_5459,N_5475);
nand U5767 (N_5767,N_5404,N_5439);
nor U5768 (N_5768,N_5503,N_5508);
nor U5769 (N_5769,N_5453,N_5531);
and U5770 (N_5770,N_5523,N_5589);
xnor U5771 (N_5771,N_5424,N_5466);
xnor U5772 (N_5772,N_5520,N_5469);
xnor U5773 (N_5773,N_5491,N_5426);
nor U5774 (N_5774,N_5410,N_5429);
or U5775 (N_5775,N_5460,N_5493);
xor U5776 (N_5776,N_5586,N_5588);
and U5777 (N_5777,N_5590,N_5426);
nand U5778 (N_5778,N_5587,N_5455);
nand U5779 (N_5779,N_5537,N_5485);
and U5780 (N_5780,N_5477,N_5578);
xnor U5781 (N_5781,N_5576,N_5463);
or U5782 (N_5782,N_5472,N_5473);
xnor U5783 (N_5783,N_5579,N_5416);
xnor U5784 (N_5784,N_5421,N_5468);
or U5785 (N_5785,N_5421,N_5549);
nor U5786 (N_5786,N_5440,N_5564);
or U5787 (N_5787,N_5557,N_5537);
xor U5788 (N_5788,N_5456,N_5536);
xor U5789 (N_5789,N_5495,N_5457);
xor U5790 (N_5790,N_5428,N_5553);
nand U5791 (N_5791,N_5444,N_5525);
nand U5792 (N_5792,N_5524,N_5523);
or U5793 (N_5793,N_5445,N_5511);
and U5794 (N_5794,N_5488,N_5431);
xnor U5795 (N_5795,N_5505,N_5570);
xor U5796 (N_5796,N_5541,N_5539);
nand U5797 (N_5797,N_5596,N_5529);
or U5798 (N_5798,N_5493,N_5441);
or U5799 (N_5799,N_5532,N_5450);
nor U5800 (N_5800,N_5646,N_5790);
xor U5801 (N_5801,N_5755,N_5642);
xnor U5802 (N_5802,N_5675,N_5655);
and U5803 (N_5803,N_5653,N_5629);
nor U5804 (N_5804,N_5616,N_5719);
or U5805 (N_5805,N_5758,N_5715);
nor U5806 (N_5806,N_5651,N_5620);
xnor U5807 (N_5807,N_5634,N_5729);
nor U5808 (N_5808,N_5659,N_5695);
or U5809 (N_5809,N_5626,N_5673);
xor U5810 (N_5810,N_5615,N_5609);
nand U5811 (N_5811,N_5681,N_5795);
nor U5812 (N_5812,N_5714,N_5747);
and U5813 (N_5813,N_5777,N_5774);
nor U5814 (N_5814,N_5627,N_5722);
nor U5815 (N_5815,N_5611,N_5754);
xnor U5816 (N_5816,N_5643,N_5772);
and U5817 (N_5817,N_5671,N_5635);
nor U5818 (N_5818,N_5640,N_5721);
nor U5819 (N_5819,N_5785,N_5760);
nor U5820 (N_5820,N_5696,N_5786);
and U5821 (N_5821,N_5607,N_5664);
or U5822 (N_5822,N_5663,N_5660);
or U5823 (N_5823,N_5776,N_5743);
nand U5824 (N_5824,N_5711,N_5728);
and U5825 (N_5825,N_5784,N_5674);
or U5826 (N_5826,N_5649,N_5689);
nor U5827 (N_5827,N_5742,N_5667);
and U5828 (N_5828,N_5628,N_5633);
and U5829 (N_5829,N_5691,N_5683);
and U5830 (N_5830,N_5676,N_5717);
and U5831 (N_5831,N_5767,N_5782);
and U5832 (N_5832,N_5704,N_5617);
and U5833 (N_5833,N_5613,N_5693);
xor U5834 (N_5834,N_5604,N_5713);
or U5835 (N_5835,N_5606,N_5708);
or U5836 (N_5836,N_5766,N_5666);
or U5837 (N_5837,N_5656,N_5623);
or U5838 (N_5838,N_5688,N_5731);
xor U5839 (N_5839,N_5770,N_5789);
and U5840 (N_5840,N_5793,N_5738);
nor U5841 (N_5841,N_5724,N_5677);
and U5842 (N_5842,N_5707,N_5727);
xnor U5843 (N_5843,N_5796,N_5661);
nor U5844 (N_5844,N_5716,N_5737);
and U5845 (N_5845,N_5602,N_5679);
nand U5846 (N_5846,N_5763,N_5712);
and U5847 (N_5847,N_5734,N_5709);
xor U5848 (N_5848,N_5736,N_5787);
nand U5849 (N_5849,N_5687,N_5775);
nor U5850 (N_5850,N_5798,N_5684);
or U5851 (N_5851,N_5749,N_5632);
or U5852 (N_5852,N_5610,N_5757);
or U5853 (N_5853,N_5750,N_5639);
xor U5854 (N_5854,N_5654,N_5745);
or U5855 (N_5855,N_5769,N_5658);
nand U5856 (N_5856,N_5703,N_5608);
nand U5857 (N_5857,N_5652,N_5601);
nand U5858 (N_5858,N_5637,N_5768);
nor U5859 (N_5859,N_5702,N_5622);
or U5860 (N_5860,N_5762,N_5759);
xor U5861 (N_5861,N_5630,N_5718);
nor U5862 (N_5862,N_5725,N_5732);
and U5863 (N_5863,N_5765,N_5624);
xnor U5864 (N_5864,N_5690,N_5698);
nand U5865 (N_5865,N_5773,N_5764);
xor U5866 (N_5866,N_5794,N_5780);
nand U5867 (N_5867,N_5779,N_5699);
or U5868 (N_5868,N_5752,N_5631);
or U5869 (N_5869,N_5603,N_5612);
xor U5870 (N_5870,N_5700,N_5706);
xnor U5871 (N_5871,N_5701,N_5791);
xnor U5872 (N_5872,N_5726,N_5621);
nand U5873 (N_5873,N_5670,N_5778);
or U5874 (N_5874,N_5665,N_5705);
xnor U5875 (N_5875,N_5710,N_5668);
and U5876 (N_5876,N_5625,N_5799);
xor U5877 (N_5877,N_5662,N_5748);
and U5878 (N_5878,N_5650,N_5685);
nand U5879 (N_5879,N_5686,N_5741);
nor U5880 (N_5880,N_5771,N_5614);
and U5881 (N_5881,N_5744,N_5723);
nor U5882 (N_5882,N_5761,N_5781);
or U5883 (N_5883,N_5648,N_5751);
nand U5884 (N_5884,N_5753,N_5638);
and U5885 (N_5885,N_5605,N_5788);
xor U5886 (N_5886,N_5735,N_5733);
and U5887 (N_5887,N_5682,N_5618);
xor U5888 (N_5888,N_5692,N_5740);
nor U5889 (N_5889,N_5644,N_5694);
or U5890 (N_5890,N_5797,N_5792);
and U5891 (N_5891,N_5783,N_5678);
nor U5892 (N_5892,N_5645,N_5730);
nand U5893 (N_5893,N_5756,N_5669);
and U5894 (N_5894,N_5720,N_5600);
xor U5895 (N_5895,N_5746,N_5641);
xnor U5896 (N_5896,N_5680,N_5672);
and U5897 (N_5897,N_5739,N_5657);
xor U5898 (N_5898,N_5619,N_5636);
and U5899 (N_5899,N_5647,N_5697);
and U5900 (N_5900,N_5730,N_5737);
xnor U5901 (N_5901,N_5607,N_5616);
nand U5902 (N_5902,N_5709,N_5778);
xnor U5903 (N_5903,N_5709,N_5708);
or U5904 (N_5904,N_5622,N_5723);
or U5905 (N_5905,N_5715,N_5781);
nor U5906 (N_5906,N_5738,N_5611);
nor U5907 (N_5907,N_5633,N_5748);
and U5908 (N_5908,N_5742,N_5680);
nor U5909 (N_5909,N_5795,N_5716);
or U5910 (N_5910,N_5617,N_5720);
xor U5911 (N_5911,N_5629,N_5672);
nor U5912 (N_5912,N_5698,N_5626);
nor U5913 (N_5913,N_5765,N_5786);
nor U5914 (N_5914,N_5602,N_5623);
xnor U5915 (N_5915,N_5751,N_5742);
and U5916 (N_5916,N_5627,N_5795);
nand U5917 (N_5917,N_5611,N_5769);
and U5918 (N_5918,N_5604,N_5754);
and U5919 (N_5919,N_5712,N_5625);
xnor U5920 (N_5920,N_5656,N_5728);
or U5921 (N_5921,N_5732,N_5657);
nand U5922 (N_5922,N_5767,N_5785);
nand U5923 (N_5923,N_5709,N_5712);
xnor U5924 (N_5924,N_5756,N_5679);
and U5925 (N_5925,N_5712,N_5751);
nor U5926 (N_5926,N_5706,N_5621);
or U5927 (N_5927,N_5795,N_5684);
xnor U5928 (N_5928,N_5785,N_5759);
or U5929 (N_5929,N_5795,N_5644);
xnor U5930 (N_5930,N_5641,N_5743);
nand U5931 (N_5931,N_5799,N_5744);
and U5932 (N_5932,N_5789,N_5635);
xnor U5933 (N_5933,N_5749,N_5791);
or U5934 (N_5934,N_5728,N_5666);
nand U5935 (N_5935,N_5660,N_5680);
nor U5936 (N_5936,N_5726,N_5676);
or U5937 (N_5937,N_5601,N_5787);
or U5938 (N_5938,N_5742,N_5740);
xor U5939 (N_5939,N_5749,N_5784);
and U5940 (N_5940,N_5799,N_5719);
or U5941 (N_5941,N_5634,N_5799);
nand U5942 (N_5942,N_5634,N_5641);
nand U5943 (N_5943,N_5728,N_5767);
nor U5944 (N_5944,N_5793,N_5773);
nor U5945 (N_5945,N_5689,N_5766);
and U5946 (N_5946,N_5716,N_5629);
or U5947 (N_5947,N_5792,N_5672);
or U5948 (N_5948,N_5652,N_5695);
nor U5949 (N_5949,N_5765,N_5648);
or U5950 (N_5950,N_5668,N_5674);
xor U5951 (N_5951,N_5739,N_5704);
xnor U5952 (N_5952,N_5651,N_5702);
and U5953 (N_5953,N_5756,N_5770);
and U5954 (N_5954,N_5730,N_5692);
or U5955 (N_5955,N_5773,N_5707);
or U5956 (N_5956,N_5715,N_5733);
nand U5957 (N_5957,N_5765,N_5603);
or U5958 (N_5958,N_5708,N_5631);
or U5959 (N_5959,N_5788,N_5786);
or U5960 (N_5960,N_5764,N_5662);
nor U5961 (N_5961,N_5672,N_5695);
nand U5962 (N_5962,N_5757,N_5761);
xnor U5963 (N_5963,N_5663,N_5610);
or U5964 (N_5964,N_5617,N_5637);
nor U5965 (N_5965,N_5728,N_5749);
or U5966 (N_5966,N_5699,N_5607);
xnor U5967 (N_5967,N_5754,N_5720);
and U5968 (N_5968,N_5755,N_5700);
xor U5969 (N_5969,N_5656,N_5614);
nor U5970 (N_5970,N_5719,N_5681);
or U5971 (N_5971,N_5712,N_5762);
nand U5972 (N_5972,N_5785,N_5645);
nor U5973 (N_5973,N_5672,N_5759);
nand U5974 (N_5974,N_5763,N_5625);
xnor U5975 (N_5975,N_5757,N_5755);
or U5976 (N_5976,N_5696,N_5780);
xnor U5977 (N_5977,N_5731,N_5609);
and U5978 (N_5978,N_5630,N_5697);
xor U5979 (N_5979,N_5706,N_5701);
nor U5980 (N_5980,N_5616,N_5721);
xor U5981 (N_5981,N_5724,N_5717);
and U5982 (N_5982,N_5713,N_5765);
nand U5983 (N_5983,N_5658,N_5688);
and U5984 (N_5984,N_5675,N_5702);
nor U5985 (N_5985,N_5607,N_5650);
xnor U5986 (N_5986,N_5633,N_5639);
nor U5987 (N_5987,N_5659,N_5676);
nor U5988 (N_5988,N_5632,N_5730);
and U5989 (N_5989,N_5656,N_5729);
and U5990 (N_5990,N_5615,N_5778);
nor U5991 (N_5991,N_5630,N_5601);
xor U5992 (N_5992,N_5701,N_5799);
or U5993 (N_5993,N_5605,N_5740);
xnor U5994 (N_5994,N_5684,N_5711);
nand U5995 (N_5995,N_5605,N_5713);
nor U5996 (N_5996,N_5776,N_5723);
xnor U5997 (N_5997,N_5624,N_5645);
nand U5998 (N_5998,N_5717,N_5698);
and U5999 (N_5999,N_5776,N_5612);
nand U6000 (N_6000,N_5879,N_5883);
xnor U6001 (N_6001,N_5919,N_5828);
or U6002 (N_6002,N_5948,N_5819);
nand U6003 (N_6003,N_5845,N_5816);
or U6004 (N_6004,N_5903,N_5848);
nand U6005 (N_6005,N_5870,N_5977);
nor U6006 (N_6006,N_5830,N_5872);
and U6007 (N_6007,N_5923,N_5986);
or U6008 (N_6008,N_5865,N_5924);
nor U6009 (N_6009,N_5899,N_5955);
or U6010 (N_6010,N_5969,N_5914);
nand U6011 (N_6011,N_5809,N_5979);
xor U6012 (N_6012,N_5889,N_5972);
and U6013 (N_6013,N_5929,N_5854);
nand U6014 (N_6014,N_5999,N_5930);
or U6015 (N_6015,N_5947,N_5911);
nor U6016 (N_6016,N_5866,N_5834);
nor U6017 (N_6017,N_5925,N_5991);
nor U6018 (N_6018,N_5805,N_5881);
nand U6019 (N_6019,N_5884,N_5811);
nor U6020 (N_6020,N_5898,N_5968);
or U6021 (N_6021,N_5803,N_5998);
nand U6022 (N_6022,N_5934,N_5994);
nand U6023 (N_6023,N_5807,N_5910);
and U6024 (N_6024,N_5992,N_5931);
nor U6025 (N_6025,N_5974,N_5840);
or U6026 (N_6026,N_5836,N_5944);
and U6027 (N_6027,N_5829,N_5863);
xnor U6028 (N_6028,N_5970,N_5943);
nand U6029 (N_6029,N_5961,N_5936);
or U6030 (N_6030,N_5984,N_5907);
nor U6031 (N_6031,N_5933,N_5942);
nor U6032 (N_6032,N_5886,N_5808);
or U6033 (N_6033,N_5843,N_5940);
nand U6034 (N_6034,N_5815,N_5952);
nor U6035 (N_6035,N_5927,N_5892);
nand U6036 (N_6036,N_5876,N_5902);
nand U6037 (N_6037,N_5856,N_5964);
or U6038 (N_6038,N_5820,N_5827);
nor U6039 (N_6039,N_5921,N_5978);
nor U6040 (N_6040,N_5855,N_5896);
xor U6041 (N_6041,N_5963,N_5966);
nor U6042 (N_6042,N_5837,N_5853);
nor U6043 (N_6043,N_5945,N_5953);
nand U6044 (N_6044,N_5922,N_5976);
and U6045 (N_6045,N_5800,N_5877);
and U6046 (N_6046,N_5965,N_5859);
or U6047 (N_6047,N_5812,N_5821);
and U6048 (N_6048,N_5960,N_5817);
and U6049 (N_6049,N_5905,N_5860);
xor U6050 (N_6050,N_5990,N_5823);
xor U6051 (N_6051,N_5871,N_5920);
nand U6052 (N_6052,N_5904,N_5842);
xnor U6053 (N_6053,N_5802,N_5841);
or U6054 (N_6054,N_5875,N_5975);
xor U6055 (N_6055,N_5838,N_5891);
nand U6056 (N_6056,N_5814,N_5826);
and U6057 (N_6057,N_5913,N_5824);
nand U6058 (N_6058,N_5868,N_5833);
and U6059 (N_6059,N_5996,N_5873);
nand U6060 (N_6060,N_5894,N_5857);
or U6061 (N_6061,N_5971,N_5980);
nor U6062 (N_6062,N_5983,N_5887);
nor U6063 (N_6063,N_5878,N_5981);
and U6064 (N_6064,N_5818,N_5989);
nor U6065 (N_6065,N_5844,N_5987);
and U6066 (N_6066,N_5852,N_5890);
or U6067 (N_6067,N_5935,N_5956);
xnor U6068 (N_6068,N_5835,N_5908);
xnor U6069 (N_6069,N_5888,N_5941);
xor U6070 (N_6070,N_5906,N_5926);
nand U6071 (N_6071,N_5849,N_5982);
xnor U6072 (N_6072,N_5831,N_5958);
nand U6073 (N_6073,N_5885,N_5967);
xor U6074 (N_6074,N_5946,N_5938);
nand U6075 (N_6075,N_5901,N_5973);
nor U6076 (N_6076,N_5850,N_5932);
xnor U6077 (N_6077,N_5916,N_5893);
nand U6078 (N_6078,N_5993,N_5851);
nand U6079 (N_6079,N_5861,N_5867);
xnor U6080 (N_6080,N_5825,N_5839);
xnor U6081 (N_6081,N_5915,N_5962);
xnor U6082 (N_6082,N_5804,N_5928);
and U6083 (N_6083,N_5806,N_5988);
and U6084 (N_6084,N_5950,N_5937);
or U6085 (N_6085,N_5939,N_5874);
xnor U6086 (N_6086,N_5951,N_5900);
nand U6087 (N_6087,N_5858,N_5957);
nor U6088 (N_6088,N_5862,N_5949);
and U6089 (N_6089,N_5810,N_5918);
xnor U6090 (N_6090,N_5864,N_5917);
nor U6091 (N_6091,N_5895,N_5909);
xor U6092 (N_6092,N_5954,N_5995);
nand U6093 (N_6093,N_5912,N_5959);
xor U6094 (N_6094,N_5822,N_5869);
xor U6095 (N_6095,N_5832,N_5846);
or U6096 (N_6096,N_5847,N_5897);
and U6097 (N_6097,N_5985,N_5882);
and U6098 (N_6098,N_5801,N_5880);
nor U6099 (N_6099,N_5997,N_5813);
and U6100 (N_6100,N_5927,N_5963);
nand U6101 (N_6101,N_5874,N_5871);
nand U6102 (N_6102,N_5936,N_5898);
nand U6103 (N_6103,N_5814,N_5827);
and U6104 (N_6104,N_5945,N_5988);
xnor U6105 (N_6105,N_5823,N_5899);
and U6106 (N_6106,N_5911,N_5923);
or U6107 (N_6107,N_5866,N_5877);
nand U6108 (N_6108,N_5983,N_5854);
or U6109 (N_6109,N_5977,N_5984);
xnor U6110 (N_6110,N_5880,N_5920);
or U6111 (N_6111,N_5804,N_5907);
and U6112 (N_6112,N_5935,N_5964);
nand U6113 (N_6113,N_5838,N_5845);
and U6114 (N_6114,N_5976,N_5820);
nor U6115 (N_6115,N_5951,N_5938);
and U6116 (N_6116,N_5884,N_5827);
and U6117 (N_6117,N_5961,N_5856);
or U6118 (N_6118,N_5823,N_5937);
and U6119 (N_6119,N_5969,N_5833);
nor U6120 (N_6120,N_5830,N_5999);
xor U6121 (N_6121,N_5903,N_5857);
and U6122 (N_6122,N_5805,N_5974);
and U6123 (N_6123,N_5975,N_5967);
nand U6124 (N_6124,N_5936,N_5882);
nor U6125 (N_6125,N_5893,N_5807);
nor U6126 (N_6126,N_5902,N_5924);
nor U6127 (N_6127,N_5818,N_5872);
nand U6128 (N_6128,N_5968,N_5960);
or U6129 (N_6129,N_5911,N_5824);
nand U6130 (N_6130,N_5964,N_5866);
nand U6131 (N_6131,N_5974,N_5835);
and U6132 (N_6132,N_5964,N_5821);
and U6133 (N_6133,N_5941,N_5825);
nor U6134 (N_6134,N_5922,N_5819);
nor U6135 (N_6135,N_5824,N_5825);
and U6136 (N_6136,N_5918,N_5916);
nor U6137 (N_6137,N_5943,N_5900);
xor U6138 (N_6138,N_5973,N_5871);
xor U6139 (N_6139,N_5904,N_5996);
nand U6140 (N_6140,N_5846,N_5957);
xnor U6141 (N_6141,N_5970,N_5803);
nor U6142 (N_6142,N_5912,N_5867);
and U6143 (N_6143,N_5917,N_5990);
xor U6144 (N_6144,N_5942,N_5902);
and U6145 (N_6145,N_5913,N_5830);
and U6146 (N_6146,N_5936,N_5813);
xor U6147 (N_6147,N_5957,N_5933);
or U6148 (N_6148,N_5986,N_5866);
nor U6149 (N_6149,N_5888,N_5825);
nor U6150 (N_6150,N_5951,N_5968);
and U6151 (N_6151,N_5853,N_5959);
xnor U6152 (N_6152,N_5820,N_5985);
nor U6153 (N_6153,N_5822,N_5897);
xor U6154 (N_6154,N_5818,N_5978);
and U6155 (N_6155,N_5888,N_5822);
nor U6156 (N_6156,N_5954,N_5882);
nand U6157 (N_6157,N_5828,N_5914);
nor U6158 (N_6158,N_5857,N_5820);
xor U6159 (N_6159,N_5914,N_5887);
or U6160 (N_6160,N_5851,N_5821);
xnor U6161 (N_6161,N_5820,N_5965);
or U6162 (N_6162,N_5989,N_5814);
nor U6163 (N_6163,N_5926,N_5882);
and U6164 (N_6164,N_5911,N_5962);
or U6165 (N_6165,N_5881,N_5856);
nand U6166 (N_6166,N_5875,N_5938);
and U6167 (N_6167,N_5832,N_5879);
xnor U6168 (N_6168,N_5948,N_5912);
and U6169 (N_6169,N_5961,N_5995);
nor U6170 (N_6170,N_5863,N_5969);
or U6171 (N_6171,N_5841,N_5816);
nor U6172 (N_6172,N_5944,N_5816);
or U6173 (N_6173,N_5814,N_5800);
and U6174 (N_6174,N_5971,N_5876);
xnor U6175 (N_6175,N_5890,N_5800);
nand U6176 (N_6176,N_5930,N_5874);
and U6177 (N_6177,N_5832,N_5844);
nor U6178 (N_6178,N_5989,N_5887);
nor U6179 (N_6179,N_5949,N_5891);
and U6180 (N_6180,N_5854,N_5995);
nand U6181 (N_6181,N_5999,N_5954);
and U6182 (N_6182,N_5853,N_5922);
and U6183 (N_6183,N_5987,N_5977);
or U6184 (N_6184,N_5806,N_5967);
xor U6185 (N_6185,N_5915,N_5882);
and U6186 (N_6186,N_5955,N_5860);
xnor U6187 (N_6187,N_5929,N_5980);
nor U6188 (N_6188,N_5900,N_5965);
xor U6189 (N_6189,N_5885,N_5922);
nor U6190 (N_6190,N_5826,N_5844);
nor U6191 (N_6191,N_5873,N_5951);
or U6192 (N_6192,N_5950,N_5860);
and U6193 (N_6193,N_5927,N_5891);
xnor U6194 (N_6194,N_5870,N_5920);
or U6195 (N_6195,N_5822,N_5894);
or U6196 (N_6196,N_5967,N_5847);
and U6197 (N_6197,N_5877,N_5996);
xor U6198 (N_6198,N_5860,N_5816);
nand U6199 (N_6199,N_5883,N_5867);
and U6200 (N_6200,N_6072,N_6032);
or U6201 (N_6201,N_6071,N_6033);
nor U6202 (N_6202,N_6146,N_6158);
nor U6203 (N_6203,N_6180,N_6073);
or U6204 (N_6204,N_6150,N_6029);
or U6205 (N_6205,N_6002,N_6186);
and U6206 (N_6206,N_6088,N_6021);
xor U6207 (N_6207,N_6095,N_6114);
or U6208 (N_6208,N_6022,N_6074);
nand U6209 (N_6209,N_6078,N_6178);
nand U6210 (N_6210,N_6182,N_6188);
xor U6211 (N_6211,N_6007,N_6037);
and U6212 (N_6212,N_6082,N_6039);
and U6213 (N_6213,N_6080,N_6132);
and U6214 (N_6214,N_6177,N_6137);
and U6215 (N_6215,N_6181,N_6164);
xnor U6216 (N_6216,N_6130,N_6166);
and U6217 (N_6217,N_6098,N_6174);
and U6218 (N_6218,N_6089,N_6165);
or U6219 (N_6219,N_6144,N_6127);
or U6220 (N_6220,N_6040,N_6016);
or U6221 (N_6221,N_6066,N_6069);
nor U6222 (N_6222,N_6169,N_6035);
nor U6223 (N_6223,N_6184,N_6000);
nand U6224 (N_6224,N_6145,N_6091);
nor U6225 (N_6225,N_6008,N_6196);
and U6226 (N_6226,N_6139,N_6172);
nand U6227 (N_6227,N_6157,N_6160);
xor U6228 (N_6228,N_6175,N_6121);
nand U6229 (N_6229,N_6170,N_6006);
xor U6230 (N_6230,N_6168,N_6135);
or U6231 (N_6231,N_6051,N_6161);
xor U6232 (N_6232,N_6063,N_6013);
xor U6233 (N_6233,N_6136,N_6119);
nor U6234 (N_6234,N_6059,N_6140);
or U6235 (N_6235,N_6142,N_6173);
and U6236 (N_6236,N_6075,N_6005);
and U6237 (N_6237,N_6024,N_6058);
xnor U6238 (N_6238,N_6067,N_6038);
nand U6239 (N_6239,N_6106,N_6162);
nor U6240 (N_6240,N_6167,N_6050);
xor U6241 (N_6241,N_6153,N_6010);
xor U6242 (N_6242,N_6195,N_6034);
and U6243 (N_6243,N_6014,N_6001);
nor U6244 (N_6244,N_6105,N_6156);
nand U6245 (N_6245,N_6122,N_6128);
or U6246 (N_6246,N_6094,N_6012);
nor U6247 (N_6247,N_6129,N_6049);
and U6248 (N_6248,N_6041,N_6102);
and U6249 (N_6249,N_6068,N_6159);
nand U6250 (N_6250,N_6133,N_6093);
and U6251 (N_6251,N_6047,N_6043);
nand U6252 (N_6252,N_6055,N_6062);
or U6253 (N_6253,N_6183,N_6061);
or U6254 (N_6254,N_6101,N_6120);
or U6255 (N_6255,N_6103,N_6107);
or U6256 (N_6256,N_6025,N_6198);
nor U6257 (N_6257,N_6116,N_6096);
and U6258 (N_6258,N_6163,N_6048);
and U6259 (N_6259,N_6185,N_6143);
nor U6260 (N_6260,N_6045,N_6019);
xnor U6261 (N_6261,N_6110,N_6018);
nor U6262 (N_6262,N_6109,N_6124);
and U6263 (N_6263,N_6065,N_6149);
xor U6264 (N_6264,N_6125,N_6070);
nor U6265 (N_6265,N_6064,N_6123);
or U6266 (N_6266,N_6134,N_6017);
xnor U6267 (N_6267,N_6042,N_6118);
xnor U6268 (N_6268,N_6176,N_6020);
or U6269 (N_6269,N_6197,N_6148);
nor U6270 (N_6270,N_6192,N_6154);
nand U6271 (N_6271,N_6044,N_6117);
nand U6272 (N_6272,N_6052,N_6108);
or U6273 (N_6273,N_6092,N_6083);
xor U6274 (N_6274,N_6115,N_6079);
xor U6275 (N_6275,N_6054,N_6031);
nand U6276 (N_6276,N_6060,N_6189);
nand U6277 (N_6277,N_6194,N_6026);
and U6278 (N_6278,N_6152,N_6009);
or U6279 (N_6279,N_6104,N_6199);
xnor U6280 (N_6280,N_6028,N_6076);
or U6281 (N_6281,N_6077,N_6081);
and U6282 (N_6282,N_6138,N_6023);
nand U6283 (N_6283,N_6151,N_6112);
xor U6284 (N_6284,N_6190,N_6030);
nor U6285 (N_6285,N_6011,N_6179);
or U6286 (N_6286,N_6191,N_6147);
or U6287 (N_6287,N_6084,N_6003);
nor U6288 (N_6288,N_6090,N_6141);
nor U6289 (N_6289,N_6046,N_6027);
xnor U6290 (N_6290,N_6085,N_6057);
nor U6291 (N_6291,N_6131,N_6113);
or U6292 (N_6292,N_6187,N_6086);
xor U6293 (N_6293,N_6004,N_6097);
or U6294 (N_6294,N_6193,N_6126);
nand U6295 (N_6295,N_6100,N_6053);
or U6296 (N_6296,N_6171,N_6036);
and U6297 (N_6297,N_6111,N_6015);
or U6298 (N_6298,N_6056,N_6155);
xnor U6299 (N_6299,N_6087,N_6099);
and U6300 (N_6300,N_6066,N_6129);
nand U6301 (N_6301,N_6198,N_6084);
nand U6302 (N_6302,N_6161,N_6068);
or U6303 (N_6303,N_6020,N_6028);
and U6304 (N_6304,N_6037,N_6087);
xnor U6305 (N_6305,N_6022,N_6015);
nand U6306 (N_6306,N_6142,N_6171);
or U6307 (N_6307,N_6070,N_6072);
or U6308 (N_6308,N_6082,N_6026);
and U6309 (N_6309,N_6116,N_6136);
nand U6310 (N_6310,N_6105,N_6174);
or U6311 (N_6311,N_6154,N_6014);
xor U6312 (N_6312,N_6048,N_6018);
nand U6313 (N_6313,N_6107,N_6143);
nand U6314 (N_6314,N_6147,N_6050);
nand U6315 (N_6315,N_6018,N_6106);
or U6316 (N_6316,N_6025,N_6104);
or U6317 (N_6317,N_6044,N_6029);
or U6318 (N_6318,N_6141,N_6178);
and U6319 (N_6319,N_6059,N_6021);
xnor U6320 (N_6320,N_6154,N_6056);
nor U6321 (N_6321,N_6064,N_6146);
and U6322 (N_6322,N_6095,N_6146);
and U6323 (N_6323,N_6175,N_6131);
or U6324 (N_6324,N_6007,N_6104);
and U6325 (N_6325,N_6103,N_6056);
nand U6326 (N_6326,N_6034,N_6078);
or U6327 (N_6327,N_6139,N_6033);
nor U6328 (N_6328,N_6185,N_6007);
nor U6329 (N_6329,N_6164,N_6196);
nor U6330 (N_6330,N_6150,N_6154);
nor U6331 (N_6331,N_6116,N_6010);
or U6332 (N_6332,N_6072,N_6103);
or U6333 (N_6333,N_6030,N_6102);
xnor U6334 (N_6334,N_6104,N_6177);
xor U6335 (N_6335,N_6036,N_6190);
nand U6336 (N_6336,N_6057,N_6033);
xnor U6337 (N_6337,N_6079,N_6178);
or U6338 (N_6338,N_6061,N_6093);
xnor U6339 (N_6339,N_6035,N_6183);
xor U6340 (N_6340,N_6142,N_6062);
and U6341 (N_6341,N_6197,N_6033);
or U6342 (N_6342,N_6101,N_6050);
nor U6343 (N_6343,N_6064,N_6055);
or U6344 (N_6344,N_6191,N_6140);
or U6345 (N_6345,N_6162,N_6151);
or U6346 (N_6346,N_6076,N_6019);
xnor U6347 (N_6347,N_6022,N_6032);
nor U6348 (N_6348,N_6061,N_6139);
xor U6349 (N_6349,N_6107,N_6004);
or U6350 (N_6350,N_6193,N_6188);
nor U6351 (N_6351,N_6093,N_6079);
or U6352 (N_6352,N_6172,N_6065);
xor U6353 (N_6353,N_6103,N_6151);
nor U6354 (N_6354,N_6072,N_6077);
xor U6355 (N_6355,N_6029,N_6178);
nand U6356 (N_6356,N_6152,N_6057);
xor U6357 (N_6357,N_6142,N_6190);
nor U6358 (N_6358,N_6077,N_6059);
and U6359 (N_6359,N_6133,N_6079);
xnor U6360 (N_6360,N_6114,N_6074);
xnor U6361 (N_6361,N_6101,N_6029);
and U6362 (N_6362,N_6155,N_6044);
nand U6363 (N_6363,N_6155,N_6158);
and U6364 (N_6364,N_6042,N_6178);
xor U6365 (N_6365,N_6100,N_6142);
or U6366 (N_6366,N_6086,N_6049);
xor U6367 (N_6367,N_6173,N_6175);
xor U6368 (N_6368,N_6014,N_6172);
xor U6369 (N_6369,N_6118,N_6125);
or U6370 (N_6370,N_6177,N_6000);
xnor U6371 (N_6371,N_6198,N_6154);
xnor U6372 (N_6372,N_6114,N_6049);
and U6373 (N_6373,N_6008,N_6178);
nand U6374 (N_6374,N_6145,N_6099);
nand U6375 (N_6375,N_6113,N_6149);
nand U6376 (N_6376,N_6171,N_6002);
nor U6377 (N_6377,N_6147,N_6193);
xor U6378 (N_6378,N_6106,N_6197);
and U6379 (N_6379,N_6035,N_6094);
nand U6380 (N_6380,N_6120,N_6004);
xnor U6381 (N_6381,N_6005,N_6043);
xor U6382 (N_6382,N_6095,N_6189);
and U6383 (N_6383,N_6007,N_6005);
nor U6384 (N_6384,N_6051,N_6092);
nor U6385 (N_6385,N_6048,N_6056);
and U6386 (N_6386,N_6009,N_6025);
and U6387 (N_6387,N_6164,N_6141);
or U6388 (N_6388,N_6050,N_6089);
and U6389 (N_6389,N_6014,N_6132);
and U6390 (N_6390,N_6098,N_6074);
and U6391 (N_6391,N_6169,N_6026);
xnor U6392 (N_6392,N_6066,N_6079);
and U6393 (N_6393,N_6194,N_6134);
or U6394 (N_6394,N_6147,N_6086);
xnor U6395 (N_6395,N_6099,N_6197);
and U6396 (N_6396,N_6150,N_6091);
nand U6397 (N_6397,N_6025,N_6180);
nor U6398 (N_6398,N_6155,N_6129);
and U6399 (N_6399,N_6160,N_6168);
xnor U6400 (N_6400,N_6353,N_6322);
xor U6401 (N_6401,N_6246,N_6315);
nand U6402 (N_6402,N_6241,N_6203);
nor U6403 (N_6403,N_6300,N_6327);
nor U6404 (N_6404,N_6253,N_6235);
nor U6405 (N_6405,N_6399,N_6341);
or U6406 (N_6406,N_6369,N_6359);
nor U6407 (N_6407,N_6375,N_6320);
nor U6408 (N_6408,N_6220,N_6256);
or U6409 (N_6409,N_6397,N_6204);
and U6410 (N_6410,N_6384,N_6213);
or U6411 (N_6411,N_6283,N_6263);
and U6412 (N_6412,N_6243,N_6351);
or U6413 (N_6413,N_6393,N_6388);
or U6414 (N_6414,N_6303,N_6221);
nand U6415 (N_6415,N_6358,N_6367);
nor U6416 (N_6416,N_6216,N_6211);
nor U6417 (N_6417,N_6293,N_6391);
nand U6418 (N_6418,N_6270,N_6224);
and U6419 (N_6419,N_6350,N_6336);
or U6420 (N_6420,N_6311,N_6222);
nor U6421 (N_6421,N_6390,N_6288);
nand U6422 (N_6422,N_6290,N_6208);
or U6423 (N_6423,N_6289,N_6250);
nor U6424 (N_6424,N_6282,N_6240);
and U6425 (N_6425,N_6279,N_6245);
nand U6426 (N_6426,N_6339,N_6382);
xnor U6427 (N_6427,N_6317,N_6378);
nand U6428 (N_6428,N_6330,N_6343);
nand U6429 (N_6429,N_6249,N_6340);
or U6430 (N_6430,N_6305,N_6365);
xor U6431 (N_6431,N_6362,N_6278);
and U6432 (N_6432,N_6325,N_6307);
nand U6433 (N_6433,N_6364,N_6247);
nand U6434 (N_6434,N_6366,N_6242);
nor U6435 (N_6435,N_6271,N_6266);
and U6436 (N_6436,N_6296,N_6237);
nor U6437 (N_6437,N_6318,N_6226);
nor U6438 (N_6438,N_6294,N_6381);
nor U6439 (N_6439,N_6217,N_6370);
or U6440 (N_6440,N_6298,N_6349);
xor U6441 (N_6441,N_6209,N_6234);
xnor U6442 (N_6442,N_6261,N_6308);
or U6443 (N_6443,N_6262,N_6368);
and U6444 (N_6444,N_6200,N_6206);
or U6445 (N_6445,N_6342,N_6387);
xor U6446 (N_6446,N_6332,N_6324);
xnor U6447 (N_6447,N_6306,N_6386);
nor U6448 (N_6448,N_6372,N_6233);
xor U6449 (N_6449,N_6319,N_6285);
nor U6450 (N_6450,N_6223,N_6281);
or U6451 (N_6451,N_6361,N_6329);
and U6452 (N_6452,N_6238,N_6265);
nand U6453 (N_6453,N_6335,N_6272);
or U6454 (N_6454,N_6257,N_6210);
nand U6455 (N_6455,N_6310,N_6302);
or U6456 (N_6456,N_6299,N_6225);
nand U6457 (N_6457,N_6385,N_6344);
and U6458 (N_6458,N_6248,N_6356);
nand U6459 (N_6459,N_6346,N_6218);
nand U6460 (N_6460,N_6323,N_6316);
nand U6461 (N_6461,N_6328,N_6398);
nor U6462 (N_6462,N_6355,N_6314);
and U6463 (N_6463,N_6352,N_6373);
or U6464 (N_6464,N_6260,N_6331);
nor U6465 (N_6465,N_6392,N_6227);
xnor U6466 (N_6466,N_6239,N_6371);
xor U6467 (N_6467,N_6276,N_6277);
xnor U6468 (N_6468,N_6333,N_6259);
or U6469 (N_6469,N_6347,N_6252);
and U6470 (N_6470,N_6377,N_6202);
and U6471 (N_6471,N_6251,N_6207);
nor U6472 (N_6472,N_6360,N_6338);
nor U6473 (N_6473,N_6254,N_6396);
xnor U6474 (N_6474,N_6354,N_6376);
xor U6475 (N_6475,N_6232,N_6212);
or U6476 (N_6476,N_6297,N_6379);
nand U6477 (N_6477,N_6287,N_6295);
nand U6478 (N_6478,N_6301,N_6214);
nand U6479 (N_6479,N_6229,N_6255);
nor U6480 (N_6480,N_6205,N_6334);
and U6481 (N_6481,N_6236,N_6275);
nand U6482 (N_6482,N_6274,N_6291);
nor U6483 (N_6483,N_6348,N_6267);
xor U6484 (N_6484,N_6312,N_6284);
or U6485 (N_6485,N_6326,N_6394);
xnor U6486 (N_6486,N_6273,N_6280);
nor U6487 (N_6487,N_6374,N_6264);
xnor U6488 (N_6488,N_6230,N_6309);
nand U6489 (N_6489,N_6286,N_6321);
nand U6490 (N_6490,N_6389,N_6258);
nand U6491 (N_6491,N_6269,N_6201);
or U6492 (N_6492,N_6345,N_6304);
or U6493 (N_6493,N_6219,N_6228);
xnor U6494 (N_6494,N_6357,N_6292);
xor U6495 (N_6495,N_6313,N_6215);
nand U6496 (N_6496,N_6383,N_6244);
or U6497 (N_6497,N_6395,N_6231);
xnor U6498 (N_6498,N_6363,N_6337);
or U6499 (N_6499,N_6268,N_6380);
nand U6500 (N_6500,N_6254,N_6226);
and U6501 (N_6501,N_6345,N_6263);
nor U6502 (N_6502,N_6345,N_6383);
nand U6503 (N_6503,N_6278,N_6377);
nor U6504 (N_6504,N_6242,N_6201);
or U6505 (N_6505,N_6260,N_6209);
xor U6506 (N_6506,N_6228,N_6225);
nand U6507 (N_6507,N_6205,N_6316);
xnor U6508 (N_6508,N_6213,N_6293);
and U6509 (N_6509,N_6395,N_6309);
and U6510 (N_6510,N_6293,N_6397);
and U6511 (N_6511,N_6299,N_6332);
nand U6512 (N_6512,N_6329,N_6241);
and U6513 (N_6513,N_6252,N_6285);
xor U6514 (N_6514,N_6374,N_6299);
and U6515 (N_6515,N_6249,N_6233);
nand U6516 (N_6516,N_6286,N_6269);
nand U6517 (N_6517,N_6399,N_6332);
and U6518 (N_6518,N_6376,N_6310);
or U6519 (N_6519,N_6365,N_6219);
xor U6520 (N_6520,N_6248,N_6347);
nand U6521 (N_6521,N_6393,N_6327);
xor U6522 (N_6522,N_6259,N_6319);
xor U6523 (N_6523,N_6278,N_6387);
nor U6524 (N_6524,N_6368,N_6373);
and U6525 (N_6525,N_6308,N_6294);
xor U6526 (N_6526,N_6218,N_6366);
nand U6527 (N_6527,N_6306,N_6379);
nor U6528 (N_6528,N_6271,N_6395);
xor U6529 (N_6529,N_6366,N_6328);
nor U6530 (N_6530,N_6341,N_6294);
nor U6531 (N_6531,N_6243,N_6241);
xor U6532 (N_6532,N_6290,N_6281);
xor U6533 (N_6533,N_6250,N_6396);
or U6534 (N_6534,N_6387,N_6334);
nor U6535 (N_6535,N_6343,N_6258);
and U6536 (N_6536,N_6300,N_6220);
nor U6537 (N_6537,N_6360,N_6315);
or U6538 (N_6538,N_6258,N_6293);
and U6539 (N_6539,N_6334,N_6309);
and U6540 (N_6540,N_6288,N_6254);
or U6541 (N_6541,N_6377,N_6329);
and U6542 (N_6542,N_6261,N_6327);
nand U6543 (N_6543,N_6386,N_6216);
and U6544 (N_6544,N_6375,N_6214);
xnor U6545 (N_6545,N_6354,N_6360);
or U6546 (N_6546,N_6236,N_6346);
nor U6547 (N_6547,N_6233,N_6218);
xor U6548 (N_6548,N_6318,N_6223);
or U6549 (N_6549,N_6323,N_6384);
nand U6550 (N_6550,N_6322,N_6395);
and U6551 (N_6551,N_6212,N_6357);
nand U6552 (N_6552,N_6208,N_6399);
nor U6553 (N_6553,N_6291,N_6380);
nand U6554 (N_6554,N_6385,N_6209);
or U6555 (N_6555,N_6208,N_6345);
xor U6556 (N_6556,N_6364,N_6272);
or U6557 (N_6557,N_6330,N_6256);
or U6558 (N_6558,N_6356,N_6224);
xnor U6559 (N_6559,N_6332,N_6278);
nand U6560 (N_6560,N_6294,N_6221);
or U6561 (N_6561,N_6326,N_6303);
xor U6562 (N_6562,N_6236,N_6381);
or U6563 (N_6563,N_6228,N_6299);
nand U6564 (N_6564,N_6386,N_6365);
nand U6565 (N_6565,N_6248,N_6210);
nor U6566 (N_6566,N_6273,N_6259);
or U6567 (N_6567,N_6299,N_6310);
xnor U6568 (N_6568,N_6343,N_6235);
xnor U6569 (N_6569,N_6369,N_6353);
or U6570 (N_6570,N_6227,N_6374);
nand U6571 (N_6571,N_6272,N_6255);
nor U6572 (N_6572,N_6248,N_6359);
or U6573 (N_6573,N_6241,N_6386);
and U6574 (N_6574,N_6300,N_6223);
nand U6575 (N_6575,N_6363,N_6222);
xor U6576 (N_6576,N_6297,N_6208);
or U6577 (N_6577,N_6302,N_6273);
xnor U6578 (N_6578,N_6345,N_6265);
or U6579 (N_6579,N_6224,N_6253);
and U6580 (N_6580,N_6258,N_6338);
or U6581 (N_6581,N_6391,N_6274);
nand U6582 (N_6582,N_6246,N_6276);
nor U6583 (N_6583,N_6229,N_6318);
and U6584 (N_6584,N_6397,N_6346);
and U6585 (N_6585,N_6204,N_6313);
nand U6586 (N_6586,N_6233,N_6323);
nor U6587 (N_6587,N_6387,N_6245);
nand U6588 (N_6588,N_6221,N_6261);
and U6589 (N_6589,N_6212,N_6247);
nor U6590 (N_6590,N_6300,N_6230);
nand U6591 (N_6591,N_6368,N_6232);
nand U6592 (N_6592,N_6280,N_6235);
nand U6593 (N_6593,N_6286,N_6363);
nor U6594 (N_6594,N_6228,N_6293);
nand U6595 (N_6595,N_6246,N_6236);
nor U6596 (N_6596,N_6385,N_6329);
and U6597 (N_6597,N_6372,N_6288);
nand U6598 (N_6598,N_6306,N_6249);
nor U6599 (N_6599,N_6280,N_6376);
nand U6600 (N_6600,N_6536,N_6426);
xor U6601 (N_6601,N_6478,N_6555);
nor U6602 (N_6602,N_6576,N_6550);
nor U6603 (N_6603,N_6499,N_6533);
nand U6604 (N_6604,N_6534,N_6589);
xor U6605 (N_6605,N_6583,N_6543);
xor U6606 (N_6606,N_6520,N_6516);
and U6607 (N_6607,N_6595,N_6406);
xnor U6608 (N_6608,N_6505,N_6409);
nor U6609 (N_6609,N_6491,N_6472);
nand U6610 (N_6610,N_6445,N_6525);
nand U6611 (N_6611,N_6489,N_6532);
xnor U6612 (N_6612,N_6514,N_6560);
nor U6613 (N_6613,N_6462,N_6488);
or U6614 (N_6614,N_6542,N_6561);
and U6615 (N_6615,N_6578,N_6402);
nor U6616 (N_6616,N_6457,N_6461);
nand U6617 (N_6617,N_6582,N_6537);
nor U6618 (N_6618,N_6401,N_6590);
xor U6619 (N_6619,N_6574,N_6530);
and U6620 (N_6620,N_6449,N_6470);
nand U6621 (N_6621,N_6458,N_6413);
and U6622 (N_6622,N_6587,N_6544);
nand U6623 (N_6623,N_6511,N_6498);
nand U6624 (N_6624,N_6464,N_6454);
or U6625 (N_6625,N_6535,N_6580);
nor U6626 (N_6626,N_6492,N_6513);
nand U6627 (N_6627,N_6549,N_6418);
xnor U6628 (N_6628,N_6540,N_6442);
nand U6629 (N_6629,N_6419,N_6433);
nand U6630 (N_6630,N_6456,N_6452);
nand U6631 (N_6631,N_6509,N_6485);
nand U6632 (N_6632,N_6477,N_6403);
nand U6633 (N_6633,N_6483,N_6588);
nand U6634 (N_6634,N_6577,N_6476);
nor U6635 (N_6635,N_6437,N_6547);
and U6636 (N_6636,N_6439,N_6598);
xor U6637 (N_6637,N_6551,N_6482);
nand U6638 (N_6638,N_6429,N_6453);
and U6639 (N_6639,N_6591,N_6436);
xnor U6640 (N_6640,N_6424,N_6447);
nor U6641 (N_6641,N_6440,N_6572);
nand U6642 (N_6642,N_6430,N_6484);
nor U6643 (N_6643,N_6480,N_6428);
or U6644 (N_6644,N_6473,N_6460);
nand U6645 (N_6645,N_6558,N_6404);
nor U6646 (N_6646,N_6508,N_6412);
nor U6647 (N_6647,N_6579,N_6502);
and U6648 (N_6648,N_6407,N_6474);
and U6649 (N_6649,N_6500,N_6564);
or U6650 (N_6650,N_6575,N_6567);
nand U6651 (N_6651,N_6446,N_6501);
and U6652 (N_6652,N_6400,N_6538);
xor U6653 (N_6653,N_6545,N_6573);
or U6654 (N_6654,N_6497,N_6463);
xnor U6655 (N_6655,N_6548,N_6469);
and U6656 (N_6656,N_6569,N_6512);
nor U6657 (N_6657,N_6443,N_6597);
or U6658 (N_6658,N_6566,N_6565);
or U6659 (N_6659,N_6559,N_6475);
nand U6660 (N_6660,N_6531,N_6425);
xnor U6661 (N_6661,N_6459,N_6570);
nand U6662 (N_6662,N_6450,N_6571);
nand U6663 (N_6663,N_6504,N_6556);
nand U6664 (N_6664,N_6427,N_6432);
and U6665 (N_6665,N_6416,N_6455);
xor U6666 (N_6666,N_6529,N_6467);
and U6667 (N_6667,N_6562,N_6546);
nand U6668 (N_6668,N_6493,N_6506);
nor U6669 (N_6669,N_6466,N_6405);
nor U6670 (N_6670,N_6522,N_6557);
or U6671 (N_6671,N_6408,N_6584);
or U6672 (N_6672,N_6441,N_6496);
xor U6673 (N_6673,N_6420,N_6594);
or U6674 (N_6674,N_6431,N_6495);
and U6675 (N_6675,N_6448,N_6423);
and U6676 (N_6676,N_6411,N_6528);
or U6677 (N_6677,N_6414,N_6465);
nand U6678 (N_6678,N_6486,N_6518);
or U6679 (N_6679,N_6494,N_6585);
or U6680 (N_6680,N_6415,N_6422);
and U6681 (N_6681,N_6521,N_6526);
xnor U6682 (N_6682,N_6438,N_6487);
nand U6683 (N_6683,N_6524,N_6596);
xnor U6684 (N_6684,N_6527,N_6417);
nor U6685 (N_6685,N_6593,N_6410);
nor U6686 (N_6686,N_6421,N_6553);
nor U6687 (N_6687,N_6599,N_6581);
or U6688 (N_6688,N_6554,N_6434);
and U6689 (N_6689,N_6541,N_6523);
nand U6690 (N_6690,N_6539,N_6586);
nor U6691 (N_6691,N_6552,N_6451);
nand U6692 (N_6692,N_6503,N_6481);
and U6693 (N_6693,N_6519,N_6515);
and U6694 (N_6694,N_6435,N_6471);
and U6695 (N_6695,N_6563,N_6490);
xnor U6696 (N_6696,N_6507,N_6444);
and U6697 (N_6697,N_6568,N_6468);
and U6698 (N_6698,N_6592,N_6479);
and U6699 (N_6699,N_6510,N_6517);
nor U6700 (N_6700,N_6401,N_6539);
or U6701 (N_6701,N_6512,N_6483);
xnor U6702 (N_6702,N_6560,N_6445);
or U6703 (N_6703,N_6570,N_6436);
and U6704 (N_6704,N_6562,N_6475);
nor U6705 (N_6705,N_6486,N_6455);
and U6706 (N_6706,N_6557,N_6545);
nand U6707 (N_6707,N_6575,N_6590);
or U6708 (N_6708,N_6415,N_6540);
or U6709 (N_6709,N_6404,N_6468);
nand U6710 (N_6710,N_6564,N_6456);
and U6711 (N_6711,N_6468,N_6478);
xor U6712 (N_6712,N_6431,N_6595);
and U6713 (N_6713,N_6404,N_6472);
nor U6714 (N_6714,N_6417,N_6587);
or U6715 (N_6715,N_6517,N_6511);
nor U6716 (N_6716,N_6569,N_6520);
or U6717 (N_6717,N_6432,N_6568);
or U6718 (N_6718,N_6512,N_6567);
xor U6719 (N_6719,N_6571,N_6579);
xnor U6720 (N_6720,N_6439,N_6449);
xnor U6721 (N_6721,N_6580,N_6531);
and U6722 (N_6722,N_6549,N_6533);
or U6723 (N_6723,N_6433,N_6403);
xnor U6724 (N_6724,N_6589,N_6441);
and U6725 (N_6725,N_6577,N_6458);
or U6726 (N_6726,N_6436,N_6481);
nor U6727 (N_6727,N_6413,N_6472);
nor U6728 (N_6728,N_6541,N_6538);
xnor U6729 (N_6729,N_6488,N_6445);
xor U6730 (N_6730,N_6568,N_6552);
and U6731 (N_6731,N_6427,N_6549);
nor U6732 (N_6732,N_6595,N_6487);
nor U6733 (N_6733,N_6468,N_6461);
nor U6734 (N_6734,N_6455,N_6531);
or U6735 (N_6735,N_6510,N_6402);
nor U6736 (N_6736,N_6567,N_6540);
nand U6737 (N_6737,N_6593,N_6400);
nor U6738 (N_6738,N_6402,N_6424);
or U6739 (N_6739,N_6513,N_6437);
nand U6740 (N_6740,N_6411,N_6401);
nor U6741 (N_6741,N_6518,N_6567);
nor U6742 (N_6742,N_6458,N_6431);
or U6743 (N_6743,N_6571,N_6531);
nand U6744 (N_6744,N_6562,N_6476);
nand U6745 (N_6745,N_6461,N_6412);
or U6746 (N_6746,N_6427,N_6469);
or U6747 (N_6747,N_6534,N_6503);
xor U6748 (N_6748,N_6417,N_6550);
nor U6749 (N_6749,N_6421,N_6429);
or U6750 (N_6750,N_6415,N_6508);
xnor U6751 (N_6751,N_6596,N_6490);
or U6752 (N_6752,N_6554,N_6506);
xor U6753 (N_6753,N_6457,N_6453);
and U6754 (N_6754,N_6498,N_6504);
or U6755 (N_6755,N_6405,N_6492);
nand U6756 (N_6756,N_6582,N_6464);
or U6757 (N_6757,N_6483,N_6473);
nand U6758 (N_6758,N_6464,N_6565);
nor U6759 (N_6759,N_6557,N_6465);
nor U6760 (N_6760,N_6429,N_6457);
or U6761 (N_6761,N_6539,N_6583);
nand U6762 (N_6762,N_6475,N_6563);
and U6763 (N_6763,N_6557,N_6445);
xnor U6764 (N_6764,N_6551,N_6438);
xor U6765 (N_6765,N_6422,N_6596);
or U6766 (N_6766,N_6468,N_6545);
nand U6767 (N_6767,N_6494,N_6531);
nor U6768 (N_6768,N_6586,N_6467);
nand U6769 (N_6769,N_6502,N_6582);
nor U6770 (N_6770,N_6590,N_6488);
nor U6771 (N_6771,N_6474,N_6442);
and U6772 (N_6772,N_6463,N_6532);
nor U6773 (N_6773,N_6493,N_6456);
or U6774 (N_6774,N_6447,N_6552);
or U6775 (N_6775,N_6566,N_6493);
or U6776 (N_6776,N_6402,N_6457);
nand U6777 (N_6777,N_6474,N_6488);
nor U6778 (N_6778,N_6493,N_6466);
nor U6779 (N_6779,N_6450,N_6594);
nand U6780 (N_6780,N_6434,N_6552);
nand U6781 (N_6781,N_6583,N_6555);
nand U6782 (N_6782,N_6550,N_6411);
nand U6783 (N_6783,N_6589,N_6595);
nand U6784 (N_6784,N_6515,N_6528);
and U6785 (N_6785,N_6440,N_6524);
and U6786 (N_6786,N_6506,N_6427);
nand U6787 (N_6787,N_6590,N_6402);
nand U6788 (N_6788,N_6491,N_6455);
nand U6789 (N_6789,N_6533,N_6571);
xor U6790 (N_6790,N_6499,N_6580);
xnor U6791 (N_6791,N_6513,N_6540);
nor U6792 (N_6792,N_6462,N_6436);
nor U6793 (N_6793,N_6514,N_6583);
nor U6794 (N_6794,N_6581,N_6480);
nand U6795 (N_6795,N_6434,N_6448);
xor U6796 (N_6796,N_6519,N_6427);
or U6797 (N_6797,N_6494,N_6421);
or U6798 (N_6798,N_6598,N_6554);
nor U6799 (N_6799,N_6580,N_6541);
or U6800 (N_6800,N_6747,N_6704);
and U6801 (N_6801,N_6653,N_6610);
and U6802 (N_6802,N_6667,N_6632);
or U6803 (N_6803,N_6606,N_6677);
nand U6804 (N_6804,N_6627,N_6728);
or U6805 (N_6805,N_6714,N_6613);
and U6806 (N_6806,N_6731,N_6718);
nand U6807 (N_6807,N_6797,N_6776);
nor U6808 (N_6808,N_6643,N_6641);
or U6809 (N_6809,N_6622,N_6758);
nand U6810 (N_6810,N_6692,N_6735);
xor U6811 (N_6811,N_6699,N_6717);
or U6812 (N_6812,N_6799,N_6617);
or U6813 (N_6813,N_6742,N_6697);
or U6814 (N_6814,N_6788,N_6631);
and U6815 (N_6815,N_6765,N_6734);
and U6816 (N_6816,N_6630,N_6693);
nand U6817 (N_6817,N_6674,N_6701);
xnor U6818 (N_6818,N_6795,N_6766);
xor U6819 (N_6819,N_6737,N_6736);
xnor U6820 (N_6820,N_6726,N_6778);
or U6821 (N_6821,N_6796,N_6724);
nand U6822 (N_6822,N_6761,N_6725);
nand U6823 (N_6823,N_6789,N_6713);
or U6824 (N_6824,N_6652,N_6715);
or U6825 (N_6825,N_6741,N_6794);
and U6826 (N_6826,N_6666,N_6780);
nor U6827 (N_6827,N_6764,N_6785);
and U6828 (N_6828,N_6711,N_6683);
nand U6829 (N_6829,N_6635,N_6675);
or U6830 (N_6830,N_6688,N_6782);
or U6831 (N_6831,N_6791,N_6605);
and U6832 (N_6832,N_6609,N_6660);
nor U6833 (N_6833,N_6712,N_6706);
and U6834 (N_6834,N_6775,N_6696);
or U6835 (N_6835,N_6619,N_6618);
and U6836 (N_6836,N_6753,N_6739);
and U6837 (N_6837,N_6624,N_6769);
or U6838 (N_6838,N_6680,N_6691);
nand U6839 (N_6839,N_6751,N_6777);
or U6840 (N_6840,N_6602,N_6626);
and U6841 (N_6841,N_6685,N_6729);
or U6842 (N_6842,N_6774,N_6621);
or U6843 (N_6843,N_6673,N_6798);
and U6844 (N_6844,N_6640,N_6601);
and U6845 (N_6845,N_6604,N_6738);
nor U6846 (N_6846,N_6745,N_6615);
and U6847 (N_6847,N_6665,N_6750);
xnor U6848 (N_6848,N_6642,N_6676);
nor U6849 (N_6849,N_6771,N_6757);
xnor U6850 (N_6850,N_6792,N_6636);
nand U6851 (N_6851,N_6648,N_6722);
and U6852 (N_6852,N_6748,N_6709);
or U6853 (N_6853,N_6721,N_6607);
xor U6854 (N_6854,N_6781,N_6754);
xnor U6855 (N_6855,N_6787,N_6708);
nor U6856 (N_6856,N_6698,N_6679);
xor U6857 (N_6857,N_6756,N_6629);
xnor U6858 (N_6858,N_6694,N_6655);
and U6859 (N_6859,N_6662,N_6647);
and U6860 (N_6860,N_6637,N_6730);
and U6861 (N_6861,N_6689,N_6657);
xor U6862 (N_6862,N_6723,N_6614);
nand U6863 (N_6863,N_6650,N_6740);
xnor U6864 (N_6864,N_6710,N_6681);
or U6865 (N_6865,N_6658,N_6608);
nor U6866 (N_6866,N_6633,N_6623);
xor U6867 (N_6867,N_6793,N_6611);
xnor U6868 (N_6868,N_6744,N_6763);
nand U6869 (N_6869,N_6671,N_6670);
or U6870 (N_6870,N_6646,N_6634);
and U6871 (N_6871,N_6755,N_6702);
xnor U6872 (N_6872,N_6684,N_6727);
nand U6873 (N_6873,N_6784,N_6656);
nand U6874 (N_6874,N_6659,N_6603);
nor U6875 (N_6875,N_6686,N_6651);
nand U6876 (N_6876,N_6687,N_6638);
or U6877 (N_6877,N_6649,N_6625);
nand U6878 (N_6878,N_6644,N_6762);
nand U6879 (N_6879,N_6672,N_6733);
or U6880 (N_6880,N_6695,N_6669);
or U6881 (N_6881,N_6783,N_6716);
and U6882 (N_6882,N_6749,N_6690);
nor U6883 (N_6883,N_6720,N_6668);
nor U6884 (N_6884,N_6700,N_6746);
or U6885 (N_6885,N_6732,N_6620);
or U6886 (N_6886,N_6663,N_6703);
and U6887 (N_6887,N_6719,N_6616);
nand U6888 (N_6888,N_6773,N_6664);
and U6889 (N_6889,N_6759,N_6779);
nor U6890 (N_6890,N_6628,N_6645);
and U6891 (N_6891,N_6678,N_6600);
and U6892 (N_6892,N_6612,N_6682);
and U6893 (N_6893,N_6768,N_6639);
xor U6894 (N_6894,N_6661,N_6770);
and U6895 (N_6895,N_6790,N_6707);
nand U6896 (N_6896,N_6786,N_6767);
xor U6897 (N_6897,N_6743,N_6752);
xor U6898 (N_6898,N_6705,N_6654);
or U6899 (N_6899,N_6760,N_6772);
nand U6900 (N_6900,N_6653,N_6768);
nand U6901 (N_6901,N_6750,N_6747);
or U6902 (N_6902,N_6600,N_6788);
nand U6903 (N_6903,N_6674,N_6616);
or U6904 (N_6904,N_6793,N_6649);
and U6905 (N_6905,N_6715,N_6635);
xor U6906 (N_6906,N_6794,N_6742);
and U6907 (N_6907,N_6642,N_6737);
xor U6908 (N_6908,N_6767,N_6710);
and U6909 (N_6909,N_6699,N_6732);
nand U6910 (N_6910,N_6774,N_6703);
and U6911 (N_6911,N_6795,N_6722);
nand U6912 (N_6912,N_6625,N_6601);
xnor U6913 (N_6913,N_6766,N_6732);
nand U6914 (N_6914,N_6675,N_6764);
and U6915 (N_6915,N_6770,N_6671);
nand U6916 (N_6916,N_6633,N_6625);
and U6917 (N_6917,N_6741,N_6637);
or U6918 (N_6918,N_6719,N_6682);
and U6919 (N_6919,N_6752,N_6740);
xor U6920 (N_6920,N_6775,N_6603);
nor U6921 (N_6921,N_6607,N_6621);
or U6922 (N_6922,N_6785,N_6760);
nor U6923 (N_6923,N_6792,N_6734);
and U6924 (N_6924,N_6640,N_6645);
xnor U6925 (N_6925,N_6664,N_6646);
nor U6926 (N_6926,N_6787,N_6714);
nor U6927 (N_6927,N_6605,N_6709);
or U6928 (N_6928,N_6773,N_6786);
xnor U6929 (N_6929,N_6661,N_6626);
nand U6930 (N_6930,N_6767,N_6784);
nand U6931 (N_6931,N_6761,N_6741);
and U6932 (N_6932,N_6637,N_6763);
or U6933 (N_6933,N_6798,N_6799);
nand U6934 (N_6934,N_6672,N_6699);
nor U6935 (N_6935,N_6699,N_6640);
and U6936 (N_6936,N_6797,N_6675);
nor U6937 (N_6937,N_6758,N_6665);
xor U6938 (N_6938,N_6772,N_6654);
nor U6939 (N_6939,N_6782,N_6716);
xor U6940 (N_6940,N_6604,N_6688);
xor U6941 (N_6941,N_6748,N_6627);
and U6942 (N_6942,N_6690,N_6632);
and U6943 (N_6943,N_6612,N_6602);
and U6944 (N_6944,N_6607,N_6702);
nand U6945 (N_6945,N_6603,N_6762);
nor U6946 (N_6946,N_6769,N_6685);
nand U6947 (N_6947,N_6617,N_6771);
and U6948 (N_6948,N_6734,N_6713);
xnor U6949 (N_6949,N_6677,N_6714);
nor U6950 (N_6950,N_6689,N_6632);
or U6951 (N_6951,N_6780,N_6782);
xor U6952 (N_6952,N_6726,N_6719);
or U6953 (N_6953,N_6731,N_6742);
and U6954 (N_6954,N_6681,N_6682);
and U6955 (N_6955,N_6760,N_6735);
xor U6956 (N_6956,N_6786,N_6779);
nand U6957 (N_6957,N_6669,N_6762);
or U6958 (N_6958,N_6753,N_6602);
and U6959 (N_6959,N_6685,N_6743);
xnor U6960 (N_6960,N_6735,N_6780);
nor U6961 (N_6961,N_6696,N_6764);
or U6962 (N_6962,N_6624,N_6695);
nor U6963 (N_6963,N_6779,N_6704);
or U6964 (N_6964,N_6739,N_6759);
nor U6965 (N_6965,N_6727,N_6719);
xnor U6966 (N_6966,N_6733,N_6613);
nor U6967 (N_6967,N_6782,N_6794);
and U6968 (N_6968,N_6604,N_6680);
or U6969 (N_6969,N_6792,N_6621);
xnor U6970 (N_6970,N_6743,N_6610);
xor U6971 (N_6971,N_6712,N_6763);
and U6972 (N_6972,N_6725,N_6670);
nand U6973 (N_6973,N_6741,N_6626);
nor U6974 (N_6974,N_6670,N_6617);
nor U6975 (N_6975,N_6755,N_6709);
nand U6976 (N_6976,N_6742,N_6698);
nor U6977 (N_6977,N_6677,N_6662);
nand U6978 (N_6978,N_6794,N_6603);
or U6979 (N_6979,N_6608,N_6700);
nand U6980 (N_6980,N_6787,N_6772);
or U6981 (N_6981,N_6687,N_6680);
nor U6982 (N_6982,N_6609,N_6645);
xor U6983 (N_6983,N_6750,N_6664);
xnor U6984 (N_6984,N_6630,N_6781);
xnor U6985 (N_6985,N_6771,N_6731);
nand U6986 (N_6986,N_6783,N_6707);
nor U6987 (N_6987,N_6771,N_6611);
or U6988 (N_6988,N_6605,N_6664);
or U6989 (N_6989,N_6710,N_6751);
nor U6990 (N_6990,N_6620,N_6752);
or U6991 (N_6991,N_6655,N_6785);
or U6992 (N_6992,N_6678,N_6642);
or U6993 (N_6993,N_6753,N_6740);
nand U6994 (N_6994,N_6683,N_6616);
or U6995 (N_6995,N_6663,N_6688);
nand U6996 (N_6996,N_6692,N_6727);
nand U6997 (N_6997,N_6756,N_6772);
xnor U6998 (N_6998,N_6603,N_6622);
or U6999 (N_6999,N_6642,N_6777);
nand U7000 (N_7000,N_6989,N_6809);
and U7001 (N_7001,N_6992,N_6973);
nor U7002 (N_7002,N_6818,N_6832);
nor U7003 (N_7003,N_6863,N_6899);
or U7004 (N_7004,N_6949,N_6843);
and U7005 (N_7005,N_6847,N_6815);
and U7006 (N_7006,N_6962,N_6806);
nor U7007 (N_7007,N_6856,N_6984);
nor U7008 (N_7008,N_6905,N_6968);
or U7009 (N_7009,N_6998,N_6945);
nand U7010 (N_7010,N_6851,N_6862);
nand U7011 (N_7011,N_6956,N_6912);
or U7012 (N_7012,N_6914,N_6835);
nand U7013 (N_7013,N_6924,N_6950);
nor U7014 (N_7014,N_6886,N_6892);
nand U7015 (N_7015,N_6814,N_6994);
and U7016 (N_7016,N_6848,N_6879);
nand U7017 (N_7017,N_6805,N_6898);
nand U7018 (N_7018,N_6845,N_6801);
xor U7019 (N_7019,N_6907,N_6811);
and U7020 (N_7020,N_6939,N_6904);
xor U7021 (N_7021,N_6834,N_6842);
or U7022 (N_7022,N_6993,N_6824);
or U7023 (N_7023,N_6893,N_6963);
nor U7024 (N_7024,N_6854,N_6894);
nand U7025 (N_7025,N_6976,N_6958);
xor U7026 (N_7026,N_6840,N_6821);
or U7027 (N_7027,N_6867,N_6920);
nand U7028 (N_7028,N_6861,N_6868);
xnor U7029 (N_7029,N_6929,N_6891);
nor U7030 (N_7030,N_6921,N_6910);
or U7031 (N_7031,N_6810,N_6819);
xnor U7032 (N_7032,N_6951,N_6823);
nor U7033 (N_7033,N_6959,N_6838);
nand U7034 (N_7034,N_6925,N_6870);
or U7035 (N_7035,N_6908,N_6931);
nand U7036 (N_7036,N_6877,N_6941);
nand U7037 (N_7037,N_6936,N_6954);
or U7038 (N_7038,N_6919,N_6804);
xnor U7039 (N_7039,N_6928,N_6858);
or U7040 (N_7040,N_6926,N_6808);
or U7041 (N_7041,N_6999,N_6857);
xnor U7042 (N_7042,N_6930,N_6952);
nand U7043 (N_7043,N_6836,N_6915);
nor U7044 (N_7044,N_6841,N_6977);
nand U7045 (N_7045,N_6803,N_6873);
nor U7046 (N_7046,N_6943,N_6986);
or U7047 (N_7047,N_6972,N_6820);
nor U7048 (N_7048,N_6800,N_6875);
nand U7049 (N_7049,N_6935,N_6982);
and U7050 (N_7050,N_6940,N_6966);
xor U7051 (N_7051,N_6846,N_6826);
and U7052 (N_7052,N_6884,N_6866);
nand U7053 (N_7053,N_6948,N_6864);
nand U7054 (N_7054,N_6860,N_6944);
xnor U7055 (N_7055,N_6980,N_6849);
or U7056 (N_7056,N_6874,N_6997);
and U7057 (N_7057,N_6885,N_6850);
xor U7058 (N_7058,N_6991,N_6871);
nor U7059 (N_7059,N_6964,N_6917);
nor U7060 (N_7060,N_6830,N_6876);
nand U7061 (N_7061,N_6996,N_6869);
nand U7062 (N_7062,N_6937,N_6988);
and U7063 (N_7063,N_6895,N_6897);
and U7064 (N_7064,N_6922,N_6923);
and U7065 (N_7065,N_6957,N_6961);
nand U7066 (N_7066,N_6970,N_6965);
xnor U7067 (N_7067,N_6896,N_6883);
nor U7068 (N_7068,N_6932,N_6967);
and U7069 (N_7069,N_6911,N_6909);
and U7070 (N_7070,N_6983,N_6837);
nand U7071 (N_7071,N_6981,N_6816);
and U7072 (N_7072,N_6844,N_6985);
and U7073 (N_7073,N_6953,N_6974);
xor U7074 (N_7074,N_6934,N_6955);
nor U7075 (N_7075,N_6995,N_6853);
or U7076 (N_7076,N_6888,N_6825);
xor U7077 (N_7077,N_6978,N_6822);
nand U7078 (N_7078,N_6969,N_6812);
nor U7079 (N_7079,N_6831,N_6880);
nor U7080 (N_7080,N_6878,N_6906);
nor U7081 (N_7081,N_6852,N_6913);
or U7082 (N_7082,N_6987,N_6828);
xnor U7083 (N_7083,N_6933,N_6975);
or U7084 (N_7084,N_6802,N_6960);
xor U7085 (N_7085,N_6890,N_6918);
nand U7086 (N_7086,N_6900,N_6817);
and U7087 (N_7087,N_6827,N_6990);
or U7088 (N_7088,N_6916,N_6901);
and U7089 (N_7089,N_6902,N_6947);
and U7090 (N_7090,N_6881,N_6872);
nor U7091 (N_7091,N_6855,N_6859);
xor U7092 (N_7092,N_6971,N_6833);
or U7093 (N_7093,N_6979,N_6865);
or U7094 (N_7094,N_6887,N_6889);
or U7095 (N_7095,N_6829,N_6807);
xnor U7096 (N_7096,N_6938,N_6927);
nand U7097 (N_7097,N_6813,N_6942);
xor U7098 (N_7098,N_6882,N_6839);
nor U7099 (N_7099,N_6946,N_6903);
and U7100 (N_7100,N_6849,N_6858);
and U7101 (N_7101,N_6862,N_6831);
xnor U7102 (N_7102,N_6983,N_6925);
and U7103 (N_7103,N_6823,N_6890);
and U7104 (N_7104,N_6903,N_6917);
or U7105 (N_7105,N_6944,N_6886);
and U7106 (N_7106,N_6865,N_6807);
and U7107 (N_7107,N_6937,N_6914);
or U7108 (N_7108,N_6996,N_6977);
nand U7109 (N_7109,N_6902,N_6839);
xnor U7110 (N_7110,N_6841,N_6945);
or U7111 (N_7111,N_6887,N_6823);
nor U7112 (N_7112,N_6924,N_6946);
xnor U7113 (N_7113,N_6952,N_6855);
xor U7114 (N_7114,N_6941,N_6919);
nand U7115 (N_7115,N_6827,N_6893);
and U7116 (N_7116,N_6954,N_6915);
nand U7117 (N_7117,N_6903,N_6864);
or U7118 (N_7118,N_6947,N_6917);
and U7119 (N_7119,N_6977,N_6870);
nand U7120 (N_7120,N_6979,N_6853);
nor U7121 (N_7121,N_6832,N_6866);
nor U7122 (N_7122,N_6920,N_6832);
xor U7123 (N_7123,N_6981,N_6941);
or U7124 (N_7124,N_6821,N_6921);
xnor U7125 (N_7125,N_6978,N_6805);
xor U7126 (N_7126,N_6878,N_6872);
or U7127 (N_7127,N_6870,N_6847);
and U7128 (N_7128,N_6880,N_6883);
nor U7129 (N_7129,N_6915,N_6934);
nor U7130 (N_7130,N_6932,N_6890);
xnor U7131 (N_7131,N_6932,N_6868);
and U7132 (N_7132,N_6909,N_6962);
or U7133 (N_7133,N_6883,N_6862);
xnor U7134 (N_7134,N_6846,N_6992);
xor U7135 (N_7135,N_6871,N_6817);
xor U7136 (N_7136,N_6827,N_6996);
or U7137 (N_7137,N_6903,N_6956);
and U7138 (N_7138,N_6940,N_6826);
nor U7139 (N_7139,N_6991,N_6939);
and U7140 (N_7140,N_6842,N_6888);
nand U7141 (N_7141,N_6835,N_6961);
and U7142 (N_7142,N_6939,N_6831);
xnor U7143 (N_7143,N_6805,N_6963);
or U7144 (N_7144,N_6911,N_6958);
nand U7145 (N_7145,N_6953,N_6834);
xnor U7146 (N_7146,N_6902,N_6925);
nand U7147 (N_7147,N_6972,N_6807);
nor U7148 (N_7148,N_6919,N_6828);
xnor U7149 (N_7149,N_6996,N_6843);
or U7150 (N_7150,N_6845,N_6881);
and U7151 (N_7151,N_6808,N_6913);
xor U7152 (N_7152,N_6954,N_6906);
and U7153 (N_7153,N_6982,N_6971);
nand U7154 (N_7154,N_6933,N_6939);
and U7155 (N_7155,N_6930,N_6909);
nor U7156 (N_7156,N_6979,N_6882);
nand U7157 (N_7157,N_6885,N_6965);
nor U7158 (N_7158,N_6977,N_6981);
nand U7159 (N_7159,N_6991,N_6906);
nor U7160 (N_7160,N_6816,N_6918);
or U7161 (N_7161,N_6914,N_6960);
and U7162 (N_7162,N_6943,N_6808);
nor U7163 (N_7163,N_6960,N_6889);
nand U7164 (N_7164,N_6974,N_6972);
nand U7165 (N_7165,N_6964,N_6941);
nand U7166 (N_7166,N_6807,N_6826);
xnor U7167 (N_7167,N_6980,N_6968);
nand U7168 (N_7168,N_6916,N_6826);
nand U7169 (N_7169,N_6849,N_6846);
nand U7170 (N_7170,N_6921,N_6876);
nand U7171 (N_7171,N_6972,N_6983);
xnor U7172 (N_7172,N_6922,N_6855);
or U7173 (N_7173,N_6998,N_6837);
or U7174 (N_7174,N_6876,N_6987);
xnor U7175 (N_7175,N_6968,N_6987);
nor U7176 (N_7176,N_6927,N_6945);
nand U7177 (N_7177,N_6971,N_6964);
nor U7178 (N_7178,N_6990,N_6813);
and U7179 (N_7179,N_6889,N_6900);
or U7180 (N_7180,N_6986,N_6859);
or U7181 (N_7181,N_6910,N_6952);
and U7182 (N_7182,N_6843,N_6907);
xnor U7183 (N_7183,N_6973,N_6824);
nand U7184 (N_7184,N_6985,N_6966);
or U7185 (N_7185,N_6933,N_6842);
nand U7186 (N_7186,N_6865,N_6841);
or U7187 (N_7187,N_6894,N_6815);
nand U7188 (N_7188,N_6851,N_6864);
xor U7189 (N_7189,N_6869,N_6947);
or U7190 (N_7190,N_6816,N_6835);
xnor U7191 (N_7191,N_6841,N_6842);
and U7192 (N_7192,N_6931,N_6819);
nor U7193 (N_7193,N_6909,N_6830);
nor U7194 (N_7194,N_6850,N_6906);
nand U7195 (N_7195,N_6952,N_6840);
or U7196 (N_7196,N_6947,N_6853);
and U7197 (N_7197,N_6837,N_6839);
nor U7198 (N_7198,N_6927,N_6904);
and U7199 (N_7199,N_6850,N_6980);
nor U7200 (N_7200,N_7063,N_7186);
nand U7201 (N_7201,N_7035,N_7144);
xor U7202 (N_7202,N_7092,N_7046);
nor U7203 (N_7203,N_7165,N_7169);
nand U7204 (N_7204,N_7051,N_7173);
nor U7205 (N_7205,N_7161,N_7196);
or U7206 (N_7206,N_7053,N_7026);
nor U7207 (N_7207,N_7099,N_7020);
and U7208 (N_7208,N_7137,N_7023);
nand U7209 (N_7209,N_7138,N_7012);
xnor U7210 (N_7210,N_7016,N_7094);
xor U7211 (N_7211,N_7000,N_7059);
nand U7212 (N_7212,N_7128,N_7028);
nand U7213 (N_7213,N_7153,N_7139);
nor U7214 (N_7214,N_7154,N_7033);
and U7215 (N_7215,N_7038,N_7042);
or U7216 (N_7216,N_7197,N_7034);
and U7217 (N_7217,N_7022,N_7057);
and U7218 (N_7218,N_7002,N_7132);
nor U7219 (N_7219,N_7114,N_7080);
nor U7220 (N_7220,N_7071,N_7179);
xnor U7221 (N_7221,N_7006,N_7069);
nor U7222 (N_7222,N_7019,N_7001);
or U7223 (N_7223,N_7040,N_7047);
nor U7224 (N_7224,N_7077,N_7118);
and U7225 (N_7225,N_7088,N_7090);
nand U7226 (N_7226,N_7122,N_7079);
or U7227 (N_7227,N_7108,N_7003);
xnor U7228 (N_7228,N_7013,N_7120);
xnor U7229 (N_7229,N_7131,N_7146);
nor U7230 (N_7230,N_7182,N_7198);
or U7231 (N_7231,N_7184,N_7039);
or U7232 (N_7232,N_7098,N_7104);
and U7233 (N_7233,N_7109,N_7135);
nor U7234 (N_7234,N_7081,N_7149);
nor U7235 (N_7235,N_7005,N_7036);
nor U7236 (N_7236,N_7067,N_7102);
nor U7237 (N_7237,N_7141,N_7155);
and U7238 (N_7238,N_7060,N_7097);
or U7239 (N_7239,N_7043,N_7119);
or U7240 (N_7240,N_7085,N_7084);
xor U7241 (N_7241,N_7107,N_7160);
xnor U7242 (N_7242,N_7152,N_7070);
nor U7243 (N_7243,N_7130,N_7110);
nor U7244 (N_7244,N_7192,N_7054);
nand U7245 (N_7245,N_7064,N_7078);
nand U7246 (N_7246,N_7166,N_7170);
nand U7247 (N_7247,N_7121,N_7162);
nand U7248 (N_7248,N_7174,N_7124);
nor U7249 (N_7249,N_7140,N_7142);
nand U7250 (N_7250,N_7103,N_7191);
nand U7251 (N_7251,N_7126,N_7089);
or U7252 (N_7252,N_7199,N_7048);
or U7253 (N_7253,N_7143,N_7076);
or U7254 (N_7254,N_7185,N_7065);
xnor U7255 (N_7255,N_7041,N_7021);
nand U7256 (N_7256,N_7148,N_7105);
nor U7257 (N_7257,N_7195,N_7189);
xor U7258 (N_7258,N_7027,N_7159);
and U7259 (N_7259,N_7129,N_7194);
nor U7260 (N_7260,N_7116,N_7113);
nand U7261 (N_7261,N_7086,N_7052);
or U7262 (N_7262,N_7018,N_7172);
or U7263 (N_7263,N_7010,N_7008);
xor U7264 (N_7264,N_7163,N_7083);
nand U7265 (N_7265,N_7150,N_7117);
or U7266 (N_7266,N_7145,N_7106);
or U7267 (N_7267,N_7111,N_7062);
xor U7268 (N_7268,N_7029,N_7125);
and U7269 (N_7269,N_7136,N_7093);
xnor U7270 (N_7270,N_7037,N_7058);
or U7271 (N_7271,N_7171,N_7100);
nand U7272 (N_7272,N_7101,N_7032);
or U7273 (N_7273,N_7112,N_7009);
and U7274 (N_7274,N_7049,N_7030);
xnor U7275 (N_7275,N_7087,N_7025);
nand U7276 (N_7276,N_7045,N_7061);
and U7277 (N_7277,N_7133,N_7127);
nand U7278 (N_7278,N_7134,N_7031);
and U7279 (N_7279,N_7183,N_7181);
xnor U7280 (N_7280,N_7044,N_7147);
and U7281 (N_7281,N_7011,N_7164);
or U7282 (N_7282,N_7187,N_7096);
xnor U7283 (N_7283,N_7072,N_7176);
xnor U7284 (N_7284,N_7014,N_7180);
nand U7285 (N_7285,N_7091,N_7050);
nand U7286 (N_7286,N_7188,N_7168);
or U7287 (N_7287,N_7074,N_7075);
xnor U7288 (N_7288,N_7178,N_7004);
nand U7289 (N_7289,N_7123,N_7066);
or U7290 (N_7290,N_7177,N_7167);
nand U7291 (N_7291,N_7175,N_7015);
nor U7292 (N_7292,N_7024,N_7056);
or U7293 (N_7293,N_7073,N_7157);
and U7294 (N_7294,N_7151,N_7055);
nor U7295 (N_7295,N_7095,N_7193);
and U7296 (N_7296,N_7068,N_7007);
xnor U7297 (N_7297,N_7190,N_7082);
nor U7298 (N_7298,N_7156,N_7017);
xnor U7299 (N_7299,N_7158,N_7115);
nand U7300 (N_7300,N_7001,N_7042);
nand U7301 (N_7301,N_7029,N_7110);
nand U7302 (N_7302,N_7022,N_7116);
nor U7303 (N_7303,N_7179,N_7116);
nor U7304 (N_7304,N_7023,N_7027);
nor U7305 (N_7305,N_7046,N_7169);
nor U7306 (N_7306,N_7046,N_7062);
nand U7307 (N_7307,N_7061,N_7031);
nor U7308 (N_7308,N_7168,N_7067);
nand U7309 (N_7309,N_7084,N_7056);
nand U7310 (N_7310,N_7148,N_7120);
nand U7311 (N_7311,N_7157,N_7142);
and U7312 (N_7312,N_7105,N_7000);
nor U7313 (N_7313,N_7159,N_7103);
xor U7314 (N_7314,N_7169,N_7068);
xnor U7315 (N_7315,N_7172,N_7156);
nor U7316 (N_7316,N_7079,N_7037);
nand U7317 (N_7317,N_7010,N_7055);
nor U7318 (N_7318,N_7119,N_7026);
xnor U7319 (N_7319,N_7087,N_7091);
nor U7320 (N_7320,N_7131,N_7047);
nand U7321 (N_7321,N_7180,N_7063);
nand U7322 (N_7322,N_7003,N_7138);
or U7323 (N_7323,N_7024,N_7023);
and U7324 (N_7324,N_7056,N_7091);
and U7325 (N_7325,N_7016,N_7084);
xnor U7326 (N_7326,N_7000,N_7023);
nand U7327 (N_7327,N_7117,N_7023);
xnor U7328 (N_7328,N_7003,N_7173);
nor U7329 (N_7329,N_7168,N_7153);
xor U7330 (N_7330,N_7151,N_7173);
or U7331 (N_7331,N_7024,N_7048);
nand U7332 (N_7332,N_7181,N_7161);
or U7333 (N_7333,N_7034,N_7108);
xnor U7334 (N_7334,N_7186,N_7107);
and U7335 (N_7335,N_7056,N_7155);
xor U7336 (N_7336,N_7044,N_7057);
nand U7337 (N_7337,N_7110,N_7191);
nand U7338 (N_7338,N_7107,N_7133);
nand U7339 (N_7339,N_7192,N_7185);
nor U7340 (N_7340,N_7084,N_7003);
or U7341 (N_7341,N_7034,N_7102);
xor U7342 (N_7342,N_7169,N_7014);
xor U7343 (N_7343,N_7143,N_7032);
or U7344 (N_7344,N_7082,N_7071);
nand U7345 (N_7345,N_7033,N_7181);
xor U7346 (N_7346,N_7185,N_7039);
xor U7347 (N_7347,N_7023,N_7173);
or U7348 (N_7348,N_7111,N_7165);
xor U7349 (N_7349,N_7196,N_7085);
xor U7350 (N_7350,N_7107,N_7111);
nand U7351 (N_7351,N_7106,N_7057);
nand U7352 (N_7352,N_7147,N_7158);
nand U7353 (N_7353,N_7187,N_7059);
nor U7354 (N_7354,N_7117,N_7199);
nor U7355 (N_7355,N_7144,N_7065);
nand U7356 (N_7356,N_7151,N_7109);
nor U7357 (N_7357,N_7186,N_7144);
and U7358 (N_7358,N_7178,N_7093);
xnor U7359 (N_7359,N_7130,N_7107);
and U7360 (N_7360,N_7079,N_7031);
or U7361 (N_7361,N_7027,N_7006);
nor U7362 (N_7362,N_7156,N_7113);
or U7363 (N_7363,N_7199,N_7038);
xnor U7364 (N_7364,N_7124,N_7186);
nand U7365 (N_7365,N_7098,N_7026);
nand U7366 (N_7366,N_7170,N_7169);
xor U7367 (N_7367,N_7017,N_7096);
nand U7368 (N_7368,N_7178,N_7113);
or U7369 (N_7369,N_7076,N_7015);
nand U7370 (N_7370,N_7001,N_7013);
nor U7371 (N_7371,N_7129,N_7045);
xnor U7372 (N_7372,N_7131,N_7052);
nor U7373 (N_7373,N_7025,N_7002);
nor U7374 (N_7374,N_7019,N_7030);
xnor U7375 (N_7375,N_7029,N_7015);
and U7376 (N_7376,N_7001,N_7072);
and U7377 (N_7377,N_7040,N_7157);
xor U7378 (N_7378,N_7109,N_7153);
or U7379 (N_7379,N_7192,N_7070);
or U7380 (N_7380,N_7181,N_7165);
xnor U7381 (N_7381,N_7058,N_7053);
xnor U7382 (N_7382,N_7051,N_7174);
nor U7383 (N_7383,N_7089,N_7030);
or U7384 (N_7384,N_7079,N_7007);
or U7385 (N_7385,N_7146,N_7055);
nand U7386 (N_7386,N_7124,N_7112);
nor U7387 (N_7387,N_7191,N_7083);
nand U7388 (N_7388,N_7182,N_7006);
nand U7389 (N_7389,N_7133,N_7162);
nand U7390 (N_7390,N_7064,N_7188);
and U7391 (N_7391,N_7081,N_7160);
and U7392 (N_7392,N_7060,N_7008);
nand U7393 (N_7393,N_7059,N_7145);
xor U7394 (N_7394,N_7146,N_7139);
xnor U7395 (N_7395,N_7166,N_7188);
xnor U7396 (N_7396,N_7004,N_7191);
and U7397 (N_7397,N_7081,N_7165);
xor U7398 (N_7398,N_7033,N_7013);
and U7399 (N_7399,N_7144,N_7040);
and U7400 (N_7400,N_7309,N_7385);
and U7401 (N_7401,N_7370,N_7339);
xnor U7402 (N_7402,N_7275,N_7217);
nand U7403 (N_7403,N_7271,N_7298);
or U7404 (N_7404,N_7238,N_7336);
and U7405 (N_7405,N_7320,N_7310);
nor U7406 (N_7406,N_7231,N_7380);
xor U7407 (N_7407,N_7297,N_7204);
or U7408 (N_7408,N_7332,N_7268);
or U7409 (N_7409,N_7304,N_7345);
or U7410 (N_7410,N_7236,N_7393);
and U7411 (N_7411,N_7224,N_7360);
nor U7412 (N_7412,N_7388,N_7299);
and U7413 (N_7413,N_7372,N_7256);
nand U7414 (N_7414,N_7364,N_7270);
nand U7415 (N_7415,N_7250,N_7350);
and U7416 (N_7416,N_7206,N_7335);
xor U7417 (N_7417,N_7211,N_7261);
nand U7418 (N_7418,N_7343,N_7296);
nor U7419 (N_7419,N_7289,N_7252);
xor U7420 (N_7420,N_7286,N_7301);
and U7421 (N_7421,N_7379,N_7284);
xnor U7422 (N_7422,N_7327,N_7306);
nor U7423 (N_7423,N_7207,N_7361);
or U7424 (N_7424,N_7242,N_7221);
nand U7425 (N_7425,N_7226,N_7315);
and U7426 (N_7426,N_7333,N_7237);
nand U7427 (N_7427,N_7347,N_7325);
and U7428 (N_7428,N_7287,N_7396);
nand U7429 (N_7429,N_7203,N_7305);
or U7430 (N_7430,N_7210,N_7258);
or U7431 (N_7431,N_7294,N_7334);
or U7432 (N_7432,N_7342,N_7265);
xor U7433 (N_7433,N_7355,N_7316);
nand U7434 (N_7434,N_7220,N_7277);
or U7435 (N_7435,N_7337,N_7240);
nand U7436 (N_7436,N_7225,N_7201);
xor U7437 (N_7437,N_7213,N_7251);
or U7438 (N_7438,N_7308,N_7389);
or U7439 (N_7439,N_7291,N_7399);
and U7440 (N_7440,N_7331,N_7373);
nand U7441 (N_7441,N_7283,N_7245);
and U7442 (N_7442,N_7216,N_7254);
nor U7443 (N_7443,N_7311,N_7382);
and U7444 (N_7444,N_7293,N_7212);
nor U7445 (N_7445,N_7313,N_7227);
or U7446 (N_7446,N_7290,N_7324);
xnor U7447 (N_7447,N_7255,N_7234);
nand U7448 (N_7448,N_7295,N_7249);
or U7449 (N_7449,N_7367,N_7264);
nand U7450 (N_7450,N_7369,N_7281);
and U7451 (N_7451,N_7377,N_7274);
nand U7452 (N_7452,N_7392,N_7241);
nand U7453 (N_7453,N_7257,N_7384);
nand U7454 (N_7454,N_7303,N_7247);
or U7455 (N_7455,N_7329,N_7346);
xor U7456 (N_7456,N_7358,N_7368);
nor U7457 (N_7457,N_7340,N_7398);
or U7458 (N_7458,N_7317,N_7349);
nand U7459 (N_7459,N_7263,N_7228);
xnor U7460 (N_7460,N_7222,N_7330);
xor U7461 (N_7461,N_7260,N_7307);
or U7462 (N_7462,N_7266,N_7302);
nand U7463 (N_7463,N_7390,N_7285);
or U7464 (N_7464,N_7282,N_7383);
nand U7465 (N_7465,N_7366,N_7279);
or U7466 (N_7466,N_7397,N_7363);
and U7467 (N_7467,N_7208,N_7344);
nor U7468 (N_7468,N_7362,N_7230);
or U7469 (N_7469,N_7280,N_7312);
and U7470 (N_7470,N_7200,N_7328);
or U7471 (N_7471,N_7338,N_7300);
or U7472 (N_7472,N_7348,N_7214);
and U7473 (N_7473,N_7394,N_7319);
nor U7474 (N_7474,N_7215,N_7357);
xnor U7475 (N_7475,N_7248,N_7314);
xnor U7476 (N_7476,N_7239,N_7223);
and U7477 (N_7477,N_7219,N_7386);
or U7478 (N_7478,N_7352,N_7387);
nor U7479 (N_7479,N_7273,N_7371);
nor U7480 (N_7480,N_7272,N_7218);
or U7481 (N_7481,N_7267,N_7326);
xor U7482 (N_7482,N_7395,N_7365);
or U7483 (N_7483,N_7292,N_7354);
nand U7484 (N_7484,N_7233,N_7321);
xnor U7485 (N_7485,N_7205,N_7278);
and U7486 (N_7486,N_7341,N_7288);
xor U7487 (N_7487,N_7262,N_7276);
xor U7488 (N_7488,N_7351,N_7318);
xor U7489 (N_7489,N_7253,N_7381);
and U7490 (N_7490,N_7235,N_7259);
xnor U7491 (N_7491,N_7232,N_7353);
nand U7492 (N_7492,N_7246,N_7376);
nand U7493 (N_7493,N_7229,N_7244);
nor U7494 (N_7494,N_7323,N_7391);
nor U7495 (N_7495,N_7378,N_7269);
or U7496 (N_7496,N_7375,N_7322);
nand U7497 (N_7497,N_7202,N_7374);
or U7498 (N_7498,N_7359,N_7356);
nor U7499 (N_7499,N_7209,N_7243);
xnor U7500 (N_7500,N_7388,N_7294);
xnor U7501 (N_7501,N_7273,N_7368);
and U7502 (N_7502,N_7230,N_7223);
nand U7503 (N_7503,N_7263,N_7384);
xor U7504 (N_7504,N_7273,N_7287);
or U7505 (N_7505,N_7367,N_7223);
nand U7506 (N_7506,N_7316,N_7281);
nand U7507 (N_7507,N_7246,N_7395);
or U7508 (N_7508,N_7351,N_7381);
or U7509 (N_7509,N_7315,N_7228);
or U7510 (N_7510,N_7281,N_7256);
nor U7511 (N_7511,N_7255,N_7250);
nand U7512 (N_7512,N_7316,N_7202);
or U7513 (N_7513,N_7206,N_7369);
and U7514 (N_7514,N_7396,N_7295);
nor U7515 (N_7515,N_7207,N_7230);
and U7516 (N_7516,N_7236,N_7307);
and U7517 (N_7517,N_7354,N_7205);
nand U7518 (N_7518,N_7251,N_7211);
or U7519 (N_7519,N_7393,N_7304);
or U7520 (N_7520,N_7355,N_7312);
or U7521 (N_7521,N_7204,N_7292);
and U7522 (N_7522,N_7347,N_7375);
nand U7523 (N_7523,N_7282,N_7267);
or U7524 (N_7524,N_7369,N_7321);
xor U7525 (N_7525,N_7273,N_7209);
and U7526 (N_7526,N_7397,N_7270);
nor U7527 (N_7527,N_7353,N_7270);
or U7528 (N_7528,N_7264,N_7353);
nor U7529 (N_7529,N_7384,N_7392);
nand U7530 (N_7530,N_7301,N_7353);
and U7531 (N_7531,N_7258,N_7220);
nor U7532 (N_7532,N_7390,N_7311);
and U7533 (N_7533,N_7250,N_7357);
nand U7534 (N_7534,N_7317,N_7208);
or U7535 (N_7535,N_7331,N_7391);
nor U7536 (N_7536,N_7258,N_7203);
xor U7537 (N_7537,N_7221,N_7206);
and U7538 (N_7538,N_7238,N_7301);
or U7539 (N_7539,N_7256,N_7244);
xor U7540 (N_7540,N_7346,N_7272);
nor U7541 (N_7541,N_7230,N_7248);
xor U7542 (N_7542,N_7330,N_7235);
xnor U7543 (N_7543,N_7240,N_7257);
nor U7544 (N_7544,N_7252,N_7224);
xnor U7545 (N_7545,N_7318,N_7288);
xnor U7546 (N_7546,N_7219,N_7334);
or U7547 (N_7547,N_7385,N_7229);
or U7548 (N_7548,N_7201,N_7229);
and U7549 (N_7549,N_7270,N_7392);
xor U7550 (N_7550,N_7261,N_7223);
nand U7551 (N_7551,N_7337,N_7326);
and U7552 (N_7552,N_7250,N_7366);
xor U7553 (N_7553,N_7245,N_7216);
and U7554 (N_7554,N_7340,N_7295);
nor U7555 (N_7555,N_7202,N_7233);
xnor U7556 (N_7556,N_7249,N_7273);
nor U7557 (N_7557,N_7314,N_7235);
nor U7558 (N_7558,N_7214,N_7280);
nor U7559 (N_7559,N_7311,N_7300);
nand U7560 (N_7560,N_7209,N_7336);
nor U7561 (N_7561,N_7205,N_7395);
nor U7562 (N_7562,N_7389,N_7372);
or U7563 (N_7563,N_7312,N_7342);
xnor U7564 (N_7564,N_7302,N_7260);
and U7565 (N_7565,N_7221,N_7251);
and U7566 (N_7566,N_7284,N_7380);
nor U7567 (N_7567,N_7311,N_7334);
and U7568 (N_7568,N_7290,N_7328);
and U7569 (N_7569,N_7387,N_7231);
xnor U7570 (N_7570,N_7259,N_7253);
xnor U7571 (N_7571,N_7261,N_7333);
or U7572 (N_7572,N_7238,N_7284);
nand U7573 (N_7573,N_7360,N_7347);
nand U7574 (N_7574,N_7356,N_7367);
nor U7575 (N_7575,N_7262,N_7365);
nand U7576 (N_7576,N_7256,N_7362);
xor U7577 (N_7577,N_7251,N_7202);
nor U7578 (N_7578,N_7287,N_7321);
or U7579 (N_7579,N_7233,N_7211);
or U7580 (N_7580,N_7352,N_7224);
and U7581 (N_7581,N_7255,N_7240);
and U7582 (N_7582,N_7356,N_7282);
nand U7583 (N_7583,N_7296,N_7229);
and U7584 (N_7584,N_7299,N_7352);
nand U7585 (N_7585,N_7223,N_7290);
and U7586 (N_7586,N_7352,N_7205);
xor U7587 (N_7587,N_7269,N_7245);
or U7588 (N_7588,N_7370,N_7201);
xor U7589 (N_7589,N_7285,N_7262);
nor U7590 (N_7590,N_7257,N_7268);
nand U7591 (N_7591,N_7217,N_7297);
nor U7592 (N_7592,N_7219,N_7355);
and U7593 (N_7593,N_7201,N_7377);
nand U7594 (N_7594,N_7201,N_7216);
nor U7595 (N_7595,N_7233,N_7291);
nor U7596 (N_7596,N_7352,N_7238);
or U7597 (N_7597,N_7264,N_7239);
and U7598 (N_7598,N_7298,N_7393);
and U7599 (N_7599,N_7303,N_7330);
xnor U7600 (N_7600,N_7542,N_7458);
nor U7601 (N_7601,N_7557,N_7413);
and U7602 (N_7602,N_7481,N_7595);
and U7603 (N_7603,N_7409,N_7568);
nand U7604 (N_7604,N_7570,N_7567);
or U7605 (N_7605,N_7441,N_7402);
nor U7606 (N_7606,N_7579,N_7505);
nand U7607 (N_7607,N_7523,N_7565);
xnor U7608 (N_7608,N_7545,N_7574);
and U7609 (N_7609,N_7411,N_7566);
xnor U7610 (N_7610,N_7527,N_7528);
and U7611 (N_7611,N_7475,N_7462);
nand U7612 (N_7612,N_7407,N_7585);
and U7613 (N_7613,N_7434,N_7455);
and U7614 (N_7614,N_7487,N_7406);
xnor U7615 (N_7615,N_7476,N_7597);
or U7616 (N_7616,N_7526,N_7492);
nand U7617 (N_7617,N_7418,N_7572);
and U7618 (N_7618,N_7591,N_7543);
and U7619 (N_7619,N_7564,N_7422);
or U7620 (N_7620,N_7581,N_7587);
xnor U7621 (N_7621,N_7414,N_7547);
nor U7622 (N_7622,N_7474,N_7541);
or U7623 (N_7623,N_7494,N_7513);
nand U7624 (N_7624,N_7436,N_7575);
nor U7625 (N_7625,N_7514,N_7596);
nand U7626 (N_7626,N_7578,N_7447);
xor U7627 (N_7627,N_7599,N_7583);
xor U7628 (N_7628,N_7460,N_7509);
xor U7629 (N_7629,N_7497,N_7424);
xnor U7630 (N_7630,N_7561,N_7582);
nor U7631 (N_7631,N_7558,N_7553);
xnor U7632 (N_7632,N_7540,N_7501);
and U7633 (N_7633,N_7469,N_7552);
nand U7634 (N_7634,N_7408,N_7534);
and U7635 (N_7635,N_7478,N_7423);
or U7636 (N_7636,N_7431,N_7464);
or U7637 (N_7637,N_7510,N_7525);
nor U7638 (N_7638,N_7521,N_7593);
xnor U7639 (N_7639,N_7446,N_7461);
or U7640 (N_7640,N_7554,N_7559);
and U7641 (N_7641,N_7508,N_7483);
xor U7642 (N_7642,N_7598,N_7479);
or U7643 (N_7643,N_7437,N_7499);
nor U7644 (N_7644,N_7556,N_7442);
nor U7645 (N_7645,N_7440,N_7531);
nor U7646 (N_7646,N_7507,N_7573);
nor U7647 (N_7647,N_7537,N_7555);
or U7648 (N_7648,N_7577,N_7400);
nand U7649 (N_7649,N_7401,N_7512);
xor U7650 (N_7650,N_7450,N_7421);
nor U7651 (N_7651,N_7480,N_7432);
xnor U7652 (N_7652,N_7562,N_7524);
and U7653 (N_7653,N_7502,N_7500);
or U7654 (N_7654,N_7457,N_7420);
nor U7655 (N_7655,N_7430,N_7425);
nor U7656 (N_7656,N_7463,N_7580);
and U7657 (N_7657,N_7491,N_7451);
nand U7658 (N_7658,N_7517,N_7466);
and U7659 (N_7659,N_7445,N_7589);
and U7660 (N_7660,N_7538,N_7576);
nor U7661 (N_7661,N_7456,N_7443);
nor U7662 (N_7662,N_7549,N_7433);
and U7663 (N_7663,N_7520,N_7560);
nand U7664 (N_7664,N_7495,N_7515);
nand U7665 (N_7665,N_7529,N_7449);
and U7666 (N_7666,N_7532,N_7438);
xor U7667 (N_7667,N_7415,N_7468);
nor U7668 (N_7668,N_7503,N_7426);
xor U7669 (N_7669,N_7496,N_7533);
or U7670 (N_7670,N_7482,N_7403);
xnor U7671 (N_7671,N_7427,N_7429);
and U7672 (N_7672,N_7488,N_7439);
nand U7673 (N_7673,N_7519,N_7546);
and U7674 (N_7674,N_7498,N_7569);
nand U7675 (N_7675,N_7536,N_7493);
and U7676 (N_7676,N_7448,N_7477);
nor U7677 (N_7677,N_7594,N_7467);
nand U7678 (N_7678,N_7419,N_7544);
xnor U7679 (N_7679,N_7530,N_7539);
or U7680 (N_7680,N_7550,N_7592);
nand U7681 (N_7681,N_7548,N_7485);
or U7682 (N_7682,N_7405,N_7586);
xnor U7683 (N_7683,N_7486,N_7459);
nand U7684 (N_7684,N_7588,N_7551);
nor U7685 (N_7685,N_7563,N_7435);
and U7686 (N_7686,N_7571,N_7504);
nor U7687 (N_7687,N_7584,N_7473);
and U7688 (N_7688,N_7511,N_7484);
and U7689 (N_7689,N_7444,N_7518);
and U7690 (N_7690,N_7522,N_7404);
nor U7691 (N_7691,N_7535,N_7506);
or U7692 (N_7692,N_7489,N_7454);
xor U7693 (N_7693,N_7516,N_7465);
nor U7694 (N_7694,N_7590,N_7428);
nor U7695 (N_7695,N_7417,N_7452);
nand U7696 (N_7696,N_7412,N_7416);
nor U7697 (N_7697,N_7471,N_7470);
and U7698 (N_7698,N_7490,N_7410);
nand U7699 (N_7699,N_7472,N_7453);
nor U7700 (N_7700,N_7437,N_7563);
xor U7701 (N_7701,N_7453,N_7482);
xnor U7702 (N_7702,N_7588,N_7526);
and U7703 (N_7703,N_7586,N_7464);
nor U7704 (N_7704,N_7410,N_7563);
xor U7705 (N_7705,N_7471,N_7537);
nor U7706 (N_7706,N_7519,N_7588);
xor U7707 (N_7707,N_7439,N_7474);
xnor U7708 (N_7708,N_7547,N_7440);
nor U7709 (N_7709,N_7482,N_7563);
xnor U7710 (N_7710,N_7525,N_7413);
xnor U7711 (N_7711,N_7426,N_7436);
and U7712 (N_7712,N_7428,N_7448);
xor U7713 (N_7713,N_7500,N_7546);
and U7714 (N_7714,N_7537,N_7581);
and U7715 (N_7715,N_7402,N_7550);
nand U7716 (N_7716,N_7586,N_7474);
nor U7717 (N_7717,N_7599,N_7451);
nor U7718 (N_7718,N_7427,N_7504);
or U7719 (N_7719,N_7564,N_7484);
nand U7720 (N_7720,N_7586,N_7579);
xor U7721 (N_7721,N_7471,N_7477);
xnor U7722 (N_7722,N_7580,N_7457);
nor U7723 (N_7723,N_7473,N_7492);
nand U7724 (N_7724,N_7438,N_7459);
nand U7725 (N_7725,N_7467,N_7472);
and U7726 (N_7726,N_7557,N_7425);
xor U7727 (N_7727,N_7530,N_7543);
nand U7728 (N_7728,N_7448,N_7533);
xor U7729 (N_7729,N_7522,N_7541);
or U7730 (N_7730,N_7512,N_7500);
nor U7731 (N_7731,N_7582,N_7439);
nor U7732 (N_7732,N_7583,N_7419);
nor U7733 (N_7733,N_7525,N_7446);
nand U7734 (N_7734,N_7412,N_7591);
nand U7735 (N_7735,N_7505,N_7551);
or U7736 (N_7736,N_7486,N_7596);
nand U7737 (N_7737,N_7458,N_7581);
xnor U7738 (N_7738,N_7414,N_7411);
nor U7739 (N_7739,N_7460,N_7505);
nand U7740 (N_7740,N_7504,N_7547);
nor U7741 (N_7741,N_7553,N_7411);
nor U7742 (N_7742,N_7586,N_7527);
nor U7743 (N_7743,N_7529,N_7523);
nor U7744 (N_7744,N_7586,N_7573);
nor U7745 (N_7745,N_7516,N_7479);
nor U7746 (N_7746,N_7599,N_7428);
or U7747 (N_7747,N_7471,N_7455);
and U7748 (N_7748,N_7481,N_7537);
nor U7749 (N_7749,N_7584,N_7457);
or U7750 (N_7750,N_7494,N_7561);
and U7751 (N_7751,N_7503,N_7482);
and U7752 (N_7752,N_7508,N_7574);
or U7753 (N_7753,N_7596,N_7551);
xnor U7754 (N_7754,N_7483,N_7411);
nor U7755 (N_7755,N_7588,N_7545);
nand U7756 (N_7756,N_7530,N_7569);
nand U7757 (N_7757,N_7594,N_7584);
nor U7758 (N_7758,N_7559,N_7496);
and U7759 (N_7759,N_7517,N_7552);
xnor U7760 (N_7760,N_7458,N_7493);
and U7761 (N_7761,N_7599,N_7598);
nor U7762 (N_7762,N_7485,N_7546);
or U7763 (N_7763,N_7542,N_7502);
nand U7764 (N_7764,N_7445,N_7401);
xnor U7765 (N_7765,N_7401,N_7568);
nand U7766 (N_7766,N_7477,N_7427);
and U7767 (N_7767,N_7417,N_7543);
and U7768 (N_7768,N_7597,N_7501);
nand U7769 (N_7769,N_7424,N_7556);
nor U7770 (N_7770,N_7535,N_7436);
nand U7771 (N_7771,N_7492,N_7545);
or U7772 (N_7772,N_7423,N_7435);
or U7773 (N_7773,N_7411,N_7492);
nand U7774 (N_7774,N_7564,N_7505);
nand U7775 (N_7775,N_7514,N_7483);
nand U7776 (N_7776,N_7550,N_7413);
nor U7777 (N_7777,N_7410,N_7576);
and U7778 (N_7778,N_7510,N_7439);
nor U7779 (N_7779,N_7584,N_7467);
or U7780 (N_7780,N_7583,N_7575);
and U7781 (N_7781,N_7421,N_7503);
nor U7782 (N_7782,N_7513,N_7530);
or U7783 (N_7783,N_7471,N_7524);
and U7784 (N_7784,N_7522,N_7422);
nand U7785 (N_7785,N_7486,N_7594);
xor U7786 (N_7786,N_7588,N_7535);
nand U7787 (N_7787,N_7500,N_7452);
or U7788 (N_7788,N_7485,N_7481);
nor U7789 (N_7789,N_7535,N_7492);
nor U7790 (N_7790,N_7552,N_7493);
and U7791 (N_7791,N_7430,N_7519);
or U7792 (N_7792,N_7456,N_7453);
xor U7793 (N_7793,N_7453,N_7433);
nand U7794 (N_7794,N_7528,N_7513);
or U7795 (N_7795,N_7561,N_7535);
and U7796 (N_7796,N_7413,N_7586);
nand U7797 (N_7797,N_7498,N_7517);
xor U7798 (N_7798,N_7460,N_7414);
nand U7799 (N_7799,N_7489,N_7506);
or U7800 (N_7800,N_7709,N_7697);
xor U7801 (N_7801,N_7747,N_7761);
xnor U7802 (N_7802,N_7618,N_7691);
nand U7803 (N_7803,N_7622,N_7721);
nand U7804 (N_7804,N_7671,N_7674);
or U7805 (N_7805,N_7648,N_7765);
and U7806 (N_7806,N_7796,N_7665);
and U7807 (N_7807,N_7694,N_7640);
nor U7808 (N_7808,N_7766,N_7693);
xor U7809 (N_7809,N_7630,N_7741);
xor U7810 (N_7810,N_7685,N_7667);
xor U7811 (N_7811,N_7773,N_7654);
xor U7812 (N_7812,N_7732,N_7713);
nand U7813 (N_7813,N_7635,N_7774);
xnor U7814 (N_7814,N_7708,N_7661);
and U7815 (N_7815,N_7743,N_7725);
xnor U7816 (N_7816,N_7601,N_7656);
nand U7817 (N_7817,N_7609,N_7620);
and U7818 (N_7818,N_7679,N_7727);
xnor U7819 (N_7819,N_7631,N_7789);
nand U7820 (N_7820,N_7730,N_7675);
and U7821 (N_7821,N_7681,N_7615);
and U7822 (N_7822,N_7722,N_7612);
nor U7823 (N_7823,N_7737,N_7670);
xor U7824 (N_7824,N_7611,N_7791);
nor U7825 (N_7825,N_7792,N_7759);
or U7826 (N_7826,N_7650,N_7775);
and U7827 (N_7827,N_7680,N_7720);
nor U7828 (N_7828,N_7718,N_7700);
nand U7829 (N_7829,N_7764,N_7702);
and U7830 (N_7830,N_7715,N_7628);
nor U7831 (N_7831,N_7632,N_7798);
xnor U7832 (N_7832,N_7657,N_7610);
or U7833 (N_7833,N_7664,N_7688);
nand U7834 (N_7834,N_7644,N_7662);
nand U7835 (N_7835,N_7782,N_7728);
or U7836 (N_7836,N_7666,N_7704);
and U7837 (N_7837,N_7642,N_7734);
or U7838 (N_7838,N_7659,N_7617);
nand U7839 (N_7839,N_7690,N_7748);
or U7840 (N_7840,N_7756,N_7677);
xor U7841 (N_7841,N_7724,N_7613);
nor U7842 (N_7842,N_7772,N_7658);
xor U7843 (N_7843,N_7699,N_7776);
xor U7844 (N_7844,N_7760,N_7768);
xnor U7845 (N_7845,N_7636,N_7784);
nor U7846 (N_7846,N_7624,N_7738);
and U7847 (N_7847,N_7653,N_7770);
nor U7848 (N_7848,N_7757,N_7625);
and U7849 (N_7849,N_7785,N_7703);
xnor U7850 (N_7850,N_7733,N_7669);
and U7851 (N_7851,N_7649,N_7746);
nand U7852 (N_7852,N_7646,N_7607);
and U7853 (N_7853,N_7602,N_7778);
nand U7854 (N_7854,N_7637,N_7729);
and U7855 (N_7855,N_7723,N_7735);
nand U7856 (N_7856,N_7626,N_7771);
or U7857 (N_7857,N_7707,N_7614);
xnor U7858 (N_7858,N_7672,N_7604);
or U7859 (N_7859,N_7797,N_7623);
xnor U7860 (N_7860,N_7783,N_7711);
and U7861 (N_7861,N_7689,N_7692);
xor U7862 (N_7862,N_7744,N_7608);
nand U7863 (N_7863,N_7714,N_7655);
and U7864 (N_7864,N_7762,N_7763);
xor U7865 (N_7865,N_7682,N_7786);
nor U7866 (N_7866,N_7780,N_7600);
nor U7867 (N_7867,N_7634,N_7710);
nor U7868 (N_7868,N_7660,N_7750);
xnor U7869 (N_7869,N_7769,N_7645);
xor U7870 (N_7870,N_7668,N_7739);
nor U7871 (N_7871,N_7736,N_7716);
and U7872 (N_7872,N_7651,N_7705);
nand U7873 (N_7873,N_7616,N_7740);
or U7874 (N_7874,N_7673,N_7621);
and U7875 (N_7875,N_7695,N_7790);
nand U7876 (N_7876,N_7638,N_7641);
nand U7877 (N_7877,N_7754,N_7749);
and U7878 (N_7878,N_7603,N_7794);
xor U7879 (N_7879,N_7643,N_7619);
or U7880 (N_7880,N_7652,N_7627);
nor U7881 (N_7881,N_7686,N_7726);
and U7882 (N_7882,N_7799,N_7781);
and U7883 (N_7883,N_7647,N_7712);
and U7884 (N_7884,N_7663,N_7717);
nor U7885 (N_7885,N_7752,N_7758);
nor U7886 (N_7886,N_7731,N_7753);
nor U7887 (N_7887,N_7687,N_7701);
xor U7888 (N_7888,N_7639,N_7788);
and U7889 (N_7889,N_7755,N_7795);
nor U7890 (N_7890,N_7676,N_7719);
nor U7891 (N_7891,N_7605,N_7793);
or U7892 (N_7892,N_7678,N_7683);
or U7893 (N_7893,N_7606,N_7684);
xor U7894 (N_7894,N_7742,N_7767);
nand U7895 (N_7895,N_7787,N_7751);
and U7896 (N_7896,N_7696,N_7633);
or U7897 (N_7897,N_7745,N_7706);
or U7898 (N_7898,N_7629,N_7698);
nand U7899 (N_7899,N_7779,N_7777);
or U7900 (N_7900,N_7744,N_7731);
or U7901 (N_7901,N_7676,N_7797);
xor U7902 (N_7902,N_7792,N_7754);
or U7903 (N_7903,N_7785,N_7758);
nor U7904 (N_7904,N_7748,N_7778);
nand U7905 (N_7905,N_7659,N_7649);
nor U7906 (N_7906,N_7611,N_7671);
or U7907 (N_7907,N_7765,N_7633);
nand U7908 (N_7908,N_7641,N_7750);
xor U7909 (N_7909,N_7737,N_7740);
nor U7910 (N_7910,N_7634,N_7730);
nor U7911 (N_7911,N_7657,N_7618);
and U7912 (N_7912,N_7631,N_7756);
and U7913 (N_7913,N_7770,N_7662);
nor U7914 (N_7914,N_7767,N_7638);
or U7915 (N_7915,N_7622,N_7618);
nand U7916 (N_7916,N_7649,N_7720);
and U7917 (N_7917,N_7785,N_7693);
nor U7918 (N_7918,N_7620,N_7611);
nor U7919 (N_7919,N_7658,N_7606);
nor U7920 (N_7920,N_7650,N_7792);
nor U7921 (N_7921,N_7616,N_7638);
nor U7922 (N_7922,N_7702,N_7720);
nor U7923 (N_7923,N_7655,N_7604);
xor U7924 (N_7924,N_7759,N_7763);
nor U7925 (N_7925,N_7732,N_7716);
xor U7926 (N_7926,N_7648,N_7664);
nor U7927 (N_7927,N_7737,N_7761);
or U7928 (N_7928,N_7795,N_7621);
nor U7929 (N_7929,N_7716,N_7705);
or U7930 (N_7930,N_7697,N_7797);
and U7931 (N_7931,N_7619,N_7710);
and U7932 (N_7932,N_7757,N_7716);
nor U7933 (N_7933,N_7649,N_7670);
and U7934 (N_7934,N_7615,N_7708);
xnor U7935 (N_7935,N_7747,N_7690);
xnor U7936 (N_7936,N_7732,N_7655);
and U7937 (N_7937,N_7711,N_7625);
nand U7938 (N_7938,N_7682,N_7668);
nand U7939 (N_7939,N_7737,N_7650);
and U7940 (N_7940,N_7767,N_7772);
nor U7941 (N_7941,N_7774,N_7719);
and U7942 (N_7942,N_7722,N_7765);
and U7943 (N_7943,N_7619,N_7753);
and U7944 (N_7944,N_7641,N_7757);
or U7945 (N_7945,N_7708,N_7702);
xnor U7946 (N_7946,N_7798,N_7732);
or U7947 (N_7947,N_7719,N_7752);
xnor U7948 (N_7948,N_7644,N_7764);
xnor U7949 (N_7949,N_7703,N_7685);
and U7950 (N_7950,N_7623,N_7741);
nor U7951 (N_7951,N_7612,N_7614);
xor U7952 (N_7952,N_7723,N_7772);
nand U7953 (N_7953,N_7620,N_7616);
xnor U7954 (N_7954,N_7780,N_7689);
xor U7955 (N_7955,N_7719,N_7748);
and U7956 (N_7956,N_7687,N_7706);
or U7957 (N_7957,N_7707,N_7718);
and U7958 (N_7958,N_7727,N_7791);
or U7959 (N_7959,N_7750,N_7733);
and U7960 (N_7960,N_7618,N_7679);
or U7961 (N_7961,N_7738,N_7718);
or U7962 (N_7962,N_7791,N_7637);
xor U7963 (N_7963,N_7675,N_7768);
and U7964 (N_7964,N_7732,N_7712);
or U7965 (N_7965,N_7626,N_7733);
and U7966 (N_7966,N_7750,N_7695);
xor U7967 (N_7967,N_7787,N_7612);
and U7968 (N_7968,N_7686,N_7752);
nor U7969 (N_7969,N_7611,N_7792);
xor U7970 (N_7970,N_7774,N_7650);
or U7971 (N_7971,N_7729,N_7751);
xor U7972 (N_7972,N_7742,N_7772);
or U7973 (N_7973,N_7616,N_7773);
xor U7974 (N_7974,N_7697,N_7700);
nand U7975 (N_7975,N_7608,N_7671);
xnor U7976 (N_7976,N_7646,N_7658);
xnor U7977 (N_7977,N_7794,N_7713);
and U7978 (N_7978,N_7676,N_7711);
xnor U7979 (N_7979,N_7682,N_7602);
and U7980 (N_7980,N_7618,N_7720);
or U7981 (N_7981,N_7754,N_7637);
nor U7982 (N_7982,N_7765,N_7759);
or U7983 (N_7983,N_7638,N_7668);
and U7984 (N_7984,N_7608,N_7767);
xor U7985 (N_7985,N_7748,N_7679);
xor U7986 (N_7986,N_7622,N_7662);
or U7987 (N_7987,N_7787,N_7670);
or U7988 (N_7988,N_7611,N_7699);
nand U7989 (N_7989,N_7667,N_7646);
or U7990 (N_7990,N_7624,N_7734);
nand U7991 (N_7991,N_7678,N_7787);
and U7992 (N_7992,N_7704,N_7791);
and U7993 (N_7993,N_7719,N_7772);
xnor U7994 (N_7994,N_7695,N_7618);
and U7995 (N_7995,N_7737,N_7792);
nor U7996 (N_7996,N_7787,N_7793);
nand U7997 (N_7997,N_7748,N_7707);
nand U7998 (N_7998,N_7652,N_7709);
and U7999 (N_7999,N_7718,N_7758);
or U8000 (N_8000,N_7815,N_7986);
nand U8001 (N_8001,N_7908,N_7967);
nand U8002 (N_8002,N_7835,N_7842);
nor U8003 (N_8003,N_7873,N_7861);
nor U8004 (N_8004,N_7858,N_7905);
nor U8005 (N_8005,N_7977,N_7935);
xnor U8006 (N_8006,N_7929,N_7919);
nand U8007 (N_8007,N_7994,N_7958);
and U8008 (N_8008,N_7846,N_7907);
nand U8009 (N_8009,N_7916,N_7979);
xnor U8010 (N_8010,N_7866,N_7889);
nor U8011 (N_8011,N_7820,N_7933);
nor U8012 (N_8012,N_7852,N_7906);
nor U8013 (N_8013,N_7829,N_7940);
xor U8014 (N_8014,N_7895,N_7938);
and U8015 (N_8015,N_7909,N_7999);
and U8016 (N_8016,N_7837,N_7839);
nor U8017 (N_8017,N_7981,N_7956);
xnor U8018 (N_8018,N_7863,N_7900);
and U8019 (N_8019,N_7893,N_7995);
xnor U8020 (N_8020,N_7985,N_7896);
xnor U8021 (N_8021,N_7973,N_7843);
nand U8022 (N_8022,N_7887,N_7879);
and U8023 (N_8023,N_7834,N_7961);
nand U8024 (N_8024,N_7899,N_7806);
and U8025 (N_8025,N_7888,N_7990);
nand U8026 (N_8026,N_7816,N_7825);
nand U8027 (N_8027,N_7821,N_7832);
or U8028 (N_8028,N_7849,N_7833);
or U8029 (N_8029,N_7865,N_7809);
nor U8030 (N_8030,N_7951,N_7871);
nand U8031 (N_8031,N_7957,N_7892);
or U8032 (N_8032,N_7841,N_7830);
and U8033 (N_8033,N_7847,N_7971);
and U8034 (N_8034,N_7913,N_7862);
and U8035 (N_8035,N_7910,N_7844);
and U8036 (N_8036,N_7886,N_7959);
or U8037 (N_8037,N_7932,N_7881);
and U8038 (N_8038,N_7931,N_7854);
or U8039 (N_8039,N_7855,N_7891);
or U8040 (N_8040,N_7805,N_7827);
xor U8041 (N_8041,N_7810,N_7975);
xnor U8042 (N_8042,N_7911,N_7992);
nor U8043 (N_8043,N_7876,N_7925);
or U8044 (N_8044,N_7914,N_7822);
or U8045 (N_8045,N_7883,N_7983);
or U8046 (N_8046,N_7955,N_7851);
xor U8047 (N_8047,N_7878,N_7978);
xor U8048 (N_8048,N_7921,N_7901);
and U8049 (N_8049,N_7944,N_7848);
or U8050 (N_8050,N_7870,N_7920);
xnor U8051 (N_8051,N_7860,N_7894);
and U8052 (N_8052,N_7924,N_7976);
nor U8053 (N_8053,N_7819,N_7853);
xnor U8054 (N_8054,N_7984,N_7996);
xnor U8055 (N_8055,N_7954,N_7812);
nor U8056 (N_8056,N_7803,N_7941);
nand U8057 (N_8057,N_7814,N_7939);
and U8058 (N_8058,N_7918,N_7942);
nand U8059 (N_8059,N_7828,N_7857);
xor U8060 (N_8060,N_7838,N_7950);
xor U8061 (N_8061,N_7903,N_7998);
or U8062 (N_8062,N_7943,N_7993);
or U8063 (N_8063,N_7937,N_7923);
or U8064 (N_8064,N_7930,N_7922);
or U8065 (N_8065,N_7946,N_7964);
and U8066 (N_8066,N_7856,N_7811);
and U8067 (N_8067,N_7884,N_7968);
xnor U8068 (N_8068,N_7991,N_7970);
nor U8069 (N_8069,N_7869,N_7836);
xor U8070 (N_8070,N_7966,N_7915);
or U8071 (N_8071,N_7867,N_7997);
or U8072 (N_8072,N_7801,N_7813);
nor U8073 (N_8073,N_7969,N_7800);
and U8074 (N_8074,N_7974,N_7912);
and U8075 (N_8075,N_7927,N_7904);
and U8076 (N_8076,N_7874,N_7972);
xnor U8077 (N_8077,N_7817,N_7936);
nor U8078 (N_8078,N_7963,N_7897);
nand U8079 (N_8079,N_7928,N_7880);
xor U8080 (N_8080,N_7890,N_7875);
xnor U8081 (N_8081,N_7831,N_7804);
or U8082 (N_8082,N_7988,N_7948);
nor U8083 (N_8083,N_7808,N_7949);
and U8084 (N_8084,N_7945,N_7980);
or U8085 (N_8085,N_7960,N_7850);
nand U8086 (N_8086,N_7864,N_7802);
and U8087 (N_8087,N_7807,N_7953);
xor U8088 (N_8088,N_7868,N_7962);
or U8089 (N_8089,N_7987,N_7823);
nor U8090 (N_8090,N_7917,N_7898);
or U8091 (N_8091,N_7902,N_7818);
or U8092 (N_8092,N_7952,N_7882);
nand U8093 (N_8093,N_7926,N_7885);
and U8094 (N_8094,N_7934,N_7989);
or U8095 (N_8095,N_7947,N_7859);
or U8096 (N_8096,N_7877,N_7840);
nor U8097 (N_8097,N_7872,N_7845);
and U8098 (N_8098,N_7826,N_7982);
xor U8099 (N_8099,N_7965,N_7824);
or U8100 (N_8100,N_7939,N_7997);
and U8101 (N_8101,N_7834,N_7914);
nand U8102 (N_8102,N_7807,N_7923);
nor U8103 (N_8103,N_7922,N_7876);
nand U8104 (N_8104,N_7825,N_7940);
or U8105 (N_8105,N_7970,N_7898);
nand U8106 (N_8106,N_7994,N_7921);
and U8107 (N_8107,N_7945,N_7929);
xor U8108 (N_8108,N_7994,N_7937);
nand U8109 (N_8109,N_7926,N_7855);
xor U8110 (N_8110,N_7924,N_7868);
nand U8111 (N_8111,N_7968,N_7975);
or U8112 (N_8112,N_7826,N_7897);
nand U8113 (N_8113,N_7840,N_7957);
and U8114 (N_8114,N_7966,N_7910);
nor U8115 (N_8115,N_7889,N_7983);
or U8116 (N_8116,N_7821,N_7927);
or U8117 (N_8117,N_7965,N_7960);
xor U8118 (N_8118,N_7886,N_7904);
nor U8119 (N_8119,N_7939,N_7885);
xor U8120 (N_8120,N_7975,N_7998);
nor U8121 (N_8121,N_7873,N_7845);
nor U8122 (N_8122,N_7813,N_7810);
nand U8123 (N_8123,N_7812,N_7867);
nor U8124 (N_8124,N_7873,N_7996);
xnor U8125 (N_8125,N_7934,N_7912);
nand U8126 (N_8126,N_7880,N_7944);
and U8127 (N_8127,N_7951,N_7997);
nand U8128 (N_8128,N_7820,N_7928);
nand U8129 (N_8129,N_7875,N_7846);
xor U8130 (N_8130,N_7837,N_7863);
nor U8131 (N_8131,N_7875,N_7866);
or U8132 (N_8132,N_7814,N_7856);
and U8133 (N_8133,N_7861,N_7951);
or U8134 (N_8134,N_7927,N_7968);
and U8135 (N_8135,N_7885,N_7918);
xor U8136 (N_8136,N_7823,N_7969);
and U8137 (N_8137,N_7839,N_7959);
and U8138 (N_8138,N_7984,N_7818);
xnor U8139 (N_8139,N_7831,N_7818);
and U8140 (N_8140,N_7823,N_7926);
xnor U8141 (N_8141,N_7905,N_7957);
or U8142 (N_8142,N_7948,N_7812);
or U8143 (N_8143,N_7970,N_7935);
and U8144 (N_8144,N_7866,N_7837);
nor U8145 (N_8145,N_7893,N_7832);
and U8146 (N_8146,N_7921,N_7808);
and U8147 (N_8147,N_7969,N_7925);
and U8148 (N_8148,N_7964,N_7936);
nand U8149 (N_8149,N_7909,N_7875);
nand U8150 (N_8150,N_7898,N_7951);
xor U8151 (N_8151,N_7918,N_7845);
nand U8152 (N_8152,N_7947,N_7959);
nor U8153 (N_8153,N_7889,N_7828);
xnor U8154 (N_8154,N_7989,N_7858);
nor U8155 (N_8155,N_7976,N_7944);
nand U8156 (N_8156,N_7806,N_7936);
nand U8157 (N_8157,N_7980,N_7935);
xor U8158 (N_8158,N_7964,N_7807);
nor U8159 (N_8159,N_7924,N_7819);
xor U8160 (N_8160,N_7862,N_7875);
nand U8161 (N_8161,N_7816,N_7977);
xnor U8162 (N_8162,N_7972,N_7959);
nor U8163 (N_8163,N_7966,N_7806);
nand U8164 (N_8164,N_7828,N_7803);
nand U8165 (N_8165,N_7931,N_7977);
nand U8166 (N_8166,N_7978,N_7969);
or U8167 (N_8167,N_7930,N_7811);
or U8168 (N_8168,N_7896,N_7867);
nor U8169 (N_8169,N_7879,N_7955);
nor U8170 (N_8170,N_7822,N_7845);
or U8171 (N_8171,N_7882,N_7986);
xor U8172 (N_8172,N_7945,N_7853);
xnor U8173 (N_8173,N_7946,N_7836);
and U8174 (N_8174,N_7891,N_7897);
or U8175 (N_8175,N_7974,N_7955);
or U8176 (N_8176,N_7814,N_7968);
xnor U8177 (N_8177,N_7822,N_7936);
and U8178 (N_8178,N_7953,N_7997);
or U8179 (N_8179,N_7963,N_7900);
and U8180 (N_8180,N_7917,N_7950);
nor U8181 (N_8181,N_7874,N_7868);
or U8182 (N_8182,N_7989,N_7855);
or U8183 (N_8183,N_7921,N_7839);
xnor U8184 (N_8184,N_7838,N_7866);
nand U8185 (N_8185,N_7991,N_7973);
nand U8186 (N_8186,N_7923,N_7927);
and U8187 (N_8187,N_7934,N_7905);
nor U8188 (N_8188,N_7904,N_7976);
xnor U8189 (N_8189,N_7860,N_7872);
or U8190 (N_8190,N_7846,N_7845);
and U8191 (N_8191,N_7810,N_7968);
nor U8192 (N_8192,N_7837,N_7913);
nor U8193 (N_8193,N_7959,N_7997);
or U8194 (N_8194,N_7992,N_7851);
and U8195 (N_8195,N_7934,N_7893);
xor U8196 (N_8196,N_7906,N_7926);
xor U8197 (N_8197,N_7822,N_7847);
xor U8198 (N_8198,N_7890,N_7818);
or U8199 (N_8199,N_7956,N_7988);
nand U8200 (N_8200,N_8046,N_8100);
xnor U8201 (N_8201,N_8121,N_8055);
nor U8202 (N_8202,N_8184,N_8125);
nor U8203 (N_8203,N_8075,N_8033);
or U8204 (N_8204,N_8109,N_8183);
and U8205 (N_8205,N_8086,N_8032);
or U8206 (N_8206,N_8164,N_8110);
and U8207 (N_8207,N_8030,N_8188);
nor U8208 (N_8208,N_8167,N_8180);
nand U8209 (N_8209,N_8060,N_8077);
nor U8210 (N_8210,N_8002,N_8087);
or U8211 (N_8211,N_8088,N_8019);
xor U8212 (N_8212,N_8064,N_8127);
xor U8213 (N_8213,N_8049,N_8138);
and U8214 (N_8214,N_8153,N_8112);
xor U8215 (N_8215,N_8156,N_8043);
and U8216 (N_8216,N_8130,N_8016);
nor U8217 (N_8217,N_8027,N_8197);
nand U8218 (N_8218,N_8158,N_8007);
nand U8219 (N_8219,N_8124,N_8120);
and U8220 (N_8220,N_8089,N_8135);
nor U8221 (N_8221,N_8067,N_8041);
nor U8222 (N_8222,N_8042,N_8003);
and U8223 (N_8223,N_8131,N_8031);
or U8224 (N_8224,N_8050,N_8160);
nand U8225 (N_8225,N_8017,N_8079);
or U8226 (N_8226,N_8009,N_8061);
nand U8227 (N_8227,N_8181,N_8013);
nand U8228 (N_8228,N_8001,N_8172);
or U8229 (N_8229,N_8119,N_8146);
nor U8230 (N_8230,N_8157,N_8150);
nor U8231 (N_8231,N_8165,N_8068);
and U8232 (N_8232,N_8014,N_8114);
or U8233 (N_8233,N_8143,N_8054);
nand U8234 (N_8234,N_8170,N_8152);
or U8235 (N_8235,N_8113,N_8045);
or U8236 (N_8236,N_8091,N_8195);
nand U8237 (N_8237,N_8021,N_8093);
or U8238 (N_8238,N_8106,N_8192);
nand U8239 (N_8239,N_8111,N_8073);
nand U8240 (N_8240,N_8166,N_8015);
xnor U8241 (N_8241,N_8047,N_8059);
or U8242 (N_8242,N_8005,N_8026);
nor U8243 (N_8243,N_8175,N_8190);
and U8244 (N_8244,N_8115,N_8147);
or U8245 (N_8245,N_8107,N_8072);
xnor U8246 (N_8246,N_8025,N_8159);
or U8247 (N_8247,N_8070,N_8076);
and U8248 (N_8248,N_8140,N_8194);
nor U8249 (N_8249,N_8022,N_8116);
and U8250 (N_8250,N_8186,N_8085);
nand U8251 (N_8251,N_8034,N_8142);
or U8252 (N_8252,N_8139,N_8044);
nand U8253 (N_8253,N_8123,N_8023);
or U8254 (N_8254,N_8191,N_8171);
nor U8255 (N_8255,N_8105,N_8010);
or U8256 (N_8256,N_8169,N_8117);
nor U8257 (N_8257,N_8092,N_8144);
nor U8258 (N_8258,N_8038,N_8168);
and U8259 (N_8259,N_8126,N_8128);
nor U8260 (N_8260,N_8199,N_8048);
and U8261 (N_8261,N_8074,N_8102);
nand U8262 (N_8262,N_8094,N_8163);
nand U8263 (N_8263,N_8040,N_8057);
and U8264 (N_8264,N_8193,N_8069);
nand U8265 (N_8265,N_8103,N_8162);
nor U8266 (N_8266,N_8006,N_8177);
nand U8267 (N_8267,N_8000,N_8136);
nor U8268 (N_8268,N_8004,N_8185);
xor U8269 (N_8269,N_8036,N_8149);
nor U8270 (N_8270,N_8118,N_8051);
xor U8271 (N_8271,N_8104,N_8062);
and U8272 (N_8272,N_8176,N_8066);
nand U8273 (N_8273,N_8098,N_8161);
nor U8274 (N_8274,N_8134,N_8024);
nor U8275 (N_8275,N_8011,N_8012);
xor U8276 (N_8276,N_8174,N_8129);
nor U8277 (N_8277,N_8178,N_8122);
or U8278 (N_8278,N_8039,N_8028);
nor U8279 (N_8279,N_8037,N_8083);
or U8280 (N_8280,N_8155,N_8052);
and U8281 (N_8281,N_8084,N_8053);
nor U8282 (N_8282,N_8065,N_8029);
nand U8283 (N_8283,N_8101,N_8090);
xor U8284 (N_8284,N_8056,N_8071);
or U8285 (N_8285,N_8078,N_8081);
or U8286 (N_8286,N_8148,N_8196);
nor U8287 (N_8287,N_8182,N_8058);
or U8288 (N_8288,N_8189,N_8133);
xor U8289 (N_8289,N_8132,N_8187);
nor U8290 (N_8290,N_8096,N_8020);
and U8291 (N_8291,N_8099,N_8018);
nor U8292 (N_8292,N_8082,N_8154);
nand U8293 (N_8293,N_8095,N_8108);
nor U8294 (N_8294,N_8035,N_8141);
or U8295 (N_8295,N_8198,N_8097);
nor U8296 (N_8296,N_8008,N_8179);
nor U8297 (N_8297,N_8063,N_8080);
nand U8298 (N_8298,N_8137,N_8145);
nor U8299 (N_8299,N_8173,N_8151);
and U8300 (N_8300,N_8121,N_8112);
nand U8301 (N_8301,N_8001,N_8169);
and U8302 (N_8302,N_8063,N_8131);
nand U8303 (N_8303,N_8147,N_8043);
nand U8304 (N_8304,N_8110,N_8142);
xnor U8305 (N_8305,N_8180,N_8056);
nand U8306 (N_8306,N_8066,N_8140);
nand U8307 (N_8307,N_8004,N_8092);
xnor U8308 (N_8308,N_8040,N_8053);
or U8309 (N_8309,N_8040,N_8158);
xnor U8310 (N_8310,N_8054,N_8107);
and U8311 (N_8311,N_8196,N_8186);
and U8312 (N_8312,N_8100,N_8101);
and U8313 (N_8313,N_8013,N_8016);
nor U8314 (N_8314,N_8190,N_8012);
and U8315 (N_8315,N_8133,N_8047);
xnor U8316 (N_8316,N_8060,N_8151);
nand U8317 (N_8317,N_8191,N_8129);
nand U8318 (N_8318,N_8075,N_8097);
and U8319 (N_8319,N_8124,N_8123);
or U8320 (N_8320,N_8182,N_8193);
and U8321 (N_8321,N_8166,N_8134);
nor U8322 (N_8322,N_8132,N_8056);
and U8323 (N_8323,N_8131,N_8199);
or U8324 (N_8324,N_8020,N_8149);
or U8325 (N_8325,N_8176,N_8159);
xnor U8326 (N_8326,N_8049,N_8000);
and U8327 (N_8327,N_8163,N_8165);
nand U8328 (N_8328,N_8035,N_8118);
or U8329 (N_8329,N_8004,N_8035);
or U8330 (N_8330,N_8161,N_8024);
nand U8331 (N_8331,N_8123,N_8052);
nor U8332 (N_8332,N_8104,N_8057);
and U8333 (N_8333,N_8150,N_8133);
and U8334 (N_8334,N_8009,N_8085);
or U8335 (N_8335,N_8163,N_8173);
nand U8336 (N_8336,N_8017,N_8077);
and U8337 (N_8337,N_8070,N_8128);
nand U8338 (N_8338,N_8027,N_8073);
and U8339 (N_8339,N_8039,N_8121);
and U8340 (N_8340,N_8195,N_8084);
or U8341 (N_8341,N_8185,N_8014);
nor U8342 (N_8342,N_8143,N_8130);
xnor U8343 (N_8343,N_8177,N_8166);
and U8344 (N_8344,N_8165,N_8186);
and U8345 (N_8345,N_8167,N_8085);
nor U8346 (N_8346,N_8133,N_8093);
xor U8347 (N_8347,N_8131,N_8082);
or U8348 (N_8348,N_8017,N_8136);
xnor U8349 (N_8349,N_8043,N_8039);
and U8350 (N_8350,N_8153,N_8141);
nand U8351 (N_8351,N_8103,N_8017);
nor U8352 (N_8352,N_8039,N_8130);
xor U8353 (N_8353,N_8166,N_8121);
nor U8354 (N_8354,N_8001,N_8185);
or U8355 (N_8355,N_8028,N_8140);
nand U8356 (N_8356,N_8155,N_8035);
or U8357 (N_8357,N_8082,N_8145);
nand U8358 (N_8358,N_8035,N_8038);
or U8359 (N_8359,N_8021,N_8136);
and U8360 (N_8360,N_8101,N_8008);
or U8361 (N_8361,N_8068,N_8051);
or U8362 (N_8362,N_8041,N_8141);
xor U8363 (N_8363,N_8128,N_8099);
or U8364 (N_8364,N_8146,N_8044);
nor U8365 (N_8365,N_8083,N_8094);
nor U8366 (N_8366,N_8125,N_8162);
xor U8367 (N_8367,N_8176,N_8075);
nand U8368 (N_8368,N_8082,N_8113);
nand U8369 (N_8369,N_8106,N_8082);
or U8370 (N_8370,N_8129,N_8141);
or U8371 (N_8371,N_8005,N_8014);
xor U8372 (N_8372,N_8032,N_8193);
xor U8373 (N_8373,N_8043,N_8182);
or U8374 (N_8374,N_8051,N_8034);
nor U8375 (N_8375,N_8035,N_8071);
and U8376 (N_8376,N_8101,N_8093);
or U8377 (N_8377,N_8165,N_8024);
nand U8378 (N_8378,N_8135,N_8184);
and U8379 (N_8379,N_8144,N_8128);
nor U8380 (N_8380,N_8130,N_8035);
nand U8381 (N_8381,N_8011,N_8029);
nand U8382 (N_8382,N_8046,N_8055);
and U8383 (N_8383,N_8120,N_8107);
xnor U8384 (N_8384,N_8068,N_8064);
xor U8385 (N_8385,N_8181,N_8176);
or U8386 (N_8386,N_8083,N_8044);
or U8387 (N_8387,N_8128,N_8059);
and U8388 (N_8388,N_8025,N_8069);
and U8389 (N_8389,N_8028,N_8080);
nand U8390 (N_8390,N_8174,N_8128);
or U8391 (N_8391,N_8016,N_8193);
or U8392 (N_8392,N_8131,N_8020);
nor U8393 (N_8393,N_8192,N_8054);
nand U8394 (N_8394,N_8000,N_8110);
xnor U8395 (N_8395,N_8123,N_8185);
nand U8396 (N_8396,N_8049,N_8156);
nor U8397 (N_8397,N_8137,N_8008);
nor U8398 (N_8398,N_8138,N_8130);
and U8399 (N_8399,N_8084,N_8178);
nor U8400 (N_8400,N_8382,N_8245);
nor U8401 (N_8401,N_8304,N_8225);
or U8402 (N_8402,N_8275,N_8386);
nand U8403 (N_8403,N_8301,N_8265);
nor U8404 (N_8404,N_8292,N_8278);
xor U8405 (N_8405,N_8374,N_8360);
nor U8406 (N_8406,N_8205,N_8237);
and U8407 (N_8407,N_8223,N_8221);
or U8408 (N_8408,N_8350,N_8238);
nand U8409 (N_8409,N_8321,N_8342);
or U8410 (N_8410,N_8282,N_8334);
nand U8411 (N_8411,N_8210,N_8220);
nor U8412 (N_8412,N_8370,N_8222);
nand U8413 (N_8413,N_8212,N_8327);
and U8414 (N_8414,N_8390,N_8291);
nor U8415 (N_8415,N_8371,N_8317);
nand U8416 (N_8416,N_8315,N_8217);
nand U8417 (N_8417,N_8219,N_8295);
xnor U8418 (N_8418,N_8293,N_8239);
nor U8419 (N_8419,N_8369,N_8358);
nand U8420 (N_8420,N_8284,N_8266);
and U8421 (N_8421,N_8272,N_8251);
and U8422 (N_8422,N_8318,N_8280);
or U8423 (N_8423,N_8394,N_8381);
nand U8424 (N_8424,N_8224,N_8269);
xor U8425 (N_8425,N_8355,N_8336);
nand U8426 (N_8426,N_8395,N_8385);
and U8427 (N_8427,N_8388,N_8380);
and U8428 (N_8428,N_8240,N_8283);
nand U8429 (N_8429,N_8201,N_8367);
or U8430 (N_8430,N_8271,N_8325);
and U8431 (N_8431,N_8285,N_8247);
nand U8432 (N_8432,N_8333,N_8242);
and U8433 (N_8433,N_8324,N_8236);
nor U8434 (N_8434,N_8302,N_8288);
nor U8435 (N_8435,N_8377,N_8303);
nor U8436 (N_8436,N_8299,N_8320);
xnor U8437 (N_8437,N_8264,N_8308);
xor U8438 (N_8438,N_8313,N_8351);
nor U8439 (N_8439,N_8379,N_8286);
and U8440 (N_8440,N_8384,N_8228);
nor U8441 (N_8441,N_8366,N_8215);
xor U8442 (N_8442,N_8345,N_8204);
xnor U8443 (N_8443,N_8289,N_8391);
xnor U8444 (N_8444,N_8259,N_8202);
or U8445 (N_8445,N_8241,N_8393);
xnor U8446 (N_8446,N_8372,N_8218);
or U8447 (N_8447,N_8263,N_8294);
xnor U8448 (N_8448,N_8352,N_8387);
xnor U8449 (N_8449,N_8314,N_8298);
and U8450 (N_8450,N_8338,N_8392);
xor U8451 (N_8451,N_8396,N_8311);
or U8452 (N_8452,N_8211,N_8214);
nor U8453 (N_8453,N_8362,N_8276);
and U8454 (N_8454,N_8312,N_8273);
and U8455 (N_8455,N_8375,N_8208);
xor U8456 (N_8456,N_8340,N_8346);
and U8457 (N_8457,N_8353,N_8328);
xnor U8458 (N_8458,N_8256,N_8364);
or U8459 (N_8459,N_8383,N_8307);
nor U8460 (N_8460,N_8207,N_8365);
nand U8461 (N_8461,N_8330,N_8234);
nor U8462 (N_8462,N_8258,N_8373);
nand U8463 (N_8463,N_8279,N_8398);
or U8464 (N_8464,N_8244,N_8248);
nand U8465 (N_8465,N_8357,N_8235);
nand U8466 (N_8466,N_8243,N_8343);
nor U8467 (N_8467,N_8354,N_8213);
nand U8468 (N_8468,N_8332,N_8230);
nor U8469 (N_8469,N_8297,N_8233);
nor U8470 (N_8470,N_8339,N_8277);
and U8471 (N_8471,N_8287,N_8376);
nor U8472 (N_8472,N_8254,N_8310);
xnor U8473 (N_8473,N_8267,N_8347);
xnor U8474 (N_8474,N_8368,N_8261);
nand U8475 (N_8475,N_8399,N_8363);
nor U8476 (N_8476,N_8356,N_8227);
xnor U8477 (N_8477,N_8257,N_8326);
or U8478 (N_8478,N_8337,N_8323);
or U8479 (N_8479,N_8232,N_8226);
xnor U8480 (N_8480,N_8335,N_8319);
xnor U8481 (N_8481,N_8270,N_8252);
nor U8482 (N_8482,N_8246,N_8200);
nor U8483 (N_8483,N_8348,N_8296);
and U8484 (N_8484,N_8389,N_8305);
nor U8485 (N_8485,N_8359,N_8361);
nand U8486 (N_8486,N_8344,N_8253);
or U8487 (N_8487,N_8231,N_8203);
or U8488 (N_8488,N_8206,N_8349);
and U8489 (N_8489,N_8378,N_8274);
nand U8490 (N_8490,N_8300,N_8209);
or U8491 (N_8491,N_8329,N_8262);
nand U8492 (N_8492,N_8309,N_8260);
or U8493 (N_8493,N_8249,N_8397);
and U8494 (N_8494,N_8316,N_8331);
or U8495 (N_8495,N_8322,N_8255);
nand U8496 (N_8496,N_8341,N_8216);
xnor U8497 (N_8497,N_8281,N_8250);
nand U8498 (N_8498,N_8290,N_8229);
nor U8499 (N_8499,N_8306,N_8268);
nor U8500 (N_8500,N_8362,N_8339);
nor U8501 (N_8501,N_8300,N_8268);
nor U8502 (N_8502,N_8383,N_8338);
xnor U8503 (N_8503,N_8327,N_8234);
or U8504 (N_8504,N_8306,N_8292);
nand U8505 (N_8505,N_8364,N_8210);
nor U8506 (N_8506,N_8278,N_8263);
nor U8507 (N_8507,N_8324,N_8263);
xor U8508 (N_8508,N_8209,N_8396);
xnor U8509 (N_8509,N_8328,N_8391);
and U8510 (N_8510,N_8377,N_8227);
nor U8511 (N_8511,N_8215,N_8279);
or U8512 (N_8512,N_8221,N_8239);
nand U8513 (N_8513,N_8298,N_8344);
or U8514 (N_8514,N_8366,N_8263);
or U8515 (N_8515,N_8222,N_8238);
or U8516 (N_8516,N_8398,N_8218);
nand U8517 (N_8517,N_8344,N_8200);
xor U8518 (N_8518,N_8359,N_8324);
or U8519 (N_8519,N_8242,N_8229);
and U8520 (N_8520,N_8282,N_8226);
nor U8521 (N_8521,N_8249,N_8263);
xnor U8522 (N_8522,N_8359,N_8261);
and U8523 (N_8523,N_8349,N_8393);
and U8524 (N_8524,N_8217,N_8306);
nor U8525 (N_8525,N_8292,N_8385);
nand U8526 (N_8526,N_8292,N_8265);
or U8527 (N_8527,N_8347,N_8274);
or U8528 (N_8528,N_8253,N_8247);
nor U8529 (N_8529,N_8232,N_8241);
and U8530 (N_8530,N_8317,N_8343);
xor U8531 (N_8531,N_8271,N_8219);
and U8532 (N_8532,N_8269,N_8339);
xnor U8533 (N_8533,N_8308,N_8212);
and U8534 (N_8534,N_8241,N_8376);
and U8535 (N_8535,N_8355,N_8251);
xnor U8536 (N_8536,N_8309,N_8335);
nand U8537 (N_8537,N_8282,N_8213);
nand U8538 (N_8538,N_8269,N_8382);
or U8539 (N_8539,N_8223,N_8306);
xnor U8540 (N_8540,N_8312,N_8265);
nor U8541 (N_8541,N_8385,N_8209);
xnor U8542 (N_8542,N_8203,N_8288);
and U8543 (N_8543,N_8295,N_8352);
xor U8544 (N_8544,N_8312,N_8207);
nor U8545 (N_8545,N_8331,N_8246);
xor U8546 (N_8546,N_8247,N_8292);
nor U8547 (N_8547,N_8365,N_8359);
and U8548 (N_8548,N_8373,N_8392);
nand U8549 (N_8549,N_8228,N_8247);
nor U8550 (N_8550,N_8330,N_8363);
nand U8551 (N_8551,N_8241,N_8224);
or U8552 (N_8552,N_8297,N_8261);
nand U8553 (N_8553,N_8311,N_8203);
nand U8554 (N_8554,N_8365,N_8256);
xnor U8555 (N_8555,N_8347,N_8378);
and U8556 (N_8556,N_8217,N_8270);
xor U8557 (N_8557,N_8262,N_8220);
and U8558 (N_8558,N_8395,N_8234);
xor U8559 (N_8559,N_8230,N_8274);
xnor U8560 (N_8560,N_8302,N_8371);
and U8561 (N_8561,N_8202,N_8352);
and U8562 (N_8562,N_8254,N_8201);
or U8563 (N_8563,N_8369,N_8285);
and U8564 (N_8564,N_8380,N_8360);
and U8565 (N_8565,N_8398,N_8377);
and U8566 (N_8566,N_8215,N_8302);
or U8567 (N_8567,N_8341,N_8203);
xnor U8568 (N_8568,N_8382,N_8384);
xnor U8569 (N_8569,N_8206,N_8240);
and U8570 (N_8570,N_8326,N_8223);
and U8571 (N_8571,N_8312,N_8344);
nor U8572 (N_8572,N_8241,N_8311);
nor U8573 (N_8573,N_8208,N_8399);
nand U8574 (N_8574,N_8287,N_8398);
and U8575 (N_8575,N_8287,N_8204);
or U8576 (N_8576,N_8290,N_8369);
nor U8577 (N_8577,N_8348,N_8391);
nand U8578 (N_8578,N_8275,N_8330);
nor U8579 (N_8579,N_8376,N_8382);
xnor U8580 (N_8580,N_8335,N_8367);
nand U8581 (N_8581,N_8304,N_8349);
xor U8582 (N_8582,N_8299,N_8349);
nor U8583 (N_8583,N_8211,N_8339);
xor U8584 (N_8584,N_8263,N_8280);
xor U8585 (N_8585,N_8233,N_8239);
xor U8586 (N_8586,N_8257,N_8375);
xnor U8587 (N_8587,N_8375,N_8232);
nor U8588 (N_8588,N_8233,N_8350);
nand U8589 (N_8589,N_8250,N_8360);
nor U8590 (N_8590,N_8366,N_8283);
nand U8591 (N_8591,N_8344,N_8394);
and U8592 (N_8592,N_8200,N_8275);
xor U8593 (N_8593,N_8315,N_8280);
or U8594 (N_8594,N_8260,N_8323);
nand U8595 (N_8595,N_8394,N_8300);
or U8596 (N_8596,N_8200,N_8282);
and U8597 (N_8597,N_8302,N_8365);
xor U8598 (N_8598,N_8357,N_8359);
and U8599 (N_8599,N_8394,N_8245);
nor U8600 (N_8600,N_8417,N_8522);
or U8601 (N_8601,N_8589,N_8455);
and U8602 (N_8602,N_8518,N_8565);
xor U8603 (N_8603,N_8468,N_8456);
nor U8604 (N_8604,N_8594,N_8496);
nor U8605 (N_8605,N_8517,N_8527);
or U8606 (N_8606,N_8436,N_8563);
nor U8607 (N_8607,N_8545,N_8407);
xnor U8608 (N_8608,N_8444,N_8543);
nand U8609 (N_8609,N_8479,N_8454);
and U8610 (N_8610,N_8464,N_8427);
nor U8611 (N_8611,N_8569,N_8449);
nor U8612 (N_8612,N_8447,N_8445);
xnor U8613 (N_8613,N_8596,N_8473);
or U8614 (N_8614,N_8423,N_8548);
and U8615 (N_8615,N_8549,N_8512);
nor U8616 (N_8616,N_8526,N_8583);
or U8617 (N_8617,N_8511,N_8421);
and U8618 (N_8618,N_8426,N_8475);
xor U8619 (N_8619,N_8520,N_8422);
nor U8620 (N_8620,N_8480,N_8439);
nor U8621 (N_8621,N_8494,N_8516);
xnor U8622 (N_8622,N_8528,N_8478);
xnor U8623 (N_8623,N_8443,N_8579);
xnor U8624 (N_8624,N_8587,N_8466);
nand U8625 (N_8625,N_8508,N_8469);
and U8626 (N_8626,N_8578,N_8585);
xnor U8627 (N_8627,N_8487,N_8428);
and U8628 (N_8628,N_8538,N_8448);
nand U8629 (N_8629,N_8539,N_8581);
xor U8630 (N_8630,N_8550,N_8547);
and U8631 (N_8631,N_8425,N_8413);
nand U8632 (N_8632,N_8523,N_8483);
xnor U8633 (N_8633,N_8577,N_8574);
or U8634 (N_8634,N_8442,N_8534);
or U8635 (N_8635,N_8403,N_8412);
and U8636 (N_8636,N_8476,N_8564);
nand U8637 (N_8637,N_8529,N_8580);
and U8638 (N_8638,N_8513,N_8459);
or U8639 (N_8639,N_8544,N_8586);
or U8640 (N_8640,N_8499,N_8558);
nand U8641 (N_8641,N_8410,N_8530);
nor U8642 (N_8642,N_8493,N_8561);
xor U8643 (N_8643,N_8429,N_8582);
xor U8644 (N_8644,N_8507,N_8562);
nand U8645 (N_8645,N_8482,N_8457);
or U8646 (N_8646,N_8572,N_8568);
nand U8647 (N_8647,N_8418,N_8595);
nor U8648 (N_8648,N_8424,N_8575);
nand U8649 (N_8649,N_8566,N_8465);
nor U8650 (N_8650,N_8438,N_8519);
and U8651 (N_8651,N_8495,N_8419);
xnor U8652 (N_8652,N_8411,N_8515);
and U8653 (N_8653,N_8584,N_8446);
and U8654 (N_8654,N_8488,N_8450);
or U8655 (N_8655,N_8540,N_8441);
or U8656 (N_8656,N_8567,N_8555);
nand U8657 (N_8657,N_8591,N_8597);
nand U8658 (N_8658,N_8431,N_8477);
or U8659 (N_8659,N_8505,N_8541);
nand U8660 (N_8660,N_8420,N_8461);
or U8661 (N_8661,N_8560,N_8551);
nor U8662 (N_8662,N_8492,N_8504);
nand U8663 (N_8663,N_8452,N_8434);
xor U8664 (N_8664,N_8481,N_8546);
or U8665 (N_8665,N_8533,N_8430);
or U8666 (N_8666,N_8532,N_8462);
nand U8667 (N_8667,N_8474,N_8451);
nor U8668 (N_8668,N_8590,N_8470);
nor U8669 (N_8669,N_8460,N_8401);
nor U8670 (N_8670,N_8571,N_8491);
nand U8671 (N_8671,N_8542,N_8593);
and U8672 (N_8672,N_8506,N_8573);
xor U8673 (N_8673,N_8524,N_8514);
and U8674 (N_8674,N_8502,N_8489);
and U8675 (N_8675,N_8435,N_8498);
xor U8676 (N_8676,N_8463,N_8556);
xor U8677 (N_8677,N_8433,N_8485);
or U8678 (N_8678,N_8453,N_8576);
nand U8679 (N_8679,N_8559,N_8432);
xor U8680 (N_8680,N_8437,N_8408);
nand U8681 (N_8681,N_8471,N_8503);
nand U8682 (N_8682,N_8592,N_8409);
or U8683 (N_8683,N_8501,N_8406);
nor U8684 (N_8684,N_8405,N_8414);
and U8685 (N_8685,N_8554,N_8552);
nor U8686 (N_8686,N_8440,N_8510);
xnor U8687 (N_8687,N_8484,N_8416);
nand U8688 (N_8688,N_8415,N_8588);
and U8689 (N_8689,N_8531,N_8402);
nor U8690 (N_8690,N_8570,N_8490);
nand U8691 (N_8691,N_8500,N_8598);
nor U8692 (N_8692,N_8497,N_8536);
or U8693 (N_8693,N_8472,N_8521);
or U8694 (N_8694,N_8486,N_8537);
xnor U8695 (N_8695,N_8553,N_8535);
xor U8696 (N_8696,N_8557,N_8458);
nor U8697 (N_8697,N_8404,N_8525);
nand U8698 (N_8698,N_8400,N_8509);
nand U8699 (N_8699,N_8467,N_8599);
nor U8700 (N_8700,N_8592,N_8564);
nor U8701 (N_8701,N_8485,N_8522);
nand U8702 (N_8702,N_8515,N_8480);
xnor U8703 (N_8703,N_8487,N_8473);
and U8704 (N_8704,N_8452,N_8441);
and U8705 (N_8705,N_8438,N_8521);
nand U8706 (N_8706,N_8430,N_8510);
or U8707 (N_8707,N_8559,N_8405);
and U8708 (N_8708,N_8449,N_8475);
xor U8709 (N_8709,N_8482,N_8519);
xor U8710 (N_8710,N_8428,N_8491);
nand U8711 (N_8711,N_8416,N_8466);
or U8712 (N_8712,N_8505,N_8483);
xnor U8713 (N_8713,N_8477,N_8503);
nor U8714 (N_8714,N_8443,N_8577);
nand U8715 (N_8715,N_8423,N_8416);
and U8716 (N_8716,N_8448,N_8460);
xnor U8717 (N_8717,N_8541,N_8597);
xor U8718 (N_8718,N_8527,N_8504);
nor U8719 (N_8719,N_8466,N_8582);
or U8720 (N_8720,N_8589,N_8484);
and U8721 (N_8721,N_8573,N_8542);
and U8722 (N_8722,N_8412,N_8446);
nand U8723 (N_8723,N_8466,N_8406);
xor U8724 (N_8724,N_8513,N_8522);
xnor U8725 (N_8725,N_8479,N_8471);
nand U8726 (N_8726,N_8557,N_8464);
nand U8727 (N_8727,N_8457,N_8416);
nor U8728 (N_8728,N_8465,N_8571);
xor U8729 (N_8729,N_8512,N_8499);
or U8730 (N_8730,N_8521,N_8487);
or U8731 (N_8731,N_8481,N_8465);
or U8732 (N_8732,N_8499,N_8536);
or U8733 (N_8733,N_8471,N_8452);
nand U8734 (N_8734,N_8444,N_8402);
nand U8735 (N_8735,N_8458,N_8510);
xor U8736 (N_8736,N_8415,N_8548);
nand U8737 (N_8737,N_8410,N_8521);
nand U8738 (N_8738,N_8553,N_8547);
xor U8739 (N_8739,N_8594,N_8472);
nor U8740 (N_8740,N_8505,N_8488);
xnor U8741 (N_8741,N_8564,N_8473);
xnor U8742 (N_8742,N_8463,N_8426);
xor U8743 (N_8743,N_8486,N_8569);
or U8744 (N_8744,N_8411,N_8437);
xnor U8745 (N_8745,N_8534,N_8408);
nor U8746 (N_8746,N_8534,N_8527);
nor U8747 (N_8747,N_8403,N_8508);
or U8748 (N_8748,N_8475,N_8529);
xor U8749 (N_8749,N_8540,N_8522);
and U8750 (N_8750,N_8477,N_8454);
xor U8751 (N_8751,N_8472,N_8460);
or U8752 (N_8752,N_8530,N_8525);
and U8753 (N_8753,N_8561,N_8586);
or U8754 (N_8754,N_8497,N_8552);
nand U8755 (N_8755,N_8589,N_8513);
nor U8756 (N_8756,N_8479,N_8510);
nand U8757 (N_8757,N_8430,N_8477);
or U8758 (N_8758,N_8485,N_8545);
nand U8759 (N_8759,N_8492,N_8519);
or U8760 (N_8760,N_8511,N_8561);
nor U8761 (N_8761,N_8405,N_8513);
and U8762 (N_8762,N_8485,N_8507);
nand U8763 (N_8763,N_8577,N_8546);
or U8764 (N_8764,N_8401,N_8420);
or U8765 (N_8765,N_8592,N_8544);
nand U8766 (N_8766,N_8531,N_8492);
xor U8767 (N_8767,N_8403,N_8407);
and U8768 (N_8768,N_8483,N_8537);
and U8769 (N_8769,N_8471,N_8415);
and U8770 (N_8770,N_8434,N_8589);
and U8771 (N_8771,N_8432,N_8437);
and U8772 (N_8772,N_8450,N_8580);
xor U8773 (N_8773,N_8437,N_8582);
or U8774 (N_8774,N_8490,N_8419);
nand U8775 (N_8775,N_8537,N_8478);
nand U8776 (N_8776,N_8508,N_8493);
nor U8777 (N_8777,N_8587,N_8477);
nor U8778 (N_8778,N_8522,N_8495);
nand U8779 (N_8779,N_8539,N_8459);
nor U8780 (N_8780,N_8443,N_8468);
xnor U8781 (N_8781,N_8437,N_8440);
and U8782 (N_8782,N_8578,N_8531);
nand U8783 (N_8783,N_8553,N_8512);
xor U8784 (N_8784,N_8434,N_8585);
nor U8785 (N_8785,N_8513,N_8508);
nand U8786 (N_8786,N_8472,N_8592);
and U8787 (N_8787,N_8552,N_8540);
nand U8788 (N_8788,N_8408,N_8423);
xor U8789 (N_8789,N_8411,N_8586);
nor U8790 (N_8790,N_8595,N_8404);
nor U8791 (N_8791,N_8432,N_8598);
and U8792 (N_8792,N_8577,N_8404);
or U8793 (N_8793,N_8486,N_8490);
or U8794 (N_8794,N_8592,N_8560);
or U8795 (N_8795,N_8451,N_8503);
nor U8796 (N_8796,N_8575,N_8404);
and U8797 (N_8797,N_8416,N_8495);
and U8798 (N_8798,N_8431,N_8496);
nand U8799 (N_8799,N_8569,N_8462);
or U8800 (N_8800,N_8698,N_8710);
xnor U8801 (N_8801,N_8657,N_8675);
nor U8802 (N_8802,N_8750,N_8606);
nand U8803 (N_8803,N_8737,N_8696);
and U8804 (N_8804,N_8795,N_8684);
nand U8805 (N_8805,N_8686,N_8605);
nand U8806 (N_8806,N_8661,N_8751);
xnor U8807 (N_8807,N_8678,N_8631);
xor U8808 (N_8808,N_8726,N_8730);
nor U8809 (N_8809,N_8702,N_8646);
or U8810 (N_8810,N_8797,N_8739);
nand U8811 (N_8811,N_8611,N_8765);
or U8812 (N_8812,N_8782,N_8786);
and U8813 (N_8813,N_8766,N_8796);
or U8814 (N_8814,N_8602,N_8798);
and U8815 (N_8815,N_8793,N_8663);
xor U8816 (N_8816,N_8719,N_8683);
nor U8817 (N_8817,N_8637,N_8682);
and U8818 (N_8818,N_8672,N_8731);
nor U8819 (N_8819,N_8764,N_8665);
and U8820 (N_8820,N_8771,N_8620);
nand U8821 (N_8821,N_8770,N_8621);
and U8822 (N_8822,N_8768,N_8775);
and U8823 (N_8823,N_8670,N_8639);
or U8824 (N_8824,N_8667,N_8741);
or U8825 (N_8825,N_8651,N_8718);
or U8826 (N_8826,N_8674,N_8788);
or U8827 (N_8827,N_8619,N_8607);
xor U8828 (N_8828,N_8688,N_8618);
nor U8829 (N_8829,N_8625,N_8627);
xor U8830 (N_8830,N_8794,N_8790);
nand U8831 (N_8831,N_8642,N_8626);
or U8832 (N_8832,N_8650,N_8753);
or U8833 (N_8833,N_8700,N_8748);
nand U8834 (N_8834,N_8769,N_8729);
xnor U8835 (N_8835,N_8640,N_8629);
xor U8836 (N_8836,N_8755,N_8761);
nor U8837 (N_8837,N_8694,N_8773);
nor U8838 (N_8838,N_8711,N_8612);
xor U8839 (N_8839,N_8638,N_8772);
and U8840 (N_8840,N_8704,N_8701);
nand U8841 (N_8841,N_8722,N_8756);
and U8842 (N_8842,N_8630,N_8655);
and U8843 (N_8843,N_8649,N_8777);
and U8844 (N_8844,N_8617,N_8656);
nand U8845 (N_8845,N_8643,N_8789);
nor U8846 (N_8846,N_8762,N_8784);
or U8847 (N_8847,N_8636,N_8624);
nand U8848 (N_8848,N_8633,N_8660);
nand U8849 (N_8849,N_8615,N_8600);
nor U8850 (N_8850,N_8743,N_8690);
nor U8851 (N_8851,N_8705,N_8634);
nand U8852 (N_8852,N_8767,N_8680);
nand U8853 (N_8853,N_8717,N_8608);
and U8854 (N_8854,N_8779,N_8783);
nor U8855 (N_8855,N_8699,N_8774);
nand U8856 (N_8856,N_8734,N_8740);
xnor U8857 (N_8857,N_8628,N_8776);
and U8858 (N_8858,N_8635,N_8644);
and U8859 (N_8859,N_8679,N_8736);
nor U8860 (N_8860,N_8623,N_8645);
or U8861 (N_8861,N_8721,N_8652);
xor U8862 (N_8862,N_8759,N_8723);
nor U8863 (N_8863,N_8780,N_8695);
and U8864 (N_8864,N_8799,N_8791);
nor U8865 (N_8865,N_8760,N_8662);
nand U8866 (N_8866,N_8744,N_8677);
nand U8867 (N_8867,N_8610,N_8714);
or U8868 (N_8868,N_8671,N_8715);
or U8869 (N_8869,N_8745,N_8632);
xnor U8870 (N_8870,N_8727,N_8720);
and U8871 (N_8871,N_8706,N_8616);
or U8872 (N_8872,N_8622,N_8747);
and U8873 (N_8873,N_8738,N_8754);
and U8874 (N_8874,N_8707,N_8654);
nor U8875 (N_8875,N_8733,N_8687);
and U8876 (N_8876,N_8692,N_8691);
nor U8877 (N_8877,N_8735,N_8658);
or U8878 (N_8878,N_8712,N_8746);
or U8879 (N_8879,N_8778,N_8659);
xnor U8880 (N_8880,N_8725,N_8693);
xnor U8881 (N_8881,N_8666,N_8732);
nor U8882 (N_8882,N_8641,N_8787);
or U8883 (N_8883,N_8604,N_8653);
nand U8884 (N_8884,N_8792,N_8647);
xnor U8885 (N_8885,N_8758,N_8708);
xor U8886 (N_8886,N_8664,N_8689);
or U8887 (N_8887,N_8781,N_8763);
and U8888 (N_8888,N_8757,N_8601);
xnor U8889 (N_8889,N_8673,N_8685);
nor U8890 (N_8890,N_8713,N_8648);
xor U8891 (N_8891,N_8676,N_8724);
xnor U8892 (N_8892,N_8681,N_8669);
or U8893 (N_8893,N_8703,N_8668);
nand U8894 (N_8894,N_8603,N_8613);
xor U8895 (N_8895,N_8614,N_8609);
and U8896 (N_8896,N_8709,N_8728);
xor U8897 (N_8897,N_8785,N_8697);
xnor U8898 (N_8898,N_8716,N_8752);
nand U8899 (N_8899,N_8749,N_8742);
nor U8900 (N_8900,N_8759,N_8672);
and U8901 (N_8901,N_8765,N_8783);
nor U8902 (N_8902,N_8794,N_8791);
or U8903 (N_8903,N_8633,N_8788);
xnor U8904 (N_8904,N_8679,N_8606);
and U8905 (N_8905,N_8774,N_8625);
or U8906 (N_8906,N_8766,N_8780);
or U8907 (N_8907,N_8773,N_8702);
nor U8908 (N_8908,N_8603,N_8716);
or U8909 (N_8909,N_8673,N_8628);
nand U8910 (N_8910,N_8745,N_8790);
nand U8911 (N_8911,N_8640,N_8675);
nor U8912 (N_8912,N_8650,N_8622);
and U8913 (N_8913,N_8798,N_8752);
nand U8914 (N_8914,N_8745,N_8742);
xnor U8915 (N_8915,N_8677,N_8680);
and U8916 (N_8916,N_8733,N_8679);
or U8917 (N_8917,N_8642,N_8654);
and U8918 (N_8918,N_8725,N_8638);
or U8919 (N_8919,N_8743,N_8622);
or U8920 (N_8920,N_8796,N_8759);
nand U8921 (N_8921,N_8762,N_8733);
xor U8922 (N_8922,N_8605,N_8676);
nor U8923 (N_8923,N_8632,N_8643);
and U8924 (N_8924,N_8734,N_8775);
nor U8925 (N_8925,N_8678,N_8691);
or U8926 (N_8926,N_8788,N_8608);
or U8927 (N_8927,N_8756,N_8603);
nor U8928 (N_8928,N_8736,N_8739);
nor U8929 (N_8929,N_8791,N_8615);
and U8930 (N_8930,N_8615,N_8724);
xnor U8931 (N_8931,N_8665,N_8787);
and U8932 (N_8932,N_8667,N_8628);
or U8933 (N_8933,N_8775,N_8670);
and U8934 (N_8934,N_8784,N_8719);
nand U8935 (N_8935,N_8731,N_8640);
nor U8936 (N_8936,N_8721,N_8616);
xnor U8937 (N_8937,N_8780,N_8616);
or U8938 (N_8938,N_8638,N_8624);
nand U8939 (N_8939,N_8651,N_8735);
or U8940 (N_8940,N_8663,N_8764);
and U8941 (N_8941,N_8792,N_8737);
xnor U8942 (N_8942,N_8663,N_8631);
xor U8943 (N_8943,N_8785,N_8616);
xnor U8944 (N_8944,N_8674,N_8665);
nor U8945 (N_8945,N_8737,N_8649);
or U8946 (N_8946,N_8758,N_8731);
nand U8947 (N_8947,N_8767,N_8742);
and U8948 (N_8948,N_8792,N_8604);
and U8949 (N_8949,N_8768,N_8669);
and U8950 (N_8950,N_8727,N_8796);
and U8951 (N_8951,N_8673,N_8627);
and U8952 (N_8952,N_8717,N_8784);
and U8953 (N_8953,N_8625,N_8729);
nand U8954 (N_8954,N_8675,N_8714);
xor U8955 (N_8955,N_8605,N_8769);
or U8956 (N_8956,N_8628,N_8605);
nand U8957 (N_8957,N_8788,N_8641);
xor U8958 (N_8958,N_8665,N_8797);
nand U8959 (N_8959,N_8721,N_8726);
or U8960 (N_8960,N_8750,N_8662);
or U8961 (N_8961,N_8646,N_8601);
or U8962 (N_8962,N_8694,N_8762);
or U8963 (N_8963,N_8704,N_8737);
nand U8964 (N_8964,N_8630,N_8724);
nand U8965 (N_8965,N_8797,N_8715);
nor U8966 (N_8966,N_8702,N_8724);
and U8967 (N_8967,N_8683,N_8760);
or U8968 (N_8968,N_8601,N_8720);
nand U8969 (N_8969,N_8658,N_8751);
xor U8970 (N_8970,N_8635,N_8767);
xnor U8971 (N_8971,N_8620,N_8718);
nor U8972 (N_8972,N_8640,N_8796);
or U8973 (N_8973,N_8606,N_8711);
and U8974 (N_8974,N_8683,N_8798);
or U8975 (N_8975,N_8768,N_8739);
xnor U8976 (N_8976,N_8634,N_8727);
xnor U8977 (N_8977,N_8712,N_8756);
nand U8978 (N_8978,N_8694,N_8774);
and U8979 (N_8979,N_8661,N_8685);
nand U8980 (N_8980,N_8709,N_8734);
or U8981 (N_8981,N_8775,N_8657);
and U8982 (N_8982,N_8718,N_8698);
nand U8983 (N_8983,N_8681,N_8793);
xor U8984 (N_8984,N_8778,N_8742);
and U8985 (N_8985,N_8718,N_8740);
and U8986 (N_8986,N_8781,N_8699);
or U8987 (N_8987,N_8635,N_8786);
or U8988 (N_8988,N_8697,N_8724);
or U8989 (N_8989,N_8686,N_8762);
nor U8990 (N_8990,N_8760,N_8661);
and U8991 (N_8991,N_8632,N_8744);
and U8992 (N_8992,N_8600,N_8709);
and U8993 (N_8993,N_8603,N_8732);
xnor U8994 (N_8994,N_8621,N_8766);
nor U8995 (N_8995,N_8677,N_8767);
xor U8996 (N_8996,N_8632,N_8728);
nor U8997 (N_8997,N_8609,N_8781);
nor U8998 (N_8998,N_8709,N_8761);
xnor U8999 (N_8999,N_8629,N_8745);
nor U9000 (N_9000,N_8960,N_8803);
nand U9001 (N_9001,N_8897,N_8836);
and U9002 (N_9002,N_8819,N_8962);
xor U9003 (N_9003,N_8988,N_8990);
or U9004 (N_9004,N_8913,N_8868);
nand U9005 (N_9005,N_8809,N_8832);
xor U9006 (N_9006,N_8939,N_8923);
nor U9007 (N_9007,N_8851,N_8919);
xnor U9008 (N_9008,N_8804,N_8818);
or U9009 (N_9009,N_8958,N_8993);
and U9010 (N_9010,N_8860,N_8973);
xnor U9011 (N_9011,N_8944,N_8937);
xnor U9012 (N_9012,N_8918,N_8894);
nor U9013 (N_9013,N_8834,N_8921);
nand U9014 (N_9014,N_8811,N_8849);
xor U9015 (N_9015,N_8967,N_8887);
or U9016 (N_9016,N_8844,N_8873);
xor U9017 (N_9017,N_8892,N_8869);
or U9018 (N_9018,N_8911,N_8852);
nor U9019 (N_9019,N_8837,N_8974);
xor U9020 (N_9020,N_8883,N_8859);
xor U9021 (N_9021,N_8905,N_8979);
or U9022 (N_9022,N_8977,N_8885);
and U9023 (N_9023,N_8968,N_8840);
nor U9024 (N_9024,N_8874,N_8828);
nor U9025 (N_9025,N_8938,N_8929);
nor U9026 (N_9026,N_8877,N_8942);
and U9027 (N_9027,N_8880,N_8889);
nand U9028 (N_9028,N_8826,N_8855);
xor U9029 (N_9029,N_8972,N_8899);
and U9030 (N_9030,N_8940,N_8825);
nand U9031 (N_9031,N_8953,N_8916);
xor U9032 (N_9032,N_8932,N_8884);
xor U9033 (N_9033,N_8846,N_8903);
nand U9034 (N_9034,N_8985,N_8965);
nor U9035 (N_9035,N_8927,N_8945);
nor U9036 (N_9036,N_8980,N_8822);
nand U9037 (N_9037,N_8975,N_8935);
nor U9038 (N_9038,N_8956,N_8802);
or U9039 (N_9039,N_8807,N_8994);
xor U9040 (N_9040,N_8806,N_8912);
xnor U9041 (N_9041,N_8814,N_8835);
and U9042 (N_9042,N_8915,N_8984);
xor U9043 (N_9043,N_8928,N_8991);
and U9044 (N_9044,N_8854,N_8815);
nand U9045 (N_9045,N_8917,N_8845);
nand U9046 (N_9046,N_8961,N_8920);
and U9047 (N_9047,N_8982,N_8999);
xor U9048 (N_9048,N_8800,N_8963);
or U9049 (N_9049,N_8908,N_8995);
nand U9050 (N_9050,N_8954,N_8981);
nand U9051 (N_9051,N_8853,N_8941);
nand U9052 (N_9052,N_8895,N_8881);
and U9053 (N_9053,N_8898,N_8914);
nand U9054 (N_9054,N_8964,N_8878);
nand U9055 (N_9055,N_8816,N_8906);
or U9056 (N_9056,N_8924,N_8862);
nand U9057 (N_9057,N_8986,N_8870);
xnor U9058 (N_9058,N_8882,N_8998);
nor U9059 (N_9059,N_8931,N_8827);
xor U9060 (N_9060,N_8933,N_8902);
xor U9061 (N_9061,N_8901,N_8970);
and U9062 (N_9062,N_8830,N_8867);
or U9063 (N_9063,N_8904,N_8847);
xor U9064 (N_9064,N_8805,N_8808);
nand U9065 (N_9065,N_8821,N_8996);
nor U9066 (N_9066,N_8813,N_8978);
nor U9067 (N_9067,N_8983,N_8875);
nor U9068 (N_9068,N_8987,N_8841);
or U9069 (N_9069,N_8997,N_8872);
and U9070 (N_9070,N_8810,N_8969);
or U9071 (N_9071,N_8820,N_8896);
and U9072 (N_9072,N_8893,N_8949);
xnor U9073 (N_9073,N_8971,N_8891);
xor U9074 (N_9074,N_8839,N_8947);
nand U9075 (N_9075,N_8966,N_8930);
or U9076 (N_9076,N_8888,N_8812);
nor U9077 (N_9077,N_8886,N_8907);
and U9078 (N_9078,N_8879,N_8861);
xor U9079 (N_9079,N_8922,N_8831);
nor U9080 (N_9080,N_8952,N_8842);
and U9081 (N_9081,N_8823,N_8946);
or U9082 (N_9082,N_8838,N_8948);
nand U9083 (N_9083,N_8909,N_8890);
nor U9084 (N_9084,N_8865,N_8848);
nand U9085 (N_9085,N_8951,N_8833);
nor U9086 (N_9086,N_8925,N_8856);
nand U9087 (N_9087,N_8959,N_8936);
xor U9088 (N_9088,N_8801,N_8817);
or U9089 (N_9089,N_8866,N_8864);
and U9090 (N_9090,N_8900,N_8955);
or U9091 (N_9091,N_8934,N_8976);
and U9092 (N_9092,N_8950,N_8943);
and U9093 (N_9093,N_8926,N_8871);
nand U9094 (N_9094,N_8957,N_8829);
and U9095 (N_9095,N_8989,N_8843);
and U9096 (N_9096,N_8850,N_8863);
and U9097 (N_9097,N_8857,N_8824);
nand U9098 (N_9098,N_8992,N_8858);
and U9099 (N_9099,N_8876,N_8910);
xnor U9100 (N_9100,N_8872,N_8972);
or U9101 (N_9101,N_8993,N_8800);
nand U9102 (N_9102,N_8947,N_8995);
xor U9103 (N_9103,N_8878,N_8908);
and U9104 (N_9104,N_8931,N_8911);
or U9105 (N_9105,N_8981,N_8800);
xnor U9106 (N_9106,N_8855,N_8899);
nand U9107 (N_9107,N_8986,N_8984);
nor U9108 (N_9108,N_8977,N_8862);
nor U9109 (N_9109,N_8994,N_8915);
xnor U9110 (N_9110,N_8917,N_8940);
xor U9111 (N_9111,N_8947,N_8973);
nor U9112 (N_9112,N_8911,N_8995);
or U9113 (N_9113,N_8885,N_8919);
or U9114 (N_9114,N_8860,N_8940);
or U9115 (N_9115,N_8805,N_8887);
nor U9116 (N_9116,N_8928,N_8863);
nand U9117 (N_9117,N_8888,N_8977);
or U9118 (N_9118,N_8940,N_8981);
and U9119 (N_9119,N_8991,N_8909);
nand U9120 (N_9120,N_8917,N_8898);
or U9121 (N_9121,N_8870,N_8928);
nand U9122 (N_9122,N_8852,N_8957);
and U9123 (N_9123,N_8807,N_8982);
xnor U9124 (N_9124,N_8889,N_8803);
xnor U9125 (N_9125,N_8828,N_8903);
and U9126 (N_9126,N_8891,N_8979);
or U9127 (N_9127,N_8879,N_8865);
nand U9128 (N_9128,N_8922,N_8948);
nor U9129 (N_9129,N_8930,N_8965);
xnor U9130 (N_9130,N_8888,N_8933);
nand U9131 (N_9131,N_8819,N_8848);
nand U9132 (N_9132,N_8946,N_8817);
and U9133 (N_9133,N_8870,N_8968);
xnor U9134 (N_9134,N_8867,N_8902);
nor U9135 (N_9135,N_8937,N_8861);
nand U9136 (N_9136,N_8958,N_8833);
or U9137 (N_9137,N_8890,N_8844);
xnor U9138 (N_9138,N_8932,N_8923);
xnor U9139 (N_9139,N_8852,N_8912);
and U9140 (N_9140,N_8820,N_8929);
or U9141 (N_9141,N_8983,N_8939);
xnor U9142 (N_9142,N_8975,N_8840);
or U9143 (N_9143,N_8938,N_8845);
nand U9144 (N_9144,N_8936,N_8910);
and U9145 (N_9145,N_8960,N_8999);
and U9146 (N_9146,N_8802,N_8822);
and U9147 (N_9147,N_8885,N_8946);
nor U9148 (N_9148,N_8911,N_8982);
nor U9149 (N_9149,N_8997,N_8894);
nand U9150 (N_9150,N_8853,N_8820);
xor U9151 (N_9151,N_8851,N_8827);
xor U9152 (N_9152,N_8903,N_8923);
or U9153 (N_9153,N_8835,N_8863);
xor U9154 (N_9154,N_8898,N_8942);
or U9155 (N_9155,N_8819,N_8813);
and U9156 (N_9156,N_8958,N_8982);
or U9157 (N_9157,N_8918,N_8829);
nand U9158 (N_9158,N_8932,N_8994);
or U9159 (N_9159,N_8966,N_8998);
nand U9160 (N_9160,N_8936,N_8827);
nor U9161 (N_9161,N_8946,N_8883);
nand U9162 (N_9162,N_8929,N_8922);
nand U9163 (N_9163,N_8896,N_8997);
and U9164 (N_9164,N_8888,N_8985);
xnor U9165 (N_9165,N_8937,N_8934);
nand U9166 (N_9166,N_8923,N_8874);
nor U9167 (N_9167,N_8862,N_8839);
xnor U9168 (N_9168,N_8860,N_8848);
xor U9169 (N_9169,N_8843,N_8938);
and U9170 (N_9170,N_8866,N_8952);
xnor U9171 (N_9171,N_8997,N_8858);
or U9172 (N_9172,N_8982,N_8925);
nor U9173 (N_9173,N_8854,N_8857);
nand U9174 (N_9174,N_8982,N_8957);
or U9175 (N_9175,N_8882,N_8952);
or U9176 (N_9176,N_8917,N_8816);
nand U9177 (N_9177,N_8841,N_8953);
nand U9178 (N_9178,N_8901,N_8828);
nand U9179 (N_9179,N_8980,N_8816);
or U9180 (N_9180,N_8824,N_8817);
and U9181 (N_9181,N_8997,N_8891);
xnor U9182 (N_9182,N_8878,N_8942);
xor U9183 (N_9183,N_8828,N_8975);
or U9184 (N_9184,N_8888,N_8935);
xnor U9185 (N_9185,N_8878,N_8809);
and U9186 (N_9186,N_8870,N_8911);
and U9187 (N_9187,N_8993,N_8862);
nand U9188 (N_9188,N_8833,N_8856);
and U9189 (N_9189,N_8916,N_8993);
nand U9190 (N_9190,N_8956,N_8877);
nand U9191 (N_9191,N_8894,N_8868);
and U9192 (N_9192,N_8936,N_8905);
nor U9193 (N_9193,N_8830,N_8819);
nand U9194 (N_9194,N_8816,N_8961);
xor U9195 (N_9195,N_8997,N_8883);
nand U9196 (N_9196,N_8896,N_8878);
nor U9197 (N_9197,N_8821,N_8935);
nor U9198 (N_9198,N_8870,N_8879);
nand U9199 (N_9199,N_8901,N_8944);
nor U9200 (N_9200,N_9078,N_9185);
and U9201 (N_9201,N_9140,N_9148);
or U9202 (N_9202,N_9014,N_9178);
xnor U9203 (N_9203,N_9172,N_9083);
nand U9204 (N_9204,N_9117,N_9171);
nor U9205 (N_9205,N_9056,N_9141);
xnor U9206 (N_9206,N_9167,N_9190);
nor U9207 (N_9207,N_9123,N_9133);
nor U9208 (N_9208,N_9081,N_9037);
nand U9209 (N_9209,N_9130,N_9033);
and U9210 (N_9210,N_9165,N_9121);
or U9211 (N_9211,N_9054,N_9176);
xor U9212 (N_9212,N_9118,N_9115);
and U9213 (N_9213,N_9045,N_9158);
nor U9214 (N_9214,N_9076,N_9057);
or U9215 (N_9215,N_9052,N_9196);
or U9216 (N_9216,N_9146,N_9098);
nor U9217 (N_9217,N_9161,N_9046);
or U9218 (N_9218,N_9139,N_9072);
or U9219 (N_9219,N_9001,N_9025);
xor U9220 (N_9220,N_9067,N_9151);
or U9221 (N_9221,N_9020,N_9122);
nor U9222 (N_9222,N_9102,N_9147);
nand U9223 (N_9223,N_9024,N_9157);
or U9224 (N_9224,N_9095,N_9050);
or U9225 (N_9225,N_9179,N_9105);
xor U9226 (N_9226,N_9053,N_9000);
and U9227 (N_9227,N_9070,N_9004);
nor U9228 (N_9228,N_9128,N_9101);
nand U9229 (N_9229,N_9064,N_9086);
and U9230 (N_9230,N_9195,N_9082);
and U9231 (N_9231,N_9041,N_9085);
nor U9232 (N_9232,N_9173,N_9048);
nor U9233 (N_9233,N_9011,N_9012);
xnor U9234 (N_9234,N_9170,N_9097);
nand U9235 (N_9235,N_9155,N_9107);
nand U9236 (N_9236,N_9092,N_9022);
nor U9237 (N_9237,N_9091,N_9084);
nand U9238 (N_9238,N_9019,N_9152);
xnor U9239 (N_9239,N_9080,N_9144);
or U9240 (N_9240,N_9132,N_9188);
xor U9241 (N_9241,N_9166,N_9163);
or U9242 (N_9242,N_9087,N_9183);
nor U9243 (N_9243,N_9169,N_9194);
nor U9244 (N_9244,N_9007,N_9029);
or U9245 (N_9245,N_9073,N_9031);
nand U9246 (N_9246,N_9017,N_9009);
and U9247 (N_9247,N_9090,N_9096);
xor U9248 (N_9248,N_9186,N_9010);
or U9249 (N_9249,N_9189,N_9005);
and U9250 (N_9250,N_9187,N_9068);
nor U9251 (N_9251,N_9023,N_9034);
nand U9252 (N_9252,N_9079,N_9168);
nand U9253 (N_9253,N_9143,N_9109);
nor U9254 (N_9254,N_9175,N_9138);
nand U9255 (N_9255,N_9063,N_9066);
nor U9256 (N_9256,N_9013,N_9184);
xor U9257 (N_9257,N_9174,N_9153);
xor U9258 (N_9258,N_9162,N_9197);
nor U9259 (N_9259,N_9192,N_9016);
and U9260 (N_9260,N_9071,N_9111);
nor U9261 (N_9261,N_9039,N_9021);
xnor U9262 (N_9262,N_9129,N_9103);
nor U9263 (N_9263,N_9149,N_9112);
xor U9264 (N_9264,N_9089,N_9027);
or U9265 (N_9265,N_9059,N_9035);
xnor U9266 (N_9266,N_9088,N_9044);
nand U9267 (N_9267,N_9145,N_9049);
nor U9268 (N_9268,N_9093,N_9164);
nor U9269 (N_9269,N_9131,N_9002);
xnor U9270 (N_9270,N_9113,N_9150);
and U9271 (N_9271,N_9110,N_9154);
or U9272 (N_9272,N_9061,N_9120);
nand U9273 (N_9273,N_9119,N_9106);
nor U9274 (N_9274,N_9199,N_9126);
xnor U9275 (N_9275,N_9055,N_9036);
or U9276 (N_9276,N_9006,N_9077);
xor U9277 (N_9277,N_9127,N_9124);
nor U9278 (N_9278,N_9062,N_9058);
nand U9279 (N_9279,N_9018,N_9181);
or U9280 (N_9280,N_9040,N_9038);
and U9281 (N_9281,N_9042,N_9043);
or U9282 (N_9282,N_9125,N_9135);
or U9283 (N_9283,N_9193,N_9159);
xor U9284 (N_9284,N_9136,N_9047);
or U9285 (N_9285,N_9026,N_9069);
and U9286 (N_9286,N_9028,N_9142);
nor U9287 (N_9287,N_9060,N_9177);
xnor U9288 (N_9288,N_9094,N_9030);
xor U9289 (N_9289,N_9032,N_9065);
nor U9290 (N_9290,N_9104,N_9100);
xor U9291 (N_9291,N_9137,N_9015);
xnor U9292 (N_9292,N_9075,N_9191);
xor U9293 (N_9293,N_9074,N_9108);
nand U9294 (N_9294,N_9099,N_9180);
nor U9295 (N_9295,N_9160,N_9114);
xor U9296 (N_9296,N_9134,N_9051);
nor U9297 (N_9297,N_9182,N_9198);
nand U9298 (N_9298,N_9156,N_9116);
xnor U9299 (N_9299,N_9008,N_9003);
or U9300 (N_9300,N_9153,N_9059);
xor U9301 (N_9301,N_9121,N_9195);
nand U9302 (N_9302,N_9074,N_9101);
nor U9303 (N_9303,N_9148,N_9001);
xnor U9304 (N_9304,N_9058,N_9063);
and U9305 (N_9305,N_9072,N_9167);
nor U9306 (N_9306,N_9040,N_9195);
nor U9307 (N_9307,N_9094,N_9041);
and U9308 (N_9308,N_9096,N_9061);
nor U9309 (N_9309,N_9058,N_9191);
xor U9310 (N_9310,N_9051,N_9025);
and U9311 (N_9311,N_9148,N_9126);
nand U9312 (N_9312,N_9116,N_9123);
and U9313 (N_9313,N_9027,N_9047);
xor U9314 (N_9314,N_9122,N_9161);
or U9315 (N_9315,N_9118,N_9019);
nor U9316 (N_9316,N_9194,N_9093);
nor U9317 (N_9317,N_9015,N_9152);
or U9318 (N_9318,N_9018,N_9025);
or U9319 (N_9319,N_9081,N_9135);
or U9320 (N_9320,N_9053,N_9199);
and U9321 (N_9321,N_9032,N_9183);
and U9322 (N_9322,N_9071,N_9187);
xor U9323 (N_9323,N_9135,N_9150);
or U9324 (N_9324,N_9048,N_9028);
or U9325 (N_9325,N_9056,N_9189);
nand U9326 (N_9326,N_9056,N_9057);
and U9327 (N_9327,N_9111,N_9147);
or U9328 (N_9328,N_9196,N_9017);
xnor U9329 (N_9329,N_9045,N_9038);
nor U9330 (N_9330,N_9035,N_9050);
nand U9331 (N_9331,N_9092,N_9021);
nor U9332 (N_9332,N_9165,N_9174);
and U9333 (N_9333,N_9081,N_9108);
xnor U9334 (N_9334,N_9145,N_9142);
and U9335 (N_9335,N_9155,N_9128);
nor U9336 (N_9336,N_9161,N_9131);
nand U9337 (N_9337,N_9142,N_9035);
or U9338 (N_9338,N_9175,N_9160);
xor U9339 (N_9339,N_9164,N_9166);
xnor U9340 (N_9340,N_9165,N_9065);
nor U9341 (N_9341,N_9121,N_9189);
xnor U9342 (N_9342,N_9162,N_9111);
xor U9343 (N_9343,N_9032,N_9121);
and U9344 (N_9344,N_9023,N_9157);
nor U9345 (N_9345,N_9158,N_9166);
and U9346 (N_9346,N_9091,N_9183);
or U9347 (N_9347,N_9074,N_9105);
nand U9348 (N_9348,N_9110,N_9119);
and U9349 (N_9349,N_9056,N_9055);
nor U9350 (N_9350,N_9026,N_9179);
nand U9351 (N_9351,N_9070,N_9194);
or U9352 (N_9352,N_9176,N_9195);
and U9353 (N_9353,N_9071,N_9195);
nor U9354 (N_9354,N_9111,N_9193);
nor U9355 (N_9355,N_9142,N_9011);
nand U9356 (N_9356,N_9160,N_9123);
and U9357 (N_9357,N_9106,N_9032);
or U9358 (N_9358,N_9179,N_9169);
nand U9359 (N_9359,N_9081,N_9054);
nor U9360 (N_9360,N_9095,N_9032);
and U9361 (N_9361,N_9179,N_9176);
or U9362 (N_9362,N_9124,N_9074);
xor U9363 (N_9363,N_9144,N_9115);
nor U9364 (N_9364,N_9041,N_9017);
and U9365 (N_9365,N_9064,N_9190);
or U9366 (N_9366,N_9102,N_9151);
or U9367 (N_9367,N_9118,N_9028);
xor U9368 (N_9368,N_9138,N_9038);
or U9369 (N_9369,N_9182,N_9014);
or U9370 (N_9370,N_9130,N_9144);
or U9371 (N_9371,N_9102,N_9153);
nor U9372 (N_9372,N_9151,N_9063);
xor U9373 (N_9373,N_9162,N_9076);
xnor U9374 (N_9374,N_9137,N_9037);
xor U9375 (N_9375,N_9129,N_9083);
nand U9376 (N_9376,N_9182,N_9199);
nand U9377 (N_9377,N_9112,N_9096);
nor U9378 (N_9378,N_9021,N_9078);
nand U9379 (N_9379,N_9106,N_9153);
xnor U9380 (N_9380,N_9147,N_9073);
and U9381 (N_9381,N_9135,N_9058);
nor U9382 (N_9382,N_9112,N_9141);
nor U9383 (N_9383,N_9124,N_9031);
nor U9384 (N_9384,N_9121,N_9031);
and U9385 (N_9385,N_9034,N_9111);
and U9386 (N_9386,N_9146,N_9002);
or U9387 (N_9387,N_9078,N_9151);
nor U9388 (N_9388,N_9062,N_9010);
nor U9389 (N_9389,N_9094,N_9034);
and U9390 (N_9390,N_9186,N_9197);
nor U9391 (N_9391,N_9117,N_9039);
xnor U9392 (N_9392,N_9037,N_9196);
or U9393 (N_9393,N_9131,N_9087);
and U9394 (N_9394,N_9043,N_9031);
and U9395 (N_9395,N_9151,N_9161);
or U9396 (N_9396,N_9165,N_9074);
nor U9397 (N_9397,N_9031,N_9094);
nand U9398 (N_9398,N_9085,N_9179);
nand U9399 (N_9399,N_9030,N_9137);
xor U9400 (N_9400,N_9321,N_9225);
xnor U9401 (N_9401,N_9351,N_9391);
xor U9402 (N_9402,N_9201,N_9278);
and U9403 (N_9403,N_9326,N_9397);
and U9404 (N_9404,N_9264,N_9339);
xnor U9405 (N_9405,N_9297,N_9323);
xnor U9406 (N_9406,N_9301,N_9227);
xor U9407 (N_9407,N_9276,N_9367);
and U9408 (N_9408,N_9237,N_9224);
nor U9409 (N_9409,N_9382,N_9275);
nand U9410 (N_9410,N_9340,N_9258);
and U9411 (N_9411,N_9289,N_9385);
or U9412 (N_9412,N_9314,N_9252);
nor U9413 (N_9413,N_9318,N_9373);
nor U9414 (N_9414,N_9344,N_9399);
xor U9415 (N_9415,N_9349,N_9380);
xnor U9416 (N_9416,N_9304,N_9346);
xnor U9417 (N_9417,N_9204,N_9300);
and U9418 (N_9418,N_9287,N_9356);
and U9419 (N_9419,N_9241,N_9214);
xor U9420 (N_9420,N_9315,N_9228);
xnor U9421 (N_9421,N_9374,N_9248);
nand U9422 (N_9422,N_9381,N_9302);
nor U9423 (N_9423,N_9250,N_9312);
nand U9424 (N_9424,N_9215,N_9370);
or U9425 (N_9425,N_9386,N_9325);
nor U9426 (N_9426,N_9369,N_9223);
and U9427 (N_9427,N_9293,N_9209);
xnor U9428 (N_9428,N_9234,N_9230);
nor U9429 (N_9429,N_9366,N_9333);
nor U9430 (N_9430,N_9308,N_9210);
xnor U9431 (N_9431,N_9244,N_9328);
xor U9432 (N_9432,N_9341,N_9238);
and U9433 (N_9433,N_9233,N_9305);
nor U9434 (N_9434,N_9246,N_9329);
or U9435 (N_9435,N_9389,N_9249);
nand U9436 (N_9436,N_9239,N_9274);
or U9437 (N_9437,N_9263,N_9288);
or U9438 (N_9438,N_9286,N_9332);
and U9439 (N_9439,N_9379,N_9217);
or U9440 (N_9440,N_9272,N_9383);
xor U9441 (N_9441,N_9222,N_9306);
nor U9442 (N_9442,N_9296,N_9218);
xor U9443 (N_9443,N_9271,N_9336);
nor U9444 (N_9444,N_9299,N_9242);
nor U9445 (N_9445,N_9394,N_9396);
nor U9446 (N_9446,N_9206,N_9282);
nor U9447 (N_9447,N_9377,N_9232);
nor U9448 (N_9448,N_9364,N_9350);
nand U9449 (N_9449,N_9281,N_9322);
xnor U9450 (N_9450,N_9208,N_9283);
nand U9451 (N_9451,N_9365,N_9345);
xor U9452 (N_9452,N_9387,N_9295);
nand U9453 (N_9453,N_9330,N_9393);
xnor U9454 (N_9454,N_9335,N_9231);
or U9455 (N_9455,N_9235,N_9324);
nor U9456 (N_9456,N_9265,N_9347);
and U9457 (N_9457,N_9202,N_9376);
nand U9458 (N_9458,N_9392,N_9372);
xnor U9459 (N_9459,N_9310,N_9256);
xor U9460 (N_9460,N_9290,N_9213);
or U9461 (N_9461,N_9334,N_9285);
nor U9462 (N_9462,N_9360,N_9257);
xnor U9463 (N_9463,N_9337,N_9268);
or U9464 (N_9464,N_9327,N_9200);
and U9465 (N_9465,N_9362,N_9375);
nand U9466 (N_9466,N_9319,N_9226);
xnor U9467 (N_9467,N_9211,N_9259);
nor U9468 (N_9468,N_9371,N_9352);
nand U9469 (N_9469,N_9358,N_9357);
nand U9470 (N_9470,N_9205,N_9273);
xnor U9471 (N_9471,N_9251,N_9359);
and U9472 (N_9472,N_9221,N_9216);
nor U9473 (N_9473,N_9388,N_9390);
nor U9474 (N_9474,N_9353,N_9331);
nand U9475 (N_9475,N_9361,N_9292);
nand U9476 (N_9476,N_9279,N_9236);
nand U9477 (N_9477,N_9270,N_9354);
xnor U9478 (N_9478,N_9253,N_9291);
nor U9479 (N_9479,N_9395,N_9245);
nand U9480 (N_9480,N_9255,N_9378);
nor U9481 (N_9481,N_9203,N_9317);
and U9482 (N_9482,N_9267,N_9316);
or U9483 (N_9483,N_9384,N_9280);
and U9484 (N_9484,N_9284,N_9368);
and U9485 (N_9485,N_9277,N_9260);
xor U9486 (N_9486,N_9220,N_9269);
and U9487 (N_9487,N_9229,N_9240);
and U9488 (N_9488,N_9298,N_9320);
nand U9489 (N_9489,N_9348,N_9262);
and U9490 (N_9490,N_9247,N_9303);
nor U9491 (N_9491,N_9313,N_9266);
nor U9492 (N_9492,N_9207,N_9355);
or U9493 (N_9493,N_9294,N_9311);
nor U9494 (N_9494,N_9342,N_9212);
and U9495 (N_9495,N_9307,N_9254);
nand U9496 (N_9496,N_9338,N_9243);
and U9497 (N_9497,N_9398,N_9309);
or U9498 (N_9498,N_9261,N_9363);
nand U9499 (N_9499,N_9343,N_9219);
and U9500 (N_9500,N_9289,N_9302);
nand U9501 (N_9501,N_9267,N_9333);
or U9502 (N_9502,N_9205,N_9381);
and U9503 (N_9503,N_9263,N_9328);
nand U9504 (N_9504,N_9231,N_9275);
or U9505 (N_9505,N_9236,N_9380);
or U9506 (N_9506,N_9259,N_9352);
and U9507 (N_9507,N_9340,N_9273);
and U9508 (N_9508,N_9257,N_9319);
nor U9509 (N_9509,N_9254,N_9341);
xor U9510 (N_9510,N_9340,N_9375);
and U9511 (N_9511,N_9249,N_9369);
xor U9512 (N_9512,N_9212,N_9375);
nand U9513 (N_9513,N_9319,N_9292);
or U9514 (N_9514,N_9365,N_9251);
and U9515 (N_9515,N_9266,N_9342);
nor U9516 (N_9516,N_9285,N_9265);
xnor U9517 (N_9517,N_9386,N_9234);
nand U9518 (N_9518,N_9302,N_9252);
or U9519 (N_9519,N_9255,N_9282);
xor U9520 (N_9520,N_9268,N_9284);
nor U9521 (N_9521,N_9378,N_9206);
or U9522 (N_9522,N_9300,N_9209);
nand U9523 (N_9523,N_9316,N_9307);
nand U9524 (N_9524,N_9293,N_9306);
nand U9525 (N_9525,N_9357,N_9373);
nand U9526 (N_9526,N_9372,N_9249);
and U9527 (N_9527,N_9304,N_9343);
xnor U9528 (N_9528,N_9372,N_9333);
and U9529 (N_9529,N_9220,N_9336);
nor U9530 (N_9530,N_9380,N_9219);
and U9531 (N_9531,N_9337,N_9368);
and U9532 (N_9532,N_9307,N_9298);
and U9533 (N_9533,N_9284,N_9316);
xor U9534 (N_9534,N_9220,N_9300);
and U9535 (N_9535,N_9369,N_9240);
or U9536 (N_9536,N_9354,N_9332);
xnor U9537 (N_9537,N_9298,N_9289);
nand U9538 (N_9538,N_9315,N_9380);
or U9539 (N_9539,N_9249,N_9323);
or U9540 (N_9540,N_9391,N_9239);
and U9541 (N_9541,N_9201,N_9386);
xnor U9542 (N_9542,N_9313,N_9288);
or U9543 (N_9543,N_9397,N_9227);
or U9544 (N_9544,N_9320,N_9205);
xor U9545 (N_9545,N_9293,N_9214);
or U9546 (N_9546,N_9377,N_9240);
nand U9547 (N_9547,N_9224,N_9338);
or U9548 (N_9548,N_9204,N_9371);
and U9549 (N_9549,N_9347,N_9252);
nand U9550 (N_9550,N_9368,N_9356);
xor U9551 (N_9551,N_9363,N_9298);
and U9552 (N_9552,N_9283,N_9297);
nand U9553 (N_9553,N_9259,N_9269);
or U9554 (N_9554,N_9201,N_9268);
or U9555 (N_9555,N_9216,N_9382);
or U9556 (N_9556,N_9307,N_9207);
xnor U9557 (N_9557,N_9284,N_9390);
or U9558 (N_9558,N_9223,N_9316);
and U9559 (N_9559,N_9379,N_9235);
xor U9560 (N_9560,N_9294,N_9328);
xor U9561 (N_9561,N_9325,N_9345);
or U9562 (N_9562,N_9374,N_9386);
nor U9563 (N_9563,N_9204,N_9233);
and U9564 (N_9564,N_9353,N_9216);
xnor U9565 (N_9565,N_9280,N_9363);
nor U9566 (N_9566,N_9275,N_9219);
nor U9567 (N_9567,N_9319,N_9242);
and U9568 (N_9568,N_9348,N_9253);
nand U9569 (N_9569,N_9396,N_9318);
and U9570 (N_9570,N_9269,N_9287);
or U9571 (N_9571,N_9254,N_9257);
nor U9572 (N_9572,N_9202,N_9227);
nor U9573 (N_9573,N_9226,N_9386);
or U9574 (N_9574,N_9283,N_9292);
and U9575 (N_9575,N_9341,N_9309);
nor U9576 (N_9576,N_9335,N_9376);
nand U9577 (N_9577,N_9342,N_9286);
xor U9578 (N_9578,N_9372,N_9297);
xor U9579 (N_9579,N_9338,N_9385);
nand U9580 (N_9580,N_9275,N_9354);
and U9581 (N_9581,N_9370,N_9277);
or U9582 (N_9582,N_9374,N_9229);
nand U9583 (N_9583,N_9383,N_9220);
nor U9584 (N_9584,N_9303,N_9360);
xnor U9585 (N_9585,N_9279,N_9207);
xor U9586 (N_9586,N_9242,N_9351);
xnor U9587 (N_9587,N_9205,N_9252);
nand U9588 (N_9588,N_9281,N_9235);
nor U9589 (N_9589,N_9250,N_9399);
xor U9590 (N_9590,N_9354,N_9262);
and U9591 (N_9591,N_9210,N_9280);
and U9592 (N_9592,N_9286,N_9359);
or U9593 (N_9593,N_9305,N_9335);
xor U9594 (N_9594,N_9389,N_9384);
xor U9595 (N_9595,N_9359,N_9249);
xnor U9596 (N_9596,N_9213,N_9234);
xor U9597 (N_9597,N_9310,N_9387);
nor U9598 (N_9598,N_9398,N_9313);
nor U9599 (N_9599,N_9228,N_9322);
or U9600 (N_9600,N_9598,N_9448);
xnor U9601 (N_9601,N_9470,N_9531);
nand U9602 (N_9602,N_9479,N_9558);
nor U9603 (N_9603,N_9570,N_9447);
xnor U9604 (N_9604,N_9476,N_9541);
nand U9605 (N_9605,N_9537,N_9547);
nand U9606 (N_9606,N_9439,N_9596);
nor U9607 (N_9607,N_9462,N_9485);
nand U9608 (N_9608,N_9508,N_9403);
nand U9609 (N_9609,N_9597,N_9407);
and U9610 (N_9610,N_9560,N_9525);
nand U9611 (N_9611,N_9506,N_9577);
xor U9612 (N_9612,N_9555,N_9416);
and U9613 (N_9613,N_9538,N_9520);
or U9614 (N_9614,N_9496,N_9551);
nand U9615 (N_9615,N_9575,N_9469);
or U9616 (N_9616,N_9491,N_9453);
nand U9617 (N_9617,N_9440,N_9595);
nor U9618 (N_9618,N_9410,N_9486);
and U9619 (N_9619,N_9489,N_9433);
or U9620 (N_9620,N_9550,N_9473);
nor U9621 (N_9621,N_9456,N_9542);
nand U9622 (N_9622,N_9580,N_9414);
nor U9623 (N_9623,N_9475,N_9499);
xnor U9624 (N_9624,N_9468,N_9408);
nand U9625 (N_9625,N_9425,N_9492);
nor U9626 (N_9626,N_9521,N_9402);
and U9627 (N_9627,N_9458,N_9553);
nand U9628 (N_9628,N_9552,N_9498);
or U9629 (N_9629,N_9406,N_9514);
or U9630 (N_9630,N_9454,N_9568);
and U9631 (N_9631,N_9554,N_9515);
and U9632 (N_9632,N_9400,N_9412);
xor U9633 (N_9633,N_9588,N_9532);
nand U9634 (N_9634,N_9452,N_9589);
xor U9635 (N_9635,N_9430,N_9565);
xor U9636 (N_9636,N_9463,N_9451);
or U9637 (N_9637,N_9441,N_9585);
xor U9638 (N_9638,N_9438,N_9420);
xor U9639 (N_9639,N_9587,N_9459);
or U9640 (N_9640,N_9417,N_9513);
xnor U9641 (N_9641,N_9471,N_9450);
or U9642 (N_9642,N_9401,N_9534);
nand U9643 (N_9643,N_9460,N_9444);
nor U9644 (N_9644,N_9427,N_9405);
nand U9645 (N_9645,N_9599,N_9527);
nand U9646 (N_9646,N_9591,N_9546);
or U9647 (N_9647,N_9467,N_9556);
or U9648 (N_9648,N_9474,N_9523);
xnor U9649 (N_9649,N_9481,N_9422);
or U9650 (N_9650,N_9497,N_9442);
xnor U9651 (N_9651,N_9483,N_9533);
and U9652 (N_9652,N_9509,N_9435);
or U9653 (N_9653,N_9413,N_9567);
nand U9654 (N_9654,N_9432,N_9529);
nand U9655 (N_9655,N_9582,N_9411);
nand U9656 (N_9656,N_9562,N_9445);
and U9657 (N_9657,N_9522,N_9524);
and U9658 (N_9658,N_9477,N_9484);
nand U9659 (N_9659,N_9429,N_9507);
and U9660 (N_9660,N_9518,N_9569);
xnor U9661 (N_9661,N_9465,N_9593);
or U9662 (N_9662,N_9519,N_9549);
nor U9663 (N_9663,N_9528,N_9584);
or U9664 (N_9664,N_9443,N_9446);
nand U9665 (N_9665,N_9510,N_9455);
and U9666 (N_9666,N_9505,N_9466);
nor U9667 (N_9667,N_9536,N_9428);
xnor U9668 (N_9668,N_9590,N_9423);
or U9669 (N_9669,N_9581,N_9490);
and U9670 (N_9670,N_9418,N_9557);
nand U9671 (N_9671,N_9431,N_9512);
or U9672 (N_9672,N_9434,N_9500);
xnor U9673 (N_9673,N_9503,N_9576);
and U9674 (N_9674,N_9566,N_9504);
xnor U9675 (N_9675,N_9586,N_9404);
nand U9676 (N_9676,N_9457,N_9495);
and U9677 (N_9677,N_9561,N_9493);
or U9678 (N_9678,N_9502,N_9594);
nor U9679 (N_9679,N_9517,N_9461);
or U9680 (N_9680,N_9449,N_9535);
and U9681 (N_9681,N_9437,N_9526);
nand U9682 (N_9682,N_9488,N_9501);
xnor U9683 (N_9683,N_9572,N_9564);
xnor U9684 (N_9684,N_9421,N_9415);
nand U9685 (N_9685,N_9487,N_9579);
xor U9686 (N_9686,N_9559,N_9592);
and U9687 (N_9687,N_9530,N_9573);
xnor U9688 (N_9688,N_9478,N_9419);
xnor U9689 (N_9689,N_9516,N_9539);
xnor U9690 (N_9690,N_9544,N_9583);
nor U9691 (N_9691,N_9578,N_9464);
nor U9692 (N_9692,N_9540,N_9574);
nor U9693 (N_9693,N_9426,N_9571);
or U9694 (N_9694,N_9511,N_9545);
nor U9695 (N_9695,N_9494,N_9436);
nand U9696 (N_9696,N_9409,N_9480);
and U9697 (N_9697,N_9472,N_9543);
nor U9698 (N_9698,N_9548,N_9424);
xor U9699 (N_9699,N_9563,N_9482);
xor U9700 (N_9700,N_9541,N_9449);
or U9701 (N_9701,N_9411,N_9595);
nand U9702 (N_9702,N_9523,N_9537);
nand U9703 (N_9703,N_9563,N_9442);
or U9704 (N_9704,N_9597,N_9562);
and U9705 (N_9705,N_9583,N_9436);
or U9706 (N_9706,N_9423,N_9509);
or U9707 (N_9707,N_9418,N_9591);
xor U9708 (N_9708,N_9534,N_9495);
and U9709 (N_9709,N_9468,N_9498);
nor U9710 (N_9710,N_9461,N_9579);
or U9711 (N_9711,N_9415,N_9401);
nor U9712 (N_9712,N_9597,N_9576);
or U9713 (N_9713,N_9570,N_9407);
and U9714 (N_9714,N_9587,N_9556);
xor U9715 (N_9715,N_9472,N_9506);
xnor U9716 (N_9716,N_9498,N_9500);
xnor U9717 (N_9717,N_9405,N_9423);
and U9718 (N_9718,N_9453,N_9484);
nand U9719 (N_9719,N_9494,N_9591);
or U9720 (N_9720,N_9483,N_9456);
nand U9721 (N_9721,N_9428,N_9578);
and U9722 (N_9722,N_9499,N_9436);
or U9723 (N_9723,N_9562,N_9580);
nor U9724 (N_9724,N_9408,N_9409);
nand U9725 (N_9725,N_9578,N_9541);
nor U9726 (N_9726,N_9420,N_9555);
nand U9727 (N_9727,N_9595,N_9555);
or U9728 (N_9728,N_9518,N_9436);
nand U9729 (N_9729,N_9464,N_9416);
and U9730 (N_9730,N_9485,N_9465);
nand U9731 (N_9731,N_9467,N_9403);
and U9732 (N_9732,N_9548,N_9538);
nor U9733 (N_9733,N_9544,N_9424);
xnor U9734 (N_9734,N_9447,N_9468);
xor U9735 (N_9735,N_9550,N_9432);
nor U9736 (N_9736,N_9543,N_9410);
nand U9737 (N_9737,N_9440,N_9598);
nand U9738 (N_9738,N_9411,N_9523);
and U9739 (N_9739,N_9462,N_9464);
nor U9740 (N_9740,N_9545,N_9474);
xnor U9741 (N_9741,N_9561,N_9485);
xor U9742 (N_9742,N_9410,N_9565);
and U9743 (N_9743,N_9405,N_9562);
nand U9744 (N_9744,N_9589,N_9414);
xor U9745 (N_9745,N_9580,N_9556);
or U9746 (N_9746,N_9495,N_9478);
or U9747 (N_9747,N_9421,N_9529);
nand U9748 (N_9748,N_9479,N_9567);
xor U9749 (N_9749,N_9527,N_9549);
nor U9750 (N_9750,N_9439,N_9532);
nand U9751 (N_9751,N_9582,N_9432);
and U9752 (N_9752,N_9520,N_9535);
and U9753 (N_9753,N_9449,N_9467);
nor U9754 (N_9754,N_9432,N_9431);
xnor U9755 (N_9755,N_9423,N_9548);
or U9756 (N_9756,N_9519,N_9575);
or U9757 (N_9757,N_9484,N_9536);
xor U9758 (N_9758,N_9516,N_9435);
or U9759 (N_9759,N_9569,N_9442);
and U9760 (N_9760,N_9426,N_9565);
and U9761 (N_9761,N_9537,N_9488);
nand U9762 (N_9762,N_9530,N_9500);
or U9763 (N_9763,N_9592,N_9423);
nand U9764 (N_9764,N_9468,N_9512);
nor U9765 (N_9765,N_9434,N_9439);
xnor U9766 (N_9766,N_9443,N_9499);
or U9767 (N_9767,N_9594,N_9441);
and U9768 (N_9768,N_9497,N_9440);
and U9769 (N_9769,N_9560,N_9469);
and U9770 (N_9770,N_9484,N_9544);
and U9771 (N_9771,N_9575,N_9489);
and U9772 (N_9772,N_9458,N_9569);
and U9773 (N_9773,N_9571,N_9557);
and U9774 (N_9774,N_9461,N_9571);
nor U9775 (N_9775,N_9461,N_9477);
nor U9776 (N_9776,N_9423,N_9407);
nand U9777 (N_9777,N_9576,N_9510);
nand U9778 (N_9778,N_9493,N_9414);
nand U9779 (N_9779,N_9499,N_9482);
nand U9780 (N_9780,N_9475,N_9567);
nor U9781 (N_9781,N_9500,N_9433);
or U9782 (N_9782,N_9436,N_9541);
and U9783 (N_9783,N_9491,N_9454);
nand U9784 (N_9784,N_9546,N_9468);
xnor U9785 (N_9785,N_9406,N_9574);
and U9786 (N_9786,N_9546,N_9438);
and U9787 (N_9787,N_9471,N_9440);
and U9788 (N_9788,N_9498,N_9535);
nand U9789 (N_9789,N_9541,N_9464);
and U9790 (N_9790,N_9599,N_9483);
nor U9791 (N_9791,N_9527,N_9486);
xnor U9792 (N_9792,N_9507,N_9569);
or U9793 (N_9793,N_9540,N_9521);
or U9794 (N_9794,N_9482,N_9414);
nor U9795 (N_9795,N_9456,N_9539);
or U9796 (N_9796,N_9578,N_9560);
xnor U9797 (N_9797,N_9421,N_9560);
xor U9798 (N_9798,N_9576,N_9582);
and U9799 (N_9799,N_9579,N_9486);
nor U9800 (N_9800,N_9621,N_9600);
xnor U9801 (N_9801,N_9775,N_9772);
xnor U9802 (N_9802,N_9611,N_9661);
xor U9803 (N_9803,N_9690,N_9734);
nand U9804 (N_9804,N_9787,N_9613);
xor U9805 (N_9805,N_9644,N_9773);
nor U9806 (N_9806,N_9752,N_9761);
nand U9807 (N_9807,N_9608,N_9601);
nand U9808 (N_9808,N_9618,N_9706);
or U9809 (N_9809,N_9643,N_9749);
nand U9810 (N_9810,N_9650,N_9623);
or U9811 (N_9811,N_9676,N_9604);
and U9812 (N_9812,N_9732,N_9740);
or U9813 (N_9813,N_9794,N_9738);
and U9814 (N_9814,N_9607,N_9663);
or U9815 (N_9815,N_9662,N_9768);
or U9816 (N_9816,N_9779,N_9656);
nor U9817 (N_9817,N_9748,N_9707);
nor U9818 (N_9818,N_9624,N_9796);
and U9819 (N_9819,N_9709,N_9784);
and U9820 (N_9820,N_9646,N_9717);
and U9821 (N_9821,N_9710,N_9770);
xnor U9822 (N_9822,N_9625,N_9627);
nor U9823 (N_9823,N_9700,N_9631);
and U9824 (N_9824,N_9799,N_9686);
or U9825 (N_9825,N_9635,N_9792);
nand U9826 (N_9826,N_9671,N_9777);
and U9827 (N_9827,N_9798,N_9719);
nand U9828 (N_9828,N_9679,N_9688);
or U9829 (N_9829,N_9733,N_9687);
or U9830 (N_9830,N_9652,N_9703);
nand U9831 (N_9831,N_9664,N_9648);
xnor U9832 (N_9832,N_9704,N_9786);
xnor U9833 (N_9833,N_9746,N_9774);
nand U9834 (N_9834,N_9753,N_9637);
xor U9835 (N_9835,N_9744,N_9682);
and U9836 (N_9836,N_9767,N_9667);
nor U9837 (N_9837,N_9653,N_9657);
xor U9838 (N_9838,N_9639,N_9736);
nand U9839 (N_9839,N_9712,N_9751);
nor U9840 (N_9840,N_9730,N_9741);
xor U9841 (N_9841,N_9689,N_9756);
and U9842 (N_9842,N_9747,N_9699);
xor U9843 (N_9843,N_9750,N_9714);
and U9844 (N_9844,N_9785,N_9616);
or U9845 (N_9845,N_9691,N_9735);
xnor U9846 (N_9846,N_9790,N_9640);
nor U9847 (N_9847,N_9698,N_9665);
nand U9848 (N_9848,N_9680,N_9612);
and U9849 (N_9849,N_9673,N_9658);
or U9850 (N_9850,N_9739,N_9702);
nor U9851 (N_9851,N_9781,N_9636);
and U9852 (N_9852,N_9668,N_9649);
or U9853 (N_9853,N_9797,N_9620);
xnor U9854 (N_9854,N_9666,N_9684);
or U9855 (N_9855,N_9766,N_9602);
or U9856 (N_9856,N_9633,N_9615);
or U9857 (N_9857,N_9638,N_9692);
or U9858 (N_9858,N_9672,N_9745);
xnor U9859 (N_9859,N_9695,N_9760);
nand U9860 (N_9860,N_9782,N_9642);
nand U9861 (N_9861,N_9681,N_9697);
nand U9862 (N_9862,N_9743,N_9725);
xor U9863 (N_9863,N_9634,N_9763);
nand U9864 (N_9864,N_9713,N_9609);
nor U9865 (N_9865,N_9742,N_9795);
or U9866 (N_9866,N_9641,N_9708);
and U9867 (N_9867,N_9783,N_9614);
xnor U9868 (N_9868,N_9701,N_9685);
and U9869 (N_9869,N_9670,N_9678);
xnor U9870 (N_9870,N_9677,N_9720);
xor U9871 (N_9871,N_9654,N_9651);
xnor U9872 (N_9872,N_9716,N_9721);
xor U9873 (N_9873,N_9696,N_9778);
xor U9874 (N_9874,N_9737,N_9674);
or U9875 (N_9875,N_9726,N_9765);
or U9876 (N_9876,N_9758,N_9769);
xor U9877 (N_9877,N_9655,N_9718);
or U9878 (N_9878,N_9729,N_9727);
xnor U9879 (N_9879,N_9728,N_9776);
or U9880 (N_9880,N_9722,N_9619);
or U9881 (N_9881,N_9780,N_9610);
nor U9882 (N_9882,N_9762,N_9793);
or U9883 (N_9883,N_9683,N_9757);
and U9884 (N_9884,N_9723,N_9705);
nor U9885 (N_9885,N_9731,N_9754);
xnor U9886 (N_9886,N_9606,N_9755);
xor U9887 (N_9887,N_9693,N_9724);
and U9888 (N_9888,N_9647,N_9632);
nand U9889 (N_9889,N_9605,N_9788);
and U9890 (N_9890,N_9629,N_9759);
and U9891 (N_9891,N_9630,N_9669);
nand U9892 (N_9892,N_9764,N_9791);
xor U9893 (N_9893,N_9789,N_9675);
nand U9894 (N_9894,N_9628,N_9622);
and U9895 (N_9895,N_9694,N_9659);
and U9896 (N_9896,N_9626,N_9715);
or U9897 (N_9897,N_9771,N_9603);
xnor U9898 (N_9898,N_9660,N_9711);
or U9899 (N_9899,N_9645,N_9617);
and U9900 (N_9900,N_9664,N_9631);
and U9901 (N_9901,N_9622,N_9644);
nand U9902 (N_9902,N_9788,N_9612);
and U9903 (N_9903,N_9673,N_9692);
and U9904 (N_9904,N_9784,N_9699);
nand U9905 (N_9905,N_9678,N_9754);
nand U9906 (N_9906,N_9786,N_9610);
or U9907 (N_9907,N_9669,N_9790);
xor U9908 (N_9908,N_9731,N_9705);
xor U9909 (N_9909,N_9766,N_9626);
and U9910 (N_9910,N_9745,N_9678);
nand U9911 (N_9911,N_9660,N_9785);
xor U9912 (N_9912,N_9683,N_9685);
and U9913 (N_9913,N_9647,N_9762);
and U9914 (N_9914,N_9646,N_9766);
and U9915 (N_9915,N_9725,N_9600);
xnor U9916 (N_9916,N_9792,N_9781);
xnor U9917 (N_9917,N_9708,N_9738);
nor U9918 (N_9918,N_9631,N_9640);
or U9919 (N_9919,N_9626,N_9734);
nor U9920 (N_9920,N_9634,N_9781);
xnor U9921 (N_9921,N_9736,N_9650);
nand U9922 (N_9922,N_9743,N_9768);
nand U9923 (N_9923,N_9714,N_9657);
or U9924 (N_9924,N_9667,N_9641);
and U9925 (N_9925,N_9698,N_9664);
or U9926 (N_9926,N_9676,N_9790);
or U9927 (N_9927,N_9744,N_9770);
xor U9928 (N_9928,N_9760,N_9631);
nand U9929 (N_9929,N_9669,N_9734);
nor U9930 (N_9930,N_9629,N_9641);
or U9931 (N_9931,N_9696,N_9634);
or U9932 (N_9932,N_9600,N_9726);
or U9933 (N_9933,N_9607,N_9625);
nor U9934 (N_9934,N_9761,N_9749);
or U9935 (N_9935,N_9698,N_9703);
and U9936 (N_9936,N_9689,N_9785);
and U9937 (N_9937,N_9791,N_9605);
nand U9938 (N_9938,N_9629,N_9624);
and U9939 (N_9939,N_9732,N_9758);
nor U9940 (N_9940,N_9701,N_9705);
xnor U9941 (N_9941,N_9743,N_9755);
nand U9942 (N_9942,N_9764,N_9748);
or U9943 (N_9943,N_9691,N_9708);
nand U9944 (N_9944,N_9641,N_9780);
and U9945 (N_9945,N_9696,N_9726);
and U9946 (N_9946,N_9737,N_9705);
and U9947 (N_9947,N_9626,N_9631);
xor U9948 (N_9948,N_9778,N_9676);
or U9949 (N_9949,N_9784,N_9681);
and U9950 (N_9950,N_9645,N_9693);
xor U9951 (N_9951,N_9746,N_9665);
nor U9952 (N_9952,N_9673,N_9698);
xor U9953 (N_9953,N_9607,N_9767);
xnor U9954 (N_9954,N_9698,N_9689);
nor U9955 (N_9955,N_9734,N_9749);
or U9956 (N_9956,N_9781,N_9738);
nand U9957 (N_9957,N_9652,N_9661);
xnor U9958 (N_9958,N_9712,N_9767);
nor U9959 (N_9959,N_9741,N_9794);
xnor U9960 (N_9960,N_9794,N_9649);
and U9961 (N_9961,N_9623,N_9656);
nand U9962 (N_9962,N_9770,N_9658);
or U9963 (N_9963,N_9707,N_9789);
nor U9964 (N_9964,N_9782,N_9780);
nor U9965 (N_9965,N_9716,N_9761);
nor U9966 (N_9966,N_9624,N_9748);
nand U9967 (N_9967,N_9636,N_9683);
or U9968 (N_9968,N_9774,N_9763);
nor U9969 (N_9969,N_9629,N_9680);
nor U9970 (N_9970,N_9682,N_9721);
xnor U9971 (N_9971,N_9604,N_9697);
nand U9972 (N_9972,N_9658,N_9742);
or U9973 (N_9973,N_9726,N_9741);
xor U9974 (N_9974,N_9644,N_9620);
and U9975 (N_9975,N_9669,N_9688);
nor U9976 (N_9976,N_9754,N_9624);
and U9977 (N_9977,N_9765,N_9701);
nand U9978 (N_9978,N_9798,N_9675);
nand U9979 (N_9979,N_9626,N_9634);
nand U9980 (N_9980,N_9728,N_9661);
and U9981 (N_9981,N_9629,N_9761);
nand U9982 (N_9982,N_9647,N_9689);
nor U9983 (N_9983,N_9758,N_9681);
nor U9984 (N_9984,N_9696,N_9790);
and U9985 (N_9985,N_9608,N_9616);
xnor U9986 (N_9986,N_9647,N_9637);
and U9987 (N_9987,N_9741,N_9686);
nor U9988 (N_9988,N_9668,N_9774);
nand U9989 (N_9989,N_9702,N_9611);
or U9990 (N_9990,N_9655,N_9785);
nand U9991 (N_9991,N_9695,N_9606);
or U9992 (N_9992,N_9689,N_9762);
nor U9993 (N_9993,N_9769,N_9768);
nand U9994 (N_9994,N_9678,N_9688);
or U9995 (N_9995,N_9641,N_9634);
and U9996 (N_9996,N_9688,N_9641);
xnor U9997 (N_9997,N_9616,N_9796);
nor U9998 (N_9998,N_9777,N_9759);
and U9999 (N_9999,N_9604,N_9741);
xnor U10000 (N_10000,N_9980,N_9848);
nand U10001 (N_10001,N_9901,N_9997);
xnor U10002 (N_10002,N_9988,N_9884);
xor U10003 (N_10003,N_9913,N_9861);
xor U10004 (N_10004,N_9916,N_9951);
nor U10005 (N_10005,N_9864,N_9829);
and U10006 (N_10006,N_9924,N_9991);
xor U10007 (N_10007,N_9813,N_9915);
nor U10008 (N_10008,N_9961,N_9985);
or U10009 (N_10009,N_9801,N_9932);
nand U10010 (N_10010,N_9954,N_9909);
and U10011 (N_10011,N_9953,N_9823);
nor U10012 (N_10012,N_9993,N_9834);
nand U10013 (N_10013,N_9802,N_9902);
and U10014 (N_10014,N_9847,N_9862);
or U10015 (N_10015,N_9850,N_9979);
nand U10016 (N_10016,N_9892,N_9874);
and U10017 (N_10017,N_9910,N_9875);
and U10018 (N_10018,N_9887,N_9812);
xor U10019 (N_10019,N_9838,N_9858);
xnor U10020 (N_10020,N_9824,N_9950);
and U10021 (N_10021,N_9831,N_9947);
nand U10022 (N_10022,N_9956,N_9878);
or U10023 (N_10023,N_9849,N_9839);
nand U10024 (N_10024,N_9925,N_9906);
nand U10025 (N_10025,N_9904,N_9805);
nand U10026 (N_10026,N_9966,N_9810);
and U10027 (N_10027,N_9994,N_9857);
nor U10028 (N_10028,N_9978,N_9845);
nor U10029 (N_10029,N_9970,N_9869);
and U10030 (N_10030,N_9856,N_9871);
nand U10031 (N_10031,N_9891,N_9975);
and U10032 (N_10032,N_9941,N_9843);
xor U10033 (N_10033,N_9957,N_9804);
xor U10034 (N_10034,N_9882,N_9827);
xor U10035 (N_10035,N_9944,N_9918);
xor U10036 (N_10036,N_9984,N_9836);
xor U10037 (N_10037,N_9952,N_9817);
nand U10038 (N_10038,N_9938,N_9934);
nor U10039 (N_10039,N_9880,N_9982);
nand U10040 (N_10040,N_9972,N_9907);
nand U10041 (N_10041,N_9999,N_9983);
and U10042 (N_10042,N_9976,N_9903);
or U10043 (N_10043,N_9911,N_9899);
nor U10044 (N_10044,N_9822,N_9897);
nor U10045 (N_10045,N_9998,N_9964);
and U10046 (N_10046,N_9940,N_9948);
xor U10047 (N_10047,N_9883,N_9808);
nand U10048 (N_10048,N_9846,N_9917);
or U10049 (N_10049,N_9922,N_9854);
or U10050 (N_10050,N_9830,N_9969);
xor U10051 (N_10051,N_9981,N_9870);
and U10052 (N_10052,N_9990,N_9895);
or U10053 (N_10053,N_9971,N_9927);
nand U10054 (N_10054,N_9877,N_9803);
or U10055 (N_10055,N_9912,N_9986);
nand U10056 (N_10056,N_9898,N_9844);
nand U10057 (N_10057,N_9885,N_9876);
or U10058 (N_10058,N_9888,N_9851);
xor U10059 (N_10059,N_9974,N_9935);
nand U10060 (N_10060,N_9958,N_9929);
xnor U10061 (N_10061,N_9818,N_9942);
nand U10062 (N_10062,N_9853,N_9908);
xnor U10063 (N_10063,N_9893,N_9968);
and U10064 (N_10064,N_9937,N_9811);
xnor U10065 (N_10065,N_9955,N_9814);
xnor U10066 (N_10066,N_9967,N_9867);
and U10067 (N_10067,N_9840,N_9946);
nor U10068 (N_10068,N_9841,N_9914);
xnor U10069 (N_10069,N_9873,N_9842);
or U10070 (N_10070,N_9890,N_9963);
and U10071 (N_10071,N_9820,N_9872);
nand U10072 (N_10072,N_9825,N_9826);
nand U10073 (N_10073,N_9800,N_9949);
or U10074 (N_10074,N_9921,N_9945);
nor U10075 (N_10075,N_9828,N_9960);
nand U10076 (N_10076,N_9933,N_9860);
nor U10077 (N_10077,N_9837,N_9859);
xnor U10078 (N_10078,N_9905,N_9943);
and U10079 (N_10079,N_9928,N_9819);
nor U10080 (N_10080,N_9992,N_9879);
nor U10081 (N_10081,N_9807,N_9931);
and U10082 (N_10082,N_9926,N_9923);
xor U10083 (N_10083,N_9835,N_9894);
or U10084 (N_10084,N_9865,N_9863);
and U10085 (N_10085,N_9806,N_9965);
nor U10086 (N_10086,N_9896,N_9833);
nor U10087 (N_10087,N_9989,N_9973);
xor U10088 (N_10088,N_9881,N_9900);
or U10089 (N_10089,N_9832,N_9919);
xnor U10090 (N_10090,N_9816,N_9889);
and U10091 (N_10091,N_9995,N_9936);
and U10092 (N_10092,N_9886,N_9821);
nand U10093 (N_10093,N_9987,N_9868);
and U10094 (N_10094,N_9977,N_9920);
or U10095 (N_10095,N_9959,N_9996);
nor U10096 (N_10096,N_9809,N_9855);
nand U10097 (N_10097,N_9930,N_9866);
nand U10098 (N_10098,N_9939,N_9815);
xnor U10099 (N_10099,N_9852,N_9962);
and U10100 (N_10100,N_9830,N_9923);
or U10101 (N_10101,N_9867,N_9923);
or U10102 (N_10102,N_9827,N_9865);
and U10103 (N_10103,N_9986,N_9858);
and U10104 (N_10104,N_9950,N_9923);
xnor U10105 (N_10105,N_9815,N_9975);
nor U10106 (N_10106,N_9882,N_9958);
xnor U10107 (N_10107,N_9992,N_9964);
nor U10108 (N_10108,N_9817,N_9945);
xnor U10109 (N_10109,N_9839,N_9935);
xnor U10110 (N_10110,N_9956,N_9884);
nand U10111 (N_10111,N_9982,N_9929);
nand U10112 (N_10112,N_9824,N_9961);
nor U10113 (N_10113,N_9897,N_9818);
or U10114 (N_10114,N_9862,N_9871);
and U10115 (N_10115,N_9885,N_9824);
xnor U10116 (N_10116,N_9802,N_9986);
or U10117 (N_10117,N_9841,N_9875);
and U10118 (N_10118,N_9967,N_9912);
and U10119 (N_10119,N_9991,N_9831);
and U10120 (N_10120,N_9935,N_9976);
or U10121 (N_10121,N_9989,N_9813);
and U10122 (N_10122,N_9929,N_9806);
and U10123 (N_10123,N_9888,N_9957);
nand U10124 (N_10124,N_9993,N_9935);
nand U10125 (N_10125,N_9967,N_9909);
and U10126 (N_10126,N_9933,N_9825);
nor U10127 (N_10127,N_9821,N_9865);
nor U10128 (N_10128,N_9851,N_9874);
nand U10129 (N_10129,N_9910,N_9918);
or U10130 (N_10130,N_9917,N_9883);
nor U10131 (N_10131,N_9862,N_9829);
nand U10132 (N_10132,N_9825,N_9932);
xor U10133 (N_10133,N_9811,N_9843);
and U10134 (N_10134,N_9956,N_9900);
xnor U10135 (N_10135,N_9950,N_9848);
nand U10136 (N_10136,N_9892,N_9944);
or U10137 (N_10137,N_9859,N_9844);
nand U10138 (N_10138,N_9974,N_9902);
or U10139 (N_10139,N_9882,N_9903);
xnor U10140 (N_10140,N_9949,N_9882);
and U10141 (N_10141,N_9877,N_9857);
nor U10142 (N_10142,N_9974,N_9908);
xnor U10143 (N_10143,N_9810,N_9941);
xnor U10144 (N_10144,N_9822,N_9847);
and U10145 (N_10145,N_9894,N_9874);
nor U10146 (N_10146,N_9828,N_9867);
nor U10147 (N_10147,N_9954,N_9830);
or U10148 (N_10148,N_9911,N_9860);
nand U10149 (N_10149,N_9864,N_9882);
nor U10150 (N_10150,N_9846,N_9960);
or U10151 (N_10151,N_9975,N_9996);
or U10152 (N_10152,N_9970,N_9894);
nor U10153 (N_10153,N_9859,N_9912);
or U10154 (N_10154,N_9894,N_9948);
or U10155 (N_10155,N_9825,N_9948);
nor U10156 (N_10156,N_9878,N_9841);
xnor U10157 (N_10157,N_9819,N_9884);
and U10158 (N_10158,N_9846,N_9841);
or U10159 (N_10159,N_9927,N_9982);
nand U10160 (N_10160,N_9933,N_9945);
xnor U10161 (N_10161,N_9805,N_9992);
nand U10162 (N_10162,N_9941,N_9841);
nand U10163 (N_10163,N_9926,N_9898);
nand U10164 (N_10164,N_9931,N_9947);
xnor U10165 (N_10165,N_9911,N_9984);
xnor U10166 (N_10166,N_9959,N_9900);
xnor U10167 (N_10167,N_9847,N_9860);
and U10168 (N_10168,N_9990,N_9884);
or U10169 (N_10169,N_9879,N_9943);
nor U10170 (N_10170,N_9839,N_9910);
nor U10171 (N_10171,N_9806,N_9902);
or U10172 (N_10172,N_9904,N_9857);
nor U10173 (N_10173,N_9951,N_9864);
nor U10174 (N_10174,N_9964,N_9865);
and U10175 (N_10175,N_9970,N_9857);
nor U10176 (N_10176,N_9870,N_9989);
xor U10177 (N_10177,N_9902,N_9851);
xor U10178 (N_10178,N_9977,N_9987);
nand U10179 (N_10179,N_9991,N_9949);
xnor U10180 (N_10180,N_9863,N_9851);
or U10181 (N_10181,N_9827,N_9976);
xnor U10182 (N_10182,N_9857,N_9825);
xnor U10183 (N_10183,N_9812,N_9817);
nor U10184 (N_10184,N_9826,N_9801);
nand U10185 (N_10185,N_9966,N_9818);
and U10186 (N_10186,N_9989,N_9921);
nor U10187 (N_10187,N_9859,N_9857);
and U10188 (N_10188,N_9951,N_9954);
and U10189 (N_10189,N_9873,N_9964);
xor U10190 (N_10190,N_9876,N_9972);
and U10191 (N_10191,N_9942,N_9848);
or U10192 (N_10192,N_9820,N_9875);
and U10193 (N_10193,N_9866,N_9924);
nand U10194 (N_10194,N_9923,N_9857);
xnor U10195 (N_10195,N_9813,N_9934);
nor U10196 (N_10196,N_9814,N_9821);
or U10197 (N_10197,N_9985,N_9940);
and U10198 (N_10198,N_9814,N_9944);
nor U10199 (N_10199,N_9871,N_9992);
nor U10200 (N_10200,N_10049,N_10123);
xor U10201 (N_10201,N_10050,N_10037);
nand U10202 (N_10202,N_10044,N_10083);
and U10203 (N_10203,N_10002,N_10052);
nand U10204 (N_10204,N_10017,N_10026);
and U10205 (N_10205,N_10032,N_10180);
and U10206 (N_10206,N_10139,N_10035);
nor U10207 (N_10207,N_10100,N_10133);
and U10208 (N_10208,N_10014,N_10195);
nor U10209 (N_10209,N_10092,N_10149);
and U10210 (N_10210,N_10169,N_10001);
nand U10211 (N_10211,N_10160,N_10068);
nor U10212 (N_10212,N_10134,N_10057);
nand U10213 (N_10213,N_10129,N_10082);
nor U10214 (N_10214,N_10010,N_10033);
or U10215 (N_10215,N_10125,N_10179);
and U10216 (N_10216,N_10110,N_10076);
or U10217 (N_10217,N_10011,N_10086);
xnor U10218 (N_10218,N_10025,N_10194);
or U10219 (N_10219,N_10174,N_10126);
or U10220 (N_10220,N_10150,N_10059);
and U10221 (N_10221,N_10113,N_10103);
nor U10222 (N_10222,N_10102,N_10114);
or U10223 (N_10223,N_10081,N_10198);
nand U10224 (N_10224,N_10043,N_10003);
xor U10225 (N_10225,N_10028,N_10094);
nor U10226 (N_10226,N_10085,N_10185);
nand U10227 (N_10227,N_10093,N_10196);
or U10228 (N_10228,N_10004,N_10173);
and U10229 (N_10229,N_10170,N_10062);
nand U10230 (N_10230,N_10140,N_10060);
xnor U10231 (N_10231,N_10005,N_10088);
xor U10232 (N_10232,N_10168,N_10029);
xor U10233 (N_10233,N_10018,N_10143);
xnor U10234 (N_10234,N_10188,N_10144);
or U10235 (N_10235,N_10090,N_10105);
nor U10236 (N_10236,N_10084,N_10159);
xor U10237 (N_10237,N_10131,N_10146);
nand U10238 (N_10238,N_10022,N_10071);
nand U10239 (N_10239,N_10053,N_10064);
and U10240 (N_10240,N_10027,N_10070);
xnor U10241 (N_10241,N_10163,N_10192);
and U10242 (N_10242,N_10075,N_10167);
and U10243 (N_10243,N_10189,N_10136);
or U10244 (N_10244,N_10184,N_10069);
or U10245 (N_10245,N_10041,N_10145);
xor U10246 (N_10246,N_10045,N_10152);
xor U10247 (N_10247,N_10137,N_10008);
nor U10248 (N_10248,N_10116,N_10165);
or U10249 (N_10249,N_10095,N_10048);
and U10250 (N_10250,N_10073,N_10074);
nand U10251 (N_10251,N_10183,N_10036);
or U10252 (N_10252,N_10106,N_10030);
or U10253 (N_10253,N_10024,N_10120);
or U10254 (N_10254,N_10007,N_10079);
xor U10255 (N_10255,N_10066,N_10199);
xnor U10256 (N_10256,N_10040,N_10181);
nor U10257 (N_10257,N_10031,N_10191);
or U10258 (N_10258,N_10063,N_10186);
or U10259 (N_10259,N_10067,N_10099);
xnor U10260 (N_10260,N_10121,N_10019);
or U10261 (N_10261,N_10111,N_10112);
xnor U10262 (N_10262,N_10177,N_10171);
xnor U10263 (N_10263,N_10020,N_10157);
nand U10264 (N_10264,N_10117,N_10096);
nor U10265 (N_10265,N_10098,N_10118);
and U10266 (N_10266,N_10142,N_10193);
and U10267 (N_10267,N_10172,N_10147);
or U10268 (N_10268,N_10166,N_10078);
xor U10269 (N_10269,N_10135,N_10176);
xnor U10270 (N_10270,N_10042,N_10023);
nor U10271 (N_10271,N_10175,N_10006);
nor U10272 (N_10272,N_10012,N_10000);
and U10273 (N_10273,N_10155,N_10108);
nand U10274 (N_10274,N_10162,N_10089);
nand U10275 (N_10275,N_10154,N_10039);
nand U10276 (N_10276,N_10130,N_10056);
xor U10277 (N_10277,N_10187,N_10128);
nor U10278 (N_10278,N_10141,N_10080);
nand U10279 (N_10279,N_10087,N_10046);
nor U10280 (N_10280,N_10101,N_10124);
or U10281 (N_10281,N_10156,N_10158);
and U10282 (N_10282,N_10051,N_10077);
or U10283 (N_10283,N_10015,N_10058);
nand U10284 (N_10284,N_10072,N_10148);
xnor U10285 (N_10285,N_10013,N_10151);
or U10286 (N_10286,N_10065,N_10061);
nand U10287 (N_10287,N_10034,N_10107);
and U10288 (N_10288,N_10021,N_10197);
nand U10289 (N_10289,N_10119,N_10054);
nor U10290 (N_10290,N_10164,N_10104);
and U10291 (N_10291,N_10122,N_10016);
xnor U10292 (N_10292,N_10190,N_10009);
xnor U10293 (N_10293,N_10115,N_10097);
nor U10294 (N_10294,N_10178,N_10109);
nand U10295 (N_10295,N_10153,N_10055);
nor U10296 (N_10296,N_10091,N_10132);
nand U10297 (N_10297,N_10161,N_10182);
and U10298 (N_10298,N_10138,N_10038);
xor U10299 (N_10299,N_10047,N_10127);
nor U10300 (N_10300,N_10166,N_10128);
xor U10301 (N_10301,N_10112,N_10024);
nand U10302 (N_10302,N_10181,N_10176);
nor U10303 (N_10303,N_10110,N_10133);
or U10304 (N_10304,N_10167,N_10124);
and U10305 (N_10305,N_10123,N_10191);
nor U10306 (N_10306,N_10008,N_10095);
xnor U10307 (N_10307,N_10132,N_10101);
and U10308 (N_10308,N_10182,N_10007);
and U10309 (N_10309,N_10060,N_10013);
xnor U10310 (N_10310,N_10196,N_10137);
xor U10311 (N_10311,N_10147,N_10184);
nor U10312 (N_10312,N_10189,N_10142);
or U10313 (N_10313,N_10011,N_10196);
and U10314 (N_10314,N_10100,N_10155);
or U10315 (N_10315,N_10084,N_10068);
xor U10316 (N_10316,N_10111,N_10163);
and U10317 (N_10317,N_10115,N_10183);
xor U10318 (N_10318,N_10005,N_10136);
nand U10319 (N_10319,N_10157,N_10056);
xor U10320 (N_10320,N_10016,N_10118);
or U10321 (N_10321,N_10128,N_10178);
or U10322 (N_10322,N_10056,N_10033);
nor U10323 (N_10323,N_10022,N_10196);
or U10324 (N_10324,N_10174,N_10110);
nand U10325 (N_10325,N_10038,N_10082);
nand U10326 (N_10326,N_10032,N_10139);
nor U10327 (N_10327,N_10041,N_10137);
xor U10328 (N_10328,N_10003,N_10101);
xnor U10329 (N_10329,N_10020,N_10152);
nor U10330 (N_10330,N_10174,N_10084);
or U10331 (N_10331,N_10165,N_10177);
nand U10332 (N_10332,N_10035,N_10100);
and U10333 (N_10333,N_10078,N_10163);
nand U10334 (N_10334,N_10127,N_10005);
nand U10335 (N_10335,N_10068,N_10109);
nand U10336 (N_10336,N_10144,N_10182);
or U10337 (N_10337,N_10059,N_10196);
and U10338 (N_10338,N_10176,N_10189);
and U10339 (N_10339,N_10122,N_10161);
xor U10340 (N_10340,N_10114,N_10095);
nor U10341 (N_10341,N_10184,N_10095);
xor U10342 (N_10342,N_10043,N_10024);
xor U10343 (N_10343,N_10190,N_10069);
and U10344 (N_10344,N_10175,N_10168);
or U10345 (N_10345,N_10092,N_10170);
xor U10346 (N_10346,N_10166,N_10132);
nand U10347 (N_10347,N_10195,N_10180);
nor U10348 (N_10348,N_10186,N_10106);
or U10349 (N_10349,N_10105,N_10077);
xor U10350 (N_10350,N_10054,N_10153);
nor U10351 (N_10351,N_10091,N_10133);
nor U10352 (N_10352,N_10061,N_10113);
xnor U10353 (N_10353,N_10128,N_10062);
nand U10354 (N_10354,N_10194,N_10046);
nand U10355 (N_10355,N_10162,N_10175);
xnor U10356 (N_10356,N_10086,N_10127);
nor U10357 (N_10357,N_10015,N_10130);
or U10358 (N_10358,N_10199,N_10187);
and U10359 (N_10359,N_10039,N_10189);
xnor U10360 (N_10360,N_10176,N_10134);
nand U10361 (N_10361,N_10108,N_10156);
or U10362 (N_10362,N_10059,N_10141);
nor U10363 (N_10363,N_10133,N_10007);
and U10364 (N_10364,N_10091,N_10004);
nor U10365 (N_10365,N_10192,N_10055);
and U10366 (N_10366,N_10172,N_10085);
and U10367 (N_10367,N_10162,N_10036);
nand U10368 (N_10368,N_10022,N_10081);
nor U10369 (N_10369,N_10143,N_10006);
nand U10370 (N_10370,N_10063,N_10105);
or U10371 (N_10371,N_10154,N_10063);
or U10372 (N_10372,N_10043,N_10037);
nand U10373 (N_10373,N_10033,N_10001);
xor U10374 (N_10374,N_10135,N_10186);
xnor U10375 (N_10375,N_10175,N_10069);
xor U10376 (N_10376,N_10025,N_10099);
or U10377 (N_10377,N_10108,N_10075);
nor U10378 (N_10378,N_10123,N_10057);
xnor U10379 (N_10379,N_10129,N_10193);
nor U10380 (N_10380,N_10045,N_10150);
nor U10381 (N_10381,N_10023,N_10151);
xor U10382 (N_10382,N_10082,N_10131);
or U10383 (N_10383,N_10099,N_10122);
nand U10384 (N_10384,N_10073,N_10186);
and U10385 (N_10385,N_10180,N_10130);
nand U10386 (N_10386,N_10029,N_10010);
and U10387 (N_10387,N_10046,N_10088);
nand U10388 (N_10388,N_10136,N_10064);
and U10389 (N_10389,N_10195,N_10181);
xnor U10390 (N_10390,N_10046,N_10023);
or U10391 (N_10391,N_10022,N_10152);
nor U10392 (N_10392,N_10171,N_10076);
xor U10393 (N_10393,N_10029,N_10150);
and U10394 (N_10394,N_10133,N_10085);
or U10395 (N_10395,N_10072,N_10133);
and U10396 (N_10396,N_10030,N_10003);
or U10397 (N_10397,N_10036,N_10126);
or U10398 (N_10398,N_10002,N_10086);
xor U10399 (N_10399,N_10157,N_10121);
and U10400 (N_10400,N_10386,N_10250);
nand U10401 (N_10401,N_10236,N_10204);
nand U10402 (N_10402,N_10328,N_10226);
nor U10403 (N_10403,N_10244,N_10373);
nor U10404 (N_10404,N_10238,N_10214);
xnor U10405 (N_10405,N_10206,N_10310);
nand U10406 (N_10406,N_10395,N_10273);
nand U10407 (N_10407,N_10257,N_10308);
and U10408 (N_10408,N_10252,N_10378);
and U10409 (N_10409,N_10247,N_10360);
nor U10410 (N_10410,N_10325,N_10279);
and U10411 (N_10411,N_10233,N_10393);
nand U10412 (N_10412,N_10202,N_10292);
and U10413 (N_10413,N_10220,N_10394);
xor U10414 (N_10414,N_10383,N_10303);
and U10415 (N_10415,N_10346,N_10242);
nor U10416 (N_10416,N_10299,N_10230);
nand U10417 (N_10417,N_10262,N_10245);
nor U10418 (N_10418,N_10267,N_10305);
or U10419 (N_10419,N_10237,N_10203);
and U10420 (N_10420,N_10352,N_10243);
or U10421 (N_10421,N_10307,N_10348);
and U10422 (N_10422,N_10336,N_10218);
nand U10423 (N_10423,N_10283,N_10340);
and U10424 (N_10424,N_10304,N_10228);
or U10425 (N_10425,N_10248,N_10370);
xnor U10426 (N_10426,N_10268,N_10358);
nor U10427 (N_10427,N_10350,N_10372);
nand U10428 (N_10428,N_10335,N_10381);
nand U10429 (N_10429,N_10210,N_10334);
nand U10430 (N_10430,N_10282,N_10391);
or U10431 (N_10431,N_10365,N_10338);
xnor U10432 (N_10432,N_10392,N_10314);
and U10433 (N_10433,N_10219,N_10294);
nand U10434 (N_10434,N_10285,N_10264);
and U10435 (N_10435,N_10270,N_10213);
and U10436 (N_10436,N_10260,N_10398);
or U10437 (N_10437,N_10315,N_10209);
or U10438 (N_10438,N_10362,N_10255);
nor U10439 (N_10439,N_10227,N_10345);
or U10440 (N_10440,N_10318,N_10229);
xor U10441 (N_10441,N_10211,N_10387);
nand U10442 (N_10442,N_10259,N_10367);
and U10443 (N_10443,N_10239,N_10256);
xor U10444 (N_10444,N_10216,N_10368);
and U10445 (N_10445,N_10297,N_10207);
nor U10446 (N_10446,N_10208,N_10385);
nor U10447 (N_10447,N_10361,N_10374);
nor U10448 (N_10448,N_10384,N_10287);
xnor U10449 (N_10449,N_10277,N_10275);
xnor U10450 (N_10450,N_10399,N_10389);
nor U10451 (N_10451,N_10309,N_10377);
or U10452 (N_10452,N_10357,N_10349);
and U10453 (N_10453,N_10326,N_10354);
nor U10454 (N_10454,N_10344,N_10313);
nor U10455 (N_10455,N_10369,N_10330);
xnor U10456 (N_10456,N_10333,N_10272);
nor U10457 (N_10457,N_10343,N_10281);
or U10458 (N_10458,N_10331,N_10397);
nor U10459 (N_10459,N_10274,N_10390);
xor U10460 (N_10460,N_10376,N_10254);
nor U10461 (N_10461,N_10311,N_10280);
or U10462 (N_10462,N_10234,N_10327);
nor U10463 (N_10463,N_10266,N_10312);
nor U10464 (N_10464,N_10251,N_10261);
nand U10465 (N_10465,N_10364,N_10271);
xor U10466 (N_10466,N_10321,N_10396);
nor U10467 (N_10467,N_10291,N_10293);
nor U10468 (N_10468,N_10356,N_10363);
xor U10469 (N_10469,N_10355,N_10359);
or U10470 (N_10470,N_10222,N_10288);
nand U10471 (N_10471,N_10205,N_10225);
nand U10472 (N_10472,N_10323,N_10380);
and U10473 (N_10473,N_10286,N_10375);
and U10474 (N_10474,N_10301,N_10235);
nand U10475 (N_10475,N_10341,N_10221);
nand U10476 (N_10476,N_10246,N_10332);
xor U10477 (N_10477,N_10290,N_10351);
or U10478 (N_10478,N_10249,N_10329);
nor U10479 (N_10479,N_10379,N_10241);
nor U10480 (N_10480,N_10296,N_10324);
xor U10481 (N_10481,N_10353,N_10265);
or U10482 (N_10482,N_10366,N_10223);
xor U10483 (N_10483,N_10322,N_10382);
or U10484 (N_10484,N_10284,N_10240);
or U10485 (N_10485,N_10231,N_10295);
nand U10486 (N_10486,N_10342,N_10388);
or U10487 (N_10487,N_10269,N_10316);
nand U10488 (N_10488,N_10258,N_10320);
or U10489 (N_10489,N_10200,N_10347);
nand U10490 (N_10490,N_10319,N_10224);
xnor U10491 (N_10491,N_10302,N_10298);
or U10492 (N_10492,N_10212,N_10215);
and U10493 (N_10493,N_10263,N_10276);
nor U10494 (N_10494,N_10317,N_10201);
xor U10495 (N_10495,N_10339,N_10289);
and U10496 (N_10496,N_10232,N_10300);
or U10497 (N_10497,N_10253,N_10371);
xnor U10498 (N_10498,N_10306,N_10217);
and U10499 (N_10499,N_10337,N_10278);
xor U10500 (N_10500,N_10308,N_10390);
xnor U10501 (N_10501,N_10244,N_10223);
and U10502 (N_10502,N_10264,N_10399);
or U10503 (N_10503,N_10201,N_10338);
or U10504 (N_10504,N_10296,N_10338);
or U10505 (N_10505,N_10314,N_10296);
nor U10506 (N_10506,N_10236,N_10325);
nand U10507 (N_10507,N_10390,N_10303);
nor U10508 (N_10508,N_10238,N_10210);
nor U10509 (N_10509,N_10250,N_10313);
nand U10510 (N_10510,N_10373,N_10387);
nand U10511 (N_10511,N_10305,N_10222);
or U10512 (N_10512,N_10368,N_10372);
nand U10513 (N_10513,N_10388,N_10233);
xor U10514 (N_10514,N_10378,N_10397);
and U10515 (N_10515,N_10233,N_10298);
nor U10516 (N_10516,N_10308,N_10301);
xor U10517 (N_10517,N_10366,N_10263);
and U10518 (N_10518,N_10375,N_10224);
xor U10519 (N_10519,N_10240,N_10350);
xnor U10520 (N_10520,N_10350,N_10368);
xor U10521 (N_10521,N_10200,N_10202);
nand U10522 (N_10522,N_10207,N_10268);
and U10523 (N_10523,N_10392,N_10237);
nand U10524 (N_10524,N_10338,N_10219);
and U10525 (N_10525,N_10304,N_10351);
xnor U10526 (N_10526,N_10356,N_10352);
nor U10527 (N_10527,N_10322,N_10383);
xnor U10528 (N_10528,N_10253,N_10316);
nand U10529 (N_10529,N_10280,N_10283);
nor U10530 (N_10530,N_10218,N_10334);
or U10531 (N_10531,N_10251,N_10274);
nor U10532 (N_10532,N_10338,N_10223);
xor U10533 (N_10533,N_10344,N_10213);
nand U10534 (N_10534,N_10295,N_10208);
xor U10535 (N_10535,N_10376,N_10369);
or U10536 (N_10536,N_10218,N_10327);
xor U10537 (N_10537,N_10273,N_10243);
xor U10538 (N_10538,N_10219,N_10226);
or U10539 (N_10539,N_10358,N_10264);
xor U10540 (N_10540,N_10224,N_10286);
nand U10541 (N_10541,N_10292,N_10332);
or U10542 (N_10542,N_10349,N_10358);
nand U10543 (N_10543,N_10277,N_10237);
xnor U10544 (N_10544,N_10343,N_10230);
and U10545 (N_10545,N_10225,N_10279);
and U10546 (N_10546,N_10273,N_10211);
and U10547 (N_10547,N_10284,N_10387);
nand U10548 (N_10548,N_10298,N_10356);
nand U10549 (N_10549,N_10270,N_10352);
or U10550 (N_10550,N_10248,N_10202);
and U10551 (N_10551,N_10318,N_10351);
and U10552 (N_10552,N_10310,N_10348);
and U10553 (N_10553,N_10288,N_10347);
xnor U10554 (N_10554,N_10331,N_10392);
or U10555 (N_10555,N_10289,N_10219);
xnor U10556 (N_10556,N_10211,N_10388);
or U10557 (N_10557,N_10379,N_10239);
nand U10558 (N_10558,N_10296,N_10284);
or U10559 (N_10559,N_10352,N_10287);
and U10560 (N_10560,N_10328,N_10257);
nor U10561 (N_10561,N_10299,N_10288);
or U10562 (N_10562,N_10311,N_10383);
nor U10563 (N_10563,N_10298,N_10359);
or U10564 (N_10564,N_10250,N_10315);
and U10565 (N_10565,N_10281,N_10245);
nand U10566 (N_10566,N_10351,N_10282);
or U10567 (N_10567,N_10398,N_10360);
xor U10568 (N_10568,N_10282,N_10399);
and U10569 (N_10569,N_10352,N_10218);
nor U10570 (N_10570,N_10349,N_10352);
and U10571 (N_10571,N_10245,N_10389);
or U10572 (N_10572,N_10277,N_10312);
and U10573 (N_10573,N_10353,N_10286);
or U10574 (N_10574,N_10216,N_10343);
and U10575 (N_10575,N_10349,N_10347);
nand U10576 (N_10576,N_10375,N_10264);
nor U10577 (N_10577,N_10329,N_10370);
xnor U10578 (N_10578,N_10233,N_10361);
xnor U10579 (N_10579,N_10224,N_10376);
nor U10580 (N_10580,N_10277,N_10215);
nand U10581 (N_10581,N_10285,N_10216);
nor U10582 (N_10582,N_10335,N_10328);
nor U10583 (N_10583,N_10322,N_10289);
or U10584 (N_10584,N_10309,N_10349);
nor U10585 (N_10585,N_10277,N_10271);
nor U10586 (N_10586,N_10305,N_10290);
nand U10587 (N_10587,N_10396,N_10324);
and U10588 (N_10588,N_10322,N_10273);
and U10589 (N_10589,N_10229,N_10321);
and U10590 (N_10590,N_10273,N_10316);
nor U10591 (N_10591,N_10248,N_10332);
nor U10592 (N_10592,N_10341,N_10301);
xnor U10593 (N_10593,N_10244,N_10257);
or U10594 (N_10594,N_10200,N_10361);
nand U10595 (N_10595,N_10379,N_10264);
xor U10596 (N_10596,N_10359,N_10364);
nor U10597 (N_10597,N_10309,N_10396);
nor U10598 (N_10598,N_10280,N_10222);
nor U10599 (N_10599,N_10324,N_10222);
xnor U10600 (N_10600,N_10585,N_10452);
nand U10601 (N_10601,N_10539,N_10472);
nor U10602 (N_10602,N_10569,N_10430);
nor U10603 (N_10603,N_10525,N_10542);
and U10604 (N_10604,N_10449,N_10405);
nand U10605 (N_10605,N_10415,N_10416);
xor U10606 (N_10606,N_10473,N_10543);
nor U10607 (N_10607,N_10445,N_10424);
xor U10608 (N_10608,N_10481,N_10514);
and U10609 (N_10609,N_10588,N_10531);
xor U10610 (N_10610,N_10412,N_10470);
nor U10611 (N_10611,N_10511,N_10437);
or U10612 (N_10612,N_10439,N_10598);
or U10613 (N_10613,N_10435,N_10597);
nor U10614 (N_10614,N_10480,N_10519);
or U10615 (N_10615,N_10518,N_10501);
or U10616 (N_10616,N_10595,N_10410);
and U10617 (N_10617,N_10419,N_10450);
xor U10618 (N_10618,N_10478,N_10546);
and U10619 (N_10619,N_10568,N_10491);
or U10620 (N_10620,N_10429,N_10565);
or U10621 (N_10621,N_10502,N_10516);
nor U10622 (N_10622,N_10469,N_10426);
and U10623 (N_10623,N_10455,N_10488);
nand U10624 (N_10624,N_10587,N_10510);
nor U10625 (N_10625,N_10497,N_10484);
and U10626 (N_10626,N_10522,N_10548);
xnor U10627 (N_10627,N_10592,N_10557);
nor U10628 (N_10628,N_10456,N_10537);
xor U10629 (N_10629,N_10536,N_10538);
nand U10630 (N_10630,N_10505,N_10549);
nor U10631 (N_10631,N_10579,N_10483);
nand U10632 (N_10632,N_10425,N_10485);
xnor U10633 (N_10633,N_10432,N_10570);
nand U10634 (N_10634,N_10513,N_10583);
nand U10635 (N_10635,N_10431,N_10494);
xnor U10636 (N_10636,N_10508,N_10457);
or U10637 (N_10637,N_10423,N_10418);
nor U10638 (N_10638,N_10413,N_10599);
or U10639 (N_10639,N_10477,N_10551);
and U10640 (N_10640,N_10500,N_10401);
xor U10641 (N_10641,N_10581,N_10409);
nor U10642 (N_10642,N_10554,N_10521);
nor U10643 (N_10643,N_10540,N_10556);
and U10644 (N_10644,N_10489,N_10560);
nor U10645 (N_10645,N_10520,N_10532);
nor U10646 (N_10646,N_10572,N_10421);
nand U10647 (N_10647,N_10553,N_10468);
xnor U10648 (N_10648,N_10461,N_10517);
xnor U10649 (N_10649,N_10467,N_10534);
xor U10650 (N_10650,N_10564,N_10594);
and U10651 (N_10651,N_10448,N_10503);
xor U10652 (N_10652,N_10411,N_10400);
xnor U10653 (N_10653,N_10582,N_10466);
nand U10654 (N_10654,N_10440,N_10465);
and U10655 (N_10655,N_10545,N_10479);
and U10656 (N_10656,N_10530,N_10577);
nor U10657 (N_10657,N_10447,N_10566);
or U10658 (N_10658,N_10561,N_10417);
nor U10659 (N_10659,N_10490,N_10506);
xor U10660 (N_10660,N_10573,N_10535);
and U10661 (N_10661,N_10575,N_10509);
nor U10662 (N_10662,N_10458,N_10471);
nor U10663 (N_10663,N_10527,N_10591);
or U10664 (N_10664,N_10451,N_10571);
and U10665 (N_10665,N_10404,N_10406);
xnor U10666 (N_10666,N_10402,N_10562);
nor U10667 (N_10667,N_10499,N_10574);
nor U10668 (N_10668,N_10563,N_10463);
nand U10669 (N_10669,N_10550,N_10475);
nand U10670 (N_10670,N_10487,N_10407);
and U10671 (N_10671,N_10524,N_10558);
and U10672 (N_10672,N_10444,N_10459);
or U10673 (N_10673,N_10441,N_10474);
xnor U10674 (N_10674,N_10462,N_10453);
or U10675 (N_10675,N_10576,N_10541);
xor U10676 (N_10676,N_10454,N_10434);
xnor U10677 (N_10677,N_10464,N_10414);
xnor U10678 (N_10678,N_10420,N_10493);
xor U10679 (N_10679,N_10504,N_10515);
or U10680 (N_10680,N_10433,N_10442);
or U10681 (N_10681,N_10559,N_10523);
and U10682 (N_10682,N_10486,N_10584);
nand U10683 (N_10683,N_10496,N_10567);
or U10684 (N_10684,N_10552,N_10446);
nor U10685 (N_10685,N_10593,N_10492);
nor U10686 (N_10686,N_10526,N_10436);
xor U10687 (N_10687,N_10555,N_10578);
or U10688 (N_10688,N_10512,N_10408);
or U10689 (N_10689,N_10460,N_10547);
nor U10690 (N_10690,N_10482,N_10427);
nor U10691 (N_10691,N_10590,N_10476);
nand U10692 (N_10692,N_10586,N_10589);
nand U10693 (N_10693,N_10443,N_10403);
or U10694 (N_10694,N_10428,N_10498);
xor U10695 (N_10695,N_10529,N_10438);
and U10696 (N_10696,N_10507,N_10528);
and U10697 (N_10697,N_10533,N_10596);
nand U10698 (N_10698,N_10422,N_10580);
nor U10699 (N_10699,N_10544,N_10495);
xnor U10700 (N_10700,N_10589,N_10590);
nand U10701 (N_10701,N_10596,N_10489);
nor U10702 (N_10702,N_10539,N_10514);
or U10703 (N_10703,N_10585,N_10549);
nand U10704 (N_10704,N_10410,N_10464);
and U10705 (N_10705,N_10434,N_10554);
nand U10706 (N_10706,N_10406,N_10563);
nor U10707 (N_10707,N_10408,N_10518);
and U10708 (N_10708,N_10460,N_10415);
or U10709 (N_10709,N_10546,N_10587);
xor U10710 (N_10710,N_10531,N_10538);
xnor U10711 (N_10711,N_10557,N_10488);
and U10712 (N_10712,N_10513,N_10534);
nand U10713 (N_10713,N_10592,N_10492);
or U10714 (N_10714,N_10438,N_10568);
and U10715 (N_10715,N_10539,N_10425);
nor U10716 (N_10716,N_10481,N_10496);
and U10717 (N_10717,N_10518,N_10444);
nand U10718 (N_10718,N_10576,N_10580);
nor U10719 (N_10719,N_10477,N_10401);
nor U10720 (N_10720,N_10476,N_10546);
nand U10721 (N_10721,N_10555,N_10400);
and U10722 (N_10722,N_10400,N_10503);
and U10723 (N_10723,N_10582,N_10551);
nor U10724 (N_10724,N_10521,N_10583);
or U10725 (N_10725,N_10427,N_10525);
or U10726 (N_10726,N_10565,N_10489);
or U10727 (N_10727,N_10558,N_10581);
nand U10728 (N_10728,N_10423,N_10540);
nor U10729 (N_10729,N_10476,N_10472);
and U10730 (N_10730,N_10466,N_10530);
nor U10731 (N_10731,N_10519,N_10447);
xnor U10732 (N_10732,N_10464,N_10470);
xor U10733 (N_10733,N_10556,N_10433);
xor U10734 (N_10734,N_10553,N_10585);
xor U10735 (N_10735,N_10578,N_10551);
or U10736 (N_10736,N_10419,N_10453);
nor U10737 (N_10737,N_10591,N_10555);
and U10738 (N_10738,N_10540,N_10419);
or U10739 (N_10739,N_10442,N_10406);
and U10740 (N_10740,N_10430,N_10496);
or U10741 (N_10741,N_10474,N_10404);
nor U10742 (N_10742,N_10578,N_10481);
or U10743 (N_10743,N_10572,N_10590);
or U10744 (N_10744,N_10426,N_10412);
nand U10745 (N_10745,N_10412,N_10409);
nor U10746 (N_10746,N_10501,N_10514);
xnor U10747 (N_10747,N_10568,N_10531);
nor U10748 (N_10748,N_10540,N_10533);
or U10749 (N_10749,N_10485,N_10450);
and U10750 (N_10750,N_10563,N_10431);
xor U10751 (N_10751,N_10412,N_10552);
or U10752 (N_10752,N_10491,N_10437);
and U10753 (N_10753,N_10469,N_10453);
nor U10754 (N_10754,N_10572,N_10538);
xnor U10755 (N_10755,N_10415,N_10492);
nor U10756 (N_10756,N_10525,N_10557);
xor U10757 (N_10757,N_10436,N_10473);
or U10758 (N_10758,N_10407,N_10540);
nand U10759 (N_10759,N_10444,N_10498);
nand U10760 (N_10760,N_10588,N_10433);
nand U10761 (N_10761,N_10588,N_10524);
xor U10762 (N_10762,N_10445,N_10556);
and U10763 (N_10763,N_10459,N_10461);
or U10764 (N_10764,N_10590,N_10419);
xor U10765 (N_10765,N_10447,N_10508);
xnor U10766 (N_10766,N_10432,N_10414);
and U10767 (N_10767,N_10591,N_10429);
nand U10768 (N_10768,N_10508,N_10459);
or U10769 (N_10769,N_10556,N_10440);
xor U10770 (N_10770,N_10411,N_10416);
and U10771 (N_10771,N_10404,N_10593);
nor U10772 (N_10772,N_10586,N_10452);
nor U10773 (N_10773,N_10472,N_10575);
and U10774 (N_10774,N_10421,N_10524);
nor U10775 (N_10775,N_10451,N_10520);
or U10776 (N_10776,N_10584,N_10414);
or U10777 (N_10777,N_10428,N_10584);
nand U10778 (N_10778,N_10566,N_10405);
nor U10779 (N_10779,N_10565,N_10566);
nand U10780 (N_10780,N_10585,N_10464);
xnor U10781 (N_10781,N_10441,N_10476);
and U10782 (N_10782,N_10419,N_10512);
and U10783 (N_10783,N_10550,N_10455);
nor U10784 (N_10784,N_10461,N_10549);
xnor U10785 (N_10785,N_10443,N_10535);
and U10786 (N_10786,N_10511,N_10464);
xor U10787 (N_10787,N_10554,N_10440);
and U10788 (N_10788,N_10434,N_10413);
nand U10789 (N_10789,N_10594,N_10494);
nor U10790 (N_10790,N_10505,N_10535);
or U10791 (N_10791,N_10543,N_10587);
and U10792 (N_10792,N_10548,N_10597);
or U10793 (N_10793,N_10548,N_10588);
xor U10794 (N_10794,N_10549,N_10482);
and U10795 (N_10795,N_10480,N_10421);
xnor U10796 (N_10796,N_10533,N_10437);
nor U10797 (N_10797,N_10408,N_10578);
xor U10798 (N_10798,N_10464,N_10445);
or U10799 (N_10799,N_10557,N_10468);
nor U10800 (N_10800,N_10631,N_10750);
nor U10801 (N_10801,N_10774,N_10657);
nor U10802 (N_10802,N_10693,N_10606);
nand U10803 (N_10803,N_10744,N_10636);
nor U10804 (N_10804,N_10764,N_10681);
or U10805 (N_10805,N_10625,N_10609);
nor U10806 (N_10806,N_10620,N_10742);
xnor U10807 (N_10807,N_10730,N_10798);
nor U10808 (N_10808,N_10710,N_10683);
and U10809 (N_10809,N_10762,N_10753);
xnor U10810 (N_10810,N_10766,N_10747);
and U10811 (N_10811,N_10752,N_10617);
nor U10812 (N_10812,N_10732,N_10667);
xnor U10813 (N_10813,N_10734,N_10663);
or U10814 (N_10814,N_10677,N_10624);
or U10815 (N_10815,N_10756,N_10645);
or U10816 (N_10816,N_10647,N_10672);
or U10817 (N_10817,N_10669,N_10623);
xnor U10818 (N_10818,N_10605,N_10694);
nor U10819 (N_10819,N_10790,N_10745);
nor U10820 (N_10820,N_10695,N_10709);
nand U10821 (N_10821,N_10748,N_10687);
and U10822 (N_10822,N_10682,N_10662);
nor U10823 (N_10823,N_10629,N_10634);
or U10824 (N_10824,N_10674,N_10728);
and U10825 (N_10825,N_10630,N_10603);
or U10826 (N_10826,N_10782,N_10699);
nor U10827 (N_10827,N_10700,N_10754);
or U10828 (N_10828,N_10763,N_10627);
nand U10829 (N_10829,N_10776,N_10641);
and U10830 (N_10830,N_10684,N_10661);
nand U10831 (N_10831,N_10670,N_10615);
and U10832 (N_10832,N_10659,N_10707);
nor U10833 (N_10833,N_10619,N_10793);
or U10834 (N_10834,N_10722,N_10607);
nor U10835 (N_10835,N_10675,N_10765);
and U10836 (N_10836,N_10711,N_10777);
or U10837 (N_10837,N_10723,N_10779);
nor U10838 (N_10838,N_10795,N_10704);
and U10839 (N_10839,N_10621,N_10755);
xnor U10840 (N_10840,N_10655,N_10688);
xnor U10841 (N_10841,N_10622,N_10712);
nor U10842 (N_10842,N_10638,N_10775);
and U10843 (N_10843,N_10676,N_10643);
nor U10844 (N_10844,N_10686,N_10769);
nor U10845 (N_10845,N_10660,N_10656);
xnor U10846 (N_10846,N_10758,N_10757);
or U10847 (N_10847,N_10652,N_10665);
and U10848 (N_10848,N_10714,N_10613);
xnor U10849 (N_10849,N_10601,N_10759);
nor U10850 (N_10850,N_10720,N_10713);
nand U10851 (N_10851,N_10740,N_10706);
or U10852 (N_10852,N_10637,N_10649);
nor U10853 (N_10853,N_10760,N_10604);
or U10854 (N_10854,N_10773,N_10696);
nor U10855 (N_10855,N_10666,N_10668);
nor U10856 (N_10856,N_10761,N_10703);
nor U10857 (N_10857,N_10751,N_10736);
xnor U10858 (N_10858,N_10626,N_10780);
nor U10859 (N_10859,N_10708,N_10653);
nand U10860 (N_10860,N_10678,N_10727);
and U10861 (N_10861,N_10729,N_10794);
and U10862 (N_10862,N_10797,N_10616);
nor U10863 (N_10863,N_10610,N_10644);
nand U10864 (N_10864,N_10799,N_10746);
nor U10865 (N_10865,N_10721,N_10783);
or U10866 (N_10866,N_10770,N_10715);
nor U10867 (N_10867,N_10771,N_10691);
xnor U10868 (N_10868,N_10784,N_10791);
xnor U10869 (N_10869,N_10731,N_10718);
or U10870 (N_10870,N_10738,N_10664);
xor U10871 (N_10871,N_10679,N_10789);
or U10872 (N_10872,N_10726,N_10608);
and U10873 (N_10873,N_10646,N_10787);
xor U10874 (N_10874,N_10689,N_10739);
or U10875 (N_10875,N_10716,N_10697);
nand U10876 (N_10876,N_10781,N_10628);
nand U10877 (N_10877,N_10658,N_10772);
nand U10878 (N_10878,N_10671,N_10611);
nand U10879 (N_10879,N_10786,N_10648);
nand U10880 (N_10880,N_10767,N_10768);
nor U10881 (N_10881,N_10680,N_10701);
nor U10882 (N_10882,N_10642,N_10602);
xor U10883 (N_10883,N_10612,N_10685);
xor U10884 (N_10884,N_10654,N_10600);
nand U10885 (N_10885,N_10651,N_10735);
nor U10886 (N_10886,N_10673,N_10733);
nor U10887 (N_10887,N_10705,N_10698);
or U10888 (N_10888,N_10749,N_10724);
or U10889 (N_10889,N_10796,N_10719);
and U10890 (N_10890,N_10635,N_10717);
or U10891 (N_10891,N_10614,N_10785);
xnor U10892 (N_10892,N_10690,N_10702);
nand U10893 (N_10893,N_10640,N_10737);
or U10894 (N_10894,N_10741,N_10639);
xnor U10895 (N_10895,N_10725,N_10778);
xor U10896 (N_10896,N_10788,N_10692);
nor U10897 (N_10897,N_10632,N_10633);
xnor U10898 (N_10898,N_10618,N_10792);
nor U10899 (N_10899,N_10650,N_10743);
or U10900 (N_10900,N_10711,N_10638);
or U10901 (N_10901,N_10758,N_10729);
nand U10902 (N_10902,N_10657,N_10660);
and U10903 (N_10903,N_10671,N_10681);
xnor U10904 (N_10904,N_10727,N_10648);
xor U10905 (N_10905,N_10681,N_10697);
nor U10906 (N_10906,N_10719,N_10707);
nor U10907 (N_10907,N_10737,N_10703);
xor U10908 (N_10908,N_10699,N_10608);
nand U10909 (N_10909,N_10725,N_10728);
nor U10910 (N_10910,N_10776,N_10645);
nor U10911 (N_10911,N_10741,N_10616);
xnor U10912 (N_10912,N_10748,N_10798);
or U10913 (N_10913,N_10606,N_10668);
xor U10914 (N_10914,N_10603,N_10751);
nor U10915 (N_10915,N_10792,N_10738);
xnor U10916 (N_10916,N_10631,N_10768);
xnor U10917 (N_10917,N_10724,N_10612);
nand U10918 (N_10918,N_10718,N_10721);
nor U10919 (N_10919,N_10627,N_10774);
and U10920 (N_10920,N_10731,N_10724);
nor U10921 (N_10921,N_10781,N_10704);
nand U10922 (N_10922,N_10650,N_10766);
or U10923 (N_10923,N_10627,N_10672);
or U10924 (N_10924,N_10732,N_10609);
nand U10925 (N_10925,N_10761,N_10706);
or U10926 (N_10926,N_10620,N_10780);
nor U10927 (N_10927,N_10629,N_10727);
nand U10928 (N_10928,N_10736,N_10684);
xor U10929 (N_10929,N_10711,N_10738);
or U10930 (N_10930,N_10756,N_10782);
and U10931 (N_10931,N_10686,N_10757);
or U10932 (N_10932,N_10634,N_10697);
nor U10933 (N_10933,N_10727,N_10610);
nand U10934 (N_10934,N_10699,N_10610);
or U10935 (N_10935,N_10762,N_10632);
and U10936 (N_10936,N_10770,N_10686);
nand U10937 (N_10937,N_10661,N_10600);
or U10938 (N_10938,N_10671,N_10713);
nand U10939 (N_10939,N_10792,N_10703);
nand U10940 (N_10940,N_10689,N_10727);
and U10941 (N_10941,N_10776,N_10613);
or U10942 (N_10942,N_10682,N_10652);
xor U10943 (N_10943,N_10791,N_10638);
nor U10944 (N_10944,N_10655,N_10788);
nand U10945 (N_10945,N_10779,N_10681);
or U10946 (N_10946,N_10644,N_10769);
and U10947 (N_10947,N_10670,N_10643);
nand U10948 (N_10948,N_10622,N_10758);
and U10949 (N_10949,N_10799,N_10661);
and U10950 (N_10950,N_10649,N_10694);
nor U10951 (N_10951,N_10670,N_10618);
xnor U10952 (N_10952,N_10764,N_10747);
xor U10953 (N_10953,N_10671,N_10799);
nor U10954 (N_10954,N_10770,N_10718);
and U10955 (N_10955,N_10604,N_10639);
nand U10956 (N_10956,N_10636,N_10730);
nand U10957 (N_10957,N_10689,N_10604);
nor U10958 (N_10958,N_10649,N_10730);
and U10959 (N_10959,N_10617,N_10757);
xnor U10960 (N_10960,N_10605,N_10751);
or U10961 (N_10961,N_10650,N_10678);
nand U10962 (N_10962,N_10769,N_10704);
nor U10963 (N_10963,N_10616,N_10641);
xnor U10964 (N_10964,N_10638,N_10750);
or U10965 (N_10965,N_10685,N_10711);
or U10966 (N_10966,N_10673,N_10745);
and U10967 (N_10967,N_10619,N_10668);
or U10968 (N_10968,N_10695,N_10738);
nand U10969 (N_10969,N_10698,N_10605);
xnor U10970 (N_10970,N_10604,N_10654);
xnor U10971 (N_10971,N_10673,N_10619);
nand U10972 (N_10972,N_10662,N_10691);
xor U10973 (N_10973,N_10747,N_10608);
nand U10974 (N_10974,N_10618,N_10650);
xnor U10975 (N_10975,N_10667,N_10734);
nor U10976 (N_10976,N_10715,N_10768);
nor U10977 (N_10977,N_10743,N_10696);
xor U10978 (N_10978,N_10682,N_10766);
and U10979 (N_10979,N_10695,N_10799);
and U10980 (N_10980,N_10746,N_10665);
nand U10981 (N_10981,N_10670,N_10693);
nor U10982 (N_10982,N_10664,N_10621);
or U10983 (N_10983,N_10616,N_10744);
nand U10984 (N_10984,N_10737,N_10612);
nand U10985 (N_10985,N_10641,N_10762);
nand U10986 (N_10986,N_10674,N_10752);
nor U10987 (N_10987,N_10743,N_10683);
nand U10988 (N_10988,N_10772,N_10729);
xor U10989 (N_10989,N_10744,N_10686);
nor U10990 (N_10990,N_10635,N_10679);
nand U10991 (N_10991,N_10653,N_10665);
or U10992 (N_10992,N_10629,N_10769);
xnor U10993 (N_10993,N_10656,N_10732);
or U10994 (N_10994,N_10741,N_10721);
nand U10995 (N_10995,N_10714,N_10642);
xor U10996 (N_10996,N_10654,N_10638);
or U10997 (N_10997,N_10724,N_10615);
nor U10998 (N_10998,N_10655,N_10760);
xor U10999 (N_10999,N_10799,N_10688);
or U11000 (N_11000,N_10867,N_10838);
and U11001 (N_11001,N_10856,N_10925);
nand U11002 (N_11002,N_10929,N_10887);
or U11003 (N_11003,N_10843,N_10970);
nor U11004 (N_11004,N_10836,N_10889);
xnor U11005 (N_11005,N_10850,N_10927);
xnor U11006 (N_11006,N_10876,N_10910);
and U11007 (N_11007,N_10989,N_10840);
or U11008 (N_11008,N_10818,N_10950);
and U11009 (N_11009,N_10827,N_10875);
nand U11010 (N_11010,N_10922,N_10801);
or U11011 (N_11011,N_10808,N_10935);
xnor U11012 (N_11012,N_10860,N_10844);
and U11013 (N_11013,N_10940,N_10972);
or U11014 (N_11014,N_10878,N_10920);
or U11015 (N_11015,N_10893,N_10924);
xor U11016 (N_11016,N_10855,N_10820);
xor U11017 (N_11017,N_10899,N_10936);
nand U11018 (N_11018,N_10859,N_10825);
nand U11019 (N_11019,N_10909,N_10905);
and U11020 (N_11020,N_10819,N_10951);
nor U11021 (N_11021,N_10985,N_10993);
nor U11022 (N_11022,N_10853,N_10866);
nand U11023 (N_11023,N_10861,N_10946);
xor U11024 (N_11024,N_10968,N_10942);
or U11025 (N_11025,N_10991,N_10952);
nor U11026 (N_11026,N_10911,N_10813);
and U11027 (N_11027,N_10858,N_10872);
nor U11028 (N_11028,N_10892,N_10849);
nand U11029 (N_11029,N_10982,N_10891);
nand U11030 (N_11030,N_10996,N_10962);
or U11031 (N_11031,N_10978,N_10971);
and U11032 (N_11032,N_10919,N_10980);
and U11033 (N_11033,N_10945,N_10958);
nand U11034 (N_11034,N_10913,N_10999);
nand U11035 (N_11035,N_10981,N_10874);
nor U11036 (N_11036,N_10883,N_10830);
xor U11037 (N_11037,N_10894,N_10865);
nand U11038 (N_11038,N_10828,N_10937);
nand U11039 (N_11039,N_10966,N_10871);
nor U11040 (N_11040,N_10926,N_10977);
xnor U11041 (N_11041,N_10886,N_10955);
nand U11042 (N_11042,N_10862,N_10897);
or U11043 (N_11043,N_10906,N_10868);
xor U11044 (N_11044,N_10890,N_10988);
and U11045 (N_11045,N_10900,N_10973);
nand U11046 (N_11046,N_10880,N_10806);
xor U11047 (N_11047,N_10815,N_10960);
nor U11048 (N_11048,N_10907,N_10834);
or U11049 (N_11049,N_10804,N_10957);
or U11050 (N_11050,N_10963,N_10863);
nor U11051 (N_11051,N_10903,N_10976);
xor U11052 (N_11052,N_10944,N_10846);
and U11053 (N_11053,N_10814,N_10812);
and U11054 (N_11054,N_10984,N_10916);
and U11055 (N_11055,N_10854,N_10967);
xor U11056 (N_11056,N_10947,N_10847);
nor U11057 (N_11057,N_10933,N_10879);
or U11058 (N_11058,N_10896,N_10932);
nor U11059 (N_11059,N_10826,N_10983);
and U11060 (N_11060,N_10802,N_10829);
or U11061 (N_11061,N_10998,N_10914);
nor U11062 (N_11062,N_10917,N_10997);
nor U11063 (N_11063,N_10965,N_10833);
nand U11064 (N_11064,N_10881,N_10869);
nand U11065 (N_11065,N_10992,N_10832);
xor U11066 (N_11066,N_10994,N_10803);
xnor U11067 (N_11067,N_10824,N_10959);
or U11068 (N_11068,N_10987,N_10974);
xnor U11069 (N_11069,N_10823,N_10953);
and U11070 (N_11070,N_10928,N_10805);
or U11071 (N_11071,N_10954,N_10943);
xnor U11072 (N_11072,N_10822,N_10870);
xnor U11073 (N_11073,N_10885,N_10845);
xnor U11074 (N_11074,N_10915,N_10882);
nor U11075 (N_11075,N_10964,N_10904);
and U11076 (N_11076,N_10831,N_10857);
nand U11077 (N_11077,N_10923,N_10841);
nor U11078 (N_11078,N_10842,N_10908);
and U11079 (N_11079,N_10956,N_10851);
xnor U11080 (N_11080,N_10888,N_10817);
xnor U11081 (N_11081,N_10821,N_10934);
xnor U11082 (N_11082,N_10939,N_10941);
or U11083 (N_11083,N_10816,N_10912);
or U11084 (N_11084,N_10807,N_10895);
nor U11085 (N_11085,N_10877,N_10837);
xnor U11086 (N_11086,N_10961,N_10986);
xor U11087 (N_11087,N_10938,N_10931);
nand U11088 (N_11088,N_10930,N_10969);
nor U11089 (N_11089,N_10811,N_10948);
and U11090 (N_11090,N_10918,N_10800);
nand U11091 (N_11091,N_10848,N_10995);
and U11092 (N_11092,N_10901,N_10835);
nand U11093 (N_11093,N_10810,N_10902);
nor U11094 (N_11094,N_10809,N_10949);
nand U11095 (N_11095,N_10979,N_10864);
and U11096 (N_11096,N_10921,N_10884);
nand U11097 (N_11097,N_10852,N_10839);
or U11098 (N_11098,N_10873,N_10975);
nor U11099 (N_11099,N_10898,N_10990);
and U11100 (N_11100,N_10955,N_10986);
or U11101 (N_11101,N_10800,N_10891);
and U11102 (N_11102,N_10928,N_10848);
nand U11103 (N_11103,N_10912,N_10823);
xor U11104 (N_11104,N_10807,N_10900);
xor U11105 (N_11105,N_10819,N_10810);
xor U11106 (N_11106,N_10951,N_10816);
nand U11107 (N_11107,N_10849,N_10935);
xor U11108 (N_11108,N_10854,N_10905);
and U11109 (N_11109,N_10945,N_10877);
xnor U11110 (N_11110,N_10937,N_10935);
nor U11111 (N_11111,N_10897,N_10933);
nand U11112 (N_11112,N_10838,N_10969);
and U11113 (N_11113,N_10856,N_10941);
and U11114 (N_11114,N_10826,N_10995);
nor U11115 (N_11115,N_10949,N_10855);
and U11116 (N_11116,N_10943,N_10946);
xor U11117 (N_11117,N_10891,N_10907);
or U11118 (N_11118,N_10811,N_10937);
and U11119 (N_11119,N_10909,N_10881);
nor U11120 (N_11120,N_10814,N_10907);
and U11121 (N_11121,N_10833,N_10901);
nand U11122 (N_11122,N_10859,N_10866);
or U11123 (N_11123,N_10939,N_10803);
xnor U11124 (N_11124,N_10943,N_10992);
or U11125 (N_11125,N_10816,N_10967);
nand U11126 (N_11126,N_10870,N_10834);
or U11127 (N_11127,N_10960,N_10944);
or U11128 (N_11128,N_10964,N_10864);
and U11129 (N_11129,N_10833,N_10943);
nand U11130 (N_11130,N_10841,N_10823);
or U11131 (N_11131,N_10802,N_10877);
nor U11132 (N_11132,N_10890,N_10849);
or U11133 (N_11133,N_10885,N_10916);
and U11134 (N_11134,N_10864,N_10836);
nor U11135 (N_11135,N_10914,N_10990);
nor U11136 (N_11136,N_10906,N_10985);
or U11137 (N_11137,N_10880,N_10997);
and U11138 (N_11138,N_10835,N_10905);
nand U11139 (N_11139,N_10977,N_10802);
and U11140 (N_11140,N_10989,N_10918);
and U11141 (N_11141,N_10887,N_10921);
nand U11142 (N_11142,N_10856,N_10800);
xor U11143 (N_11143,N_10918,N_10893);
nand U11144 (N_11144,N_10873,N_10835);
nor U11145 (N_11145,N_10863,N_10938);
nor U11146 (N_11146,N_10828,N_10991);
or U11147 (N_11147,N_10836,N_10844);
xnor U11148 (N_11148,N_10886,N_10879);
and U11149 (N_11149,N_10890,N_10882);
nor U11150 (N_11150,N_10801,N_10860);
nand U11151 (N_11151,N_10912,N_10879);
nand U11152 (N_11152,N_10961,N_10892);
or U11153 (N_11153,N_10976,N_10871);
nand U11154 (N_11154,N_10821,N_10956);
or U11155 (N_11155,N_10986,N_10817);
nor U11156 (N_11156,N_10941,N_10921);
nand U11157 (N_11157,N_10903,N_10893);
and U11158 (N_11158,N_10905,N_10857);
nand U11159 (N_11159,N_10903,N_10945);
or U11160 (N_11160,N_10824,N_10969);
and U11161 (N_11161,N_10830,N_10938);
xor U11162 (N_11162,N_10870,N_10980);
and U11163 (N_11163,N_10996,N_10819);
xor U11164 (N_11164,N_10911,N_10828);
or U11165 (N_11165,N_10831,N_10897);
nand U11166 (N_11166,N_10999,N_10946);
and U11167 (N_11167,N_10836,N_10946);
nor U11168 (N_11168,N_10881,N_10888);
or U11169 (N_11169,N_10933,N_10952);
nor U11170 (N_11170,N_10890,N_10818);
and U11171 (N_11171,N_10809,N_10981);
xnor U11172 (N_11172,N_10880,N_10924);
xnor U11173 (N_11173,N_10899,N_10850);
nand U11174 (N_11174,N_10939,N_10814);
and U11175 (N_11175,N_10968,N_10977);
xor U11176 (N_11176,N_10850,N_10978);
and U11177 (N_11177,N_10815,N_10973);
nand U11178 (N_11178,N_10895,N_10864);
and U11179 (N_11179,N_10860,N_10969);
nor U11180 (N_11180,N_10805,N_10975);
nand U11181 (N_11181,N_10848,N_10973);
xor U11182 (N_11182,N_10928,N_10861);
nand U11183 (N_11183,N_10828,N_10869);
or U11184 (N_11184,N_10961,N_10957);
or U11185 (N_11185,N_10937,N_10874);
nor U11186 (N_11186,N_10935,N_10978);
and U11187 (N_11187,N_10952,N_10966);
xor U11188 (N_11188,N_10983,N_10858);
nor U11189 (N_11189,N_10894,N_10940);
nand U11190 (N_11190,N_10878,N_10998);
and U11191 (N_11191,N_10985,N_10806);
nor U11192 (N_11192,N_10882,N_10965);
nand U11193 (N_11193,N_10883,N_10942);
and U11194 (N_11194,N_10847,N_10936);
xor U11195 (N_11195,N_10959,N_10945);
and U11196 (N_11196,N_10872,N_10928);
and U11197 (N_11197,N_10831,N_10824);
or U11198 (N_11198,N_10898,N_10811);
or U11199 (N_11199,N_10895,N_10873);
nor U11200 (N_11200,N_11174,N_11115);
or U11201 (N_11201,N_11089,N_11167);
or U11202 (N_11202,N_11016,N_11077);
or U11203 (N_11203,N_11147,N_11145);
and U11204 (N_11204,N_11153,N_11197);
nor U11205 (N_11205,N_11086,N_11176);
xor U11206 (N_11206,N_11012,N_11002);
nand U11207 (N_11207,N_11046,N_11148);
nor U11208 (N_11208,N_11155,N_11004);
xnor U11209 (N_11209,N_11065,N_11068);
nand U11210 (N_11210,N_11047,N_11175);
nor U11211 (N_11211,N_11049,N_11194);
nand U11212 (N_11212,N_11029,N_11063);
nor U11213 (N_11213,N_11187,N_11157);
and U11214 (N_11214,N_11100,N_11191);
and U11215 (N_11215,N_11126,N_11052);
xor U11216 (N_11216,N_11195,N_11113);
or U11217 (N_11217,N_11005,N_11120);
xnor U11218 (N_11218,N_11097,N_11121);
xnor U11219 (N_11219,N_11081,N_11160);
nor U11220 (N_11220,N_11088,N_11026);
and U11221 (N_11221,N_11102,N_11050);
or U11222 (N_11222,N_11041,N_11098);
xor U11223 (N_11223,N_11107,N_11030);
and U11224 (N_11224,N_11158,N_11130);
and U11225 (N_11225,N_11165,N_11171);
nor U11226 (N_11226,N_11177,N_11183);
xnor U11227 (N_11227,N_11020,N_11122);
xor U11228 (N_11228,N_11142,N_11064);
and U11229 (N_11229,N_11062,N_11186);
and U11230 (N_11230,N_11132,N_11109);
nor U11231 (N_11231,N_11076,N_11179);
xnor U11232 (N_11232,N_11078,N_11092);
nor U11233 (N_11233,N_11090,N_11127);
nand U11234 (N_11234,N_11173,N_11161);
and U11235 (N_11235,N_11074,N_11119);
nand U11236 (N_11236,N_11034,N_11083);
nand U11237 (N_11237,N_11071,N_11116);
nand U11238 (N_11238,N_11022,N_11163);
and U11239 (N_11239,N_11110,N_11140);
nand U11240 (N_11240,N_11015,N_11018);
or U11241 (N_11241,N_11024,N_11061);
nor U11242 (N_11242,N_11133,N_11036);
nor U11243 (N_11243,N_11150,N_11079);
nand U11244 (N_11244,N_11131,N_11073);
nor U11245 (N_11245,N_11108,N_11139);
and U11246 (N_11246,N_11111,N_11181);
nand U11247 (N_11247,N_11105,N_11008);
nand U11248 (N_11248,N_11025,N_11045);
nand U11249 (N_11249,N_11058,N_11027);
xor U11250 (N_11250,N_11196,N_11067);
xnor U11251 (N_11251,N_11040,N_11048);
or U11252 (N_11252,N_11124,N_11137);
xor U11253 (N_11253,N_11159,N_11057);
and U11254 (N_11254,N_11136,N_11118);
and U11255 (N_11255,N_11072,N_11085);
nor U11256 (N_11256,N_11093,N_11006);
xnor U11257 (N_11257,N_11135,N_11128);
xor U11258 (N_11258,N_11070,N_11184);
nand U11259 (N_11259,N_11117,N_11189);
nand U11260 (N_11260,N_11129,N_11146);
nand U11261 (N_11261,N_11134,N_11055);
or U11262 (N_11262,N_11039,N_11023);
nand U11263 (N_11263,N_11170,N_11031);
nand U11264 (N_11264,N_11001,N_11101);
and U11265 (N_11265,N_11185,N_11180);
nand U11266 (N_11266,N_11125,N_11141);
nand U11267 (N_11267,N_11028,N_11192);
or U11268 (N_11268,N_11014,N_11051);
or U11269 (N_11269,N_11053,N_11190);
and U11270 (N_11270,N_11042,N_11151);
nand U11271 (N_11271,N_11094,N_11037);
or U11272 (N_11272,N_11099,N_11054);
nor U11273 (N_11273,N_11080,N_11075);
nor U11274 (N_11274,N_11096,N_11000);
xnor U11275 (N_11275,N_11017,N_11019);
nand U11276 (N_11276,N_11033,N_11084);
nor U11277 (N_11277,N_11114,N_11172);
nand U11278 (N_11278,N_11193,N_11103);
and U11279 (N_11279,N_11168,N_11009);
and U11280 (N_11280,N_11007,N_11152);
or U11281 (N_11281,N_11199,N_11038);
or U11282 (N_11282,N_11082,N_11156);
or U11283 (N_11283,N_11011,N_11044);
nand U11284 (N_11284,N_11091,N_11138);
nand U11285 (N_11285,N_11149,N_11169);
or U11286 (N_11286,N_11104,N_11154);
or U11287 (N_11287,N_11164,N_11043);
xor U11288 (N_11288,N_11013,N_11188);
xnor U11289 (N_11289,N_11144,N_11123);
xor U11290 (N_11290,N_11032,N_11143);
and U11291 (N_11291,N_11021,N_11095);
nor U11292 (N_11292,N_11059,N_11178);
or U11293 (N_11293,N_11003,N_11056);
nand U11294 (N_11294,N_11198,N_11069);
xnor U11295 (N_11295,N_11010,N_11162);
and U11296 (N_11296,N_11106,N_11035);
or U11297 (N_11297,N_11060,N_11066);
or U11298 (N_11298,N_11087,N_11166);
nor U11299 (N_11299,N_11112,N_11182);
or U11300 (N_11300,N_11057,N_11042);
nand U11301 (N_11301,N_11029,N_11182);
or U11302 (N_11302,N_11158,N_11095);
xor U11303 (N_11303,N_11019,N_11035);
and U11304 (N_11304,N_11071,N_11166);
xor U11305 (N_11305,N_11130,N_11109);
nor U11306 (N_11306,N_11071,N_11019);
and U11307 (N_11307,N_11074,N_11027);
or U11308 (N_11308,N_11014,N_11030);
or U11309 (N_11309,N_11007,N_11039);
xor U11310 (N_11310,N_11078,N_11166);
nor U11311 (N_11311,N_11179,N_11101);
or U11312 (N_11312,N_11078,N_11069);
nand U11313 (N_11313,N_11176,N_11155);
or U11314 (N_11314,N_11095,N_11068);
xnor U11315 (N_11315,N_11091,N_11152);
nor U11316 (N_11316,N_11126,N_11086);
and U11317 (N_11317,N_11153,N_11168);
nor U11318 (N_11318,N_11048,N_11160);
and U11319 (N_11319,N_11051,N_11016);
xnor U11320 (N_11320,N_11168,N_11074);
nor U11321 (N_11321,N_11153,N_11172);
nor U11322 (N_11322,N_11122,N_11109);
nor U11323 (N_11323,N_11095,N_11034);
nor U11324 (N_11324,N_11006,N_11146);
nand U11325 (N_11325,N_11152,N_11183);
nor U11326 (N_11326,N_11087,N_11093);
and U11327 (N_11327,N_11052,N_11060);
and U11328 (N_11328,N_11123,N_11014);
and U11329 (N_11329,N_11177,N_11165);
or U11330 (N_11330,N_11049,N_11155);
xor U11331 (N_11331,N_11007,N_11022);
xor U11332 (N_11332,N_11017,N_11193);
nor U11333 (N_11333,N_11125,N_11028);
and U11334 (N_11334,N_11146,N_11115);
or U11335 (N_11335,N_11077,N_11179);
and U11336 (N_11336,N_11023,N_11134);
and U11337 (N_11337,N_11063,N_11051);
xnor U11338 (N_11338,N_11174,N_11134);
nor U11339 (N_11339,N_11126,N_11056);
or U11340 (N_11340,N_11095,N_11129);
nor U11341 (N_11341,N_11190,N_11027);
and U11342 (N_11342,N_11179,N_11072);
or U11343 (N_11343,N_11094,N_11011);
and U11344 (N_11344,N_11041,N_11103);
or U11345 (N_11345,N_11055,N_11161);
nor U11346 (N_11346,N_11131,N_11093);
xor U11347 (N_11347,N_11071,N_11014);
nor U11348 (N_11348,N_11110,N_11133);
and U11349 (N_11349,N_11037,N_11060);
or U11350 (N_11350,N_11093,N_11180);
or U11351 (N_11351,N_11016,N_11140);
nand U11352 (N_11352,N_11001,N_11181);
nand U11353 (N_11353,N_11002,N_11056);
xor U11354 (N_11354,N_11120,N_11087);
xor U11355 (N_11355,N_11176,N_11081);
and U11356 (N_11356,N_11073,N_11151);
xnor U11357 (N_11357,N_11127,N_11185);
and U11358 (N_11358,N_11091,N_11177);
and U11359 (N_11359,N_11127,N_11084);
and U11360 (N_11360,N_11119,N_11115);
and U11361 (N_11361,N_11005,N_11164);
and U11362 (N_11362,N_11059,N_11189);
nor U11363 (N_11363,N_11056,N_11195);
xor U11364 (N_11364,N_11042,N_11030);
xnor U11365 (N_11365,N_11081,N_11111);
xnor U11366 (N_11366,N_11176,N_11078);
or U11367 (N_11367,N_11066,N_11169);
xnor U11368 (N_11368,N_11014,N_11050);
nand U11369 (N_11369,N_11115,N_11074);
nand U11370 (N_11370,N_11140,N_11080);
nor U11371 (N_11371,N_11076,N_11117);
xnor U11372 (N_11372,N_11082,N_11137);
and U11373 (N_11373,N_11159,N_11155);
and U11374 (N_11374,N_11155,N_11051);
xnor U11375 (N_11375,N_11164,N_11056);
nor U11376 (N_11376,N_11031,N_11065);
and U11377 (N_11377,N_11046,N_11169);
nor U11378 (N_11378,N_11177,N_11082);
xnor U11379 (N_11379,N_11067,N_11197);
nor U11380 (N_11380,N_11042,N_11058);
and U11381 (N_11381,N_11161,N_11127);
nor U11382 (N_11382,N_11144,N_11163);
or U11383 (N_11383,N_11116,N_11006);
nor U11384 (N_11384,N_11178,N_11099);
nand U11385 (N_11385,N_11194,N_11178);
or U11386 (N_11386,N_11075,N_11079);
and U11387 (N_11387,N_11198,N_11163);
xnor U11388 (N_11388,N_11089,N_11134);
or U11389 (N_11389,N_11161,N_11175);
or U11390 (N_11390,N_11088,N_11103);
nand U11391 (N_11391,N_11175,N_11162);
xnor U11392 (N_11392,N_11154,N_11184);
nor U11393 (N_11393,N_11033,N_11175);
xor U11394 (N_11394,N_11060,N_11047);
xor U11395 (N_11395,N_11063,N_11044);
and U11396 (N_11396,N_11107,N_11196);
and U11397 (N_11397,N_11169,N_11157);
nor U11398 (N_11398,N_11002,N_11118);
nor U11399 (N_11399,N_11021,N_11134);
or U11400 (N_11400,N_11299,N_11337);
and U11401 (N_11401,N_11227,N_11201);
and U11402 (N_11402,N_11333,N_11334);
xor U11403 (N_11403,N_11292,N_11336);
nor U11404 (N_11404,N_11380,N_11236);
nand U11405 (N_11405,N_11377,N_11341);
and U11406 (N_11406,N_11396,N_11259);
nand U11407 (N_11407,N_11237,N_11373);
nor U11408 (N_11408,N_11247,N_11260);
xor U11409 (N_11409,N_11381,N_11244);
nor U11410 (N_11410,N_11270,N_11379);
xnor U11411 (N_11411,N_11399,N_11367);
or U11412 (N_11412,N_11328,N_11343);
nor U11413 (N_11413,N_11229,N_11219);
or U11414 (N_11414,N_11209,N_11254);
nand U11415 (N_11415,N_11382,N_11233);
nand U11416 (N_11416,N_11262,N_11305);
or U11417 (N_11417,N_11307,N_11295);
nor U11418 (N_11418,N_11222,N_11374);
nor U11419 (N_11419,N_11365,N_11360);
and U11420 (N_11420,N_11204,N_11293);
nor U11421 (N_11421,N_11207,N_11356);
and U11422 (N_11422,N_11398,N_11226);
nand U11423 (N_11423,N_11287,N_11298);
or U11424 (N_11424,N_11281,N_11251);
or U11425 (N_11425,N_11368,N_11327);
xnor U11426 (N_11426,N_11267,N_11339);
xor U11427 (N_11427,N_11364,N_11257);
or U11428 (N_11428,N_11317,N_11218);
xor U11429 (N_11429,N_11275,N_11375);
xnor U11430 (N_11430,N_11344,N_11216);
nand U11431 (N_11431,N_11350,N_11280);
nor U11432 (N_11432,N_11303,N_11314);
xor U11433 (N_11433,N_11323,N_11348);
and U11434 (N_11434,N_11369,N_11345);
nor U11435 (N_11435,N_11290,N_11351);
nand U11436 (N_11436,N_11325,N_11383);
and U11437 (N_11437,N_11385,N_11200);
xnor U11438 (N_11438,N_11234,N_11363);
or U11439 (N_11439,N_11310,N_11318);
and U11440 (N_11440,N_11221,N_11230);
and U11441 (N_11441,N_11372,N_11215);
nor U11442 (N_11442,N_11352,N_11296);
xnor U11443 (N_11443,N_11249,N_11346);
xor U11444 (N_11444,N_11300,N_11258);
and U11445 (N_11445,N_11246,N_11277);
xor U11446 (N_11446,N_11313,N_11302);
nand U11447 (N_11447,N_11212,N_11265);
xnor U11448 (N_11448,N_11252,N_11268);
nor U11449 (N_11449,N_11248,N_11271);
and U11450 (N_11450,N_11205,N_11269);
nand U11451 (N_11451,N_11357,N_11322);
or U11452 (N_11452,N_11340,N_11211);
and U11453 (N_11453,N_11255,N_11387);
or U11454 (N_11454,N_11371,N_11304);
or U11455 (N_11455,N_11203,N_11206);
nand U11456 (N_11456,N_11208,N_11388);
xnor U11457 (N_11457,N_11243,N_11370);
nor U11458 (N_11458,N_11354,N_11319);
xor U11459 (N_11459,N_11253,N_11395);
nor U11460 (N_11460,N_11291,N_11288);
nand U11461 (N_11461,N_11332,N_11239);
and U11462 (N_11462,N_11272,N_11225);
and U11463 (N_11463,N_11338,N_11263);
and U11464 (N_11464,N_11342,N_11311);
or U11465 (N_11465,N_11347,N_11312);
or U11466 (N_11466,N_11231,N_11355);
nor U11467 (N_11467,N_11389,N_11235);
or U11468 (N_11468,N_11286,N_11316);
and U11469 (N_11469,N_11261,N_11294);
nand U11470 (N_11470,N_11210,N_11386);
xnor U11471 (N_11471,N_11220,N_11264);
xor U11472 (N_11472,N_11378,N_11279);
or U11473 (N_11473,N_11393,N_11326);
and U11474 (N_11474,N_11362,N_11306);
xnor U11475 (N_11475,N_11394,N_11320);
and U11476 (N_11476,N_11353,N_11232);
nor U11477 (N_11477,N_11289,N_11217);
nand U11478 (N_11478,N_11242,N_11321);
or U11479 (N_11479,N_11285,N_11329);
or U11480 (N_11480,N_11276,N_11390);
and U11481 (N_11481,N_11241,N_11213);
or U11482 (N_11482,N_11361,N_11392);
nor U11483 (N_11483,N_11278,N_11349);
and U11484 (N_11484,N_11250,N_11282);
nand U11485 (N_11485,N_11245,N_11359);
or U11486 (N_11486,N_11274,N_11330);
nand U11487 (N_11487,N_11391,N_11324);
and U11488 (N_11488,N_11228,N_11284);
xor U11489 (N_11489,N_11223,N_11308);
nand U11490 (N_11490,N_11240,N_11224);
xor U11491 (N_11491,N_11301,N_11335);
nand U11492 (N_11492,N_11358,N_11331);
xnor U11493 (N_11493,N_11376,N_11297);
nor U11494 (N_11494,N_11309,N_11256);
xor U11495 (N_11495,N_11202,N_11315);
xnor U11496 (N_11496,N_11273,N_11238);
xor U11497 (N_11497,N_11366,N_11283);
or U11498 (N_11498,N_11384,N_11397);
or U11499 (N_11499,N_11266,N_11214);
nor U11500 (N_11500,N_11306,N_11205);
xor U11501 (N_11501,N_11378,N_11301);
xnor U11502 (N_11502,N_11358,N_11320);
and U11503 (N_11503,N_11235,N_11219);
and U11504 (N_11504,N_11318,N_11266);
nand U11505 (N_11505,N_11253,N_11203);
nand U11506 (N_11506,N_11317,N_11207);
nor U11507 (N_11507,N_11354,N_11259);
nor U11508 (N_11508,N_11375,N_11246);
nand U11509 (N_11509,N_11394,N_11369);
nor U11510 (N_11510,N_11222,N_11236);
and U11511 (N_11511,N_11299,N_11320);
or U11512 (N_11512,N_11201,N_11390);
and U11513 (N_11513,N_11252,N_11303);
and U11514 (N_11514,N_11291,N_11262);
nand U11515 (N_11515,N_11210,N_11296);
nor U11516 (N_11516,N_11219,N_11398);
nand U11517 (N_11517,N_11384,N_11357);
nand U11518 (N_11518,N_11249,N_11211);
xor U11519 (N_11519,N_11295,N_11277);
and U11520 (N_11520,N_11213,N_11358);
or U11521 (N_11521,N_11379,N_11263);
xor U11522 (N_11522,N_11284,N_11232);
and U11523 (N_11523,N_11397,N_11399);
or U11524 (N_11524,N_11301,N_11247);
or U11525 (N_11525,N_11303,N_11276);
or U11526 (N_11526,N_11252,N_11305);
nor U11527 (N_11527,N_11343,N_11210);
nor U11528 (N_11528,N_11204,N_11358);
xnor U11529 (N_11529,N_11255,N_11374);
and U11530 (N_11530,N_11237,N_11239);
or U11531 (N_11531,N_11280,N_11249);
nor U11532 (N_11532,N_11317,N_11372);
or U11533 (N_11533,N_11351,N_11207);
and U11534 (N_11534,N_11385,N_11271);
and U11535 (N_11535,N_11259,N_11324);
xnor U11536 (N_11536,N_11358,N_11282);
xor U11537 (N_11537,N_11295,N_11258);
or U11538 (N_11538,N_11389,N_11338);
and U11539 (N_11539,N_11225,N_11277);
and U11540 (N_11540,N_11233,N_11214);
and U11541 (N_11541,N_11346,N_11340);
and U11542 (N_11542,N_11297,N_11205);
nand U11543 (N_11543,N_11254,N_11398);
nand U11544 (N_11544,N_11373,N_11239);
nor U11545 (N_11545,N_11212,N_11226);
nand U11546 (N_11546,N_11317,N_11391);
nor U11547 (N_11547,N_11244,N_11209);
nand U11548 (N_11548,N_11202,N_11301);
nand U11549 (N_11549,N_11272,N_11320);
and U11550 (N_11550,N_11245,N_11211);
and U11551 (N_11551,N_11276,N_11353);
nand U11552 (N_11552,N_11284,N_11283);
xnor U11553 (N_11553,N_11360,N_11246);
nand U11554 (N_11554,N_11355,N_11391);
nor U11555 (N_11555,N_11296,N_11388);
or U11556 (N_11556,N_11377,N_11271);
nor U11557 (N_11557,N_11356,N_11393);
xnor U11558 (N_11558,N_11259,N_11245);
nand U11559 (N_11559,N_11359,N_11356);
and U11560 (N_11560,N_11201,N_11399);
xor U11561 (N_11561,N_11360,N_11201);
or U11562 (N_11562,N_11261,N_11325);
nand U11563 (N_11563,N_11280,N_11200);
nor U11564 (N_11564,N_11218,N_11341);
nand U11565 (N_11565,N_11336,N_11335);
nor U11566 (N_11566,N_11223,N_11341);
and U11567 (N_11567,N_11361,N_11280);
xor U11568 (N_11568,N_11261,N_11302);
nor U11569 (N_11569,N_11273,N_11302);
or U11570 (N_11570,N_11298,N_11361);
nor U11571 (N_11571,N_11366,N_11209);
or U11572 (N_11572,N_11293,N_11349);
nor U11573 (N_11573,N_11270,N_11279);
xor U11574 (N_11574,N_11204,N_11286);
and U11575 (N_11575,N_11385,N_11222);
nand U11576 (N_11576,N_11364,N_11312);
and U11577 (N_11577,N_11290,N_11354);
nor U11578 (N_11578,N_11334,N_11268);
nand U11579 (N_11579,N_11280,N_11291);
xnor U11580 (N_11580,N_11295,N_11347);
nand U11581 (N_11581,N_11398,N_11224);
nand U11582 (N_11582,N_11340,N_11359);
and U11583 (N_11583,N_11359,N_11391);
nand U11584 (N_11584,N_11349,N_11273);
nor U11585 (N_11585,N_11351,N_11324);
or U11586 (N_11586,N_11302,N_11244);
or U11587 (N_11587,N_11247,N_11241);
and U11588 (N_11588,N_11208,N_11242);
and U11589 (N_11589,N_11250,N_11225);
xnor U11590 (N_11590,N_11395,N_11375);
or U11591 (N_11591,N_11260,N_11233);
or U11592 (N_11592,N_11305,N_11219);
xor U11593 (N_11593,N_11200,N_11270);
and U11594 (N_11594,N_11203,N_11321);
and U11595 (N_11595,N_11365,N_11255);
and U11596 (N_11596,N_11328,N_11394);
and U11597 (N_11597,N_11228,N_11336);
xor U11598 (N_11598,N_11242,N_11361);
nand U11599 (N_11599,N_11360,N_11250);
and U11600 (N_11600,N_11517,N_11475);
xnor U11601 (N_11601,N_11546,N_11556);
and U11602 (N_11602,N_11555,N_11433);
and U11603 (N_11603,N_11508,N_11470);
and U11604 (N_11604,N_11516,N_11495);
nand U11605 (N_11605,N_11551,N_11493);
xor U11606 (N_11606,N_11531,N_11590);
and U11607 (N_11607,N_11409,N_11592);
xnor U11608 (N_11608,N_11498,N_11418);
or U11609 (N_11609,N_11423,N_11539);
nor U11610 (N_11610,N_11404,N_11532);
nand U11611 (N_11611,N_11594,N_11442);
xnor U11612 (N_11612,N_11459,N_11501);
nand U11613 (N_11613,N_11510,N_11488);
xnor U11614 (N_11614,N_11579,N_11564);
and U11615 (N_11615,N_11439,N_11525);
nor U11616 (N_11616,N_11481,N_11467);
nand U11617 (N_11617,N_11521,N_11453);
nand U11618 (N_11618,N_11548,N_11573);
nor U11619 (N_11619,N_11407,N_11430);
or U11620 (N_11620,N_11526,N_11458);
xor U11621 (N_11621,N_11503,N_11499);
and U11622 (N_11622,N_11565,N_11588);
or U11623 (N_11623,N_11447,N_11455);
and U11624 (N_11624,N_11586,N_11544);
xor U11625 (N_11625,N_11450,N_11511);
or U11626 (N_11626,N_11401,N_11572);
and U11627 (N_11627,N_11578,N_11554);
and U11628 (N_11628,N_11575,N_11449);
nand U11629 (N_11629,N_11529,N_11599);
nor U11630 (N_11630,N_11413,N_11483);
or U11631 (N_11631,N_11568,N_11491);
and U11632 (N_11632,N_11584,N_11534);
nor U11633 (N_11633,N_11474,N_11598);
and U11634 (N_11634,N_11591,N_11436);
or U11635 (N_11635,N_11435,N_11597);
or U11636 (N_11636,N_11497,N_11445);
or U11637 (N_11637,N_11570,N_11490);
and U11638 (N_11638,N_11560,N_11500);
or U11639 (N_11639,N_11464,N_11469);
xor U11640 (N_11640,N_11402,N_11550);
and U11641 (N_11641,N_11567,N_11563);
or U11642 (N_11642,N_11415,N_11509);
nor U11643 (N_11643,N_11535,N_11471);
or U11644 (N_11644,N_11593,N_11460);
xor U11645 (N_11645,N_11577,N_11443);
xnor U11646 (N_11646,N_11446,N_11482);
xor U11647 (N_11647,N_11477,N_11537);
nor U11648 (N_11648,N_11422,N_11561);
xnor U11649 (N_11649,N_11486,N_11566);
and U11650 (N_11650,N_11496,N_11533);
xor U11651 (N_11651,N_11519,N_11411);
or U11652 (N_11652,N_11466,N_11538);
xnor U11653 (N_11653,N_11494,N_11473);
nand U11654 (N_11654,N_11476,N_11426);
nor U11655 (N_11655,N_11456,N_11434);
or U11656 (N_11656,N_11558,N_11523);
nand U11657 (N_11657,N_11425,N_11513);
nand U11658 (N_11658,N_11540,N_11595);
or U11659 (N_11659,N_11541,N_11427);
nor U11660 (N_11660,N_11428,N_11549);
and U11661 (N_11661,N_11569,N_11574);
xnor U11662 (N_11662,N_11408,N_11462);
and U11663 (N_11663,N_11557,N_11457);
or U11664 (N_11664,N_11547,N_11429);
or U11665 (N_11665,N_11410,N_11441);
or U11666 (N_11666,N_11484,N_11504);
or U11667 (N_11667,N_11530,N_11472);
nand U11668 (N_11668,N_11528,N_11485);
nor U11669 (N_11669,N_11465,N_11412);
nand U11670 (N_11670,N_11507,N_11543);
nor U11671 (N_11671,N_11542,N_11559);
xor U11672 (N_11672,N_11438,N_11502);
or U11673 (N_11673,N_11562,N_11479);
nor U11674 (N_11674,N_11587,N_11431);
nand U11675 (N_11675,N_11416,N_11581);
nor U11676 (N_11676,N_11478,N_11576);
nor U11677 (N_11677,N_11520,N_11440);
or U11678 (N_11678,N_11421,N_11536);
or U11679 (N_11679,N_11403,N_11506);
nor U11680 (N_11680,N_11454,N_11489);
or U11681 (N_11681,N_11463,N_11524);
xnor U11682 (N_11682,N_11444,N_11596);
and U11683 (N_11683,N_11571,N_11514);
xor U11684 (N_11684,N_11589,N_11405);
or U11685 (N_11685,N_11552,N_11518);
xnor U11686 (N_11686,N_11492,N_11505);
nor U11687 (N_11687,N_11553,N_11582);
and U11688 (N_11688,N_11451,N_11448);
xor U11689 (N_11689,N_11522,N_11580);
xor U11690 (N_11690,N_11515,N_11468);
xor U11691 (N_11691,N_11400,N_11583);
or U11692 (N_11692,N_11487,N_11545);
or U11693 (N_11693,N_11432,N_11461);
nor U11694 (N_11694,N_11414,N_11480);
nand U11695 (N_11695,N_11417,N_11452);
and U11696 (N_11696,N_11424,N_11527);
nor U11697 (N_11697,N_11585,N_11437);
xor U11698 (N_11698,N_11512,N_11419);
xor U11699 (N_11699,N_11420,N_11406);
and U11700 (N_11700,N_11493,N_11452);
nor U11701 (N_11701,N_11584,N_11501);
nand U11702 (N_11702,N_11521,N_11470);
and U11703 (N_11703,N_11596,N_11541);
nand U11704 (N_11704,N_11548,N_11524);
or U11705 (N_11705,N_11400,N_11447);
nand U11706 (N_11706,N_11535,N_11554);
nor U11707 (N_11707,N_11560,N_11438);
nor U11708 (N_11708,N_11553,N_11460);
xnor U11709 (N_11709,N_11400,N_11540);
and U11710 (N_11710,N_11438,N_11450);
or U11711 (N_11711,N_11579,N_11408);
nand U11712 (N_11712,N_11560,N_11495);
nor U11713 (N_11713,N_11447,N_11468);
nand U11714 (N_11714,N_11452,N_11499);
nor U11715 (N_11715,N_11459,N_11487);
or U11716 (N_11716,N_11573,N_11577);
or U11717 (N_11717,N_11598,N_11478);
and U11718 (N_11718,N_11497,N_11482);
xnor U11719 (N_11719,N_11568,N_11558);
or U11720 (N_11720,N_11563,N_11424);
nor U11721 (N_11721,N_11464,N_11579);
or U11722 (N_11722,N_11464,N_11509);
nand U11723 (N_11723,N_11506,N_11400);
xnor U11724 (N_11724,N_11439,N_11519);
xor U11725 (N_11725,N_11521,N_11577);
or U11726 (N_11726,N_11512,N_11544);
xor U11727 (N_11727,N_11523,N_11550);
nand U11728 (N_11728,N_11491,N_11412);
or U11729 (N_11729,N_11488,N_11405);
xor U11730 (N_11730,N_11593,N_11524);
nand U11731 (N_11731,N_11586,N_11430);
or U11732 (N_11732,N_11447,N_11544);
or U11733 (N_11733,N_11489,N_11451);
or U11734 (N_11734,N_11416,N_11559);
or U11735 (N_11735,N_11581,N_11461);
nor U11736 (N_11736,N_11412,N_11476);
nor U11737 (N_11737,N_11466,N_11571);
or U11738 (N_11738,N_11535,N_11457);
nand U11739 (N_11739,N_11591,N_11578);
nor U11740 (N_11740,N_11498,N_11568);
nand U11741 (N_11741,N_11426,N_11513);
nand U11742 (N_11742,N_11587,N_11477);
xor U11743 (N_11743,N_11420,N_11513);
or U11744 (N_11744,N_11547,N_11422);
and U11745 (N_11745,N_11547,N_11540);
xnor U11746 (N_11746,N_11508,N_11462);
and U11747 (N_11747,N_11572,N_11435);
nor U11748 (N_11748,N_11594,N_11491);
or U11749 (N_11749,N_11439,N_11477);
and U11750 (N_11750,N_11421,N_11434);
nand U11751 (N_11751,N_11568,N_11419);
xnor U11752 (N_11752,N_11468,N_11525);
nor U11753 (N_11753,N_11446,N_11503);
or U11754 (N_11754,N_11430,N_11517);
and U11755 (N_11755,N_11469,N_11590);
and U11756 (N_11756,N_11422,N_11420);
xor U11757 (N_11757,N_11589,N_11436);
and U11758 (N_11758,N_11469,N_11568);
nor U11759 (N_11759,N_11504,N_11528);
and U11760 (N_11760,N_11501,N_11426);
xor U11761 (N_11761,N_11536,N_11541);
xor U11762 (N_11762,N_11505,N_11494);
or U11763 (N_11763,N_11507,N_11489);
and U11764 (N_11764,N_11564,N_11410);
nor U11765 (N_11765,N_11403,N_11538);
nor U11766 (N_11766,N_11577,N_11520);
or U11767 (N_11767,N_11486,N_11405);
xor U11768 (N_11768,N_11413,N_11597);
nor U11769 (N_11769,N_11439,N_11475);
and U11770 (N_11770,N_11510,N_11588);
nand U11771 (N_11771,N_11412,N_11475);
or U11772 (N_11772,N_11544,N_11416);
nor U11773 (N_11773,N_11566,N_11437);
or U11774 (N_11774,N_11473,N_11593);
nand U11775 (N_11775,N_11460,N_11569);
nand U11776 (N_11776,N_11513,N_11414);
nand U11777 (N_11777,N_11463,N_11548);
xnor U11778 (N_11778,N_11552,N_11563);
nand U11779 (N_11779,N_11503,N_11555);
xor U11780 (N_11780,N_11451,N_11513);
nand U11781 (N_11781,N_11405,N_11540);
or U11782 (N_11782,N_11532,N_11570);
and U11783 (N_11783,N_11411,N_11548);
xor U11784 (N_11784,N_11401,N_11545);
or U11785 (N_11785,N_11509,N_11590);
and U11786 (N_11786,N_11477,N_11517);
xnor U11787 (N_11787,N_11536,N_11450);
or U11788 (N_11788,N_11564,N_11530);
nor U11789 (N_11789,N_11411,N_11521);
nand U11790 (N_11790,N_11402,N_11422);
or U11791 (N_11791,N_11563,N_11586);
xor U11792 (N_11792,N_11456,N_11513);
or U11793 (N_11793,N_11544,N_11497);
xor U11794 (N_11794,N_11400,N_11451);
or U11795 (N_11795,N_11502,N_11520);
nand U11796 (N_11796,N_11500,N_11483);
and U11797 (N_11797,N_11565,N_11594);
nor U11798 (N_11798,N_11520,N_11459);
and U11799 (N_11799,N_11486,N_11449);
xor U11800 (N_11800,N_11621,N_11602);
and U11801 (N_11801,N_11610,N_11798);
nor U11802 (N_11802,N_11634,N_11763);
and U11803 (N_11803,N_11734,N_11785);
or U11804 (N_11804,N_11764,N_11788);
xnor U11805 (N_11805,N_11779,N_11636);
xnor U11806 (N_11806,N_11727,N_11666);
or U11807 (N_11807,N_11743,N_11725);
nand U11808 (N_11808,N_11781,N_11792);
xnor U11809 (N_11809,N_11657,N_11627);
or U11810 (N_11810,N_11651,N_11638);
nand U11811 (N_11811,N_11662,N_11643);
xor U11812 (N_11812,N_11770,N_11726);
nor U11813 (N_11813,N_11695,N_11758);
xnor U11814 (N_11814,N_11768,N_11609);
nand U11815 (N_11815,N_11612,N_11647);
or U11816 (N_11816,N_11654,N_11720);
nor U11817 (N_11817,N_11697,N_11639);
nand U11818 (N_11818,N_11687,N_11671);
nand U11819 (N_11819,N_11692,N_11616);
nor U11820 (N_11820,N_11652,N_11756);
xnor U11821 (N_11821,N_11633,N_11776);
and U11822 (N_11822,N_11696,N_11645);
nor U11823 (N_11823,N_11767,N_11759);
nand U11824 (N_11824,N_11716,N_11748);
nand U11825 (N_11825,N_11678,N_11786);
and U11826 (N_11826,N_11630,N_11656);
nand U11827 (N_11827,N_11714,N_11685);
or U11828 (N_11828,N_11746,N_11774);
nor U11829 (N_11829,N_11607,N_11659);
xor U11830 (N_11830,N_11673,N_11670);
and U11831 (N_11831,N_11637,N_11700);
and U11832 (N_11832,N_11782,N_11740);
and U11833 (N_11833,N_11711,N_11628);
xor U11834 (N_11834,N_11623,N_11729);
nor U11835 (N_11835,N_11731,N_11603);
nor U11836 (N_11836,N_11622,N_11618);
nor U11837 (N_11837,N_11613,N_11706);
xnor U11838 (N_11838,N_11699,N_11715);
or U11839 (N_11839,N_11723,N_11669);
nor U11840 (N_11840,N_11744,N_11762);
xor U11841 (N_11841,N_11619,N_11739);
nand U11842 (N_11842,N_11611,N_11676);
nor U11843 (N_11843,N_11795,N_11680);
nor U11844 (N_11844,N_11772,N_11717);
nor U11845 (N_11845,N_11661,N_11705);
and U11846 (N_11846,N_11753,N_11644);
and U11847 (N_11847,N_11665,N_11766);
and U11848 (N_11848,N_11732,N_11682);
or U11849 (N_11849,N_11642,N_11690);
nor U11850 (N_11850,N_11784,N_11658);
nor U11851 (N_11851,N_11605,N_11641);
and U11852 (N_11852,N_11624,N_11655);
or U11853 (N_11853,N_11601,N_11640);
nor U11854 (N_11854,N_11718,N_11600);
or U11855 (N_11855,N_11620,N_11778);
or U11856 (N_11856,N_11684,N_11672);
nor U11857 (N_11857,N_11686,N_11736);
nand U11858 (N_11858,N_11789,N_11797);
nand U11859 (N_11859,N_11708,N_11660);
nor U11860 (N_11860,N_11614,N_11701);
nand U11861 (N_11861,N_11664,N_11649);
nor U11862 (N_11862,N_11667,N_11787);
nor U11863 (N_11863,N_11741,N_11760);
xnor U11864 (N_11864,N_11750,N_11689);
or U11865 (N_11865,N_11745,N_11653);
or U11866 (N_11866,N_11757,N_11625);
xor U11867 (N_11867,N_11698,N_11681);
nor U11868 (N_11868,N_11771,N_11721);
nand U11869 (N_11869,N_11773,N_11742);
nor U11870 (N_11870,N_11783,N_11626);
or U11871 (N_11871,N_11604,N_11713);
xor U11872 (N_11872,N_11775,N_11793);
or U11873 (N_11873,N_11761,N_11606);
nor U11874 (N_11874,N_11608,N_11769);
xor U11875 (N_11875,N_11765,N_11799);
and U11876 (N_11876,N_11728,N_11648);
nor U11877 (N_11877,N_11703,N_11615);
nand U11878 (N_11878,N_11790,N_11617);
or U11879 (N_11879,N_11733,N_11693);
or U11880 (N_11880,N_11719,N_11791);
xor U11881 (N_11881,N_11710,N_11688);
or U11882 (N_11882,N_11683,N_11752);
and U11883 (N_11883,N_11777,N_11694);
nor U11884 (N_11884,N_11675,N_11755);
nand U11885 (N_11885,N_11677,N_11632);
nand U11886 (N_11886,N_11674,N_11724);
nor U11887 (N_11887,N_11738,N_11796);
nor U11888 (N_11888,N_11679,N_11709);
nand U11889 (N_11889,N_11794,N_11730);
nand U11890 (N_11890,N_11704,N_11712);
and U11891 (N_11891,N_11691,N_11780);
xor U11892 (N_11892,N_11668,N_11629);
xor U11893 (N_11893,N_11702,N_11737);
nand U11894 (N_11894,N_11631,N_11749);
or U11895 (N_11895,N_11751,N_11646);
nor U11896 (N_11896,N_11722,N_11747);
xnor U11897 (N_11897,N_11650,N_11707);
xnor U11898 (N_11898,N_11635,N_11663);
nor U11899 (N_11899,N_11735,N_11754);
nor U11900 (N_11900,N_11719,N_11735);
or U11901 (N_11901,N_11794,N_11665);
nor U11902 (N_11902,N_11680,N_11622);
or U11903 (N_11903,N_11688,N_11766);
xnor U11904 (N_11904,N_11666,N_11792);
nor U11905 (N_11905,N_11697,N_11692);
or U11906 (N_11906,N_11631,N_11645);
and U11907 (N_11907,N_11646,N_11788);
nor U11908 (N_11908,N_11787,N_11768);
or U11909 (N_11909,N_11768,N_11704);
or U11910 (N_11910,N_11792,N_11679);
nand U11911 (N_11911,N_11677,N_11790);
nor U11912 (N_11912,N_11754,N_11739);
nor U11913 (N_11913,N_11622,N_11743);
or U11914 (N_11914,N_11764,N_11769);
xor U11915 (N_11915,N_11785,N_11704);
nor U11916 (N_11916,N_11718,N_11686);
or U11917 (N_11917,N_11736,N_11622);
xnor U11918 (N_11918,N_11733,N_11785);
and U11919 (N_11919,N_11627,N_11640);
or U11920 (N_11920,N_11679,N_11684);
or U11921 (N_11921,N_11790,N_11668);
xnor U11922 (N_11922,N_11715,N_11733);
nand U11923 (N_11923,N_11702,N_11606);
nand U11924 (N_11924,N_11700,N_11791);
and U11925 (N_11925,N_11799,N_11676);
and U11926 (N_11926,N_11607,N_11693);
and U11927 (N_11927,N_11622,N_11645);
nor U11928 (N_11928,N_11648,N_11609);
nor U11929 (N_11929,N_11735,N_11790);
nor U11930 (N_11930,N_11649,N_11702);
xor U11931 (N_11931,N_11770,N_11600);
nor U11932 (N_11932,N_11725,N_11735);
xor U11933 (N_11933,N_11623,N_11793);
nand U11934 (N_11934,N_11762,N_11681);
nand U11935 (N_11935,N_11730,N_11742);
or U11936 (N_11936,N_11727,N_11732);
nor U11937 (N_11937,N_11648,N_11606);
xnor U11938 (N_11938,N_11762,N_11791);
nor U11939 (N_11939,N_11709,N_11742);
xnor U11940 (N_11940,N_11694,N_11611);
nor U11941 (N_11941,N_11604,N_11629);
xnor U11942 (N_11942,N_11728,N_11770);
xor U11943 (N_11943,N_11683,N_11661);
xnor U11944 (N_11944,N_11749,N_11600);
and U11945 (N_11945,N_11730,N_11668);
nor U11946 (N_11946,N_11620,N_11796);
nor U11947 (N_11947,N_11729,N_11781);
xnor U11948 (N_11948,N_11622,N_11642);
nand U11949 (N_11949,N_11715,N_11685);
and U11950 (N_11950,N_11729,N_11660);
nor U11951 (N_11951,N_11720,N_11684);
nor U11952 (N_11952,N_11741,N_11711);
and U11953 (N_11953,N_11740,N_11643);
nor U11954 (N_11954,N_11758,N_11703);
nand U11955 (N_11955,N_11636,N_11687);
nand U11956 (N_11956,N_11735,N_11684);
and U11957 (N_11957,N_11750,N_11738);
xor U11958 (N_11958,N_11677,N_11665);
nor U11959 (N_11959,N_11699,N_11669);
nand U11960 (N_11960,N_11726,N_11774);
nor U11961 (N_11961,N_11742,N_11725);
nand U11962 (N_11962,N_11728,N_11647);
and U11963 (N_11963,N_11670,N_11628);
nand U11964 (N_11964,N_11770,N_11664);
nand U11965 (N_11965,N_11728,N_11687);
nand U11966 (N_11966,N_11626,N_11650);
and U11967 (N_11967,N_11603,N_11712);
and U11968 (N_11968,N_11729,N_11618);
nor U11969 (N_11969,N_11765,N_11621);
or U11970 (N_11970,N_11687,N_11600);
xnor U11971 (N_11971,N_11778,N_11671);
and U11972 (N_11972,N_11748,N_11699);
xnor U11973 (N_11973,N_11623,N_11732);
or U11974 (N_11974,N_11622,N_11655);
nand U11975 (N_11975,N_11760,N_11625);
nor U11976 (N_11976,N_11727,N_11790);
or U11977 (N_11977,N_11622,N_11757);
and U11978 (N_11978,N_11621,N_11638);
and U11979 (N_11979,N_11672,N_11675);
or U11980 (N_11980,N_11780,N_11676);
xnor U11981 (N_11981,N_11673,N_11700);
nor U11982 (N_11982,N_11647,N_11763);
nor U11983 (N_11983,N_11613,N_11641);
nor U11984 (N_11984,N_11735,N_11779);
or U11985 (N_11985,N_11671,N_11713);
and U11986 (N_11986,N_11642,N_11648);
nor U11987 (N_11987,N_11752,N_11756);
nand U11988 (N_11988,N_11636,N_11603);
xnor U11989 (N_11989,N_11713,N_11721);
and U11990 (N_11990,N_11763,N_11604);
nor U11991 (N_11991,N_11764,N_11713);
nand U11992 (N_11992,N_11729,N_11703);
nor U11993 (N_11993,N_11731,N_11794);
nand U11994 (N_11994,N_11739,N_11658);
xor U11995 (N_11995,N_11645,N_11705);
nand U11996 (N_11996,N_11729,N_11670);
nor U11997 (N_11997,N_11624,N_11616);
or U11998 (N_11998,N_11707,N_11662);
nand U11999 (N_11999,N_11736,N_11709);
and U12000 (N_12000,N_11932,N_11831);
or U12001 (N_12001,N_11843,N_11865);
xnor U12002 (N_12002,N_11827,N_11954);
nand U12003 (N_12003,N_11918,N_11888);
and U12004 (N_12004,N_11876,N_11858);
nor U12005 (N_12005,N_11812,N_11874);
nor U12006 (N_12006,N_11961,N_11962);
nor U12007 (N_12007,N_11811,N_11863);
nor U12008 (N_12008,N_11956,N_11845);
or U12009 (N_12009,N_11909,N_11927);
or U12010 (N_12010,N_11853,N_11809);
nor U12011 (N_12011,N_11913,N_11866);
nor U12012 (N_12012,N_11902,N_11930);
nor U12013 (N_12013,N_11835,N_11971);
nand U12014 (N_12014,N_11905,N_11878);
and U12015 (N_12015,N_11993,N_11982);
or U12016 (N_12016,N_11979,N_11875);
and U12017 (N_12017,N_11841,N_11818);
xnor U12018 (N_12018,N_11872,N_11969);
or U12019 (N_12019,N_11936,N_11973);
nor U12020 (N_12020,N_11937,N_11912);
nand U12021 (N_12021,N_11908,N_11907);
or U12022 (N_12022,N_11972,N_11931);
nand U12023 (N_12023,N_11800,N_11990);
nand U12024 (N_12024,N_11964,N_11922);
or U12025 (N_12025,N_11824,N_11934);
xnor U12026 (N_12026,N_11994,N_11946);
or U12027 (N_12027,N_11816,N_11830);
or U12028 (N_12028,N_11923,N_11940);
and U12029 (N_12029,N_11917,N_11986);
xor U12030 (N_12030,N_11895,N_11883);
or U12031 (N_12031,N_11920,N_11857);
nor U12032 (N_12032,N_11911,N_11861);
and U12033 (N_12033,N_11980,N_11896);
nand U12034 (N_12034,N_11886,N_11882);
xnor U12035 (N_12035,N_11869,N_11846);
or U12036 (N_12036,N_11868,N_11996);
nor U12037 (N_12037,N_11915,N_11806);
nand U12038 (N_12038,N_11885,N_11814);
or U12039 (N_12039,N_11807,N_11856);
nor U12040 (N_12040,N_11832,N_11897);
nand U12041 (N_12041,N_11975,N_11823);
xor U12042 (N_12042,N_11847,N_11995);
and U12043 (N_12043,N_11985,N_11963);
nand U12044 (N_12044,N_11839,N_11810);
nand U12045 (N_12045,N_11953,N_11851);
or U12046 (N_12046,N_11850,N_11826);
nor U12047 (N_12047,N_11881,N_11855);
nor U12048 (N_12048,N_11877,N_11989);
xnor U12049 (N_12049,N_11849,N_11828);
xnor U12050 (N_12050,N_11898,N_11991);
nor U12051 (N_12051,N_11801,N_11862);
xor U12052 (N_12052,N_11992,N_11948);
or U12053 (N_12053,N_11904,N_11943);
nor U12054 (N_12054,N_11804,N_11891);
xnor U12055 (N_12055,N_11852,N_11935);
xnor U12056 (N_12056,N_11997,N_11802);
and U12057 (N_12057,N_11929,N_11871);
and U12058 (N_12058,N_11941,N_11813);
and U12059 (N_12059,N_11938,N_11834);
or U12060 (N_12060,N_11844,N_11970);
xor U12061 (N_12061,N_11854,N_11819);
or U12062 (N_12062,N_11822,N_11833);
xor U12063 (N_12063,N_11999,N_11951);
or U12064 (N_12064,N_11981,N_11817);
nand U12065 (N_12065,N_11884,N_11949);
xor U12066 (N_12066,N_11960,N_11958);
nand U12067 (N_12067,N_11890,N_11837);
and U12068 (N_12068,N_11906,N_11836);
nand U12069 (N_12069,N_11910,N_11880);
and U12070 (N_12070,N_11914,N_11959);
and U12071 (N_12071,N_11947,N_11860);
nand U12072 (N_12072,N_11892,N_11899);
xor U12073 (N_12073,N_11848,N_11903);
nand U12074 (N_12074,N_11829,N_11955);
and U12075 (N_12075,N_11950,N_11939);
nor U12076 (N_12076,N_11803,N_11901);
xor U12077 (N_12077,N_11998,N_11820);
and U12078 (N_12078,N_11842,N_11919);
xor U12079 (N_12079,N_11983,N_11952);
nand U12080 (N_12080,N_11967,N_11870);
nor U12081 (N_12081,N_11900,N_11887);
nor U12082 (N_12082,N_11942,N_11879);
xor U12083 (N_12083,N_11925,N_11815);
xor U12084 (N_12084,N_11987,N_11957);
nand U12085 (N_12085,N_11838,N_11924);
and U12086 (N_12086,N_11821,N_11988);
xnor U12087 (N_12087,N_11825,N_11928);
nor U12088 (N_12088,N_11808,N_11864);
and U12089 (N_12089,N_11968,N_11926);
or U12090 (N_12090,N_11984,N_11944);
xnor U12091 (N_12091,N_11894,N_11966);
xnor U12092 (N_12092,N_11893,N_11916);
or U12093 (N_12093,N_11974,N_11976);
nor U12094 (N_12094,N_11867,N_11965);
xnor U12095 (N_12095,N_11921,N_11977);
and U12096 (N_12096,N_11840,N_11933);
xor U12097 (N_12097,N_11859,N_11805);
and U12098 (N_12098,N_11945,N_11873);
xnor U12099 (N_12099,N_11978,N_11889);
xor U12100 (N_12100,N_11937,N_11862);
or U12101 (N_12101,N_11921,N_11934);
xor U12102 (N_12102,N_11851,N_11905);
xnor U12103 (N_12103,N_11939,N_11907);
xnor U12104 (N_12104,N_11906,N_11803);
or U12105 (N_12105,N_11959,N_11859);
xnor U12106 (N_12106,N_11943,N_11907);
nand U12107 (N_12107,N_11835,N_11983);
nand U12108 (N_12108,N_11891,N_11937);
nor U12109 (N_12109,N_11871,N_11879);
or U12110 (N_12110,N_11897,N_11997);
and U12111 (N_12111,N_11927,N_11918);
or U12112 (N_12112,N_11932,N_11893);
xor U12113 (N_12113,N_11956,N_11801);
nor U12114 (N_12114,N_11875,N_11984);
and U12115 (N_12115,N_11980,N_11919);
xor U12116 (N_12116,N_11878,N_11812);
or U12117 (N_12117,N_11946,N_11821);
nand U12118 (N_12118,N_11927,N_11924);
xor U12119 (N_12119,N_11871,N_11829);
nor U12120 (N_12120,N_11900,N_11960);
nand U12121 (N_12121,N_11867,N_11910);
or U12122 (N_12122,N_11979,N_11921);
nand U12123 (N_12123,N_11869,N_11856);
nor U12124 (N_12124,N_11964,N_11832);
or U12125 (N_12125,N_11923,N_11885);
or U12126 (N_12126,N_11850,N_11925);
xor U12127 (N_12127,N_11800,N_11898);
nor U12128 (N_12128,N_11974,N_11966);
xor U12129 (N_12129,N_11863,N_11959);
xnor U12130 (N_12130,N_11978,N_11971);
nor U12131 (N_12131,N_11920,N_11954);
and U12132 (N_12132,N_11841,N_11933);
nor U12133 (N_12133,N_11911,N_11824);
xnor U12134 (N_12134,N_11850,N_11836);
or U12135 (N_12135,N_11972,N_11881);
nand U12136 (N_12136,N_11930,N_11969);
nor U12137 (N_12137,N_11841,N_11836);
nand U12138 (N_12138,N_11983,N_11842);
and U12139 (N_12139,N_11955,N_11920);
xor U12140 (N_12140,N_11966,N_11865);
nor U12141 (N_12141,N_11882,N_11939);
and U12142 (N_12142,N_11989,N_11980);
nor U12143 (N_12143,N_11829,N_11864);
and U12144 (N_12144,N_11836,N_11802);
and U12145 (N_12145,N_11939,N_11975);
xnor U12146 (N_12146,N_11807,N_11953);
or U12147 (N_12147,N_11943,N_11911);
xnor U12148 (N_12148,N_11860,N_11935);
or U12149 (N_12149,N_11959,N_11899);
and U12150 (N_12150,N_11951,N_11854);
and U12151 (N_12151,N_11975,N_11859);
or U12152 (N_12152,N_11916,N_11988);
or U12153 (N_12153,N_11952,N_11803);
xnor U12154 (N_12154,N_11843,N_11827);
xor U12155 (N_12155,N_11912,N_11903);
nand U12156 (N_12156,N_11832,N_11872);
nand U12157 (N_12157,N_11843,N_11940);
and U12158 (N_12158,N_11990,N_11994);
nor U12159 (N_12159,N_11978,N_11963);
xnor U12160 (N_12160,N_11891,N_11918);
or U12161 (N_12161,N_11827,N_11900);
xnor U12162 (N_12162,N_11838,N_11894);
nand U12163 (N_12163,N_11857,N_11845);
and U12164 (N_12164,N_11845,N_11930);
nand U12165 (N_12165,N_11883,N_11816);
nor U12166 (N_12166,N_11852,N_11861);
or U12167 (N_12167,N_11968,N_11893);
and U12168 (N_12168,N_11845,N_11863);
nor U12169 (N_12169,N_11834,N_11922);
or U12170 (N_12170,N_11834,N_11965);
nand U12171 (N_12171,N_11967,N_11969);
or U12172 (N_12172,N_11924,N_11891);
nor U12173 (N_12173,N_11896,N_11901);
and U12174 (N_12174,N_11972,N_11983);
and U12175 (N_12175,N_11813,N_11995);
nor U12176 (N_12176,N_11955,N_11877);
and U12177 (N_12177,N_11995,N_11940);
nand U12178 (N_12178,N_11878,N_11907);
nor U12179 (N_12179,N_11945,N_11809);
or U12180 (N_12180,N_11955,N_11891);
and U12181 (N_12181,N_11823,N_11888);
and U12182 (N_12182,N_11910,N_11881);
xnor U12183 (N_12183,N_11866,N_11920);
and U12184 (N_12184,N_11833,N_11930);
nor U12185 (N_12185,N_11857,N_11918);
xor U12186 (N_12186,N_11971,N_11915);
nor U12187 (N_12187,N_11879,N_11976);
or U12188 (N_12188,N_11820,N_11928);
or U12189 (N_12189,N_11860,N_11834);
or U12190 (N_12190,N_11876,N_11934);
nand U12191 (N_12191,N_11842,N_11877);
nand U12192 (N_12192,N_11882,N_11918);
nor U12193 (N_12193,N_11889,N_11944);
xor U12194 (N_12194,N_11928,N_11837);
nand U12195 (N_12195,N_11905,N_11861);
xnor U12196 (N_12196,N_11938,N_11921);
or U12197 (N_12197,N_11994,N_11982);
and U12198 (N_12198,N_11904,N_11802);
or U12199 (N_12199,N_11908,N_11966);
nand U12200 (N_12200,N_12026,N_12028);
and U12201 (N_12201,N_12017,N_12152);
or U12202 (N_12202,N_12104,N_12058);
nand U12203 (N_12203,N_12176,N_12053);
xnor U12204 (N_12204,N_12154,N_12137);
nor U12205 (N_12205,N_12052,N_12096);
or U12206 (N_12206,N_12078,N_12118);
nor U12207 (N_12207,N_12165,N_12110);
nand U12208 (N_12208,N_12044,N_12039);
nor U12209 (N_12209,N_12196,N_12088);
and U12210 (N_12210,N_12198,N_12151);
nor U12211 (N_12211,N_12109,N_12159);
or U12212 (N_12212,N_12068,N_12032);
nand U12213 (N_12213,N_12021,N_12150);
xor U12214 (N_12214,N_12130,N_12171);
or U12215 (N_12215,N_12116,N_12157);
xor U12216 (N_12216,N_12036,N_12147);
nand U12217 (N_12217,N_12010,N_12190);
nand U12218 (N_12218,N_12120,N_12013);
xnor U12219 (N_12219,N_12061,N_12112);
or U12220 (N_12220,N_12169,N_12046);
nand U12221 (N_12221,N_12059,N_12091);
xor U12222 (N_12222,N_12014,N_12107);
nor U12223 (N_12223,N_12106,N_12144);
nand U12224 (N_12224,N_12136,N_12166);
and U12225 (N_12225,N_12023,N_12015);
nand U12226 (N_12226,N_12134,N_12108);
and U12227 (N_12227,N_12094,N_12125);
xor U12228 (N_12228,N_12089,N_12082);
nor U12229 (N_12229,N_12191,N_12161);
and U12230 (N_12230,N_12189,N_12079);
nor U12231 (N_12231,N_12073,N_12183);
or U12232 (N_12232,N_12076,N_12135);
nor U12233 (N_12233,N_12143,N_12133);
nor U12234 (N_12234,N_12123,N_12177);
nor U12235 (N_12235,N_12004,N_12060);
and U12236 (N_12236,N_12156,N_12007);
or U12237 (N_12237,N_12139,N_12128);
xnor U12238 (N_12238,N_12074,N_12000);
or U12239 (N_12239,N_12031,N_12069);
and U12240 (N_12240,N_12077,N_12100);
or U12241 (N_12241,N_12054,N_12083);
xor U12242 (N_12242,N_12018,N_12034);
xnor U12243 (N_12243,N_12081,N_12194);
and U12244 (N_12244,N_12111,N_12199);
nor U12245 (N_12245,N_12178,N_12142);
or U12246 (N_12246,N_12181,N_12168);
xor U12247 (N_12247,N_12114,N_12001);
or U12248 (N_12248,N_12048,N_12187);
xnor U12249 (N_12249,N_12050,N_12188);
nor U12250 (N_12250,N_12124,N_12092);
nor U12251 (N_12251,N_12121,N_12006);
and U12252 (N_12252,N_12155,N_12072);
nor U12253 (N_12253,N_12167,N_12038);
xnor U12254 (N_12254,N_12027,N_12024);
nor U12255 (N_12255,N_12115,N_12041);
nand U12256 (N_12256,N_12186,N_12005);
or U12257 (N_12257,N_12160,N_12097);
xor U12258 (N_12258,N_12179,N_12148);
xor U12259 (N_12259,N_12063,N_12117);
xnor U12260 (N_12260,N_12016,N_12003);
nor U12261 (N_12261,N_12062,N_12030);
xnor U12262 (N_12262,N_12129,N_12174);
nand U12263 (N_12263,N_12011,N_12085);
nor U12264 (N_12264,N_12101,N_12009);
xnor U12265 (N_12265,N_12035,N_12019);
xnor U12266 (N_12266,N_12057,N_12126);
and U12267 (N_12267,N_12029,N_12040);
nor U12268 (N_12268,N_12158,N_12193);
or U12269 (N_12269,N_12051,N_12055);
nand U12270 (N_12270,N_12087,N_12025);
or U12271 (N_12271,N_12163,N_12037);
and U12272 (N_12272,N_12197,N_12105);
xnor U12273 (N_12273,N_12182,N_12008);
nor U12274 (N_12274,N_12012,N_12095);
nand U12275 (N_12275,N_12127,N_12084);
nor U12276 (N_12276,N_12002,N_12043);
xnor U12277 (N_12277,N_12149,N_12192);
and U12278 (N_12278,N_12138,N_12047);
nand U12279 (N_12279,N_12103,N_12071);
xor U12280 (N_12280,N_12064,N_12070);
nand U12281 (N_12281,N_12122,N_12145);
xor U12282 (N_12282,N_12173,N_12146);
or U12283 (N_12283,N_12172,N_12153);
and U12284 (N_12284,N_12098,N_12184);
xnor U12285 (N_12285,N_12056,N_12132);
nand U12286 (N_12286,N_12119,N_12141);
and U12287 (N_12287,N_12065,N_12042);
xnor U12288 (N_12288,N_12075,N_12045);
nand U12289 (N_12289,N_12099,N_12102);
and U12290 (N_12290,N_12020,N_12067);
nand U12291 (N_12291,N_12090,N_12113);
xor U12292 (N_12292,N_12170,N_12022);
or U12293 (N_12293,N_12140,N_12162);
or U12294 (N_12294,N_12195,N_12185);
and U12295 (N_12295,N_12180,N_12086);
nand U12296 (N_12296,N_12066,N_12131);
and U12297 (N_12297,N_12164,N_12049);
nor U12298 (N_12298,N_12175,N_12093);
nand U12299 (N_12299,N_12080,N_12033);
nor U12300 (N_12300,N_12117,N_12126);
xnor U12301 (N_12301,N_12034,N_12164);
xor U12302 (N_12302,N_12179,N_12185);
xor U12303 (N_12303,N_12067,N_12072);
or U12304 (N_12304,N_12092,N_12110);
nor U12305 (N_12305,N_12013,N_12156);
and U12306 (N_12306,N_12042,N_12134);
nor U12307 (N_12307,N_12196,N_12016);
nand U12308 (N_12308,N_12096,N_12069);
nand U12309 (N_12309,N_12076,N_12159);
xor U12310 (N_12310,N_12158,N_12175);
or U12311 (N_12311,N_12141,N_12035);
and U12312 (N_12312,N_12176,N_12128);
nor U12313 (N_12313,N_12151,N_12107);
nor U12314 (N_12314,N_12085,N_12070);
and U12315 (N_12315,N_12113,N_12167);
nor U12316 (N_12316,N_12133,N_12081);
or U12317 (N_12317,N_12146,N_12186);
or U12318 (N_12318,N_12022,N_12193);
and U12319 (N_12319,N_12195,N_12058);
and U12320 (N_12320,N_12144,N_12157);
xnor U12321 (N_12321,N_12112,N_12153);
and U12322 (N_12322,N_12096,N_12152);
nor U12323 (N_12323,N_12042,N_12082);
nand U12324 (N_12324,N_12007,N_12122);
xnor U12325 (N_12325,N_12049,N_12017);
and U12326 (N_12326,N_12004,N_12175);
and U12327 (N_12327,N_12121,N_12031);
nand U12328 (N_12328,N_12185,N_12000);
nor U12329 (N_12329,N_12039,N_12046);
and U12330 (N_12330,N_12157,N_12044);
and U12331 (N_12331,N_12099,N_12189);
or U12332 (N_12332,N_12128,N_12022);
nand U12333 (N_12333,N_12145,N_12112);
nor U12334 (N_12334,N_12032,N_12034);
nor U12335 (N_12335,N_12019,N_12096);
or U12336 (N_12336,N_12046,N_12195);
and U12337 (N_12337,N_12019,N_12031);
nand U12338 (N_12338,N_12197,N_12171);
nor U12339 (N_12339,N_12048,N_12106);
nor U12340 (N_12340,N_12011,N_12098);
xnor U12341 (N_12341,N_12166,N_12010);
nor U12342 (N_12342,N_12134,N_12084);
nand U12343 (N_12343,N_12008,N_12140);
nor U12344 (N_12344,N_12059,N_12177);
nor U12345 (N_12345,N_12031,N_12101);
nor U12346 (N_12346,N_12119,N_12143);
nor U12347 (N_12347,N_12136,N_12172);
xnor U12348 (N_12348,N_12072,N_12008);
nand U12349 (N_12349,N_12106,N_12011);
nand U12350 (N_12350,N_12129,N_12068);
or U12351 (N_12351,N_12043,N_12126);
nand U12352 (N_12352,N_12114,N_12044);
or U12353 (N_12353,N_12062,N_12072);
nand U12354 (N_12354,N_12046,N_12098);
or U12355 (N_12355,N_12029,N_12000);
and U12356 (N_12356,N_12156,N_12050);
or U12357 (N_12357,N_12032,N_12013);
nand U12358 (N_12358,N_12160,N_12108);
nor U12359 (N_12359,N_12115,N_12051);
xor U12360 (N_12360,N_12087,N_12102);
xnor U12361 (N_12361,N_12195,N_12140);
nor U12362 (N_12362,N_12121,N_12107);
nand U12363 (N_12363,N_12025,N_12183);
nand U12364 (N_12364,N_12020,N_12089);
xnor U12365 (N_12365,N_12144,N_12059);
and U12366 (N_12366,N_12038,N_12002);
nand U12367 (N_12367,N_12159,N_12148);
or U12368 (N_12368,N_12196,N_12046);
or U12369 (N_12369,N_12005,N_12001);
nand U12370 (N_12370,N_12028,N_12110);
or U12371 (N_12371,N_12101,N_12124);
or U12372 (N_12372,N_12144,N_12167);
nor U12373 (N_12373,N_12003,N_12020);
xor U12374 (N_12374,N_12015,N_12039);
xnor U12375 (N_12375,N_12009,N_12161);
nor U12376 (N_12376,N_12012,N_12122);
or U12377 (N_12377,N_12109,N_12117);
nand U12378 (N_12378,N_12195,N_12149);
and U12379 (N_12379,N_12008,N_12077);
and U12380 (N_12380,N_12025,N_12122);
nand U12381 (N_12381,N_12166,N_12043);
nor U12382 (N_12382,N_12107,N_12087);
and U12383 (N_12383,N_12180,N_12062);
and U12384 (N_12384,N_12064,N_12099);
and U12385 (N_12385,N_12035,N_12140);
nor U12386 (N_12386,N_12146,N_12094);
xor U12387 (N_12387,N_12079,N_12148);
xor U12388 (N_12388,N_12087,N_12010);
nor U12389 (N_12389,N_12023,N_12075);
and U12390 (N_12390,N_12048,N_12121);
or U12391 (N_12391,N_12193,N_12181);
nand U12392 (N_12392,N_12166,N_12062);
nor U12393 (N_12393,N_12021,N_12195);
or U12394 (N_12394,N_12111,N_12109);
and U12395 (N_12395,N_12079,N_12186);
nor U12396 (N_12396,N_12097,N_12132);
and U12397 (N_12397,N_12123,N_12074);
nor U12398 (N_12398,N_12132,N_12021);
xor U12399 (N_12399,N_12177,N_12009);
and U12400 (N_12400,N_12239,N_12309);
nor U12401 (N_12401,N_12210,N_12338);
nor U12402 (N_12402,N_12231,N_12328);
and U12403 (N_12403,N_12234,N_12261);
nand U12404 (N_12404,N_12284,N_12362);
nand U12405 (N_12405,N_12256,N_12283);
nand U12406 (N_12406,N_12297,N_12312);
or U12407 (N_12407,N_12357,N_12258);
and U12408 (N_12408,N_12219,N_12390);
and U12409 (N_12409,N_12385,N_12295);
nor U12410 (N_12410,N_12388,N_12293);
nand U12411 (N_12411,N_12236,N_12369);
or U12412 (N_12412,N_12350,N_12339);
nand U12413 (N_12413,N_12399,N_12370);
nor U12414 (N_12414,N_12241,N_12202);
nand U12415 (N_12415,N_12319,N_12215);
xnor U12416 (N_12416,N_12200,N_12213);
and U12417 (N_12417,N_12227,N_12310);
or U12418 (N_12418,N_12279,N_12228);
or U12419 (N_12419,N_12320,N_12230);
or U12420 (N_12420,N_12377,N_12305);
and U12421 (N_12421,N_12367,N_12285);
or U12422 (N_12422,N_12307,N_12243);
nand U12423 (N_12423,N_12220,N_12380);
nand U12424 (N_12424,N_12308,N_12291);
xor U12425 (N_12425,N_12366,N_12379);
nor U12426 (N_12426,N_12334,N_12251);
nand U12427 (N_12427,N_12317,N_12269);
or U12428 (N_12428,N_12206,N_12209);
nand U12429 (N_12429,N_12267,N_12292);
nor U12430 (N_12430,N_12356,N_12257);
and U12431 (N_12431,N_12363,N_12347);
and U12432 (N_12432,N_12337,N_12351);
or U12433 (N_12433,N_12325,N_12371);
or U12434 (N_12434,N_12264,N_12315);
nand U12435 (N_12435,N_12259,N_12298);
xnor U12436 (N_12436,N_12262,N_12216);
or U12437 (N_12437,N_12286,N_12232);
xnor U12438 (N_12438,N_12300,N_12349);
xor U12439 (N_12439,N_12278,N_12266);
and U12440 (N_12440,N_12276,N_12393);
nor U12441 (N_12441,N_12205,N_12341);
or U12442 (N_12442,N_12247,N_12391);
nand U12443 (N_12443,N_12288,N_12384);
nor U12444 (N_12444,N_12280,N_12224);
nor U12445 (N_12445,N_12395,N_12277);
and U12446 (N_12446,N_12218,N_12360);
and U12447 (N_12447,N_12252,N_12263);
nand U12448 (N_12448,N_12354,N_12306);
nor U12449 (N_12449,N_12389,N_12212);
and U12450 (N_12450,N_12394,N_12348);
xor U12451 (N_12451,N_12359,N_12346);
xor U12452 (N_12452,N_12233,N_12235);
nor U12453 (N_12453,N_12222,N_12274);
or U12454 (N_12454,N_12343,N_12345);
and U12455 (N_12455,N_12270,N_12253);
and U12456 (N_12456,N_12381,N_12301);
nor U12457 (N_12457,N_12245,N_12373);
xnor U12458 (N_12458,N_12323,N_12226);
nand U12459 (N_12459,N_12392,N_12335);
or U12460 (N_12460,N_12217,N_12229);
or U12461 (N_12461,N_12322,N_12327);
or U12462 (N_12462,N_12299,N_12340);
xnor U12463 (N_12463,N_12324,N_12376);
and U12464 (N_12464,N_12225,N_12248);
nor U12465 (N_12465,N_12275,N_12353);
xor U12466 (N_12466,N_12282,N_12303);
nor U12467 (N_12467,N_12221,N_12290);
nor U12468 (N_12468,N_12204,N_12246);
xor U12469 (N_12469,N_12260,N_12387);
nand U12470 (N_12470,N_12240,N_12208);
xnor U12471 (N_12471,N_12313,N_12254);
xor U12472 (N_12472,N_12333,N_12365);
nand U12473 (N_12473,N_12326,N_12368);
nand U12474 (N_12474,N_12355,N_12203);
and U12475 (N_12475,N_12302,N_12265);
nand U12476 (N_12476,N_12398,N_12294);
xnor U12477 (N_12477,N_12255,N_12383);
and U12478 (N_12478,N_12314,N_12242);
nor U12479 (N_12479,N_12268,N_12375);
nand U12480 (N_12480,N_12364,N_12304);
and U12481 (N_12481,N_12223,N_12372);
nand U12482 (N_12482,N_12331,N_12238);
nand U12483 (N_12483,N_12358,N_12397);
nor U12484 (N_12484,N_12361,N_12396);
nor U12485 (N_12485,N_12329,N_12296);
nand U12486 (N_12486,N_12336,N_12271);
and U12487 (N_12487,N_12237,N_12386);
and U12488 (N_12488,N_12316,N_12211);
xor U12489 (N_12489,N_12272,N_12374);
nor U12490 (N_12490,N_12378,N_12249);
or U12491 (N_12491,N_12287,N_12214);
nor U12492 (N_12492,N_12273,N_12244);
and U12493 (N_12493,N_12318,N_12332);
nor U12494 (N_12494,N_12281,N_12382);
or U12495 (N_12495,N_12344,N_12207);
xnor U12496 (N_12496,N_12342,N_12352);
and U12497 (N_12497,N_12250,N_12311);
nand U12498 (N_12498,N_12330,N_12201);
and U12499 (N_12499,N_12289,N_12321);
and U12500 (N_12500,N_12348,N_12318);
xor U12501 (N_12501,N_12363,N_12374);
or U12502 (N_12502,N_12310,N_12355);
and U12503 (N_12503,N_12373,N_12233);
nor U12504 (N_12504,N_12332,N_12319);
xor U12505 (N_12505,N_12244,N_12304);
nand U12506 (N_12506,N_12363,N_12371);
and U12507 (N_12507,N_12330,N_12349);
nand U12508 (N_12508,N_12386,N_12304);
or U12509 (N_12509,N_12395,N_12359);
nor U12510 (N_12510,N_12232,N_12281);
nand U12511 (N_12511,N_12374,N_12334);
and U12512 (N_12512,N_12309,N_12221);
or U12513 (N_12513,N_12324,N_12396);
nor U12514 (N_12514,N_12257,N_12351);
nand U12515 (N_12515,N_12364,N_12290);
xor U12516 (N_12516,N_12353,N_12386);
or U12517 (N_12517,N_12252,N_12376);
xnor U12518 (N_12518,N_12215,N_12342);
nand U12519 (N_12519,N_12276,N_12216);
and U12520 (N_12520,N_12243,N_12215);
or U12521 (N_12521,N_12297,N_12210);
nor U12522 (N_12522,N_12361,N_12389);
and U12523 (N_12523,N_12311,N_12252);
and U12524 (N_12524,N_12346,N_12364);
nor U12525 (N_12525,N_12267,N_12306);
and U12526 (N_12526,N_12303,N_12337);
xnor U12527 (N_12527,N_12294,N_12289);
and U12528 (N_12528,N_12262,N_12348);
nor U12529 (N_12529,N_12201,N_12254);
nor U12530 (N_12530,N_12325,N_12343);
nand U12531 (N_12531,N_12229,N_12376);
or U12532 (N_12532,N_12345,N_12229);
and U12533 (N_12533,N_12212,N_12231);
and U12534 (N_12534,N_12266,N_12365);
or U12535 (N_12535,N_12363,N_12266);
xor U12536 (N_12536,N_12289,N_12395);
nand U12537 (N_12537,N_12252,N_12207);
and U12538 (N_12538,N_12346,N_12394);
nand U12539 (N_12539,N_12275,N_12280);
nor U12540 (N_12540,N_12295,N_12246);
nor U12541 (N_12541,N_12205,N_12219);
nor U12542 (N_12542,N_12289,N_12280);
nand U12543 (N_12543,N_12216,N_12271);
nor U12544 (N_12544,N_12373,N_12355);
and U12545 (N_12545,N_12295,N_12315);
or U12546 (N_12546,N_12333,N_12335);
nor U12547 (N_12547,N_12211,N_12342);
xor U12548 (N_12548,N_12263,N_12385);
nand U12549 (N_12549,N_12202,N_12281);
nand U12550 (N_12550,N_12262,N_12270);
or U12551 (N_12551,N_12362,N_12348);
or U12552 (N_12552,N_12209,N_12307);
and U12553 (N_12553,N_12290,N_12391);
and U12554 (N_12554,N_12286,N_12301);
or U12555 (N_12555,N_12227,N_12274);
nor U12556 (N_12556,N_12207,N_12205);
nand U12557 (N_12557,N_12299,N_12257);
or U12558 (N_12558,N_12233,N_12264);
xnor U12559 (N_12559,N_12360,N_12248);
nor U12560 (N_12560,N_12344,N_12366);
and U12561 (N_12561,N_12223,N_12204);
xnor U12562 (N_12562,N_12296,N_12231);
nor U12563 (N_12563,N_12270,N_12365);
xor U12564 (N_12564,N_12377,N_12292);
nor U12565 (N_12565,N_12257,N_12242);
nor U12566 (N_12566,N_12266,N_12248);
and U12567 (N_12567,N_12283,N_12383);
and U12568 (N_12568,N_12277,N_12218);
nor U12569 (N_12569,N_12339,N_12256);
nand U12570 (N_12570,N_12229,N_12228);
nor U12571 (N_12571,N_12346,N_12380);
xnor U12572 (N_12572,N_12278,N_12237);
xnor U12573 (N_12573,N_12344,N_12382);
xor U12574 (N_12574,N_12378,N_12330);
nand U12575 (N_12575,N_12243,N_12288);
nor U12576 (N_12576,N_12282,N_12269);
nor U12577 (N_12577,N_12329,N_12391);
or U12578 (N_12578,N_12248,N_12365);
and U12579 (N_12579,N_12355,N_12225);
or U12580 (N_12580,N_12211,N_12224);
and U12581 (N_12581,N_12213,N_12265);
nand U12582 (N_12582,N_12254,N_12269);
nor U12583 (N_12583,N_12245,N_12209);
xnor U12584 (N_12584,N_12287,N_12235);
and U12585 (N_12585,N_12315,N_12246);
nor U12586 (N_12586,N_12219,N_12334);
nand U12587 (N_12587,N_12260,N_12277);
and U12588 (N_12588,N_12255,N_12251);
or U12589 (N_12589,N_12204,N_12279);
or U12590 (N_12590,N_12279,N_12252);
and U12591 (N_12591,N_12219,N_12283);
xnor U12592 (N_12592,N_12301,N_12314);
or U12593 (N_12593,N_12281,N_12304);
nor U12594 (N_12594,N_12294,N_12389);
or U12595 (N_12595,N_12236,N_12312);
or U12596 (N_12596,N_12317,N_12326);
nand U12597 (N_12597,N_12333,N_12315);
xnor U12598 (N_12598,N_12219,N_12267);
and U12599 (N_12599,N_12289,N_12242);
and U12600 (N_12600,N_12500,N_12506);
and U12601 (N_12601,N_12460,N_12549);
xor U12602 (N_12602,N_12538,N_12548);
nor U12603 (N_12603,N_12450,N_12486);
nor U12604 (N_12604,N_12503,N_12529);
nor U12605 (N_12605,N_12512,N_12598);
or U12606 (N_12606,N_12514,N_12513);
or U12607 (N_12607,N_12413,N_12508);
nand U12608 (N_12608,N_12577,N_12579);
nor U12609 (N_12609,N_12440,N_12449);
xnor U12610 (N_12610,N_12541,N_12414);
nor U12611 (N_12611,N_12583,N_12596);
xor U12612 (N_12612,N_12404,N_12443);
nand U12613 (N_12613,N_12494,N_12571);
and U12614 (N_12614,N_12478,N_12573);
nand U12615 (N_12615,N_12422,N_12570);
xnor U12616 (N_12616,N_12477,N_12578);
nand U12617 (N_12617,N_12431,N_12590);
nor U12618 (N_12618,N_12417,N_12472);
nor U12619 (N_12619,N_12565,N_12507);
and U12620 (N_12620,N_12562,N_12447);
nor U12621 (N_12621,N_12425,N_12516);
and U12622 (N_12622,N_12484,N_12581);
and U12623 (N_12623,N_12521,N_12458);
and U12624 (N_12624,N_12533,N_12580);
xnor U12625 (N_12625,N_12424,N_12461);
and U12626 (N_12626,N_12444,N_12589);
nand U12627 (N_12627,N_12591,N_12531);
xnor U12628 (N_12628,N_12402,N_12466);
xor U12629 (N_12629,N_12409,N_12434);
or U12630 (N_12630,N_12524,N_12481);
xor U12631 (N_12631,N_12445,N_12437);
nor U12632 (N_12632,N_12552,N_12593);
nor U12633 (N_12633,N_12423,N_12496);
nor U12634 (N_12634,N_12530,N_12525);
xor U12635 (N_12635,N_12483,N_12459);
xor U12636 (N_12636,N_12490,N_12534);
or U12637 (N_12637,N_12476,N_12420);
and U12638 (N_12638,N_12535,N_12451);
or U12639 (N_12639,N_12557,N_12493);
and U12640 (N_12640,N_12546,N_12527);
or U12641 (N_12641,N_12412,N_12592);
and U12642 (N_12642,N_12569,N_12563);
nor U12643 (N_12643,N_12501,N_12401);
or U12644 (N_12644,N_12595,N_12482);
and U12645 (N_12645,N_12470,N_12543);
nand U12646 (N_12646,N_12474,N_12553);
or U12647 (N_12647,N_12411,N_12561);
nor U12648 (N_12648,N_12597,N_12436);
nand U12649 (N_12649,N_12406,N_12442);
or U12650 (N_12650,N_12502,N_12454);
or U12651 (N_12651,N_12403,N_12537);
and U12652 (N_12652,N_12519,N_12480);
xor U12653 (N_12653,N_12469,N_12489);
xnor U12654 (N_12654,N_12439,N_12463);
nor U12655 (N_12655,N_12455,N_12560);
xnor U12656 (N_12656,N_12457,N_12576);
nor U12657 (N_12657,N_12433,N_12429);
and U12658 (N_12658,N_12498,N_12567);
or U12659 (N_12659,N_12479,N_12419);
and U12660 (N_12660,N_12599,N_12415);
nand U12661 (N_12661,N_12555,N_12491);
xnor U12662 (N_12662,N_12471,N_12566);
and U12663 (N_12663,N_12568,N_12526);
xnor U12664 (N_12664,N_12550,N_12467);
or U12665 (N_12665,N_12408,N_12544);
nor U12666 (N_12666,N_12556,N_12400);
nor U12667 (N_12667,N_12421,N_12430);
nand U12668 (N_12668,N_12473,N_12574);
nand U12669 (N_12669,N_12585,N_12536);
and U12670 (N_12670,N_12588,N_12492);
and U12671 (N_12671,N_12426,N_12559);
nand U12672 (N_12672,N_12464,N_12594);
nor U12673 (N_12673,N_12584,N_12509);
xor U12674 (N_12674,N_12495,N_12446);
nor U12675 (N_12675,N_12462,N_12582);
and U12676 (N_12676,N_12539,N_12407);
and U12677 (N_12677,N_12518,N_12572);
nor U12678 (N_12678,N_12547,N_12427);
xnor U12679 (N_12679,N_12448,N_12558);
nor U12680 (N_12680,N_12545,N_12586);
nor U12681 (N_12681,N_12453,N_12488);
and U12682 (N_12682,N_12410,N_12428);
xor U12683 (N_12683,N_12418,N_12564);
or U12684 (N_12684,N_12468,N_12499);
nand U12685 (N_12685,N_12432,N_12511);
and U12686 (N_12686,N_12528,N_12485);
nor U12687 (N_12687,N_12515,N_12522);
xnor U12688 (N_12688,N_12435,N_12405);
nor U12689 (N_12689,N_12554,N_12465);
nand U12690 (N_12690,N_12497,N_12540);
or U12691 (N_12691,N_12542,N_12452);
nand U12692 (N_12692,N_12504,N_12520);
or U12693 (N_12693,N_12517,N_12587);
or U12694 (N_12694,N_12438,N_12575);
and U12695 (N_12695,N_12510,N_12456);
nand U12696 (N_12696,N_12416,N_12487);
and U12697 (N_12697,N_12532,N_12441);
nand U12698 (N_12698,N_12475,N_12505);
or U12699 (N_12699,N_12523,N_12551);
xnor U12700 (N_12700,N_12556,N_12423);
xor U12701 (N_12701,N_12585,N_12463);
xnor U12702 (N_12702,N_12459,N_12508);
nand U12703 (N_12703,N_12520,N_12531);
nor U12704 (N_12704,N_12568,N_12480);
and U12705 (N_12705,N_12454,N_12497);
nand U12706 (N_12706,N_12458,N_12546);
nor U12707 (N_12707,N_12533,N_12513);
and U12708 (N_12708,N_12472,N_12545);
nand U12709 (N_12709,N_12492,N_12448);
nor U12710 (N_12710,N_12416,N_12423);
nand U12711 (N_12711,N_12407,N_12552);
or U12712 (N_12712,N_12596,N_12472);
and U12713 (N_12713,N_12523,N_12572);
nand U12714 (N_12714,N_12574,N_12519);
nand U12715 (N_12715,N_12443,N_12464);
nor U12716 (N_12716,N_12474,N_12403);
or U12717 (N_12717,N_12408,N_12502);
or U12718 (N_12718,N_12531,N_12550);
and U12719 (N_12719,N_12595,N_12419);
nor U12720 (N_12720,N_12407,N_12408);
and U12721 (N_12721,N_12446,N_12549);
nor U12722 (N_12722,N_12472,N_12580);
and U12723 (N_12723,N_12567,N_12581);
and U12724 (N_12724,N_12421,N_12534);
nor U12725 (N_12725,N_12495,N_12515);
or U12726 (N_12726,N_12479,N_12439);
and U12727 (N_12727,N_12564,N_12509);
or U12728 (N_12728,N_12565,N_12480);
and U12729 (N_12729,N_12540,N_12492);
and U12730 (N_12730,N_12556,N_12590);
or U12731 (N_12731,N_12403,N_12542);
or U12732 (N_12732,N_12535,N_12412);
nor U12733 (N_12733,N_12523,N_12564);
nor U12734 (N_12734,N_12506,N_12540);
nand U12735 (N_12735,N_12417,N_12491);
or U12736 (N_12736,N_12538,N_12495);
or U12737 (N_12737,N_12444,N_12569);
and U12738 (N_12738,N_12522,N_12548);
nand U12739 (N_12739,N_12542,N_12417);
nand U12740 (N_12740,N_12429,N_12591);
or U12741 (N_12741,N_12586,N_12400);
nand U12742 (N_12742,N_12417,N_12524);
xor U12743 (N_12743,N_12591,N_12419);
nand U12744 (N_12744,N_12515,N_12470);
or U12745 (N_12745,N_12483,N_12598);
or U12746 (N_12746,N_12511,N_12545);
nand U12747 (N_12747,N_12542,N_12582);
and U12748 (N_12748,N_12504,N_12416);
and U12749 (N_12749,N_12543,N_12408);
nor U12750 (N_12750,N_12466,N_12492);
nand U12751 (N_12751,N_12521,N_12497);
or U12752 (N_12752,N_12523,N_12558);
or U12753 (N_12753,N_12409,N_12478);
or U12754 (N_12754,N_12457,N_12531);
and U12755 (N_12755,N_12424,N_12433);
or U12756 (N_12756,N_12531,N_12484);
nor U12757 (N_12757,N_12461,N_12430);
nor U12758 (N_12758,N_12543,N_12573);
and U12759 (N_12759,N_12437,N_12508);
and U12760 (N_12760,N_12408,N_12415);
or U12761 (N_12761,N_12548,N_12553);
xnor U12762 (N_12762,N_12538,N_12421);
xnor U12763 (N_12763,N_12451,N_12590);
and U12764 (N_12764,N_12532,N_12597);
nor U12765 (N_12765,N_12483,N_12495);
nand U12766 (N_12766,N_12402,N_12534);
nand U12767 (N_12767,N_12518,N_12441);
and U12768 (N_12768,N_12462,N_12471);
nor U12769 (N_12769,N_12454,N_12588);
or U12770 (N_12770,N_12496,N_12448);
and U12771 (N_12771,N_12400,N_12537);
nand U12772 (N_12772,N_12425,N_12536);
and U12773 (N_12773,N_12423,N_12552);
and U12774 (N_12774,N_12482,N_12481);
and U12775 (N_12775,N_12522,N_12567);
or U12776 (N_12776,N_12594,N_12549);
nand U12777 (N_12777,N_12460,N_12542);
nand U12778 (N_12778,N_12595,N_12556);
xnor U12779 (N_12779,N_12426,N_12560);
nor U12780 (N_12780,N_12558,N_12490);
or U12781 (N_12781,N_12555,N_12565);
xor U12782 (N_12782,N_12448,N_12553);
and U12783 (N_12783,N_12469,N_12533);
nor U12784 (N_12784,N_12417,N_12448);
and U12785 (N_12785,N_12418,N_12489);
xor U12786 (N_12786,N_12536,N_12591);
nand U12787 (N_12787,N_12496,N_12559);
or U12788 (N_12788,N_12509,N_12553);
xnor U12789 (N_12789,N_12509,N_12434);
nor U12790 (N_12790,N_12598,N_12574);
and U12791 (N_12791,N_12496,N_12408);
nand U12792 (N_12792,N_12462,N_12506);
or U12793 (N_12793,N_12540,N_12488);
nand U12794 (N_12794,N_12546,N_12540);
or U12795 (N_12795,N_12420,N_12498);
xnor U12796 (N_12796,N_12524,N_12577);
or U12797 (N_12797,N_12574,N_12418);
and U12798 (N_12798,N_12469,N_12523);
nand U12799 (N_12799,N_12538,N_12539);
and U12800 (N_12800,N_12798,N_12736);
and U12801 (N_12801,N_12719,N_12694);
and U12802 (N_12802,N_12684,N_12771);
xnor U12803 (N_12803,N_12784,N_12654);
or U12804 (N_12804,N_12650,N_12613);
and U12805 (N_12805,N_12661,N_12738);
and U12806 (N_12806,N_12621,N_12689);
xor U12807 (N_12807,N_12646,N_12769);
or U12808 (N_12808,N_12751,N_12609);
nand U12809 (N_12809,N_12634,N_12705);
xor U12810 (N_12810,N_12747,N_12628);
and U12811 (N_12811,N_12642,N_12753);
nor U12812 (N_12812,N_12627,N_12727);
and U12813 (N_12813,N_12795,N_12778);
nand U12814 (N_12814,N_12721,N_12725);
or U12815 (N_12815,N_12764,N_12672);
and U12816 (N_12816,N_12787,N_12611);
nand U12817 (N_12817,N_12712,N_12757);
and U12818 (N_12818,N_12639,N_12667);
nand U12819 (N_12819,N_12754,N_12765);
or U12820 (N_12820,N_12700,N_12744);
or U12821 (N_12821,N_12709,N_12641);
nand U12822 (N_12822,N_12732,N_12624);
nor U12823 (N_12823,N_12691,N_12740);
and U12824 (N_12824,N_12663,N_12723);
nor U12825 (N_12825,N_12632,N_12671);
or U12826 (N_12826,N_12640,N_12616);
or U12827 (N_12827,N_12713,N_12633);
nor U12828 (N_12828,N_12733,N_12674);
or U12829 (N_12829,N_12786,N_12707);
and U12830 (N_12830,N_12711,N_12706);
nand U12831 (N_12831,N_12749,N_12734);
and U12832 (N_12832,N_12750,N_12683);
or U12833 (N_12833,N_12767,N_12729);
xnor U12834 (N_12834,N_12682,N_12792);
or U12835 (N_12835,N_12741,N_12715);
nand U12836 (N_12836,N_12619,N_12657);
and U12837 (N_12837,N_12755,N_12653);
xnor U12838 (N_12838,N_12791,N_12774);
and U12839 (N_12839,N_12612,N_12703);
and U12840 (N_12840,N_12745,N_12673);
xnor U12841 (N_12841,N_12600,N_12796);
or U12842 (N_12842,N_12675,N_12676);
and U12843 (N_12843,N_12680,N_12759);
or U12844 (N_12844,N_12763,N_12724);
nor U12845 (N_12845,N_12647,N_12697);
nor U12846 (N_12846,N_12776,N_12644);
or U12847 (N_12847,N_12752,N_12625);
xor U12848 (N_12848,N_12690,N_12766);
xor U12849 (N_12849,N_12716,N_12743);
or U12850 (N_12850,N_12665,N_12620);
xnor U12851 (N_12851,N_12636,N_12678);
or U12852 (N_12852,N_12652,N_12735);
and U12853 (N_12853,N_12702,N_12748);
nor U12854 (N_12854,N_12722,N_12648);
nand U12855 (N_12855,N_12658,N_12762);
xnor U12856 (N_12856,N_12651,N_12622);
nor U12857 (N_12857,N_12602,N_12629);
or U12858 (N_12858,N_12742,N_12617);
nor U12859 (N_12859,N_12699,N_12794);
or U12860 (N_12860,N_12758,N_12601);
nor U12861 (N_12861,N_12698,N_12696);
and U12862 (N_12862,N_12614,N_12788);
or U12863 (N_12863,N_12693,N_12610);
nor U12864 (N_12864,N_12685,N_12710);
nor U12865 (N_12865,N_12679,N_12789);
or U12866 (N_12866,N_12649,N_12777);
or U12867 (N_12867,N_12793,N_12605);
and U12868 (N_12868,N_12688,N_12692);
xnor U12869 (N_12869,N_12608,N_12643);
or U12870 (N_12870,N_12714,N_12645);
xor U12871 (N_12871,N_12677,N_12604);
nand U12872 (N_12872,N_12772,N_12607);
nand U12873 (N_12873,N_12695,N_12780);
nand U12874 (N_12874,N_12668,N_12701);
and U12875 (N_12875,N_12664,N_12618);
or U12876 (N_12876,N_12718,N_12662);
nor U12877 (N_12877,N_12631,N_12785);
xor U12878 (N_12878,N_12708,N_12756);
nor U12879 (N_12879,N_12730,N_12635);
xor U12880 (N_12880,N_12775,N_12681);
and U12881 (N_12881,N_12660,N_12773);
xor U12882 (N_12882,N_12687,N_12728);
xor U12883 (N_12883,N_12746,N_12603);
nor U12884 (N_12884,N_12656,N_12781);
nand U12885 (N_12885,N_12626,N_12630);
nand U12886 (N_12886,N_12638,N_12739);
and U12887 (N_12887,N_12726,N_12770);
and U12888 (N_12888,N_12615,N_12637);
and U12889 (N_12889,N_12606,N_12704);
nand U12890 (N_12890,N_12737,N_12670);
or U12891 (N_12891,N_12666,N_12779);
and U12892 (N_12892,N_12797,N_12761);
or U12893 (N_12893,N_12782,N_12720);
or U12894 (N_12894,N_12717,N_12760);
nand U12895 (N_12895,N_12783,N_12790);
nor U12896 (N_12896,N_12655,N_12686);
nor U12897 (N_12897,N_12799,N_12623);
and U12898 (N_12898,N_12731,N_12669);
nand U12899 (N_12899,N_12659,N_12768);
and U12900 (N_12900,N_12627,N_12689);
nor U12901 (N_12901,N_12799,N_12706);
nor U12902 (N_12902,N_12630,N_12770);
and U12903 (N_12903,N_12669,N_12624);
or U12904 (N_12904,N_12731,N_12787);
or U12905 (N_12905,N_12697,N_12756);
nor U12906 (N_12906,N_12719,N_12780);
and U12907 (N_12907,N_12645,N_12619);
and U12908 (N_12908,N_12653,N_12671);
nand U12909 (N_12909,N_12655,N_12762);
nand U12910 (N_12910,N_12700,N_12786);
xnor U12911 (N_12911,N_12618,N_12658);
and U12912 (N_12912,N_12779,N_12736);
or U12913 (N_12913,N_12699,N_12686);
or U12914 (N_12914,N_12657,N_12648);
or U12915 (N_12915,N_12649,N_12695);
nor U12916 (N_12916,N_12745,N_12601);
or U12917 (N_12917,N_12749,N_12700);
and U12918 (N_12918,N_12663,N_12669);
and U12919 (N_12919,N_12653,N_12739);
xor U12920 (N_12920,N_12714,N_12610);
and U12921 (N_12921,N_12690,N_12760);
or U12922 (N_12922,N_12721,N_12773);
or U12923 (N_12923,N_12624,N_12799);
xor U12924 (N_12924,N_12619,N_12670);
and U12925 (N_12925,N_12699,N_12677);
and U12926 (N_12926,N_12683,N_12641);
nor U12927 (N_12927,N_12711,N_12677);
and U12928 (N_12928,N_12781,N_12738);
nor U12929 (N_12929,N_12617,N_12759);
nand U12930 (N_12930,N_12744,N_12787);
xor U12931 (N_12931,N_12700,N_12717);
nor U12932 (N_12932,N_12672,N_12678);
and U12933 (N_12933,N_12733,N_12697);
nor U12934 (N_12934,N_12796,N_12715);
nor U12935 (N_12935,N_12793,N_12661);
xor U12936 (N_12936,N_12752,N_12664);
nor U12937 (N_12937,N_12737,N_12723);
nor U12938 (N_12938,N_12676,N_12727);
or U12939 (N_12939,N_12779,N_12777);
nand U12940 (N_12940,N_12636,N_12719);
xnor U12941 (N_12941,N_12722,N_12750);
or U12942 (N_12942,N_12745,N_12699);
nand U12943 (N_12943,N_12696,N_12739);
xor U12944 (N_12944,N_12670,N_12685);
xnor U12945 (N_12945,N_12749,N_12747);
nor U12946 (N_12946,N_12601,N_12772);
or U12947 (N_12947,N_12724,N_12752);
or U12948 (N_12948,N_12789,N_12652);
xnor U12949 (N_12949,N_12666,N_12725);
and U12950 (N_12950,N_12780,N_12777);
and U12951 (N_12951,N_12743,N_12656);
and U12952 (N_12952,N_12772,N_12738);
nor U12953 (N_12953,N_12681,N_12759);
nand U12954 (N_12954,N_12658,N_12683);
and U12955 (N_12955,N_12737,N_12780);
nor U12956 (N_12956,N_12737,N_12658);
nor U12957 (N_12957,N_12676,N_12654);
nor U12958 (N_12958,N_12789,N_12616);
and U12959 (N_12959,N_12651,N_12743);
nand U12960 (N_12960,N_12663,N_12729);
or U12961 (N_12961,N_12765,N_12744);
or U12962 (N_12962,N_12621,N_12725);
nor U12963 (N_12963,N_12674,N_12662);
nor U12964 (N_12964,N_12702,N_12627);
or U12965 (N_12965,N_12727,N_12635);
xnor U12966 (N_12966,N_12652,N_12613);
and U12967 (N_12967,N_12696,N_12700);
and U12968 (N_12968,N_12640,N_12615);
nand U12969 (N_12969,N_12795,N_12639);
nor U12970 (N_12970,N_12741,N_12636);
and U12971 (N_12971,N_12734,N_12608);
nand U12972 (N_12972,N_12719,N_12687);
or U12973 (N_12973,N_12635,N_12691);
and U12974 (N_12974,N_12608,N_12659);
xor U12975 (N_12975,N_12606,N_12772);
xnor U12976 (N_12976,N_12605,N_12762);
and U12977 (N_12977,N_12644,N_12786);
xnor U12978 (N_12978,N_12767,N_12758);
nor U12979 (N_12979,N_12738,N_12634);
nor U12980 (N_12980,N_12660,N_12751);
nand U12981 (N_12981,N_12776,N_12627);
xnor U12982 (N_12982,N_12780,N_12735);
xor U12983 (N_12983,N_12685,N_12752);
or U12984 (N_12984,N_12726,N_12685);
nor U12985 (N_12985,N_12780,N_12715);
or U12986 (N_12986,N_12793,N_12705);
xnor U12987 (N_12987,N_12704,N_12727);
nor U12988 (N_12988,N_12645,N_12667);
nor U12989 (N_12989,N_12645,N_12675);
nand U12990 (N_12990,N_12779,N_12707);
nand U12991 (N_12991,N_12635,N_12673);
nand U12992 (N_12992,N_12620,N_12614);
xor U12993 (N_12993,N_12795,N_12711);
or U12994 (N_12994,N_12766,N_12765);
nor U12995 (N_12995,N_12768,N_12681);
nor U12996 (N_12996,N_12678,N_12601);
nand U12997 (N_12997,N_12700,N_12707);
nand U12998 (N_12998,N_12698,N_12707);
nor U12999 (N_12999,N_12668,N_12694);
xor U13000 (N_13000,N_12892,N_12941);
nor U13001 (N_13001,N_12928,N_12825);
nand U13002 (N_13002,N_12979,N_12803);
xnor U13003 (N_13003,N_12809,N_12867);
nor U13004 (N_13004,N_12985,N_12870);
or U13005 (N_13005,N_12991,N_12893);
or U13006 (N_13006,N_12835,N_12926);
nor U13007 (N_13007,N_12831,N_12869);
or U13008 (N_13008,N_12921,N_12883);
nor U13009 (N_13009,N_12800,N_12833);
xnor U13010 (N_13010,N_12801,N_12912);
nand U13011 (N_13011,N_12992,N_12860);
nand U13012 (N_13012,N_12842,N_12838);
and U13013 (N_13013,N_12956,N_12876);
and U13014 (N_13014,N_12938,N_12850);
nand U13015 (N_13015,N_12899,N_12964);
xnor U13016 (N_13016,N_12861,N_12829);
or U13017 (N_13017,N_12816,N_12874);
and U13018 (N_13018,N_12868,N_12898);
nor U13019 (N_13019,N_12837,N_12997);
nand U13020 (N_13020,N_12887,N_12931);
nand U13021 (N_13021,N_12966,N_12805);
or U13022 (N_13022,N_12836,N_12970);
xor U13023 (N_13023,N_12902,N_12946);
nor U13024 (N_13024,N_12895,N_12917);
or U13025 (N_13025,N_12882,N_12986);
nand U13026 (N_13026,N_12952,N_12930);
nor U13027 (N_13027,N_12854,N_12989);
xor U13028 (N_13028,N_12936,N_12821);
or U13029 (N_13029,N_12859,N_12840);
xnor U13030 (N_13030,N_12843,N_12885);
nand U13031 (N_13031,N_12954,N_12958);
nor U13032 (N_13032,N_12851,N_12877);
and U13033 (N_13033,N_12819,N_12813);
or U13034 (N_13034,N_12848,N_12914);
and U13035 (N_13035,N_12897,N_12967);
or U13036 (N_13036,N_12804,N_12849);
xor U13037 (N_13037,N_12891,N_12965);
nand U13038 (N_13038,N_12846,N_12910);
nor U13039 (N_13039,N_12960,N_12920);
nor U13040 (N_13040,N_12904,N_12820);
and U13041 (N_13041,N_12907,N_12886);
nor U13042 (N_13042,N_12969,N_12839);
nor U13043 (N_13043,N_12934,N_12915);
nor U13044 (N_13044,N_12929,N_12943);
xor U13045 (N_13045,N_12865,N_12890);
or U13046 (N_13046,N_12974,N_12913);
nor U13047 (N_13047,N_12932,N_12852);
nor U13048 (N_13048,N_12900,N_12808);
xor U13049 (N_13049,N_12984,N_12949);
nand U13050 (N_13050,N_12968,N_12948);
xnor U13051 (N_13051,N_12935,N_12975);
and U13052 (N_13052,N_12944,N_12995);
nand U13053 (N_13053,N_12845,N_12810);
and U13054 (N_13054,N_12872,N_12866);
xnor U13055 (N_13055,N_12828,N_12862);
xnor U13056 (N_13056,N_12863,N_12924);
or U13057 (N_13057,N_12972,N_12856);
or U13058 (N_13058,N_12918,N_12812);
nor U13059 (N_13059,N_12871,N_12841);
xnor U13060 (N_13060,N_12853,N_12879);
nor U13061 (N_13061,N_12971,N_12880);
or U13062 (N_13062,N_12977,N_12806);
xnor U13063 (N_13063,N_12826,N_12927);
nand U13064 (N_13064,N_12888,N_12951);
nand U13065 (N_13065,N_12978,N_12981);
nor U13066 (N_13066,N_12873,N_12996);
nor U13067 (N_13067,N_12823,N_12802);
nand U13068 (N_13068,N_12909,N_12963);
or U13069 (N_13069,N_12844,N_12811);
or U13070 (N_13070,N_12940,N_12994);
or U13071 (N_13071,N_12822,N_12933);
and U13072 (N_13072,N_12947,N_12824);
xor U13073 (N_13073,N_12923,N_12896);
nand U13074 (N_13074,N_12942,N_12911);
and U13075 (N_13075,N_12999,N_12864);
and U13076 (N_13076,N_12959,N_12827);
or U13077 (N_13077,N_12919,N_12906);
and U13078 (N_13078,N_12973,N_12957);
nor U13079 (N_13079,N_12855,N_12884);
or U13080 (N_13080,N_12807,N_12818);
and U13081 (N_13081,N_12953,N_12987);
nand U13082 (N_13082,N_12905,N_12814);
nand U13083 (N_13083,N_12939,N_12815);
nor U13084 (N_13084,N_12908,N_12830);
xnor U13085 (N_13085,N_12982,N_12955);
xor U13086 (N_13086,N_12903,N_12901);
nand U13087 (N_13087,N_12878,N_12834);
and U13088 (N_13088,N_12857,N_12998);
and U13089 (N_13089,N_12980,N_12962);
xor U13090 (N_13090,N_12983,N_12925);
and U13091 (N_13091,N_12993,N_12945);
and U13092 (N_13092,N_12937,N_12875);
xnor U13093 (N_13093,N_12832,N_12922);
nor U13094 (N_13094,N_12858,N_12990);
and U13095 (N_13095,N_12847,N_12988);
or U13096 (N_13096,N_12916,N_12881);
nor U13097 (N_13097,N_12961,N_12817);
and U13098 (N_13098,N_12894,N_12950);
nor U13099 (N_13099,N_12976,N_12889);
xnor U13100 (N_13100,N_12945,N_12870);
nand U13101 (N_13101,N_12809,N_12876);
nor U13102 (N_13102,N_12904,N_12969);
xnor U13103 (N_13103,N_12883,N_12985);
or U13104 (N_13104,N_12923,N_12801);
or U13105 (N_13105,N_12933,N_12924);
or U13106 (N_13106,N_12904,N_12810);
and U13107 (N_13107,N_12881,N_12899);
nand U13108 (N_13108,N_12843,N_12986);
or U13109 (N_13109,N_12828,N_12968);
and U13110 (N_13110,N_12969,N_12821);
xor U13111 (N_13111,N_12864,N_12877);
or U13112 (N_13112,N_12892,N_12856);
xor U13113 (N_13113,N_12942,N_12997);
and U13114 (N_13114,N_12866,N_12960);
and U13115 (N_13115,N_12818,N_12906);
nand U13116 (N_13116,N_12900,N_12978);
and U13117 (N_13117,N_12982,N_12939);
and U13118 (N_13118,N_12871,N_12913);
nand U13119 (N_13119,N_12885,N_12951);
or U13120 (N_13120,N_12997,N_12816);
nand U13121 (N_13121,N_12913,N_12846);
nor U13122 (N_13122,N_12802,N_12990);
xor U13123 (N_13123,N_12921,N_12938);
or U13124 (N_13124,N_12905,N_12902);
nor U13125 (N_13125,N_12817,N_12922);
xor U13126 (N_13126,N_12923,N_12867);
nand U13127 (N_13127,N_12864,N_12870);
nor U13128 (N_13128,N_12932,N_12839);
or U13129 (N_13129,N_12961,N_12913);
nor U13130 (N_13130,N_12995,N_12830);
and U13131 (N_13131,N_12995,N_12971);
nand U13132 (N_13132,N_12820,N_12864);
or U13133 (N_13133,N_12853,N_12990);
xor U13134 (N_13134,N_12959,N_12991);
and U13135 (N_13135,N_12853,N_12900);
and U13136 (N_13136,N_12990,N_12810);
nor U13137 (N_13137,N_12961,N_12975);
and U13138 (N_13138,N_12898,N_12801);
nand U13139 (N_13139,N_12835,N_12881);
and U13140 (N_13140,N_12929,N_12966);
xnor U13141 (N_13141,N_12896,N_12911);
or U13142 (N_13142,N_12945,N_12885);
or U13143 (N_13143,N_12898,N_12981);
or U13144 (N_13144,N_12833,N_12992);
nor U13145 (N_13145,N_12900,N_12855);
xnor U13146 (N_13146,N_12937,N_12979);
or U13147 (N_13147,N_12926,N_12967);
nor U13148 (N_13148,N_12806,N_12821);
xor U13149 (N_13149,N_12937,N_12954);
xnor U13150 (N_13150,N_12986,N_12947);
and U13151 (N_13151,N_12986,N_12894);
nand U13152 (N_13152,N_12975,N_12973);
nor U13153 (N_13153,N_12866,N_12890);
or U13154 (N_13154,N_12971,N_12879);
or U13155 (N_13155,N_12993,N_12965);
and U13156 (N_13156,N_12963,N_12990);
nand U13157 (N_13157,N_12996,N_12833);
nor U13158 (N_13158,N_12861,N_12969);
nor U13159 (N_13159,N_12809,N_12934);
xor U13160 (N_13160,N_12840,N_12968);
xor U13161 (N_13161,N_12965,N_12937);
or U13162 (N_13162,N_12843,N_12873);
or U13163 (N_13163,N_12973,N_12803);
xnor U13164 (N_13164,N_12829,N_12855);
nand U13165 (N_13165,N_12899,N_12810);
and U13166 (N_13166,N_12836,N_12837);
xor U13167 (N_13167,N_12918,N_12910);
or U13168 (N_13168,N_12833,N_12955);
nor U13169 (N_13169,N_12822,N_12985);
xnor U13170 (N_13170,N_12878,N_12842);
nor U13171 (N_13171,N_12839,N_12940);
nand U13172 (N_13172,N_12851,N_12926);
nand U13173 (N_13173,N_12992,N_12994);
xnor U13174 (N_13174,N_12880,N_12853);
or U13175 (N_13175,N_12872,N_12940);
xnor U13176 (N_13176,N_12949,N_12985);
and U13177 (N_13177,N_12995,N_12840);
xor U13178 (N_13178,N_12862,N_12838);
and U13179 (N_13179,N_12856,N_12982);
nand U13180 (N_13180,N_12983,N_12914);
nor U13181 (N_13181,N_12961,N_12825);
or U13182 (N_13182,N_12837,N_12975);
nor U13183 (N_13183,N_12953,N_12977);
or U13184 (N_13184,N_12862,N_12891);
and U13185 (N_13185,N_12989,N_12807);
and U13186 (N_13186,N_12811,N_12803);
xnor U13187 (N_13187,N_12950,N_12882);
nor U13188 (N_13188,N_12997,N_12960);
nand U13189 (N_13189,N_12835,N_12830);
nand U13190 (N_13190,N_12892,N_12827);
and U13191 (N_13191,N_12933,N_12956);
and U13192 (N_13192,N_12822,N_12998);
nand U13193 (N_13193,N_12887,N_12888);
or U13194 (N_13194,N_12923,N_12837);
nand U13195 (N_13195,N_12819,N_12947);
and U13196 (N_13196,N_12808,N_12902);
and U13197 (N_13197,N_12865,N_12834);
or U13198 (N_13198,N_12892,N_12922);
nor U13199 (N_13199,N_12959,N_12924);
nor U13200 (N_13200,N_13163,N_13114);
or U13201 (N_13201,N_13112,N_13030);
or U13202 (N_13202,N_13170,N_13109);
nor U13203 (N_13203,N_13049,N_13097);
and U13204 (N_13204,N_13015,N_13157);
and U13205 (N_13205,N_13037,N_13003);
or U13206 (N_13206,N_13180,N_13052);
xnor U13207 (N_13207,N_13048,N_13077);
nor U13208 (N_13208,N_13140,N_13043);
and U13209 (N_13209,N_13176,N_13073);
and U13210 (N_13210,N_13064,N_13158);
or U13211 (N_13211,N_13034,N_13189);
or U13212 (N_13212,N_13136,N_13104);
xnor U13213 (N_13213,N_13022,N_13094);
nand U13214 (N_13214,N_13076,N_13081);
or U13215 (N_13215,N_13124,N_13012);
nand U13216 (N_13216,N_13070,N_13035);
and U13217 (N_13217,N_13145,N_13149);
nand U13218 (N_13218,N_13010,N_13053);
or U13219 (N_13219,N_13093,N_13131);
xor U13220 (N_13220,N_13181,N_13006);
nand U13221 (N_13221,N_13045,N_13100);
and U13222 (N_13222,N_13166,N_13126);
nand U13223 (N_13223,N_13067,N_13001);
nand U13224 (N_13224,N_13098,N_13167);
nor U13225 (N_13225,N_13085,N_13113);
and U13226 (N_13226,N_13177,N_13080);
or U13227 (N_13227,N_13123,N_13040);
nor U13228 (N_13228,N_13134,N_13032);
xnor U13229 (N_13229,N_13150,N_13153);
nand U13230 (N_13230,N_13156,N_13074);
and U13231 (N_13231,N_13143,N_13106);
or U13232 (N_13232,N_13091,N_13054);
nand U13233 (N_13233,N_13146,N_13172);
and U13234 (N_13234,N_13198,N_13063);
nor U13235 (N_13235,N_13026,N_13038);
and U13236 (N_13236,N_13033,N_13041);
nand U13237 (N_13237,N_13116,N_13023);
nor U13238 (N_13238,N_13118,N_13155);
and U13239 (N_13239,N_13183,N_13174);
and U13240 (N_13240,N_13028,N_13092);
xnor U13241 (N_13241,N_13182,N_13195);
or U13242 (N_13242,N_13083,N_13152);
or U13243 (N_13243,N_13193,N_13161);
or U13244 (N_13244,N_13141,N_13095);
nor U13245 (N_13245,N_13160,N_13105);
and U13246 (N_13246,N_13059,N_13039);
nor U13247 (N_13247,N_13154,N_13197);
nand U13248 (N_13248,N_13187,N_13107);
nand U13249 (N_13249,N_13178,N_13191);
or U13250 (N_13250,N_13021,N_13142);
nor U13251 (N_13251,N_13108,N_13016);
xnor U13252 (N_13252,N_13027,N_13075);
and U13253 (N_13253,N_13065,N_13139);
and U13254 (N_13254,N_13007,N_13014);
xnor U13255 (N_13255,N_13057,N_13066);
xor U13256 (N_13256,N_13084,N_13137);
or U13257 (N_13257,N_13068,N_13175);
nand U13258 (N_13258,N_13096,N_13024);
nand U13259 (N_13259,N_13044,N_13078);
nor U13260 (N_13260,N_13121,N_13151);
nand U13261 (N_13261,N_13031,N_13135);
nor U13262 (N_13262,N_13060,N_13162);
nor U13263 (N_13263,N_13088,N_13199);
xor U13264 (N_13264,N_13058,N_13055);
and U13265 (N_13265,N_13130,N_13000);
and U13266 (N_13266,N_13169,N_13050);
and U13267 (N_13267,N_13129,N_13046);
nand U13268 (N_13268,N_13103,N_13190);
and U13269 (N_13269,N_13029,N_13013);
nand U13270 (N_13270,N_13144,N_13062);
and U13271 (N_13271,N_13079,N_13019);
and U13272 (N_13272,N_13165,N_13099);
or U13273 (N_13273,N_13017,N_13005);
and U13274 (N_13274,N_13072,N_13011);
and U13275 (N_13275,N_13002,N_13008);
nand U13276 (N_13276,N_13087,N_13186);
nor U13277 (N_13277,N_13061,N_13082);
and U13278 (N_13278,N_13125,N_13171);
or U13279 (N_13279,N_13122,N_13133);
nand U13280 (N_13280,N_13117,N_13025);
nand U13281 (N_13281,N_13119,N_13089);
nand U13282 (N_13282,N_13090,N_13128);
nand U13283 (N_13283,N_13168,N_13159);
and U13284 (N_13284,N_13110,N_13196);
nand U13285 (N_13285,N_13069,N_13148);
nor U13286 (N_13286,N_13132,N_13086);
nor U13287 (N_13287,N_13179,N_13185);
and U13288 (N_13288,N_13036,N_13138);
xor U13289 (N_13289,N_13047,N_13127);
and U13290 (N_13290,N_13164,N_13004);
nand U13291 (N_13291,N_13009,N_13120);
nor U13292 (N_13292,N_13071,N_13115);
or U13293 (N_13293,N_13102,N_13056);
or U13294 (N_13294,N_13188,N_13184);
xor U13295 (N_13295,N_13051,N_13111);
nor U13296 (N_13296,N_13018,N_13101);
nand U13297 (N_13297,N_13020,N_13042);
xnor U13298 (N_13298,N_13147,N_13192);
nand U13299 (N_13299,N_13194,N_13173);
nand U13300 (N_13300,N_13071,N_13092);
nand U13301 (N_13301,N_13058,N_13173);
xnor U13302 (N_13302,N_13150,N_13066);
nand U13303 (N_13303,N_13193,N_13090);
nor U13304 (N_13304,N_13063,N_13157);
or U13305 (N_13305,N_13147,N_13177);
and U13306 (N_13306,N_13132,N_13051);
or U13307 (N_13307,N_13022,N_13167);
xnor U13308 (N_13308,N_13084,N_13046);
nor U13309 (N_13309,N_13037,N_13036);
xnor U13310 (N_13310,N_13056,N_13121);
or U13311 (N_13311,N_13100,N_13044);
and U13312 (N_13312,N_13158,N_13087);
and U13313 (N_13313,N_13056,N_13067);
or U13314 (N_13314,N_13007,N_13029);
nor U13315 (N_13315,N_13037,N_13034);
or U13316 (N_13316,N_13105,N_13003);
xor U13317 (N_13317,N_13005,N_13097);
nor U13318 (N_13318,N_13033,N_13005);
and U13319 (N_13319,N_13188,N_13077);
and U13320 (N_13320,N_13177,N_13130);
or U13321 (N_13321,N_13014,N_13024);
nand U13322 (N_13322,N_13000,N_13149);
xor U13323 (N_13323,N_13034,N_13169);
xnor U13324 (N_13324,N_13161,N_13098);
or U13325 (N_13325,N_13111,N_13008);
and U13326 (N_13326,N_13100,N_13030);
nand U13327 (N_13327,N_13092,N_13099);
nand U13328 (N_13328,N_13094,N_13037);
nand U13329 (N_13329,N_13080,N_13091);
and U13330 (N_13330,N_13199,N_13024);
nor U13331 (N_13331,N_13017,N_13062);
nor U13332 (N_13332,N_13093,N_13103);
or U13333 (N_13333,N_13130,N_13002);
and U13334 (N_13334,N_13122,N_13149);
nand U13335 (N_13335,N_13075,N_13085);
nor U13336 (N_13336,N_13106,N_13160);
nand U13337 (N_13337,N_13125,N_13043);
and U13338 (N_13338,N_13054,N_13052);
and U13339 (N_13339,N_13165,N_13011);
and U13340 (N_13340,N_13196,N_13042);
or U13341 (N_13341,N_13068,N_13106);
and U13342 (N_13342,N_13177,N_13167);
nand U13343 (N_13343,N_13117,N_13068);
and U13344 (N_13344,N_13142,N_13026);
or U13345 (N_13345,N_13011,N_13144);
or U13346 (N_13346,N_13149,N_13123);
nand U13347 (N_13347,N_13155,N_13083);
nor U13348 (N_13348,N_13149,N_13052);
nand U13349 (N_13349,N_13025,N_13087);
and U13350 (N_13350,N_13032,N_13000);
nand U13351 (N_13351,N_13041,N_13167);
or U13352 (N_13352,N_13087,N_13003);
xor U13353 (N_13353,N_13042,N_13074);
nand U13354 (N_13354,N_13074,N_13164);
xnor U13355 (N_13355,N_13010,N_13047);
xor U13356 (N_13356,N_13195,N_13174);
nand U13357 (N_13357,N_13114,N_13066);
or U13358 (N_13358,N_13003,N_13022);
nand U13359 (N_13359,N_13163,N_13093);
xor U13360 (N_13360,N_13167,N_13009);
and U13361 (N_13361,N_13177,N_13081);
or U13362 (N_13362,N_13018,N_13092);
and U13363 (N_13363,N_13195,N_13156);
or U13364 (N_13364,N_13074,N_13178);
nand U13365 (N_13365,N_13195,N_13172);
nor U13366 (N_13366,N_13018,N_13185);
nand U13367 (N_13367,N_13174,N_13086);
xnor U13368 (N_13368,N_13007,N_13172);
nor U13369 (N_13369,N_13162,N_13043);
nor U13370 (N_13370,N_13045,N_13152);
xnor U13371 (N_13371,N_13093,N_13065);
nor U13372 (N_13372,N_13083,N_13150);
xnor U13373 (N_13373,N_13078,N_13048);
xor U13374 (N_13374,N_13121,N_13023);
and U13375 (N_13375,N_13035,N_13110);
nor U13376 (N_13376,N_13185,N_13000);
nand U13377 (N_13377,N_13048,N_13132);
nand U13378 (N_13378,N_13079,N_13052);
xnor U13379 (N_13379,N_13101,N_13187);
or U13380 (N_13380,N_13147,N_13055);
xnor U13381 (N_13381,N_13178,N_13032);
or U13382 (N_13382,N_13135,N_13090);
or U13383 (N_13383,N_13168,N_13082);
xnor U13384 (N_13384,N_13150,N_13019);
or U13385 (N_13385,N_13188,N_13024);
nor U13386 (N_13386,N_13176,N_13015);
nor U13387 (N_13387,N_13155,N_13015);
and U13388 (N_13388,N_13113,N_13114);
xor U13389 (N_13389,N_13104,N_13172);
and U13390 (N_13390,N_13098,N_13122);
xor U13391 (N_13391,N_13024,N_13166);
or U13392 (N_13392,N_13187,N_13165);
or U13393 (N_13393,N_13062,N_13042);
nand U13394 (N_13394,N_13143,N_13059);
nand U13395 (N_13395,N_13080,N_13142);
or U13396 (N_13396,N_13032,N_13001);
or U13397 (N_13397,N_13006,N_13140);
and U13398 (N_13398,N_13024,N_13026);
nor U13399 (N_13399,N_13095,N_13074);
nor U13400 (N_13400,N_13319,N_13266);
and U13401 (N_13401,N_13343,N_13308);
or U13402 (N_13402,N_13248,N_13390);
and U13403 (N_13403,N_13225,N_13320);
nor U13404 (N_13404,N_13312,N_13217);
or U13405 (N_13405,N_13322,N_13286);
nor U13406 (N_13406,N_13384,N_13282);
nand U13407 (N_13407,N_13336,N_13358);
nor U13408 (N_13408,N_13380,N_13270);
and U13409 (N_13409,N_13366,N_13246);
nor U13410 (N_13410,N_13351,N_13313);
nor U13411 (N_13411,N_13391,N_13207);
nor U13412 (N_13412,N_13259,N_13284);
xnor U13413 (N_13413,N_13359,N_13298);
and U13414 (N_13414,N_13299,N_13377);
and U13415 (N_13415,N_13360,N_13334);
nor U13416 (N_13416,N_13387,N_13317);
and U13417 (N_13417,N_13382,N_13329);
and U13418 (N_13418,N_13353,N_13311);
or U13419 (N_13419,N_13243,N_13200);
nor U13420 (N_13420,N_13350,N_13293);
nor U13421 (N_13421,N_13258,N_13242);
nor U13422 (N_13422,N_13237,N_13279);
xnor U13423 (N_13423,N_13398,N_13328);
nand U13424 (N_13424,N_13345,N_13367);
or U13425 (N_13425,N_13342,N_13307);
or U13426 (N_13426,N_13295,N_13208);
nor U13427 (N_13427,N_13302,N_13327);
xnor U13428 (N_13428,N_13333,N_13206);
and U13429 (N_13429,N_13362,N_13203);
or U13430 (N_13430,N_13238,N_13300);
nand U13431 (N_13431,N_13253,N_13277);
nand U13432 (N_13432,N_13297,N_13287);
and U13433 (N_13433,N_13271,N_13230);
nand U13434 (N_13434,N_13325,N_13304);
and U13435 (N_13435,N_13249,N_13301);
and U13436 (N_13436,N_13397,N_13318);
nor U13437 (N_13437,N_13372,N_13370);
nand U13438 (N_13438,N_13375,N_13252);
nand U13439 (N_13439,N_13289,N_13294);
xor U13440 (N_13440,N_13251,N_13264);
nor U13441 (N_13441,N_13232,N_13393);
or U13442 (N_13442,N_13261,N_13234);
nor U13443 (N_13443,N_13202,N_13278);
or U13444 (N_13444,N_13290,N_13226);
nand U13445 (N_13445,N_13247,N_13254);
xor U13446 (N_13446,N_13223,N_13315);
nor U13447 (N_13447,N_13354,N_13331);
nor U13448 (N_13448,N_13385,N_13386);
and U13449 (N_13449,N_13235,N_13396);
nor U13450 (N_13450,N_13292,N_13296);
nand U13451 (N_13451,N_13369,N_13352);
nand U13452 (N_13452,N_13365,N_13240);
and U13453 (N_13453,N_13269,N_13285);
xnor U13454 (N_13454,N_13273,N_13337);
nor U13455 (N_13455,N_13291,N_13338);
xnor U13456 (N_13456,N_13250,N_13321);
or U13457 (N_13457,N_13229,N_13383);
nor U13458 (N_13458,N_13378,N_13257);
xnor U13459 (N_13459,N_13316,N_13389);
nor U13460 (N_13460,N_13205,N_13239);
nor U13461 (N_13461,N_13394,N_13222);
xor U13462 (N_13462,N_13262,N_13233);
nand U13463 (N_13463,N_13283,N_13255);
xnor U13464 (N_13464,N_13218,N_13212);
or U13465 (N_13465,N_13306,N_13310);
xor U13466 (N_13466,N_13215,N_13260);
or U13467 (N_13467,N_13355,N_13267);
nand U13468 (N_13468,N_13373,N_13201);
and U13469 (N_13469,N_13280,N_13341);
and U13470 (N_13470,N_13347,N_13231);
and U13471 (N_13471,N_13241,N_13314);
and U13472 (N_13472,N_13213,N_13346);
or U13473 (N_13473,N_13356,N_13395);
nor U13474 (N_13474,N_13348,N_13281);
or U13475 (N_13475,N_13276,N_13349);
xnor U13476 (N_13476,N_13228,N_13361);
nor U13477 (N_13477,N_13244,N_13274);
nor U13478 (N_13478,N_13357,N_13335);
nand U13479 (N_13479,N_13209,N_13275);
or U13480 (N_13480,N_13392,N_13268);
and U13481 (N_13481,N_13363,N_13371);
or U13482 (N_13482,N_13210,N_13256);
or U13483 (N_13483,N_13379,N_13344);
or U13484 (N_13484,N_13265,N_13221);
nand U13485 (N_13485,N_13303,N_13211);
or U13486 (N_13486,N_13339,N_13340);
nand U13487 (N_13487,N_13381,N_13374);
xnor U13488 (N_13488,N_13263,N_13368);
nand U13489 (N_13489,N_13227,N_13305);
xor U13490 (N_13490,N_13204,N_13216);
nor U13491 (N_13491,N_13245,N_13323);
and U13492 (N_13492,N_13214,N_13220);
xor U13493 (N_13493,N_13309,N_13376);
or U13494 (N_13494,N_13272,N_13288);
and U13495 (N_13495,N_13324,N_13332);
nor U13496 (N_13496,N_13399,N_13330);
nor U13497 (N_13497,N_13364,N_13326);
and U13498 (N_13498,N_13219,N_13224);
or U13499 (N_13499,N_13388,N_13236);
xnor U13500 (N_13500,N_13283,N_13300);
or U13501 (N_13501,N_13298,N_13272);
nand U13502 (N_13502,N_13233,N_13325);
xor U13503 (N_13503,N_13242,N_13274);
and U13504 (N_13504,N_13282,N_13320);
xnor U13505 (N_13505,N_13200,N_13373);
nand U13506 (N_13506,N_13360,N_13303);
and U13507 (N_13507,N_13212,N_13309);
nor U13508 (N_13508,N_13391,N_13383);
nand U13509 (N_13509,N_13215,N_13345);
and U13510 (N_13510,N_13333,N_13233);
or U13511 (N_13511,N_13346,N_13317);
nor U13512 (N_13512,N_13236,N_13277);
nor U13513 (N_13513,N_13331,N_13391);
and U13514 (N_13514,N_13325,N_13314);
nand U13515 (N_13515,N_13240,N_13235);
nand U13516 (N_13516,N_13338,N_13202);
xnor U13517 (N_13517,N_13365,N_13353);
xor U13518 (N_13518,N_13241,N_13332);
xnor U13519 (N_13519,N_13369,N_13311);
and U13520 (N_13520,N_13277,N_13258);
or U13521 (N_13521,N_13384,N_13348);
nand U13522 (N_13522,N_13218,N_13237);
nor U13523 (N_13523,N_13356,N_13219);
nand U13524 (N_13524,N_13355,N_13257);
or U13525 (N_13525,N_13239,N_13243);
or U13526 (N_13526,N_13253,N_13222);
nand U13527 (N_13527,N_13345,N_13387);
or U13528 (N_13528,N_13257,N_13281);
and U13529 (N_13529,N_13368,N_13271);
nor U13530 (N_13530,N_13291,N_13289);
or U13531 (N_13531,N_13367,N_13314);
nor U13532 (N_13532,N_13244,N_13228);
and U13533 (N_13533,N_13351,N_13226);
nor U13534 (N_13534,N_13266,N_13262);
or U13535 (N_13535,N_13391,N_13334);
and U13536 (N_13536,N_13266,N_13364);
and U13537 (N_13537,N_13285,N_13257);
or U13538 (N_13538,N_13395,N_13321);
and U13539 (N_13539,N_13345,N_13366);
xnor U13540 (N_13540,N_13327,N_13378);
nor U13541 (N_13541,N_13211,N_13316);
nand U13542 (N_13542,N_13388,N_13288);
xnor U13543 (N_13543,N_13285,N_13376);
and U13544 (N_13544,N_13319,N_13276);
and U13545 (N_13545,N_13233,N_13240);
and U13546 (N_13546,N_13316,N_13266);
xor U13547 (N_13547,N_13218,N_13366);
xnor U13548 (N_13548,N_13232,N_13271);
and U13549 (N_13549,N_13236,N_13385);
xor U13550 (N_13550,N_13298,N_13213);
nor U13551 (N_13551,N_13262,N_13393);
xnor U13552 (N_13552,N_13260,N_13212);
or U13553 (N_13553,N_13276,N_13231);
xnor U13554 (N_13554,N_13214,N_13279);
and U13555 (N_13555,N_13219,N_13373);
nor U13556 (N_13556,N_13270,N_13379);
or U13557 (N_13557,N_13304,N_13323);
or U13558 (N_13558,N_13201,N_13257);
nor U13559 (N_13559,N_13346,N_13292);
or U13560 (N_13560,N_13286,N_13317);
and U13561 (N_13561,N_13372,N_13371);
nand U13562 (N_13562,N_13271,N_13389);
nor U13563 (N_13563,N_13298,N_13212);
xnor U13564 (N_13564,N_13304,N_13246);
and U13565 (N_13565,N_13217,N_13270);
xnor U13566 (N_13566,N_13224,N_13282);
and U13567 (N_13567,N_13398,N_13229);
nand U13568 (N_13568,N_13234,N_13231);
nand U13569 (N_13569,N_13232,N_13296);
and U13570 (N_13570,N_13386,N_13352);
nor U13571 (N_13571,N_13358,N_13351);
or U13572 (N_13572,N_13301,N_13217);
nor U13573 (N_13573,N_13296,N_13337);
xor U13574 (N_13574,N_13202,N_13389);
or U13575 (N_13575,N_13383,N_13377);
nor U13576 (N_13576,N_13205,N_13304);
and U13577 (N_13577,N_13371,N_13203);
or U13578 (N_13578,N_13308,N_13217);
or U13579 (N_13579,N_13201,N_13330);
or U13580 (N_13580,N_13248,N_13283);
and U13581 (N_13581,N_13292,N_13383);
nand U13582 (N_13582,N_13284,N_13390);
nand U13583 (N_13583,N_13316,N_13224);
or U13584 (N_13584,N_13235,N_13332);
and U13585 (N_13585,N_13269,N_13209);
nor U13586 (N_13586,N_13336,N_13376);
xnor U13587 (N_13587,N_13385,N_13266);
xnor U13588 (N_13588,N_13243,N_13285);
nor U13589 (N_13589,N_13241,N_13313);
or U13590 (N_13590,N_13340,N_13337);
xnor U13591 (N_13591,N_13271,N_13250);
nand U13592 (N_13592,N_13333,N_13326);
or U13593 (N_13593,N_13259,N_13223);
nor U13594 (N_13594,N_13204,N_13340);
and U13595 (N_13595,N_13394,N_13217);
nand U13596 (N_13596,N_13250,N_13384);
nand U13597 (N_13597,N_13342,N_13228);
and U13598 (N_13598,N_13316,N_13208);
xor U13599 (N_13599,N_13361,N_13212);
nor U13600 (N_13600,N_13587,N_13410);
and U13601 (N_13601,N_13519,N_13491);
or U13602 (N_13602,N_13549,N_13465);
nand U13603 (N_13603,N_13454,N_13516);
or U13604 (N_13604,N_13506,N_13414);
nand U13605 (N_13605,N_13492,N_13495);
nor U13606 (N_13606,N_13566,N_13541);
nand U13607 (N_13607,N_13422,N_13479);
nand U13608 (N_13608,N_13542,N_13552);
nand U13609 (N_13609,N_13559,N_13538);
nand U13610 (N_13610,N_13494,N_13515);
xor U13611 (N_13611,N_13427,N_13534);
xor U13612 (N_13612,N_13527,N_13579);
xor U13613 (N_13613,N_13416,N_13503);
xor U13614 (N_13614,N_13407,N_13502);
nor U13615 (N_13615,N_13562,N_13509);
xnor U13616 (N_13616,N_13412,N_13486);
nand U13617 (N_13617,N_13499,N_13592);
or U13618 (N_13618,N_13467,N_13547);
xnor U13619 (N_13619,N_13569,N_13565);
nand U13620 (N_13620,N_13507,N_13472);
or U13621 (N_13621,N_13482,N_13554);
or U13622 (N_13622,N_13432,N_13484);
xor U13623 (N_13623,N_13449,N_13403);
xnor U13624 (N_13624,N_13537,N_13535);
nor U13625 (N_13625,N_13557,N_13582);
and U13626 (N_13626,N_13460,N_13525);
xor U13627 (N_13627,N_13511,N_13452);
and U13628 (N_13628,N_13590,N_13585);
nor U13629 (N_13629,N_13483,N_13532);
nand U13630 (N_13630,N_13470,N_13555);
xor U13631 (N_13631,N_13424,N_13481);
xnor U13632 (N_13632,N_13560,N_13567);
or U13633 (N_13633,N_13433,N_13469);
nor U13634 (N_13634,N_13531,N_13437);
or U13635 (N_13635,N_13501,N_13448);
nor U13636 (N_13636,N_13426,N_13533);
xor U13637 (N_13637,N_13419,N_13443);
and U13638 (N_13638,N_13488,N_13423);
nand U13639 (N_13639,N_13468,N_13480);
or U13640 (N_13640,N_13584,N_13505);
nand U13641 (N_13641,N_13508,N_13447);
nand U13642 (N_13642,N_13456,N_13586);
and U13643 (N_13643,N_13487,N_13445);
xor U13644 (N_13644,N_13477,N_13524);
xor U13645 (N_13645,N_13597,N_13438);
xor U13646 (N_13646,N_13421,N_13400);
and U13647 (N_13647,N_13520,N_13466);
xor U13648 (N_13648,N_13420,N_13459);
and U13649 (N_13649,N_13510,N_13498);
xor U13650 (N_13650,N_13588,N_13404);
and U13651 (N_13651,N_13446,N_13530);
nor U13652 (N_13652,N_13455,N_13595);
and U13653 (N_13653,N_13573,N_13551);
and U13654 (N_13654,N_13553,N_13496);
nor U13655 (N_13655,N_13593,N_13409);
or U13656 (N_13656,N_13471,N_13493);
and U13657 (N_13657,N_13429,N_13478);
or U13658 (N_13658,N_13563,N_13457);
xnor U13659 (N_13659,N_13439,N_13546);
and U13660 (N_13660,N_13473,N_13529);
and U13661 (N_13661,N_13474,N_13425);
nor U13662 (N_13662,N_13489,N_13434);
nand U13663 (N_13663,N_13451,N_13512);
or U13664 (N_13664,N_13568,N_13581);
nor U13665 (N_13665,N_13517,N_13476);
xor U13666 (N_13666,N_13522,N_13575);
or U13667 (N_13667,N_13526,N_13596);
nor U13668 (N_13668,N_13572,N_13539);
nor U13669 (N_13669,N_13543,N_13415);
xor U13670 (N_13670,N_13558,N_13536);
or U13671 (N_13671,N_13594,N_13570);
xnor U13672 (N_13672,N_13436,N_13523);
nand U13673 (N_13673,N_13580,N_13556);
and U13674 (N_13674,N_13442,N_13408);
nor U13675 (N_13675,N_13458,N_13513);
nor U13676 (N_13676,N_13561,N_13453);
or U13677 (N_13677,N_13548,N_13577);
nand U13678 (N_13678,N_13406,N_13576);
xor U13679 (N_13679,N_13440,N_13540);
and U13680 (N_13680,N_13462,N_13402);
or U13681 (N_13681,N_13591,N_13528);
and U13682 (N_13682,N_13544,N_13504);
or U13683 (N_13683,N_13461,N_13405);
or U13684 (N_13684,N_13464,N_13430);
or U13685 (N_13685,N_13411,N_13441);
and U13686 (N_13686,N_13583,N_13521);
nor U13687 (N_13687,N_13571,N_13578);
or U13688 (N_13688,N_13589,N_13545);
nand U13689 (N_13689,N_13431,N_13413);
or U13690 (N_13690,N_13564,N_13417);
or U13691 (N_13691,N_13490,N_13497);
nor U13692 (N_13692,N_13428,N_13500);
or U13693 (N_13693,N_13574,N_13401);
nand U13694 (N_13694,N_13599,N_13450);
nand U13695 (N_13695,N_13475,N_13444);
nor U13696 (N_13696,N_13418,N_13485);
or U13697 (N_13697,N_13598,N_13518);
nand U13698 (N_13698,N_13514,N_13463);
xnor U13699 (N_13699,N_13550,N_13435);
nand U13700 (N_13700,N_13450,N_13571);
xnor U13701 (N_13701,N_13526,N_13571);
and U13702 (N_13702,N_13403,N_13522);
nor U13703 (N_13703,N_13445,N_13447);
and U13704 (N_13704,N_13584,N_13428);
or U13705 (N_13705,N_13465,N_13599);
and U13706 (N_13706,N_13458,N_13453);
xnor U13707 (N_13707,N_13580,N_13520);
nor U13708 (N_13708,N_13465,N_13438);
nor U13709 (N_13709,N_13457,N_13444);
and U13710 (N_13710,N_13496,N_13493);
nand U13711 (N_13711,N_13427,N_13541);
nor U13712 (N_13712,N_13436,N_13426);
and U13713 (N_13713,N_13495,N_13493);
nor U13714 (N_13714,N_13580,N_13554);
xnor U13715 (N_13715,N_13527,N_13430);
nor U13716 (N_13716,N_13587,N_13580);
nand U13717 (N_13717,N_13509,N_13405);
nand U13718 (N_13718,N_13488,N_13466);
nand U13719 (N_13719,N_13462,N_13497);
nor U13720 (N_13720,N_13568,N_13536);
or U13721 (N_13721,N_13480,N_13530);
xor U13722 (N_13722,N_13548,N_13469);
nand U13723 (N_13723,N_13403,N_13509);
nand U13724 (N_13724,N_13451,N_13588);
xnor U13725 (N_13725,N_13458,N_13421);
nand U13726 (N_13726,N_13535,N_13500);
nand U13727 (N_13727,N_13551,N_13400);
nor U13728 (N_13728,N_13485,N_13516);
nor U13729 (N_13729,N_13557,N_13410);
nand U13730 (N_13730,N_13486,N_13529);
nand U13731 (N_13731,N_13560,N_13535);
xor U13732 (N_13732,N_13593,N_13532);
xnor U13733 (N_13733,N_13557,N_13482);
and U13734 (N_13734,N_13425,N_13487);
and U13735 (N_13735,N_13505,N_13588);
or U13736 (N_13736,N_13522,N_13401);
xor U13737 (N_13737,N_13428,N_13410);
nand U13738 (N_13738,N_13413,N_13489);
xor U13739 (N_13739,N_13451,N_13561);
nand U13740 (N_13740,N_13556,N_13429);
or U13741 (N_13741,N_13498,N_13548);
xor U13742 (N_13742,N_13427,N_13432);
and U13743 (N_13743,N_13486,N_13508);
or U13744 (N_13744,N_13553,N_13576);
or U13745 (N_13745,N_13451,N_13418);
nand U13746 (N_13746,N_13463,N_13536);
nor U13747 (N_13747,N_13444,N_13509);
xor U13748 (N_13748,N_13437,N_13575);
nand U13749 (N_13749,N_13548,N_13456);
and U13750 (N_13750,N_13458,N_13415);
or U13751 (N_13751,N_13467,N_13418);
nor U13752 (N_13752,N_13442,N_13527);
nor U13753 (N_13753,N_13538,N_13432);
nor U13754 (N_13754,N_13466,N_13536);
xnor U13755 (N_13755,N_13550,N_13404);
nor U13756 (N_13756,N_13523,N_13448);
nor U13757 (N_13757,N_13526,N_13510);
nand U13758 (N_13758,N_13552,N_13490);
nor U13759 (N_13759,N_13569,N_13571);
or U13760 (N_13760,N_13596,N_13516);
nand U13761 (N_13761,N_13537,N_13422);
nand U13762 (N_13762,N_13477,N_13567);
and U13763 (N_13763,N_13445,N_13584);
nor U13764 (N_13764,N_13458,N_13538);
or U13765 (N_13765,N_13467,N_13552);
nor U13766 (N_13766,N_13533,N_13485);
or U13767 (N_13767,N_13568,N_13408);
and U13768 (N_13768,N_13440,N_13462);
or U13769 (N_13769,N_13535,N_13502);
nand U13770 (N_13770,N_13519,N_13477);
or U13771 (N_13771,N_13426,N_13493);
xor U13772 (N_13772,N_13459,N_13471);
and U13773 (N_13773,N_13541,N_13537);
and U13774 (N_13774,N_13415,N_13526);
xor U13775 (N_13775,N_13496,N_13579);
nor U13776 (N_13776,N_13413,N_13545);
or U13777 (N_13777,N_13409,N_13587);
nand U13778 (N_13778,N_13556,N_13481);
nor U13779 (N_13779,N_13476,N_13448);
xnor U13780 (N_13780,N_13598,N_13495);
and U13781 (N_13781,N_13541,N_13410);
xnor U13782 (N_13782,N_13518,N_13559);
or U13783 (N_13783,N_13573,N_13505);
xnor U13784 (N_13784,N_13475,N_13524);
nand U13785 (N_13785,N_13421,N_13498);
or U13786 (N_13786,N_13426,N_13523);
nand U13787 (N_13787,N_13489,N_13427);
nor U13788 (N_13788,N_13539,N_13559);
and U13789 (N_13789,N_13512,N_13423);
or U13790 (N_13790,N_13514,N_13586);
or U13791 (N_13791,N_13554,N_13478);
and U13792 (N_13792,N_13497,N_13509);
xnor U13793 (N_13793,N_13512,N_13461);
xor U13794 (N_13794,N_13520,N_13488);
xnor U13795 (N_13795,N_13544,N_13581);
xnor U13796 (N_13796,N_13567,N_13408);
nand U13797 (N_13797,N_13592,N_13550);
and U13798 (N_13798,N_13513,N_13572);
xnor U13799 (N_13799,N_13531,N_13414);
nor U13800 (N_13800,N_13747,N_13601);
nand U13801 (N_13801,N_13730,N_13626);
xor U13802 (N_13802,N_13680,N_13761);
and U13803 (N_13803,N_13683,N_13740);
and U13804 (N_13804,N_13785,N_13640);
and U13805 (N_13805,N_13631,N_13779);
nand U13806 (N_13806,N_13604,N_13764);
nand U13807 (N_13807,N_13789,N_13718);
and U13808 (N_13808,N_13731,N_13629);
nor U13809 (N_13809,N_13630,N_13754);
and U13810 (N_13810,N_13797,N_13732);
xor U13811 (N_13811,N_13669,N_13671);
nand U13812 (N_13812,N_13697,N_13651);
nor U13813 (N_13813,N_13649,N_13733);
nor U13814 (N_13814,N_13663,N_13796);
xor U13815 (N_13815,N_13682,N_13793);
or U13816 (N_13816,N_13638,N_13742);
nor U13817 (N_13817,N_13798,N_13790);
and U13818 (N_13818,N_13757,N_13695);
and U13819 (N_13819,N_13759,N_13643);
and U13820 (N_13820,N_13679,N_13622);
nand U13821 (N_13821,N_13737,N_13636);
nor U13822 (N_13822,N_13709,N_13784);
and U13823 (N_13823,N_13620,N_13749);
or U13824 (N_13824,N_13750,N_13788);
nand U13825 (N_13825,N_13723,N_13687);
xor U13826 (N_13826,N_13613,N_13600);
nor U13827 (N_13827,N_13662,N_13748);
xor U13828 (N_13828,N_13675,N_13642);
or U13829 (N_13829,N_13603,N_13625);
xor U13830 (N_13830,N_13717,N_13650);
and U13831 (N_13831,N_13678,N_13736);
nand U13832 (N_13832,N_13724,N_13701);
xnor U13833 (N_13833,N_13794,N_13741);
nor U13834 (N_13834,N_13602,N_13783);
and U13835 (N_13835,N_13692,N_13777);
xor U13836 (N_13836,N_13743,N_13693);
xnor U13837 (N_13837,N_13677,N_13707);
xor U13838 (N_13838,N_13756,N_13714);
xor U13839 (N_13839,N_13791,N_13763);
xnor U13840 (N_13840,N_13619,N_13735);
xnor U13841 (N_13841,N_13658,N_13728);
or U13842 (N_13842,N_13653,N_13664);
and U13843 (N_13843,N_13726,N_13702);
nand U13844 (N_13844,N_13667,N_13713);
nand U13845 (N_13845,N_13769,N_13795);
nor U13846 (N_13846,N_13772,N_13617);
nand U13847 (N_13847,N_13673,N_13684);
nand U13848 (N_13848,N_13610,N_13786);
and U13849 (N_13849,N_13751,N_13778);
nand U13850 (N_13850,N_13771,N_13628);
and U13851 (N_13851,N_13689,N_13746);
and U13852 (N_13852,N_13627,N_13612);
or U13853 (N_13853,N_13725,N_13787);
nor U13854 (N_13854,N_13632,N_13699);
or U13855 (N_13855,N_13755,N_13607);
xor U13856 (N_13856,N_13688,N_13660);
xnor U13857 (N_13857,N_13666,N_13654);
nor U13858 (N_13858,N_13608,N_13776);
and U13859 (N_13859,N_13729,N_13656);
and U13860 (N_13860,N_13722,N_13690);
nand U13861 (N_13861,N_13681,N_13655);
or U13862 (N_13862,N_13739,N_13611);
or U13863 (N_13863,N_13659,N_13606);
or U13864 (N_13864,N_13645,N_13674);
nand U13865 (N_13865,N_13652,N_13657);
nor U13866 (N_13866,N_13760,N_13727);
and U13867 (N_13867,N_13721,N_13708);
or U13868 (N_13868,N_13686,N_13644);
xor U13869 (N_13869,N_13694,N_13792);
nand U13870 (N_13870,N_13661,N_13646);
or U13871 (N_13871,N_13648,N_13704);
nand U13872 (N_13872,N_13665,N_13711);
xnor U13873 (N_13873,N_13780,N_13799);
and U13874 (N_13874,N_13781,N_13621);
and U13875 (N_13875,N_13765,N_13676);
and U13876 (N_13876,N_13647,N_13720);
nand U13877 (N_13877,N_13634,N_13753);
nor U13878 (N_13878,N_13696,N_13782);
nor U13879 (N_13879,N_13623,N_13672);
xor U13880 (N_13880,N_13758,N_13624);
nand U13881 (N_13881,N_13716,N_13715);
nand U13882 (N_13882,N_13706,N_13734);
nor U13883 (N_13883,N_13609,N_13770);
nor U13884 (N_13884,N_13712,N_13641);
and U13885 (N_13885,N_13698,N_13705);
nand U13886 (N_13886,N_13639,N_13637);
nand U13887 (N_13887,N_13635,N_13775);
and U13888 (N_13888,N_13616,N_13691);
nor U13889 (N_13889,N_13767,N_13766);
and U13890 (N_13890,N_13668,N_13719);
nor U13891 (N_13891,N_13685,N_13744);
nand U13892 (N_13892,N_13605,N_13738);
nand U13893 (N_13893,N_13703,N_13618);
or U13894 (N_13894,N_13773,N_13762);
nor U13895 (N_13895,N_13710,N_13633);
or U13896 (N_13896,N_13774,N_13615);
nor U13897 (N_13897,N_13752,N_13614);
nor U13898 (N_13898,N_13670,N_13768);
nor U13899 (N_13899,N_13745,N_13700);
or U13900 (N_13900,N_13789,N_13683);
nor U13901 (N_13901,N_13627,N_13654);
nand U13902 (N_13902,N_13773,N_13714);
or U13903 (N_13903,N_13752,N_13749);
or U13904 (N_13904,N_13704,N_13719);
and U13905 (N_13905,N_13641,N_13640);
and U13906 (N_13906,N_13669,N_13678);
nand U13907 (N_13907,N_13761,N_13688);
and U13908 (N_13908,N_13643,N_13606);
nor U13909 (N_13909,N_13680,N_13717);
nor U13910 (N_13910,N_13765,N_13622);
nand U13911 (N_13911,N_13791,N_13675);
or U13912 (N_13912,N_13655,N_13614);
xor U13913 (N_13913,N_13707,N_13744);
or U13914 (N_13914,N_13675,N_13666);
or U13915 (N_13915,N_13682,N_13687);
xor U13916 (N_13916,N_13765,N_13789);
nand U13917 (N_13917,N_13730,N_13685);
nor U13918 (N_13918,N_13693,N_13725);
xnor U13919 (N_13919,N_13635,N_13797);
nand U13920 (N_13920,N_13738,N_13796);
and U13921 (N_13921,N_13763,N_13732);
or U13922 (N_13922,N_13790,N_13687);
and U13923 (N_13923,N_13644,N_13697);
nand U13924 (N_13924,N_13644,N_13693);
nor U13925 (N_13925,N_13636,N_13718);
nor U13926 (N_13926,N_13660,N_13721);
or U13927 (N_13927,N_13691,N_13633);
xnor U13928 (N_13928,N_13686,N_13798);
or U13929 (N_13929,N_13740,N_13711);
nand U13930 (N_13930,N_13676,N_13678);
xor U13931 (N_13931,N_13752,N_13698);
and U13932 (N_13932,N_13615,N_13694);
nor U13933 (N_13933,N_13686,N_13717);
or U13934 (N_13934,N_13721,N_13780);
and U13935 (N_13935,N_13646,N_13743);
or U13936 (N_13936,N_13620,N_13669);
nor U13937 (N_13937,N_13758,N_13715);
or U13938 (N_13938,N_13794,N_13685);
nand U13939 (N_13939,N_13601,N_13653);
or U13940 (N_13940,N_13768,N_13785);
nand U13941 (N_13941,N_13617,N_13640);
nor U13942 (N_13942,N_13742,N_13657);
nor U13943 (N_13943,N_13714,N_13640);
or U13944 (N_13944,N_13765,N_13701);
nand U13945 (N_13945,N_13609,N_13792);
nand U13946 (N_13946,N_13788,N_13772);
and U13947 (N_13947,N_13772,N_13699);
or U13948 (N_13948,N_13607,N_13601);
nand U13949 (N_13949,N_13705,N_13779);
and U13950 (N_13950,N_13706,N_13697);
or U13951 (N_13951,N_13742,N_13752);
nand U13952 (N_13952,N_13797,N_13686);
nand U13953 (N_13953,N_13677,N_13761);
xor U13954 (N_13954,N_13644,N_13735);
and U13955 (N_13955,N_13784,N_13658);
nor U13956 (N_13956,N_13744,N_13668);
nor U13957 (N_13957,N_13640,N_13724);
or U13958 (N_13958,N_13654,N_13782);
or U13959 (N_13959,N_13608,N_13758);
xnor U13960 (N_13960,N_13651,N_13664);
nor U13961 (N_13961,N_13656,N_13606);
xor U13962 (N_13962,N_13733,N_13743);
and U13963 (N_13963,N_13743,N_13661);
nor U13964 (N_13964,N_13781,N_13618);
and U13965 (N_13965,N_13791,N_13654);
nor U13966 (N_13966,N_13617,N_13739);
or U13967 (N_13967,N_13623,N_13636);
or U13968 (N_13968,N_13711,N_13758);
xor U13969 (N_13969,N_13701,N_13602);
and U13970 (N_13970,N_13781,N_13685);
and U13971 (N_13971,N_13748,N_13760);
and U13972 (N_13972,N_13739,N_13707);
nand U13973 (N_13973,N_13622,N_13680);
or U13974 (N_13974,N_13649,N_13688);
nand U13975 (N_13975,N_13627,N_13740);
or U13976 (N_13976,N_13722,N_13620);
xor U13977 (N_13977,N_13638,N_13678);
and U13978 (N_13978,N_13713,N_13629);
nand U13979 (N_13979,N_13668,N_13625);
nand U13980 (N_13980,N_13637,N_13675);
xnor U13981 (N_13981,N_13675,N_13796);
or U13982 (N_13982,N_13716,N_13776);
or U13983 (N_13983,N_13779,N_13716);
nand U13984 (N_13984,N_13626,N_13630);
xnor U13985 (N_13985,N_13738,N_13677);
xor U13986 (N_13986,N_13692,N_13639);
xor U13987 (N_13987,N_13708,N_13725);
or U13988 (N_13988,N_13649,N_13703);
and U13989 (N_13989,N_13658,N_13788);
xnor U13990 (N_13990,N_13713,N_13733);
xor U13991 (N_13991,N_13619,N_13671);
and U13992 (N_13992,N_13618,N_13799);
or U13993 (N_13993,N_13616,N_13631);
xor U13994 (N_13994,N_13798,N_13720);
nor U13995 (N_13995,N_13655,N_13652);
nand U13996 (N_13996,N_13732,N_13766);
nand U13997 (N_13997,N_13604,N_13610);
nand U13998 (N_13998,N_13658,N_13743);
nand U13999 (N_13999,N_13697,N_13731);
or U14000 (N_14000,N_13994,N_13928);
nor U14001 (N_14001,N_13986,N_13855);
or U14002 (N_14002,N_13875,N_13912);
or U14003 (N_14003,N_13806,N_13882);
nand U14004 (N_14004,N_13831,N_13987);
or U14005 (N_14005,N_13958,N_13979);
nand U14006 (N_14006,N_13990,N_13863);
nand U14007 (N_14007,N_13949,N_13918);
nand U14008 (N_14008,N_13982,N_13872);
nand U14009 (N_14009,N_13942,N_13884);
xor U14010 (N_14010,N_13812,N_13866);
and U14011 (N_14011,N_13953,N_13825);
xnor U14012 (N_14012,N_13888,N_13814);
or U14013 (N_14013,N_13818,N_13943);
or U14014 (N_14014,N_13807,N_13985);
and U14015 (N_14015,N_13952,N_13995);
nor U14016 (N_14016,N_13864,N_13964);
nor U14017 (N_14017,N_13852,N_13996);
nand U14018 (N_14018,N_13902,N_13908);
and U14019 (N_14019,N_13824,N_13898);
xnor U14020 (N_14020,N_13926,N_13878);
or U14021 (N_14021,N_13983,N_13838);
xnor U14022 (N_14022,N_13896,N_13873);
nand U14023 (N_14023,N_13847,N_13925);
or U14024 (N_14024,N_13885,N_13800);
nand U14025 (N_14025,N_13922,N_13936);
nand U14026 (N_14026,N_13955,N_13886);
nor U14027 (N_14027,N_13808,N_13978);
xnor U14028 (N_14028,N_13843,N_13981);
and U14029 (N_14029,N_13932,N_13883);
nor U14030 (N_14030,N_13803,N_13837);
or U14031 (N_14031,N_13931,N_13862);
nor U14032 (N_14032,N_13934,N_13881);
or U14033 (N_14033,N_13917,N_13962);
or U14034 (N_14034,N_13961,N_13867);
xnor U14035 (N_14035,N_13820,N_13841);
or U14036 (N_14036,N_13856,N_13822);
nand U14037 (N_14037,N_13945,N_13868);
nor U14038 (N_14038,N_13998,N_13933);
xor U14039 (N_14039,N_13944,N_13966);
or U14040 (N_14040,N_13924,N_13997);
and U14041 (N_14041,N_13907,N_13861);
xor U14042 (N_14042,N_13810,N_13965);
or U14043 (N_14043,N_13938,N_13920);
or U14044 (N_14044,N_13858,N_13816);
xnor U14045 (N_14045,N_13891,N_13980);
or U14046 (N_14046,N_13963,N_13969);
or U14047 (N_14047,N_13999,N_13840);
xnor U14048 (N_14048,N_13839,N_13951);
or U14049 (N_14049,N_13857,N_13874);
and U14050 (N_14050,N_13832,N_13870);
nand U14051 (N_14051,N_13984,N_13830);
xnor U14052 (N_14052,N_13801,N_13959);
nor U14053 (N_14053,N_13915,N_13971);
nor U14054 (N_14054,N_13890,N_13941);
or U14055 (N_14055,N_13992,N_13901);
xnor U14056 (N_14056,N_13865,N_13836);
and U14057 (N_14057,N_13827,N_13853);
or U14058 (N_14058,N_13876,N_13970);
nor U14059 (N_14059,N_13906,N_13960);
xnor U14060 (N_14060,N_13976,N_13948);
nor U14061 (N_14061,N_13802,N_13826);
nand U14062 (N_14062,N_13887,N_13821);
and U14063 (N_14063,N_13929,N_13919);
nor U14064 (N_14064,N_13916,N_13911);
and U14065 (N_14065,N_13974,N_13921);
nand U14066 (N_14066,N_13954,N_13939);
or U14067 (N_14067,N_13849,N_13975);
and U14068 (N_14068,N_13900,N_13813);
nor U14069 (N_14069,N_13889,N_13817);
and U14070 (N_14070,N_13879,N_13850);
nor U14071 (N_14071,N_13835,N_13991);
nand U14072 (N_14072,N_13950,N_13809);
nand U14073 (N_14073,N_13804,N_13935);
and U14074 (N_14074,N_13904,N_13897);
nand U14075 (N_14075,N_13895,N_13909);
nand U14076 (N_14076,N_13927,N_13811);
and U14077 (N_14077,N_13823,N_13844);
nand U14078 (N_14078,N_13869,N_13968);
xnor U14079 (N_14079,N_13957,N_13805);
nand U14080 (N_14080,N_13977,N_13940);
nor U14081 (N_14081,N_13946,N_13892);
and U14082 (N_14082,N_13989,N_13967);
nor U14083 (N_14083,N_13988,N_13846);
nand U14084 (N_14084,N_13842,N_13956);
xnor U14085 (N_14085,N_13845,N_13923);
and U14086 (N_14086,N_13914,N_13851);
nor U14087 (N_14087,N_13848,N_13937);
and U14088 (N_14088,N_13910,N_13877);
nor U14089 (N_14089,N_13834,N_13871);
or U14090 (N_14090,N_13815,N_13854);
xnor U14091 (N_14091,N_13819,N_13930);
nand U14092 (N_14092,N_13899,N_13860);
nand U14093 (N_14093,N_13859,N_13829);
and U14094 (N_14094,N_13913,N_13894);
nor U14095 (N_14095,N_13903,N_13972);
nand U14096 (N_14096,N_13893,N_13947);
or U14097 (N_14097,N_13973,N_13833);
or U14098 (N_14098,N_13880,N_13905);
nor U14099 (N_14099,N_13828,N_13993);
and U14100 (N_14100,N_13904,N_13802);
nor U14101 (N_14101,N_13866,N_13805);
or U14102 (N_14102,N_13975,N_13912);
nor U14103 (N_14103,N_13929,N_13909);
and U14104 (N_14104,N_13950,N_13921);
and U14105 (N_14105,N_13921,N_13801);
nand U14106 (N_14106,N_13852,N_13865);
nor U14107 (N_14107,N_13905,N_13902);
nand U14108 (N_14108,N_13932,N_13878);
nor U14109 (N_14109,N_13946,N_13949);
xnor U14110 (N_14110,N_13833,N_13870);
and U14111 (N_14111,N_13905,N_13973);
nor U14112 (N_14112,N_13923,N_13980);
xor U14113 (N_14113,N_13994,N_13867);
or U14114 (N_14114,N_13930,N_13990);
and U14115 (N_14115,N_13917,N_13832);
and U14116 (N_14116,N_13984,N_13833);
or U14117 (N_14117,N_13999,N_13886);
or U14118 (N_14118,N_13843,N_13974);
nand U14119 (N_14119,N_13985,N_13894);
and U14120 (N_14120,N_13889,N_13914);
xor U14121 (N_14121,N_13825,N_13879);
nor U14122 (N_14122,N_13923,N_13912);
and U14123 (N_14123,N_13893,N_13920);
or U14124 (N_14124,N_13960,N_13929);
nand U14125 (N_14125,N_13811,N_13967);
and U14126 (N_14126,N_13925,N_13986);
nand U14127 (N_14127,N_13918,N_13828);
xor U14128 (N_14128,N_13805,N_13951);
xor U14129 (N_14129,N_13818,N_13979);
xor U14130 (N_14130,N_13897,N_13905);
nor U14131 (N_14131,N_13916,N_13984);
xnor U14132 (N_14132,N_13836,N_13902);
nand U14133 (N_14133,N_13954,N_13826);
nor U14134 (N_14134,N_13884,N_13965);
and U14135 (N_14135,N_13975,N_13995);
or U14136 (N_14136,N_13993,N_13818);
or U14137 (N_14137,N_13972,N_13957);
or U14138 (N_14138,N_13884,N_13845);
and U14139 (N_14139,N_13919,N_13890);
and U14140 (N_14140,N_13802,N_13900);
nor U14141 (N_14141,N_13981,N_13882);
and U14142 (N_14142,N_13979,N_13977);
or U14143 (N_14143,N_13996,N_13994);
and U14144 (N_14144,N_13846,N_13819);
nand U14145 (N_14145,N_13976,N_13803);
and U14146 (N_14146,N_13993,N_13881);
nand U14147 (N_14147,N_13881,N_13991);
nand U14148 (N_14148,N_13801,N_13976);
nor U14149 (N_14149,N_13893,N_13849);
nor U14150 (N_14150,N_13850,N_13901);
or U14151 (N_14151,N_13848,N_13980);
nor U14152 (N_14152,N_13870,N_13885);
nor U14153 (N_14153,N_13844,N_13954);
nor U14154 (N_14154,N_13943,N_13975);
xor U14155 (N_14155,N_13804,N_13852);
xnor U14156 (N_14156,N_13925,N_13905);
nor U14157 (N_14157,N_13940,N_13934);
nor U14158 (N_14158,N_13942,N_13984);
xor U14159 (N_14159,N_13879,N_13811);
xnor U14160 (N_14160,N_13858,N_13936);
nor U14161 (N_14161,N_13863,N_13813);
nand U14162 (N_14162,N_13866,N_13932);
and U14163 (N_14163,N_13808,N_13818);
xnor U14164 (N_14164,N_13960,N_13859);
and U14165 (N_14165,N_13921,N_13843);
and U14166 (N_14166,N_13943,N_13862);
and U14167 (N_14167,N_13985,N_13901);
xor U14168 (N_14168,N_13936,N_13918);
or U14169 (N_14169,N_13948,N_13946);
nor U14170 (N_14170,N_13867,N_13822);
nor U14171 (N_14171,N_13991,N_13934);
or U14172 (N_14172,N_13960,N_13908);
or U14173 (N_14173,N_13960,N_13869);
or U14174 (N_14174,N_13821,N_13956);
and U14175 (N_14175,N_13915,N_13870);
xor U14176 (N_14176,N_13824,N_13950);
and U14177 (N_14177,N_13861,N_13902);
xor U14178 (N_14178,N_13953,N_13972);
xor U14179 (N_14179,N_13952,N_13842);
and U14180 (N_14180,N_13917,N_13968);
nor U14181 (N_14181,N_13863,N_13903);
nor U14182 (N_14182,N_13932,N_13944);
nand U14183 (N_14183,N_13858,N_13962);
and U14184 (N_14184,N_13867,N_13816);
or U14185 (N_14185,N_13873,N_13990);
or U14186 (N_14186,N_13909,N_13857);
nand U14187 (N_14187,N_13902,N_13800);
or U14188 (N_14188,N_13942,N_13875);
nor U14189 (N_14189,N_13961,N_13862);
or U14190 (N_14190,N_13924,N_13892);
nor U14191 (N_14191,N_13834,N_13931);
or U14192 (N_14192,N_13953,N_13995);
nor U14193 (N_14193,N_13858,N_13981);
nor U14194 (N_14194,N_13827,N_13878);
or U14195 (N_14195,N_13968,N_13882);
and U14196 (N_14196,N_13818,N_13978);
and U14197 (N_14197,N_13894,N_13982);
nand U14198 (N_14198,N_13904,N_13995);
xor U14199 (N_14199,N_13922,N_13876);
nand U14200 (N_14200,N_14046,N_14132);
or U14201 (N_14201,N_14045,N_14092);
and U14202 (N_14202,N_14177,N_14015);
xnor U14203 (N_14203,N_14061,N_14077);
nor U14204 (N_14204,N_14039,N_14073);
and U14205 (N_14205,N_14145,N_14110);
nand U14206 (N_14206,N_14172,N_14125);
nor U14207 (N_14207,N_14066,N_14161);
xor U14208 (N_14208,N_14118,N_14042);
xor U14209 (N_14209,N_14026,N_14184);
or U14210 (N_14210,N_14129,N_14011);
nor U14211 (N_14211,N_14059,N_14179);
or U14212 (N_14212,N_14079,N_14148);
nor U14213 (N_14213,N_14126,N_14101);
xnor U14214 (N_14214,N_14174,N_14183);
and U14215 (N_14215,N_14016,N_14117);
and U14216 (N_14216,N_14030,N_14072);
nor U14217 (N_14217,N_14084,N_14180);
nor U14218 (N_14218,N_14080,N_14107);
xnor U14219 (N_14219,N_14078,N_14008);
xor U14220 (N_14220,N_14071,N_14181);
nand U14221 (N_14221,N_14195,N_14143);
or U14222 (N_14222,N_14095,N_14043);
nor U14223 (N_14223,N_14113,N_14038);
nor U14224 (N_14224,N_14168,N_14051);
and U14225 (N_14225,N_14152,N_14105);
xor U14226 (N_14226,N_14048,N_14050);
and U14227 (N_14227,N_14150,N_14186);
or U14228 (N_14228,N_14182,N_14196);
xor U14229 (N_14229,N_14022,N_14058);
or U14230 (N_14230,N_14147,N_14023);
nor U14231 (N_14231,N_14106,N_14185);
nand U14232 (N_14232,N_14169,N_14197);
nand U14233 (N_14233,N_14010,N_14131);
or U14234 (N_14234,N_14173,N_14193);
or U14235 (N_14235,N_14018,N_14053);
nand U14236 (N_14236,N_14031,N_14122);
xnor U14237 (N_14237,N_14153,N_14109);
or U14238 (N_14238,N_14124,N_14114);
xnor U14239 (N_14239,N_14149,N_14088);
nor U14240 (N_14240,N_14004,N_14190);
or U14241 (N_14241,N_14093,N_14067);
nor U14242 (N_14242,N_14094,N_14069);
xnor U14243 (N_14243,N_14020,N_14134);
and U14244 (N_14244,N_14044,N_14056);
nor U14245 (N_14245,N_14108,N_14194);
or U14246 (N_14246,N_14017,N_14191);
nand U14247 (N_14247,N_14086,N_14036);
or U14248 (N_14248,N_14176,N_14060);
and U14249 (N_14249,N_14006,N_14189);
or U14250 (N_14250,N_14139,N_14116);
nor U14251 (N_14251,N_14001,N_14064);
nand U14252 (N_14252,N_14014,N_14141);
and U14253 (N_14253,N_14121,N_14054);
xnor U14254 (N_14254,N_14009,N_14024);
and U14255 (N_14255,N_14175,N_14033);
nor U14256 (N_14256,N_14019,N_14133);
nand U14257 (N_14257,N_14076,N_14000);
and U14258 (N_14258,N_14055,N_14170);
or U14259 (N_14259,N_14021,N_14063);
nor U14260 (N_14260,N_14085,N_14104);
and U14261 (N_14261,N_14035,N_14074);
nand U14262 (N_14262,N_14041,N_14070);
nand U14263 (N_14263,N_14178,N_14112);
and U14264 (N_14264,N_14089,N_14111);
and U14265 (N_14265,N_14167,N_14140);
xnor U14266 (N_14266,N_14130,N_14096);
nand U14267 (N_14267,N_14159,N_14075);
nand U14268 (N_14268,N_14119,N_14187);
nand U14269 (N_14269,N_14083,N_14013);
nand U14270 (N_14270,N_14100,N_14137);
or U14271 (N_14271,N_14047,N_14003);
nor U14272 (N_14272,N_14155,N_14103);
nand U14273 (N_14273,N_14025,N_14120);
xnor U14274 (N_14274,N_14007,N_14040);
xor U14275 (N_14275,N_14034,N_14082);
xor U14276 (N_14276,N_14171,N_14068);
nor U14277 (N_14277,N_14049,N_14123);
xor U14278 (N_14278,N_14087,N_14163);
nand U14279 (N_14279,N_14142,N_14127);
or U14280 (N_14280,N_14029,N_14005);
xnor U14281 (N_14281,N_14097,N_14027);
nor U14282 (N_14282,N_14012,N_14156);
nor U14283 (N_14283,N_14052,N_14188);
nor U14284 (N_14284,N_14165,N_14164);
xor U14285 (N_14285,N_14198,N_14065);
xnor U14286 (N_14286,N_14157,N_14002);
xor U14287 (N_14287,N_14160,N_14154);
xnor U14288 (N_14288,N_14199,N_14057);
and U14289 (N_14289,N_14028,N_14098);
nor U14290 (N_14290,N_14115,N_14144);
or U14291 (N_14291,N_14192,N_14166);
nand U14292 (N_14292,N_14081,N_14135);
nand U14293 (N_14293,N_14102,N_14136);
nor U14294 (N_14294,N_14146,N_14091);
nand U14295 (N_14295,N_14037,N_14062);
and U14296 (N_14296,N_14138,N_14158);
and U14297 (N_14297,N_14162,N_14151);
and U14298 (N_14298,N_14032,N_14099);
or U14299 (N_14299,N_14090,N_14128);
nor U14300 (N_14300,N_14099,N_14132);
and U14301 (N_14301,N_14001,N_14065);
nand U14302 (N_14302,N_14172,N_14134);
and U14303 (N_14303,N_14042,N_14107);
nand U14304 (N_14304,N_14078,N_14177);
and U14305 (N_14305,N_14012,N_14115);
nand U14306 (N_14306,N_14095,N_14156);
and U14307 (N_14307,N_14004,N_14065);
xor U14308 (N_14308,N_14085,N_14094);
and U14309 (N_14309,N_14024,N_14126);
and U14310 (N_14310,N_14041,N_14170);
nand U14311 (N_14311,N_14090,N_14120);
xnor U14312 (N_14312,N_14099,N_14157);
and U14313 (N_14313,N_14170,N_14050);
and U14314 (N_14314,N_14110,N_14173);
nor U14315 (N_14315,N_14020,N_14064);
or U14316 (N_14316,N_14065,N_14194);
xor U14317 (N_14317,N_14002,N_14178);
nand U14318 (N_14318,N_14117,N_14186);
nand U14319 (N_14319,N_14152,N_14068);
and U14320 (N_14320,N_14129,N_14050);
and U14321 (N_14321,N_14048,N_14173);
and U14322 (N_14322,N_14156,N_14010);
or U14323 (N_14323,N_14012,N_14076);
and U14324 (N_14324,N_14176,N_14086);
nor U14325 (N_14325,N_14020,N_14037);
or U14326 (N_14326,N_14192,N_14022);
xnor U14327 (N_14327,N_14155,N_14128);
or U14328 (N_14328,N_14025,N_14133);
nand U14329 (N_14329,N_14064,N_14030);
xnor U14330 (N_14330,N_14168,N_14039);
nand U14331 (N_14331,N_14131,N_14188);
nand U14332 (N_14332,N_14110,N_14139);
xor U14333 (N_14333,N_14071,N_14000);
nand U14334 (N_14334,N_14117,N_14142);
and U14335 (N_14335,N_14189,N_14057);
or U14336 (N_14336,N_14114,N_14092);
nor U14337 (N_14337,N_14032,N_14041);
and U14338 (N_14338,N_14049,N_14087);
or U14339 (N_14339,N_14129,N_14045);
and U14340 (N_14340,N_14186,N_14183);
or U14341 (N_14341,N_14020,N_14057);
or U14342 (N_14342,N_14117,N_14088);
nor U14343 (N_14343,N_14094,N_14133);
or U14344 (N_14344,N_14053,N_14100);
xnor U14345 (N_14345,N_14187,N_14182);
or U14346 (N_14346,N_14054,N_14074);
xor U14347 (N_14347,N_14152,N_14155);
xnor U14348 (N_14348,N_14096,N_14191);
nand U14349 (N_14349,N_14111,N_14123);
xnor U14350 (N_14350,N_14044,N_14167);
and U14351 (N_14351,N_14093,N_14007);
xor U14352 (N_14352,N_14000,N_14035);
and U14353 (N_14353,N_14121,N_14155);
nor U14354 (N_14354,N_14107,N_14192);
xor U14355 (N_14355,N_14146,N_14044);
nor U14356 (N_14356,N_14145,N_14004);
nand U14357 (N_14357,N_14053,N_14060);
xnor U14358 (N_14358,N_14193,N_14050);
nand U14359 (N_14359,N_14164,N_14152);
nand U14360 (N_14360,N_14098,N_14110);
xnor U14361 (N_14361,N_14173,N_14078);
or U14362 (N_14362,N_14048,N_14008);
and U14363 (N_14363,N_14084,N_14018);
nor U14364 (N_14364,N_14031,N_14017);
nor U14365 (N_14365,N_14010,N_14146);
or U14366 (N_14366,N_14101,N_14022);
nor U14367 (N_14367,N_14139,N_14024);
xnor U14368 (N_14368,N_14083,N_14049);
xor U14369 (N_14369,N_14075,N_14085);
or U14370 (N_14370,N_14129,N_14126);
nand U14371 (N_14371,N_14089,N_14010);
or U14372 (N_14372,N_14130,N_14010);
xnor U14373 (N_14373,N_14136,N_14101);
nor U14374 (N_14374,N_14095,N_14096);
nand U14375 (N_14375,N_14009,N_14033);
and U14376 (N_14376,N_14047,N_14127);
and U14377 (N_14377,N_14012,N_14191);
nor U14378 (N_14378,N_14022,N_14028);
or U14379 (N_14379,N_14019,N_14091);
and U14380 (N_14380,N_14048,N_14010);
nor U14381 (N_14381,N_14113,N_14105);
or U14382 (N_14382,N_14100,N_14180);
or U14383 (N_14383,N_14191,N_14090);
nor U14384 (N_14384,N_14184,N_14039);
nor U14385 (N_14385,N_14075,N_14031);
nor U14386 (N_14386,N_14135,N_14196);
or U14387 (N_14387,N_14112,N_14083);
xor U14388 (N_14388,N_14132,N_14093);
xor U14389 (N_14389,N_14098,N_14118);
or U14390 (N_14390,N_14142,N_14008);
nor U14391 (N_14391,N_14027,N_14093);
and U14392 (N_14392,N_14140,N_14104);
or U14393 (N_14393,N_14084,N_14131);
nor U14394 (N_14394,N_14090,N_14041);
nand U14395 (N_14395,N_14074,N_14148);
and U14396 (N_14396,N_14037,N_14023);
or U14397 (N_14397,N_14172,N_14182);
nand U14398 (N_14398,N_14185,N_14089);
nand U14399 (N_14399,N_14124,N_14128);
or U14400 (N_14400,N_14223,N_14329);
and U14401 (N_14401,N_14280,N_14203);
and U14402 (N_14402,N_14265,N_14228);
and U14403 (N_14403,N_14248,N_14397);
and U14404 (N_14404,N_14244,N_14285);
nand U14405 (N_14405,N_14281,N_14217);
or U14406 (N_14406,N_14387,N_14344);
nand U14407 (N_14407,N_14235,N_14355);
or U14408 (N_14408,N_14332,N_14300);
or U14409 (N_14409,N_14342,N_14345);
nor U14410 (N_14410,N_14314,N_14295);
xor U14411 (N_14411,N_14252,N_14386);
xor U14412 (N_14412,N_14319,N_14219);
xor U14413 (N_14413,N_14350,N_14242);
nand U14414 (N_14414,N_14239,N_14211);
or U14415 (N_14415,N_14218,N_14269);
or U14416 (N_14416,N_14233,N_14322);
and U14417 (N_14417,N_14277,N_14230);
or U14418 (N_14418,N_14288,N_14255);
or U14419 (N_14419,N_14356,N_14226);
nand U14420 (N_14420,N_14245,N_14385);
nor U14421 (N_14421,N_14290,N_14257);
and U14422 (N_14422,N_14351,N_14298);
and U14423 (N_14423,N_14343,N_14282);
nor U14424 (N_14424,N_14380,N_14313);
and U14425 (N_14425,N_14250,N_14394);
xnor U14426 (N_14426,N_14354,N_14278);
nor U14427 (N_14427,N_14320,N_14232);
or U14428 (N_14428,N_14297,N_14229);
or U14429 (N_14429,N_14370,N_14327);
and U14430 (N_14430,N_14365,N_14212);
nor U14431 (N_14431,N_14268,N_14373);
and U14432 (N_14432,N_14309,N_14306);
and U14433 (N_14433,N_14213,N_14367);
nor U14434 (N_14434,N_14305,N_14347);
xnor U14435 (N_14435,N_14393,N_14287);
nor U14436 (N_14436,N_14270,N_14358);
xor U14437 (N_14437,N_14384,N_14346);
and U14438 (N_14438,N_14307,N_14312);
nor U14439 (N_14439,N_14237,N_14264);
and U14440 (N_14440,N_14272,N_14204);
and U14441 (N_14441,N_14392,N_14341);
and U14442 (N_14442,N_14321,N_14304);
nor U14443 (N_14443,N_14366,N_14378);
nand U14444 (N_14444,N_14353,N_14263);
nor U14445 (N_14445,N_14205,N_14396);
and U14446 (N_14446,N_14241,N_14202);
xor U14447 (N_14447,N_14208,N_14337);
or U14448 (N_14448,N_14249,N_14227);
nor U14449 (N_14449,N_14390,N_14294);
and U14450 (N_14450,N_14225,N_14299);
xor U14451 (N_14451,N_14286,N_14262);
nor U14452 (N_14452,N_14231,N_14361);
nand U14453 (N_14453,N_14301,N_14359);
or U14454 (N_14454,N_14325,N_14383);
xor U14455 (N_14455,N_14224,N_14243);
nand U14456 (N_14456,N_14238,N_14357);
and U14457 (N_14457,N_14210,N_14234);
and U14458 (N_14458,N_14381,N_14362);
nand U14459 (N_14459,N_14256,N_14247);
nand U14460 (N_14460,N_14308,N_14291);
xnor U14461 (N_14461,N_14363,N_14283);
nor U14462 (N_14462,N_14330,N_14258);
nand U14463 (N_14463,N_14302,N_14303);
nor U14464 (N_14464,N_14376,N_14316);
nand U14465 (N_14465,N_14275,N_14382);
or U14466 (N_14466,N_14273,N_14324);
and U14467 (N_14467,N_14310,N_14331);
xor U14468 (N_14468,N_14289,N_14377);
and U14469 (N_14469,N_14292,N_14352);
nor U14470 (N_14470,N_14260,N_14334);
nand U14471 (N_14471,N_14279,N_14240);
xor U14472 (N_14472,N_14220,N_14389);
or U14473 (N_14473,N_14338,N_14293);
nor U14474 (N_14474,N_14221,N_14388);
xnor U14475 (N_14475,N_14251,N_14375);
xnor U14476 (N_14476,N_14391,N_14399);
and U14477 (N_14477,N_14271,N_14214);
nor U14478 (N_14478,N_14222,N_14317);
nor U14479 (N_14479,N_14209,N_14254);
xor U14480 (N_14480,N_14369,N_14335);
or U14481 (N_14481,N_14318,N_14236);
or U14482 (N_14482,N_14216,N_14328);
or U14483 (N_14483,N_14261,N_14276);
nor U14484 (N_14484,N_14326,N_14348);
nand U14485 (N_14485,N_14215,N_14395);
or U14486 (N_14486,N_14340,N_14259);
and U14487 (N_14487,N_14266,N_14207);
and U14488 (N_14488,N_14371,N_14284);
and U14489 (N_14489,N_14246,N_14368);
and U14490 (N_14490,N_14253,N_14374);
or U14491 (N_14491,N_14379,N_14336);
nor U14492 (N_14492,N_14201,N_14315);
xor U14493 (N_14493,N_14349,N_14206);
or U14494 (N_14494,N_14398,N_14200);
or U14495 (N_14495,N_14364,N_14339);
nor U14496 (N_14496,N_14323,N_14333);
and U14497 (N_14497,N_14274,N_14360);
and U14498 (N_14498,N_14372,N_14311);
or U14499 (N_14499,N_14267,N_14296);
nor U14500 (N_14500,N_14293,N_14223);
and U14501 (N_14501,N_14380,N_14292);
and U14502 (N_14502,N_14212,N_14250);
nor U14503 (N_14503,N_14273,N_14296);
and U14504 (N_14504,N_14342,N_14304);
or U14505 (N_14505,N_14306,N_14276);
nand U14506 (N_14506,N_14375,N_14353);
xor U14507 (N_14507,N_14262,N_14343);
xnor U14508 (N_14508,N_14203,N_14224);
xnor U14509 (N_14509,N_14342,N_14253);
or U14510 (N_14510,N_14321,N_14250);
xnor U14511 (N_14511,N_14395,N_14374);
nor U14512 (N_14512,N_14376,N_14384);
nand U14513 (N_14513,N_14376,N_14240);
nand U14514 (N_14514,N_14373,N_14336);
and U14515 (N_14515,N_14214,N_14260);
and U14516 (N_14516,N_14247,N_14273);
xor U14517 (N_14517,N_14390,N_14324);
xnor U14518 (N_14518,N_14274,N_14364);
nand U14519 (N_14519,N_14283,N_14259);
nand U14520 (N_14520,N_14304,N_14306);
nand U14521 (N_14521,N_14255,N_14239);
nand U14522 (N_14522,N_14398,N_14392);
and U14523 (N_14523,N_14355,N_14290);
xnor U14524 (N_14524,N_14272,N_14277);
xor U14525 (N_14525,N_14254,N_14267);
or U14526 (N_14526,N_14309,N_14228);
xor U14527 (N_14527,N_14277,N_14237);
nor U14528 (N_14528,N_14335,N_14264);
nand U14529 (N_14529,N_14282,N_14270);
nand U14530 (N_14530,N_14319,N_14295);
nand U14531 (N_14531,N_14269,N_14287);
or U14532 (N_14532,N_14207,N_14367);
and U14533 (N_14533,N_14251,N_14329);
or U14534 (N_14534,N_14386,N_14378);
and U14535 (N_14535,N_14363,N_14219);
nand U14536 (N_14536,N_14312,N_14209);
and U14537 (N_14537,N_14235,N_14217);
nand U14538 (N_14538,N_14207,N_14365);
xor U14539 (N_14539,N_14271,N_14285);
nand U14540 (N_14540,N_14378,N_14211);
and U14541 (N_14541,N_14265,N_14394);
nand U14542 (N_14542,N_14249,N_14362);
nand U14543 (N_14543,N_14339,N_14314);
nand U14544 (N_14544,N_14318,N_14202);
nor U14545 (N_14545,N_14312,N_14248);
and U14546 (N_14546,N_14340,N_14313);
nand U14547 (N_14547,N_14245,N_14281);
nor U14548 (N_14548,N_14264,N_14340);
and U14549 (N_14549,N_14380,N_14278);
nor U14550 (N_14550,N_14232,N_14336);
xor U14551 (N_14551,N_14257,N_14204);
and U14552 (N_14552,N_14268,N_14204);
nand U14553 (N_14553,N_14244,N_14345);
or U14554 (N_14554,N_14260,N_14220);
or U14555 (N_14555,N_14335,N_14268);
nand U14556 (N_14556,N_14214,N_14204);
or U14557 (N_14557,N_14383,N_14228);
nor U14558 (N_14558,N_14236,N_14276);
and U14559 (N_14559,N_14358,N_14289);
nand U14560 (N_14560,N_14340,N_14362);
and U14561 (N_14561,N_14225,N_14384);
xnor U14562 (N_14562,N_14295,N_14248);
and U14563 (N_14563,N_14389,N_14310);
and U14564 (N_14564,N_14307,N_14351);
and U14565 (N_14565,N_14235,N_14264);
or U14566 (N_14566,N_14269,N_14278);
and U14567 (N_14567,N_14209,N_14396);
or U14568 (N_14568,N_14305,N_14204);
nand U14569 (N_14569,N_14316,N_14348);
xnor U14570 (N_14570,N_14346,N_14310);
or U14571 (N_14571,N_14362,N_14304);
or U14572 (N_14572,N_14213,N_14293);
xnor U14573 (N_14573,N_14268,N_14235);
and U14574 (N_14574,N_14228,N_14307);
nand U14575 (N_14575,N_14304,N_14285);
or U14576 (N_14576,N_14313,N_14395);
and U14577 (N_14577,N_14350,N_14335);
nor U14578 (N_14578,N_14376,N_14336);
and U14579 (N_14579,N_14373,N_14234);
or U14580 (N_14580,N_14397,N_14388);
or U14581 (N_14581,N_14216,N_14267);
and U14582 (N_14582,N_14280,N_14306);
nor U14583 (N_14583,N_14342,N_14243);
nand U14584 (N_14584,N_14250,N_14288);
nand U14585 (N_14585,N_14357,N_14296);
or U14586 (N_14586,N_14238,N_14233);
nor U14587 (N_14587,N_14394,N_14303);
nand U14588 (N_14588,N_14341,N_14373);
nand U14589 (N_14589,N_14223,N_14270);
and U14590 (N_14590,N_14209,N_14349);
xnor U14591 (N_14591,N_14241,N_14303);
nor U14592 (N_14592,N_14317,N_14373);
or U14593 (N_14593,N_14327,N_14396);
or U14594 (N_14594,N_14220,N_14215);
nor U14595 (N_14595,N_14205,N_14327);
xnor U14596 (N_14596,N_14324,N_14227);
xnor U14597 (N_14597,N_14363,N_14333);
and U14598 (N_14598,N_14254,N_14265);
nand U14599 (N_14599,N_14252,N_14350);
xor U14600 (N_14600,N_14575,N_14516);
and U14601 (N_14601,N_14520,N_14579);
nor U14602 (N_14602,N_14517,N_14463);
and U14603 (N_14603,N_14522,N_14481);
nor U14604 (N_14604,N_14596,N_14503);
nand U14605 (N_14605,N_14582,N_14421);
xnor U14606 (N_14606,N_14493,N_14598);
nor U14607 (N_14607,N_14453,N_14411);
xnor U14608 (N_14608,N_14537,N_14477);
or U14609 (N_14609,N_14494,N_14490);
or U14610 (N_14610,N_14542,N_14551);
nor U14611 (N_14611,N_14590,N_14573);
nand U14612 (N_14612,N_14489,N_14416);
and U14613 (N_14613,N_14508,N_14450);
and U14614 (N_14614,N_14580,N_14595);
xnor U14615 (N_14615,N_14548,N_14514);
nand U14616 (N_14616,N_14418,N_14402);
and U14617 (N_14617,N_14465,N_14563);
or U14618 (N_14618,N_14518,N_14586);
or U14619 (N_14619,N_14510,N_14547);
nand U14620 (N_14620,N_14435,N_14445);
and U14621 (N_14621,N_14535,N_14546);
and U14622 (N_14622,N_14506,N_14419);
nand U14623 (N_14623,N_14544,N_14485);
nand U14624 (N_14624,N_14429,N_14521);
xor U14625 (N_14625,N_14552,N_14472);
or U14626 (N_14626,N_14570,N_14425);
nor U14627 (N_14627,N_14519,N_14467);
nand U14628 (N_14628,N_14484,N_14457);
and U14629 (N_14629,N_14536,N_14427);
and U14630 (N_14630,N_14559,N_14462);
nor U14631 (N_14631,N_14431,N_14599);
nand U14632 (N_14632,N_14515,N_14476);
or U14633 (N_14633,N_14561,N_14422);
or U14634 (N_14634,N_14513,N_14434);
or U14635 (N_14635,N_14432,N_14415);
xor U14636 (N_14636,N_14451,N_14577);
nand U14637 (N_14637,N_14576,N_14486);
nor U14638 (N_14638,N_14562,N_14446);
and U14639 (N_14639,N_14567,N_14504);
or U14640 (N_14640,N_14498,N_14524);
and U14641 (N_14641,N_14528,N_14568);
xnor U14642 (N_14642,N_14420,N_14554);
xor U14643 (N_14643,N_14461,N_14400);
nor U14644 (N_14644,N_14594,N_14491);
nand U14645 (N_14645,N_14479,N_14557);
nand U14646 (N_14646,N_14505,N_14483);
and U14647 (N_14647,N_14525,N_14458);
or U14648 (N_14648,N_14540,N_14409);
nand U14649 (N_14649,N_14584,N_14482);
nand U14650 (N_14650,N_14452,N_14478);
and U14651 (N_14651,N_14589,N_14456);
or U14652 (N_14652,N_14593,N_14556);
or U14653 (N_14653,N_14473,N_14541);
and U14654 (N_14654,N_14440,N_14549);
and U14655 (N_14655,N_14558,N_14469);
or U14656 (N_14656,N_14454,N_14588);
xnor U14657 (N_14657,N_14401,N_14436);
nand U14658 (N_14658,N_14474,N_14449);
nor U14659 (N_14659,N_14480,N_14414);
nor U14660 (N_14660,N_14550,N_14464);
and U14661 (N_14661,N_14443,N_14511);
xnor U14662 (N_14662,N_14499,N_14587);
nor U14663 (N_14663,N_14459,N_14428);
xor U14664 (N_14664,N_14532,N_14531);
nand U14665 (N_14665,N_14533,N_14555);
nand U14666 (N_14666,N_14527,N_14408);
and U14667 (N_14667,N_14572,N_14412);
xor U14668 (N_14668,N_14496,N_14404);
nor U14669 (N_14669,N_14410,N_14539);
and U14670 (N_14670,N_14403,N_14437);
nor U14671 (N_14671,N_14553,N_14569);
xor U14672 (N_14672,N_14574,N_14471);
nand U14673 (N_14673,N_14438,N_14413);
xor U14674 (N_14674,N_14545,N_14501);
nor U14675 (N_14675,N_14442,N_14475);
nor U14676 (N_14676,N_14488,N_14592);
and U14677 (N_14677,N_14460,N_14581);
or U14678 (N_14678,N_14406,N_14500);
nand U14679 (N_14679,N_14507,N_14526);
or U14680 (N_14680,N_14433,N_14466);
and U14681 (N_14681,N_14566,N_14405);
xnor U14682 (N_14682,N_14441,N_14495);
and U14683 (N_14683,N_14523,N_14560);
and U14684 (N_14684,N_14407,N_14417);
and U14685 (N_14685,N_14530,N_14468);
or U14686 (N_14686,N_14487,N_14543);
and U14687 (N_14687,N_14591,N_14512);
xnor U14688 (N_14688,N_14597,N_14447);
nor U14689 (N_14689,N_14444,N_14448);
and U14690 (N_14690,N_14502,N_14585);
xor U14691 (N_14691,N_14470,N_14424);
and U14692 (N_14692,N_14564,N_14439);
or U14693 (N_14693,N_14538,N_14534);
xor U14694 (N_14694,N_14571,N_14565);
nand U14695 (N_14695,N_14509,N_14455);
xor U14696 (N_14696,N_14497,N_14430);
or U14697 (N_14697,N_14578,N_14423);
and U14698 (N_14698,N_14492,N_14529);
nand U14699 (N_14699,N_14426,N_14583);
xnor U14700 (N_14700,N_14591,N_14500);
nor U14701 (N_14701,N_14543,N_14578);
xnor U14702 (N_14702,N_14496,N_14590);
and U14703 (N_14703,N_14490,N_14485);
or U14704 (N_14704,N_14569,N_14477);
xnor U14705 (N_14705,N_14596,N_14480);
nor U14706 (N_14706,N_14573,N_14551);
and U14707 (N_14707,N_14430,N_14484);
or U14708 (N_14708,N_14478,N_14501);
nor U14709 (N_14709,N_14582,N_14455);
or U14710 (N_14710,N_14460,N_14446);
or U14711 (N_14711,N_14594,N_14529);
nand U14712 (N_14712,N_14453,N_14594);
xnor U14713 (N_14713,N_14417,N_14590);
nand U14714 (N_14714,N_14581,N_14432);
xor U14715 (N_14715,N_14429,N_14534);
nand U14716 (N_14716,N_14571,N_14591);
nand U14717 (N_14717,N_14476,N_14542);
xnor U14718 (N_14718,N_14529,N_14445);
and U14719 (N_14719,N_14547,N_14590);
xor U14720 (N_14720,N_14443,N_14528);
or U14721 (N_14721,N_14439,N_14455);
or U14722 (N_14722,N_14458,N_14558);
xor U14723 (N_14723,N_14437,N_14453);
and U14724 (N_14724,N_14420,N_14561);
nor U14725 (N_14725,N_14527,N_14487);
or U14726 (N_14726,N_14481,N_14472);
nor U14727 (N_14727,N_14573,N_14509);
nand U14728 (N_14728,N_14452,N_14599);
nand U14729 (N_14729,N_14439,N_14507);
and U14730 (N_14730,N_14472,N_14586);
and U14731 (N_14731,N_14510,N_14414);
nor U14732 (N_14732,N_14441,N_14467);
or U14733 (N_14733,N_14418,N_14515);
and U14734 (N_14734,N_14535,N_14483);
and U14735 (N_14735,N_14495,N_14432);
xnor U14736 (N_14736,N_14570,N_14526);
xor U14737 (N_14737,N_14587,N_14560);
nand U14738 (N_14738,N_14409,N_14541);
nor U14739 (N_14739,N_14408,N_14568);
nor U14740 (N_14740,N_14462,N_14538);
nand U14741 (N_14741,N_14455,N_14410);
or U14742 (N_14742,N_14443,N_14561);
or U14743 (N_14743,N_14592,N_14476);
nand U14744 (N_14744,N_14564,N_14485);
nand U14745 (N_14745,N_14471,N_14571);
xnor U14746 (N_14746,N_14422,N_14447);
and U14747 (N_14747,N_14494,N_14515);
or U14748 (N_14748,N_14503,N_14556);
xnor U14749 (N_14749,N_14597,N_14450);
and U14750 (N_14750,N_14533,N_14438);
and U14751 (N_14751,N_14531,N_14429);
or U14752 (N_14752,N_14498,N_14436);
and U14753 (N_14753,N_14475,N_14421);
and U14754 (N_14754,N_14544,N_14458);
nor U14755 (N_14755,N_14533,N_14531);
or U14756 (N_14756,N_14484,N_14593);
or U14757 (N_14757,N_14453,N_14464);
or U14758 (N_14758,N_14519,N_14507);
nor U14759 (N_14759,N_14580,N_14555);
nor U14760 (N_14760,N_14594,N_14579);
xnor U14761 (N_14761,N_14449,N_14532);
nand U14762 (N_14762,N_14402,N_14541);
nand U14763 (N_14763,N_14511,N_14514);
nand U14764 (N_14764,N_14588,N_14543);
nand U14765 (N_14765,N_14596,N_14598);
or U14766 (N_14766,N_14505,N_14508);
and U14767 (N_14767,N_14462,N_14580);
and U14768 (N_14768,N_14494,N_14412);
and U14769 (N_14769,N_14443,N_14446);
nor U14770 (N_14770,N_14537,N_14565);
nor U14771 (N_14771,N_14446,N_14584);
or U14772 (N_14772,N_14402,N_14442);
and U14773 (N_14773,N_14597,N_14574);
xnor U14774 (N_14774,N_14490,N_14532);
nor U14775 (N_14775,N_14428,N_14441);
and U14776 (N_14776,N_14460,N_14405);
xor U14777 (N_14777,N_14426,N_14445);
or U14778 (N_14778,N_14402,N_14414);
and U14779 (N_14779,N_14445,N_14486);
or U14780 (N_14780,N_14461,N_14478);
xor U14781 (N_14781,N_14553,N_14525);
or U14782 (N_14782,N_14511,N_14480);
xor U14783 (N_14783,N_14485,N_14435);
and U14784 (N_14784,N_14443,N_14590);
nand U14785 (N_14785,N_14583,N_14432);
nor U14786 (N_14786,N_14496,N_14572);
and U14787 (N_14787,N_14493,N_14435);
nand U14788 (N_14788,N_14551,N_14483);
nand U14789 (N_14789,N_14479,N_14452);
or U14790 (N_14790,N_14566,N_14584);
and U14791 (N_14791,N_14567,N_14412);
nand U14792 (N_14792,N_14521,N_14456);
xnor U14793 (N_14793,N_14443,N_14484);
nor U14794 (N_14794,N_14582,N_14441);
nor U14795 (N_14795,N_14562,N_14472);
nor U14796 (N_14796,N_14536,N_14570);
xor U14797 (N_14797,N_14411,N_14515);
nor U14798 (N_14798,N_14541,N_14532);
nand U14799 (N_14799,N_14561,N_14486);
and U14800 (N_14800,N_14641,N_14784);
or U14801 (N_14801,N_14686,N_14718);
and U14802 (N_14802,N_14668,N_14735);
xor U14803 (N_14803,N_14617,N_14780);
nand U14804 (N_14804,N_14707,N_14645);
nand U14805 (N_14805,N_14748,N_14727);
nand U14806 (N_14806,N_14665,N_14675);
xnor U14807 (N_14807,N_14717,N_14737);
nand U14808 (N_14808,N_14782,N_14650);
xnor U14809 (N_14809,N_14740,N_14722);
nand U14810 (N_14810,N_14746,N_14772);
and U14811 (N_14811,N_14794,N_14638);
xnor U14812 (N_14812,N_14630,N_14776);
and U14813 (N_14813,N_14756,N_14655);
or U14814 (N_14814,N_14758,N_14741);
or U14815 (N_14815,N_14683,N_14747);
or U14816 (N_14816,N_14702,N_14607);
or U14817 (N_14817,N_14708,N_14723);
xor U14818 (N_14818,N_14629,N_14695);
or U14819 (N_14819,N_14761,N_14713);
nor U14820 (N_14820,N_14681,N_14777);
nand U14821 (N_14821,N_14688,N_14640);
or U14822 (N_14822,N_14628,N_14646);
and U14823 (N_14823,N_14786,N_14647);
nand U14824 (N_14824,N_14743,N_14687);
xor U14825 (N_14825,N_14604,N_14738);
or U14826 (N_14826,N_14745,N_14651);
nor U14827 (N_14827,N_14724,N_14728);
nand U14828 (N_14828,N_14609,N_14676);
nor U14829 (N_14829,N_14790,N_14616);
nand U14830 (N_14830,N_14669,N_14771);
xnor U14831 (N_14831,N_14781,N_14779);
nor U14832 (N_14832,N_14754,N_14678);
xor U14833 (N_14833,N_14685,N_14760);
nor U14834 (N_14834,N_14763,N_14765);
nor U14835 (N_14835,N_14635,N_14689);
nor U14836 (N_14836,N_14769,N_14697);
or U14837 (N_14837,N_14749,N_14742);
or U14838 (N_14838,N_14666,N_14672);
or U14839 (N_14839,N_14632,N_14658);
xor U14840 (N_14840,N_14710,N_14648);
and U14841 (N_14841,N_14625,N_14791);
xor U14842 (N_14842,N_14671,N_14732);
nor U14843 (N_14843,N_14799,N_14762);
or U14844 (N_14844,N_14634,N_14706);
nor U14845 (N_14845,N_14736,N_14701);
nor U14846 (N_14846,N_14788,N_14690);
nor U14847 (N_14847,N_14659,N_14792);
or U14848 (N_14848,N_14775,N_14611);
nand U14849 (N_14849,N_14642,N_14751);
xor U14850 (N_14850,N_14661,N_14637);
nand U14851 (N_14851,N_14730,N_14753);
nor U14852 (N_14852,N_14627,N_14692);
nor U14853 (N_14853,N_14606,N_14673);
nor U14854 (N_14854,N_14764,N_14608);
or U14855 (N_14855,N_14798,N_14662);
nand U14856 (N_14856,N_14752,N_14783);
nor U14857 (N_14857,N_14739,N_14795);
nor U14858 (N_14858,N_14660,N_14789);
nor U14859 (N_14859,N_14601,N_14774);
and U14860 (N_14860,N_14773,N_14704);
nand U14861 (N_14861,N_14750,N_14694);
and U14862 (N_14862,N_14664,N_14652);
nor U14863 (N_14863,N_14677,N_14602);
or U14864 (N_14864,N_14711,N_14684);
or U14865 (N_14865,N_14721,N_14613);
nor U14866 (N_14866,N_14605,N_14654);
nand U14867 (N_14867,N_14623,N_14663);
or U14868 (N_14868,N_14680,N_14759);
nor U14869 (N_14869,N_14649,N_14703);
or U14870 (N_14870,N_14719,N_14767);
nor U14871 (N_14871,N_14633,N_14778);
or U14872 (N_14872,N_14653,N_14624);
xnor U14873 (N_14873,N_14643,N_14696);
nand U14874 (N_14874,N_14656,N_14715);
xor U14875 (N_14875,N_14714,N_14705);
nor U14876 (N_14876,N_14700,N_14644);
and U14877 (N_14877,N_14631,N_14709);
nand U14878 (N_14878,N_14619,N_14612);
xnor U14879 (N_14879,N_14618,N_14725);
and U14880 (N_14880,N_14793,N_14614);
xnor U14881 (N_14881,N_14766,N_14639);
or U14882 (N_14882,N_14636,N_14670);
and U14883 (N_14883,N_14734,N_14720);
nor U14884 (N_14884,N_14768,N_14716);
xnor U14885 (N_14885,N_14744,N_14674);
or U14886 (N_14886,N_14615,N_14731);
nor U14887 (N_14887,N_14729,N_14682);
xnor U14888 (N_14888,N_14699,N_14693);
nand U14889 (N_14889,N_14620,N_14785);
nor U14890 (N_14890,N_14621,N_14610);
nand U14891 (N_14891,N_14770,N_14757);
and U14892 (N_14892,N_14755,N_14679);
xor U14893 (N_14893,N_14603,N_14726);
or U14894 (N_14894,N_14787,N_14733);
xnor U14895 (N_14895,N_14600,N_14626);
and U14896 (N_14896,N_14667,N_14712);
nor U14897 (N_14897,N_14657,N_14691);
nor U14898 (N_14898,N_14797,N_14698);
and U14899 (N_14899,N_14796,N_14622);
or U14900 (N_14900,N_14711,N_14730);
nor U14901 (N_14901,N_14685,N_14788);
xor U14902 (N_14902,N_14613,N_14755);
nor U14903 (N_14903,N_14710,N_14776);
xor U14904 (N_14904,N_14637,N_14607);
xnor U14905 (N_14905,N_14750,N_14728);
nand U14906 (N_14906,N_14662,N_14760);
nor U14907 (N_14907,N_14758,N_14749);
nand U14908 (N_14908,N_14691,N_14755);
and U14909 (N_14909,N_14620,N_14700);
and U14910 (N_14910,N_14682,N_14714);
xor U14911 (N_14911,N_14664,N_14766);
or U14912 (N_14912,N_14697,N_14611);
or U14913 (N_14913,N_14668,N_14644);
nor U14914 (N_14914,N_14763,N_14653);
and U14915 (N_14915,N_14672,N_14776);
xnor U14916 (N_14916,N_14771,N_14635);
and U14917 (N_14917,N_14771,N_14674);
xnor U14918 (N_14918,N_14700,N_14664);
nand U14919 (N_14919,N_14603,N_14650);
and U14920 (N_14920,N_14602,N_14633);
nand U14921 (N_14921,N_14668,N_14667);
xor U14922 (N_14922,N_14613,N_14724);
xor U14923 (N_14923,N_14799,N_14789);
nor U14924 (N_14924,N_14642,N_14785);
nand U14925 (N_14925,N_14771,N_14726);
nor U14926 (N_14926,N_14784,N_14738);
or U14927 (N_14927,N_14764,N_14657);
nor U14928 (N_14928,N_14650,N_14724);
or U14929 (N_14929,N_14615,N_14795);
nor U14930 (N_14930,N_14638,N_14641);
or U14931 (N_14931,N_14786,N_14719);
nor U14932 (N_14932,N_14648,N_14673);
or U14933 (N_14933,N_14637,N_14742);
or U14934 (N_14934,N_14657,N_14789);
nand U14935 (N_14935,N_14667,N_14709);
nor U14936 (N_14936,N_14620,N_14671);
nand U14937 (N_14937,N_14692,N_14787);
nand U14938 (N_14938,N_14618,N_14748);
and U14939 (N_14939,N_14666,N_14646);
or U14940 (N_14940,N_14721,N_14682);
nor U14941 (N_14941,N_14702,N_14615);
xor U14942 (N_14942,N_14765,N_14772);
or U14943 (N_14943,N_14635,N_14624);
xor U14944 (N_14944,N_14716,N_14749);
nor U14945 (N_14945,N_14780,N_14763);
or U14946 (N_14946,N_14779,N_14698);
nand U14947 (N_14947,N_14728,N_14773);
xnor U14948 (N_14948,N_14701,N_14605);
or U14949 (N_14949,N_14661,N_14601);
and U14950 (N_14950,N_14723,N_14644);
xor U14951 (N_14951,N_14620,N_14708);
nand U14952 (N_14952,N_14661,N_14626);
nor U14953 (N_14953,N_14667,N_14797);
or U14954 (N_14954,N_14791,N_14675);
or U14955 (N_14955,N_14608,N_14760);
nor U14956 (N_14956,N_14674,N_14769);
or U14957 (N_14957,N_14784,N_14719);
or U14958 (N_14958,N_14625,N_14793);
nand U14959 (N_14959,N_14751,N_14754);
and U14960 (N_14960,N_14795,N_14750);
and U14961 (N_14961,N_14724,N_14742);
or U14962 (N_14962,N_14701,N_14692);
or U14963 (N_14963,N_14621,N_14609);
or U14964 (N_14964,N_14730,N_14775);
nor U14965 (N_14965,N_14767,N_14626);
xor U14966 (N_14966,N_14656,N_14641);
nor U14967 (N_14967,N_14739,N_14777);
and U14968 (N_14968,N_14626,N_14786);
nand U14969 (N_14969,N_14603,N_14700);
and U14970 (N_14970,N_14608,N_14626);
xnor U14971 (N_14971,N_14639,N_14774);
nor U14972 (N_14972,N_14648,N_14681);
nor U14973 (N_14973,N_14798,N_14622);
xnor U14974 (N_14974,N_14748,N_14794);
or U14975 (N_14975,N_14771,N_14649);
and U14976 (N_14976,N_14630,N_14702);
or U14977 (N_14977,N_14648,N_14626);
nand U14978 (N_14978,N_14646,N_14754);
xnor U14979 (N_14979,N_14761,N_14668);
nand U14980 (N_14980,N_14728,N_14791);
or U14981 (N_14981,N_14710,N_14747);
nor U14982 (N_14982,N_14786,N_14645);
nor U14983 (N_14983,N_14699,N_14629);
nor U14984 (N_14984,N_14658,N_14657);
or U14985 (N_14985,N_14608,N_14685);
and U14986 (N_14986,N_14610,N_14753);
nand U14987 (N_14987,N_14796,N_14780);
and U14988 (N_14988,N_14655,N_14686);
nand U14989 (N_14989,N_14730,N_14606);
xor U14990 (N_14990,N_14780,N_14651);
nor U14991 (N_14991,N_14631,N_14719);
xnor U14992 (N_14992,N_14751,N_14641);
nand U14993 (N_14993,N_14789,N_14787);
nor U14994 (N_14994,N_14664,N_14657);
or U14995 (N_14995,N_14631,N_14639);
nor U14996 (N_14996,N_14757,N_14661);
xor U14997 (N_14997,N_14730,N_14700);
and U14998 (N_14998,N_14788,N_14676);
or U14999 (N_14999,N_14606,N_14648);
nand U15000 (N_15000,N_14847,N_14981);
and U15001 (N_15001,N_14883,N_14818);
or U15002 (N_15002,N_14925,N_14899);
nor U15003 (N_15003,N_14909,N_14838);
nand U15004 (N_15004,N_14931,N_14846);
and U15005 (N_15005,N_14831,N_14837);
xor U15006 (N_15006,N_14940,N_14815);
and U15007 (N_15007,N_14907,N_14912);
xor U15008 (N_15008,N_14811,N_14957);
or U15009 (N_15009,N_14984,N_14880);
xnor U15010 (N_15010,N_14827,N_14858);
nand U15011 (N_15011,N_14968,N_14994);
nand U15012 (N_15012,N_14840,N_14870);
nand U15013 (N_15013,N_14897,N_14844);
nand U15014 (N_15014,N_14945,N_14872);
xor U15015 (N_15015,N_14895,N_14871);
and U15016 (N_15016,N_14856,N_14990);
nor U15017 (N_15017,N_14970,N_14973);
nand U15018 (N_15018,N_14841,N_14851);
or U15019 (N_15019,N_14930,N_14857);
or U15020 (N_15020,N_14867,N_14891);
nor U15021 (N_15021,N_14999,N_14836);
nor U15022 (N_15022,N_14866,N_14989);
xnor U15023 (N_15023,N_14876,N_14890);
nor U15024 (N_15024,N_14963,N_14887);
xor U15025 (N_15025,N_14939,N_14821);
nand U15026 (N_15026,N_14881,N_14896);
xnor U15027 (N_15027,N_14991,N_14860);
xnor U15028 (N_15028,N_14974,N_14959);
and U15029 (N_15029,N_14921,N_14893);
nand U15030 (N_15030,N_14910,N_14900);
or U15031 (N_15031,N_14975,N_14853);
or U15032 (N_15032,N_14908,N_14806);
xnor U15033 (N_15033,N_14972,N_14822);
nor U15034 (N_15034,N_14993,N_14809);
nand U15035 (N_15035,N_14926,N_14960);
nor U15036 (N_15036,N_14804,N_14979);
nand U15037 (N_15037,N_14835,N_14850);
xnor U15038 (N_15038,N_14862,N_14944);
nand U15039 (N_15039,N_14854,N_14934);
xnor U15040 (N_15040,N_14885,N_14919);
nor U15041 (N_15041,N_14958,N_14976);
xnor U15042 (N_15042,N_14929,N_14848);
and U15043 (N_15043,N_14879,N_14828);
and U15044 (N_15044,N_14961,N_14859);
or U15045 (N_15045,N_14898,N_14807);
nor U15046 (N_15046,N_14852,N_14955);
nand U15047 (N_15047,N_14820,N_14942);
nand U15048 (N_15048,N_14892,N_14923);
nand U15049 (N_15049,N_14875,N_14980);
xnor U15050 (N_15050,N_14877,N_14878);
and U15051 (N_15051,N_14915,N_14842);
or U15052 (N_15052,N_14916,N_14810);
and U15053 (N_15053,N_14800,N_14918);
or U15054 (N_15054,N_14834,N_14932);
nor U15055 (N_15055,N_14819,N_14953);
nand U15056 (N_15056,N_14965,N_14829);
or U15057 (N_15057,N_14951,N_14987);
or U15058 (N_15058,N_14861,N_14967);
and U15059 (N_15059,N_14969,N_14845);
nor U15060 (N_15060,N_14826,N_14914);
nand U15061 (N_15061,N_14920,N_14865);
nor U15062 (N_15062,N_14855,N_14882);
nor U15063 (N_15063,N_14902,N_14833);
xnor U15064 (N_15064,N_14935,N_14928);
nand U15065 (N_15065,N_14873,N_14943);
and U15066 (N_15066,N_14813,N_14849);
or U15067 (N_15067,N_14997,N_14808);
nor U15068 (N_15068,N_14906,N_14864);
and U15069 (N_15069,N_14941,N_14801);
and U15070 (N_15070,N_14888,N_14956);
or U15071 (N_15071,N_14904,N_14814);
and U15072 (N_15072,N_14830,N_14863);
and U15073 (N_15073,N_14917,N_14982);
xnor U15074 (N_15074,N_14823,N_14817);
nand U15075 (N_15075,N_14913,N_14927);
xnor U15076 (N_15076,N_14983,N_14946);
or U15077 (N_15077,N_14868,N_14985);
nand U15078 (N_15078,N_14839,N_14971);
and U15079 (N_15079,N_14978,N_14824);
or U15080 (N_15080,N_14950,N_14947);
or U15081 (N_15081,N_14924,N_14911);
nand U15082 (N_15082,N_14889,N_14894);
or U15083 (N_15083,N_14998,N_14962);
xnor U15084 (N_15084,N_14964,N_14825);
and U15085 (N_15085,N_14903,N_14901);
nor U15086 (N_15086,N_14803,N_14884);
nand U15087 (N_15087,N_14843,N_14874);
and U15088 (N_15088,N_14938,N_14954);
xnor U15089 (N_15089,N_14933,N_14952);
nand U15090 (N_15090,N_14992,N_14812);
or U15091 (N_15091,N_14937,N_14995);
and U15092 (N_15092,N_14832,N_14988);
nand U15093 (N_15093,N_14966,N_14977);
and U15094 (N_15094,N_14886,N_14986);
xnor U15095 (N_15095,N_14905,N_14996);
nand U15096 (N_15096,N_14805,N_14816);
nor U15097 (N_15097,N_14869,N_14802);
and U15098 (N_15098,N_14949,N_14948);
xnor U15099 (N_15099,N_14922,N_14936);
or U15100 (N_15100,N_14943,N_14828);
nor U15101 (N_15101,N_14893,N_14820);
and U15102 (N_15102,N_14945,N_14882);
or U15103 (N_15103,N_14863,N_14971);
xor U15104 (N_15104,N_14969,N_14834);
and U15105 (N_15105,N_14843,N_14933);
nor U15106 (N_15106,N_14948,N_14890);
xor U15107 (N_15107,N_14948,N_14835);
or U15108 (N_15108,N_14910,N_14947);
nor U15109 (N_15109,N_14844,N_14970);
or U15110 (N_15110,N_14818,N_14927);
nand U15111 (N_15111,N_14974,N_14872);
or U15112 (N_15112,N_14819,N_14952);
or U15113 (N_15113,N_14842,N_14883);
nor U15114 (N_15114,N_14847,N_14987);
xnor U15115 (N_15115,N_14939,N_14887);
nor U15116 (N_15116,N_14890,N_14867);
or U15117 (N_15117,N_14983,N_14989);
xor U15118 (N_15118,N_14903,N_14987);
nor U15119 (N_15119,N_14983,N_14861);
and U15120 (N_15120,N_14997,N_14882);
nor U15121 (N_15121,N_14821,N_14964);
or U15122 (N_15122,N_14945,N_14893);
xor U15123 (N_15123,N_14806,N_14965);
and U15124 (N_15124,N_14953,N_14853);
or U15125 (N_15125,N_14877,N_14906);
or U15126 (N_15126,N_14847,N_14820);
nand U15127 (N_15127,N_14841,N_14919);
xnor U15128 (N_15128,N_14864,N_14894);
nor U15129 (N_15129,N_14935,N_14842);
xnor U15130 (N_15130,N_14866,N_14843);
nand U15131 (N_15131,N_14951,N_14939);
nor U15132 (N_15132,N_14876,N_14982);
nor U15133 (N_15133,N_14988,N_14923);
nand U15134 (N_15134,N_14909,N_14999);
or U15135 (N_15135,N_14993,N_14896);
or U15136 (N_15136,N_14812,N_14868);
nor U15137 (N_15137,N_14823,N_14845);
xnor U15138 (N_15138,N_14851,N_14940);
and U15139 (N_15139,N_14866,N_14807);
nand U15140 (N_15140,N_14951,N_14974);
xnor U15141 (N_15141,N_14861,N_14988);
nand U15142 (N_15142,N_14999,N_14993);
xor U15143 (N_15143,N_14890,N_14844);
nand U15144 (N_15144,N_14835,N_14817);
nor U15145 (N_15145,N_14828,N_14816);
or U15146 (N_15146,N_14804,N_14872);
xnor U15147 (N_15147,N_14823,N_14981);
nand U15148 (N_15148,N_14897,N_14976);
and U15149 (N_15149,N_14985,N_14945);
nor U15150 (N_15150,N_14898,N_14976);
nor U15151 (N_15151,N_14850,N_14983);
and U15152 (N_15152,N_14896,N_14954);
xor U15153 (N_15153,N_14915,N_14885);
or U15154 (N_15154,N_14943,N_14949);
xor U15155 (N_15155,N_14836,N_14828);
or U15156 (N_15156,N_14934,N_14931);
nand U15157 (N_15157,N_14928,N_14888);
and U15158 (N_15158,N_14889,N_14967);
nor U15159 (N_15159,N_14805,N_14947);
nor U15160 (N_15160,N_14806,N_14844);
nor U15161 (N_15161,N_14867,N_14847);
and U15162 (N_15162,N_14840,N_14849);
and U15163 (N_15163,N_14930,N_14905);
nand U15164 (N_15164,N_14965,N_14971);
and U15165 (N_15165,N_14867,N_14868);
xor U15166 (N_15166,N_14876,N_14879);
nor U15167 (N_15167,N_14936,N_14894);
xor U15168 (N_15168,N_14873,N_14874);
or U15169 (N_15169,N_14923,N_14941);
nor U15170 (N_15170,N_14888,N_14880);
or U15171 (N_15171,N_14828,N_14923);
nand U15172 (N_15172,N_14805,N_14895);
xor U15173 (N_15173,N_14832,N_14862);
xor U15174 (N_15174,N_14973,N_14845);
xnor U15175 (N_15175,N_14988,N_14956);
and U15176 (N_15176,N_14885,N_14851);
and U15177 (N_15177,N_14826,N_14988);
or U15178 (N_15178,N_14874,N_14930);
xor U15179 (N_15179,N_14876,N_14815);
nor U15180 (N_15180,N_14927,N_14940);
or U15181 (N_15181,N_14996,N_14958);
nand U15182 (N_15182,N_14858,N_14996);
nand U15183 (N_15183,N_14888,N_14986);
nor U15184 (N_15184,N_14928,N_14987);
nand U15185 (N_15185,N_14801,N_14983);
and U15186 (N_15186,N_14999,N_14935);
and U15187 (N_15187,N_14889,N_14901);
nor U15188 (N_15188,N_14841,N_14855);
and U15189 (N_15189,N_14978,N_14922);
xor U15190 (N_15190,N_14971,N_14819);
or U15191 (N_15191,N_14921,N_14920);
nor U15192 (N_15192,N_14823,N_14968);
nor U15193 (N_15193,N_14805,N_14817);
nand U15194 (N_15194,N_14964,N_14883);
nand U15195 (N_15195,N_14870,N_14937);
nand U15196 (N_15196,N_14936,N_14899);
nor U15197 (N_15197,N_14858,N_14990);
or U15198 (N_15198,N_14836,N_14958);
nor U15199 (N_15199,N_14852,N_14973);
nor U15200 (N_15200,N_15190,N_15106);
or U15201 (N_15201,N_15000,N_15136);
nand U15202 (N_15202,N_15186,N_15109);
and U15203 (N_15203,N_15161,N_15128);
xnor U15204 (N_15204,N_15076,N_15168);
nor U15205 (N_15205,N_15146,N_15165);
nor U15206 (N_15206,N_15097,N_15108);
and U15207 (N_15207,N_15145,N_15044);
and U15208 (N_15208,N_15127,N_15079);
and U15209 (N_15209,N_15035,N_15039);
nor U15210 (N_15210,N_15199,N_15123);
nand U15211 (N_15211,N_15131,N_15029);
and U15212 (N_15212,N_15071,N_15081);
xor U15213 (N_15213,N_15173,N_15115);
and U15214 (N_15214,N_15132,N_15111);
nand U15215 (N_15215,N_15171,N_15080);
xor U15216 (N_15216,N_15107,N_15021);
nand U15217 (N_15217,N_15036,N_15058);
and U15218 (N_15218,N_15195,N_15129);
nand U15219 (N_15219,N_15117,N_15158);
and U15220 (N_15220,N_15082,N_15012);
xor U15221 (N_15221,N_15051,N_15143);
nor U15222 (N_15222,N_15042,N_15091);
xnor U15223 (N_15223,N_15053,N_15007);
nor U15224 (N_15224,N_15118,N_15162);
and U15225 (N_15225,N_15142,N_15032);
nand U15226 (N_15226,N_15175,N_15178);
or U15227 (N_15227,N_15038,N_15164);
and U15228 (N_15228,N_15031,N_15122);
nand U15229 (N_15229,N_15126,N_15169);
and U15230 (N_15230,N_15069,N_15119);
xnor U15231 (N_15231,N_15144,N_15019);
or U15232 (N_15232,N_15047,N_15015);
and U15233 (N_15233,N_15022,N_15088);
or U15234 (N_15234,N_15043,N_15141);
xnor U15235 (N_15235,N_15084,N_15137);
xnor U15236 (N_15236,N_15054,N_15060);
nand U15237 (N_15237,N_15074,N_15152);
or U15238 (N_15238,N_15189,N_15033);
and U15239 (N_15239,N_15011,N_15147);
nand U15240 (N_15240,N_15180,N_15159);
nor U15241 (N_15241,N_15188,N_15066);
or U15242 (N_15242,N_15055,N_15177);
xor U15243 (N_15243,N_15027,N_15110);
xnor U15244 (N_15244,N_15174,N_15016);
and U15245 (N_15245,N_15020,N_15090);
xnor U15246 (N_15246,N_15198,N_15150);
and U15247 (N_15247,N_15098,N_15050);
xor U15248 (N_15248,N_15017,N_15046);
and U15249 (N_15249,N_15006,N_15056);
nor U15250 (N_15250,N_15133,N_15155);
and U15251 (N_15251,N_15005,N_15170);
nor U15252 (N_15252,N_15166,N_15193);
nand U15253 (N_15253,N_15078,N_15135);
and U15254 (N_15254,N_15028,N_15105);
nand U15255 (N_15255,N_15037,N_15116);
nor U15256 (N_15256,N_15120,N_15181);
nand U15257 (N_15257,N_15153,N_15184);
nor U15258 (N_15258,N_15160,N_15094);
xnor U15259 (N_15259,N_15085,N_15089);
xor U15260 (N_15260,N_15083,N_15003);
nand U15261 (N_15261,N_15052,N_15059);
nand U15262 (N_15262,N_15067,N_15179);
and U15263 (N_15263,N_15099,N_15040);
nand U15264 (N_15264,N_15064,N_15148);
nor U15265 (N_15265,N_15086,N_15065);
and U15266 (N_15266,N_15063,N_15187);
and U15267 (N_15267,N_15048,N_15196);
and U15268 (N_15268,N_15096,N_15001);
xor U15269 (N_15269,N_15172,N_15041);
or U15270 (N_15270,N_15114,N_15100);
nand U15271 (N_15271,N_15124,N_15139);
and U15272 (N_15272,N_15194,N_15182);
xnor U15273 (N_15273,N_15026,N_15121);
xnor U15274 (N_15274,N_15034,N_15072);
nor U15275 (N_15275,N_15025,N_15024);
nor U15276 (N_15276,N_15014,N_15192);
xnor U15277 (N_15277,N_15004,N_15008);
and U15278 (N_15278,N_15068,N_15030);
xnor U15279 (N_15279,N_15087,N_15185);
xnor U15280 (N_15280,N_15061,N_15009);
nand U15281 (N_15281,N_15125,N_15103);
nand U15282 (N_15282,N_15093,N_15130);
or U15283 (N_15283,N_15101,N_15102);
nand U15284 (N_15284,N_15057,N_15138);
xnor U15285 (N_15285,N_15073,N_15167);
xnor U15286 (N_15286,N_15112,N_15070);
xnor U15287 (N_15287,N_15077,N_15176);
and U15288 (N_15288,N_15163,N_15092);
or U15289 (N_15289,N_15113,N_15154);
nor U15290 (N_15290,N_15140,N_15095);
xnor U15291 (N_15291,N_15010,N_15045);
and U15292 (N_15292,N_15191,N_15157);
and U15293 (N_15293,N_15075,N_15149);
xor U15294 (N_15294,N_15156,N_15062);
and U15295 (N_15295,N_15018,N_15013);
nor U15296 (N_15296,N_15151,N_15023);
and U15297 (N_15297,N_15104,N_15134);
xnor U15298 (N_15298,N_15197,N_15002);
or U15299 (N_15299,N_15049,N_15183);
xnor U15300 (N_15300,N_15040,N_15108);
and U15301 (N_15301,N_15028,N_15053);
nand U15302 (N_15302,N_15186,N_15181);
nand U15303 (N_15303,N_15194,N_15005);
and U15304 (N_15304,N_15021,N_15174);
or U15305 (N_15305,N_15127,N_15157);
xor U15306 (N_15306,N_15193,N_15029);
nor U15307 (N_15307,N_15093,N_15066);
xor U15308 (N_15308,N_15061,N_15141);
nor U15309 (N_15309,N_15022,N_15035);
and U15310 (N_15310,N_15193,N_15031);
xor U15311 (N_15311,N_15021,N_15061);
and U15312 (N_15312,N_15060,N_15123);
nand U15313 (N_15313,N_15172,N_15051);
and U15314 (N_15314,N_15154,N_15005);
or U15315 (N_15315,N_15029,N_15039);
xor U15316 (N_15316,N_15060,N_15129);
nor U15317 (N_15317,N_15045,N_15044);
nor U15318 (N_15318,N_15190,N_15041);
and U15319 (N_15319,N_15171,N_15026);
and U15320 (N_15320,N_15135,N_15013);
nand U15321 (N_15321,N_15073,N_15193);
and U15322 (N_15322,N_15168,N_15196);
or U15323 (N_15323,N_15102,N_15074);
nand U15324 (N_15324,N_15161,N_15064);
or U15325 (N_15325,N_15175,N_15187);
nor U15326 (N_15326,N_15180,N_15118);
xor U15327 (N_15327,N_15160,N_15121);
xnor U15328 (N_15328,N_15197,N_15017);
or U15329 (N_15329,N_15196,N_15082);
nor U15330 (N_15330,N_15157,N_15007);
or U15331 (N_15331,N_15145,N_15004);
xor U15332 (N_15332,N_15141,N_15182);
or U15333 (N_15333,N_15090,N_15091);
nand U15334 (N_15334,N_15171,N_15002);
or U15335 (N_15335,N_15172,N_15062);
and U15336 (N_15336,N_15154,N_15047);
and U15337 (N_15337,N_15049,N_15169);
or U15338 (N_15338,N_15173,N_15175);
and U15339 (N_15339,N_15031,N_15142);
nor U15340 (N_15340,N_15070,N_15041);
nor U15341 (N_15341,N_15170,N_15164);
xnor U15342 (N_15342,N_15174,N_15190);
or U15343 (N_15343,N_15188,N_15171);
xor U15344 (N_15344,N_15017,N_15008);
xnor U15345 (N_15345,N_15006,N_15176);
or U15346 (N_15346,N_15079,N_15069);
xor U15347 (N_15347,N_15174,N_15037);
nor U15348 (N_15348,N_15071,N_15152);
nor U15349 (N_15349,N_15024,N_15129);
and U15350 (N_15350,N_15015,N_15179);
and U15351 (N_15351,N_15020,N_15041);
nand U15352 (N_15352,N_15014,N_15129);
xnor U15353 (N_15353,N_15069,N_15151);
nand U15354 (N_15354,N_15086,N_15150);
nor U15355 (N_15355,N_15191,N_15178);
nand U15356 (N_15356,N_15021,N_15008);
xor U15357 (N_15357,N_15178,N_15129);
nand U15358 (N_15358,N_15148,N_15168);
and U15359 (N_15359,N_15159,N_15009);
or U15360 (N_15360,N_15013,N_15158);
xnor U15361 (N_15361,N_15067,N_15167);
xor U15362 (N_15362,N_15063,N_15073);
nand U15363 (N_15363,N_15162,N_15122);
nand U15364 (N_15364,N_15168,N_15188);
and U15365 (N_15365,N_15012,N_15151);
and U15366 (N_15366,N_15165,N_15170);
or U15367 (N_15367,N_15079,N_15121);
nor U15368 (N_15368,N_15137,N_15164);
xnor U15369 (N_15369,N_15140,N_15164);
nor U15370 (N_15370,N_15164,N_15003);
xor U15371 (N_15371,N_15010,N_15025);
or U15372 (N_15372,N_15070,N_15029);
or U15373 (N_15373,N_15067,N_15118);
xor U15374 (N_15374,N_15194,N_15031);
nand U15375 (N_15375,N_15089,N_15024);
nand U15376 (N_15376,N_15183,N_15001);
or U15377 (N_15377,N_15033,N_15072);
nor U15378 (N_15378,N_15055,N_15199);
or U15379 (N_15379,N_15181,N_15067);
nor U15380 (N_15380,N_15058,N_15063);
or U15381 (N_15381,N_15134,N_15173);
or U15382 (N_15382,N_15082,N_15199);
or U15383 (N_15383,N_15103,N_15113);
and U15384 (N_15384,N_15153,N_15019);
xnor U15385 (N_15385,N_15012,N_15103);
or U15386 (N_15386,N_15192,N_15039);
xnor U15387 (N_15387,N_15078,N_15055);
nor U15388 (N_15388,N_15133,N_15048);
nand U15389 (N_15389,N_15027,N_15091);
xnor U15390 (N_15390,N_15191,N_15087);
or U15391 (N_15391,N_15092,N_15191);
and U15392 (N_15392,N_15075,N_15067);
and U15393 (N_15393,N_15142,N_15088);
or U15394 (N_15394,N_15153,N_15180);
and U15395 (N_15395,N_15005,N_15138);
xor U15396 (N_15396,N_15076,N_15140);
nand U15397 (N_15397,N_15010,N_15012);
xor U15398 (N_15398,N_15185,N_15090);
or U15399 (N_15399,N_15145,N_15188);
or U15400 (N_15400,N_15223,N_15201);
nand U15401 (N_15401,N_15287,N_15346);
or U15402 (N_15402,N_15311,N_15353);
xnor U15403 (N_15403,N_15345,N_15277);
xnor U15404 (N_15404,N_15377,N_15384);
nand U15405 (N_15405,N_15338,N_15273);
and U15406 (N_15406,N_15249,N_15343);
nor U15407 (N_15407,N_15313,N_15212);
xnor U15408 (N_15408,N_15297,N_15284);
nand U15409 (N_15409,N_15381,N_15315);
and U15410 (N_15410,N_15302,N_15283);
and U15411 (N_15411,N_15375,N_15299);
and U15412 (N_15412,N_15348,N_15392);
xor U15413 (N_15413,N_15253,N_15232);
xor U15414 (N_15414,N_15324,N_15389);
nand U15415 (N_15415,N_15307,N_15390);
xnor U15416 (N_15416,N_15263,N_15241);
or U15417 (N_15417,N_15300,N_15340);
or U15418 (N_15418,N_15296,N_15228);
and U15419 (N_15419,N_15293,N_15396);
or U15420 (N_15420,N_15280,N_15366);
nand U15421 (N_15421,N_15398,N_15336);
or U15422 (N_15422,N_15252,N_15383);
nor U15423 (N_15423,N_15222,N_15248);
nand U15424 (N_15424,N_15327,N_15351);
nor U15425 (N_15425,N_15380,N_15225);
and U15426 (N_15426,N_15367,N_15231);
and U15427 (N_15427,N_15372,N_15285);
or U15428 (N_15428,N_15272,N_15339);
or U15429 (N_15429,N_15294,N_15274);
or U15430 (N_15430,N_15303,N_15275);
or U15431 (N_15431,N_15288,N_15255);
xnor U15432 (N_15432,N_15312,N_15266);
nand U15433 (N_15433,N_15226,N_15318);
xor U15434 (N_15434,N_15350,N_15230);
nor U15435 (N_15435,N_15358,N_15354);
nor U15436 (N_15436,N_15251,N_15238);
xor U15437 (N_15437,N_15298,N_15295);
xor U15438 (N_15438,N_15257,N_15363);
nand U15439 (N_15439,N_15268,N_15221);
and U15440 (N_15440,N_15322,N_15271);
or U15441 (N_15441,N_15216,N_15301);
or U15442 (N_15442,N_15364,N_15250);
nor U15443 (N_15443,N_15305,N_15229);
or U15444 (N_15444,N_15362,N_15369);
nand U15445 (N_15445,N_15335,N_15304);
xnor U15446 (N_15446,N_15206,N_15355);
nor U15447 (N_15447,N_15334,N_15244);
and U15448 (N_15448,N_15368,N_15376);
nand U15449 (N_15449,N_15349,N_15326);
nand U15450 (N_15450,N_15208,N_15330);
and U15451 (N_15451,N_15281,N_15373);
or U15452 (N_15452,N_15374,N_15388);
xnor U15453 (N_15453,N_15234,N_15314);
xor U15454 (N_15454,N_15309,N_15344);
nand U15455 (N_15455,N_15306,N_15397);
nor U15456 (N_15456,N_15323,N_15211);
nor U15457 (N_15457,N_15292,N_15245);
and U15458 (N_15458,N_15331,N_15360);
nand U15459 (N_15459,N_15240,N_15207);
or U15460 (N_15460,N_15329,N_15276);
or U15461 (N_15461,N_15317,N_15260);
and U15462 (N_15462,N_15218,N_15290);
nor U15463 (N_15463,N_15379,N_15254);
xnor U15464 (N_15464,N_15246,N_15264);
nand U15465 (N_15465,N_15205,N_15370);
nand U15466 (N_15466,N_15382,N_15356);
xnor U15467 (N_15467,N_15332,N_15333);
xnor U15468 (N_15468,N_15395,N_15261);
or U15469 (N_15469,N_15267,N_15239);
nand U15470 (N_15470,N_15394,N_15278);
nor U15471 (N_15471,N_15385,N_15219);
and U15472 (N_15472,N_15365,N_15308);
and U15473 (N_15473,N_15359,N_15224);
xnor U15474 (N_15474,N_15237,N_15204);
xor U15475 (N_15475,N_15227,N_15242);
nor U15476 (N_15476,N_15259,N_15291);
nand U15477 (N_15477,N_15282,N_15347);
nand U15478 (N_15478,N_15203,N_15217);
or U15479 (N_15479,N_15391,N_15399);
nand U15480 (N_15480,N_15341,N_15378);
nor U15481 (N_15481,N_15200,N_15202);
xnor U15482 (N_15482,N_15321,N_15220);
nor U15483 (N_15483,N_15265,N_15215);
or U15484 (N_15484,N_15352,N_15279);
nand U15485 (N_15485,N_15342,N_15337);
nand U15486 (N_15486,N_15270,N_15316);
or U15487 (N_15487,N_15236,N_15310);
and U15488 (N_15488,N_15357,N_15289);
or U15489 (N_15489,N_15233,N_15243);
or U15490 (N_15490,N_15210,N_15214);
nand U15491 (N_15491,N_15262,N_15286);
and U15492 (N_15492,N_15269,N_15256);
xor U15493 (N_15493,N_15209,N_15361);
and U15494 (N_15494,N_15320,N_15393);
nand U15495 (N_15495,N_15213,N_15325);
or U15496 (N_15496,N_15386,N_15258);
and U15497 (N_15497,N_15387,N_15235);
nor U15498 (N_15498,N_15371,N_15319);
nand U15499 (N_15499,N_15328,N_15247);
xor U15500 (N_15500,N_15382,N_15203);
nand U15501 (N_15501,N_15255,N_15383);
and U15502 (N_15502,N_15389,N_15257);
nor U15503 (N_15503,N_15382,N_15292);
xnor U15504 (N_15504,N_15244,N_15267);
xor U15505 (N_15505,N_15376,N_15234);
xor U15506 (N_15506,N_15291,N_15233);
nor U15507 (N_15507,N_15284,N_15356);
nor U15508 (N_15508,N_15252,N_15289);
nand U15509 (N_15509,N_15200,N_15395);
and U15510 (N_15510,N_15329,N_15259);
xnor U15511 (N_15511,N_15386,N_15332);
and U15512 (N_15512,N_15208,N_15379);
xor U15513 (N_15513,N_15268,N_15312);
and U15514 (N_15514,N_15326,N_15366);
and U15515 (N_15515,N_15220,N_15361);
or U15516 (N_15516,N_15223,N_15224);
and U15517 (N_15517,N_15277,N_15237);
nand U15518 (N_15518,N_15304,N_15217);
or U15519 (N_15519,N_15284,N_15347);
xnor U15520 (N_15520,N_15388,N_15264);
and U15521 (N_15521,N_15313,N_15390);
xor U15522 (N_15522,N_15265,N_15303);
nor U15523 (N_15523,N_15381,N_15324);
xnor U15524 (N_15524,N_15396,N_15383);
xor U15525 (N_15525,N_15306,N_15280);
nand U15526 (N_15526,N_15372,N_15312);
nor U15527 (N_15527,N_15273,N_15254);
or U15528 (N_15528,N_15394,N_15248);
xor U15529 (N_15529,N_15229,N_15318);
nor U15530 (N_15530,N_15381,N_15389);
and U15531 (N_15531,N_15233,N_15266);
nor U15532 (N_15532,N_15294,N_15367);
and U15533 (N_15533,N_15257,N_15333);
or U15534 (N_15534,N_15270,N_15207);
nand U15535 (N_15535,N_15391,N_15278);
nor U15536 (N_15536,N_15320,N_15218);
nand U15537 (N_15537,N_15306,N_15240);
nor U15538 (N_15538,N_15378,N_15250);
nor U15539 (N_15539,N_15213,N_15241);
or U15540 (N_15540,N_15339,N_15252);
nor U15541 (N_15541,N_15227,N_15351);
and U15542 (N_15542,N_15207,N_15310);
and U15543 (N_15543,N_15367,N_15241);
or U15544 (N_15544,N_15279,N_15280);
or U15545 (N_15545,N_15310,N_15353);
xnor U15546 (N_15546,N_15329,N_15272);
nor U15547 (N_15547,N_15236,N_15309);
or U15548 (N_15548,N_15378,N_15330);
nor U15549 (N_15549,N_15321,N_15277);
and U15550 (N_15550,N_15275,N_15254);
and U15551 (N_15551,N_15238,N_15285);
nor U15552 (N_15552,N_15223,N_15297);
nand U15553 (N_15553,N_15214,N_15220);
or U15554 (N_15554,N_15245,N_15325);
xor U15555 (N_15555,N_15202,N_15258);
nand U15556 (N_15556,N_15325,N_15308);
xnor U15557 (N_15557,N_15316,N_15368);
or U15558 (N_15558,N_15357,N_15378);
nand U15559 (N_15559,N_15255,N_15214);
xnor U15560 (N_15560,N_15362,N_15326);
nor U15561 (N_15561,N_15285,N_15346);
nor U15562 (N_15562,N_15265,N_15223);
or U15563 (N_15563,N_15382,N_15208);
xnor U15564 (N_15564,N_15270,N_15352);
nor U15565 (N_15565,N_15307,N_15335);
and U15566 (N_15566,N_15308,N_15204);
and U15567 (N_15567,N_15366,N_15224);
and U15568 (N_15568,N_15287,N_15367);
and U15569 (N_15569,N_15304,N_15328);
or U15570 (N_15570,N_15382,N_15273);
or U15571 (N_15571,N_15297,N_15374);
nor U15572 (N_15572,N_15366,N_15259);
xor U15573 (N_15573,N_15365,N_15220);
and U15574 (N_15574,N_15387,N_15247);
and U15575 (N_15575,N_15365,N_15271);
xor U15576 (N_15576,N_15215,N_15345);
nand U15577 (N_15577,N_15396,N_15367);
nor U15578 (N_15578,N_15332,N_15225);
nor U15579 (N_15579,N_15308,N_15338);
xor U15580 (N_15580,N_15377,N_15356);
xor U15581 (N_15581,N_15329,N_15253);
nand U15582 (N_15582,N_15267,N_15302);
and U15583 (N_15583,N_15211,N_15302);
xnor U15584 (N_15584,N_15381,N_15348);
nor U15585 (N_15585,N_15259,N_15370);
nor U15586 (N_15586,N_15256,N_15386);
and U15587 (N_15587,N_15386,N_15246);
and U15588 (N_15588,N_15238,N_15232);
nand U15589 (N_15589,N_15222,N_15230);
and U15590 (N_15590,N_15247,N_15306);
or U15591 (N_15591,N_15284,N_15331);
or U15592 (N_15592,N_15319,N_15350);
and U15593 (N_15593,N_15390,N_15392);
and U15594 (N_15594,N_15251,N_15211);
nand U15595 (N_15595,N_15377,N_15218);
xor U15596 (N_15596,N_15315,N_15241);
xor U15597 (N_15597,N_15369,N_15381);
nand U15598 (N_15598,N_15341,N_15314);
nand U15599 (N_15599,N_15394,N_15333);
nand U15600 (N_15600,N_15516,N_15498);
xor U15601 (N_15601,N_15438,N_15435);
or U15602 (N_15602,N_15460,N_15479);
nor U15603 (N_15603,N_15509,N_15573);
or U15604 (N_15604,N_15547,N_15536);
nand U15605 (N_15605,N_15402,N_15477);
xnor U15606 (N_15606,N_15462,N_15428);
xnor U15607 (N_15607,N_15565,N_15576);
nand U15608 (N_15608,N_15440,N_15587);
nor U15609 (N_15609,N_15458,N_15415);
and U15610 (N_15610,N_15468,N_15599);
or U15611 (N_15611,N_15544,N_15420);
nor U15612 (N_15612,N_15452,N_15581);
or U15613 (N_15613,N_15523,N_15430);
and U15614 (N_15614,N_15524,N_15489);
nand U15615 (N_15615,N_15531,N_15474);
and U15616 (N_15616,N_15476,N_15480);
xor U15617 (N_15617,N_15589,N_15448);
nand U15618 (N_15618,N_15541,N_15493);
nand U15619 (N_15619,N_15583,N_15443);
xor U15620 (N_15620,N_15478,N_15575);
xor U15621 (N_15621,N_15567,N_15537);
nand U15622 (N_15622,N_15511,N_15557);
and U15623 (N_15623,N_15491,N_15554);
or U15624 (N_15624,N_15564,N_15595);
xor U15625 (N_15625,N_15426,N_15513);
or U15626 (N_15626,N_15505,N_15504);
nor U15627 (N_15627,N_15475,N_15563);
xnor U15628 (N_15628,N_15441,N_15529);
xor U15629 (N_15629,N_15558,N_15465);
nor U15630 (N_15630,N_15409,N_15432);
or U15631 (N_15631,N_15562,N_15507);
and U15632 (N_15632,N_15407,N_15429);
xor U15633 (N_15633,N_15455,N_15467);
nor U15634 (N_15634,N_15483,N_15528);
xor U15635 (N_15635,N_15423,N_15419);
or U15636 (N_15636,N_15470,N_15431);
and U15637 (N_15637,N_15539,N_15450);
and U15638 (N_15638,N_15406,N_15457);
nand U15639 (N_15639,N_15514,N_15540);
nor U15640 (N_15640,N_15456,N_15579);
nand U15641 (N_15641,N_15515,N_15453);
xnor U15642 (N_15642,N_15552,N_15550);
xor U15643 (N_15643,N_15488,N_15592);
nand U15644 (N_15644,N_15466,N_15593);
and U15645 (N_15645,N_15520,N_15538);
or U15646 (N_15646,N_15532,N_15427);
xnor U15647 (N_15647,N_15444,N_15588);
xnor U15648 (N_15648,N_15495,N_15416);
and U15649 (N_15649,N_15425,N_15445);
nand U15650 (N_15650,N_15551,N_15446);
and U15651 (N_15651,N_15424,N_15501);
and U15652 (N_15652,N_15598,N_15586);
nand U15653 (N_15653,N_15522,N_15512);
nor U15654 (N_15654,N_15451,N_15405);
nor U15655 (N_15655,N_15421,N_15545);
nor U15656 (N_15656,N_15559,N_15482);
xor U15657 (N_15657,N_15418,N_15502);
nor U15658 (N_15658,N_15526,N_15543);
or U15659 (N_15659,N_15571,N_15459);
nand U15660 (N_15660,N_15481,N_15473);
nor U15661 (N_15661,N_15411,N_15553);
xnor U15662 (N_15662,N_15584,N_15401);
and U15663 (N_15663,N_15591,N_15503);
or U15664 (N_15664,N_15410,N_15590);
nor U15665 (N_15665,N_15580,N_15497);
nand U15666 (N_15666,N_15408,N_15561);
or U15667 (N_15667,N_15454,N_15496);
nor U15668 (N_15668,N_15484,N_15414);
xor U15669 (N_15669,N_15578,N_15490);
nand U15670 (N_15670,N_15548,N_15560);
nor U15671 (N_15671,N_15403,N_15471);
nor U15672 (N_15672,N_15527,N_15597);
nand U15673 (N_15673,N_15542,N_15525);
and U15674 (N_15674,N_15499,N_15422);
and U15675 (N_15675,N_15517,N_15472);
nand U15676 (N_15676,N_15506,N_15500);
and U15677 (N_15677,N_15461,N_15485);
nand U15678 (N_15678,N_15530,N_15447);
nand U15679 (N_15679,N_15568,N_15510);
nor U15680 (N_15680,N_15464,N_15596);
nand U15681 (N_15681,N_15439,N_15549);
nand U15682 (N_15682,N_15492,N_15486);
nor U15683 (N_15683,N_15463,N_15582);
nand U15684 (N_15684,N_15469,N_15572);
nor U15685 (N_15685,N_15494,N_15555);
nand U15686 (N_15686,N_15487,N_15518);
or U15687 (N_15687,N_15508,N_15437);
or U15688 (N_15688,N_15519,N_15569);
nand U15689 (N_15689,N_15413,N_15556);
xnor U15690 (N_15690,N_15546,N_15449);
and U15691 (N_15691,N_15574,N_15570);
and U15692 (N_15692,N_15404,N_15417);
nand U15693 (N_15693,N_15436,N_15594);
xnor U15694 (N_15694,N_15412,N_15585);
or U15695 (N_15695,N_15566,N_15433);
nor U15696 (N_15696,N_15442,N_15577);
or U15697 (N_15697,N_15534,N_15533);
xnor U15698 (N_15698,N_15434,N_15400);
nor U15699 (N_15699,N_15521,N_15535);
and U15700 (N_15700,N_15516,N_15563);
nor U15701 (N_15701,N_15584,N_15576);
xor U15702 (N_15702,N_15590,N_15538);
nor U15703 (N_15703,N_15507,N_15424);
nor U15704 (N_15704,N_15510,N_15539);
xnor U15705 (N_15705,N_15445,N_15430);
nor U15706 (N_15706,N_15545,N_15475);
nor U15707 (N_15707,N_15593,N_15589);
xnor U15708 (N_15708,N_15449,N_15555);
nand U15709 (N_15709,N_15539,N_15560);
or U15710 (N_15710,N_15481,N_15599);
xor U15711 (N_15711,N_15530,N_15437);
nor U15712 (N_15712,N_15456,N_15429);
nand U15713 (N_15713,N_15425,N_15593);
or U15714 (N_15714,N_15583,N_15501);
and U15715 (N_15715,N_15545,N_15461);
nand U15716 (N_15716,N_15415,N_15467);
nor U15717 (N_15717,N_15489,N_15558);
nand U15718 (N_15718,N_15508,N_15472);
and U15719 (N_15719,N_15555,N_15568);
or U15720 (N_15720,N_15421,N_15576);
nor U15721 (N_15721,N_15457,N_15525);
nand U15722 (N_15722,N_15545,N_15409);
or U15723 (N_15723,N_15489,N_15497);
and U15724 (N_15724,N_15582,N_15507);
nor U15725 (N_15725,N_15561,N_15551);
or U15726 (N_15726,N_15482,N_15470);
or U15727 (N_15727,N_15526,N_15444);
or U15728 (N_15728,N_15481,N_15562);
nand U15729 (N_15729,N_15536,N_15474);
nor U15730 (N_15730,N_15420,N_15547);
xor U15731 (N_15731,N_15475,N_15550);
nand U15732 (N_15732,N_15479,N_15583);
nand U15733 (N_15733,N_15432,N_15478);
xor U15734 (N_15734,N_15414,N_15581);
or U15735 (N_15735,N_15544,N_15585);
nor U15736 (N_15736,N_15490,N_15401);
or U15737 (N_15737,N_15597,N_15528);
or U15738 (N_15738,N_15504,N_15450);
xnor U15739 (N_15739,N_15498,N_15433);
xnor U15740 (N_15740,N_15595,N_15402);
and U15741 (N_15741,N_15524,N_15419);
nor U15742 (N_15742,N_15552,N_15526);
and U15743 (N_15743,N_15566,N_15546);
and U15744 (N_15744,N_15587,N_15551);
nor U15745 (N_15745,N_15438,N_15543);
or U15746 (N_15746,N_15422,N_15411);
nand U15747 (N_15747,N_15505,N_15521);
nand U15748 (N_15748,N_15440,N_15426);
or U15749 (N_15749,N_15549,N_15567);
nand U15750 (N_15750,N_15596,N_15581);
or U15751 (N_15751,N_15485,N_15556);
or U15752 (N_15752,N_15481,N_15569);
nor U15753 (N_15753,N_15434,N_15475);
and U15754 (N_15754,N_15521,N_15448);
nor U15755 (N_15755,N_15419,N_15530);
nor U15756 (N_15756,N_15418,N_15524);
and U15757 (N_15757,N_15457,N_15577);
or U15758 (N_15758,N_15488,N_15554);
or U15759 (N_15759,N_15499,N_15401);
nand U15760 (N_15760,N_15562,N_15414);
or U15761 (N_15761,N_15487,N_15590);
or U15762 (N_15762,N_15447,N_15439);
or U15763 (N_15763,N_15503,N_15401);
nor U15764 (N_15764,N_15463,N_15584);
nor U15765 (N_15765,N_15547,N_15518);
nand U15766 (N_15766,N_15529,N_15481);
nor U15767 (N_15767,N_15518,N_15457);
nand U15768 (N_15768,N_15468,N_15416);
nor U15769 (N_15769,N_15432,N_15521);
and U15770 (N_15770,N_15579,N_15557);
or U15771 (N_15771,N_15563,N_15450);
and U15772 (N_15772,N_15417,N_15435);
or U15773 (N_15773,N_15529,N_15588);
or U15774 (N_15774,N_15544,N_15550);
or U15775 (N_15775,N_15483,N_15515);
and U15776 (N_15776,N_15559,N_15553);
nand U15777 (N_15777,N_15449,N_15541);
xnor U15778 (N_15778,N_15430,N_15415);
nand U15779 (N_15779,N_15572,N_15436);
and U15780 (N_15780,N_15498,N_15442);
and U15781 (N_15781,N_15512,N_15500);
xnor U15782 (N_15782,N_15425,N_15437);
and U15783 (N_15783,N_15449,N_15450);
xor U15784 (N_15784,N_15458,N_15581);
or U15785 (N_15785,N_15429,N_15428);
xnor U15786 (N_15786,N_15580,N_15574);
xor U15787 (N_15787,N_15477,N_15518);
nor U15788 (N_15788,N_15452,N_15471);
and U15789 (N_15789,N_15597,N_15495);
and U15790 (N_15790,N_15470,N_15568);
xor U15791 (N_15791,N_15417,N_15518);
xor U15792 (N_15792,N_15414,N_15534);
xnor U15793 (N_15793,N_15421,N_15475);
or U15794 (N_15794,N_15553,N_15474);
and U15795 (N_15795,N_15497,N_15453);
nor U15796 (N_15796,N_15446,N_15481);
and U15797 (N_15797,N_15578,N_15465);
nor U15798 (N_15798,N_15502,N_15412);
or U15799 (N_15799,N_15456,N_15590);
xnor U15800 (N_15800,N_15723,N_15751);
nor U15801 (N_15801,N_15617,N_15687);
and U15802 (N_15802,N_15729,N_15636);
nand U15803 (N_15803,N_15733,N_15655);
nand U15804 (N_15804,N_15743,N_15613);
xor U15805 (N_15805,N_15667,N_15782);
xnor U15806 (N_15806,N_15759,N_15600);
or U15807 (N_15807,N_15770,N_15649);
or U15808 (N_15808,N_15766,N_15702);
and U15809 (N_15809,N_15719,N_15607);
nor U15810 (N_15810,N_15640,N_15626);
nor U15811 (N_15811,N_15608,N_15638);
nor U15812 (N_15812,N_15749,N_15740);
nand U15813 (N_15813,N_15665,N_15648);
or U15814 (N_15814,N_15634,N_15788);
or U15815 (N_15815,N_15656,N_15601);
or U15816 (N_15816,N_15642,N_15658);
and U15817 (N_15817,N_15605,N_15778);
and U15818 (N_15818,N_15795,N_15761);
and U15819 (N_15819,N_15675,N_15669);
or U15820 (N_15820,N_15639,N_15706);
nand U15821 (N_15821,N_15701,N_15700);
and U15822 (N_15822,N_15690,N_15726);
and U15823 (N_15823,N_15753,N_15609);
nor U15824 (N_15824,N_15629,N_15791);
xor U15825 (N_15825,N_15750,N_15731);
or U15826 (N_15826,N_15610,N_15628);
or U15827 (N_15827,N_15627,N_15757);
or U15828 (N_15828,N_15620,N_15670);
xor U15829 (N_15829,N_15727,N_15752);
and U15830 (N_15830,N_15790,N_15739);
nor U15831 (N_15831,N_15737,N_15654);
nor U15832 (N_15832,N_15754,N_15748);
nor U15833 (N_15833,N_15738,N_15683);
xnor U15834 (N_15834,N_15728,N_15619);
nand U15835 (N_15835,N_15714,N_15674);
and U15836 (N_15836,N_15779,N_15784);
xnor U15837 (N_15837,N_15664,N_15744);
or U15838 (N_15838,N_15780,N_15708);
nor U15839 (N_15839,N_15765,N_15732);
xor U15840 (N_15840,N_15792,N_15688);
nor U15841 (N_15841,N_15705,N_15604);
xnor U15842 (N_15842,N_15709,N_15786);
or U15843 (N_15843,N_15773,N_15746);
and U15844 (N_15844,N_15696,N_15735);
or U15845 (N_15845,N_15734,N_15794);
and U15846 (N_15846,N_15633,N_15760);
and U15847 (N_15847,N_15685,N_15614);
nand U15848 (N_15848,N_15755,N_15684);
or U15849 (N_15849,N_15637,N_15769);
and U15850 (N_15850,N_15793,N_15711);
xnor U15851 (N_15851,N_15603,N_15776);
or U15852 (N_15852,N_15623,N_15615);
or U15853 (N_15853,N_15771,N_15797);
nand U15854 (N_15854,N_15673,N_15643);
xnor U15855 (N_15855,N_15611,N_15678);
nor U15856 (N_15856,N_15736,N_15622);
or U15857 (N_15857,N_15682,N_15710);
nor U15858 (N_15858,N_15653,N_15718);
or U15859 (N_15859,N_15606,N_15630);
nand U15860 (N_15860,N_15689,N_15713);
xnor U15861 (N_15861,N_15679,N_15796);
xor U15862 (N_15862,N_15712,N_15652);
or U15863 (N_15863,N_15695,N_15767);
xor U15864 (N_15864,N_15798,N_15616);
xor U15865 (N_15865,N_15745,N_15602);
or U15866 (N_15866,N_15661,N_15676);
nor U15867 (N_15867,N_15768,N_15624);
and U15868 (N_15868,N_15730,N_15707);
nor U15869 (N_15869,N_15686,N_15666);
nand U15870 (N_15870,N_15677,N_15758);
and U15871 (N_15871,N_15672,N_15742);
xor U15872 (N_15872,N_15631,N_15644);
and U15873 (N_15873,N_15618,N_15646);
nor U15874 (N_15874,N_15612,N_15625);
nand U15875 (N_15875,N_15651,N_15785);
nand U15876 (N_15876,N_15699,N_15663);
xnor U15877 (N_15877,N_15645,N_15756);
nor U15878 (N_15878,N_15647,N_15775);
nor U15879 (N_15879,N_15722,N_15635);
xnor U15880 (N_15880,N_15741,N_15662);
nor U15881 (N_15881,N_15660,N_15783);
and U15882 (N_15882,N_15697,N_15692);
nor U15883 (N_15883,N_15659,N_15703);
nor U15884 (N_15884,N_15680,N_15787);
xor U15885 (N_15885,N_15720,N_15799);
nand U15886 (N_15886,N_15657,N_15693);
nor U15887 (N_15887,N_15641,N_15781);
nand U15888 (N_15888,N_15694,N_15621);
nand U15889 (N_15889,N_15671,N_15762);
or U15890 (N_15890,N_15717,N_15704);
xor U15891 (N_15891,N_15789,N_15650);
nand U15892 (N_15892,N_15668,N_15691);
and U15893 (N_15893,N_15698,N_15725);
xor U15894 (N_15894,N_15774,N_15777);
nor U15895 (N_15895,N_15724,N_15716);
nor U15896 (N_15896,N_15747,N_15721);
or U15897 (N_15897,N_15632,N_15772);
or U15898 (N_15898,N_15763,N_15681);
nor U15899 (N_15899,N_15715,N_15764);
xnor U15900 (N_15900,N_15684,N_15795);
nor U15901 (N_15901,N_15795,N_15724);
nor U15902 (N_15902,N_15779,N_15679);
nor U15903 (N_15903,N_15770,N_15646);
nor U15904 (N_15904,N_15620,N_15791);
nand U15905 (N_15905,N_15759,N_15613);
or U15906 (N_15906,N_15766,N_15799);
or U15907 (N_15907,N_15721,N_15623);
nor U15908 (N_15908,N_15704,N_15655);
or U15909 (N_15909,N_15612,N_15606);
nand U15910 (N_15910,N_15644,N_15606);
nor U15911 (N_15911,N_15703,N_15704);
nand U15912 (N_15912,N_15659,N_15773);
or U15913 (N_15913,N_15677,N_15630);
nand U15914 (N_15914,N_15630,N_15696);
or U15915 (N_15915,N_15659,N_15709);
xnor U15916 (N_15916,N_15601,N_15787);
and U15917 (N_15917,N_15649,N_15768);
or U15918 (N_15918,N_15737,N_15607);
and U15919 (N_15919,N_15730,N_15724);
nor U15920 (N_15920,N_15712,N_15644);
and U15921 (N_15921,N_15654,N_15775);
and U15922 (N_15922,N_15798,N_15653);
nor U15923 (N_15923,N_15681,N_15687);
or U15924 (N_15924,N_15620,N_15771);
or U15925 (N_15925,N_15771,N_15734);
nor U15926 (N_15926,N_15606,N_15731);
nor U15927 (N_15927,N_15717,N_15644);
or U15928 (N_15928,N_15624,N_15735);
and U15929 (N_15929,N_15728,N_15719);
xnor U15930 (N_15930,N_15793,N_15751);
and U15931 (N_15931,N_15771,N_15695);
and U15932 (N_15932,N_15664,N_15616);
xnor U15933 (N_15933,N_15723,N_15715);
and U15934 (N_15934,N_15720,N_15674);
or U15935 (N_15935,N_15616,N_15649);
nand U15936 (N_15936,N_15744,N_15718);
nor U15937 (N_15937,N_15683,N_15741);
or U15938 (N_15938,N_15618,N_15611);
nor U15939 (N_15939,N_15798,N_15737);
xor U15940 (N_15940,N_15790,N_15636);
xor U15941 (N_15941,N_15784,N_15623);
or U15942 (N_15942,N_15734,N_15743);
and U15943 (N_15943,N_15612,N_15757);
and U15944 (N_15944,N_15694,N_15692);
xor U15945 (N_15945,N_15746,N_15726);
or U15946 (N_15946,N_15718,N_15763);
or U15947 (N_15947,N_15612,N_15602);
nor U15948 (N_15948,N_15719,N_15735);
xor U15949 (N_15949,N_15680,N_15602);
nand U15950 (N_15950,N_15742,N_15628);
and U15951 (N_15951,N_15606,N_15627);
nor U15952 (N_15952,N_15665,N_15689);
and U15953 (N_15953,N_15678,N_15764);
nor U15954 (N_15954,N_15733,N_15612);
nand U15955 (N_15955,N_15714,N_15759);
nand U15956 (N_15956,N_15746,N_15775);
and U15957 (N_15957,N_15799,N_15697);
or U15958 (N_15958,N_15793,N_15647);
nand U15959 (N_15959,N_15672,N_15712);
nor U15960 (N_15960,N_15651,N_15661);
xnor U15961 (N_15961,N_15668,N_15657);
nor U15962 (N_15962,N_15789,N_15780);
nand U15963 (N_15963,N_15710,N_15642);
nand U15964 (N_15964,N_15690,N_15724);
nor U15965 (N_15965,N_15723,N_15780);
nand U15966 (N_15966,N_15738,N_15669);
or U15967 (N_15967,N_15753,N_15798);
or U15968 (N_15968,N_15750,N_15707);
and U15969 (N_15969,N_15771,N_15609);
nand U15970 (N_15970,N_15703,N_15694);
nor U15971 (N_15971,N_15780,N_15674);
and U15972 (N_15972,N_15752,N_15780);
xor U15973 (N_15973,N_15754,N_15723);
nand U15974 (N_15974,N_15649,N_15648);
nand U15975 (N_15975,N_15790,N_15737);
nor U15976 (N_15976,N_15690,N_15774);
or U15977 (N_15977,N_15766,N_15705);
and U15978 (N_15978,N_15704,N_15665);
or U15979 (N_15979,N_15785,N_15615);
nor U15980 (N_15980,N_15639,N_15606);
nand U15981 (N_15981,N_15702,N_15763);
and U15982 (N_15982,N_15713,N_15612);
or U15983 (N_15983,N_15759,N_15797);
or U15984 (N_15984,N_15781,N_15700);
and U15985 (N_15985,N_15769,N_15666);
or U15986 (N_15986,N_15684,N_15679);
nor U15987 (N_15987,N_15727,N_15631);
nor U15988 (N_15988,N_15698,N_15792);
or U15989 (N_15989,N_15718,N_15645);
and U15990 (N_15990,N_15761,N_15669);
or U15991 (N_15991,N_15753,N_15658);
or U15992 (N_15992,N_15789,N_15692);
or U15993 (N_15993,N_15752,N_15732);
nand U15994 (N_15994,N_15638,N_15698);
nand U15995 (N_15995,N_15648,N_15702);
or U15996 (N_15996,N_15642,N_15774);
nor U15997 (N_15997,N_15659,N_15603);
nand U15998 (N_15998,N_15768,N_15746);
nand U15999 (N_15999,N_15715,N_15667);
xor U16000 (N_16000,N_15856,N_15972);
nand U16001 (N_16001,N_15868,N_15839);
nand U16002 (N_16002,N_15887,N_15941);
xor U16003 (N_16003,N_15876,N_15869);
and U16004 (N_16004,N_15872,N_15873);
xor U16005 (N_16005,N_15926,N_15965);
nor U16006 (N_16006,N_15935,N_15999);
nand U16007 (N_16007,N_15843,N_15893);
nand U16008 (N_16008,N_15950,N_15900);
nand U16009 (N_16009,N_15801,N_15924);
nor U16010 (N_16010,N_15824,N_15975);
or U16011 (N_16011,N_15855,N_15960);
nand U16012 (N_16012,N_15894,N_15979);
nor U16013 (N_16013,N_15936,N_15806);
xor U16014 (N_16014,N_15823,N_15804);
or U16015 (N_16015,N_15827,N_15838);
xor U16016 (N_16016,N_15857,N_15957);
xnor U16017 (N_16017,N_15969,N_15939);
and U16018 (N_16018,N_15962,N_15896);
or U16019 (N_16019,N_15910,N_15877);
and U16020 (N_16020,N_15889,N_15967);
xnor U16021 (N_16021,N_15891,N_15840);
nand U16022 (N_16022,N_15912,N_15892);
and U16023 (N_16023,N_15860,N_15819);
nand U16024 (N_16024,N_15955,N_15833);
nand U16025 (N_16025,N_15992,N_15805);
nand U16026 (N_16026,N_15818,N_15940);
or U16027 (N_16027,N_15928,N_15997);
nor U16028 (N_16028,N_15832,N_15858);
and U16029 (N_16029,N_15919,N_15879);
nor U16030 (N_16030,N_15987,N_15983);
nor U16031 (N_16031,N_15849,N_15809);
xor U16032 (N_16032,N_15985,N_15874);
nand U16033 (N_16033,N_15851,N_15841);
nand U16034 (N_16034,N_15852,N_15954);
nor U16035 (N_16035,N_15817,N_15977);
nand U16036 (N_16036,N_15995,N_15808);
xnor U16037 (N_16037,N_15811,N_15971);
nor U16038 (N_16038,N_15885,N_15844);
or U16039 (N_16039,N_15883,N_15929);
and U16040 (N_16040,N_15937,N_15813);
xnor U16041 (N_16041,N_15945,N_15864);
nand U16042 (N_16042,N_15904,N_15836);
nor U16043 (N_16043,N_15907,N_15800);
or U16044 (N_16044,N_15964,N_15895);
and U16045 (N_16045,N_15993,N_15988);
and U16046 (N_16046,N_15916,N_15932);
nor U16047 (N_16047,N_15989,N_15944);
or U16048 (N_16048,N_15853,N_15897);
or U16049 (N_16049,N_15807,N_15842);
or U16050 (N_16050,N_15922,N_15903);
nor U16051 (N_16051,N_15847,N_15854);
nor U16052 (N_16052,N_15942,N_15834);
nor U16053 (N_16053,N_15923,N_15915);
nor U16054 (N_16054,N_15933,N_15970);
and U16055 (N_16055,N_15990,N_15850);
nand U16056 (N_16056,N_15810,N_15870);
or U16057 (N_16057,N_15973,N_15996);
xor U16058 (N_16058,N_15948,N_15921);
nand U16059 (N_16059,N_15902,N_15927);
xnor U16060 (N_16060,N_15835,N_15898);
and U16061 (N_16061,N_15884,N_15946);
nor U16062 (N_16062,N_15815,N_15875);
xor U16063 (N_16063,N_15865,N_15830);
nand U16064 (N_16064,N_15866,N_15822);
xnor U16065 (N_16065,N_15963,N_15871);
xnor U16066 (N_16066,N_15998,N_15953);
and U16067 (N_16067,N_15821,N_15982);
nand U16068 (N_16068,N_15931,N_15981);
nand U16069 (N_16069,N_15816,N_15909);
nor U16070 (N_16070,N_15930,N_15829);
nand U16071 (N_16071,N_15846,N_15925);
nor U16072 (N_16072,N_15952,N_15863);
or U16073 (N_16073,N_15826,N_15888);
xor U16074 (N_16074,N_15867,N_15917);
xnor U16075 (N_16075,N_15901,N_15938);
and U16076 (N_16076,N_15980,N_15802);
and U16077 (N_16077,N_15947,N_15880);
nand U16078 (N_16078,N_15913,N_15920);
or U16079 (N_16079,N_15994,N_15848);
nor U16080 (N_16080,N_15978,N_15803);
nand U16081 (N_16081,N_15845,N_15984);
nor U16082 (N_16082,N_15914,N_15828);
and U16083 (N_16083,N_15820,N_15991);
and U16084 (N_16084,N_15934,N_15958);
and U16085 (N_16085,N_15886,N_15890);
nor U16086 (N_16086,N_15831,N_15951);
xor U16087 (N_16087,N_15814,N_15905);
nand U16088 (N_16088,N_15899,N_15918);
and U16089 (N_16089,N_15906,N_15949);
or U16090 (N_16090,N_15956,N_15976);
and U16091 (N_16091,N_15961,N_15968);
or U16092 (N_16092,N_15837,N_15878);
or U16093 (N_16093,N_15974,N_15862);
or U16094 (N_16094,N_15825,N_15861);
nand U16095 (N_16095,N_15812,N_15908);
and U16096 (N_16096,N_15859,N_15911);
xor U16097 (N_16097,N_15966,N_15881);
nand U16098 (N_16098,N_15959,N_15882);
xnor U16099 (N_16099,N_15986,N_15943);
or U16100 (N_16100,N_15804,N_15969);
nand U16101 (N_16101,N_15884,N_15987);
nand U16102 (N_16102,N_15969,N_15849);
nor U16103 (N_16103,N_15867,N_15877);
or U16104 (N_16104,N_15948,N_15930);
or U16105 (N_16105,N_15947,N_15803);
or U16106 (N_16106,N_15991,N_15847);
and U16107 (N_16107,N_15960,N_15806);
nand U16108 (N_16108,N_15859,N_15890);
or U16109 (N_16109,N_15929,N_15957);
and U16110 (N_16110,N_15909,N_15972);
or U16111 (N_16111,N_15992,N_15928);
and U16112 (N_16112,N_15915,N_15937);
nand U16113 (N_16113,N_15836,N_15968);
and U16114 (N_16114,N_15937,N_15908);
or U16115 (N_16115,N_15870,N_15942);
nand U16116 (N_16116,N_15826,N_15887);
or U16117 (N_16117,N_15903,N_15952);
xnor U16118 (N_16118,N_15941,N_15811);
nand U16119 (N_16119,N_15850,N_15903);
xor U16120 (N_16120,N_15864,N_15874);
nor U16121 (N_16121,N_15934,N_15868);
xor U16122 (N_16122,N_15952,N_15940);
and U16123 (N_16123,N_15961,N_15848);
nor U16124 (N_16124,N_15884,N_15992);
and U16125 (N_16125,N_15993,N_15840);
nor U16126 (N_16126,N_15800,N_15943);
and U16127 (N_16127,N_15871,N_15804);
xor U16128 (N_16128,N_15961,N_15870);
nor U16129 (N_16129,N_15903,N_15877);
xnor U16130 (N_16130,N_15852,N_15986);
or U16131 (N_16131,N_15813,N_15999);
xor U16132 (N_16132,N_15868,N_15955);
xor U16133 (N_16133,N_15939,N_15855);
nand U16134 (N_16134,N_15923,N_15966);
and U16135 (N_16135,N_15803,N_15867);
and U16136 (N_16136,N_15989,N_15932);
or U16137 (N_16137,N_15853,N_15891);
nor U16138 (N_16138,N_15819,N_15895);
nand U16139 (N_16139,N_15993,N_15871);
nand U16140 (N_16140,N_15867,N_15946);
nand U16141 (N_16141,N_15928,N_15801);
nand U16142 (N_16142,N_15897,N_15912);
nand U16143 (N_16143,N_15972,N_15935);
and U16144 (N_16144,N_15967,N_15923);
and U16145 (N_16145,N_15985,N_15812);
xor U16146 (N_16146,N_15885,N_15915);
and U16147 (N_16147,N_15988,N_15826);
nand U16148 (N_16148,N_15809,N_15829);
or U16149 (N_16149,N_15932,N_15993);
and U16150 (N_16150,N_15863,N_15987);
and U16151 (N_16151,N_15818,N_15971);
or U16152 (N_16152,N_15982,N_15988);
xnor U16153 (N_16153,N_15803,N_15919);
or U16154 (N_16154,N_15841,N_15986);
or U16155 (N_16155,N_15922,N_15956);
and U16156 (N_16156,N_15865,N_15982);
nor U16157 (N_16157,N_15836,N_15874);
nor U16158 (N_16158,N_15835,N_15822);
xnor U16159 (N_16159,N_15907,N_15910);
xnor U16160 (N_16160,N_15992,N_15845);
and U16161 (N_16161,N_15991,N_15815);
nor U16162 (N_16162,N_15845,N_15958);
and U16163 (N_16163,N_15833,N_15934);
or U16164 (N_16164,N_15830,N_15866);
or U16165 (N_16165,N_15930,N_15831);
nand U16166 (N_16166,N_15814,N_15962);
xnor U16167 (N_16167,N_15897,N_15961);
and U16168 (N_16168,N_15951,N_15959);
xnor U16169 (N_16169,N_15818,N_15807);
and U16170 (N_16170,N_15984,N_15930);
nand U16171 (N_16171,N_15833,N_15860);
xor U16172 (N_16172,N_15871,N_15923);
nor U16173 (N_16173,N_15864,N_15820);
nor U16174 (N_16174,N_15971,N_15867);
nor U16175 (N_16175,N_15812,N_15990);
xor U16176 (N_16176,N_15904,N_15896);
and U16177 (N_16177,N_15844,N_15874);
nor U16178 (N_16178,N_15882,N_15888);
or U16179 (N_16179,N_15877,N_15932);
or U16180 (N_16180,N_15815,N_15953);
nand U16181 (N_16181,N_15944,N_15972);
xnor U16182 (N_16182,N_15974,N_15848);
xnor U16183 (N_16183,N_15826,N_15960);
nor U16184 (N_16184,N_15947,N_15931);
and U16185 (N_16185,N_15825,N_15829);
and U16186 (N_16186,N_15947,N_15856);
nor U16187 (N_16187,N_15845,N_15837);
nand U16188 (N_16188,N_15804,N_15924);
nor U16189 (N_16189,N_15949,N_15905);
nor U16190 (N_16190,N_15970,N_15841);
and U16191 (N_16191,N_15953,N_15839);
nand U16192 (N_16192,N_15850,N_15936);
xnor U16193 (N_16193,N_15837,N_15849);
nor U16194 (N_16194,N_15855,N_15997);
nor U16195 (N_16195,N_15964,N_15956);
xnor U16196 (N_16196,N_15822,N_15862);
or U16197 (N_16197,N_15923,N_15919);
xnor U16198 (N_16198,N_15981,N_15860);
xor U16199 (N_16199,N_15933,N_15962);
nand U16200 (N_16200,N_16030,N_16097);
nand U16201 (N_16201,N_16194,N_16181);
nand U16202 (N_16202,N_16076,N_16034);
or U16203 (N_16203,N_16058,N_16071);
and U16204 (N_16204,N_16153,N_16118);
nor U16205 (N_16205,N_16074,N_16197);
xnor U16206 (N_16206,N_16063,N_16135);
xor U16207 (N_16207,N_16137,N_16077);
and U16208 (N_16208,N_16022,N_16041);
nor U16209 (N_16209,N_16141,N_16019);
xor U16210 (N_16210,N_16003,N_16116);
or U16211 (N_16211,N_16112,N_16053);
xor U16212 (N_16212,N_16007,N_16160);
and U16213 (N_16213,N_16104,N_16059);
nor U16214 (N_16214,N_16027,N_16047);
and U16215 (N_16215,N_16146,N_16064);
and U16216 (N_16216,N_16023,N_16017);
and U16217 (N_16217,N_16015,N_16098);
xor U16218 (N_16218,N_16109,N_16073);
and U16219 (N_16219,N_16067,N_16111);
xnor U16220 (N_16220,N_16102,N_16176);
and U16221 (N_16221,N_16149,N_16081);
nand U16222 (N_16222,N_16052,N_16139);
xor U16223 (N_16223,N_16179,N_16048);
or U16224 (N_16224,N_16157,N_16156);
nand U16225 (N_16225,N_16188,N_16178);
xor U16226 (N_16226,N_16050,N_16129);
nor U16227 (N_16227,N_16173,N_16126);
nor U16228 (N_16228,N_16091,N_16164);
nor U16229 (N_16229,N_16080,N_16183);
and U16230 (N_16230,N_16026,N_16079);
nor U16231 (N_16231,N_16083,N_16100);
xor U16232 (N_16232,N_16094,N_16168);
nor U16233 (N_16233,N_16087,N_16046);
nor U16234 (N_16234,N_16029,N_16088);
nor U16235 (N_16235,N_16170,N_16195);
and U16236 (N_16236,N_16001,N_16128);
and U16237 (N_16237,N_16175,N_16006);
xnor U16238 (N_16238,N_16166,N_16145);
and U16239 (N_16239,N_16103,N_16082);
nor U16240 (N_16240,N_16171,N_16038);
xnor U16241 (N_16241,N_16158,N_16016);
xor U16242 (N_16242,N_16042,N_16099);
xnor U16243 (N_16243,N_16165,N_16199);
nand U16244 (N_16244,N_16096,N_16024);
or U16245 (N_16245,N_16152,N_16115);
or U16246 (N_16246,N_16093,N_16189);
nor U16247 (N_16247,N_16085,N_16033);
nor U16248 (N_16248,N_16070,N_16054);
nor U16249 (N_16249,N_16198,N_16185);
xnor U16250 (N_16250,N_16132,N_16119);
nor U16251 (N_16251,N_16035,N_16114);
and U16252 (N_16252,N_16133,N_16108);
or U16253 (N_16253,N_16084,N_16174);
nand U16254 (N_16254,N_16127,N_16075);
and U16255 (N_16255,N_16043,N_16037);
nand U16256 (N_16256,N_16028,N_16013);
nor U16257 (N_16257,N_16177,N_16147);
nor U16258 (N_16258,N_16123,N_16196);
nand U16259 (N_16259,N_16182,N_16140);
nand U16260 (N_16260,N_16009,N_16186);
and U16261 (N_16261,N_16092,N_16187);
nor U16262 (N_16262,N_16122,N_16131);
nor U16263 (N_16263,N_16072,N_16142);
xnor U16264 (N_16264,N_16056,N_16036);
nand U16265 (N_16265,N_16089,N_16014);
or U16266 (N_16266,N_16130,N_16044);
nand U16267 (N_16267,N_16032,N_16154);
xnor U16268 (N_16268,N_16120,N_16068);
and U16269 (N_16269,N_16025,N_16113);
nor U16270 (N_16270,N_16057,N_16125);
or U16271 (N_16271,N_16010,N_16004);
and U16272 (N_16272,N_16107,N_16143);
and U16273 (N_16273,N_16138,N_16169);
nor U16274 (N_16274,N_16061,N_16151);
nand U16275 (N_16275,N_16095,N_16163);
nor U16276 (N_16276,N_16172,N_16192);
or U16277 (N_16277,N_16090,N_16106);
nand U16278 (N_16278,N_16191,N_16021);
and U16279 (N_16279,N_16051,N_16162);
or U16280 (N_16280,N_16144,N_16066);
or U16281 (N_16281,N_16049,N_16062);
nand U16282 (N_16282,N_16124,N_16008);
nor U16283 (N_16283,N_16105,N_16180);
and U16284 (N_16284,N_16148,N_16134);
and U16285 (N_16285,N_16002,N_16159);
nand U16286 (N_16286,N_16078,N_16184);
nand U16287 (N_16287,N_16045,N_16086);
and U16288 (N_16288,N_16018,N_16117);
nor U16289 (N_16289,N_16121,N_16110);
and U16290 (N_16290,N_16069,N_16040);
or U16291 (N_16291,N_16136,N_16000);
xnor U16292 (N_16292,N_16161,N_16060);
or U16293 (N_16293,N_16055,N_16011);
xor U16294 (N_16294,N_16193,N_16012);
or U16295 (N_16295,N_16031,N_16020);
or U16296 (N_16296,N_16167,N_16065);
nand U16297 (N_16297,N_16101,N_16155);
or U16298 (N_16298,N_16190,N_16150);
nor U16299 (N_16299,N_16039,N_16005);
nor U16300 (N_16300,N_16073,N_16074);
xor U16301 (N_16301,N_16005,N_16086);
nor U16302 (N_16302,N_16181,N_16055);
nor U16303 (N_16303,N_16132,N_16092);
nand U16304 (N_16304,N_16156,N_16110);
nor U16305 (N_16305,N_16066,N_16120);
xnor U16306 (N_16306,N_16116,N_16076);
xor U16307 (N_16307,N_16133,N_16192);
nor U16308 (N_16308,N_16106,N_16073);
nor U16309 (N_16309,N_16120,N_16072);
xnor U16310 (N_16310,N_16177,N_16012);
nand U16311 (N_16311,N_16051,N_16166);
nor U16312 (N_16312,N_16106,N_16159);
or U16313 (N_16313,N_16016,N_16168);
and U16314 (N_16314,N_16077,N_16078);
xnor U16315 (N_16315,N_16121,N_16096);
or U16316 (N_16316,N_16099,N_16037);
or U16317 (N_16317,N_16112,N_16051);
and U16318 (N_16318,N_16071,N_16154);
and U16319 (N_16319,N_16029,N_16175);
nor U16320 (N_16320,N_16046,N_16162);
or U16321 (N_16321,N_16044,N_16171);
and U16322 (N_16322,N_16150,N_16032);
and U16323 (N_16323,N_16004,N_16006);
xnor U16324 (N_16324,N_16138,N_16022);
xnor U16325 (N_16325,N_16087,N_16088);
nor U16326 (N_16326,N_16087,N_16082);
nor U16327 (N_16327,N_16066,N_16177);
or U16328 (N_16328,N_16135,N_16023);
nand U16329 (N_16329,N_16033,N_16149);
nor U16330 (N_16330,N_16153,N_16036);
or U16331 (N_16331,N_16000,N_16157);
and U16332 (N_16332,N_16068,N_16161);
and U16333 (N_16333,N_16149,N_16000);
or U16334 (N_16334,N_16155,N_16198);
nor U16335 (N_16335,N_16051,N_16024);
nor U16336 (N_16336,N_16187,N_16148);
nor U16337 (N_16337,N_16003,N_16159);
xnor U16338 (N_16338,N_16100,N_16107);
and U16339 (N_16339,N_16171,N_16198);
xnor U16340 (N_16340,N_16144,N_16091);
and U16341 (N_16341,N_16058,N_16030);
or U16342 (N_16342,N_16031,N_16116);
and U16343 (N_16343,N_16008,N_16007);
or U16344 (N_16344,N_16111,N_16186);
or U16345 (N_16345,N_16170,N_16029);
and U16346 (N_16346,N_16133,N_16169);
xor U16347 (N_16347,N_16109,N_16039);
nor U16348 (N_16348,N_16124,N_16119);
nand U16349 (N_16349,N_16198,N_16136);
and U16350 (N_16350,N_16120,N_16032);
and U16351 (N_16351,N_16066,N_16173);
and U16352 (N_16352,N_16176,N_16057);
and U16353 (N_16353,N_16024,N_16179);
xnor U16354 (N_16354,N_16196,N_16155);
and U16355 (N_16355,N_16093,N_16135);
nand U16356 (N_16356,N_16176,N_16109);
or U16357 (N_16357,N_16099,N_16104);
nand U16358 (N_16358,N_16015,N_16037);
nand U16359 (N_16359,N_16120,N_16186);
xnor U16360 (N_16360,N_16010,N_16174);
xor U16361 (N_16361,N_16176,N_16111);
or U16362 (N_16362,N_16088,N_16165);
nand U16363 (N_16363,N_16191,N_16070);
xnor U16364 (N_16364,N_16072,N_16069);
or U16365 (N_16365,N_16172,N_16140);
xor U16366 (N_16366,N_16133,N_16186);
or U16367 (N_16367,N_16084,N_16035);
and U16368 (N_16368,N_16066,N_16199);
or U16369 (N_16369,N_16170,N_16042);
or U16370 (N_16370,N_16008,N_16064);
nor U16371 (N_16371,N_16108,N_16056);
nand U16372 (N_16372,N_16174,N_16171);
nand U16373 (N_16373,N_16190,N_16113);
or U16374 (N_16374,N_16073,N_16184);
nor U16375 (N_16375,N_16085,N_16088);
and U16376 (N_16376,N_16002,N_16026);
xor U16377 (N_16377,N_16177,N_16079);
or U16378 (N_16378,N_16058,N_16121);
nand U16379 (N_16379,N_16072,N_16184);
and U16380 (N_16380,N_16122,N_16070);
or U16381 (N_16381,N_16002,N_16021);
nor U16382 (N_16382,N_16102,N_16050);
nor U16383 (N_16383,N_16053,N_16143);
nand U16384 (N_16384,N_16114,N_16176);
nand U16385 (N_16385,N_16018,N_16090);
nor U16386 (N_16386,N_16084,N_16040);
nand U16387 (N_16387,N_16053,N_16179);
and U16388 (N_16388,N_16047,N_16194);
and U16389 (N_16389,N_16180,N_16077);
or U16390 (N_16390,N_16154,N_16072);
nor U16391 (N_16391,N_16177,N_16129);
or U16392 (N_16392,N_16073,N_16015);
nand U16393 (N_16393,N_16093,N_16054);
nand U16394 (N_16394,N_16142,N_16095);
or U16395 (N_16395,N_16110,N_16068);
and U16396 (N_16396,N_16073,N_16126);
or U16397 (N_16397,N_16139,N_16035);
nor U16398 (N_16398,N_16170,N_16004);
or U16399 (N_16399,N_16144,N_16140);
or U16400 (N_16400,N_16316,N_16251);
and U16401 (N_16401,N_16368,N_16322);
nor U16402 (N_16402,N_16265,N_16320);
or U16403 (N_16403,N_16239,N_16375);
xor U16404 (N_16404,N_16225,N_16308);
or U16405 (N_16405,N_16240,N_16396);
or U16406 (N_16406,N_16291,N_16285);
nor U16407 (N_16407,N_16301,N_16259);
xor U16408 (N_16408,N_16202,N_16398);
xor U16409 (N_16409,N_16312,N_16311);
xor U16410 (N_16410,N_16217,N_16223);
xnor U16411 (N_16411,N_16277,N_16354);
xnor U16412 (N_16412,N_16255,N_16208);
xnor U16413 (N_16413,N_16374,N_16342);
or U16414 (N_16414,N_16226,N_16349);
or U16415 (N_16415,N_16343,N_16260);
and U16416 (N_16416,N_16245,N_16262);
xor U16417 (N_16417,N_16231,N_16282);
xor U16418 (N_16418,N_16362,N_16356);
and U16419 (N_16419,N_16336,N_16234);
xnor U16420 (N_16420,N_16203,N_16298);
or U16421 (N_16421,N_16325,N_16244);
nand U16422 (N_16422,N_16317,N_16241);
xor U16423 (N_16423,N_16272,N_16377);
nand U16424 (N_16424,N_16395,N_16273);
nor U16425 (N_16425,N_16366,N_16289);
or U16426 (N_16426,N_16337,N_16220);
nor U16427 (N_16427,N_16254,N_16328);
or U16428 (N_16428,N_16399,N_16383);
or U16429 (N_16429,N_16352,N_16313);
or U16430 (N_16430,N_16393,N_16266);
nor U16431 (N_16431,N_16380,N_16249);
and U16432 (N_16432,N_16387,N_16237);
and U16433 (N_16433,N_16267,N_16390);
xnor U16434 (N_16434,N_16307,N_16309);
nand U16435 (N_16435,N_16385,N_16269);
and U16436 (N_16436,N_16286,N_16274);
xnor U16437 (N_16437,N_16351,N_16391);
nor U16438 (N_16438,N_16229,N_16324);
nor U16439 (N_16439,N_16278,N_16252);
xnor U16440 (N_16440,N_16389,N_16315);
and U16441 (N_16441,N_16341,N_16388);
or U16442 (N_16442,N_16303,N_16364);
or U16443 (N_16443,N_16215,N_16357);
or U16444 (N_16444,N_16279,N_16264);
or U16445 (N_16445,N_16297,N_16238);
or U16446 (N_16446,N_16372,N_16292);
xor U16447 (N_16447,N_16201,N_16263);
or U16448 (N_16448,N_16360,N_16230);
xor U16449 (N_16449,N_16211,N_16228);
nor U16450 (N_16450,N_16331,N_16200);
xnor U16451 (N_16451,N_16280,N_16296);
and U16452 (N_16452,N_16378,N_16250);
and U16453 (N_16453,N_16361,N_16365);
xor U16454 (N_16454,N_16386,N_16310);
nand U16455 (N_16455,N_16379,N_16258);
or U16456 (N_16456,N_16353,N_16276);
and U16457 (N_16457,N_16243,N_16384);
nor U16458 (N_16458,N_16204,N_16275);
or U16459 (N_16459,N_16306,N_16283);
nand U16460 (N_16460,N_16305,N_16344);
nand U16461 (N_16461,N_16300,N_16261);
and U16462 (N_16462,N_16367,N_16346);
or U16463 (N_16463,N_16340,N_16246);
nor U16464 (N_16464,N_16293,N_16358);
and U16465 (N_16465,N_16330,N_16381);
and U16466 (N_16466,N_16212,N_16394);
nand U16467 (N_16467,N_16271,N_16221);
and U16468 (N_16468,N_16326,N_16222);
nor U16469 (N_16469,N_16319,N_16206);
and U16470 (N_16470,N_16235,N_16270);
and U16471 (N_16471,N_16248,N_16247);
xor U16472 (N_16472,N_16294,N_16207);
xor U16473 (N_16473,N_16257,N_16332);
nand U16474 (N_16474,N_16314,N_16288);
nand U16475 (N_16475,N_16232,N_16302);
xor U16476 (N_16476,N_16339,N_16209);
nand U16477 (N_16477,N_16355,N_16345);
xor U16478 (N_16478,N_16338,N_16347);
nand U16479 (N_16479,N_16335,N_16350);
nor U16480 (N_16480,N_16321,N_16256);
and U16481 (N_16481,N_16371,N_16397);
or U16482 (N_16482,N_16327,N_16376);
nor U16483 (N_16483,N_16236,N_16216);
or U16484 (N_16484,N_16290,N_16287);
xnor U16485 (N_16485,N_16373,N_16370);
xnor U16486 (N_16486,N_16382,N_16268);
nor U16487 (N_16487,N_16334,N_16284);
nor U16488 (N_16488,N_16218,N_16253);
nor U16489 (N_16489,N_16318,N_16323);
and U16490 (N_16490,N_16299,N_16210);
and U16491 (N_16491,N_16369,N_16304);
nor U16492 (N_16492,N_16205,N_16219);
xnor U16493 (N_16493,N_16227,N_16224);
xnor U16494 (N_16494,N_16329,N_16233);
nand U16495 (N_16495,N_16242,N_16359);
nand U16496 (N_16496,N_16392,N_16348);
nor U16497 (N_16497,N_16333,N_16213);
nor U16498 (N_16498,N_16214,N_16281);
xnor U16499 (N_16499,N_16295,N_16363);
nand U16500 (N_16500,N_16384,N_16321);
xor U16501 (N_16501,N_16377,N_16376);
nand U16502 (N_16502,N_16284,N_16384);
or U16503 (N_16503,N_16280,N_16243);
xnor U16504 (N_16504,N_16276,N_16294);
nand U16505 (N_16505,N_16381,N_16232);
and U16506 (N_16506,N_16343,N_16370);
nand U16507 (N_16507,N_16283,N_16334);
nor U16508 (N_16508,N_16386,N_16347);
xnor U16509 (N_16509,N_16305,N_16206);
nand U16510 (N_16510,N_16210,N_16394);
nor U16511 (N_16511,N_16358,N_16215);
nand U16512 (N_16512,N_16346,N_16396);
nor U16513 (N_16513,N_16217,N_16274);
nor U16514 (N_16514,N_16385,N_16272);
xor U16515 (N_16515,N_16317,N_16350);
xor U16516 (N_16516,N_16247,N_16312);
and U16517 (N_16517,N_16223,N_16317);
nor U16518 (N_16518,N_16229,N_16392);
nor U16519 (N_16519,N_16250,N_16233);
nor U16520 (N_16520,N_16200,N_16293);
or U16521 (N_16521,N_16203,N_16268);
nand U16522 (N_16522,N_16396,N_16215);
or U16523 (N_16523,N_16225,N_16329);
or U16524 (N_16524,N_16245,N_16378);
or U16525 (N_16525,N_16222,N_16299);
and U16526 (N_16526,N_16331,N_16298);
nand U16527 (N_16527,N_16381,N_16287);
xor U16528 (N_16528,N_16260,N_16355);
xnor U16529 (N_16529,N_16294,N_16332);
or U16530 (N_16530,N_16292,N_16255);
xnor U16531 (N_16531,N_16312,N_16262);
and U16532 (N_16532,N_16245,N_16292);
nor U16533 (N_16533,N_16201,N_16292);
nor U16534 (N_16534,N_16346,N_16279);
or U16535 (N_16535,N_16213,N_16206);
nor U16536 (N_16536,N_16236,N_16333);
nand U16537 (N_16537,N_16293,N_16252);
nand U16538 (N_16538,N_16371,N_16318);
nand U16539 (N_16539,N_16337,N_16252);
nor U16540 (N_16540,N_16232,N_16268);
or U16541 (N_16541,N_16334,N_16338);
nand U16542 (N_16542,N_16366,N_16346);
nor U16543 (N_16543,N_16222,N_16343);
nor U16544 (N_16544,N_16236,N_16386);
and U16545 (N_16545,N_16335,N_16258);
and U16546 (N_16546,N_16254,N_16236);
and U16547 (N_16547,N_16267,N_16323);
xor U16548 (N_16548,N_16385,N_16225);
nand U16549 (N_16549,N_16214,N_16292);
nor U16550 (N_16550,N_16243,N_16349);
nor U16551 (N_16551,N_16270,N_16269);
xor U16552 (N_16552,N_16223,N_16268);
xnor U16553 (N_16553,N_16389,N_16349);
or U16554 (N_16554,N_16333,N_16267);
or U16555 (N_16555,N_16272,N_16362);
nand U16556 (N_16556,N_16392,N_16327);
nor U16557 (N_16557,N_16375,N_16253);
or U16558 (N_16558,N_16217,N_16322);
or U16559 (N_16559,N_16257,N_16206);
xor U16560 (N_16560,N_16359,N_16274);
nand U16561 (N_16561,N_16322,N_16246);
nor U16562 (N_16562,N_16212,N_16369);
nand U16563 (N_16563,N_16249,N_16331);
or U16564 (N_16564,N_16234,N_16274);
xor U16565 (N_16565,N_16398,N_16277);
xnor U16566 (N_16566,N_16239,N_16344);
and U16567 (N_16567,N_16295,N_16312);
nand U16568 (N_16568,N_16304,N_16360);
nor U16569 (N_16569,N_16259,N_16290);
nor U16570 (N_16570,N_16292,N_16341);
and U16571 (N_16571,N_16314,N_16302);
xor U16572 (N_16572,N_16222,N_16223);
or U16573 (N_16573,N_16219,N_16270);
and U16574 (N_16574,N_16388,N_16394);
xor U16575 (N_16575,N_16200,N_16247);
xor U16576 (N_16576,N_16359,N_16299);
nor U16577 (N_16577,N_16223,N_16360);
or U16578 (N_16578,N_16326,N_16338);
nor U16579 (N_16579,N_16374,N_16345);
xor U16580 (N_16580,N_16303,N_16343);
nand U16581 (N_16581,N_16334,N_16262);
or U16582 (N_16582,N_16339,N_16395);
nand U16583 (N_16583,N_16219,N_16328);
or U16584 (N_16584,N_16287,N_16373);
xnor U16585 (N_16585,N_16373,N_16302);
nor U16586 (N_16586,N_16389,N_16270);
or U16587 (N_16587,N_16338,N_16302);
nand U16588 (N_16588,N_16276,N_16334);
or U16589 (N_16589,N_16291,N_16387);
or U16590 (N_16590,N_16255,N_16303);
xnor U16591 (N_16591,N_16370,N_16372);
nand U16592 (N_16592,N_16264,N_16286);
and U16593 (N_16593,N_16271,N_16329);
or U16594 (N_16594,N_16292,N_16377);
nor U16595 (N_16595,N_16275,N_16365);
nand U16596 (N_16596,N_16251,N_16321);
nor U16597 (N_16597,N_16227,N_16376);
nor U16598 (N_16598,N_16338,N_16309);
xor U16599 (N_16599,N_16333,N_16201);
and U16600 (N_16600,N_16475,N_16537);
and U16601 (N_16601,N_16561,N_16512);
nor U16602 (N_16602,N_16487,N_16424);
nor U16603 (N_16603,N_16555,N_16465);
nand U16604 (N_16604,N_16458,N_16550);
and U16605 (N_16605,N_16434,N_16562);
or U16606 (N_16606,N_16502,N_16430);
xor U16607 (N_16607,N_16538,N_16428);
or U16608 (N_16608,N_16417,N_16489);
and U16609 (N_16609,N_16484,N_16589);
nor U16610 (N_16610,N_16548,N_16482);
or U16611 (N_16611,N_16407,N_16477);
nor U16612 (N_16612,N_16557,N_16564);
nand U16613 (N_16613,N_16420,N_16520);
nor U16614 (N_16614,N_16490,N_16419);
xnor U16615 (N_16615,N_16497,N_16574);
and U16616 (N_16616,N_16421,N_16583);
nor U16617 (N_16617,N_16585,N_16597);
and U16618 (N_16618,N_16534,N_16441);
or U16619 (N_16619,N_16485,N_16568);
nand U16620 (N_16620,N_16542,N_16570);
xor U16621 (N_16621,N_16586,N_16546);
or U16622 (N_16622,N_16540,N_16456);
nor U16623 (N_16623,N_16529,N_16478);
nand U16624 (N_16624,N_16523,N_16422);
nand U16625 (N_16625,N_16514,N_16535);
or U16626 (N_16626,N_16525,N_16599);
and U16627 (N_16627,N_16431,N_16413);
nand U16628 (N_16628,N_16544,N_16435);
nor U16629 (N_16629,N_16594,N_16440);
and U16630 (N_16630,N_16416,N_16590);
xor U16631 (N_16631,N_16518,N_16469);
xor U16632 (N_16632,N_16439,N_16414);
and U16633 (N_16633,N_16449,N_16498);
nand U16634 (N_16634,N_16411,N_16553);
nand U16635 (N_16635,N_16543,N_16495);
nor U16636 (N_16636,N_16558,N_16426);
and U16637 (N_16637,N_16576,N_16578);
nand U16638 (N_16638,N_16532,N_16447);
xor U16639 (N_16639,N_16471,N_16486);
nor U16640 (N_16640,N_16410,N_16507);
nand U16641 (N_16641,N_16462,N_16463);
and U16642 (N_16642,N_16563,N_16479);
and U16643 (N_16643,N_16443,N_16457);
nor U16644 (N_16644,N_16432,N_16521);
and U16645 (N_16645,N_16598,N_16517);
or U16646 (N_16646,N_16404,N_16433);
or U16647 (N_16647,N_16595,N_16587);
or U16648 (N_16648,N_16400,N_16581);
nand U16649 (N_16649,N_16519,N_16437);
xnor U16650 (N_16650,N_16592,N_16472);
nand U16651 (N_16651,N_16405,N_16536);
nor U16652 (N_16652,N_16442,N_16531);
nor U16653 (N_16653,N_16505,N_16588);
or U16654 (N_16654,N_16539,N_16425);
nor U16655 (N_16655,N_16418,N_16541);
xnor U16656 (N_16656,N_16448,N_16453);
and U16657 (N_16657,N_16466,N_16459);
and U16658 (N_16658,N_16455,N_16513);
nor U16659 (N_16659,N_16470,N_16481);
or U16660 (N_16660,N_16533,N_16580);
or U16661 (N_16661,N_16504,N_16451);
nand U16662 (N_16662,N_16577,N_16450);
nor U16663 (N_16663,N_16579,N_16454);
nand U16664 (N_16664,N_16509,N_16423);
nor U16665 (N_16665,N_16567,N_16545);
and U16666 (N_16666,N_16510,N_16569);
and U16667 (N_16667,N_16412,N_16566);
and U16668 (N_16668,N_16552,N_16584);
or U16669 (N_16669,N_16503,N_16565);
nand U16670 (N_16670,N_16596,N_16491);
nor U16671 (N_16671,N_16494,N_16460);
nand U16672 (N_16672,N_16492,N_16427);
nand U16673 (N_16673,N_16429,N_16508);
or U16674 (N_16674,N_16476,N_16445);
nand U16675 (N_16675,N_16483,N_16515);
and U16676 (N_16676,N_16572,N_16530);
xnor U16677 (N_16677,N_16461,N_16573);
or U16678 (N_16678,N_16403,N_16524);
and U16679 (N_16679,N_16528,N_16408);
nand U16680 (N_16680,N_16500,N_16559);
nand U16681 (N_16681,N_16593,N_16493);
xor U16682 (N_16682,N_16409,N_16549);
nand U16683 (N_16683,N_16452,N_16496);
and U16684 (N_16684,N_16402,N_16551);
nor U16685 (N_16685,N_16474,N_16480);
or U16686 (N_16686,N_16556,N_16499);
nor U16687 (N_16687,N_16527,N_16560);
and U16688 (N_16688,N_16406,N_16571);
and U16689 (N_16689,N_16501,N_16446);
and U16690 (N_16690,N_16438,N_16473);
nand U16691 (N_16691,N_16516,N_16444);
and U16692 (N_16692,N_16436,N_16506);
or U16693 (N_16693,N_16547,N_16464);
or U16694 (N_16694,N_16575,N_16488);
nor U16695 (N_16695,N_16468,N_16582);
or U16696 (N_16696,N_16401,N_16467);
or U16697 (N_16697,N_16591,N_16511);
nand U16698 (N_16698,N_16554,N_16415);
xnor U16699 (N_16699,N_16522,N_16526);
and U16700 (N_16700,N_16516,N_16400);
xnor U16701 (N_16701,N_16566,N_16503);
nor U16702 (N_16702,N_16505,N_16448);
nor U16703 (N_16703,N_16432,N_16491);
or U16704 (N_16704,N_16594,N_16447);
or U16705 (N_16705,N_16417,N_16580);
nor U16706 (N_16706,N_16588,N_16496);
and U16707 (N_16707,N_16552,N_16557);
nor U16708 (N_16708,N_16412,N_16447);
and U16709 (N_16709,N_16598,N_16501);
or U16710 (N_16710,N_16558,N_16463);
xor U16711 (N_16711,N_16436,N_16482);
nor U16712 (N_16712,N_16478,N_16531);
xor U16713 (N_16713,N_16489,N_16406);
nand U16714 (N_16714,N_16561,N_16547);
and U16715 (N_16715,N_16595,N_16406);
xnor U16716 (N_16716,N_16412,N_16460);
nor U16717 (N_16717,N_16519,N_16456);
nand U16718 (N_16718,N_16455,N_16474);
or U16719 (N_16719,N_16571,N_16451);
nor U16720 (N_16720,N_16461,N_16547);
nand U16721 (N_16721,N_16493,N_16412);
nand U16722 (N_16722,N_16567,N_16401);
xnor U16723 (N_16723,N_16579,N_16599);
nand U16724 (N_16724,N_16453,N_16554);
nand U16725 (N_16725,N_16450,N_16526);
nand U16726 (N_16726,N_16556,N_16506);
nor U16727 (N_16727,N_16439,N_16545);
xor U16728 (N_16728,N_16586,N_16598);
and U16729 (N_16729,N_16470,N_16432);
xnor U16730 (N_16730,N_16452,N_16498);
nand U16731 (N_16731,N_16428,N_16572);
nand U16732 (N_16732,N_16575,N_16493);
xnor U16733 (N_16733,N_16576,N_16584);
or U16734 (N_16734,N_16480,N_16401);
nor U16735 (N_16735,N_16467,N_16432);
xor U16736 (N_16736,N_16589,N_16485);
and U16737 (N_16737,N_16492,N_16521);
xor U16738 (N_16738,N_16497,N_16403);
and U16739 (N_16739,N_16407,N_16591);
nor U16740 (N_16740,N_16478,N_16508);
nand U16741 (N_16741,N_16439,N_16521);
or U16742 (N_16742,N_16471,N_16409);
nand U16743 (N_16743,N_16533,N_16503);
and U16744 (N_16744,N_16462,N_16543);
xnor U16745 (N_16745,N_16432,N_16414);
nand U16746 (N_16746,N_16502,N_16482);
or U16747 (N_16747,N_16469,N_16564);
or U16748 (N_16748,N_16568,N_16596);
nand U16749 (N_16749,N_16538,N_16590);
and U16750 (N_16750,N_16440,N_16400);
or U16751 (N_16751,N_16540,N_16466);
and U16752 (N_16752,N_16499,N_16571);
or U16753 (N_16753,N_16455,N_16508);
nor U16754 (N_16754,N_16560,N_16438);
nor U16755 (N_16755,N_16461,N_16566);
nand U16756 (N_16756,N_16515,N_16524);
xor U16757 (N_16757,N_16407,N_16485);
or U16758 (N_16758,N_16480,N_16435);
nor U16759 (N_16759,N_16582,N_16453);
or U16760 (N_16760,N_16425,N_16583);
nand U16761 (N_16761,N_16422,N_16492);
xnor U16762 (N_16762,N_16426,N_16511);
xor U16763 (N_16763,N_16498,N_16497);
nor U16764 (N_16764,N_16513,N_16408);
nor U16765 (N_16765,N_16412,N_16497);
and U16766 (N_16766,N_16460,N_16565);
or U16767 (N_16767,N_16435,N_16567);
or U16768 (N_16768,N_16411,N_16563);
or U16769 (N_16769,N_16533,N_16467);
nand U16770 (N_16770,N_16452,N_16492);
xnor U16771 (N_16771,N_16584,N_16469);
or U16772 (N_16772,N_16542,N_16453);
nand U16773 (N_16773,N_16593,N_16484);
or U16774 (N_16774,N_16599,N_16524);
or U16775 (N_16775,N_16497,N_16459);
and U16776 (N_16776,N_16468,N_16565);
xnor U16777 (N_16777,N_16447,N_16402);
and U16778 (N_16778,N_16470,N_16450);
and U16779 (N_16779,N_16412,N_16486);
nand U16780 (N_16780,N_16470,N_16525);
xnor U16781 (N_16781,N_16502,N_16509);
nand U16782 (N_16782,N_16570,N_16411);
nor U16783 (N_16783,N_16515,N_16486);
nor U16784 (N_16784,N_16446,N_16554);
xnor U16785 (N_16785,N_16543,N_16498);
and U16786 (N_16786,N_16444,N_16554);
nor U16787 (N_16787,N_16552,N_16492);
xnor U16788 (N_16788,N_16492,N_16491);
nor U16789 (N_16789,N_16460,N_16432);
nor U16790 (N_16790,N_16574,N_16410);
or U16791 (N_16791,N_16475,N_16523);
or U16792 (N_16792,N_16570,N_16534);
nor U16793 (N_16793,N_16570,N_16491);
or U16794 (N_16794,N_16444,N_16495);
nand U16795 (N_16795,N_16572,N_16570);
and U16796 (N_16796,N_16561,N_16553);
nand U16797 (N_16797,N_16478,N_16588);
nor U16798 (N_16798,N_16418,N_16548);
and U16799 (N_16799,N_16439,N_16482);
and U16800 (N_16800,N_16731,N_16791);
nor U16801 (N_16801,N_16683,N_16698);
xnor U16802 (N_16802,N_16672,N_16738);
or U16803 (N_16803,N_16736,N_16623);
nor U16804 (N_16804,N_16705,N_16647);
and U16805 (N_16805,N_16638,N_16628);
nor U16806 (N_16806,N_16675,N_16745);
xor U16807 (N_16807,N_16720,N_16733);
or U16808 (N_16808,N_16786,N_16663);
nand U16809 (N_16809,N_16740,N_16766);
nand U16810 (N_16810,N_16709,N_16783);
xor U16811 (N_16811,N_16637,N_16797);
or U16812 (N_16812,N_16689,N_16760);
nor U16813 (N_16813,N_16613,N_16771);
xor U16814 (N_16814,N_16798,N_16643);
or U16815 (N_16815,N_16608,N_16601);
xnor U16816 (N_16816,N_16715,N_16767);
nor U16817 (N_16817,N_16655,N_16653);
nand U16818 (N_16818,N_16617,N_16735);
xnor U16819 (N_16819,N_16790,N_16614);
xor U16820 (N_16820,N_16780,N_16724);
and U16821 (N_16821,N_16743,N_16606);
nand U16822 (N_16822,N_16764,N_16659);
nand U16823 (N_16823,N_16769,N_16629);
nor U16824 (N_16824,N_16772,N_16691);
nor U16825 (N_16825,N_16710,N_16702);
xor U16826 (N_16826,N_16749,N_16762);
nand U16827 (N_16827,N_16602,N_16773);
nand U16828 (N_16828,N_16630,N_16604);
or U16829 (N_16829,N_16678,N_16714);
nor U16830 (N_16830,N_16716,N_16666);
or U16831 (N_16831,N_16632,N_16779);
nor U16832 (N_16832,N_16744,N_16785);
or U16833 (N_16833,N_16670,N_16778);
or U16834 (N_16834,N_16770,N_16753);
nand U16835 (N_16835,N_16685,N_16750);
and U16836 (N_16836,N_16758,N_16642);
xor U16837 (N_16837,N_16761,N_16667);
or U16838 (N_16838,N_16686,N_16603);
nor U16839 (N_16839,N_16665,N_16730);
and U16840 (N_16840,N_16616,N_16631);
nand U16841 (N_16841,N_16793,N_16746);
xor U16842 (N_16842,N_16656,N_16694);
nand U16843 (N_16843,N_16671,N_16765);
and U16844 (N_16844,N_16679,N_16742);
nand U16845 (N_16845,N_16695,N_16756);
nor U16846 (N_16846,N_16607,N_16657);
nand U16847 (N_16847,N_16704,N_16737);
or U16848 (N_16848,N_16649,N_16621);
xnor U16849 (N_16849,N_16781,N_16741);
and U16850 (N_16850,N_16755,N_16759);
or U16851 (N_16851,N_16725,N_16640);
nand U16852 (N_16852,N_16687,N_16624);
xor U16853 (N_16853,N_16754,N_16696);
and U16854 (N_16854,N_16639,N_16795);
nor U16855 (N_16855,N_16774,N_16703);
nand U16856 (N_16856,N_16697,N_16747);
xnor U16857 (N_16857,N_16728,N_16626);
and U16858 (N_16858,N_16644,N_16717);
nor U16859 (N_16859,N_16719,N_16751);
nor U16860 (N_16860,N_16723,N_16713);
and U16861 (N_16861,N_16684,N_16796);
and U16862 (N_16862,N_16775,N_16726);
or U16863 (N_16863,N_16768,N_16700);
xor U16864 (N_16864,N_16650,N_16712);
and U16865 (N_16865,N_16622,N_16763);
or U16866 (N_16866,N_16784,N_16633);
xnor U16867 (N_16867,N_16636,N_16611);
and U16868 (N_16868,N_16708,N_16727);
or U16869 (N_16869,N_16618,N_16619);
or U16870 (N_16870,N_16699,N_16799);
nand U16871 (N_16871,N_16688,N_16635);
nor U16872 (N_16872,N_16701,N_16794);
nor U16873 (N_16873,N_16661,N_16748);
or U16874 (N_16874,N_16722,N_16729);
and U16875 (N_16875,N_16707,N_16680);
nor U16876 (N_16876,N_16777,N_16711);
and U16877 (N_16877,N_16641,N_16648);
xnor U16878 (N_16878,N_16627,N_16662);
xnor U16879 (N_16879,N_16757,N_16693);
xnor U16880 (N_16880,N_16739,N_16706);
xnor U16881 (N_16881,N_16787,N_16625);
or U16882 (N_16882,N_16674,N_16654);
and U16883 (N_16883,N_16776,N_16664);
nor U16884 (N_16884,N_16752,N_16732);
or U16885 (N_16885,N_16620,N_16721);
and U16886 (N_16886,N_16692,N_16677);
or U16887 (N_16887,N_16609,N_16634);
nor U16888 (N_16888,N_16610,N_16682);
xor U16889 (N_16889,N_16668,N_16652);
or U16890 (N_16890,N_16646,N_16658);
nor U16891 (N_16891,N_16660,N_16734);
nand U16892 (N_16892,N_16789,N_16681);
nand U16893 (N_16893,N_16669,N_16792);
nand U16894 (N_16894,N_16615,N_16788);
nor U16895 (N_16895,N_16645,N_16600);
nor U16896 (N_16896,N_16718,N_16782);
xor U16897 (N_16897,N_16690,N_16676);
nor U16898 (N_16898,N_16651,N_16612);
xnor U16899 (N_16899,N_16673,N_16605);
and U16900 (N_16900,N_16615,N_16632);
nand U16901 (N_16901,N_16795,N_16723);
nor U16902 (N_16902,N_16694,N_16732);
or U16903 (N_16903,N_16635,N_16676);
or U16904 (N_16904,N_16779,N_16740);
nand U16905 (N_16905,N_16783,N_16656);
and U16906 (N_16906,N_16622,N_16609);
xor U16907 (N_16907,N_16731,N_16760);
nand U16908 (N_16908,N_16701,N_16607);
or U16909 (N_16909,N_16690,N_16654);
and U16910 (N_16910,N_16774,N_16666);
and U16911 (N_16911,N_16714,N_16725);
xnor U16912 (N_16912,N_16681,N_16743);
or U16913 (N_16913,N_16681,N_16649);
or U16914 (N_16914,N_16682,N_16696);
or U16915 (N_16915,N_16700,N_16749);
and U16916 (N_16916,N_16651,N_16796);
nand U16917 (N_16917,N_16622,N_16649);
xor U16918 (N_16918,N_16700,N_16697);
nand U16919 (N_16919,N_16650,N_16603);
nor U16920 (N_16920,N_16736,N_16635);
nor U16921 (N_16921,N_16757,N_16658);
xor U16922 (N_16922,N_16691,N_16716);
or U16923 (N_16923,N_16670,N_16709);
xnor U16924 (N_16924,N_16614,N_16757);
or U16925 (N_16925,N_16642,N_16760);
nor U16926 (N_16926,N_16766,N_16732);
and U16927 (N_16927,N_16782,N_16747);
nand U16928 (N_16928,N_16788,N_16609);
and U16929 (N_16929,N_16763,N_16776);
and U16930 (N_16930,N_16613,N_16703);
nor U16931 (N_16931,N_16763,N_16755);
or U16932 (N_16932,N_16697,N_16716);
nand U16933 (N_16933,N_16626,N_16693);
nor U16934 (N_16934,N_16732,N_16615);
nor U16935 (N_16935,N_16680,N_16741);
or U16936 (N_16936,N_16764,N_16626);
nor U16937 (N_16937,N_16641,N_16626);
and U16938 (N_16938,N_16712,N_16685);
and U16939 (N_16939,N_16698,N_16701);
and U16940 (N_16940,N_16784,N_16765);
or U16941 (N_16941,N_16790,N_16666);
nand U16942 (N_16942,N_16618,N_16796);
nor U16943 (N_16943,N_16727,N_16667);
xnor U16944 (N_16944,N_16607,N_16764);
and U16945 (N_16945,N_16605,N_16601);
or U16946 (N_16946,N_16604,N_16602);
xnor U16947 (N_16947,N_16653,N_16776);
nand U16948 (N_16948,N_16685,N_16779);
or U16949 (N_16949,N_16797,N_16760);
nor U16950 (N_16950,N_16600,N_16727);
and U16951 (N_16951,N_16619,N_16718);
and U16952 (N_16952,N_16639,N_16647);
nor U16953 (N_16953,N_16626,N_16776);
nand U16954 (N_16954,N_16790,N_16655);
and U16955 (N_16955,N_16645,N_16604);
and U16956 (N_16956,N_16655,N_16732);
or U16957 (N_16957,N_16604,N_16753);
xnor U16958 (N_16958,N_16601,N_16611);
nand U16959 (N_16959,N_16683,N_16621);
nor U16960 (N_16960,N_16689,N_16704);
nor U16961 (N_16961,N_16684,N_16650);
or U16962 (N_16962,N_16612,N_16769);
and U16963 (N_16963,N_16787,N_16773);
or U16964 (N_16964,N_16617,N_16689);
nand U16965 (N_16965,N_16602,N_16697);
or U16966 (N_16966,N_16712,N_16644);
and U16967 (N_16967,N_16753,N_16687);
nand U16968 (N_16968,N_16746,N_16771);
nand U16969 (N_16969,N_16723,N_16654);
nor U16970 (N_16970,N_16657,N_16648);
and U16971 (N_16971,N_16730,N_16747);
nor U16972 (N_16972,N_16729,N_16650);
nand U16973 (N_16973,N_16620,N_16763);
and U16974 (N_16974,N_16743,N_16692);
or U16975 (N_16975,N_16794,N_16648);
or U16976 (N_16976,N_16760,N_16622);
nand U16977 (N_16977,N_16628,N_16782);
and U16978 (N_16978,N_16699,N_16617);
nor U16979 (N_16979,N_16705,N_16664);
nor U16980 (N_16980,N_16766,N_16692);
nand U16981 (N_16981,N_16782,N_16798);
nor U16982 (N_16982,N_16661,N_16690);
or U16983 (N_16983,N_16670,N_16683);
and U16984 (N_16984,N_16608,N_16677);
or U16985 (N_16985,N_16737,N_16605);
nor U16986 (N_16986,N_16614,N_16727);
nor U16987 (N_16987,N_16742,N_16745);
xnor U16988 (N_16988,N_16749,N_16667);
nor U16989 (N_16989,N_16628,N_16773);
nand U16990 (N_16990,N_16787,N_16703);
or U16991 (N_16991,N_16750,N_16639);
or U16992 (N_16992,N_16731,N_16774);
nand U16993 (N_16993,N_16773,N_16784);
nor U16994 (N_16994,N_16664,N_16620);
nor U16995 (N_16995,N_16780,N_16769);
xor U16996 (N_16996,N_16713,N_16714);
nor U16997 (N_16997,N_16694,N_16759);
xnor U16998 (N_16998,N_16765,N_16679);
and U16999 (N_16999,N_16601,N_16724);
or U17000 (N_17000,N_16897,N_16801);
or U17001 (N_17001,N_16853,N_16888);
nand U17002 (N_17002,N_16970,N_16951);
nor U17003 (N_17003,N_16894,N_16930);
nor U17004 (N_17004,N_16993,N_16833);
nand U17005 (N_17005,N_16845,N_16906);
nand U17006 (N_17006,N_16882,N_16928);
and U17007 (N_17007,N_16898,N_16890);
nand U17008 (N_17008,N_16839,N_16827);
and U17009 (N_17009,N_16844,N_16875);
nor U17010 (N_17010,N_16931,N_16869);
or U17011 (N_17011,N_16901,N_16848);
xor U17012 (N_17012,N_16988,N_16958);
or U17013 (N_17013,N_16900,N_16960);
or U17014 (N_17014,N_16999,N_16914);
nor U17015 (N_17015,N_16824,N_16977);
nor U17016 (N_17016,N_16813,N_16817);
or U17017 (N_17017,N_16852,N_16926);
xnor U17018 (N_17018,N_16902,N_16811);
and U17019 (N_17019,N_16805,N_16866);
or U17020 (N_17020,N_16837,N_16807);
nor U17021 (N_17021,N_16870,N_16963);
nand U17022 (N_17022,N_16818,N_16985);
and U17023 (N_17023,N_16821,N_16909);
xnor U17024 (N_17024,N_16995,N_16978);
xor U17025 (N_17025,N_16893,N_16877);
nand U17026 (N_17026,N_16983,N_16940);
or U17027 (N_17027,N_16861,N_16980);
nor U17028 (N_17028,N_16952,N_16874);
and U17029 (N_17029,N_16913,N_16990);
xnor U17030 (N_17030,N_16810,N_16871);
xor U17031 (N_17031,N_16966,N_16804);
and U17032 (N_17032,N_16984,N_16962);
xnor U17033 (N_17033,N_16904,N_16922);
nor U17034 (N_17034,N_16806,N_16856);
and U17035 (N_17035,N_16889,N_16864);
nor U17036 (N_17036,N_16907,N_16994);
or U17037 (N_17037,N_16920,N_16800);
or U17038 (N_17038,N_16903,N_16849);
or U17039 (N_17039,N_16857,N_16938);
or U17040 (N_17040,N_16973,N_16905);
nand U17041 (N_17041,N_16921,N_16934);
and U17042 (N_17042,N_16974,N_16803);
and U17043 (N_17043,N_16885,N_16823);
or U17044 (N_17044,N_16825,N_16954);
and U17045 (N_17045,N_16808,N_16965);
nand U17046 (N_17046,N_16826,N_16935);
and U17047 (N_17047,N_16834,N_16955);
xnor U17048 (N_17048,N_16918,N_16891);
xnor U17049 (N_17049,N_16986,N_16989);
nand U17050 (N_17050,N_16956,N_16937);
nand U17051 (N_17051,N_16859,N_16911);
nor U17052 (N_17052,N_16863,N_16923);
or U17053 (N_17053,N_16860,N_16941);
xnor U17054 (N_17054,N_16814,N_16868);
nor U17055 (N_17055,N_16987,N_16899);
nor U17056 (N_17056,N_16933,N_16841);
nand U17057 (N_17057,N_16915,N_16981);
xor U17058 (N_17058,N_16831,N_16846);
and U17059 (N_17059,N_16946,N_16816);
or U17060 (N_17060,N_16982,N_16924);
xor U17061 (N_17061,N_16892,N_16847);
nand U17062 (N_17062,N_16881,N_16832);
nand U17063 (N_17063,N_16997,N_16916);
or U17064 (N_17064,N_16815,N_16925);
xnor U17065 (N_17065,N_16820,N_16876);
and U17066 (N_17066,N_16880,N_16991);
nor U17067 (N_17067,N_16842,N_16838);
and U17068 (N_17068,N_16959,N_16828);
or U17069 (N_17069,N_16979,N_16975);
xor U17070 (N_17070,N_16961,N_16957);
nand U17071 (N_17071,N_16865,N_16953);
nor U17072 (N_17072,N_16919,N_16992);
or U17073 (N_17073,N_16878,N_16887);
nand U17074 (N_17074,N_16829,N_16917);
nor U17075 (N_17075,N_16939,N_16929);
and U17076 (N_17076,N_16886,N_16969);
and U17077 (N_17077,N_16858,N_16950);
or U17078 (N_17078,N_16884,N_16872);
xnor U17079 (N_17079,N_16843,N_16867);
nand U17080 (N_17080,N_16972,N_16895);
and U17081 (N_17081,N_16836,N_16947);
or U17082 (N_17082,N_16840,N_16927);
nand U17083 (N_17083,N_16809,N_16910);
nand U17084 (N_17084,N_16976,N_16851);
or U17085 (N_17085,N_16971,N_16862);
nand U17086 (N_17086,N_16822,N_16948);
xor U17087 (N_17087,N_16998,N_16855);
nor U17088 (N_17088,N_16996,N_16873);
xnor U17089 (N_17089,N_16964,N_16944);
and U17090 (N_17090,N_16850,N_16819);
or U17091 (N_17091,N_16854,N_16967);
nand U17092 (N_17092,N_16883,N_16879);
or U17093 (N_17093,N_16945,N_16896);
nor U17094 (N_17094,N_16912,N_16835);
xnor U17095 (N_17095,N_16942,N_16943);
and U17096 (N_17096,N_16812,N_16968);
or U17097 (N_17097,N_16802,N_16949);
xor U17098 (N_17098,N_16932,N_16936);
or U17099 (N_17099,N_16908,N_16830);
nand U17100 (N_17100,N_16820,N_16856);
nor U17101 (N_17101,N_16819,N_16828);
nand U17102 (N_17102,N_16807,N_16806);
xor U17103 (N_17103,N_16840,N_16936);
or U17104 (N_17104,N_16971,N_16939);
and U17105 (N_17105,N_16994,N_16872);
nor U17106 (N_17106,N_16983,N_16987);
nor U17107 (N_17107,N_16906,N_16901);
xnor U17108 (N_17108,N_16801,N_16841);
nor U17109 (N_17109,N_16834,N_16979);
or U17110 (N_17110,N_16919,N_16822);
nand U17111 (N_17111,N_16838,N_16833);
xor U17112 (N_17112,N_16882,N_16813);
xnor U17113 (N_17113,N_16935,N_16932);
xnor U17114 (N_17114,N_16893,N_16914);
xnor U17115 (N_17115,N_16911,N_16839);
xor U17116 (N_17116,N_16811,N_16926);
nor U17117 (N_17117,N_16982,N_16978);
or U17118 (N_17118,N_16896,N_16964);
and U17119 (N_17119,N_16856,N_16975);
or U17120 (N_17120,N_16883,N_16988);
and U17121 (N_17121,N_16810,N_16881);
nand U17122 (N_17122,N_16827,N_16867);
or U17123 (N_17123,N_16946,N_16848);
and U17124 (N_17124,N_16871,N_16863);
nand U17125 (N_17125,N_16916,N_16893);
or U17126 (N_17126,N_16842,N_16888);
or U17127 (N_17127,N_16882,N_16805);
or U17128 (N_17128,N_16899,N_16992);
nor U17129 (N_17129,N_16921,N_16833);
xor U17130 (N_17130,N_16963,N_16879);
nor U17131 (N_17131,N_16863,N_16891);
nor U17132 (N_17132,N_16863,N_16921);
xnor U17133 (N_17133,N_16840,N_16871);
nor U17134 (N_17134,N_16882,N_16895);
nor U17135 (N_17135,N_16878,N_16845);
nand U17136 (N_17136,N_16928,N_16805);
xnor U17137 (N_17137,N_16945,N_16803);
nor U17138 (N_17138,N_16868,N_16925);
and U17139 (N_17139,N_16969,N_16966);
nand U17140 (N_17140,N_16891,N_16875);
nand U17141 (N_17141,N_16808,N_16927);
xor U17142 (N_17142,N_16956,N_16823);
xnor U17143 (N_17143,N_16964,N_16887);
nand U17144 (N_17144,N_16933,N_16833);
and U17145 (N_17145,N_16994,N_16877);
xnor U17146 (N_17146,N_16991,N_16872);
or U17147 (N_17147,N_16953,N_16874);
nand U17148 (N_17148,N_16827,N_16920);
and U17149 (N_17149,N_16943,N_16816);
nor U17150 (N_17150,N_16992,N_16867);
or U17151 (N_17151,N_16847,N_16890);
or U17152 (N_17152,N_16934,N_16813);
nor U17153 (N_17153,N_16938,N_16812);
nor U17154 (N_17154,N_16872,N_16948);
nor U17155 (N_17155,N_16811,N_16845);
xor U17156 (N_17156,N_16957,N_16833);
nand U17157 (N_17157,N_16864,N_16962);
nor U17158 (N_17158,N_16868,N_16844);
nand U17159 (N_17159,N_16860,N_16980);
nand U17160 (N_17160,N_16949,N_16824);
xor U17161 (N_17161,N_16842,N_16859);
xor U17162 (N_17162,N_16903,N_16993);
xnor U17163 (N_17163,N_16890,N_16929);
and U17164 (N_17164,N_16818,N_16923);
xor U17165 (N_17165,N_16958,N_16836);
and U17166 (N_17166,N_16892,N_16920);
and U17167 (N_17167,N_16836,N_16898);
xnor U17168 (N_17168,N_16852,N_16939);
or U17169 (N_17169,N_16884,N_16915);
nand U17170 (N_17170,N_16854,N_16809);
xor U17171 (N_17171,N_16835,N_16906);
or U17172 (N_17172,N_16888,N_16895);
nand U17173 (N_17173,N_16923,N_16982);
nor U17174 (N_17174,N_16840,N_16868);
or U17175 (N_17175,N_16816,N_16937);
or U17176 (N_17176,N_16839,N_16939);
or U17177 (N_17177,N_16874,N_16880);
or U17178 (N_17178,N_16825,N_16984);
and U17179 (N_17179,N_16957,N_16980);
or U17180 (N_17180,N_16996,N_16952);
nor U17181 (N_17181,N_16938,N_16988);
xnor U17182 (N_17182,N_16933,N_16817);
or U17183 (N_17183,N_16948,N_16814);
and U17184 (N_17184,N_16900,N_16856);
and U17185 (N_17185,N_16883,N_16969);
nand U17186 (N_17186,N_16896,N_16841);
and U17187 (N_17187,N_16931,N_16875);
or U17188 (N_17188,N_16926,N_16923);
nand U17189 (N_17189,N_16890,N_16959);
or U17190 (N_17190,N_16849,N_16951);
and U17191 (N_17191,N_16967,N_16952);
nor U17192 (N_17192,N_16814,N_16823);
or U17193 (N_17193,N_16918,N_16846);
nand U17194 (N_17194,N_16895,N_16971);
and U17195 (N_17195,N_16869,N_16920);
nand U17196 (N_17196,N_16971,N_16833);
nand U17197 (N_17197,N_16835,N_16970);
or U17198 (N_17198,N_16933,N_16877);
nor U17199 (N_17199,N_16961,N_16825);
nor U17200 (N_17200,N_17022,N_17063);
and U17201 (N_17201,N_17042,N_17127);
xnor U17202 (N_17202,N_17006,N_17033);
and U17203 (N_17203,N_17057,N_17090);
nand U17204 (N_17204,N_17171,N_17140);
nor U17205 (N_17205,N_17094,N_17038);
nand U17206 (N_17206,N_17186,N_17051);
nand U17207 (N_17207,N_17052,N_17074);
xor U17208 (N_17208,N_17112,N_17153);
nand U17209 (N_17209,N_17134,N_17172);
or U17210 (N_17210,N_17187,N_17149);
nor U17211 (N_17211,N_17174,N_17141);
xnor U17212 (N_17212,N_17159,N_17080);
xnor U17213 (N_17213,N_17079,N_17078);
nor U17214 (N_17214,N_17059,N_17055);
nor U17215 (N_17215,N_17076,N_17054);
and U17216 (N_17216,N_17124,N_17101);
and U17217 (N_17217,N_17144,N_17178);
nand U17218 (N_17218,N_17156,N_17026);
or U17219 (N_17219,N_17177,N_17087);
and U17220 (N_17220,N_17182,N_17043);
and U17221 (N_17221,N_17049,N_17196);
or U17222 (N_17222,N_17130,N_17040);
and U17223 (N_17223,N_17041,N_17192);
and U17224 (N_17224,N_17065,N_17106);
nand U17225 (N_17225,N_17166,N_17167);
nand U17226 (N_17226,N_17120,N_17082);
and U17227 (N_17227,N_17136,N_17012);
xnor U17228 (N_17228,N_17143,N_17176);
nor U17229 (N_17229,N_17035,N_17058);
or U17230 (N_17230,N_17173,N_17077);
nand U17231 (N_17231,N_17137,N_17021);
or U17232 (N_17232,N_17095,N_17123);
xor U17233 (N_17233,N_17142,N_17061);
nand U17234 (N_17234,N_17111,N_17110);
xnor U17235 (N_17235,N_17066,N_17088);
nand U17236 (N_17236,N_17083,N_17016);
or U17237 (N_17237,N_17104,N_17183);
nor U17238 (N_17238,N_17064,N_17185);
nor U17239 (N_17239,N_17036,N_17010);
nor U17240 (N_17240,N_17170,N_17070);
and U17241 (N_17241,N_17086,N_17019);
nor U17242 (N_17242,N_17004,N_17007);
or U17243 (N_17243,N_17068,N_17030);
and U17244 (N_17244,N_17138,N_17188);
nor U17245 (N_17245,N_17168,N_17018);
nor U17246 (N_17246,N_17028,N_17005);
nor U17247 (N_17247,N_17089,N_17114);
xor U17248 (N_17248,N_17152,N_17072);
xor U17249 (N_17249,N_17103,N_17027);
xor U17250 (N_17250,N_17069,N_17048);
and U17251 (N_17251,N_17118,N_17133);
or U17252 (N_17252,N_17148,N_17116);
xor U17253 (N_17253,N_17017,N_17175);
or U17254 (N_17254,N_17093,N_17097);
xnor U17255 (N_17255,N_17034,N_17025);
nor U17256 (N_17256,N_17013,N_17160);
nor U17257 (N_17257,N_17115,N_17084);
and U17258 (N_17258,N_17009,N_17139);
or U17259 (N_17259,N_17107,N_17045);
xnor U17260 (N_17260,N_17117,N_17102);
and U17261 (N_17261,N_17191,N_17169);
or U17262 (N_17262,N_17125,N_17121);
xor U17263 (N_17263,N_17031,N_17197);
xnor U17264 (N_17264,N_17008,N_17047);
or U17265 (N_17265,N_17091,N_17000);
nand U17266 (N_17266,N_17128,N_17014);
nand U17267 (N_17267,N_17085,N_17155);
nand U17268 (N_17268,N_17195,N_17062);
and U17269 (N_17269,N_17193,N_17180);
xor U17270 (N_17270,N_17029,N_17067);
nor U17271 (N_17271,N_17151,N_17164);
and U17272 (N_17272,N_17092,N_17131);
nor U17273 (N_17273,N_17179,N_17161);
nor U17274 (N_17274,N_17060,N_17020);
xnor U17275 (N_17275,N_17126,N_17075);
or U17276 (N_17276,N_17135,N_17184);
nor U17277 (N_17277,N_17129,N_17100);
nor U17278 (N_17278,N_17150,N_17099);
xor U17279 (N_17279,N_17157,N_17044);
nor U17280 (N_17280,N_17113,N_17181);
and U17281 (N_17281,N_17015,N_17109);
and U17282 (N_17282,N_17037,N_17096);
or U17283 (N_17283,N_17073,N_17198);
nand U17284 (N_17284,N_17163,N_17199);
nor U17285 (N_17285,N_17053,N_17002);
nor U17286 (N_17286,N_17122,N_17108);
nor U17287 (N_17287,N_17132,N_17190);
and U17288 (N_17288,N_17194,N_17162);
or U17289 (N_17289,N_17003,N_17032);
and U17290 (N_17290,N_17154,N_17046);
and U17291 (N_17291,N_17146,N_17119);
nand U17292 (N_17292,N_17081,N_17158);
or U17293 (N_17293,N_17145,N_17071);
and U17294 (N_17294,N_17039,N_17165);
nor U17295 (N_17295,N_17024,N_17001);
xnor U17296 (N_17296,N_17147,N_17011);
xor U17297 (N_17297,N_17098,N_17056);
nor U17298 (N_17298,N_17189,N_17105);
or U17299 (N_17299,N_17050,N_17023);
or U17300 (N_17300,N_17176,N_17118);
and U17301 (N_17301,N_17133,N_17125);
or U17302 (N_17302,N_17056,N_17003);
or U17303 (N_17303,N_17165,N_17187);
xnor U17304 (N_17304,N_17117,N_17156);
xnor U17305 (N_17305,N_17071,N_17181);
nor U17306 (N_17306,N_17010,N_17199);
or U17307 (N_17307,N_17099,N_17139);
and U17308 (N_17308,N_17148,N_17093);
xor U17309 (N_17309,N_17141,N_17136);
nor U17310 (N_17310,N_17031,N_17157);
or U17311 (N_17311,N_17096,N_17188);
or U17312 (N_17312,N_17195,N_17117);
nor U17313 (N_17313,N_17195,N_17097);
xnor U17314 (N_17314,N_17073,N_17098);
xnor U17315 (N_17315,N_17084,N_17028);
nor U17316 (N_17316,N_17041,N_17096);
nor U17317 (N_17317,N_17123,N_17025);
xnor U17318 (N_17318,N_17032,N_17122);
xor U17319 (N_17319,N_17175,N_17041);
and U17320 (N_17320,N_17091,N_17069);
nor U17321 (N_17321,N_17048,N_17172);
and U17322 (N_17322,N_17019,N_17024);
nand U17323 (N_17323,N_17195,N_17054);
or U17324 (N_17324,N_17036,N_17143);
xnor U17325 (N_17325,N_17066,N_17022);
xnor U17326 (N_17326,N_17020,N_17052);
nand U17327 (N_17327,N_17007,N_17038);
nor U17328 (N_17328,N_17087,N_17143);
xnor U17329 (N_17329,N_17132,N_17153);
nand U17330 (N_17330,N_17121,N_17102);
or U17331 (N_17331,N_17147,N_17007);
or U17332 (N_17332,N_17136,N_17128);
nand U17333 (N_17333,N_17008,N_17145);
and U17334 (N_17334,N_17018,N_17078);
nand U17335 (N_17335,N_17190,N_17155);
nand U17336 (N_17336,N_17019,N_17115);
xor U17337 (N_17337,N_17074,N_17043);
nand U17338 (N_17338,N_17198,N_17087);
xor U17339 (N_17339,N_17098,N_17024);
nor U17340 (N_17340,N_17166,N_17113);
nor U17341 (N_17341,N_17100,N_17135);
xnor U17342 (N_17342,N_17011,N_17071);
nand U17343 (N_17343,N_17170,N_17131);
xor U17344 (N_17344,N_17155,N_17102);
nand U17345 (N_17345,N_17133,N_17097);
or U17346 (N_17346,N_17169,N_17170);
and U17347 (N_17347,N_17158,N_17079);
or U17348 (N_17348,N_17135,N_17161);
nand U17349 (N_17349,N_17164,N_17040);
nor U17350 (N_17350,N_17054,N_17071);
nand U17351 (N_17351,N_17042,N_17015);
nand U17352 (N_17352,N_17195,N_17183);
nand U17353 (N_17353,N_17049,N_17170);
nand U17354 (N_17354,N_17028,N_17179);
and U17355 (N_17355,N_17134,N_17033);
nand U17356 (N_17356,N_17046,N_17152);
xor U17357 (N_17357,N_17145,N_17053);
and U17358 (N_17358,N_17132,N_17044);
or U17359 (N_17359,N_17154,N_17148);
or U17360 (N_17360,N_17058,N_17000);
nor U17361 (N_17361,N_17081,N_17058);
nor U17362 (N_17362,N_17126,N_17053);
nand U17363 (N_17363,N_17176,N_17172);
and U17364 (N_17364,N_17199,N_17136);
xor U17365 (N_17365,N_17038,N_17196);
nand U17366 (N_17366,N_17155,N_17169);
and U17367 (N_17367,N_17163,N_17049);
nor U17368 (N_17368,N_17050,N_17029);
and U17369 (N_17369,N_17119,N_17130);
nand U17370 (N_17370,N_17020,N_17065);
nor U17371 (N_17371,N_17090,N_17175);
and U17372 (N_17372,N_17188,N_17091);
nor U17373 (N_17373,N_17189,N_17188);
or U17374 (N_17374,N_17099,N_17085);
xor U17375 (N_17375,N_17104,N_17199);
nor U17376 (N_17376,N_17118,N_17107);
nand U17377 (N_17377,N_17104,N_17151);
nor U17378 (N_17378,N_17027,N_17090);
and U17379 (N_17379,N_17028,N_17023);
nor U17380 (N_17380,N_17063,N_17100);
nor U17381 (N_17381,N_17102,N_17144);
nand U17382 (N_17382,N_17005,N_17167);
or U17383 (N_17383,N_17141,N_17120);
xor U17384 (N_17384,N_17033,N_17035);
nor U17385 (N_17385,N_17179,N_17117);
nand U17386 (N_17386,N_17055,N_17047);
xnor U17387 (N_17387,N_17062,N_17171);
xnor U17388 (N_17388,N_17037,N_17147);
and U17389 (N_17389,N_17008,N_17035);
and U17390 (N_17390,N_17080,N_17182);
nor U17391 (N_17391,N_17152,N_17156);
nand U17392 (N_17392,N_17076,N_17056);
nand U17393 (N_17393,N_17021,N_17106);
and U17394 (N_17394,N_17181,N_17013);
or U17395 (N_17395,N_17064,N_17017);
nor U17396 (N_17396,N_17126,N_17138);
and U17397 (N_17397,N_17118,N_17095);
or U17398 (N_17398,N_17124,N_17187);
and U17399 (N_17399,N_17045,N_17194);
and U17400 (N_17400,N_17336,N_17203);
or U17401 (N_17401,N_17208,N_17379);
or U17402 (N_17402,N_17325,N_17353);
nor U17403 (N_17403,N_17289,N_17321);
or U17404 (N_17404,N_17307,N_17284);
nor U17405 (N_17405,N_17395,N_17250);
or U17406 (N_17406,N_17339,N_17391);
nand U17407 (N_17407,N_17311,N_17270);
nor U17408 (N_17408,N_17310,N_17285);
xnor U17409 (N_17409,N_17388,N_17207);
or U17410 (N_17410,N_17381,N_17322);
nor U17411 (N_17411,N_17282,N_17300);
or U17412 (N_17412,N_17362,N_17387);
or U17413 (N_17413,N_17314,N_17241);
and U17414 (N_17414,N_17224,N_17398);
nand U17415 (N_17415,N_17291,N_17371);
nor U17416 (N_17416,N_17305,N_17326);
or U17417 (N_17417,N_17374,N_17292);
and U17418 (N_17418,N_17301,N_17239);
nor U17419 (N_17419,N_17397,N_17227);
and U17420 (N_17420,N_17271,N_17363);
and U17421 (N_17421,N_17378,N_17373);
and U17422 (N_17422,N_17308,N_17390);
nand U17423 (N_17423,N_17313,N_17380);
nor U17424 (N_17424,N_17204,N_17280);
or U17425 (N_17425,N_17389,N_17244);
xor U17426 (N_17426,N_17396,N_17214);
nor U17427 (N_17427,N_17294,N_17201);
nor U17428 (N_17428,N_17357,N_17318);
nor U17429 (N_17429,N_17399,N_17315);
nand U17430 (N_17430,N_17283,N_17333);
and U17431 (N_17431,N_17320,N_17365);
xor U17432 (N_17432,N_17354,N_17229);
or U17433 (N_17433,N_17202,N_17332);
nand U17434 (N_17434,N_17223,N_17225);
nand U17435 (N_17435,N_17238,N_17236);
nand U17436 (N_17436,N_17264,N_17200);
nand U17437 (N_17437,N_17242,N_17359);
nand U17438 (N_17438,N_17298,N_17377);
xor U17439 (N_17439,N_17222,N_17232);
xor U17440 (N_17440,N_17327,N_17205);
or U17441 (N_17441,N_17376,N_17209);
xor U17442 (N_17442,N_17274,N_17356);
nand U17443 (N_17443,N_17275,N_17216);
nand U17444 (N_17444,N_17266,N_17392);
or U17445 (N_17445,N_17256,N_17361);
nor U17446 (N_17446,N_17290,N_17394);
and U17447 (N_17447,N_17324,N_17375);
nor U17448 (N_17448,N_17263,N_17257);
nor U17449 (N_17449,N_17258,N_17323);
and U17450 (N_17450,N_17329,N_17364);
or U17451 (N_17451,N_17243,N_17296);
xnor U17452 (N_17452,N_17338,N_17249);
or U17453 (N_17453,N_17267,N_17383);
nor U17454 (N_17454,N_17293,N_17386);
or U17455 (N_17455,N_17279,N_17348);
and U17456 (N_17456,N_17215,N_17355);
nor U17457 (N_17457,N_17342,N_17385);
or U17458 (N_17458,N_17273,N_17233);
or U17459 (N_17459,N_17299,N_17262);
nor U17460 (N_17460,N_17316,N_17228);
nand U17461 (N_17461,N_17295,N_17220);
nor U17462 (N_17462,N_17345,N_17245);
and U17463 (N_17463,N_17328,N_17281);
or U17464 (N_17464,N_17303,N_17234);
or U17465 (N_17465,N_17360,N_17272);
nor U17466 (N_17466,N_17340,N_17370);
or U17467 (N_17467,N_17297,N_17287);
xnor U17468 (N_17468,N_17247,N_17212);
nor U17469 (N_17469,N_17358,N_17335);
nand U17470 (N_17470,N_17350,N_17278);
xor U17471 (N_17471,N_17260,N_17251);
nand U17472 (N_17472,N_17211,N_17382);
or U17473 (N_17473,N_17206,N_17237);
nand U17474 (N_17474,N_17366,N_17304);
and U17475 (N_17475,N_17312,N_17240);
and U17476 (N_17476,N_17226,N_17319);
and U17477 (N_17477,N_17255,N_17330);
nand U17478 (N_17478,N_17331,N_17218);
xnor U17479 (N_17479,N_17230,N_17252);
nor U17480 (N_17480,N_17265,N_17346);
xor U17481 (N_17481,N_17372,N_17367);
nor U17482 (N_17482,N_17259,N_17341);
and U17483 (N_17483,N_17231,N_17317);
nor U17484 (N_17484,N_17349,N_17351);
and U17485 (N_17485,N_17253,N_17337);
and U17486 (N_17486,N_17302,N_17369);
xnor U17487 (N_17487,N_17393,N_17235);
nor U17488 (N_17488,N_17254,N_17248);
or U17489 (N_17489,N_17269,N_17276);
xnor U17490 (N_17490,N_17213,N_17210);
or U17491 (N_17491,N_17261,N_17268);
nand U17492 (N_17492,N_17384,N_17347);
and U17493 (N_17493,N_17352,N_17344);
nor U17494 (N_17494,N_17219,N_17288);
nor U17495 (N_17495,N_17306,N_17368);
xnor U17496 (N_17496,N_17246,N_17343);
xnor U17497 (N_17497,N_17334,N_17217);
nor U17498 (N_17498,N_17286,N_17277);
xnor U17499 (N_17499,N_17309,N_17221);
xor U17500 (N_17500,N_17228,N_17257);
or U17501 (N_17501,N_17277,N_17366);
nor U17502 (N_17502,N_17220,N_17360);
or U17503 (N_17503,N_17297,N_17277);
and U17504 (N_17504,N_17222,N_17298);
xor U17505 (N_17505,N_17385,N_17357);
xor U17506 (N_17506,N_17387,N_17371);
and U17507 (N_17507,N_17262,N_17225);
nand U17508 (N_17508,N_17397,N_17236);
nor U17509 (N_17509,N_17348,N_17344);
xnor U17510 (N_17510,N_17354,N_17293);
and U17511 (N_17511,N_17333,N_17316);
xnor U17512 (N_17512,N_17269,N_17202);
nand U17513 (N_17513,N_17326,N_17373);
nand U17514 (N_17514,N_17234,N_17285);
and U17515 (N_17515,N_17368,N_17360);
nor U17516 (N_17516,N_17269,N_17384);
or U17517 (N_17517,N_17394,N_17333);
and U17518 (N_17518,N_17245,N_17231);
nor U17519 (N_17519,N_17391,N_17314);
and U17520 (N_17520,N_17399,N_17235);
and U17521 (N_17521,N_17210,N_17386);
and U17522 (N_17522,N_17252,N_17384);
and U17523 (N_17523,N_17355,N_17323);
nand U17524 (N_17524,N_17291,N_17307);
and U17525 (N_17525,N_17346,N_17364);
or U17526 (N_17526,N_17308,N_17288);
and U17527 (N_17527,N_17261,N_17259);
nand U17528 (N_17528,N_17371,N_17297);
nand U17529 (N_17529,N_17235,N_17266);
nand U17530 (N_17530,N_17237,N_17330);
and U17531 (N_17531,N_17343,N_17215);
nand U17532 (N_17532,N_17212,N_17347);
nor U17533 (N_17533,N_17229,N_17327);
and U17534 (N_17534,N_17347,N_17397);
or U17535 (N_17535,N_17258,N_17315);
nand U17536 (N_17536,N_17376,N_17293);
or U17537 (N_17537,N_17212,N_17310);
xnor U17538 (N_17538,N_17251,N_17328);
or U17539 (N_17539,N_17222,N_17379);
xnor U17540 (N_17540,N_17393,N_17232);
and U17541 (N_17541,N_17347,N_17298);
xor U17542 (N_17542,N_17344,N_17364);
xnor U17543 (N_17543,N_17381,N_17240);
or U17544 (N_17544,N_17208,N_17393);
nand U17545 (N_17545,N_17270,N_17317);
nand U17546 (N_17546,N_17266,N_17225);
nand U17547 (N_17547,N_17264,N_17347);
and U17548 (N_17548,N_17277,N_17258);
and U17549 (N_17549,N_17330,N_17379);
xnor U17550 (N_17550,N_17242,N_17231);
and U17551 (N_17551,N_17366,N_17268);
and U17552 (N_17552,N_17269,N_17399);
nor U17553 (N_17553,N_17364,N_17372);
nand U17554 (N_17554,N_17356,N_17268);
nand U17555 (N_17555,N_17347,N_17360);
nand U17556 (N_17556,N_17378,N_17322);
and U17557 (N_17557,N_17299,N_17349);
and U17558 (N_17558,N_17261,N_17349);
xor U17559 (N_17559,N_17285,N_17210);
xnor U17560 (N_17560,N_17395,N_17237);
nor U17561 (N_17561,N_17241,N_17349);
nand U17562 (N_17562,N_17267,N_17241);
nand U17563 (N_17563,N_17239,N_17362);
or U17564 (N_17564,N_17229,N_17331);
xor U17565 (N_17565,N_17301,N_17318);
and U17566 (N_17566,N_17363,N_17249);
nand U17567 (N_17567,N_17376,N_17292);
nor U17568 (N_17568,N_17329,N_17272);
xor U17569 (N_17569,N_17289,N_17214);
xor U17570 (N_17570,N_17326,N_17268);
nand U17571 (N_17571,N_17215,N_17373);
and U17572 (N_17572,N_17352,N_17327);
nor U17573 (N_17573,N_17242,N_17370);
and U17574 (N_17574,N_17217,N_17319);
nor U17575 (N_17575,N_17286,N_17222);
or U17576 (N_17576,N_17322,N_17200);
nand U17577 (N_17577,N_17332,N_17249);
nand U17578 (N_17578,N_17208,N_17236);
nand U17579 (N_17579,N_17332,N_17354);
nor U17580 (N_17580,N_17371,N_17374);
or U17581 (N_17581,N_17345,N_17249);
nand U17582 (N_17582,N_17256,N_17359);
nor U17583 (N_17583,N_17360,N_17306);
nand U17584 (N_17584,N_17215,N_17323);
and U17585 (N_17585,N_17288,N_17206);
or U17586 (N_17586,N_17281,N_17255);
xor U17587 (N_17587,N_17361,N_17276);
and U17588 (N_17588,N_17330,N_17376);
and U17589 (N_17589,N_17273,N_17287);
and U17590 (N_17590,N_17266,N_17262);
xor U17591 (N_17591,N_17319,N_17341);
nor U17592 (N_17592,N_17378,N_17281);
nand U17593 (N_17593,N_17225,N_17375);
and U17594 (N_17594,N_17229,N_17350);
nor U17595 (N_17595,N_17301,N_17252);
and U17596 (N_17596,N_17357,N_17270);
xor U17597 (N_17597,N_17385,N_17311);
or U17598 (N_17598,N_17348,N_17205);
xor U17599 (N_17599,N_17392,N_17377);
xnor U17600 (N_17600,N_17425,N_17423);
nor U17601 (N_17601,N_17469,N_17545);
xor U17602 (N_17602,N_17592,N_17435);
and U17603 (N_17603,N_17552,N_17526);
or U17604 (N_17604,N_17563,N_17447);
nor U17605 (N_17605,N_17465,N_17557);
and U17606 (N_17606,N_17427,N_17582);
nand U17607 (N_17607,N_17504,N_17599);
or U17608 (N_17608,N_17416,N_17574);
nand U17609 (N_17609,N_17419,N_17551);
and U17610 (N_17610,N_17512,N_17494);
nor U17611 (N_17611,N_17430,N_17481);
nor U17612 (N_17612,N_17542,N_17418);
and U17613 (N_17613,N_17451,N_17410);
or U17614 (N_17614,N_17426,N_17495);
or U17615 (N_17615,N_17468,N_17517);
nor U17616 (N_17616,N_17450,N_17490);
and U17617 (N_17617,N_17420,N_17522);
nand U17618 (N_17618,N_17521,N_17562);
or U17619 (N_17619,N_17500,N_17487);
nand U17620 (N_17620,N_17421,N_17409);
nand U17621 (N_17621,N_17444,N_17520);
nor U17622 (N_17622,N_17580,N_17448);
and U17623 (N_17623,N_17530,N_17493);
or U17624 (N_17624,N_17525,N_17588);
or U17625 (N_17625,N_17422,N_17483);
nor U17626 (N_17626,N_17445,N_17463);
and U17627 (N_17627,N_17598,N_17453);
or U17628 (N_17628,N_17477,N_17591);
or U17629 (N_17629,N_17498,N_17597);
xnor U17630 (N_17630,N_17514,N_17533);
nor U17631 (N_17631,N_17449,N_17476);
nand U17632 (N_17632,N_17524,N_17559);
nor U17633 (N_17633,N_17475,N_17497);
xor U17634 (N_17634,N_17527,N_17470);
nand U17635 (N_17635,N_17415,N_17540);
or U17636 (N_17636,N_17529,N_17446);
nor U17637 (N_17637,N_17431,N_17489);
nand U17638 (N_17638,N_17414,N_17561);
and U17639 (N_17639,N_17596,N_17471);
xnor U17640 (N_17640,N_17429,N_17515);
xor U17641 (N_17641,N_17488,N_17438);
and U17642 (N_17642,N_17452,N_17464);
or U17643 (N_17643,N_17546,N_17523);
nand U17644 (N_17644,N_17560,N_17543);
nand U17645 (N_17645,N_17442,N_17575);
or U17646 (N_17646,N_17456,N_17455);
nand U17647 (N_17647,N_17434,N_17405);
nor U17648 (N_17648,N_17459,N_17579);
and U17649 (N_17649,N_17467,N_17486);
and U17650 (N_17650,N_17538,N_17554);
xnor U17651 (N_17651,N_17516,N_17432);
or U17652 (N_17652,N_17403,N_17590);
or U17653 (N_17653,N_17458,N_17581);
nor U17654 (N_17654,N_17466,N_17576);
or U17655 (N_17655,N_17539,N_17553);
or U17656 (N_17656,N_17411,N_17479);
xor U17657 (N_17657,N_17535,N_17491);
or U17658 (N_17658,N_17485,N_17555);
and U17659 (N_17659,N_17566,N_17564);
xnor U17660 (N_17660,N_17549,N_17482);
nor U17661 (N_17661,N_17472,N_17457);
nand U17662 (N_17662,N_17462,N_17583);
xnor U17663 (N_17663,N_17528,N_17428);
xnor U17664 (N_17664,N_17417,N_17473);
nand U17665 (N_17665,N_17508,N_17503);
xnor U17666 (N_17666,N_17499,N_17502);
and U17667 (N_17667,N_17400,N_17439);
nor U17668 (N_17668,N_17407,N_17461);
xnor U17669 (N_17669,N_17454,N_17547);
nand U17670 (N_17670,N_17507,N_17505);
nand U17671 (N_17671,N_17511,N_17437);
xnor U17672 (N_17672,N_17584,N_17565);
nor U17673 (N_17673,N_17593,N_17406);
or U17674 (N_17674,N_17550,N_17402);
nor U17675 (N_17675,N_17509,N_17587);
nor U17676 (N_17676,N_17424,N_17460);
nand U17677 (N_17677,N_17440,N_17401);
and U17678 (N_17678,N_17501,N_17518);
nand U17679 (N_17679,N_17578,N_17513);
nor U17680 (N_17680,N_17408,N_17443);
and U17681 (N_17681,N_17492,N_17571);
xnor U17682 (N_17682,N_17436,N_17537);
or U17683 (N_17683,N_17506,N_17484);
and U17684 (N_17684,N_17572,N_17570);
nor U17685 (N_17685,N_17474,N_17510);
xor U17686 (N_17686,N_17412,N_17433);
nand U17687 (N_17687,N_17594,N_17544);
nor U17688 (N_17688,N_17589,N_17534);
or U17689 (N_17689,N_17531,N_17536);
nor U17690 (N_17690,N_17532,N_17541);
nand U17691 (N_17691,N_17478,N_17573);
xnor U17692 (N_17692,N_17441,N_17568);
xnor U17693 (N_17693,N_17413,N_17548);
and U17694 (N_17694,N_17480,N_17519);
nor U17695 (N_17695,N_17558,N_17556);
xnor U17696 (N_17696,N_17585,N_17595);
and U17697 (N_17697,N_17586,N_17567);
nor U17698 (N_17698,N_17404,N_17569);
xnor U17699 (N_17699,N_17496,N_17577);
xnor U17700 (N_17700,N_17506,N_17565);
xor U17701 (N_17701,N_17527,N_17492);
or U17702 (N_17702,N_17504,N_17431);
or U17703 (N_17703,N_17428,N_17429);
and U17704 (N_17704,N_17513,N_17403);
nor U17705 (N_17705,N_17569,N_17485);
xnor U17706 (N_17706,N_17575,N_17505);
nor U17707 (N_17707,N_17473,N_17468);
nor U17708 (N_17708,N_17461,N_17532);
or U17709 (N_17709,N_17426,N_17492);
xnor U17710 (N_17710,N_17444,N_17407);
or U17711 (N_17711,N_17590,N_17518);
xnor U17712 (N_17712,N_17591,N_17520);
and U17713 (N_17713,N_17453,N_17476);
xnor U17714 (N_17714,N_17569,N_17516);
nor U17715 (N_17715,N_17488,N_17457);
or U17716 (N_17716,N_17589,N_17586);
nor U17717 (N_17717,N_17510,N_17505);
and U17718 (N_17718,N_17513,N_17588);
nor U17719 (N_17719,N_17408,N_17583);
nand U17720 (N_17720,N_17519,N_17432);
and U17721 (N_17721,N_17529,N_17482);
nor U17722 (N_17722,N_17596,N_17435);
xor U17723 (N_17723,N_17509,N_17550);
or U17724 (N_17724,N_17598,N_17479);
and U17725 (N_17725,N_17406,N_17466);
xnor U17726 (N_17726,N_17553,N_17513);
or U17727 (N_17727,N_17473,N_17586);
nand U17728 (N_17728,N_17559,N_17534);
xor U17729 (N_17729,N_17564,N_17495);
or U17730 (N_17730,N_17500,N_17586);
nor U17731 (N_17731,N_17555,N_17464);
nor U17732 (N_17732,N_17522,N_17575);
nor U17733 (N_17733,N_17558,N_17435);
xnor U17734 (N_17734,N_17555,N_17583);
nand U17735 (N_17735,N_17534,N_17449);
nand U17736 (N_17736,N_17446,N_17452);
nor U17737 (N_17737,N_17553,N_17511);
xor U17738 (N_17738,N_17472,N_17517);
nor U17739 (N_17739,N_17506,N_17554);
xor U17740 (N_17740,N_17560,N_17576);
nand U17741 (N_17741,N_17555,N_17542);
and U17742 (N_17742,N_17444,N_17589);
nor U17743 (N_17743,N_17430,N_17564);
and U17744 (N_17744,N_17488,N_17510);
nor U17745 (N_17745,N_17572,N_17565);
nand U17746 (N_17746,N_17492,N_17511);
nor U17747 (N_17747,N_17494,N_17495);
nor U17748 (N_17748,N_17422,N_17597);
or U17749 (N_17749,N_17523,N_17501);
or U17750 (N_17750,N_17467,N_17474);
nor U17751 (N_17751,N_17453,N_17409);
and U17752 (N_17752,N_17447,N_17457);
xnor U17753 (N_17753,N_17494,N_17565);
or U17754 (N_17754,N_17590,N_17572);
and U17755 (N_17755,N_17496,N_17473);
nor U17756 (N_17756,N_17504,N_17426);
or U17757 (N_17757,N_17575,N_17446);
xnor U17758 (N_17758,N_17448,N_17470);
xor U17759 (N_17759,N_17539,N_17526);
or U17760 (N_17760,N_17552,N_17478);
or U17761 (N_17761,N_17424,N_17509);
and U17762 (N_17762,N_17570,N_17463);
nand U17763 (N_17763,N_17557,N_17582);
nor U17764 (N_17764,N_17496,N_17451);
nand U17765 (N_17765,N_17486,N_17574);
or U17766 (N_17766,N_17520,N_17484);
nand U17767 (N_17767,N_17585,N_17454);
xnor U17768 (N_17768,N_17552,N_17544);
or U17769 (N_17769,N_17485,N_17406);
nor U17770 (N_17770,N_17524,N_17537);
or U17771 (N_17771,N_17567,N_17496);
and U17772 (N_17772,N_17543,N_17541);
or U17773 (N_17773,N_17498,N_17559);
xor U17774 (N_17774,N_17498,N_17505);
or U17775 (N_17775,N_17444,N_17506);
nor U17776 (N_17776,N_17541,N_17594);
xor U17777 (N_17777,N_17473,N_17530);
nand U17778 (N_17778,N_17490,N_17409);
or U17779 (N_17779,N_17525,N_17511);
or U17780 (N_17780,N_17532,N_17477);
nor U17781 (N_17781,N_17510,N_17517);
xor U17782 (N_17782,N_17591,N_17434);
or U17783 (N_17783,N_17533,N_17442);
nor U17784 (N_17784,N_17424,N_17459);
xnor U17785 (N_17785,N_17458,N_17498);
nor U17786 (N_17786,N_17485,N_17499);
xnor U17787 (N_17787,N_17445,N_17593);
or U17788 (N_17788,N_17522,N_17412);
nor U17789 (N_17789,N_17487,N_17585);
nand U17790 (N_17790,N_17437,N_17543);
xnor U17791 (N_17791,N_17567,N_17497);
or U17792 (N_17792,N_17518,N_17583);
or U17793 (N_17793,N_17524,N_17575);
or U17794 (N_17794,N_17474,N_17478);
or U17795 (N_17795,N_17487,N_17481);
xnor U17796 (N_17796,N_17558,N_17504);
nand U17797 (N_17797,N_17558,N_17421);
or U17798 (N_17798,N_17445,N_17446);
and U17799 (N_17799,N_17563,N_17566);
nand U17800 (N_17800,N_17734,N_17794);
nor U17801 (N_17801,N_17781,N_17659);
nor U17802 (N_17802,N_17658,N_17647);
xnor U17803 (N_17803,N_17788,N_17751);
or U17804 (N_17804,N_17614,N_17780);
nand U17805 (N_17805,N_17676,N_17645);
nand U17806 (N_17806,N_17673,N_17782);
xnor U17807 (N_17807,N_17619,N_17705);
nor U17808 (N_17808,N_17696,N_17632);
nand U17809 (N_17809,N_17616,N_17725);
nor U17810 (N_17810,N_17642,N_17654);
or U17811 (N_17811,N_17764,N_17664);
nor U17812 (N_17812,N_17680,N_17748);
or U17813 (N_17813,N_17694,N_17608);
xor U17814 (N_17814,N_17776,N_17739);
or U17815 (N_17815,N_17762,N_17674);
nand U17816 (N_17816,N_17718,N_17760);
and U17817 (N_17817,N_17677,N_17749);
or U17818 (N_17818,N_17672,N_17693);
xnor U17819 (N_17819,N_17766,N_17600);
and U17820 (N_17820,N_17754,N_17629);
and U17821 (N_17821,N_17774,N_17669);
xor U17822 (N_17822,N_17612,N_17628);
and U17823 (N_17823,N_17602,N_17643);
and U17824 (N_17824,N_17688,N_17757);
or U17825 (N_17825,N_17615,N_17714);
xor U17826 (N_17826,N_17796,N_17732);
nand U17827 (N_17827,N_17722,N_17706);
xnor U17828 (N_17828,N_17752,N_17657);
xor U17829 (N_17829,N_17624,N_17667);
nor U17830 (N_17830,N_17661,N_17641);
nor U17831 (N_17831,N_17770,N_17731);
xnor U17832 (N_17832,N_17763,N_17604);
nand U17833 (N_17833,N_17772,N_17735);
nand U17834 (N_17834,N_17791,N_17789);
nand U17835 (N_17835,N_17793,N_17610);
nor U17836 (N_17836,N_17713,N_17700);
xnor U17837 (N_17837,N_17708,N_17753);
nor U17838 (N_17838,N_17797,N_17773);
nand U17839 (N_17839,N_17799,N_17779);
or U17840 (N_17840,N_17698,N_17765);
or U17841 (N_17841,N_17768,N_17778);
nor U17842 (N_17842,N_17792,N_17790);
nor U17843 (N_17843,N_17702,N_17671);
xor U17844 (N_17844,N_17606,N_17704);
xor U17845 (N_17845,N_17717,N_17710);
or U17846 (N_17846,N_17729,N_17775);
and U17847 (N_17847,N_17728,N_17730);
nor U17848 (N_17848,N_17678,N_17670);
and U17849 (N_17849,N_17742,N_17715);
nor U17850 (N_17850,N_17777,N_17611);
or U17851 (N_17851,N_17787,N_17721);
and U17852 (N_17852,N_17648,N_17785);
and U17853 (N_17853,N_17656,N_17724);
nand U17854 (N_17854,N_17607,N_17755);
or U17855 (N_17855,N_17738,N_17625);
xor U17856 (N_17856,N_17783,N_17691);
nand U17857 (N_17857,N_17741,N_17795);
nor U17858 (N_17858,N_17651,N_17746);
nor U17859 (N_17859,N_17621,N_17712);
nor U17860 (N_17860,N_17767,N_17639);
or U17861 (N_17861,N_17727,N_17613);
nor U17862 (N_17862,N_17736,N_17737);
nor U17863 (N_17863,N_17650,N_17709);
xor U17864 (N_17864,N_17784,N_17726);
nor U17865 (N_17865,N_17720,N_17638);
or U17866 (N_17866,N_17744,N_17740);
xor U17867 (N_17867,N_17769,N_17689);
xor U17868 (N_17868,N_17675,N_17630);
nor U17869 (N_17869,N_17653,N_17666);
or U17870 (N_17870,N_17684,N_17701);
nand U17871 (N_17871,N_17679,N_17634);
xnor U17872 (N_17872,N_17605,N_17685);
or U17873 (N_17873,N_17652,N_17637);
or U17874 (N_17874,N_17750,N_17601);
nor U17875 (N_17875,N_17771,N_17761);
nand U17876 (N_17876,N_17699,N_17626);
and U17877 (N_17877,N_17723,N_17646);
or U17878 (N_17878,N_17745,N_17786);
xnor U17879 (N_17879,N_17660,N_17603);
nand U17880 (N_17880,N_17695,N_17686);
and U17881 (N_17881,N_17620,N_17665);
or U17882 (N_17882,N_17703,N_17663);
nand U17883 (N_17883,N_17733,N_17707);
nor U17884 (N_17884,N_17682,N_17655);
and U17885 (N_17885,N_17662,N_17617);
nand U17886 (N_17886,N_17622,N_17623);
nand U17887 (N_17887,N_17681,N_17668);
nand U17888 (N_17888,N_17758,N_17743);
and U17889 (N_17889,N_17644,N_17711);
xnor U17890 (N_17890,N_17618,N_17609);
nand U17891 (N_17891,N_17798,N_17683);
xnor U17892 (N_17892,N_17627,N_17649);
nor U17893 (N_17893,N_17633,N_17635);
nand U17894 (N_17894,N_17697,N_17690);
xor U17895 (N_17895,N_17640,N_17636);
or U17896 (N_17896,N_17631,N_17756);
and U17897 (N_17897,N_17687,N_17759);
nand U17898 (N_17898,N_17719,N_17692);
xnor U17899 (N_17899,N_17716,N_17747);
nor U17900 (N_17900,N_17623,N_17735);
or U17901 (N_17901,N_17608,N_17799);
nand U17902 (N_17902,N_17748,N_17734);
xor U17903 (N_17903,N_17630,N_17694);
or U17904 (N_17904,N_17692,N_17712);
nor U17905 (N_17905,N_17749,N_17761);
or U17906 (N_17906,N_17685,N_17672);
nand U17907 (N_17907,N_17749,N_17721);
and U17908 (N_17908,N_17788,N_17752);
and U17909 (N_17909,N_17799,N_17654);
and U17910 (N_17910,N_17767,N_17772);
nor U17911 (N_17911,N_17686,N_17747);
nand U17912 (N_17912,N_17682,N_17794);
xnor U17913 (N_17913,N_17637,N_17765);
or U17914 (N_17914,N_17701,N_17672);
nand U17915 (N_17915,N_17670,N_17654);
nor U17916 (N_17916,N_17636,N_17781);
or U17917 (N_17917,N_17711,N_17688);
nor U17918 (N_17918,N_17669,N_17611);
and U17919 (N_17919,N_17705,N_17719);
xnor U17920 (N_17920,N_17681,N_17750);
nor U17921 (N_17921,N_17666,N_17603);
nand U17922 (N_17922,N_17699,N_17799);
nand U17923 (N_17923,N_17609,N_17660);
nand U17924 (N_17924,N_17645,N_17772);
or U17925 (N_17925,N_17680,N_17670);
and U17926 (N_17926,N_17795,N_17784);
nor U17927 (N_17927,N_17732,N_17641);
nor U17928 (N_17928,N_17718,N_17677);
or U17929 (N_17929,N_17721,N_17647);
or U17930 (N_17930,N_17754,N_17687);
xnor U17931 (N_17931,N_17664,N_17744);
xor U17932 (N_17932,N_17795,N_17652);
xor U17933 (N_17933,N_17796,N_17729);
and U17934 (N_17934,N_17754,N_17605);
and U17935 (N_17935,N_17701,N_17648);
nor U17936 (N_17936,N_17732,N_17766);
xor U17937 (N_17937,N_17692,N_17774);
nand U17938 (N_17938,N_17776,N_17719);
nand U17939 (N_17939,N_17681,N_17786);
or U17940 (N_17940,N_17747,N_17783);
or U17941 (N_17941,N_17665,N_17768);
and U17942 (N_17942,N_17702,N_17749);
nand U17943 (N_17943,N_17660,N_17659);
xor U17944 (N_17944,N_17730,N_17742);
xor U17945 (N_17945,N_17674,N_17627);
xor U17946 (N_17946,N_17619,N_17662);
and U17947 (N_17947,N_17629,N_17646);
and U17948 (N_17948,N_17622,N_17621);
nor U17949 (N_17949,N_17708,N_17653);
nand U17950 (N_17950,N_17660,N_17681);
nand U17951 (N_17951,N_17706,N_17726);
or U17952 (N_17952,N_17661,N_17720);
nand U17953 (N_17953,N_17634,N_17676);
nor U17954 (N_17954,N_17772,N_17648);
nor U17955 (N_17955,N_17702,N_17729);
nand U17956 (N_17956,N_17733,N_17666);
nor U17957 (N_17957,N_17607,N_17667);
xor U17958 (N_17958,N_17726,N_17698);
or U17959 (N_17959,N_17772,N_17635);
xnor U17960 (N_17960,N_17770,N_17616);
and U17961 (N_17961,N_17682,N_17764);
and U17962 (N_17962,N_17647,N_17723);
xor U17963 (N_17963,N_17705,N_17733);
and U17964 (N_17964,N_17767,N_17682);
xor U17965 (N_17965,N_17679,N_17624);
xnor U17966 (N_17966,N_17635,N_17623);
nand U17967 (N_17967,N_17683,N_17656);
xnor U17968 (N_17968,N_17780,N_17750);
xnor U17969 (N_17969,N_17741,N_17791);
nand U17970 (N_17970,N_17738,N_17646);
nand U17971 (N_17971,N_17741,N_17602);
nor U17972 (N_17972,N_17794,N_17766);
nand U17973 (N_17973,N_17650,N_17737);
nor U17974 (N_17974,N_17731,N_17798);
nor U17975 (N_17975,N_17787,N_17723);
xnor U17976 (N_17976,N_17703,N_17761);
xnor U17977 (N_17977,N_17781,N_17725);
xnor U17978 (N_17978,N_17763,N_17712);
nor U17979 (N_17979,N_17657,N_17704);
xnor U17980 (N_17980,N_17680,N_17603);
nand U17981 (N_17981,N_17797,N_17765);
xor U17982 (N_17982,N_17695,N_17648);
or U17983 (N_17983,N_17638,N_17648);
or U17984 (N_17984,N_17658,N_17695);
nor U17985 (N_17985,N_17744,N_17769);
nand U17986 (N_17986,N_17794,N_17602);
xor U17987 (N_17987,N_17740,N_17642);
and U17988 (N_17988,N_17670,N_17711);
nand U17989 (N_17989,N_17719,N_17732);
nor U17990 (N_17990,N_17705,N_17672);
and U17991 (N_17991,N_17777,N_17700);
xnor U17992 (N_17992,N_17623,N_17753);
or U17993 (N_17993,N_17796,N_17631);
nor U17994 (N_17994,N_17621,N_17744);
xor U17995 (N_17995,N_17720,N_17706);
and U17996 (N_17996,N_17771,N_17711);
xnor U17997 (N_17997,N_17771,N_17622);
nor U17998 (N_17998,N_17737,N_17608);
nor U17999 (N_17999,N_17625,N_17615);
nand U18000 (N_18000,N_17864,N_17837);
and U18001 (N_18001,N_17899,N_17995);
and U18002 (N_18002,N_17931,N_17926);
nand U18003 (N_18003,N_17889,N_17829);
or U18004 (N_18004,N_17904,N_17934);
xor U18005 (N_18005,N_17944,N_17838);
nand U18006 (N_18006,N_17978,N_17930);
and U18007 (N_18007,N_17900,N_17824);
or U18008 (N_18008,N_17848,N_17923);
or U18009 (N_18009,N_17855,N_17828);
and U18010 (N_18010,N_17884,N_17928);
nor U18011 (N_18011,N_17981,N_17826);
and U18012 (N_18012,N_17892,N_17808);
nand U18013 (N_18013,N_17968,N_17887);
or U18014 (N_18014,N_17856,N_17844);
nand U18015 (N_18015,N_17911,N_17810);
nor U18016 (N_18016,N_17945,N_17953);
nor U18017 (N_18017,N_17922,N_17893);
and U18018 (N_18018,N_17852,N_17959);
nor U18019 (N_18019,N_17835,N_17890);
and U18020 (N_18020,N_17989,N_17999);
and U18021 (N_18021,N_17806,N_17840);
xnor U18022 (N_18022,N_17876,N_17952);
nand U18023 (N_18023,N_17992,N_17818);
or U18024 (N_18024,N_17976,N_17918);
and U18025 (N_18025,N_17958,N_17822);
xnor U18026 (N_18026,N_17813,N_17935);
and U18027 (N_18027,N_17817,N_17932);
nand U18028 (N_18028,N_17871,N_17929);
xnor U18029 (N_18029,N_17907,N_17815);
nor U18030 (N_18030,N_17846,N_17843);
nor U18031 (N_18031,N_17853,N_17860);
or U18032 (N_18032,N_17803,N_17927);
and U18033 (N_18033,N_17994,N_17885);
or U18034 (N_18034,N_17820,N_17975);
or U18035 (N_18035,N_17964,N_17880);
and U18036 (N_18036,N_17888,N_17913);
xor U18037 (N_18037,N_17969,N_17894);
nor U18038 (N_18038,N_17903,N_17939);
nor U18039 (N_18039,N_17960,N_17827);
or U18040 (N_18040,N_17863,N_17906);
nand U18041 (N_18041,N_17874,N_17951);
and U18042 (N_18042,N_17883,N_17854);
xnor U18043 (N_18043,N_17983,N_17825);
xor U18044 (N_18044,N_17972,N_17850);
xnor U18045 (N_18045,N_17823,N_17910);
nor U18046 (N_18046,N_17950,N_17861);
or U18047 (N_18047,N_17800,N_17857);
and U18048 (N_18048,N_17970,N_17819);
xor U18049 (N_18049,N_17802,N_17984);
xnor U18050 (N_18050,N_17915,N_17809);
or U18051 (N_18051,N_17988,N_17933);
nand U18052 (N_18052,N_17886,N_17921);
nor U18053 (N_18053,N_17916,N_17971);
nor U18054 (N_18054,N_17963,N_17908);
xor U18055 (N_18055,N_17973,N_17901);
and U18056 (N_18056,N_17961,N_17949);
xnor U18057 (N_18057,N_17875,N_17805);
nor U18058 (N_18058,N_17867,N_17862);
or U18059 (N_18059,N_17858,N_17896);
xnor U18060 (N_18060,N_17993,N_17940);
xnor U18061 (N_18061,N_17909,N_17836);
nor U18062 (N_18062,N_17925,N_17847);
and U18063 (N_18063,N_17845,N_17991);
or U18064 (N_18064,N_17987,N_17842);
and U18065 (N_18065,N_17905,N_17966);
or U18066 (N_18066,N_17865,N_17879);
nor U18067 (N_18067,N_17917,N_17996);
and U18068 (N_18068,N_17801,N_17980);
xnor U18069 (N_18069,N_17891,N_17998);
nand U18070 (N_18070,N_17841,N_17869);
nand U18071 (N_18071,N_17956,N_17866);
nand U18072 (N_18072,N_17873,N_17821);
or U18073 (N_18073,N_17965,N_17912);
and U18074 (N_18074,N_17974,N_17982);
nor U18075 (N_18075,N_17954,N_17881);
or U18076 (N_18076,N_17849,N_17859);
and U18077 (N_18077,N_17943,N_17877);
or U18078 (N_18078,N_17962,N_17990);
xnor U18079 (N_18079,N_17902,N_17897);
and U18080 (N_18080,N_17924,N_17979);
nand U18081 (N_18081,N_17872,N_17895);
and U18082 (N_18082,N_17833,N_17919);
xnor U18083 (N_18083,N_17834,N_17977);
or U18084 (N_18084,N_17816,N_17814);
nor U18085 (N_18085,N_17985,N_17967);
nand U18086 (N_18086,N_17812,N_17807);
nand U18087 (N_18087,N_17804,N_17811);
and U18088 (N_18088,N_17947,N_17868);
nor U18089 (N_18089,N_17878,N_17948);
nand U18090 (N_18090,N_17938,N_17832);
nor U18091 (N_18091,N_17851,N_17920);
nand U18092 (N_18092,N_17898,N_17936);
and U18093 (N_18093,N_17957,N_17955);
or U18094 (N_18094,N_17882,N_17914);
nor U18095 (N_18095,N_17941,N_17942);
and U18096 (N_18096,N_17839,N_17830);
nor U18097 (N_18097,N_17870,N_17997);
xor U18098 (N_18098,N_17946,N_17937);
nand U18099 (N_18099,N_17986,N_17831);
and U18100 (N_18100,N_17832,N_17952);
xor U18101 (N_18101,N_17914,N_17854);
nand U18102 (N_18102,N_17965,N_17843);
nand U18103 (N_18103,N_17879,N_17938);
nand U18104 (N_18104,N_17821,N_17884);
or U18105 (N_18105,N_17813,N_17942);
and U18106 (N_18106,N_17887,N_17999);
xnor U18107 (N_18107,N_17978,N_17876);
or U18108 (N_18108,N_17818,N_17856);
or U18109 (N_18109,N_17813,N_17997);
and U18110 (N_18110,N_17830,N_17980);
and U18111 (N_18111,N_17958,N_17911);
or U18112 (N_18112,N_17844,N_17974);
and U18113 (N_18113,N_17982,N_17984);
nand U18114 (N_18114,N_17837,N_17802);
and U18115 (N_18115,N_17809,N_17845);
xnor U18116 (N_18116,N_17810,N_17876);
nor U18117 (N_18117,N_17830,N_17983);
nor U18118 (N_18118,N_17969,N_17827);
xor U18119 (N_18119,N_17804,N_17974);
and U18120 (N_18120,N_17992,N_17803);
nand U18121 (N_18121,N_17971,N_17881);
xnor U18122 (N_18122,N_17941,N_17847);
and U18123 (N_18123,N_17820,N_17972);
and U18124 (N_18124,N_17958,N_17931);
nor U18125 (N_18125,N_17981,N_17873);
xnor U18126 (N_18126,N_17810,N_17852);
xnor U18127 (N_18127,N_17937,N_17847);
nand U18128 (N_18128,N_17864,N_17875);
and U18129 (N_18129,N_17900,N_17929);
and U18130 (N_18130,N_17826,N_17851);
nand U18131 (N_18131,N_17885,N_17829);
or U18132 (N_18132,N_17828,N_17804);
or U18133 (N_18133,N_17983,N_17804);
xnor U18134 (N_18134,N_17854,N_17889);
xnor U18135 (N_18135,N_17838,N_17874);
and U18136 (N_18136,N_17897,N_17914);
or U18137 (N_18137,N_17901,N_17939);
and U18138 (N_18138,N_17977,N_17918);
nor U18139 (N_18139,N_17894,N_17922);
and U18140 (N_18140,N_17954,N_17990);
nor U18141 (N_18141,N_17945,N_17848);
or U18142 (N_18142,N_17870,N_17957);
nand U18143 (N_18143,N_17943,N_17971);
and U18144 (N_18144,N_17813,N_17808);
and U18145 (N_18145,N_17922,N_17850);
and U18146 (N_18146,N_17868,N_17985);
nor U18147 (N_18147,N_17848,N_17941);
nor U18148 (N_18148,N_17933,N_17951);
or U18149 (N_18149,N_17843,N_17909);
xor U18150 (N_18150,N_17884,N_17832);
nand U18151 (N_18151,N_17897,N_17802);
nor U18152 (N_18152,N_17836,N_17966);
nor U18153 (N_18153,N_17894,N_17990);
xor U18154 (N_18154,N_17964,N_17858);
and U18155 (N_18155,N_17934,N_17946);
xor U18156 (N_18156,N_17988,N_17895);
nor U18157 (N_18157,N_17856,N_17944);
nor U18158 (N_18158,N_17974,N_17922);
xor U18159 (N_18159,N_17969,N_17941);
and U18160 (N_18160,N_17897,N_17806);
or U18161 (N_18161,N_17911,N_17927);
or U18162 (N_18162,N_17963,N_17926);
or U18163 (N_18163,N_17963,N_17869);
and U18164 (N_18164,N_17998,N_17970);
and U18165 (N_18165,N_17885,N_17862);
and U18166 (N_18166,N_17826,N_17865);
or U18167 (N_18167,N_17831,N_17954);
nand U18168 (N_18168,N_17987,N_17993);
nor U18169 (N_18169,N_17803,N_17953);
nand U18170 (N_18170,N_17866,N_17939);
nor U18171 (N_18171,N_17971,N_17818);
nor U18172 (N_18172,N_17902,N_17831);
or U18173 (N_18173,N_17929,N_17999);
and U18174 (N_18174,N_17840,N_17980);
nor U18175 (N_18175,N_17960,N_17910);
or U18176 (N_18176,N_17857,N_17815);
nor U18177 (N_18177,N_17997,N_17956);
nor U18178 (N_18178,N_17925,N_17965);
and U18179 (N_18179,N_17852,N_17916);
and U18180 (N_18180,N_17801,N_17865);
nand U18181 (N_18181,N_17930,N_17987);
and U18182 (N_18182,N_17990,N_17829);
and U18183 (N_18183,N_17824,N_17883);
xor U18184 (N_18184,N_17843,N_17995);
nor U18185 (N_18185,N_17814,N_17823);
nand U18186 (N_18186,N_17859,N_17980);
xor U18187 (N_18187,N_17803,N_17997);
nand U18188 (N_18188,N_17818,N_17875);
nand U18189 (N_18189,N_17979,N_17956);
and U18190 (N_18190,N_17824,N_17845);
xor U18191 (N_18191,N_17807,N_17930);
or U18192 (N_18192,N_17963,N_17876);
nor U18193 (N_18193,N_17983,N_17916);
nor U18194 (N_18194,N_17864,N_17971);
xor U18195 (N_18195,N_17975,N_17849);
and U18196 (N_18196,N_17864,N_17865);
or U18197 (N_18197,N_17912,N_17809);
nor U18198 (N_18198,N_17993,N_17871);
xor U18199 (N_18199,N_17997,N_17908);
nand U18200 (N_18200,N_18038,N_18177);
xor U18201 (N_18201,N_18188,N_18164);
nand U18202 (N_18202,N_18071,N_18116);
or U18203 (N_18203,N_18157,N_18155);
and U18204 (N_18204,N_18152,N_18101);
or U18205 (N_18205,N_18007,N_18107);
nand U18206 (N_18206,N_18161,N_18032);
nor U18207 (N_18207,N_18045,N_18193);
nor U18208 (N_18208,N_18115,N_18044);
nor U18209 (N_18209,N_18004,N_18066);
nand U18210 (N_18210,N_18112,N_18118);
xor U18211 (N_18211,N_18182,N_18048);
nor U18212 (N_18212,N_18108,N_18176);
nand U18213 (N_18213,N_18133,N_18034);
nor U18214 (N_18214,N_18012,N_18099);
xnor U18215 (N_18215,N_18005,N_18073);
and U18216 (N_18216,N_18078,N_18162);
nor U18217 (N_18217,N_18196,N_18185);
nor U18218 (N_18218,N_18030,N_18106);
nor U18219 (N_18219,N_18061,N_18100);
xnor U18220 (N_18220,N_18173,N_18065);
and U18221 (N_18221,N_18136,N_18156);
or U18222 (N_18222,N_18120,N_18001);
or U18223 (N_18223,N_18130,N_18060);
and U18224 (N_18224,N_18077,N_18062);
or U18225 (N_18225,N_18085,N_18175);
nand U18226 (N_18226,N_18083,N_18141);
nor U18227 (N_18227,N_18017,N_18058);
or U18228 (N_18228,N_18080,N_18160);
nor U18229 (N_18229,N_18070,N_18178);
nand U18230 (N_18230,N_18103,N_18137);
nor U18231 (N_18231,N_18006,N_18190);
and U18232 (N_18232,N_18138,N_18015);
xor U18233 (N_18233,N_18184,N_18019);
xor U18234 (N_18234,N_18072,N_18020);
nor U18235 (N_18235,N_18154,N_18117);
or U18236 (N_18236,N_18081,N_18129);
and U18237 (N_18237,N_18104,N_18131);
nor U18238 (N_18238,N_18194,N_18110);
nor U18239 (N_18239,N_18195,N_18169);
nand U18240 (N_18240,N_18187,N_18093);
nor U18241 (N_18241,N_18009,N_18109);
and U18242 (N_18242,N_18135,N_18046);
and U18243 (N_18243,N_18165,N_18150);
and U18244 (N_18244,N_18170,N_18147);
and U18245 (N_18245,N_18124,N_18163);
and U18246 (N_18246,N_18097,N_18172);
or U18247 (N_18247,N_18088,N_18047);
xnor U18248 (N_18248,N_18091,N_18128);
xnor U18249 (N_18249,N_18181,N_18033);
nand U18250 (N_18250,N_18000,N_18086);
and U18251 (N_18251,N_18010,N_18064);
nor U18252 (N_18252,N_18122,N_18022);
or U18253 (N_18253,N_18043,N_18145);
nor U18254 (N_18254,N_18158,N_18036);
or U18255 (N_18255,N_18197,N_18037);
and U18256 (N_18256,N_18183,N_18199);
nor U18257 (N_18257,N_18011,N_18042);
and U18258 (N_18258,N_18014,N_18031);
or U18259 (N_18259,N_18139,N_18180);
and U18260 (N_18260,N_18035,N_18192);
or U18261 (N_18261,N_18089,N_18167);
and U18262 (N_18262,N_18049,N_18179);
and U18263 (N_18263,N_18016,N_18113);
xnor U18264 (N_18264,N_18053,N_18121);
nor U18265 (N_18265,N_18084,N_18025);
nor U18266 (N_18266,N_18008,N_18144);
nor U18267 (N_18267,N_18082,N_18052);
and U18268 (N_18268,N_18125,N_18114);
and U18269 (N_18269,N_18198,N_18095);
xor U18270 (N_18270,N_18067,N_18098);
xor U18271 (N_18271,N_18096,N_18132);
and U18272 (N_18272,N_18076,N_18140);
or U18273 (N_18273,N_18051,N_18143);
nor U18274 (N_18274,N_18087,N_18151);
and U18275 (N_18275,N_18050,N_18123);
nor U18276 (N_18276,N_18126,N_18168);
and U18277 (N_18277,N_18102,N_18148);
xor U18278 (N_18278,N_18039,N_18159);
nor U18279 (N_18279,N_18023,N_18057);
nand U18280 (N_18280,N_18149,N_18027);
nor U18281 (N_18281,N_18191,N_18054);
or U18282 (N_18282,N_18079,N_18146);
nand U18283 (N_18283,N_18127,N_18018);
or U18284 (N_18284,N_18171,N_18068);
nor U18285 (N_18285,N_18013,N_18092);
nand U18286 (N_18286,N_18111,N_18134);
or U18287 (N_18287,N_18075,N_18186);
xor U18288 (N_18288,N_18074,N_18142);
nor U18289 (N_18289,N_18055,N_18002);
and U18290 (N_18290,N_18056,N_18153);
xor U18291 (N_18291,N_18041,N_18029);
nor U18292 (N_18292,N_18026,N_18063);
nor U18293 (N_18293,N_18189,N_18094);
or U18294 (N_18294,N_18059,N_18119);
or U18295 (N_18295,N_18105,N_18024);
and U18296 (N_18296,N_18069,N_18028);
xor U18297 (N_18297,N_18040,N_18003);
or U18298 (N_18298,N_18166,N_18021);
xor U18299 (N_18299,N_18090,N_18174);
nand U18300 (N_18300,N_18154,N_18179);
or U18301 (N_18301,N_18144,N_18130);
nand U18302 (N_18302,N_18084,N_18068);
xor U18303 (N_18303,N_18140,N_18067);
nor U18304 (N_18304,N_18162,N_18141);
or U18305 (N_18305,N_18042,N_18047);
or U18306 (N_18306,N_18144,N_18092);
nor U18307 (N_18307,N_18028,N_18056);
nand U18308 (N_18308,N_18054,N_18076);
xor U18309 (N_18309,N_18148,N_18086);
and U18310 (N_18310,N_18056,N_18146);
nand U18311 (N_18311,N_18009,N_18144);
or U18312 (N_18312,N_18087,N_18178);
or U18313 (N_18313,N_18030,N_18183);
or U18314 (N_18314,N_18033,N_18071);
nor U18315 (N_18315,N_18064,N_18053);
nand U18316 (N_18316,N_18035,N_18193);
or U18317 (N_18317,N_18130,N_18032);
nand U18318 (N_18318,N_18156,N_18120);
nor U18319 (N_18319,N_18160,N_18035);
nor U18320 (N_18320,N_18023,N_18075);
and U18321 (N_18321,N_18055,N_18152);
xor U18322 (N_18322,N_18052,N_18170);
xor U18323 (N_18323,N_18173,N_18159);
xnor U18324 (N_18324,N_18139,N_18038);
xnor U18325 (N_18325,N_18087,N_18046);
xor U18326 (N_18326,N_18081,N_18105);
nor U18327 (N_18327,N_18185,N_18031);
and U18328 (N_18328,N_18026,N_18153);
nor U18329 (N_18329,N_18196,N_18109);
or U18330 (N_18330,N_18061,N_18199);
nor U18331 (N_18331,N_18017,N_18198);
or U18332 (N_18332,N_18030,N_18107);
and U18333 (N_18333,N_18160,N_18138);
and U18334 (N_18334,N_18140,N_18011);
xor U18335 (N_18335,N_18004,N_18106);
and U18336 (N_18336,N_18195,N_18081);
nand U18337 (N_18337,N_18085,N_18084);
nand U18338 (N_18338,N_18021,N_18109);
and U18339 (N_18339,N_18078,N_18145);
nand U18340 (N_18340,N_18167,N_18176);
nor U18341 (N_18341,N_18095,N_18119);
nor U18342 (N_18342,N_18000,N_18097);
nor U18343 (N_18343,N_18170,N_18111);
and U18344 (N_18344,N_18062,N_18151);
or U18345 (N_18345,N_18036,N_18042);
nand U18346 (N_18346,N_18194,N_18011);
nor U18347 (N_18347,N_18153,N_18097);
and U18348 (N_18348,N_18117,N_18155);
nand U18349 (N_18349,N_18129,N_18113);
nand U18350 (N_18350,N_18171,N_18053);
or U18351 (N_18351,N_18065,N_18147);
or U18352 (N_18352,N_18155,N_18030);
and U18353 (N_18353,N_18145,N_18044);
nor U18354 (N_18354,N_18115,N_18128);
and U18355 (N_18355,N_18154,N_18194);
nor U18356 (N_18356,N_18055,N_18063);
nand U18357 (N_18357,N_18018,N_18039);
or U18358 (N_18358,N_18101,N_18163);
and U18359 (N_18359,N_18085,N_18108);
nand U18360 (N_18360,N_18169,N_18171);
nand U18361 (N_18361,N_18111,N_18143);
or U18362 (N_18362,N_18193,N_18140);
nor U18363 (N_18363,N_18128,N_18044);
or U18364 (N_18364,N_18030,N_18188);
nand U18365 (N_18365,N_18019,N_18101);
nor U18366 (N_18366,N_18000,N_18156);
xnor U18367 (N_18367,N_18139,N_18003);
nor U18368 (N_18368,N_18017,N_18148);
nor U18369 (N_18369,N_18136,N_18025);
or U18370 (N_18370,N_18122,N_18101);
xor U18371 (N_18371,N_18162,N_18086);
or U18372 (N_18372,N_18023,N_18092);
or U18373 (N_18373,N_18027,N_18187);
or U18374 (N_18374,N_18051,N_18079);
xnor U18375 (N_18375,N_18105,N_18077);
and U18376 (N_18376,N_18113,N_18017);
nand U18377 (N_18377,N_18016,N_18081);
nand U18378 (N_18378,N_18025,N_18198);
xnor U18379 (N_18379,N_18112,N_18144);
nand U18380 (N_18380,N_18167,N_18154);
xnor U18381 (N_18381,N_18149,N_18023);
and U18382 (N_18382,N_18036,N_18100);
or U18383 (N_18383,N_18128,N_18071);
and U18384 (N_18384,N_18001,N_18118);
nand U18385 (N_18385,N_18077,N_18048);
nor U18386 (N_18386,N_18071,N_18035);
or U18387 (N_18387,N_18099,N_18136);
or U18388 (N_18388,N_18130,N_18047);
nand U18389 (N_18389,N_18064,N_18030);
xnor U18390 (N_18390,N_18096,N_18187);
or U18391 (N_18391,N_18101,N_18076);
or U18392 (N_18392,N_18075,N_18036);
nand U18393 (N_18393,N_18071,N_18073);
and U18394 (N_18394,N_18038,N_18154);
nor U18395 (N_18395,N_18002,N_18042);
nor U18396 (N_18396,N_18062,N_18095);
or U18397 (N_18397,N_18034,N_18197);
nand U18398 (N_18398,N_18184,N_18023);
or U18399 (N_18399,N_18141,N_18038);
and U18400 (N_18400,N_18217,N_18319);
or U18401 (N_18401,N_18362,N_18234);
or U18402 (N_18402,N_18389,N_18395);
xor U18403 (N_18403,N_18317,N_18321);
nand U18404 (N_18404,N_18260,N_18235);
nand U18405 (N_18405,N_18279,N_18365);
nor U18406 (N_18406,N_18352,N_18375);
nor U18407 (N_18407,N_18351,N_18367);
and U18408 (N_18408,N_18378,N_18383);
or U18409 (N_18409,N_18361,N_18392);
nand U18410 (N_18410,N_18364,N_18278);
nand U18411 (N_18411,N_18307,N_18230);
nand U18412 (N_18412,N_18220,N_18311);
xnor U18413 (N_18413,N_18388,N_18303);
xnor U18414 (N_18414,N_18323,N_18272);
nand U18415 (N_18415,N_18338,N_18283);
nor U18416 (N_18416,N_18293,N_18329);
nor U18417 (N_18417,N_18216,N_18332);
nand U18418 (N_18418,N_18238,N_18369);
nand U18419 (N_18419,N_18245,N_18267);
nor U18420 (N_18420,N_18243,N_18259);
and U18421 (N_18421,N_18219,N_18231);
nor U18422 (N_18422,N_18398,N_18337);
xor U18423 (N_18423,N_18377,N_18273);
and U18424 (N_18424,N_18228,N_18394);
xnor U18425 (N_18425,N_18294,N_18281);
and U18426 (N_18426,N_18254,N_18203);
and U18427 (N_18427,N_18384,N_18300);
and U18428 (N_18428,N_18232,N_18318);
xor U18429 (N_18429,N_18380,N_18236);
and U18430 (N_18430,N_18315,N_18265);
nand U18431 (N_18431,N_18268,N_18206);
and U18432 (N_18432,N_18366,N_18233);
and U18433 (N_18433,N_18257,N_18313);
or U18434 (N_18434,N_18240,N_18340);
or U18435 (N_18435,N_18269,N_18286);
nand U18436 (N_18436,N_18348,N_18325);
or U18437 (N_18437,N_18356,N_18310);
nand U18438 (N_18438,N_18393,N_18358);
nor U18439 (N_18439,N_18306,N_18224);
xnor U18440 (N_18440,N_18251,N_18344);
or U18441 (N_18441,N_18295,N_18334);
and U18442 (N_18442,N_18371,N_18290);
nand U18443 (N_18443,N_18255,N_18386);
and U18444 (N_18444,N_18374,N_18350);
and U18445 (N_18445,N_18397,N_18354);
nor U18446 (N_18446,N_18221,N_18284);
xnor U18447 (N_18447,N_18343,N_18368);
xor U18448 (N_18448,N_18320,N_18201);
nand U18449 (N_18449,N_18305,N_18285);
and U18450 (N_18450,N_18353,N_18248);
nor U18451 (N_18451,N_18212,N_18274);
or U18452 (N_18452,N_18357,N_18253);
nand U18453 (N_18453,N_18381,N_18261);
nor U18454 (N_18454,N_18227,N_18211);
or U18455 (N_18455,N_18247,N_18333);
and U18456 (N_18456,N_18205,N_18302);
nor U18457 (N_18457,N_18359,N_18326);
and U18458 (N_18458,N_18347,N_18207);
nand U18459 (N_18459,N_18363,N_18342);
or U18460 (N_18460,N_18387,N_18244);
or U18461 (N_18461,N_18289,N_18266);
or U18462 (N_18462,N_18271,N_18297);
nand U18463 (N_18463,N_18209,N_18264);
nand U18464 (N_18464,N_18258,N_18200);
and U18465 (N_18465,N_18213,N_18301);
xor U18466 (N_18466,N_18246,N_18276);
or U18467 (N_18467,N_18336,N_18280);
nor U18468 (N_18468,N_18331,N_18382);
xor U18469 (N_18469,N_18339,N_18298);
and U18470 (N_18470,N_18291,N_18250);
and U18471 (N_18471,N_18391,N_18328);
and U18472 (N_18472,N_18242,N_18379);
and U18473 (N_18473,N_18324,N_18215);
nor U18474 (N_18474,N_18222,N_18208);
xnor U18475 (N_18475,N_18288,N_18335);
and U18476 (N_18476,N_18322,N_18316);
nor U18477 (N_18477,N_18370,N_18218);
xnor U18478 (N_18478,N_18210,N_18355);
nand U18479 (N_18479,N_18262,N_18390);
and U18480 (N_18480,N_18396,N_18330);
nand U18481 (N_18481,N_18341,N_18308);
and U18482 (N_18482,N_18360,N_18275);
xnor U18483 (N_18483,N_18204,N_18252);
xor U18484 (N_18484,N_18296,N_18226);
or U18485 (N_18485,N_18263,N_18214);
nor U18486 (N_18486,N_18277,N_18327);
xnor U18487 (N_18487,N_18287,N_18282);
and U18488 (N_18488,N_18345,N_18202);
xnor U18489 (N_18489,N_18229,N_18312);
nor U18490 (N_18490,N_18399,N_18373);
nand U18491 (N_18491,N_18372,N_18256);
and U18492 (N_18492,N_18223,N_18270);
nand U18493 (N_18493,N_18349,N_18309);
xor U18494 (N_18494,N_18314,N_18385);
and U18495 (N_18495,N_18299,N_18304);
xor U18496 (N_18496,N_18346,N_18225);
and U18497 (N_18497,N_18237,N_18249);
and U18498 (N_18498,N_18241,N_18376);
xnor U18499 (N_18499,N_18292,N_18239);
nor U18500 (N_18500,N_18362,N_18342);
xnor U18501 (N_18501,N_18358,N_18344);
and U18502 (N_18502,N_18260,N_18393);
nand U18503 (N_18503,N_18206,N_18314);
or U18504 (N_18504,N_18363,N_18356);
nor U18505 (N_18505,N_18303,N_18358);
nor U18506 (N_18506,N_18388,N_18366);
nor U18507 (N_18507,N_18205,N_18347);
xnor U18508 (N_18508,N_18226,N_18262);
nor U18509 (N_18509,N_18267,N_18222);
nor U18510 (N_18510,N_18347,N_18247);
nand U18511 (N_18511,N_18388,N_18314);
nand U18512 (N_18512,N_18303,N_18376);
xnor U18513 (N_18513,N_18277,N_18238);
and U18514 (N_18514,N_18223,N_18314);
and U18515 (N_18515,N_18257,N_18336);
or U18516 (N_18516,N_18272,N_18280);
and U18517 (N_18517,N_18315,N_18370);
or U18518 (N_18518,N_18280,N_18234);
xnor U18519 (N_18519,N_18398,N_18336);
nand U18520 (N_18520,N_18354,N_18201);
nand U18521 (N_18521,N_18389,N_18362);
or U18522 (N_18522,N_18352,N_18233);
nand U18523 (N_18523,N_18222,N_18223);
and U18524 (N_18524,N_18368,N_18364);
or U18525 (N_18525,N_18373,N_18367);
xnor U18526 (N_18526,N_18236,N_18244);
xor U18527 (N_18527,N_18346,N_18304);
nand U18528 (N_18528,N_18359,N_18231);
nor U18529 (N_18529,N_18225,N_18324);
nor U18530 (N_18530,N_18297,N_18389);
or U18531 (N_18531,N_18362,N_18375);
nor U18532 (N_18532,N_18385,N_18316);
or U18533 (N_18533,N_18263,N_18341);
nand U18534 (N_18534,N_18306,N_18356);
and U18535 (N_18535,N_18245,N_18279);
xor U18536 (N_18536,N_18387,N_18290);
nor U18537 (N_18537,N_18391,N_18330);
xor U18538 (N_18538,N_18218,N_18286);
or U18539 (N_18539,N_18375,N_18274);
and U18540 (N_18540,N_18366,N_18282);
and U18541 (N_18541,N_18311,N_18269);
nand U18542 (N_18542,N_18391,N_18271);
nor U18543 (N_18543,N_18391,N_18215);
and U18544 (N_18544,N_18274,N_18300);
and U18545 (N_18545,N_18243,N_18220);
xnor U18546 (N_18546,N_18289,N_18206);
nand U18547 (N_18547,N_18272,N_18397);
nand U18548 (N_18548,N_18356,N_18276);
nor U18549 (N_18549,N_18354,N_18229);
and U18550 (N_18550,N_18249,N_18330);
nor U18551 (N_18551,N_18331,N_18283);
nand U18552 (N_18552,N_18223,N_18291);
nand U18553 (N_18553,N_18279,N_18295);
nand U18554 (N_18554,N_18255,N_18210);
or U18555 (N_18555,N_18211,N_18369);
nand U18556 (N_18556,N_18393,N_18202);
or U18557 (N_18557,N_18250,N_18260);
xnor U18558 (N_18558,N_18239,N_18241);
and U18559 (N_18559,N_18367,N_18251);
nand U18560 (N_18560,N_18294,N_18398);
xnor U18561 (N_18561,N_18326,N_18253);
or U18562 (N_18562,N_18221,N_18235);
nor U18563 (N_18563,N_18378,N_18320);
nor U18564 (N_18564,N_18284,N_18224);
or U18565 (N_18565,N_18282,N_18203);
or U18566 (N_18566,N_18276,N_18321);
nor U18567 (N_18567,N_18322,N_18369);
and U18568 (N_18568,N_18342,N_18275);
nand U18569 (N_18569,N_18270,N_18221);
xor U18570 (N_18570,N_18208,N_18241);
xor U18571 (N_18571,N_18208,N_18229);
or U18572 (N_18572,N_18223,N_18304);
and U18573 (N_18573,N_18278,N_18265);
or U18574 (N_18574,N_18360,N_18230);
and U18575 (N_18575,N_18358,N_18259);
nor U18576 (N_18576,N_18262,N_18221);
xor U18577 (N_18577,N_18311,N_18366);
nor U18578 (N_18578,N_18305,N_18326);
xnor U18579 (N_18579,N_18383,N_18355);
or U18580 (N_18580,N_18342,N_18220);
nand U18581 (N_18581,N_18351,N_18317);
and U18582 (N_18582,N_18396,N_18358);
or U18583 (N_18583,N_18243,N_18355);
or U18584 (N_18584,N_18211,N_18253);
xor U18585 (N_18585,N_18274,N_18227);
nand U18586 (N_18586,N_18394,N_18287);
nor U18587 (N_18587,N_18276,N_18270);
or U18588 (N_18588,N_18206,N_18344);
nor U18589 (N_18589,N_18290,N_18269);
nor U18590 (N_18590,N_18321,N_18340);
or U18591 (N_18591,N_18299,N_18312);
nor U18592 (N_18592,N_18333,N_18380);
and U18593 (N_18593,N_18209,N_18332);
and U18594 (N_18594,N_18227,N_18290);
nand U18595 (N_18595,N_18318,N_18243);
nor U18596 (N_18596,N_18379,N_18357);
xnor U18597 (N_18597,N_18249,N_18383);
nand U18598 (N_18598,N_18351,N_18272);
xor U18599 (N_18599,N_18291,N_18264);
nand U18600 (N_18600,N_18434,N_18586);
and U18601 (N_18601,N_18407,N_18461);
xor U18602 (N_18602,N_18472,N_18563);
nand U18603 (N_18603,N_18424,N_18414);
nor U18604 (N_18604,N_18541,N_18455);
and U18605 (N_18605,N_18439,N_18533);
and U18606 (N_18606,N_18475,N_18494);
xor U18607 (N_18607,N_18408,N_18505);
or U18608 (N_18608,N_18430,N_18474);
or U18609 (N_18609,N_18592,N_18404);
and U18610 (N_18610,N_18555,N_18564);
or U18611 (N_18611,N_18545,N_18552);
or U18612 (N_18612,N_18512,N_18402);
nor U18613 (N_18613,N_18460,N_18478);
or U18614 (N_18614,N_18427,N_18553);
nor U18615 (N_18615,N_18489,N_18433);
nor U18616 (N_18616,N_18508,N_18510);
nor U18617 (N_18617,N_18464,N_18535);
nor U18618 (N_18618,N_18543,N_18567);
or U18619 (N_18619,N_18495,N_18569);
nand U18620 (N_18620,N_18480,N_18518);
and U18621 (N_18621,N_18463,N_18446);
xnor U18622 (N_18622,N_18536,N_18487);
or U18623 (N_18623,N_18524,N_18591);
nand U18624 (N_18624,N_18438,N_18457);
nor U18625 (N_18625,N_18447,N_18528);
or U18626 (N_18626,N_18484,N_18595);
nor U18627 (N_18627,N_18453,N_18443);
and U18628 (N_18628,N_18576,N_18465);
nor U18629 (N_18629,N_18468,N_18514);
nand U18630 (N_18630,N_18405,N_18415);
nand U18631 (N_18631,N_18582,N_18467);
nand U18632 (N_18632,N_18578,N_18483);
or U18633 (N_18633,N_18515,N_18527);
nand U18634 (N_18634,N_18575,N_18561);
xor U18635 (N_18635,N_18406,N_18470);
xor U18636 (N_18636,N_18519,N_18585);
nor U18637 (N_18637,N_18462,N_18425);
or U18638 (N_18638,N_18416,N_18566);
nand U18639 (N_18639,N_18598,N_18412);
or U18640 (N_18640,N_18431,N_18549);
nor U18641 (N_18641,N_18511,N_18444);
or U18642 (N_18642,N_18471,N_18459);
or U18643 (N_18643,N_18499,N_18491);
or U18644 (N_18644,N_18570,N_18449);
xnor U18645 (N_18645,N_18400,N_18458);
xnor U18646 (N_18646,N_18452,N_18419);
or U18647 (N_18647,N_18502,N_18454);
and U18648 (N_18648,N_18476,N_18559);
nand U18649 (N_18649,N_18557,N_18507);
nand U18650 (N_18650,N_18413,N_18574);
xor U18651 (N_18651,N_18403,N_18426);
xor U18652 (N_18652,N_18448,N_18479);
xor U18653 (N_18653,N_18498,N_18579);
and U18654 (N_18654,N_18581,N_18445);
nand U18655 (N_18655,N_18565,N_18584);
xor U18656 (N_18656,N_18485,N_18548);
and U18657 (N_18657,N_18544,N_18437);
and U18658 (N_18658,N_18554,N_18521);
xnor U18659 (N_18659,N_18594,N_18547);
or U18660 (N_18660,N_18421,N_18436);
xnor U18661 (N_18661,N_18560,N_18440);
xnor U18662 (N_18662,N_18532,N_18423);
or U18663 (N_18663,N_18525,N_18422);
xnor U18664 (N_18664,N_18546,N_18597);
nand U18665 (N_18665,N_18593,N_18517);
or U18666 (N_18666,N_18473,N_18537);
nor U18667 (N_18667,N_18435,N_18506);
nor U18668 (N_18668,N_18520,N_18530);
nor U18669 (N_18669,N_18500,N_18599);
and U18670 (N_18670,N_18588,N_18516);
nor U18671 (N_18671,N_18420,N_18497);
or U18672 (N_18672,N_18428,N_18432);
nor U18673 (N_18673,N_18587,N_18469);
nor U18674 (N_18674,N_18523,N_18529);
or U18675 (N_18675,N_18558,N_18450);
nor U18676 (N_18676,N_18493,N_18504);
xor U18677 (N_18677,N_18481,N_18522);
nand U18678 (N_18678,N_18571,N_18409);
or U18679 (N_18679,N_18596,N_18482);
and U18680 (N_18680,N_18531,N_18417);
nand U18681 (N_18681,N_18441,N_18456);
nand U18682 (N_18682,N_18490,N_18418);
or U18683 (N_18683,N_18501,N_18477);
nand U18684 (N_18684,N_18492,N_18429);
xnor U18685 (N_18685,N_18551,N_18401);
nand U18686 (N_18686,N_18580,N_18488);
or U18687 (N_18687,N_18539,N_18503);
and U18688 (N_18688,N_18572,N_18573);
xnor U18689 (N_18689,N_18550,N_18589);
or U18690 (N_18690,N_18451,N_18562);
nor U18691 (N_18691,N_18411,N_18509);
nor U18692 (N_18692,N_18466,N_18534);
and U18693 (N_18693,N_18442,N_18513);
nand U18694 (N_18694,N_18540,N_18590);
xnor U18695 (N_18695,N_18568,N_18556);
nor U18696 (N_18696,N_18583,N_18410);
nand U18697 (N_18697,N_18538,N_18542);
and U18698 (N_18698,N_18496,N_18577);
or U18699 (N_18699,N_18486,N_18526);
xnor U18700 (N_18700,N_18596,N_18571);
nor U18701 (N_18701,N_18490,N_18590);
and U18702 (N_18702,N_18405,N_18569);
and U18703 (N_18703,N_18464,N_18533);
xnor U18704 (N_18704,N_18486,N_18467);
nor U18705 (N_18705,N_18426,N_18566);
nand U18706 (N_18706,N_18496,N_18590);
xnor U18707 (N_18707,N_18542,N_18587);
and U18708 (N_18708,N_18412,N_18528);
xnor U18709 (N_18709,N_18577,N_18531);
nor U18710 (N_18710,N_18566,N_18558);
xnor U18711 (N_18711,N_18595,N_18530);
and U18712 (N_18712,N_18538,N_18530);
nand U18713 (N_18713,N_18423,N_18467);
nand U18714 (N_18714,N_18483,N_18479);
or U18715 (N_18715,N_18510,N_18556);
xor U18716 (N_18716,N_18407,N_18483);
nand U18717 (N_18717,N_18482,N_18513);
xor U18718 (N_18718,N_18462,N_18422);
and U18719 (N_18719,N_18496,N_18588);
or U18720 (N_18720,N_18551,N_18490);
xor U18721 (N_18721,N_18498,N_18438);
and U18722 (N_18722,N_18558,N_18452);
or U18723 (N_18723,N_18528,N_18525);
and U18724 (N_18724,N_18440,N_18485);
nor U18725 (N_18725,N_18491,N_18409);
or U18726 (N_18726,N_18571,N_18566);
or U18727 (N_18727,N_18502,N_18469);
or U18728 (N_18728,N_18501,N_18529);
and U18729 (N_18729,N_18512,N_18467);
nor U18730 (N_18730,N_18463,N_18578);
nor U18731 (N_18731,N_18451,N_18415);
nor U18732 (N_18732,N_18482,N_18451);
or U18733 (N_18733,N_18478,N_18406);
nor U18734 (N_18734,N_18471,N_18504);
xnor U18735 (N_18735,N_18573,N_18497);
nor U18736 (N_18736,N_18438,N_18518);
nand U18737 (N_18737,N_18478,N_18566);
and U18738 (N_18738,N_18468,N_18596);
nor U18739 (N_18739,N_18410,N_18408);
xor U18740 (N_18740,N_18403,N_18544);
nand U18741 (N_18741,N_18411,N_18499);
nor U18742 (N_18742,N_18482,N_18414);
nand U18743 (N_18743,N_18515,N_18560);
xnor U18744 (N_18744,N_18508,N_18506);
and U18745 (N_18745,N_18592,N_18401);
xor U18746 (N_18746,N_18491,N_18484);
nor U18747 (N_18747,N_18559,N_18525);
or U18748 (N_18748,N_18464,N_18524);
and U18749 (N_18749,N_18593,N_18541);
nand U18750 (N_18750,N_18542,N_18507);
or U18751 (N_18751,N_18492,N_18485);
nor U18752 (N_18752,N_18483,N_18544);
and U18753 (N_18753,N_18537,N_18402);
xor U18754 (N_18754,N_18408,N_18519);
or U18755 (N_18755,N_18594,N_18578);
nand U18756 (N_18756,N_18504,N_18469);
nor U18757 (N_18757,N_18499,N_18576);
xnor U18758 (N_18758,N_18536,N_18583);
and U18759 (N_18759,N_18424,N_18402);
xor U18760 (N_18760,N_18596,N_18515);
or U18761 (N_18761,N_18582,N_18524);
nor U18762 (N_18762,N_18426,N_18424);
nor U18763 (N_18763,N_18515,N_18497);
xor U18764 (N_18764,N_18462,N_18526);
xor U18765 (N_18765,N_18485,N_18528);
and U18766 (N_18766,N_18543,N_18405);
nand U18767 (N_18767,N_18496,N_18490);
nor U18768 (N_18768,N_18408,N_18594);
and U18769 (N_18769,N_18597,N_18509);
and U18770 (N_18770,N_18437,N_18594);
nor U18771 (N_18771,N_18463,N_18512);
nor U18772 (N_18772,N_18530,N_18401);
or U18773 (N_18773,N_18527,N_18484);
nand U18774 (N_18774,N_18588,N_18568);
xnor U18775 (N_18775,N_18495,N_18570);
and U18776 (N_18776,N_18409,N_18434);
or U18777 (N_18777,N_18439,N_18592);
and U18778 (N_18778,N_18538,N_18453);
and U18779 (N_18779,N_18560,N_18409);
nor U18780 (N_18780,N_18562,N_18566);
and U18781 (N_18781,N_18594,N_18462);
nand U18782 (N_18782,N_18456,N_18513);
or U18783 (N_18783,N_18560,N_18457);
nor U18784 (N_18784,N_18579,N_18540);
and U18785 (N_18785,N_18400,N_18576);
xor U18786 (N_18786,N_18590,N_18427);
and U18787 (N_18787,N_18456,N_18400);
and U18788 (N_18788,N_18416,N_18466);
xor U18789 (N_18789,N_18481,N_18471);
nor U18790 (N_18790,N_18498,N_18489);
and U18791 (N_18791,N_18597,N_18476);
and U18792 (N_18792,N_18472,N_18514);
xor U18793 (N_18793,N_18581,N_18470);
nand U18794 (N_18794,N_18561,N_18436);
or U18795 (N_18795,N_18442,N_18597);
nand U18796 (N_18796,N_18482,N_18478);
and U18797 (N_18797,N_18411,N_18417);
xnor U18798 (N_18798,N_18416,N_18580);
and U18799 (N_18799,N_18443,N_18488);
nand U18800 (N_18800,N_18790,N_18600);
nor U18801 (N_18801,N_18638,N_18749);
and U18802 (N_18802,N_18617,N_18640);
xor U18803 (N_18803,N_18721,N_18667);
nor U18804 (N_18804,N_18767,N_18697);
xnor U18805 (N_18805,N_18733,N_18687);
xnor U18806 (N_18806,N_18689,N_18745);
or U18807 (N_18807,N_18742,N_18743);
and U18808 (N_18808,N_18609,N_18608);
or U18809 (N_18809,N_18644,N_18741);
or U18810 (N_18810,N_18761,N_18695);
nor U18811 (N_18811,N_18684,N_18610);
xor U18812 (N_18812,N_18662,N_18646);
and U18813 (N_18813,N_18624,N_18645);
or U18814 (N_18814,N_18722,N_18788);
and U18815 (N_18815,N_18717,N_18602);
nand U18816 (N_18816,N_18792,N_18731);
or U18817 (N_18817,N_18630,N_18639);
xnor U18818 (N_18818,N_18704,N_18700);
nand U18819 (N_18819,N_18746,N_18701);
and U18820 (N_18820,N_18772,N_18784);
and U18821 (N_18821,N_18744,N_18654);
nor U18822 (N_18822,N_18737,N_18757);
and U18823 (N_18823,N_18711,N_18778);
nor U18824 (N_18824,N_18751,N_18773);
nor U18825 (N_18825,N_18604,N_18637);
xor U18826 (N_18826,N_18777,N_18780);
or U18827 (N_18827,N_18791,N_18677);
nor U18828 (N_18828,N_18696,N_18621);
nand U18829 (N_18829,N_18754,N_18682);
and U18830 (N_18830,N_18642,N_18668);
nand U18831 (N_18831,N_18719,N_18653);
nor U18832 (N_18832,N_18631,N_18774);
nor U18833 (N_18833,N_18724,N_18634);
and U18834 (N_18834,N_18736,N_18699);
and U18835 (N_18835,N_18750,N_18636);
and U18836 (N_18836,N_18673,N_18688);
or U18837 (N_18837,N_18715,N_18762);
nor U18838 (N_18838,N_18669,N_18718);
xor U18839 (N_18839,N_18649,N_18607);
and U18840 (N_18840,N_18633,N_18785);
and U18841 (N_18841,N_18755,N_18707);
and U18842 (N_18842,N_18635,N_18680);
nor U18843 (N_18843,N_18692,N_18665);
xnor U18844 (N_18844,N_18759,N_18789);
nand U18845 (N_18845,N_18660,N_18740);
nor U18846 (N_18846,N_18694,N_18647);
xnor U18847 (N_18847,N_18601,N_18614);
or U18848 (N_18848,N_18656,N_18686);
and U18849 (N_18849,N_18760,N_18620);
nor U18850 (N_18850,N_18655,N_18752);
xor U18851 (N_18851,N_18611,N_18613);
nor U18852 (N_18852,N_18712,N_18781);
xnor U18853 (N_18853,N_18782,N_18651);
or U18854 (N_18854,N_18674,N_18765);
or U18855 (N_18855,N_18658,N_18670);
or U18856 (N_18856,N_18771,N_18678);
nand U18857 (N_18857,N_18727,N_18675);
and U18858 (N_18858,N_18626,N_18641);
xor U18859 (N_18859,N_18720,N_18714);
xor U18860 (N_18860,N_18768,N_18723);
and U18861 (N_18861,N_18779,N_18632);
xor U18862 (N_18862,N_18628,N_18713);
and U18863 (N_18863,N_18683,N_18786);
or U18864 (N_18864,N_18787,N_18763);
xnor U18865 (N_18865,N_18769,N_18698);
nor U18866 (N_18866,N_18739,N_18685);
or U18867 (N_18867,N_18738,N_18730);
xnor U18868 (N_18868,N_18766,N_18661);
nor U18869 (N_18869,N_18625,N_18663);
xor U18870 (N_18870,N_18770,N_18706);
nand U18871 (N_18871,N_18664,N_18709);
or U18872 (N_18872,N_18690,N_18659);
nor U18873 (N_18873,N_18679,N_18783);
xor U18874 (N_18874,N_18794,N_18796);
nand U18875 (N_18875,N_18756,N_18622);
xnor U18876 (N_18876,N_18612,N_18623);
nand U18877 (N_18877,N_18618,N_18648);
and U18878 (N_18878,N_18676,N_18708);
nor U18879 (N_18879,N_18799,N_18776);
or U18880 (N_18880,N_18734,N_18728);
nand U18881 (N_18881,N_18764,N_18729);
nor U18882 (N_18882,N_18710,N_18797);
xnor U18883 (N_18883,N_18693,N_18643);
nor U18884 (N_18884,N_18726,N_18748);
nor U18885 (N_18885,N_18605,N_18652);
and U18886 (N_18886,N_18603,N_18629);
nand U18887 (N_18887,N_18758,N_18657);
or U18888 (N_18888,N_18798,N_18725);
or U18889 (N_18889,N_18702,N_18672);
or U18890 (N_18890,N_18627,N_18671);
or U18891 (N_18891,N_18650,N_18747);
xor U18892 (N_18892,N_18775,N_18606);
nand U18893 (N_18893,N_18666,N_18703);
xor U18894 (N_18894,N_18753,N_18735);
nand U18895 (N_18895,N_18795,N_18619);
xor U18896 (N_18896,N_18615,N_18616);
xnor U18897 (N_18897,N_18691,N_18793);
and U18898 (N_18898,N_18732,N_18681);
nor U18899 (N_18899,N_18705,N_18716);
xor U18900 (N_18900,N_18726,N_18793);
and U18901 (N_18901,N_18638,N_18685);
nand U18902 (N_18902,N_18784,N_18728);
nand U18903 (N_18903,N_18756,N_18738);
nand U18904 (N_18904,N_18653,N_18619);
nor U18905 (N_18905,N_18712,N_18707);
nor U18906 (N_18906,N_18606,N_18789);
and U18907 (N_18907,N_18725,N_18661);
xnor U18908 (N_18908,N_18622,N_18602);
xnor U18909 (N_18909,N_18605,N_18740);
nand U18910 (N_18910,N_18710,N_18640);
or U18911 (N_18911,N_18769,N_18781);
and U18912 (N_18912,N_18782,N_18698);
nor U18913 (N_18913,N_18783,N_18717);
or U18914 (N_18914,N_18712,N_18646);
and U18915 (N_18915,N_18758,N_18603);
or U18916 (N_18916,N_18777,N_18611);
nor U18917 (N_18917,N_18627,N_18654);
xor U18918 (N_18918,N_18680,N_18750);
nand U18919 (N_18919,N_18609,N_18644);
xor U18920 (N_18920,N_18709,N_18784);
or U18921 (N_18921,N_18652,N_18642);
nor U18922 (N_18922,N_18752,N_18677);
or U18923 (N_18923,N_18659,N_18706);
xor U18924 (N_18924,N_18778,N_18642);
nand U18925 (N_18925,N_18679,N_18604);
or U18926 (N_18926,N_18639,N_18734);
or U18927 (N_18927,N_18723,N_18634);
and U18928 (N_18928,N_18620,N_18694);
nor U18929 (N_18929,N_18694,N_18653);
and U18930 (N_18930,N_18662,N_18764);
nor U18931 (N_18931,N_18658,N_18628);
nand U18932 (N_18932,N_18731,N_18620);
and U18933 (N_18933,N_18637,N_18623);
xor U18934 (N_18934,N_18725,N_18711);
nor U18935 (N_18935,N_18613,N_18739);
or U18936 (N_18936,N_18618,N_18604);
nand U18937 (N_18937,N_18743,N_18739);
and U18938 (N_18938,N_18646,N_18730);
or U18939 (N_18939,N_18745,N_18624);
nand U18940 (N_18940,N_18635,N_18704);
nand U18941 (N_18941,N_18672,N_18699);
xor U18942 (N_18942,N_18610,N_18629);
nor U18943 (N_18943,N_18641,N_18727);
or U18944 (N_18944,N_18771,N_18762);
nor U18945 (N_18945,N_18771,N_18782);
and U18946 (N_18946,N_18634,N_18752);
and U18947 (N_18947,N_18787,N_18605);
xor U18948 (N_18948,N_18742,N_18612);
or U18949 (N_18949,N_18757,N_18623);
or U18950 (N_18950,N_18681,N_18713);
nor U18951 (N_18951,N_18661,N_18791);
xor U18952 (N_18952,N_18677,N_18757);
and U18953 (N_18953,N_18621,N_18784);
xor U18954 (N_18954,N_18661,N_18750);
xnor U18955 (N_18955,N_18773,N_18664);
or U18956 (N_18956,N_18749,N_18698);
and U18957 (N_18957,N_18621,N_18741);
nand U18958 (N_18958,N_18783,N_18709);
nand U18959 (N_18959,N_18680,N_18684);
or U18960 (N_18960,N_18726,N_18609);
and U18961 (N_18961,N_18632,N_18796);
xor U18962 (N_18962,N_18609,N_18704);
nand U18963 (N_18963,N_18655,N_18626);
nand U18964 (N_18964,N_18604,N_18636);
xor U18965 (N_18965,N_18770,N_18767);
nand U18966 (N_18966,N_18720,N_18601);
nand U18967 (N_18967,N_18763,N_18767);
and U18968 (N_18968,N_18647,N_18790);
or U18969 (N_18969,N_18642,N_18753);
and U18970 (N_18970,N_18671,N_18716);
or U18971 (N_18971,N_18611,N_18797);
and U18972 (N_18972,N_18643,N_18750);
nand U18973 (N_18973,N_18714,N_18719);
xor U18974 (N_18974,N_18784,N_18654);
and U18975 (N_18975,N_18704,N_18621);
nand U18976 (N_18976,N_18713,N_18649);
or U18977 (N_18977,N_18685,N_18778);
xnor U18978 (N_18978,N_18661,N_18665);
xor U18979 (N_18979,N_18648,N_18709);
or U18980 (N_18980,N_18710,N_18634);
or U18981 (N_18981,N_18798,N_18702);
or U18982 (N_18982,N_18761,N_18706);
or U18983 (N_18983,N_18727,N_18625);
or U18984 (N_18984,N_18723,N_18737);
xor U18985 (N_18985,N_18636,N_18792);
xnor U18986 (N_18986,N_18699,N_18714);
or U18987 (N_18987,N_18782,N_18649);
or U18988 (N_18988,N_18767,N_18631);
xor U18989 (N_18989,N_18624,N_18677);
nor U18990 (N_18990,N_18626,N_18767);
nand U18991 (N_18991,N_18665,N_18738);
and U18992 (N_18992,N_18644,N_18752);
and U18993 (N_18993,N_18693,N_18600);
or U18994 (N_18994,N_18738,N_18787);
or U18995 (N_18995,N_18678,N_18741);
xor U18996 (N_18996,N_18735,N_18608);
xor U18997 (N_18997,N_18702,N_18720);
or U18998 (N_18998,N_18628,N_18675);
nor U18999 (N_18999,N_18723,N_18620);
and U19000 (N_19000,N_18950,N_18842);
nand U19001 (N_19001,N_18951,N_18955);
and U19002 (N_19002,N_18820,N_18922);
nor U19003 (N_19003,N_18884,N_18947);
or U19004 (N_19004,N_18813,N_18850);
and U19005 (N_19005,N_18986,N_18910);
and U19006 (N_19006,N_18983,N_18969);
and U19007 (N_19007,N_18989,N_18901);
or U19008 (N_19008,N_18988,N_18994);
and U19009 (N_19009,N_18918,N_18911);
nor U19010 (N_19010,N_18900,N_18875);
nand U19011 (N_19011,N_18970,N_18872);
or U19012 (N_19012,N_18887,N_18948);
and U19013 (N_19013,N_18980,N_18973);
xnor U19014 (N_19014,N_18956,N_18972);
nor U19015 (N_19015,N_18830,N_18805);
nor U19016 (N_19016,N_18822,N_18844);
nand U19017 (N_19017,N_18971,N_18981);
xor U19018 (N_19018,N_18954,N_18839);
nor U19019 (N_19019,N_18936,N_18942);
or U19020 (N_19020,N_18898,N_18831);
and U19021 (N_19021,N_18808,N_18840);
nand U19022 (N_19022,N_18926,N_18941);
nor U19023 (N_19023,N_18874,N_18801);
nand U19024 (N_19024,N_18843,N_18987);
xnor U19025 (N_19025,N_18802,N_18979);
xnor U19026 (N_19026,N_18883,N_18919);
or U19027 (N_19027,N_18930,N_18902);
and U19028 (N_19028,N_18885,N_18834);
nor U19029 (N_19029,N_18803,N_18865);
xnor U19030 (N_19030,N_18832,N_18997);
and U19031 (N_19031,N_18877,N_18828);
and U19032 (N_19032,N_18846,N_18996);
or U19033 (N_19033,N_18929,N_18867);
xnor U19034 (N_19034,N_18823,N_18953);
xnor U19035 (N_19035,N_18928,N_18824);
and U19036 (N_19036,N_18838,N_18860);
nor U19037 (N_19037,N_18825,N_18976);
nand U19038 (N_19038,N_18886,N_18896);
nand U19039 (N_19039,N_18882,N_18890);
and U19040 (N_19040,N_18871,N_18811);
nand U19041 (N_19041,N_18892,N_18909);
nand U19042 (N_19042,N_18849,N_18836);
or U19043 (N_19043,N_18920,N_18934);
nor U19044 (N_19044,N_18982,N_18949);
or U19045 (N_19045,N_18946,N_18961);
xor U19046 (N_19046,N_18837,N_18863);
xnor U19047 (N_19047,N_18833,N_18881);
nand U19048 (N_19048,N_18998,N_18880);
xor U19049 (N_19049,N_18895,N_18957);
nor U19050 (N_19050,N_18852,N_18935);
and U19051 (N_19051,N_18856,N_18894);
or U19052 (N_19052,N_18974,N_18853);
xnor U19053 (N_19053,N_18905,N_18829);
nand U19054 (N_19054,N_18995,N_18845);
nor U19055 (N_19055,N_18873,N_18870);
nor U19056 (N_19056,N_18962,N_18876);
nor U19057 (N_19057,N_18903,N_18923);
or U19058 (N_19058,N_18807,N_18945);
and U19059 (N_19059,N_18848,N_18964);
and U19060 (N_19060,N_18924,N_18993);
and U19061 (N_19061,N_18819,N_18812);
or U19062 (N_19062,N_18931,N_18809);
xnor U19063 (N_19063,N_18815,N_18921);
or U19064 (N_19064,N_18851,N_18861);
and U19065 (N_19065,N_18913,N_18897);
or U19066 (N_19066,N_18917,N_18933);
or U19067 (N_19067,N_18963,N_18810);
nand U19068 (N_19068,N_18868,N_18916);
nand U19069 (N_19069,N_18859,N_18857);
and U19070 (N_19070,N_18943,N_18878);
and U19071 (N_19071,N_18965,N_18893);
xnor U19072 (N_19072,N_18817,N_18835);
nor U19073 (N_19073,N_18907,N_18952);
xnor U19074 (N_19074,N_18866,N_18814);
or U19075 (N_19075,N_18827,N_18966);
or U19076 (N_19076,N_18991,N_18944);
or U19077 (N_19077,N_18899,N_18938);
xor U19078 (N_19078,N_18800,N_18858);
xor U19079 (N_19079,N_18915,N_18959);
and U19080 (N_19080,N_18940,N_18854);
and U19081 (N_19081,N_18927,N_18960);
and U19082 (N_19082,N_18891,N_18806);
or U19083 (N_19083,N_18932,N_18804);
xnor U19084 (N_19084,N_18862,N_18985);
or U19085 (N_19085,N_18906,N_18821);
nor U19086 (N_19086,N_18816,N_18990);
xor U19087 (N_19087,N_18818,N_18826);
or U19088 (N_19088,N_18889,N_18908);
and U19089 (N_19089,N_18958,N_18869);
nand U19090 (N_19090,N_18925,N_18968);
nor U19091 (N_19091,N_18937,N_18939);
xor U19092 (N_19092,N_18904,N_18984);
or U19093 (N_19093,N_18967,N_18999);
xnor U19094 (N_19094,N_18855,N_18978);
xnor U19095 (N_19095,N_18912,N_18992);
nand U19096 (N_19096,N_18914,N_18864);
nand U19097 (N_19097,N_18847,N_18888);
or U19098 (N_19098,N_18879,N_18977);
or U19099 (N_19099,N_18841,N_18975);
nand U19100 (N_19100,N_18904,N_18803);
nand U19101 (N_19101,N_18922,N_18843);
xnor U19102 (N_19102,N_18996,N_18998);
xor U19103 (N_19103,N_18878,N_18836);
nor U19104 (N_19104,N_18977,N_18848);
xnor U19105 (N_19105,N_18851,N_18843);
nor U19106 (N_19106,N_18946,N_18984);
nor U19107 (N_19107,N_18862,N_18847);
nor U19108 (N_19108,N_18817,N_18866);
and U19109 (N_19109,N_18999,N_18995);
or U19110 (N_19110,N_18839,N_18868);
or U19111 (N_19111,N_18886,N_18884);
or U19112 (N_19112,N_18805,N_18892);
xnor U19113 (N_19113,N_18902,N_18816);
nor U19114 (N_19114,N_18969,N_18938);
and U19115 (N_19115,N_18923,N_18884);
nor U19116 (N_19116,N_18999,N_18941);
xor U19117 (N_19117,N_18802,N_18814);
or U19118 (N_19118,N_18945,N_18866);
nor U19119 (N_19119,N_18971,N_18897);
xor U19120 (N_19120,N_18857,N_18988);
and U19121 (N_19121,N_18917,N_18949);
xnor U19122 (N_19122,N_18836,N_18918);
xor U19123 (N_19123,N_18958,N_18830);
and U19124 (N_19124,N_18886,N_18999);
nor U19125 (N_19125,N_18983,N_18984);
nand U19126 (N_19126,N_18929,N_18925);
nor U19127 (N_19127,N_18864,N_18842);
xnor U19128 (N_19128,N_18863,N_18880);
xor U19129 (N_19129,N_18833,N_18957);
or U19130 (N_19130,N_18899,N_18887);
nand U19131 (N_19131,N_18908,N_18866);
and U19132 (N_19132,N_18834,N_18941);
or U19133 (N_19133,N_18931,N_18829);
or U19134 (N_19134,N_18869,N_18933);
nand U19135 (N_19135,N_18804,N_18818);
nand U19136 (N_19136,N_18820,N_18826);
nand U19137 (N_19137,N_18801,N_18845);
xor U19138 (N_19138,N_18917,N_18800);
or U19139 (N_19139,N_18910,N_18868);
nor U19140 (N_19140,N_18922,N_18800);
and U19141 (N_19141,N_18814,N_18938);
nor U19142 (N_19142,N_18906,N_18924);
xor U19143 (N_19143,N_18883,N_18953);
and U19144 (N_19144,N_18865,N_18820);
xor U19145 (N_19145,N_18815,N_18971);
xnor U19146 (N_19146,N_18891,N_18808);
nand U19147 (N_19147,N_18868,N_18882);
and U19148 (N_19148,N_18995,N_18806);
nor U19149 (N_19149,N_18926,N_18855);
and U19150 (N_19150,N_18882,N_18915);
xor U19151 (N_19151,N_18948,N_18826);
and U19152 (N_19152,N_18986,N_18889);
xor U19153 (N_19153,N_18902,N_18973);
and U19154 (N_19154,N_18890,N_18985);
and U19155 (N_19155,N_18971,N_18919);
xor U19156 (N_19156,N_18829,N_18899);
nor U19157 (N_19157,N_18906,N_18937);
xnor U19158 (N_19158,N_18948,N_18838);
and U19159 (N_19159,N_18909,N_18970);
xnor U19160 (N_19160,N_18985,N_18821);
and U19161 (N_19161,N_18823,N_18986);
xor U19162 (N_19162,N_18902,N_18958);
nand U19163 (N_19163,N_18942,N_18808);
xnor U19164 (N_19164,N_18846,N_18901);
nor U19165 (N_19165,N_18821,N_18871);
and U19166 (N_19166,N_18843,N_18854);
or U19167 (N_19167,N_18818,N_18887);
nand U19168 (N_19168,N_18890,N_18911);
xnor U19169 (N_19169,N_18965,N_18928);
nand U19170 (N_19170,N_18834,N_18857);
nand U19171 (N_19171,N_18939,N_18903);
xnor U19172 (N_19172,N_18870,N_18855);
or U19173 (N_19173,N_18916,N_18805);
and U19174 (N_19174,N_18808,N_18916);
or U19175 (N_19175,N_18869,N_18821);
nor U19176 (N_19176,N_18948,N_18980);
and U19177 (N_19177,N_18896,N_18918);
and U19178 (N_19178,N_18942,N_18938);
or U19179 (N_19179,N_18963,N_18897);
xnor U19180 (N_19180,N_18973,N_18854);
xor U19181 (N_19181,N_18841,N_18967);
or U19182 (N_19182,N_18958,N_18866);
or U19183 (N_19183,N_18978,N_18919);
or U19184 (N_19184,N_18920,N_18808);
xnor U19185 (N_19185,N_18928,N_18862);
and U19186 (N_19186,N_18954,N_18819);
nand U19187 (N_19187,N_18876,N_18815);
and U19188 (N_19188,N_18980,N_18938);
and U19189 (N_19189,N_18913,N_18885);
nor U19190 (N_19190,N_18890,N_18893);
and U19191 (N_19191,N_18943,N_18950);
or U19192 (N_19192,N_18891,N_18909);
nand U19193 (N_19193,N_18858,N_18811);
nor U19194 (N_19194,N_18822,N_18883);
nand U19195 (N_19195,N_18924,N_18874);
or U19196 (N_19196,N_18809,N_18865);
and U19197 (N_19197,N_18893,N_18987);
nand U19198 (N_19198,N_18907,N_18982);
or U19199 (N_19199,N_18813,N_18862);
nand U19200 (N_19200,N_19098,N_19070);
and U19201 (N_19201,N_19127,N_19102);
and U19202 (N_19202,N_19179,N_19160);
or U19203 (N_19203,N_19085,N_19073);
nand U19204 (N_19204,N_19185,N_19199);
and U19205 (N_19205,N_19065,N_19133);
nand U19206 (N_19206,N_19049,N_19155);
or U19207 (N_19207,N_19142,N_19119);
or U19208 (N_19208,N_19064,N_19174);
nor U19209 (N_19209,N_19161,N_19031);
nand U19210 (N_19210,N_19099,N_19191);
nand U19211 (N_19211,N_19158,N_19072);
or U19212 (N_19212,N_19112,N_19030);
nor U19213 (N_19213,N_19106,N_19092);
xnor U19214 (N_19214,N_19175,N_19146);
nor U19215 (N_19215,N_19132,N_19068);
and U19216 (N_19216,N_19004,N_19143);
nand U19217 (N_19217,N_19008,N_19192);
or U19218 (N_19218,N_19184,N_19122);
nor U19219 (N_19219,N_19013,N_19087);
xnor U19220 (N_19220,N_19080,N_19017);
and U19221 (N_19221,N_19164,N_19025);
xor U19222 (N_19222,N_19169,N_19003);
nand U19223 (N_19223,N_19009,N_19015);
or U19224 (N_19224,N_19168,N_19172);
nor U19225 (N_19225,N_19136,N_19043);
or U19226 (N_19226,N_19019,N_19089);
nand U19227 (N_19227,N_19007,N_19055);
or U19228 (N_19228,N_19110,N_19113);
nand U19229 (N_19229,N_19181,N_19189);
xor U19230 (N_19230,N_19152,N_19062);
and U19231 (N_19231,N_19145,N_19103);
or U19232 (N_19232,N_19141,N_19157);
or U19233 (N_19233,N_19120,N_19183);
or U19234 (N_19234,N_19006,N_19100);
nor U19235 (N_19235,N_19050,N_19057);
xor U19236 (N_19236,N_19014,N_19176);
nand U19237 (N_19237,N_19170,N_19052);
or U19238 (N_19238,N_19066,N_19107);
xnor U19239 (N_19239,N_19163,N_19059);
xor U19240 (N_19240,N_19097,N_19048);
and U19241 (N_19241,N_19045,N_19056);
nand U19242 (N_19242,N_19010,N_19134);
or U19243 (N_19243,N_19190,N_19069);
nand U19244 (N_19244,N_19151,N_19038);
nor U19245 (N_19245,N_19011,N_19091);
and U19246 (N_19246,N_19074,N_19028);
and U19247 (N_19247,N_19126,N_19021);
xnor U19248 (N_19248,N_19178,N_19076);
xor U19249 (N_19249,N_19083,N_19090);
nand U19250 (N_19250,N_19117,N_19000);
or U19251 (N_19251,N_19118,N_19124);
nand U19252 (N_19252,N_19108,N_19188);
xnor U19253 (N_19253,N_19159,N_19002);
nor U19254 (N_19254,N_19144,N_19153);
or U19255 (N_19255,N_19040,N_19104);
nand U19256 (N_19256,N_19034,N_19033);
and U19257 (N_19257,N_19075,N_19139);
and U19258 (N_19258,N_19061,N_19032);
xor U19259 (N_19259,N_19005,N_19114);
or U19260 (N_19260,N_19081,N_19037);
nor U19261 (N_19261,N_19029,N_19166);
xor U19262 (N_19262,N_19173,N_19054);
nand U19263 (N_19263,N_19084,N_19047);
or U19264 (N_19264,N_19194,N_19041);
xor U19265 (N_19265,N_19165,N_19078);
or U19266 (N_19266,N_19135,N_19149);
nor U19267 (N_19267,N_19111,N_19042);
or U19268 (N_19268,N_19186,N_19067);
nor U19269 (N_19269,N_19058,N_19128);
nand U19270 (N_19270,N_19177,N_19046);
nand U19271 (N_19271,N_19150,N_19137);
nor U19272 (N_19272,N_19079,N_19167);
nor U19273 (N_19273,N_19086,N_19154);
xor U19274 (N_19274,N_19129,N_19116);
nand U19275 (N_19275,N_19182,N_19121);
nand U19276 (N_19276,N_19138,N_19060);
and U19277 (N_19277,N_19077,N_19171);
and U19278 (N_19278,N_19082,N_19096);
xor U19279 (N_19279,N_19094,N_19039);
xnor U19280 (N_19280,N_19016,N_19012);
xor U19281 (N_19281,N_19044,N_19187);
and U19282 (N_19282,N_19093,N_19095);
or U19283 (N_19283,N_19140,N_19053);
xor U19284 (N_19284,N_19035,N_19156);
nand U19285 (N_19285,N_19148,N_19115);
xor U19286 (N_19286,N_19162,N_19022);
and U19287 (N_19287,N_19023,N_19147);
or U19288 (N_19288,N_19036,N_19125);
xor U19289 (N_19289,N_19105,N_19088);
and U19290 (N_19290,N_19197,N_19026);
xor U19291 (N_19291,N_19131,N_19109);
xnor U19292 (N_19292,N_19027,N_19196);
or U19293 (N_19293,N_19063,N_19051);
nand U19294 (N_19294,N_19198,N_19193);
nor U19295 (N_19295,N_19130,N_19018);
nor U19296 (N_19296,N_19024,N_19123);
nand U19297 (N_19297,N_19195,N_19001);
xnor U19298 (N_19298,N_19101,N_19180);
nor U19299 (N_19299,N_19020,N_19071);
or U19300 (N_19300,N_19153,N_19059);
xnor U19301 (N_19301,N_19035,N_19177);
nand U19302 (N_19302,N_19024,N_19191);
xnor U19303 (N_19303,N_19049,N_19116);
xnor U19304 (N_19304,N_19064,N_19046);
or U19305 (N_19305,N_19100,N_19102);
nand U19306 (N_19306,N_19113,N_19168);
and U19307 (N_19307,N_19007,N_19063);
nand U19308 (N_19308,N_19103,N_19133);
and U19309 (N_19309,N_19192,N_19062);
nor U19310 (N_19310,N_19165,N_19048);
and U19311 (N_19311,N_19043,N_19132);
xnor U19312 (N_19312,N_19124,N_19171);
or U19313 (N_19313,N_19180,N_19154);
nor U19314 (N_19314,N_19073,N_19026);
nor U19315 (N_19315,N_19075,N_19099);
or U19316 (N_19316,N_19086,N_19199);
xnor U19317 (N_19317,N_19060,N_19041);
nor U19318 (N_19318,N_19144,N_19111);
nand U19319 (N_19319,N_19148,N_19180);
nor U19320 (N_19320,N_19098,N_19146);
and U19321 (N_19321,N_19146,N_19117);
or U19322 (N_19322,N_19179,N_19153);
nand U19323 (N_19323,N_19005,N_19072);
and U19324 (N_19324,N_19073,N_19117);
and U19325 (N_19325,N_19088,N_19027);
or U19326 (N_19326,N_19074,N_19067);
and U19327 (N_19327,N_19024,N_19000);
nor U19328 (N_19328,N_19161,N_19192);
nor U19329 (N_19329,N_19138,N_19110);
nor U19330 (N_19330,N_19154,N_19149);
xnor U19331 (N_19331,N_19117,N_19188);
xor U19332 (N_19332,N_19143,N_19072);
and U19333 (N_19333,N_19048,N_19195);
xnor U19334 (N_19334,N_19021,N_19109);
nor U19335 (N_19335,N_19073,N_19034);
xor U19336 (N_19336,N_19144,N_19083);
or U19337 (N_19337,N_19003,N_19005);
or U19338 (N_19338,N_19198,N_19155);
and U19339 (N_19339,N_19044,N_19061);
nand U19340 (N_19340,N_19090,N_19061);
nor U19341 (N_19341,N_19110,N_19162);
nor U19342 (N_19342,N_19035,N_19070);
and U19343 (N_19343,N_19187,N_19117);
and U19344 (N_19344,N_19138,N_19165);
and U19345 (N_19345,N_19192,N_19101);
nor U19346 (N_19346,N_19148,N_19024);
nor U19347 (N_19347,N_19002,N_19197);
and U19348 (N_19348,N_19052,N_19156);
nand U19349 (N_19349,N_19155,N_19101);
nor U19350 (N_19350,N_19072,N_19017);
or U19351 (N_19351,N_19021,N_19180);
nand U19352 (N_19352,N_19026,N_19195);
xnor U19353 (N_19353,N_19075,N_19061);
xor U19354 (N_19354,N_19054,N_19127);
or U19355 (N_19355,N_19018,N_19194);
and U19356 (N_19356,N_19128,N_19029);
nand U19357 (N_19357,N_19169,N_19096);
and U19358 (N_19358,N_19074,N_19049);
and U19359 (N_19359,N_19184,N_19190);
nand U19360 (N_19360,N_19075,N_19040);
and U19361 (N_19361,N_19191,N_19153);
nand U19362 (N_19362,N_19010,N_19122);
or U19363 (N_19363,N_19070,N_19156);
and U19364 (N_19364,N_19046,N_19060);
nor U19365 (N_19365,N_19051,N_19030);
nand U19366 (N_19366,N_19153,N_19076);
nand U19367 (N_19367,N_19120,N_19059);
nand U19368 (N_19368,N_19067,N_19172);
nor U19369 (N_19369,N_19153,N_19089);
nand U19370 (N_19370,N_19180,N_19111);
and U19371 (N_19371,N_19044,N_19110);
or U19372 (N_19372,N_19044,N_19113);
and U19373 (N_19373,N_19087,N_19086);
or U19374 (N_19374,N_19197,N_19044);
nor U19375 (N_19375,N_19093,N_19120);
or U19376 (N_19376,N_19081,N_19156);
xnor U19377 (N_19377,N_19025,N_19037);
and U19378 (N_19378,N_19130,N_19120);
nand U19379 (N_19379,N_19174,N_19065);
nor U19380 (N_19380,N_19188,N_19109);
and U19381 (N_19381,N_19070,N_19130);
nand U19382 (N_19382,N_19010,N_19021);
or U19383 (N_19383,N_19178,N_19175);
nand U19384 (N_19384,N_19150,N_19062);
nand U19385 (N_19385,N_19137,N_19035);
and U19386 (N_19386,N_19052,N_19178);
nand U19387 (N_19387,N_19088,N_19099);
xor U19388 (N_19388,N_19147,N_19019);
or U19389 (N_19389,N_19072,N_19069);
xnor U19390 (N_19390,N_19091,N_19141);
xor U19391 (N_19391,N_19139,N_19111);
or U19392 (N_19392,N_19196,N_19008);
and U19393 (N_19393,N_19021,N_19149);
nor U19394 (N_19394,N_19002,N_19113);
and U19395 (N_19395,N_19001,N_19130);
and U19396 (N_19396,N_19170,N_19067);
nand U19397 (N_19397,N_19179,N_19198);
nor U19398 (N_19398,N_19016,N_19014);
xnor U19399 (N_19399,N_19157,N_19110);
nor U19400 (N_19400,N_19375,N_19246);
nand U19401 (N_19401,N_19309,N_19254);
or U19402 (N_19402,N_19312,N_19392);
and U19403 (N_19403,N_19331,N_19255);
and U19404 (N_19404,N_19295,N_19276);
nor U19405 (N_19405,N_19332,N_19274);
nand U19406 (N_19406,N_19279,N_19310);
xnor U19407 (N_19407,N_19380,N_19341);
nor U19408 (N_19408,N_19225,N_19318);
nand U19409 (N_19409,N_19371,N_19241);
or U19410 (N_19410,N_19242,N_19352);
nor U19411 (N_19411,N_19298,N_19201);
nor U19412 (N_19412,N_19303,N_19258);
nand U19413 (N_19413,N_19206,N_19278);
nor U19414 (N_19414,N_19243,N_19395);
and U19415 (N_19415,N_19337,N_19256);
xor U19416 (N_19416,N_19347,N_19372);
or U19417 (N_19417,N_19314,N_19288);
nand U19418 (N_19418,N_19384,N_19245);
xnor U19419 (N_19419,N_19308,N_19270);
xor U19420 (N_19420,N_19263,N_19269);
nor U19421 (N_19421,N_19397,N_19284);
xnor U19422 (N_19422,N_19396,N_19369);
nand U19423 (N_19423,N_19348,N_19210);
nand U19424 (N_19424,N_19358,N_19239);
and U19425 (N_19425,N_19253,N_19232);
nand U19426 (N_19426,N_19217,N_19379);
xor U19427 (N_19427,N_19368,N_19351);
xor U19428 (N_19428,N_19214,N_19361);
nor U19429 (N_19429,N_19311,N_19363);
xor U19430 (N_19430,N_19299,N_19355);
xnor U19431 (N_19431,N_19327,N_19229);
nand U19432 (N_19432,N_19207,N_19302);
and U19433 (N_19433,N_19297,N_19307);
xor U19434 (N_19434,N_19359,N_19356);
xnor U19435 (N_19435,N_19353,N_19261);
nor U19436 (N_19436,N_19399,N_19296);
xor U19437 (N_19437,N_19320,N_19285);
and U19438 (N_19438,N_19280,N_19268);
or U19439 (N_19439,N_19224,N_19326);
and U19440 (N_19440,N_19293,N_19215);
nor U19441 (N_19441,N_19267,N_19333);
nor U19442 (N_19442,N_19281,N_19360);
nor U19443 (N_19443,N_19354,N_19202);
and U19444 (N_19444,N_19248,N_19230);
or U19445 (N_19445,N_19389,N_19370);
or U19446 (N_19446,N_19286,N_19291);
or U19447 (N_19447,N_19329,N_19391);
or U19448 (N_19448,N_19235,N_19316);
or U19449 (N_19449,N_19367,N_19237);
or U19450 (N_19450,N_19381,N_19234);
nor U19451 (N_19451,N_19238,N_19287);
nand U19452 (N_19452,N_19350,N_19301);
and U19453 (N_19453,N_19273,N_19342);
and U19454 (N_19454,N_19374,N_19240);
nor U19455 (N_19455,N_19362,N_19349);
nor U19456 (N_19456,N_19218,N_19227);
nand U19457 (N_19457,N_19305,N_19275);
or U19458 (N_19458,N_19338,N_19244);
or U19459 (N_19459,N_19364,N_19213);
or U19460 (N_19460,N_19336,N_19300);
nand U19461 (N_19461,N_19339,N_19211);
xor U19462 (N_19462,N_19335,N_19265);
xor U19463 (N_19463,N_19344,N_19260);
nor U19464 (N_19464,N_19304,N_19387);
nor U19465 (N_19465,N_19233,N_19283);
and U19466 (N_19466,N_19306,N_19289);
xnor U19467 (N_19467,N_19220,N_19203);
and U19468 (N_19468,N_19266,N_19200);
nand U19469 (N_19469,N_19334,N_19208);
nand U19470 (N_19470,N_19290,N_19385);
or U19471 (N_19471,N_19315,N_19328);
nand U19472 (N_19472,N_19377,N_19272);
or U19473 (N_19473,N_19259,N_19393);
and U19474 (N_19474,N_19282,N_19346);
or U19475 (N_19475,N_19228,N_19236);
and U19476 (N_19476,N_19204,N_19271);
xnor U19477 (N_19477,N_19257,N_19345);
or U19478 (N_19478,N_19249,N_19205);
or U19479 (N_19479,N_19366,N_19330);
xnor U19480 (N_19480,N_19231,N_19365);
xnor U19481 (N_19481,N_19398,N_19394);
nor U19482 (N_19482,N_19388,N_19212);
or U19483 (N_19483,N_19390,N_19219);
and U19484 (N_19484,N_19292,N_19386);
and U19485 (N_19485,N_19264,N_19343);
or U19486 (N_19486,N_19382,N_19322);
nor U19487 (N_19487,N_19324,N_19247);
nand U19488 (N_19488,N_19373,N_19319);
nand U19489 (N_19489,N_19262,N_19340);
xnor U19490 (N_19490,N_19323,N_19277);
or U19491 (N_19491,N_19376,N_19252);
or U19492 (N_19492,N_19383,N_19313);
and U19493 (N_19493,N_19321,N_19317);
nand U19494 (N_19494,N_19222,N_19251);
nor U19495 (N_19495,N_19250,N_19325);
nor U19496 (N_19496,N_19223,N_19294);
or U19497 (N_19497,N_19378,N_19216);
and U19498 (N_19498,N_19221,N_19226);
nand U19499 (N_19499,N_19357,N_19209);
or U19500 (N_19500,N_19385,N_19314);
nand U19501 (N_19501,N_19240,N_19309);
and U19502 (N_19502,N_19383,N_19213);
or U19503 (N_19503,N_19373,N_19259);
and U19504 (N_19504,N_19388,N_19204);
xnor U19505 (N_19505,N_19292,N_19217);
xnor U19506 (N_19506,N_19347,N_19240);
nand U19507 (N_19507,N_19268,N_19362);
or U19508 (N_19508,N_19354,N_19252);
or U19509 (N_19509,N_19365,N_19271);
nor U19510 (N_19510,N_19229,N_19231);
or U19511 (N_19511,N_19268,N_19391);
or U19512 (N_19512,N_19355,N_19374);
and U19513 (N_19513,N_19307,N_19238);
xor U19514 (N_19514,N_19203,N_19206);
or U19515 (N_19515,N_19252,N_19316);
nor U19516 (N_19516,N_19364,N_19334);
or U19517 (N_19517,N_19255,N_19225);
nand U19518 (N_19518,N_19251,N_19377);
nor U19519 (N_19519,N_19240,N_19210);
xnor U19520 (N_19520,N_19259,N_19360);
or U19521 (N_19521,N_19227,N_19310);
and U19522 (N_19522,N_19390,N_19290);
nand U19523 (N_19523,N_19341,N_19326);
nor U19524 (N_19524,N_19201,N_19305);
or U19525 (N_19525,N_19259,N_19279);
or U19526 (N_19526,N_19379,N_19283);
xor U19527 (N_19527,N_19225,N_19358);
and U19528 (N_19528,N_19318,N_19204);
xnor U19529 (N_19529,N_19324,N_19311);
or U19530 (N_19530,N_19242,N_19280);
nor U19531 (N_19531,N_19232,N_19338);
nand U19532 (N_19532,N_19302,N_19273);
nand U19533 (N_19533,N_19377,N_19322);
nor U19534 (N_19534,N_19249,N_19280);
nor U19535 (N_19535,N_19291,N_19225);
nor U19536 (N_19536,N_19356,N_19257);
or U19537 (N_19537,N_19316,N_19364);
nor U19538 (N_19538,N_19377,N_19210);
and U19539 (N_19539,N_19394,N_19267);
nand U19540 (N_19540,N_19359,N_19220);
and U19541 (N_19541,N_19320,N_19202);
nand U19542 (N_19542,N_19232,N_19259);
xor U19543 (N_19543,N_19254,N_19384);
and U19544 (N_19544,N_19350,N_19295);
or U19545 (N_19545,N_19260,N_19220);
or U19546 (N_19546,N_19348,N_19309);
nor U19547 (N_19547,N_19329,N_19245);
xnor U19548 (N_19548,N_19279,N_19224);
nand U19549 (N_19549,N_19337,N_19227);
nor U19550 (N_19550,N_19207,N_19282);
xnor U19551 (N_19551,N_19330,N_19342);
or U19552 (N_19552,N_19331,N_19392);
nand U19553 (N_19553,N_19285,N_19392);
xnor U19554 (N_19554,N_19379,N_19227);
xnor U19555 (N_19555,N_19266,N_19217);
xnor U19556 (N_19556,N_19396,N_19249);
nand U19557 (N_19557,N_19218,N_19241);
xnor U19558 (N_19558,N_19348,N_19295);
xor U19559 (N_19559,N_19390,N_19380);
or U19560 (N_19560,N_19213,N_19263);
or U19561 (N_19561,N_19298,N_19241);
or U19562 (N_19562,N_19344,N_19396);
nor U19563 (N_19563,N_19201,N_19293);
nor U19564 (N_19564,N_19322,N_19292);
xor U19565 (N_19565,N_19371,N_19373);
nor U19566 (N_19566,N_19224,N_19312);
nand U19567 (N_19567,N_19336,N_19302);
or U19568 (N_19568,N_19392,N_19399);
or U19569 (N_19569,N_19227,N_19312);
and U19570 (N_19570,N_19222,N_19361);
xor U19571 (N_19571,N_19312,N_19219);
or U19572 (N_19572,N_19213,N_19205);
xnor U19573 (N_19573,N_19281,N_19354);
nor U19574 (N_19574,N_19387,N_19388);
nor U19575 (N_19575,N_19299,N_19357);
and U19576 (N_19576,N_19371,N_19303);
nor U19577 (N_19577,N_19212,N_19392);
nor U19578 (N_19578,N_19353,N_19345);
xnor U19579 (N_19579,N_19335,N_19369);
nand U19580 (N_19580,N_19349,N_19205);
and U19581 (N_19581,N_19357,N_19358);
nand U19582 (N_19582,N_19289,N_19297);
or U19583 (N_19583,N_19387,N_19390);
nor U19584 (N_19584,N_19387,N_19222);
or U19585 (N_19585,N_19354,N_19261);
nor U19586 (N_19586,N_19212,N_19234);
or U19587 (N_19587,N_19359,N_19316);
xor U19588 (N_19588,N_19217,N_19368);
xnor U19589 (N_19589,N_19293,N_19362);
nand U19590 (N_19590,N_19213,N_19221);
xnor U19591 (N_19591,N_19226,N_19278);
and U19592 (N_19592,N_19255,N_19200);
xor U19593 (N_19593,N_19346,N_19381);
or U19594 (N_19594,N_19235,N_19268);
nand U19595 (N_19595,N_19291,N_19369);
or U19596 (N_19596,N_19365,N_19204);
or U19597 (N_19597,N_19214,N_19298);
and U19598 (N_19598,N_19399,N_19360);
and U19599 (N_19599,N_19323,N_19228);
and U19600 (N_19600,N_19418,N_19464);
or U19601 (N_19601,N_19560,N_19448);
or U19602 (N_19602,N_19439,N_19518);
nand U19603 (N_19603,N_19444,N_19477);
and U19604 (N_19604,N_19409,N_19534);
or U19605 (N_19605,N_19451,N_19524);
nand U19606 (N_19606,N_19580,N_19460);
and U19607 (N_19607,N_19501,N_19581);
nor U19608 (N_19608,N_19592,N_19566);
or U19609 (N_19609,N_19495,N_19473);
nor U19610 (N_19610,N_19480,N_19453);
xor U19611 (N_19611,N_19508,N_19487);
nor U19612 (N_19612,N_19526,N_19541);
xor U19613 (N_19613,N_19522,N_19571);
xor U19614 (N_19614,N_19591,N_19491);
nand U19615 (N_19615,N_19520,N_19567);
nand U19616 (N_19616,N_19528,N_19457);
nand U19617 (N_19617,N_19586,N_19596);
or U19618 (N_19618,N_19481,N_19552);
nand U19619 (N_19619,N_19406,N_19450);
and U19620 (N_19620,N_19465,N_19462);
xor U19621 (N_19621,N_19499,N_19562);
or U19622 (N_19622,N_19527,N_19594);
xor U19623 (N_19623,N_19437,N_19543);
and U19624 (N_19624,N_19428,N_19443);
nand U19625 (N_19625,N_19503,N_19532);
and U19626 (N_19626,N_19599,N_19576);
or U19627 (N_19627,N_19589,N_19430);
and U19628 (N_19628,N_19549,N_19420);
and U19629 (N_19629,N_19521,N_19459);
or U19630 (N_19630,N_19584,N_19400);
nand U19631 (N_19631,N_19598,N_19575);
and U19632 (N_19632,N_19490,N_19475);
nor U19633 (N_19633,N_19431,N_19429);
or U19634 (N_19634,N_19468,N_19425);
xor U19635 (N_19635,N_19569,N_19454);
nor U19636 (N_19636,N_19561,N_19514);
xor U19637 (N_19637,N_19590,N_19519);
or U19638 (N_19638,N_19433,N_19593);
nand U19639 (N_19639,N_19463,N_19531);
nor U19640 (N_19640,N_19414,N_19403);
and U19641 (N_19641,N_19492,N_19548);
xnor U19642 (N_19642,N_19578,N_19452);
xor U19643 (N_19643,N_19595,N_19563);
xnor U19644 (N_19644,N_19557,N_19408);
or U19645 (N_19645,N_19523,N_19556);
nor U19646 (N_19646,N_19427,N_19485);
nor U19647 (N_19647,N_19411,N_19506);
nand U19648 (N_19648,N_19479,N_19585);
or U19649 (N_19649,N_19547,N_19512);
or U19650 (N_19650,N_19441,N_19546);
nand U19651 (N_19651,N_19456,N_19401);
or U19652 (N_19652,N_19410,N_19505);
nor U19653 (N_19653,N_19516,N_19417);
and U19654 (N_19654,N_19407,N_19500);
nand U19655 (N_19655,N_19570,N_19517);
nand U19656 (N_19656,N_19436,N_19474);
nand U19657 (N_19657,N_19572,N_19419);
xor U19658 (N_19658,N_19486,N_19497);
nor U19659 (N_19659,N_19461,N_19402);
and U19660 (N_19660,N_19515,N_19542);
and U19661 (N_19661,N_19537,N_19536);
nand U19662 (N_19662,N_19488,N_19551);
xor U19663 (N_19663,N_19447,N_19413);
nor U19664 (N_19664,N_19513,N_19545);
and U19665 (N_19665,N_19559,N_19533);
xor U19666 (N_19666,N_19458,N_19434);
or U19667 (N_19667,N_19442,N_19525);
and U19668 (N_19668,N_19424,N_19511);
nor U19669 (N_19669,N_19412,N_19432);
and U19670 (N_19670,N_19577,N_19482);
nor U19671 (N_19671,N_19493,N_19574);
nand U19672 (N_19672,N_19573,N_19404);
xnor U19673 (N_19673,N_19540,N_19466);
nand U19674 (N_19674,N_19416,N_19455);
nand U19675 (N_19675,N_19483,N_19494);
and U19676 (N_19676,N_19449,N_19415);
or U19677 (N_19677,N_19467,N_19564);
nand U19678 (N_19678,N_19509,N_19507);
nand U19679 (N_19679,N_19446,N_19553);
nor U19680 (N_19680,N_19568,N_19469);
and U19681 (N_19681,N_19535,N_19472);
or U19682 (N_19682,N_19440,N_19587);
xnor U19683 (N_19683,N_19496,N_19529);
or U19684 (N_19684,N_19558,N_19405);
nor U19685 (N_19685,N_19445,N_19422);
nand U19686 (N_19686,N_19583,N_19554);
nor U19687 (N_19687,N_19565,N_19582);
xor U19688 (N_19688,N_19421,N_19489);
or U19689 (N_19689,N_19502,N_19435);
xnor U19690 (N_19690,N_19423,N_19478);
nand U19691 (N_19691,N_19438,N_19544);
or U19692 (N_19692,N_19539,N_19579);
and U19693 (N_19693,N_19588,N_19484);
nand U19694 (N_19694,N_19538,N_19426);
and U19695 (N_19695,N_19476,N_19550);
and U19696 (N_19696,N_19504,N_19530);
xnor U19697 (N_19697,N_19498,N_19597);
nand U19698 (N_19698,N_19555,N_19471);
xor U19699 (N_19699,N_19470,N_19510);
or U19700 (N_19700,N_19457,N_19530);
nor U19701 (N_19701,N_19574,N_19579);
and U19702 (N_19702,N_19449,N_19537);
xnor U19703 (N_19703,N_19512,N_19502);
nor U19704 (N_19704,N_19537,N_19551);
or U19705 (N_19705,N_19529,N_19498);
xnor U19706 (N_19706,N_19501,N_19510);
nor U19707 (N_19707,N_19401,N_19574);
or U19708 (N_19708,N_19553,N_19489);
xor U19709 (N_19709,N_19589,N_19466);
nand U19710 (N_19710,N_19465,N_19404);
xor U19711 (N_19711,N_19592,N_19405);
or U19712 (N_19712,N_19465,N_19553);
nor U19713 (N_19713,N_19446,N_19556);
xnor U19714 (N_19714,N_19514,N_19556);
nand U19715 (N_19715,N_19514,N_19565);
nand U19716 (N_19716,N_19598,N_19552);
or U19717 (N_19717,N_19572,N_19422);
or U19718 (N_19718,N_19475,N_19535);
nand U19719 (N_19719,N_19563,N_19562);
or U19720 (N_19720,N_19472,N_19563);
xor U19721 (N_19721,N_19513,N_19479);
xnor U19722 (N_19722,N_19537,N_19459);
and U19723 (N_19723,N_19568,N_19434);
nor U19724 (N_19724,N_19508,N_19546);
xnor U19725 (N_19725,N_19414,N_19540);
nor U19726 (N_19726,N_19517,N_19405);
xor U19727 (N_19727,N_19433,N_19556);
nor U19728 (N_19728,N_19516,N_19597);
and U19729 (N_19729,N_19430,N_19417);
nor U19730 (N_19730,N_19482,N_19458);
or U19731 (N_19731,N_19502,N_19440);
or U19732 (N_19732,N_19488,N_19413);
nor U19733 (N_19733,N_19523,N_19445);
and U19734 (N_19734,N_19400,N_19433);
and U19735 (N_19735,N_19417,N_19536);
nor U19736 (N_19736,N_19427,N_19497);
and U19737 (N_19737,N_19594,N_19513);
and U19738 (N_19738,N_19541,N_19536);
and U19739 (N_19739,N_19586,N_19540);
or U19740 (N_19740,N_19513,N_19536);
and U19741 (N_19741,N_19451,N_19582);
nor U19742 (N_19742,N_19460,N_19586);
nand U19743 (N_19743,N_19549,N_19557);
xnor U19744 (N_19744,N_19407,N_19436);
and U19745 (N_19745,N_19521,N_19584);
xor U19746 (N_19746,N_19418,N_19447);
and U19747 (N_19747,N_19562,N_19482);
or U19748 (N_19748,N_19526,N_19476);
and U19749 (N_19749,N_19404,N_19481);
xor U19750 (N_19750,N_19510,N_19438);
nor U19751 (N_19751,N_19590,N_19483);
xnor U19752 (N_19752,N_19567,N_19552);
or U19753 (N_19753,N_19469,N_19465);
nor U19754 (N_19754,N_19427,N_19402);
xnor U19755 (N_19755,N_19503,N_19400);
and U19756 (N_19756,N_19456,N_19533);
nor U19757 (N_19757,N_19503,N_19428);
nand U19758 (N_19758,N_19418,N_19566);
nor U19759 (N_19759,N_19518,N_19419);
xnor U19760 (N_19760,N_19400,N_19539);
nor U19761 (N_19761,N_19487,N_19496);
xor U19762 (N_19762,N_19467,N_19494);
and U19763 (N_19763,N_19536,N_19563);
or U19764 (N_19764,N_19530,N_19589);
or U19765 (N_19765,N_19574,N_19441);
nor U19766 (N_19766,N_19531,N_19427);
xnor U19767 (N_19767,N_19418,N_19554);
nand U19768 (N_19768,N_19523,N_19570);
and U19769 (N_19769,N_19563,N_19430);
nand U19770 (N_19770,N_19404,N_19467);
or U19771 (N_19771,N_19412,N_19475);
nand U19772 (N_19772,N_19597,N_19570);
nand U19773 (N_19773,N_19595,N_19508);
nor U19774 (N_19774,N_19449,N_19591);
or U19775 (N_19775,N_19557,N_19481);
and U19776 (N_19776,N_19531,N_19533);
nor U19777 (N_19777,N_19488,N_19467);
nor U19778 (N_19778,N_19535,N_19500);
nor U19779 (N_19779,N_19571,N_19437);
nand U19780 (N_19780,N_19543,N_19597);
nor U19781 (N_19781,N_19469,N_19442);
xnor U19782 (N_19782,N_19586,N_19529);
xor U19783 (N_19783,N_19523,N_19548);
and U19784 (N_19784,N_19441,N_19436);
and U19785 (N_19785,N_19495,N_19413);
and U19786 (N_19786,N_19586,N_19512);
xor U19787 (N_19787,N_19507,N_19413);
xor U19788 (N_19788,N_19526,N_19438);
xor U19789 (N_19789,N_19593,N_19549);
nand U19790 (N_19790,N_19577,N_19521);
or U19791 (N_19791,N_19461,N_19463);
nand U19792 (N_19792,N_19416,N_19501);
nand U19793 (N_19793,N_19478,N_19450);
or U19794 (N_19794,N_19529,N_19576);
or U19795 (N_19795,N_19439,N_19467);
xnor U19796 (N_19796,N_19560,N_19490);
or U19797 (N_19797,N_19576,N_19537);
nor U19798 (N_19798,N_19435,N_19539);
nand U19799 (N_19799,N_19561,N_19443);
nand U19800 (N_19800,N_19732,N_19749);
nand U19801 (N_19801,N_19683,N_19662);
nor U19802 (N_19802,N_19611,N_19601);
and U19803 (N_19803,N_19633,N_19747);
and U19804 (N_19804,N_19628,N_19769);
nand U19805 (N_19805,N_19705,N_19794);
nor U19806 (N_19806,N_19674,N_19698);
nor U19807 (N_19807,N_19721,N_19695);
nand U19808 (N_19808,N_19709,N_19603);
or U19809 (N_19809,N_19667,N_19750);
nor U19810 (N_19810,N_19668,N_19745);
and U19811 (N_19811,N_19651,N_19771);
nor U19812 (N_19812,N_19758,N_19743);
xor U19813 (N_19813,N_19626,N_19620);
nand U19814 (N_19814,N_19707,N_19708);
xnor U19815 (N_19815,N_19661,N_19751);
xnor U19816 (N_19816,N_19756,N_19777);
and U19817 (N_19817,N_19609,N_19676);
and U19818 (N_19818,N_19710,N_19605);
nand U19819 (N_19819,N_19752,N_19635);
or U19820 (N_19820,N_19785,N_19740);
nand U19821 (N_19821,N_19627,N_19711);
or U19822 (N_19822,N_19730,N_19697);
and U19823 (N_19823,N_19719,N_19658);
or U19824 (N_19824,N_19770,N_19700);
nor U19825 (N_19825,N_19656,N_19786);
and U19826 (N_19826,N_19696,N_19655);
or U19827 (N_19827,N_19755,N_19727);
nor U19828 (N_19828,N_19704,N_19797);
or U19829 (N_19829,N_19670,N_19693);
nor U19830 (N_19830,N_19678,N_19671);
nand U19831 (N_19831,N_19681,N_19734);
xor U19832 (N_19832,N_19746,N_19614);
and U19833 (N_19833,N_19766,N_19684);
and U19834 (N_19834,N_19741,N_19663);
or U19835 (N_19835,N_19629,N_19692);
or U19836 (N_19836,N_19619,N_19694);
xnor U19837 (N_19837,N_19660,N_19604);
nor U19838 (N_19838,N_19654,N_19716);
nand U19839 (N_19839,N_19636,N_19653);
and U19840 (N_19840,N_19677,N_19788);
xnor U19841 (N_19841,N_19600,N_19647);
or U19842 (N_19842,N_19613,N_19648);
xor U19843 (N_19843,N_19650,N_19793);
or U19844 (N_19844,N_19720,N_19713);
and U19845 (N_19845,N_19608,N_19634);
or U19846 (N_19846,N_19682,N_19623);
nor U19847 (N_19847,N_19624,N_19606);
xnor U19848 (N_19848,N_19737,N_19642);
nor U19849 (N_19849,N_19767,N_19691);
or U19850 (N_19850,N_19726,N_19754);
and U19851 (N_19851,N_19657,N_19773);
nand U19852 (N_19852,N_19665,N_19679);
nand U19853 (N_19853,N_19744,N_19664);
or U19854 (N_19854,N_19798,N_19715);
and U19855 (N_19855,N_19783,N_19618);
nand U19856 (N_19856,N_19718,N_19617);
or U19857 (N_19857,N_19729,N_19612);
and U19858 (N_19858,N_19790,N_19622);
and U19859 (N_19859,N_19703,N_19637);
xor U19860 (N_19860,N_19687,N_19640);
or U19861 (N_19861,N_19759,N_19760);
or U19862 (N_19862,N_19779,N_19616);
or U19863 (N_19863,N_19602,N_19776);
nand U19864 (N_19864,N_19725,N_19645);
nand U19865 (N_19865,N_19625,N_19630);
nor U19866 (N_19866,N_19717,N_19736);
xnor U19867 (N_19867,N_19652,N_19791);
xnor U19868 (N_19868,N_19762,N_19761);
nor U19869 (N_19869,N_19792,N_19675);
nor U19870 (N_19870,N_19795,N_19796);
or U19871 (N_19871,N_19780,N_19772);
xnor U19872 (N_19872,N_19673,N_19757);
nor U19873 (N_19873,N_19739,N_19778);
or U19874 (N_19874,N_19702,N_19723);
xnor U19875 (N_19875,N_19753,N_19722);
or U19876 (N_19876,N_19643,N_19712);
nor U19877 (N_19877,N_19775,N_19659);
and U19878 (N_19878,N_19672,N_19666);
or U19879 (N_19879,N_19699,N_19669);
and U19880 (N_19880,N_19714,N_19686);
nand U19881 (N_19881,N_19685,N_19765);
nor U19882 (N_19882,N_19689,N_19631);
nand U19883 (N_19883,N_19644,N_19615);
nor U19884 (N_19884,N_19641,N_19632);
nand U19885 (N_19885,N_19774,N_19610);
or U19886 (N_19886,N_19781,N_19784);
xnor U19887 (N_19887,N_19639,N_19706);
or U19888 (N_19888,N_19621,N_19638);
nand U19889 (N_19889,N_19735,N_19607);
nor U19890 (N_19890,N_19733,N_19724);
and U19891 (N_19891,N_19768,N_19731);
nor U19892 (N_19892,N_19680,N_19690);
nor U19893 (N_19893,N_19799,N_19763);
or U19894 (N_19894,N_19688,N_19789);
and U19895 (N_19895,N_19748,N_19649);
or U19896 (N_19896,N_19782,N_19646);
nand U19897 (N_19897,N_19738,N_19728);
xnor U19898 (N_19898,N_19742,N_19764);
nand U19899 (N_19899,N_19701,N_19787);
xnor U19900 (N_19900,N_19703,N_19778);
and U19901 (N_19901,N_19749,N_19713);
xnor U19902 (N_19902,N_19797,N_19606);
nor U19903 (N_19903,N_19620,N_19642);
nor U19904 (N_19904,N_19763,N_19764);
and U19905 (N_19905,N_19784,N_19610);
or U19906 (N_19906,N_19675,N_19706);
xor U19907 (N_19907,N_19736,N_19769);
nor U19908 (N_19908,N_19604,N_19735);
nand U19909 (N_19909,N_19613,N_19759);
xnor U19910 (N_19910,N_19792,N_19713);
nor U19911 (N_19911,N_19728,N_19797);
xnor U19912 (N_19912,N_19641,N_19758);
and U19913 (N_19913,N_19639,N_19783);
nor U19914 (N_19914,N_19725,N_19608);
nor U19915 (N_19915,N_19663,N_19681);
nand U19916 (N_19916,N_19644,N_19719);
xnor U19917 (N_19917,N_19791,N_19650);
xor U19918 (N_19918,N_19775,N_19643);
and U19919 (N_19919,N_19612,N_19775);
nand U19920 (N_19920,N_19784,N_19765);
or U19921 (N_19921,N_19740,N_19675);
xnor U19922 (N_19922,N_19622,N_19621);
nand U19923 (N_19923,N_19754,N_19752);
nand U19924 (N_19924,N_19766,N_19612);
xnor U19925 (N_19925,N_19618,N_19748);
nor U19926 (N_19926,N_19752,N_19776);
nand U19927 (N_19927,N_19613,N_19610);
nor U19928 (N_19928,N_19735,N_19728);
and U19929 (N_19929,N_19674,N_19777);
or U19930 (N_19930,N_19665,N_19720);
nand U19931 (N_19931,N_19673,N_19615);
or U19932 (N_19932,N_19725,N_19614);
xnor U19933 (N_19933,N_19634,N_19644);
or U19934 (N_19934,N_19679,N_19799);
nand U19935 (N_19935,N_19735,N_19697);
nor U19936 (N_19936,N_19620,N_19780);
or U19937 (N_19937,N_19782,N_19666);
nor U19938 (N_19938,N_19774,N_19705);
xor U19939 (N_19939,N_19637,N_19664);
xnor U19940 (N_19940,N_19602,N_19604);
nand U19941 (N_19941,N_19686,N_19761);
nor U19942 (N_19942,N_19783,N_19616);
nand U19943 (N_19943,N_19791,N_19705);
xor U19944 (N_19944,N_19661,N_19635);
nor U19945 (N_19945,N_19742,N_19758);
xor U19946 (N_19946,N_19613,N_19702);
and U19947 (N_19947,N_19653,N_19789);
xor U19948 (N_19948,N_19686,N_19645);
nor U19949 (N_19949,N_19649,N_19671);
nand U19950 (N_19950,N_19686,N_19692);
nor U19951 (N_19951,N_19659,N_19738);
nor U19952 (N_19952,N_19650,N_19624);
nor U19953 (N_19953,N_19787,N_19731);
and U19954 (N_19954,N_19635,N_19796);
nand U19955 (N_19955,N_19777,N_19608);
and U19956 (N_19956,N_19655,N_19609);
and U19957 (N_19957,N_19739,N_19742);
nor U19958 (N_19958,N_19795,N_19635);
xor U19959 (N_19959,N_19706,N_19714);
and U19960 (N_19960,N_19609,N_19664);
xnor U19961 (N_19961,N_19672,N_19713);
xor U19962 (N_19962,N_19797,N_19691);
xor U19963 (N_19963,N_19773,N_19687);
nand U19964 (N_19964,N_19693,N_19629);
xnor U19965 (N_19965,N_19669,N_19782);
nand U19966 (N_19966,N_19767,N_19792);
xor U19967 (N_19967,N_19696,N_19744);
and U19968 (N_19968,N_19783,N_19725);
or U19969 (N_19969,N_19722,N_19651);
or U19970 (N_19970,N_19692,N_19642);
xor U19971 (N_19971,N_19702,N_19781);
nor U19972 (N_19972,N_19792,N_19718);
and U19973 (N_19973,N_19687,N_19677);
xnor U19974 (N_19974,N_19734,N_19626);
nor U19975 (N_19975,N_19725,N_19715);
or U19976 (N_19976,N_19601,N_19605);
or U19977 (N_19977,N_19770,N_19723);
nor U19978 (N_19978,N_19647,N_19787);
xor U19979 (N_19979,N_19646,N_19799);
nand U19980 (N_19980,N_19772,N_19768);
or U19981 (N_19981,N_19644,N_19621);
nand U19982 (N_19982,N_19601,N_19620);
or U19983 (N_19983,N_19684,N_19644);
xnor U19984 (N_19984,N_19755,N_19643);
and U19985 (N_19985,N_19686,N_19608);
nor U19986 (N_19986,N_19616,N_19670);
nor U19987 (N_19987,N_19658,N_19648);
or U19988 (N_19988,N_19623,N_19697);
nand U19989 (N_19989,N_19674,N_19732);
nand U19990 (N_19990,N_19727,N_19711);
nor U19991 (N_19991,N_19711,N_19754);
or U19992 (N_19992,N_19720,N_19751);
or U19993 (N_19993,N_19669,N_19698);
xor U19994 (N_19994,N_19600,N_19678);
nor U19995 (N_19995,N_19618,N_19605);
or U19996 (N_19996,N_19741,N_19624);
nand U19997 (N_19997,N_19693,N_19720);
xor U19998 (N_19998,N_19752,N_19641);
nand U19999 (N_19999,N_19667,N_19751);
nor UO_0 (O_0,N_19849,N_19941);
nand UO_1 (O_1,N_19850,N_19863);
or UO_2 (O_2,N_19883,N_19948);
nor UO_3 (O_3,N_19989,N_19930);
nand UO_4 (O_4,N_19890,N_19981);
and UO_5 (O_5,N_19983,N_19834);
and UO_6 (O_6,N_19928,N_19964);
and UO_7 (O_7,N_19996,N_19902);
nor UO_8 (O_8,N_19921,N_19975);
and UO_9 (O_9,N_19829,N_19841);
or UO_10 (O_10,N_19857,N_19959);
xnor UO_11 (O_11,N_19917,N_19876);
nand UO_12 (O_12,N_19873,N_19938);
nor UO_13 (O_13,N_19925,N_19889);
nand UO_14 (O_14,N_19808,N_19820);
and UO_15 (O_15,N_19960,N_19985);
xnor UO_16 (O_16,N_19991,N_19942);
nand UO_17 (O_17,N_19828,N_19832);
nor UO_18 (O_18,N_19887,N_19897);
or UO_19 (O_19,N_19817,N_19931);
xnor UO_20 (O_20,N_19997,N_19870);
nand UO_21 (O_21,N_19842,N_19864);
or UO_22 (O_22,N_19944,N_19804);
and UO_23 (O_23,N_19911,N_19818);
and UO_24 (O_24,N_19933,N_19967);
nand UO_25 (O_25,N_19935,N_19845);
xnor UO_26 (O_26,N_19939,N_19812);
and UO_27 (O_27,N_19823,N_19894);
nor UO_28 (O_28,N_19885,N_19888);
nand UO_29 (O_29,N_19958,N_19833);
nand UO_30 (O_30,N_19977,N_19801);
nand UO_31 (O_31,N_19908,N_19835);
or UO_32 (O_32,N_19811,N_19910);
or UO_33 (O_33,N_19966,N_19866);
nor UO_34 (O_34,N_19836,N_19970);
nand UO_35 (O_35,N_19956,N_19816);
xor UO_36 (O_36,N_19871,N_19974);
xor UO_37 (O_37,N_19809,N_19950);
nor UO_38 (O_38,N_19862,N_19874);
and UO_39 (O_39,N_19949,N_19893);
nor UO_40 (O_40,N_19813,N_19830);
or UO_41 (O_41,N_19877,N_19962);
nand UO_42 (O_42,N_19853,N_19847);
or UO_43 (O_43,N_19851,N_19838);
nand UO_44 (O_44,N_19969,N_19951);
nor UO_45 (O_45,N_19980,N_19856);
or UO_46 (O_46,N_19920,N_19892);
nand UO_47 (O_47,N_19802,N_19927);
nor UO_48 (O_48,N_19867,N_19819);
or UO_49 (O_49,N_19932,N_19971);
nor UO_50 (O_50,N_19831,N_19859);
nor UO_51 (O_51,N_19805,N_19900);
nand UO_52 (O_52,N_19840,N_19903);
nor UO_53 (O_53,N_19855,N_19872);
and UO_54 (O_54,N_19986,N_19993);
xnor UO_55 (O_55,N_19987,N_19963);
xnor UO_56 (O_56,N_19968,N_19940);
or UO_57 (O_57,N_19926,N_19976);
and UO_58 (O_58,N_19878,N_19946);
xnor UO_59 (O_59,N_19898,N_19848);
nand UO_60 (O_60,N_19806,N_19943);
or UO_61 (O_61,N_19965,N_19923);
or UO_62 (O_62,N_19879,N_19837);
and UO_63 (O_63,N_19899,N_19884);
nor UO_64 (O_64,N_19904,N_19839);
nand UO_65 (O_65,N_19922,N_19998);
xor UO_66 (O_66,N_19973,N_19881);
or UO_67 (O_67,N_19882,N_19843);
nand UO_68 (O_68,N_19852,N_19909);
nand UO_69 (O_69,N_19988,N_19982);
and UO_70 (O_70,N_19978,N_19961);
nor UO_71 (O_71,N_19995,N_19905);
nand UO_72 (O_72,N_19822,N_19957);
or UO_73 (O_73,N_19854,N_19844);
and UO_74 (O_74,N_19918,N_19929);
xor UO_75 (O_75,N_19992,N_19936);
nor UO_76 (O_76,N_19803,N_19947);
and UO_77 (O_77,N_19924,N_19846);
nand UO_78 (O_78,N_19821,N_19990);
and UO_79 (O_79,N_19875,N_19972);
nand UO_80 (O_80,N_19827,N_19999);
nor UO_81 (O_81,N_19861,N_19916);
or UO_82 (O_82,N_19886,N_19868);
xnor UO_83 (O_83,N_19814,N_19869);
nand UO_84 (O_84,N_19858,N_19979);
or UO_85 (O_85,N_19954,N_19895);
and UO_86 (O_86,N_19824,N_19953);
nor UO_87 (O_87,N_19906,N_19901);
nor UO_88 (O_88,N_19800,N_19934);
nand UO_89 (O_89,N_19915,N_19825);
xnor UO_90 (O_90,N_19914,N_19807);
xnor UO_91 (O_91,N_19912,N_19994);
xnor UO_92 (O_92,N_19815,N_19880);
nand UO_93 (O_93,N_19984,N_19913);
and UO_94 (O_94,N_19826,N_19860);
or UO_95 (O_95,N_19919,N_19937);
nand UO_96 (O_96,N_19896,N_19810);
and UO_97 (O_97,N_19891,N_19945);
and UO_98 (O_98,N_19907,N_19952);
xnor UO_99 (O_99,N_19865,N_19955);
nor UO_100 (O_100,N_19865,N_19954);
or UO_101 (O_101,N_19931,N_19964);
or UO_102 (O_102,N_19819,N_19888);
or UO_103 (O_103,N_19988,N_19882);
nand UO_104 (O_104,N_19955,N_19939);
or UO_105 (O_105,N_19957,N_19982);
nor UO_106 (O_106,N_19983,N_19837);
and UO_107 (O_107,N_19835,N_19911);
and UO_108 (O_108,N_19903,N_19989);
xor UO_109 (O_109,N_19907,N_19826);
xnor UO_110 (O_110,N_19986,N_19932);
or UO_111 (O_111,N_19920,N_19813);
or UO_112 (O_112,N_19832,N_19830);
nand UO_113 (O_113,N_19976,N_19858);
xnor UO_114 (O_114,N_19949,N_19812);
nand UO_115 (O_115,N_19862,N_19914);
nand UO_116 (O_116,N_19990,N_19827);
nand UO_117 (O_117,N_19850,N_19947);
nor UO_118 (O_118,N_19834,N_19871);
or UO_119 (O_119,N_19865,N_19842);
xnor UO_120 (O_120,N_19880,N_19968);
or UO_121 (O_121,N_19859,N_19926);
nand UO_122 (O_122,N_19899,N_19978);
nor UO_123 (O_123,N_19931,N_19958);
xnor UO_124 (O_124,N_19899,N_19807);
nand UO_125 (O_125,N_19885,N_19941);
nor UO_126 (O_126,N_19922,N_19819);
and UO_127 (O_127,N_19870,N_19842);
nand UO_128 (O_128,N_19865,N_19851);
or UO_129 (O_129,N_19973,N_19804);
nor UO_130 (O_130,N_19970,N_19810);
xnor UO_131 (O_131,N_19888,N_19983);
nand UO_132 (O_132,N_19878,N_19820);
nor UO_133 (O_133,N_19889,N_19837);
nand UO_134 (O_134,N_19891,N_19931);
nand UO_135 (O_135,N_19864,N_19965);
nor UO_136 (O_136,N_19909,N_19974);
or UO_137 (O_137,N_19888,N_19863);
nor UO_138 (O_138,N_19980,N_19839);
xor UO_139 (O_139,N_19930,N_19997);
xor UO_140 (O_140,N_19949,N_19927);
or UO_141 (O_141,N_19807,N_19923);
nor UO_142 (O_142,N_19825,N_19936);
or UO_143 (O_143,N_19993,N_19983);
xor UO_144 (O_144,N_19977,N_19826);
and UO_145 (O_145,N_19906,N_19879);
or UO_146 (O_146,N_19921,N_19909);
nor UO_147 (O_147,N_19878,N_19973);
nor UO_148 (O_148,N_19928,N_19833);
or UO_149 (O_149,N_19843,N_19973);
nand UO_150 (O_150,N_19974,N_19920);
and UO_151 (O_151,N_19872,N_19820);
or UO_152 (O_152,N_19957,N_19875);
nand UO_153 (O_153,N_19833,N_19861);
nor UO_154 (O_154,N_19896,N_19822);
xnor UO_155 (O_155,N_19880,N_19832);
and UO_156 (O_156,N_19930,N_19857);
or UO_157 (O_157,N_19964,N_19835);
xor UO_158 (O_158,N_19842,N_19951);
and UO_159 (O_159,N_19903,N_19810);
or UO_160 (O_160,N_19956,N_19970);
or UO_161 (O_161,N_19963,N_19813);
xnor UO_162 (O_162,N_19951,N_19805);
or UO_163 (O_163,N_19916,N_19975);
nand UO_164 (O_164,N_19953,N_19835);
and UO_165 (O_165,N_19969,N_19863);
nand UO_166 (O_166,N_19969,N_19994);
xor UO_167 (O_167,N_19969,N_19832);
and UO_168 (O_168,N_19950,N_19907);
nor UO_169 (O_169,N_19812,N_19948);
or UO_170 (O_170,N_19955,N_19837);
nand UO_171 (O_171,N_19968,N_19886);
nor UO_172 (O_172,N_19858,N_19962);
or UO_173 (O_173,N_19842,N_19944);
and UO_174 (O_174,N_19891,N_19930);
or UO_175 (O_175,N_19801,N_19878);
xor UO_176 (O_176,N_19942,N_19869);
and UO_177 (O_177,N_19957,N_19959);
and UO_178 (O_178,N_19982,N_19944);
xor UO_179 (O_179,N_19952,N_19923);
nand UO_180 (O_180,N_19927,N_19881);
or UO_181 (O_181,N_19946,N_19944);
or UO_182 (O_182,N_19951,N_19962);
and UO_183 (O_183,N_19948,N_19916);
nor UO_184 (O_184,N_19818,N_19985);
nor UO_185 (O_185,N_19898,N_19802);
or UO_186 (O_186,N_19881,N_19922);
and UO_187 (O_187,N_19969,N_19829);
or UO_188 (O_188,N_19972,N_19834);
nor UO_189 (O_189,N_19961,N_19895);
xnor UO_190 (O_190,N_19835,N_19868);
nand UO_191 (O_191,N_19805,N_19815);
nor UO_192 (O_192,N_19908,N_19985);
nand UO_193 (O_193,N_19816,N_19916);
xor UO_194 (O_194,N_19882,N_19811);
or UO_195 (O_195,N_19968,N_19975);
xnor UO_196 (O_196,N_19858,N_19852);
and UO_197 (O_197,N_19964,N_19924);
or UO_198 (O_198,N_19821,N_19993);
xor UO_199 (O_199,N_19923,N_19811);
nor UO_200 (O_200,N_19863,N_19975);
or UO_201 (O_201,N_19816,N_19844);
or UO_202 (O_202,N_19866,N_19962);
nor UO_203 (O_203,N_19807,N_19927);
nand UO_204 (O_204,N_19905,N_19886);
nor UO_205 (O_205,N_19985,N_19950);
and UO_206 (O_206,N_19812,N_19850);
nor UO_207 (O_207,N_19993,N_19845);
nor UO_208 (O_208,N_19986,N_19867);
or UO_209 (O_209,N_19993,N_19991);
nand UO_210 (O_210,N_19975,N_19873);
or UO_211 (O_211,N_19802,N_19922);
nand UO_212 (O_212,N_19965,N_19803);
xnor UO_213 (O_213,N_19929,N_19980);
nand UO_214 (O_214,N_19919,N_19902);
or UO_215 (O_215,N_19953,N_19812);
nor UO_216 (O_216,N_19997,N_19932);
xor UO_217 (O_217,N_19908,N_19910);
nand UO_218 (O_218,N_19951,N_19862);
nor UO_219 (O_219,N_19824,N_19962);
and UO_220 (O_220,N_19851,N_19886);
xnor UO_221 (O_221,N_19803,N_19969);
and UO_222 (O_222,N_19885,N_19954);
and UO_223 (O_223,N_19899,N_19972);
xnor UO_224 (O_224,N_19828,N_19998);
xnor UO_225 (O_225,N_19842,N_19857);
nand UO_226 (O_226,N_19921,N_19933);
and UO_227 (O_227,N_19865,N_19812);
nand UO_228 (O_228,N_19972,N_19864);
nand UO_229 (O_229,N_19881,N_19852);
xor UO_230 (O_230,N_19904,N_19977);
nor UO_231 (O_231,N_19983,N_19934);
nand UO_232 (O_232,N_19840,N_19833);
nor UO_233 (O_233,N_19932,N_19995);
nor UO_234 (O_234,N_19888,N_19880);
nor UO_235 (O_235,N_19800,N_19906);
xnor UO_236 (O_236,N_19943,N_19956);
xor UO_237 (O_237,N_19865,N_19809);
nor UO_238 (O_238,N_19842,N_19929);
or UO_239 (O_239,N_19930,N_19905);
nor UO_240 (O_240,N_19961,N_19886);
nand UO_241 (O_241,N_19963,N_19908);
and UO_242 (O_242,N_19978,N_19920);
and UO_243 (O_243,N_19991,N_19857);
nor UO_244 (O_244,N_19804,N_19942);
or UO_245 (O_245,N_19878,N_19999);
nor UO_246 (O_246,N_19887,N_19920);
or UO_247 (O_247,N_19810,N_19817);
and UO_248 (O_248,N_19874,N_19894);
nor UO_249 (O_249,N_19924,N_19999);
nand UO_250 (O_250,N_19883,N_19800);
nor UO_251 (O_251,N_19865,N_19846);
nand UO_252 (O_252,N_19823,N_19863);
or UO_253 (O_253,N_19893,N_19912);
or UO_254 (O_254,N_19883,N_19905);
xor UO_255 (O_255,N_19887,N_19867);
nand UO_256 (O_256,N_19878,N_19844);
xnor UO_257 (O_257,N_19866,N_19818);
nor UO_258 (O_258,N_19949,N_19807);
nand UO_259 (O_259,N_19875,N_19822);
and UO_260 (O_260,N_19972,N_19901);
xor UO_261 (O_261,N_19859,N_19937);
or UO_262 (O_262,N_19934,N_19856);
nand UO_263 (O_263,N_19846,N_19896);
xor UO_264 (O_264,N_19945,N_19913);
xnor UO_265 (O_265,N_19935,N_19968);
nor UO_266 (O_266,N_19873,N_19891);
nand UO_267 (O_267,N_19952,N_19848);
or UO_268 (O_268,N_19853,N_19992);
xnor UO_269 (O_269,N_19934,N_19892);
or UO_270 (O_270,N_19980,N_19941);
and UO_271 (O_271,N_19990,N_19801);
and UO_272 (O_272,N_19925,N_19934);
nor UO_273 (O_273,N_19895,N_19853);
and UO_274 (O_274,N_19897,N_19991);
nor UO_275 (O_275,N_19801,N_19936);
or UO_276 (O_276,N_19866,N_19811);
or UO_277 (O_277,N_19833,N_19874);
xor UO_278 (O_278,N_19867,N_19836);
nor UO_279 (O_279,N_19805,N_19909);
or UO_280 (O_280,N_19991,N_19895);
xnor UO_281 (O_281,N_19852,N_19916);
or UO_282 (O_282,N_19913,N_19818);
or UO_283 (O_283,N_19938,N_19985);
nand UO_284 (O_284,N_19941,N_19831);
xor UO_285 (O_285,N_19820,N_19910);
nor UO_286 (O_286,N_19977,N_19936);
nor UO_287 (O_287,N_19840,N_19950);
xor UO_288 (O_288,N_19974,N_19916);
xnor UO_289 (O_289,N_19969,N_19894);
or UO_290 (O_290,N_19971,N_19933);
nand UO_291 (O_291,N_19993,N_19931);
nor UO_292 (O_292,N_19906,N_19973);
and UO_293 (O_293,N_19826,N_19925);
or UO_294 (O_294,N_19823,N_19955);
xnor UO_295 (O_295,N_19806,N_19849);
nand UO_296 (O_296,N_19862,N_19898);
xor UO_297 (O_297,N_19831,N_19841);
and UO_298 (O_298,N_19850,N_19849);
and UO_299 (O_299,N_19854,N_19875);
or UO_300 (O_300,N_19948,N_19881);
or UO_301 (O_301,N_19848,N_19842);
and UO_302 (O_302,N_19950,N_19810);
xnor UO_303 (O_303,N_19962,N_19838);
nand UO_304 (O_304,N_19889,N_19979);
or UO_305 (O_305,N_19945,N_19941);
or UO_306 (O_306,N_19816,N_19859);
or UO_307 (O_307,N_19961,N_19869);
nand UO_308 (O_308,N_19926,N_19805);
nand UO_309 (O_309,N_19917,N_19830);
nand UO_310 (O_310,N_19974,N_19816);
nand UO_311 (O_311,N_19971,N_19824);
or UO_312 (O_312,N_19994,N_19867);
or UO_313 (O_313,N_19965,N_19841);
nand UO_314 (O_314,N_19929,N_19931);
nand UO_315 (O_315,N_19995,N_19947);
and UO_316 (O_316,N_19900,N_19948);
xor UO_317 (O_317,N_19820,N_19888);
or UO_318 (O_318,N_19999,N_19913);
and UO_319 (O_319,N_19931,N_19814);
nor UO_320 (O_320,N_19893,N_19945);
nor UO_321 (O_321,N_19826,N_19916);
and UO_322 (O_322,N_19979,N_19818);
and UO_323 (O_323,N_19987,N_19997);
nand UO_324 (O_324,N_19834,N_19838);
nand UO_325 (O_325,N_19935,N_19843);
or UO_326 (O_326,N_19915,N_19997);
nand UO_327 (O_327,N_19896,N_19837);
xor UO_328 (O_328,N_19968,N_19872);
xnor UO_329 (O_329,N_19952,N_19917);
or UO_330 (O_330,N_19859,N_19815);
or UO_331 (O_331,N_19855,N_19825);
nand UO_332 (O_332,N_19911,N_19951);
nand UO_333 (O_333,N_19940,N_19915);
nor UO_334 (O_334,N_19871,N_19845);
nor UO_335 (O_335,N_19934,N_19826);
or UO_336 (O_336,N_19941,N_19963);
or UO_337 (O_337,N_19924,N_19821);
or UO_338 (O_338,N_19998,N_19849);
nand UO_339 (O_339,N_19858,N_19946);
xor UO_340 (O_340,N_19984,N_19931);
nor UO_341 (O_341,N_19990,N_19878);
or UO_342 (O_342,N_19821,N_19964);
nor UO_343 (O_343,N_19997,N_19948);
nand UO_344 (O_344,N_19968,N_19908);
and UO_345 (O_345,N_19848,N_19986);
xor UO_346 (O_346,N_19822,N_19900);
xnor UO_347 (O_347,N_19841,N_19847);
or UO_348 (O_348,N_19987,N_19880);
or UO_349 (O_349,N_19835,N_19828);
nand UO_350 (O_350,N_19957,N_19933);
nand UO_351 (O_351,N_19812,N_19843);
nor UO_352 (O_352,N_19951,N_19846);
or UO_353 (O_353,N_19871,N_19912);
nand UO_354 (O_354,N_19958,N_19962);
nand UO_355 (O_355,N_19880,N_19807);
and UO_356 (O_356,N_19925,N_19851);
nor UO_357 (O_357,N_19967,N_19969);
or UO_358 (O_358,N_19930,N_19921);
xnor UO_359 (O_359,N_19890,N_19825);
and UO_360 (O_360,N_19834,N_19971);
nor UO_361 (O_361,N_19806,N_19861);
xor UO_362 (O_362,N_19933,N_19986);
nand UO_363 (O_363,N_19982,N_19918);
nor UO_364 (O_364,N_19867,N_19879);
or UO_365 (O_365,N_19805,N_19831);
nor UO_366 (O_366,N_19988,N_19952);
nor UO_367 (O_367,N_19840,N_19941);
and UO_368 (O_368,N_19847,N_19987);
and UO_369 (O_369,N_19947,N_19894);
xor UO_370 (O_370,N_19841,N_19996);
or UO_371 (O_371,N_19972,N_19955);
nor UO_372 (O_372,N_19967,N_19941);
xor UO_373 (O_373,N_19829,N_19885);
nand UO_374 (O_374,N_19994,N_19827);
nand UO_375 (O_375,N_19972,N_19931);
or UO_376 (O_376,N_19977,N_19851);
xnor UO_377 (O_377,N_19917,N_19839);
nand UO_378 (O_378,N_19942,N_19914);
xor UO_379 (O_379,N_19820,N_19936);
or UO_380 (O_380,N_19823,N_19845);
xnor UO_381 (O_381,N_19947,N_19927);
nand UO_382 (O_382,N_19869,N_19894);
xnor UO_383 (O_383,N_19948,N_19924);
xor UO_384 (O_384,N_19803,N_19872);
nor UO_385 (O_385,N_19865,N_19883);
and UO_386 (O_386,N_19843,N_19940);
and UO_387 (O_387,N_19900,N_19979);
nor UO_388 (O_388,N_19837,N_19912);
and UO_389 (O_389,N_19881,N_19997);
nor UO_390 (O_390,N_19924,N_19830);
xnor UO_391 (O_391,N_19995,N_19815);
xnor UO_392 (O_392,N_19963,N_19822);
xor UO_393 (O_393,N_19830,N_19900);
nor UO_394 (O_394,N_19868,N_19940);
or UO_395 (O_395,N_19846,N_19890);
nor UO_396 (O_396,N_19885,N_19881);
nand UO_397 (O_397,N_19839,N_19984);
or UO_398 (O_398,N_19999,N_19985);
and UO_399 (O_399,N_19938,N_19980);
or UO_400 (O_400,N_19998,N_19996);
nand UO_401 (O_401,N_19840,N_19825);
or UO_402 (O_402,N_19913,N_19964);
or UO_403 (O_403,N_19995,N_19891);
or UO_404 (O_404,N_19939,N_19801);
nor UO_405 (O_405,N_19972,N_19962);
or UO_406 (O_406,N_19892,N_19878);
nand UO_407 (O_407,N_19859,N_19956);
and UO_408 (O_408,N_19893,N_19881);
nand UO_409 (O_409,N_19800,N_19844);
xnor UO_410 (O_410,N_19855,N_19868);
nand UO_411 (O_411,N_19910,N_19840);
and UO_412 (O_412,N_19872,N_19951);
xnor UO_413 (O_413,N_19827,N_19972);
and UO_414 (O_414,N_19841,N_19969);
nor UO_415 (O_415,N_19959,N_19925);
nand UO_416 (O_416,N_19855,N_19880);
nand UO_417 (O_417,N_19823,N_19861);
xnor UO_418 (O_418,N_19940,N_19809);
and UO_419 (O_419,N_19988,N_19870);
and UO_420 (O_420,N_19924,N_19841);
or UO_421 (O_421,N_19844,N_19847);
and UO_422 (O_422,N_19846,N_19969);
nand UO_423 (O_423,N_19980,N_19920);
xor UO_424 (O_424,N_19901,N_19827);
xor UO_425 (O_425,N_19878,N_19921);
or UO_426 (O_426,N_19852,N_19866);
or UO_427 (O_427,N_19863,N_19875);
nor UO_428 (O_428,N_19952,N_19821);
nor UO_429 (O_429,N_19918,N_19978);
xor UO_430 (O_430,N_19961,N_19897);
nand UO_431 (O_431,N_19867,N_19999);
nand UO_432 (O_432,N_19934,N_19968);
or UO_433 (O_433,N_19818,N_19896);
nor UO_434 (O_434,N_19832,N_19862);
xnor UO_435 (O_435,N_19898,N_19965);
nor UO_436 (O_436,N_19925,N_19830);
and UO_437 (O_437,N_19903,N_19993);
xor UO_438 (O_438,N_19853,N_19826);
xor UO_439 (O_439,N_19971,N_19805);
nor UO_440 (O_440,N_19966,N_19847);
and UO_441 (O_441,N_19834,N_19918);
nand UO_442 (O_442,N_19936,N_19953);
xnor UO_443 (O_443,N_19821,N_19917);
nand UO_444 (O_444,N_19976,N_19969);
or UO_445 (O_445,N_19901,N_19966);
xnor UO_446 (O_446,N_19862,N_19916);
or UO_447 (O_447,N_19984,N_19966);
or UO_448 (O_448,N_19938,N_19813);
or UO_449 (O_449,N_19896,N_19931);
or UO_450 (O_450,N_19838,N_19928);
and UO_451 (O_451,N_19991,N_19884);
and UO_452 (O_452,N_19885,N_19902);
xnor UO_453 (O_453,N_19863,N_19920);
nor UO_454 (O_454,N_19893,N_19980);
nand UO_455 (O_455,N_19878,N_19870);
and UO_456 (O_456,N_19818,N_19875);
nand UO_457 (O_457,N_19996,N_19967);
xor UO_458 (O_458,N_19961,N_19884);
nand UO_459 (O_459,N_19878,N_19868);
and UO_460 (O_460,N_19919,N_19846);
nor UO_461 (O_461,N_19804,N_19928);
xor UO_462 (O_462,N_19830,N_19971);
nor UO_463 (O_463,N_19822,N_19919);
nand UO_464 (O_464,N_19927,N_19945);
xnor UO_465 (O_465,N_19901,N_19840);
nor UO_466 (O_466,N_19800,N_19917);
nor UO_467 (O_467,N_19857,N_19896);
nand UO_468 (O_468,N_19899,N_19857);
nor UO_469 (O_469,N_19834,N_19901);
and UO_470 (O_470,N_19963,N_19918);
nor UO_471 (O_471,N_19885,N_19997);
and UO_472 (O_472,N_19972,N_19914);
xnor UO_473 (O_473,N_19824,N_19981);
nor UO_474 (O_474,N_19836,N_19839);
nand UO_475 (O_475,N_19930,N_19927);
or UO_476 (O_476,N_19810,N_19846);
xnor UO_477 (O_477,N_19922,N_19889);
xnor UO_478 (O_478,N_19867,N_19817);
xor UO_479 (O_479,N_19892,N_19862);
nand UO_480 (O_480,N_19875,N_19894);
or UO_481 (O_481,N_19899,N_19973);
nand UO_482 (O_482,N_19844,N_19907);
nand UO_483 (O_483,N_19823,N_19962);
nand UO_484 (O_484,N_19883,N_19946);
and UO_485 (O_485,N_19804,N_19910);
nand UO_486 (O_486,N_19894,N_19961);
nor UO_487 (O_487,N_19998,N_19980);
and UO_488 (O_488,N_19821,N_19864);
nand UO_489 (O_489,N_19927,N_19909);
or UO_490 (O_490,N_19804,N_19947);
and UO_491 (O_491,N_19892,N_19944);
and UO_492 (O_492,N_19924,N_19976);
or UO_493 (O_493,N_19886,N_19801);
nand UO_494 (O_494,N_19851,N_19821);
or UO_495 (O_495,N_19976,N_19876);
and UO_496 (O_496,N_19900,N_19976);
nor UO_497 (O_497,N_19993,N_19801);
nand UO_498 (O_498,N_19868,N_19958);
xor UO_499 (O_499,N_19969,N_19928);
or UO_500 (O_500,N_19858,N_19974);
and UO_501 (O_501,N_19853,N_19979);
and UO_502 (O_502,N_19872,N_19853);
nand UO_503 (O_503,N_19845,N_19895);
and UO_504 (O_504,N_19873,N_19882);
nand UO_505 (O_505,N_19858,N_19838);
nor UO_506 (O_506,N_19932,N_19904);
nand UO_507 (O_507,N_19831,N_19813);
nor UO_508 (O_508,N_19813,N_19944);
or UO_509 (O_509,N_19820,N_19860);
nor UO_510 (O_510,N_19861,N_19810);
nand UO_511 (O_511,N_19846,N_19917);
or UO_512 (O_512,N_19899,N_19887);
or UO_513 (O_513,N_19887,N_19957);
nand UO_514 (O_514,N_19806,N_19877);
nor UO_515 (O_515,N_19918,N_19969);
nand UO_516 (O_516,N_19967,N_19805);
nor UO_517 (O_517,N_19928,N_19817);
xor UO_518 (O_518,N_19910,N_19930);
nor UO_519 (O_519,N_19810,N_19936);
or UO_520 (O_520,N_19831,N_19855);
and UO_521 (O_521,N_19961,N_19814);
nand UO_522 (O_522,N_19894,N_19816);
and UO_523 (O_523,N_19867,N_19970);
nor UO_524 (O_524,N_19834,N_19848);
or UO_525 (O_525,N_19879,N_19905);
and UO_526 (O_526,N_19847,N_19843);
nand UO_527 (O_527,N_19872,N_19896);
xor UO_528 (O_528,N_19839,N_19864);
or UO_529 (O_529,N_19844,N_19976);
nor UO_530 (O_530,N_19969,N_19822);
nor UO_531 (O_531,N_19821,N_19802);
xnor UO_532 (O_532,N_19872,N_19813);
nor UO_533 (O_533,N_19926,N_19973);
or UO_534 (O_534,N_19956,N_19841);
nand UO_535 (O_535,N_19940,N_19953);
and UO_536 (O_536,N_19940,N_19966);
nor UO_537 (O_537,N_19952,N_19950);
xor UO_538 (O_538,N_19919,N_19901);
or UO_539 (O_539,N_19843,N_19811);
nor UO_540 (O_540,N_19973,N_19909);
and UO_541 (O_541,N_19819,N_19838);
and UO_542 (O_542,N_19836,N_19933);
nor UO_543 (O_543,N_19935,N_19898);
and UO_544 (O_544,N_19948,N_19830);
xnor UO_545 (O_545,N_19806,N_19901);
or UO_546 (O_546,N_19947,N_19985);
and UO_547 (O_547,N_19819,N_19812);
xnor UO_548 (O_548,N_19807,N_19926);
or UO_549 (O_549,N_19984,N_19812);
nor UO_550 (O_550,N_19885,N_19809);
or UO_551 (O_551,N_19946,N_19934);
nand UO_552 (O_552,N_19900,N_19810);
nor UO_553 (O_553,N_19809,N_19847);
xnor UO_554 (O_554,N_19882,N_19807);
nor UO_555 (O_555,N_19857,N_19945);
and UO_556 (O_556,N_19814,N_19965);
xor UO_557 (O_557,N_19947,N_19961);
nor UO_558 (O_558,N_19808,N_19852);
nor UO_559 (O_559,N_19805,N_19892);
xnor UO_560 (O_560,N_19925,N_19954);
nor UO_561 (O_561,N_19983,N_19820);
nor UO_562 (O_562,N_19847,N_19926);
nand UO_563 (O_563,N_19820,N_19830);
nor UO_564 (O_564,N_19825,N_19858);
nor UO_565 (O_565,N_19922,N_19986);
xnor UO_566 (O_566,N_19907,N_19873);
nand UO_567 (O_567,N_19856,N_19917);
xnor UO_568 (O_568,N_19836,N_19896);
nand UO_569 (O_569,N_19934,N_19984);
or UO_570 (O_570,N_19873,N_19957);
nand UO_571 (O_571,N_19921,N_19811);
and UO_572 (O_572,N_19957,N_19813);
or UO_573 (O_573,N_19943,N_19983);
nor UO_574 (O_574,N_19984,N_19861);
or UO_575 (O_575,N_19984,N_19885);
xor UO_576 (O_576,N_19829,N_19860);
nor UO_577 (O_577,N_19927,N_19899);
and UO_578 (O_578,N_19983,N_19914);
or UO_579 (O_579,N_19943,N_19872);
nand UO_580 (O_580,N_19990,N_19967);
nor UO_581 (O_581,N_19898,N_19842);
and UO_582 (O_582,N_19924,N_19909);
nor UO_583 (O_583,N_19909,N_19989);
and UO_584 (O_584,N_19918,N_19904);
nand UO_585 (O_585,N_19925,N_19961);
nand UO_586 (O_586,N_19801,N_19973);
xor UO_587 (O_587,N_19823,N_19996);
and UO_588 (O_588,N_19953,N_19932);
nor UO_589 (O_589,N_19809,N_19819);
nand UO_590 (O_590,N_19970,N_19820);
xor UO_591 (O_591,N_19922,N_19886);
nor UO_592 (O_592,N_19812,N_19886);
xor UO_593 (O_593,N_19818,N_19914);
and UO_594 (O_594,N_19936,N_19861);
and UO_595 (O_595,N_19869,N_19871);
and UO_596 (O_596,N_19929,N_19904);
or UO_597 (O_597,N_19897,N_19855);
nor UO_598 (O_598,N_19868,N_19870);
nand UO_599 (O_599,N_19865,N_19978);
and UO_600 (O_600,N_19988,N_19900);
or UO_601 (O_601,N_19861,N_19847);
nand UO_602 (O_602,N_19818,N_19945);
xnor UO_603 (O_603,N_19937,N_19996);
nor UO_604 (O_604,N_19970,N_19859);
or UO_605 (O_605,N_19872,N_19994);
xor UO_606 (O_606,N_19877,N_19970);
nor UO_607 (O_607,N_19967,N_19868);
xor UO_608 (O_608,N_19885,N_19966);
or UO_609 (O_609,N_19909,N_19979);
xnor UO_610 (O_610,N_19876,N_19871);
xnor UO_611 (O_611,N_19990,N_19883);
and UO_612 (O_612,N_19821,N_19980);
nor UO_613 (O_613,N_19862,N_19950);
and UO_614 (O_614,N_19856,N_19893);
xnor UO_615 (O_615,N_19975,N_19853);
and UO_616 (O_616,N_19862,N_19881);
or UO_617 (O_617,N_19969,N_19973);
xnor UO_618 (O_618,N_19931,N_19912);
nand UO_619 (O_619,N_19855,N_19973);
and UO_620 (O_620,N_19957,N_19892);
nand UO_621 (O_621,N_19911,N_19919);
and UO_622 (O_622,N_19857,N_19833);
nor UO_623 (O_623,N_19941,N_19949);
xor UO_624 (O_624,N_19981,N_19920);
and UO_625 (O_625,N_19916,N_19912);
or UO_626 (O_626,N_19841,N_19852);
nand UO_627 (O_627,N_19874,N_19910);
nor UO_628 (O_628,N_19978,N_19870);
and UO_629 (O_629,N_19977,N_19840);
and UO_630 (O_630,N_19900,N_19963);
xnor UO_631 (O_631,N_19947,N_19946);
nor UO_632 (O_632,N_19838,N_19803);
nor UO_633 (O_633,N_19862,N_19993);
and UO_634 (O_634,N_19922,N_19984);
nand UO_635 (O_635,N_19851,N_19948);
or UO_636 (O_636,N_19979,N_19825);
nor UO_637 (O_637,N_19920,N_19881);
or UO_638 (O_638,N_19976,N_19885);
nor UO_639 (O_639,N_19936,N_19837);
nand UO_640 (O_640,N_19955,N_19802);
and UO_641 (O_641,N_19843,N_19948);
xnor UO_642 (O_642,N_19980,N_19943);
nand UO_643 (O_643,N_19962,N_19851);
or UO_644 (O_644,N_19808,N_19965);
xor UO_645 (O_645,N_19800,N_19854);
and UO_646 (O_646,N_19969,N_19931);
or UO_647 (O_647,N_19854,N_19923);
nor UO_648 (O_648,N_19842,N_19899);
or UO_649 (O_649,N_19918,N_19878);
xnor UO_650 (O_650,N_19954,N_19923);
and UO_651 (O_651,N_19901,N_19848);
nor UO_652 (O_652,N_19932,N_19814);
or UO_653 (O_653,N_19913,N_19879);
or UO_654 (O_654,N_19965,N_19954);
or UO_655 (O_655,N_19998,N_19876);
nand UO_656 (O_656,N_19804,N_19957);
and UO_657 (O_657,N_19973,N_19895);
nand UO_658 (O_658,N_19974,N_19943);
nor UO_659 (O_659,N_19906,N_19948);
or UO_660 (O_660,N_19876,N_19856);
and UO_661 (O_661,N_19910,N_19894);
and UO_662 (O_662,N_19928,N_19900);
nand UO_663 (O_663,N_19873,N_19834);
xor UO_664 (O_664,N_19908,N_19991);
nor UO_665 (O_665,N_19935,N_19937);
nor UO_666 (O_666,N_19939,N_19852);
xor UO_667 (O_667,N_19937,N_19946);
xnor UO_668 (O_668,N_19848,N_19977);
nor UO_669 (O_669,N_19979,N_19997);
and UO_670 (O_670,N_19926,N_19841);
xnor UO_671 (O_671,N_19944,N_19876);
or UO_672 (O_672,N_19928,N_19864);
or UO_673 (O_673,N_19891,N_19850);
nand UO_674 (O_674,N_19930,N_19957);
nor UO_675 (O_675,N_19997,N_19856);
nand UO_676 (O_676,N_19941,N_19932);
nand UO_677 (O_677,N_19957,N_19899);
nand UO_678 (O_678,N_19863,N_19870);
or UO_679 (O_679,N_19942,N_19939);
nor UO_680 (O_680,N_19844,N_19824);
nand UO_681 (O_681,N_19989,N_19842);
nor UO_682 (O_682,N_19800,N_19919);
and UO_683 (O_683,N_19858,N_19951);
nand UO_684 (O_684,N_19987,N_19829);
or UO_685 (O_685,N_19978,N_19821);
or UO_686 (O_686,N_19906,N_19838);
xor UO_687 (O_687,N_19989,N_19844);
xnor UO_688 (O_688,N_19941,N_19924);
xor UO_689 (O_689,N_19903,N_19918);
nor UO_690 (O_690,N_19983,N_19897);
nor UO_691 (O_691,N_19880,N_19849);
or UO_692 (O_692,N_19999,N_19938);
nand UO_693 (O_693,N_19824,N_19886);
or UO_694 (O_694,N_19998,N_19912);
xnor UO_695 (O_695,N_19858,N_19812);
xor UO_696 (O_696,N_19826,N_19856);
or UO_697 (O_697,N_19810,N_19914);
nand UO_698 (O_698,N_19803,N_19967);
nand UO_699 (O_699,N_19922,N_19882);
nor UO_700 (O_700,N_19956,N_19927);
nor UO_701 (O_701,N_19941,N_19826);
nor UO_702 (O_702,N_19934,N_19915);
and UO_703 (O_703,N_19871,N_19842);
or UO_704 (O_704,N_19912,N_19862);
nand UO_705 (O_705,N_19832,N_19831);
or UO_706 (O_706,N_19948,N_19942);
nor UO_707 (O_707,N_19851,N_19958);
or UO_708 (O_708,N_19855,N_19893);
and UO_709 (O_709,N_19899,N_19981);
nand UO_710 (O_710,N_19918,N_19900);
nand UO_711 (O_711,N_19848,N_19835);
nor UO_712 (O_712,N_19929,N_19802);
xor UO_713 (O_713,N_19946,N_19817);
or UO_714 (O_714,N_19886,N_19893);
nor UO_715 (O_715,N_19910,N_19973);
xnor UO_716 (O_716,N_19901,N_19832);
nor UO_717 (O_717,N_19865,N_19860);
nor UO_718 (O_718,N_19959,N_19902);
and UO_719 (O_719,N_19875,N_19904);
xor UO_720 (O_720,N_19831,N_19850);
nand UO_721 (O_721,N_19815,N_19947);
nand UO_722 (O_722,N_19834,N_19854);
xor UO_723 (O_723,N_19908,N_19863);
nand UO_724 (O_724,N_19907,N_19806);
or UO_725 (O_725,N_19977,N_19895);
or UO_726 (O_726,N_19978,N_19898);
nand UO_727 (O_727,N_19901,N_19990);
or UO_728 (O_728,N_19965,N_19978);
nor UO_729 (O_729,N_19922,N_19899);
xor UO_730 (O_730,N_19891,N_19815);
or UO_731 (O_731,N_19842,N_19823);
nand UO_732 (O_732,N_19838,N_19988);
nor UO_733 (O_733,N_19910,N_19889);
nand UO_734 (O_734,N_19821,N_19889);
or UO_735 (O_735,N_19873,N_19923);
xnor UO_736 (O_736,N_19855,N_19997);
and UO_737 (O_737,N_19855,N_19885);
nor UO_738 (O_738,N_19820,N_19831);
nand UO_739 (O_739,N_19865,N_19995);
nand UO_740 (O_740,N_19954,N_19852);
nor UO_741 (O_741,N_19987,N_19894);
nor UO_742 (O_742,N_19801,N_19810);
and UO_743 (O_743,N_19852,N_19981);
nand UO_744 (O_744,N_19950,N_19828);
nor UO_745 (O_745,N_19964,N_19825);
and UO_746 (O_746,N_19853,N_19953);
xor UO_747 (O_747,N_19841,N_19814);
nor UO_748 (O_748,N_19957,N_19895);
xnor UO_749 (O_749,N_19976,N_19837);
and UO_750 (O_750,N_19955,N_19971);
or UO_751 (O_751,N_19886,N_19935);
nor UO_752 (O_752,N_19947,N_19855);
xnor UO_753 (O_753,N_19834,N_19942);
or UO_754 (O_754,N_19870,N_19902);
nor UO_755 (O_755,N_19812,N_19839);
xnor UO_756 (O_756,N_19988,N_19802);
nand UO_757 (O_757,N_19915,N_19928);
nand UO_758 (O_758,N_19970,N_19813);
and UO_759 (O_759,N_19954,N_19876);
or UO_760 (O_760,N_19935,N_19891);
nor UO_761 (O_761,N_19828,N_19922);
xor UO_762 (O_762,N_19936,N_19821);
and UO_763 (O_763,N_19940,N_19913);
nand UO_764 (O_764,N_19890,N_19940);
and UO_765 (O_765,N_19968,N_19978);
and UO_766 (O_766,N_19878,N_19876);
xor UO_767 (O_767,N_19939,N_19993);
or UO_768 (O_768,N_19993,N_19834);
or UO_769 (O_769,N_19805,N_19879);
or UO_770 (O_770,N_19892,N_19937);
or UO_771 (O_771,N_19835,N_19954);
nand UO_772 (O_772,N_19988,N_19897);
xnor UO_773 (O_773,N_19979,N_19879);
and UO_774 (O_774,N_19909,N_19965);
and UO_775 (O_775,N_19909,N_19803);
and UO_776 (O_776,N_19831,N_19907);
nor UO_777 (O_777,N_19868,N_19845);
nand UO_778 (O_778,N_19840,N_19899);
nor UO_779 (O_779,N_19801,N_19830);
nor UO_780 (O_780,N_19805,N_19847);
and UO_781 (O_781,N_19854,N_19868);
nor UO_782 (O_782,N_19881,N_19866);
or UO_783 (O_783,N_19806,N_19856);
and UO_784 (O_784,N_19998,N_19987);
or UO_785 (O_785,N_19906,N_19902);
nand UO_786 (O_786,N_19850,N_19906);
and UO_787 (O_787,N_19875,N_19998);
and UO_788 (O_788,N_19994,N_19819);
nor UO_789 (O_789,N_19908,N_19872);
xnor UO_790 (O_790,N_19903,N_19927);
nand UO_791 (O_791,N_19877,N_19880);
or UO_792 (O_792,N_19971,N_19991);
xnor UO_793 (O_793,N_19850,N_19967);
or UO_794 (O_794,N_19821,N_19815);
and UO_795 (O_795,N_19898,N_19876);
and UO_796 (O_796,N_19947,N_19840);
nand UO_797 (O_797,N_19834,N_19949);
and UO_798 (O_798,N_19866,N_19888);
xnor UO_799 (O_799,N_19808,N_19954);
nand UO_800 (O_800,N_19979,N_19987);
nand UO_801 (O_801,N_19852,N_19989);
xnor UO_802 (O_802,N_19927,N_19905);
or UO_803 (O_803,N_19884,N_19881);
nor UO_804 (O_804,N_19917,N_19978);
xnor UO_805 (O_805,N_19882,N_19916);
and UO_806 (O_806,N_19998,N_19850);
or UO_807 (O_807,N_19970,N_19946);
or UO_808 (O_808,N_19982,N_19892);
xor UO_809 (O_809,N_19849,N_19915);
and UO_810 (O_810,N_19962,N_19995);
nand UO_811 (O_811,N_19942,N_19851);
nor UO_812 (O_812,N_19861,N_19851);
xnor UO_813 (O_813,N_19950,N_19839);
xor UO_814 (O_814,N_19930,N_19901);
and UO_815 (O_815,N_19912,N_19936);
nand UO_816 (O_816,N_19948,N_19982);
nand UO_817 (O_817,N_19941,N_19813);
or UO_818 (O_818,N_19873,N_19897);
or UO_819 (O_819,N_19911,N_19945);
and UO_820 (O_820,N_19971,N_19884);
xnor UO_821 (O_821,N_19851,N_19829);
xor UO_822 (O_822,N_19845,N_19919);
or UO_823 (O_823,N_19949,N_19808);
and UO_824 (O_824,N_19940,N_19861);
and UO_825 (O_825,N_19971,N_19906);
and UO_826 (O_826,N_19971,N_19888);
or UO_827 (O_827,N_19853,N_19962);
nand UO_828 (O_828,N_19830,N_19979);
or UO_829 (O_829,N_19885,N_19853);
and UO_830 (O_830,N_19861,N_19944);
and UO_831 (O_831,N_19900,N_19914);
and UO_832 (O_832,N_19858,N_19926);
nor UO_833 (O_833,N_19973,N_19846);
xnor UO_834 (O_834,N_19817,N_19811);
nor UO_835 (O_835,N_19984,N_19950);
nand UO_836 (O_836,N_19883,N_19900);
or UO_837 (O_837,N_19823,N_19804);
nand UO_838 (O_838,N_19826,N_19830);
and UO_839 (O_839,N_19836,N_19901);
or UO_840 (O_840,N_19915,N_19802);
or UO_841 (O_841,N_19910,N_19865);
and UO_842 (O_842,N_19815,N_19983);
or UO_843 (O_843,N_19914,N_19986);
nand UO_844 (O_844,N_19893,N_19815);
xor UO_845 (O_845,N_19936,N_19900);
nand UO_846 (O_846,N_19826,N_19818);
nor UO_847 (O_847,N_19833,N_19854);
xor UO_848 (O_848,N_19841,N_19983);
xnor UO_849 (O_849,N_19854,N_19896);
nand UO_850 (O_850,N_19927,N_19832);
xor UO_851 (O_851,N_19897,N_19880);
and UO_852 (O_852,N_19835,N_19893);
nor UO_853 (O_853,N_19834,N_19889);
or UO_854 (O_854,N_19921,N_19820);
xor UO_855 (O_855,N_19957,N_19940);
xnor UO_856 (O_856,N_19999,N_19948);
or UO_857 (O_857,N_19811,N_19806);
xor UO_858 (O_858,N_19810,N_19831);
xor UO_859 (O_859,N_19972,N_19809);
and UO_860 (O_860,N_19854,N_19912);
or UO_861 (O_861,N_19908,N_19969);
xnor UO_862 (O_862,N_19883,N_19880);
and UO_863 (O_863,N_19845,N_19975);
and UO_864 (O_864,N_19972,N_19985);
nand UO_865 (O_865,N_19841,N_19931);
xor UO_866 (O_866,N_19868,N_19823);
or UO_867 (O_867,N_19821,N_19855);
nand UO_868 (O_868,N_19909,N_19868);
xor UO_869 (O_869,N_19911,N_19967);
and UO_870 (O_870,N_19804,N_19981);
and UO_871 (O_871,N_19875,N_19993);
and UO_872 (O_872,N_19938,N_19852);
xor UO_873 (O_873,N_19801,N_19808);
and UO_874 (O_874,N_19979,N_19842);
nand UO_875 (O_875,N_19844,N_19906);
xor UO_876 (O_876,N_19910,N_19937);
nand UO_877 (O_877,N_19968,N_19806);
nor UO_878 (O_878,N_19899,N_19992);
nand UO_879 (O_879,N_19837,N_19932);
and UO_880 (O_880,N_19839,N_19828);
and UO_881 (O_881,N_19887,N_19878);
nand UO_882 (O_882,N_19884,N_19806);
nand UO_883 (O_883,N_19966,N_19879);
and UO_884 (O_884,N_19989,N_19913);
and UO_885 (O_885,N_19909,N_19944);
and UO_886 (O_886,N_19955,N_19828);
nor UO_887 (O_887,N_19882,N_19826);
nand UO_888 (O_888,N_19873,N_19910);
or UO_889 (O_889,N_19915,N_19816);
or UO_890 (O_890,N_19802,N_19854);
nand UO_891 (O_891,N_19975,N_19876);
nor UO_892 (O_892,N_19992,N_19806);
and UO_893 (O_893,N_19818,N_19824);
nand UO_894 (O_894,N_19893,N_19986);
or UO_895 (O_895,N_19986,N_19960);
nand UO_896 (O_896,N_19838,N_19855);
nand UO_897 (O_897,N_19811,N_19927);
or UO_898 (O_898,N_19910,N_19866);
nor UO_899 (O_899,N_19953,N_19928);
nor UO_900 (O_900,N_19933,N_19819);
or UO_901 (O_901,N_19908,N_19948);
nor UO_902 (O_902,N_19880,N_19868);
xor UO_903 (O_903,N_19912,N_19833);
and UO_904 (O_904,N_19995,N_19979);
xor UO_905 (O_905,N_19888,N_19902);
xnor UO_906 (O_906,N_19894,N_19859);
or UO_907 (O_907,N_19936,N_19978);
or UO_908 (O_908,N_19873,N_19880);
and UO_909 (O_909,N_19814,N_19881);
nor UO_910 (O_910,N_19903,N_19883);
xnor UO_911 (O_911,N_19882,N_19942);
or UO_912 (O_912,N_19908,N_19972);
xnor UO_913 (O_913,N_19836,N_19888);
nor UO_914 (O_914,N_19822,N_19994);
or UO_915 (O_915,N_19874,N_19892);
or UO_916 (O_916,N_19935,N_19975);
and UO_917 (O_917,N_19933,N_19938);
xor UO_918 (O_918,N_19860,N_19868);
nor UO_919 (O_919,N_19944,N_19908);
and UO_920 (O_920,N_19849,N_19960);
nor UO_921 (O_921,N_19888,N_19846);
nand UO_922 (O_922,N_19927,N_19966);
or UO_923 (O_923,N_19904,N_19970);
nor UO_924 (O_924,N_19807,N_19900);
and UO_925 (O_925,N_19805,N_19974);
nor UO_926 (O_926,N_19885,N_19821);
nor UO_927 (O_927,N_19802,N_19841);
nand UO_928 (O_928,N_19988,N_19956);
xnor UO_929 (O_929,N_19836,N_19899);
nand UO_930 (O_930,N_19903,N_19991);
nor UO_931 (O_931,N_19949,N_19980);
xnor UO_932 (O_932,N_19981,N_19811);
or UO_933 (O_933,N_19941,N_19903);
and UO_934 (O_934,N_19955,N_19858);
nand UO_935 (O_935,N_19804,N_19881);
nor UO_936 (O_936,N_19854,N_19918);
nand UO_937 (O_937,N_19819,N_19801);
and UO_938 (O_938,N_19872,N_19875);
and UO_939 (O_939,N_19801,N_19875);
nor UO_940 (O_940,N_19881,N_19825);
xnor UO_941 (O_941,N_19884,N_19879);
and UO_942 (O_942,N_19949,N_19860);
or UO_943 (O_943,N_19842,N_19850);
xnor UO_944 (O_944,N_19881,N_19829);
and UO_945 (O_945,N_19850,N_19974);
and UO_946 (O_946,N_19897,N_19810);
or UO_947 (O_947,N_19924,N_19842);
nor UO_948 (O_948,N_19817,N_19824);
or UO_949 (O_949,N_19924,N_19940);
or UO_950 (O_950,N_19999,N_19813);
nor UO_951 (O_951,N_19947,N_19983);
nand UO_952 (O_952,N_19874,N_19850);
xnor UO_953 (O_953,N_19995,N_19824);
or UO_954 (O_954,N_19940,N_19901);
nand UO_955 (O_955,N_19963,N_19826);
nand UO_956 (O_956,N_19968,N_19989);
xor UO_957 (O_957,N_19953,N_19868);
and UO_958 (O_958,N_19917,N_19900);
and UO_959 (O_959,N_19950,N_19803);
xnor UO_960 (O_960,N_19964,N_19936);
or UO_961 (O_961,N_19906,N_19830);
or UO_962 (O_962,N_19800,N_19843);
and UO_963 (O_963,N_19817,N_19802);
or UO_964 (O_964,N_19804,N_19997);
xor UO_965 (O_965,N_19803,N_19884);
nor UO_966 (O_966,N_19996,N_19835);
nand UO_967 (O_967,N_19922,N_19968);
xor UO_968 (O_968,N_19837,N_19935);
nand UO_969 (O_969,N_19886,N_19909);
xor UO_970 (O_970,N_19974,N_19915);
and UO_971 (O_971,N_19946,N_19910);
nand UO_972 (O_972,N_19974,N_19924);
nor UO_973 (O_973,N_19903,N_19922);
xnor UO_974 (O_974,N_19809,N_19914);
xnor UO_975 (O_975,N_19982,N_19914);
xnor UO_976 (O_976,N_19922,N_19896);
nand UO_977 (O_977,N_19923,N_19853);
nand UO_978 (O_978,N_19847,N_19925);
nand UO_979 (O_979,N_19933,N_19990);
or UO_980 (O_980,N_19950,N_19928);
nor UO_981 (O_981,N_19871,N_19821);
xor UO_982 (O_982,N_19901,N_19855);
nor UO_983 (O_983,N_19862,N_19915);
and UO_984 (O_984,N_19972,N_19801);
or UO_985 (O_985,N_19827,N_19830);
nor UO_986 (O_986,N_19966,N_19924);
and UO_987 (O_987,N_19800,N_19858);
nand UO_988 (O_988,N_19983,N_19939);
xnor UO_989 (O_989,N_19874,N_19997);
and UO_990 (O_990,N_19975,N_19949);
or UO_991 (O_991,N_19816,N_19983);
xnor UO_992 (O_992,N_19825,N_19917);
or UO_993 (O_993,N_19886,N_19897);
and UO_994 (O_994,N_19886,N_19855);
and UO_995 (O_995,N_19839,N_19831);
nor UO_996 (O_996,N_19908,N_19822);
or UO_997 (O_997,N_19971,N_19814);
nand UO_998 (O_998,N_19943,N_19893);
or UO_999 (O_999,N_19902,N_19857);
and UO_1000 (O_1000,N_19867,N_19822);
nor UO_1001 (O_1001,N_19802,N_19917);
and UO_1002 (O_1002,N_19933,N_19912);
xnor UO_1003 (O_1003,N_19863,N_19824);
or UO_1004 (O_1004,N_19812,N_19913);
and UO_1005 (O_1005,N_19886,N_19984);
or UO_1006 (O_1006,N_19970,N_19834);
or UO_1007 (O_1007,N_19874,N_19856);
xor UO_1008 (O_1008,N_19811,N_19920);
and UO_1009 (O_1009,N_19852,N_19859);
xor UO_1010 (O_1010,N_19897,N_19805);
nand UO_1011 (O_1011,N_19887,N_19848);
and UO_1012 (O_1012,N_19919,N_19958);
nand UO_1013 (O_1013,N_19914,N_19923);
or UO_1014 (O_1014,N_19953,N_19943);
and UO_1015 (O_1015,N_19984,N_19823);
nand UO_1016 (O_1016,N_19960,N_19896);
or UO_1017 (O_1017,N_19907,N_19918);
nor UO_1018 (O_1018,N_19939,N_19941);
xnor UO_1019 (O_1019,N_19842,N_19995);
and UO_1020 (O_1020,N_19880,N_19963);
xor UO_1021 (O_1021,N_19961,N_19870);
and UO_1022 (O_1022,N_19809,N_19932);
nor UO_1023 (O_1023,N_19808,N_19882);
xor UO_1024 (O_1024,N_19987,N_19904);
nor UO_1025 (O_1025,N_19845,N_19915);
or UO_1026 (O_1026,N_19878,N_19938);
nand UO_1027 (O_1027,N_19822,N_19814);
nand UO_1028 (O_1028,N_19848,N_19818);
or UO_1029 (O_1029,N_19884,N_19932);
or UO_1030 (O_1030,N_19887,N_19959);
and UO_1031 (O_1031,N_19829,N_19804);
xor UO_1032 (O_1032,N_19986,N_19972);
xor UO_1033 (O_1033,N_19945,N_19948);
nor UO_1034 (O_1034,N_19972,N_19831);
and UO_1035 (O_1035,N_19828,N_19936);
xor UO_1036 (O_1036,N_19851,N_19806);
and UO_1037 (O_1037,N_19987,N_19913);
nand UO_1038 (O_1038,N_19818,N_19820);
nand UO_1039 (O_1039,N_19909,N_19985);
and UO_1040 (O_1040,N_19949,N_19895);
nand UO_1041 (O_1041,N_19942,N_19806);
or UO_1042 (O_1042,N_19972,N_19807);
nor UO_1043 (O_1043,N_19932,N_19852);
xnor UO_1044 (O_1044,N_19908,N_19983);
nand UO_1045 (O_1045,N_19840,N_19971);
nor UO_1046 (O_1046,N_19991,N_19842);
nor UO_1047 (O_1047,N_19808,N_19883);
nor UO_1048 (O_1048,N_19971,N_19986);
xnor UO_1049 (O_1049,N_19987,N_19967);
nand UO_1050 (O_1050,N_19950,N_19992);
nor UO_1051 (O_1051,N_19849,N_19974);
nor UO_1052 (O_1052,N_19913,N_19898);
nand UO_1053 (O_1053,N_19919,N_19984);
and UO_1054 (O_1054,N_19968,N_19823);
and UO_1055 (O_1055,N_19836,N_19991);
nor UO_1056 (O_1056,N_19928,N_19934);
nand UO_1057 (O_1057,N_19869,N_19892);
xor UO_1058 (O_1058,N_19880,N_19954);
nor UO_1059 (O_1059,N_19970,N_19804);
and UO_1060 (O_1060,N_19986,N_19835);
or UO_1061 (O_1061,N_19823,N_19884);
nand UO_1062 (O_1062,N_19917,N_19968);
nand UO_1063 (O_1063,N_19870,N_19856);
xor UO_1064 (O_1064,N_19967,N_19977);
nand UO_1065 (O_1065,N_19822,N_19899);
nand UO_1066 (O_1066,N_19819,N_19916);
or UO_1067 (O_1067,N_19887,N_19974);
xnor UO_1068 (O_1068,N_19951,N_19956);
or UO_1069 (O_1069,N_19921,N_19860);
nand UO_1070 (O_1070,N_19925,N_19836);
or UO_1071 (O_1071,N_19851,N_19950);
nor UO_1072 (O_1072,N_19867,N_19862);
or UO_1073 (O_1073,N_19814,N_19940);
nand UO_1074 (O_1074,N_19931,N_19894);
xor UO_1075 (O_1075,N_19819,N_19833);
or UO_1076 (O_1076,N_19847,N_19934);
or UO_1077 (O_1077,N_19924,N_19954);
nand UO_1078 (O_1078,N_19975,N_19800);
nand UO_1079 (O_1079,N_19971,N_19836);
or UO_1080 (O_1080,N_19879,N_19972);
nor UO_1081 (O_1081,N_19984,N_19876);
xor UO_1082 (O_1082,N_19929,N_19825);
and UO_1083 (O_1083,N_19936,N_19939);
nor UO_1084 (O_1084,N_19812,N_19894);
nand UO_1085 (O_1085,N_19981,N_19950);
nor UO_1086 (O_1086,N_19940,N_19993);
nand UO_1087 (O_1087,N_19871,N_19924);
or UO_1088 (O_1088,N_19939,N_19961);
nor UO_1089 (O_1089,N_19891,N_19837);
or UO_1090 (O_1090,N_19979,N_19950);
and UO_1091 (O_1091,N_19867,N_19821);
and UO_1092 (O_1092,N_19804,N_19921);
nor UO_1093 (O_1093,N_19990,N_19806);
nor UO_1094 (O_1094,N_19853,N_19916);
and UO_1095 (O_1095,N_19936,N_19902);
and UO_1096 (O_1096,N_19839,N_19993);
or UO_1097 (O_1097,N_19899,N_19963);
or UO_1098 (O_1098,N_19824,N_19832);
nand UO_1099 (O_1099,N_19984,N_19895);
xnor UO_1100 (O_1100,N_19802,N_19813);
xor UO_1101 (O_1101,N_19838,N_19823);
or UO_1102 (O_1102,N_19897,N_19800);
nand UO_1103 (O_1103,N_19997,N_19817);
nor UO_1104 (O_1104,N_19911,N_19859);
or UO_1105 (O_1105,N_19964,N_19830);
nand UO_1106 (O_1106,N_19874,N_19887);
xor UO_1107 (O_1107,N_19838,N_19876);
xnor UO_1108 (O_1108,N_19935,N_19841);
or UO_1109 (O_1109,N_19994,N_19946);
nand UO_1110 (O_1110,N_19897,N_19831);
nand UO_1111 (O_1111,N_19986,N_19819);
and UO_1112 (O_1112,N_19857,N_19843);
xnor UO_1113 (O_1113,N_19886,N_19890);
xor UO_1114 (O_1114,N_19816,N_19807);
or UO_1115 (O_1115,N_19867,N_19947);
and UO_1116 (O_1116,N_19903,N_19881);
nor UO_1117 (O_1117,N_19885,N_19800);
or UO_1118 (O_1118,N_19910,N_19846);
nor UO_1119 (O_1119,N_19890,N_19859);
or UO_1120 (O_1120,N_19867,N_19950);
or UO_1121 (O_1121,N_19967,N_19920);
and UO_1122 (O_1122,N_19859,N_19849);
and UO_1123 (O_1123,N_19843,N_19877);
xor UO_1124 (O_1124,N_19954,N_19917);
nor UO_1125 (O_1125,N_19846,N_19837);
nor UO_1126 (O_1126,N_19988,N_19930);
nand UO_1127 (O_1127,N_19992,N_19985);
or UO_1128 (O_1128,N_19879,N_19892);
nand UO_1129 (O_1129,N_19824,N_19830);
and UO_1130 (O_1130,N_19945,N_19835);
or UO_1131 (O_1131,N_19840,N_19824);
xnor UO_1132 (O_1132,N_19906,N_19835);
xor UO_1133 (O_1133,N_19920,N_19875);
nand UO_1134 (O_1134,N_19986,N_19934);
nor UO_1135 (O_1135,N_19839,N_19880);
or UO_1136 (O_1136,N_19956,N_19964);
nor UO_1137 (O_1137,N_19948,N_19904);
nor UO_1138 (O_1138,N_19844,N_19801);
nand UO_1139 (O_1139,N_19841,N_19928);
or UO_1140 (O_1140,N_19885,N_19856);
or UO_1141 (O_1141,N_19929,N_19829);
nor UO_1142 (O_1142,N_19805,N_19959);
nor UO_1143 (O_1143,N_19903,N_19968);
and UO_1144 (O_1144,N_19942,N_19905);
nand UO_1145 (O_1145,N_19930,N_19808);
nand UO_1146 (O_1146,N_19808,N_19884);
xor UO_1147 (O_1147,N_19969,N_19896);
xnor UO_1148 (O_1148,N_19938,N_19950);
nor UO_1149 (O_1149,N_19909,N_19942);
nand UO_1150 (O_1150,N_19852,N_19847);
xnor UO_1151 (O_1151,N_19930,N_19809);
and UO_1152 (O_1152,N_19804,N_19922);
nand UO_1153 (O_1153,N_19977,N_19886);
and UO_1154 (O_1154,N_19899,N_19854);
nor UO_1155 (O_1155,N_19917,N_19838);
nor UO_1156 (O_1156,N_19901,N_19893);
nand UO_1157 (O_1157,N_19930,N_19883);
nor UO_1158 (O_1158,N_19923,N_19868);
or UO_1159 (O_1159,N_19999,N_19954);
and UO_1160 (O_1160,N_19907,N_19864);
nand UO_1161 (O_1161,N_19920,N_19951);
nand UO_1162 (O_1162,N_19983,N_19812);
and UO_1163 (O_1163,N_19848,N_19968);
nand UO_1164 (O_1164,N_19914,N_19932);
and UO_1165 (O_1165,N_19868,N_19806);
or UO_1166 (O_1166,N_19917,N_19885);
and UO_1167 (O_1167,N_19895,N_19976);
nand UO_1168 (O_1168,N_19957,N_19847);
xnor UO_1169 (O_1169,N_19996,N_19880);
nor UO_1170 (O_1170,N_19985,N_19878);
nor UO_1171 (O_1171,N_19987,N_19832);
and UO_1172 (O_1172,N_19893,N_19819);
nand UO_1173 (O_1173,N_19851,N_19921);
nor UO_1174 (O_1174,N_19958,N_19882);
or UO_1175 (O_1175,N_19950,N_19960);
nand UO_1176 (O_1176,N_19966,N_19986);
or UO_1177 (O_1177,N_19954,N_19803);
nor UO_1178 (O_1178,N_19876,N_19993);
or UO_1179 (O_1179,N_19971,N_19870);
nor UO_1180 (O_1180,N_19996,N_19952);
nor UO_1181 (O_1181,N_19801,N_19820);
nor UO_1182 (O_1182,N_19949,N_19953);
and UO_1183 (O_1183,N_19947,N_19814);
xor UO_1184 (O_1184,N_19989,N_19949);
or UO_1185 (O_1185,N_19926,N_19825);
nand UO_1186 (O_1186,N_19894,N_19814);
nor UO_1187 (O_1187,N_19849,N_19919);
and UO_1188 (O_1188,N_19831,N_19827);
nand UO_1189 (O_1189,N_19986,N_19802);
or UO_1190 (O_1190,N_19941,N_19825);
or UO_1191 (O_1191,N_19850,N_19841);
xor UO_1192 (O_1192,N_19905,N_19902);
or UO_1193 (O_1193,N_19846,N_19871);
nand UO_1194 (O_1194,N_19962,N_19907);
and UO_1195 (O_1195,N_19815,N_19921);
and UO_1196 (O_1196,N_19844,N_19839);
nand UO_1197 (O_1197,N_19949,N_19916);
xnor UO_1198 (O_1198,N_19849,N_19818);
and UO_1199 (O_1199,N_19889,N_19946);
nor UO_1200 (O_1200,N_19819,N_19830);
nor UO_1201 (O_1201,N_19809,N_19913);
nand UO_1202 (O_1202,N_19913,N_19947);
and UO_1203 (O_1203,N_19877,N_19858);
or UO_1204 (O_1204,N_19885,N_19926);
nor UO_1205 (O_1205,N_19965,N_19974);
and UO_1206 (O_1206,N_19983,N_19924);
nor UO_1207 (O_1207,N_19942,N_19896);
xor UO_1208 (O_1208,N_19993,N_19829);
and UO_1209 (O_1209,N_19896,N_19875);
and UO_1210 (O_1210,N_19964,N_19965);
xor UO_1211 (O_1211,N_19905,N_19896);
nor UO_1212 (O_1212,N_19939,N_19915);
or UO_1213 (O_1213,N_19902,N_19941);
or UO_1214 (O_1214,N_19934,N_19897);
xnor UO_1215 (O_1215,N_19839,N_19979);
or UO_1216 (O_1216,N_19874,N_19896);
and UO_1217 (O_1217,N_19825,N_19818);
nor UO_1218 (O_1218,N_19989,N_19826);
nand UO_1219 (O_1219,N_19989,N_19827);
nand UO_1220 (O_1220,N_19886,N_19962);
xnor UO_1221 (O_1221,N_19838,N_19840);
nor UO_1222 (O_1222,N_19872,N_19833);
xor UO_1223 (O_1223,N_19822,N_19962);
nand UO_1224 (O_1224,N_19998,N_19897);
nand UO_1225 (O_1225,N_19835,N_19818);
nor UO_1226 (O_1226,N_19816,N_19847);
and UO_1227 (O_1227,N_19896,N_19832);
or UO_1228 (O_1228,N_19893,N_19948);
nand UO_1229 (O_1229,N_19879,N_19823);
or UO_1230 (O_1230,N_19954,N_19843);
and UO_1231 (O_1231,N_19945,N_19906);
nor UO_1232 (O_1232,N_19802,N_19865);
xnor UO_1233 (O_1233,N_19936,N_19835);
or UO_1234 (O_1234,N_19913,N_19959);
xnor UO_1235 (O_1235,N_19811,N_19914);
nand UO_1236 (O_1236,N_19856,N_19970);
and UO_1237 (O_1237,N_19997,N_19998);
or UO_1238 (O_1238,N_19880,N_19910);
and UO_1239 (O_1239,N_19941,N_19960);
xnor UO_1240 (O_1240,N_19967,N_19936);
nor UO_1241 (O_1241,N_19822,N_19857);
or UO_1242 (O_1242,N_19995,N_19884);
and UO_1243 (O_1243,N_19827,N_19992);
or UO_1244 (O_1244,N_19968,N_19950);
xor UO_1245 (O_1245,N_19884,N_19853);
and UO_1246 (O_1246,N_19951,N_19855);
and UO_1247 (O_1247,N_19913,N_19800);
or UO_1248 (O_1248,N_19817,N_19980);
and UO_1249 (O_1249,N_19872,N_19847);
nand UO_1250 (O_1250,N_19911,N_19806);
nand UO_1251 (O_1251,N_19993,N_19982);
nor UO_1252 (O_1252,N_19980,N_19985);
nor UO_1253 (O_1253,N_19944,N_19864);
and UO_1254 (O_1254,N_19876,N_19964);
nand UO_1255 (O_1255,N_19917,N_19823);
nand UO_1256 (O_1256,N_19931,N_19965);
nor UO_1257 (O_1257,N_19893,N_19834);
nand UO_1258 (O_1258,N_19939,N_19984);
nand UO_1259 (O_1259,N_19995,N_19907);
xnor UO_1260 (O_1260,N_19811,N_19971);
or UO_1261 (O_1261,N_19817,N_19823);
and UO_1262 (O_1262,N_19900,N_19884);
xnor UO_1263 (O_1263,N_19882,N_19869);
nand UO_1264 (O_1264,N_19891,N_19951);
nand UO_1265 (O_1265,N_19957,N_19914);
or UO_1266 (O_1266,N_19800,N_19955);
nor UO_1267 (O_1267,N_19843,N_19874);
or UO_1268 (O_1268,N_19843,N_19833);
and UO_1269 (O_1269,N_19895,N_19875);
nor UO_1270 (O_1270,N_19999,N_19859);
nor UO_1271 (O_1271,N_19817,N_19951);
or UO_1272 (O_1272,N_19868,N_19827);
nor UO_1273 (O_1273,N_19821,N_19960);
or UO_1274 (O_1274,N_19896,N_19941);
and UO_1275 (O_1275,N_19932,N_19908);
nor UO_1276 (O_1276,N_19860,N_19942);
nor UO_1277 (O_1277,N_19924,N_19827);
and UO_1278 (O_1278,N_19850,N_19811);
nand UO_1279 (O_1279,N_19998,N_19953);
nor UO_1280 (O_1280,N_19817,N_19988);
or UO_1281 (O_1281,N_19898,N_19880);
or UO_1282 (O_1282,N_19901,N_19883);
or UO_1283 (O_1283,N_19816,N_19923);
xor UO_1284 (O_1284,N_19895,N_19840);
and UO_1285 (O_1285,N_19874,N_19815);
or UO_1286 (O_1286,N_19804,N_19822);
nand UO_1287 (O_1287,N_19946,N_19966);
or UO_1288 (O_1288,N_19817,N_19869);
xnor UO_1289 (O_1289,N_19919,N_19810);
or UO_1290 (O_1290,N_19953,N_19941);
nand UO_1291 (O_1291,N_19901,N_19984);
xnor UO_1292 (O_1292,N_19863,N_19921);
nor UO_1293 (O_1293,N_19957,N_19926);
nor UO_1294 (O_1294,N_19917,N_19869);
nand UO_1295 (O_1295,N_19900,N_19920);
or UO_1296 (O_1296,N_19902,N_19832);
nor UO_1297 (O_1297,N_19888,N_19862);
or UO_1298 (O_1298,N_19943,N_19984);
or UO_1299 (O_1299,N_19869,N_19946);
nand UO_1300 (O_1300,N_19955,N_19825);
and UO_1301 (O_1301,N_19908,N_19950);
nand UO_1302 (O_1302,N_19978,N_19877);
nor UO_1303 (O_1303,N_19838,N_19833);
and UO_1304 (O_1304,N_19942,N_19965);
nor UO_1305 (O_1305,N_19801,N_19922);
and UO_1306 (O_1306,N_19913,N_19805);
xor UO_1307 (O_1307,N_19883,N_19973);
nand UO_1308 (O_1308,N_19933,N_19969);
nand UO_1309 (O_1309,N_19902,N_19931);
nand UO_1310 (O_1310,N_19861,N_19961);
xor UO_1311 (O_1311,N_19807,N_19960);
nand UO_1312 (O_1312,N_19828,N_19975);
xnor UO_1313 (O_1313,N_19951,N_19812);
nand UO_1314 (O_1314,N_19875,N_19923);
nor UO_1315 (O_1315,N_19820,N_19898);
nand UO_1316 (O_1316,N_19934,N_19916);
nor UO_1317 (O_1317,N_19889,N_19904);
nor UO_1318 (O_1318,N_19975,N_19906);
and UO_1319 (O_1319,N_19927,N_19917);
xor UO_1320 (O_1320,N_19958,N_19982);
nand UO_1321 (O_1321,N_19811,N_19970);
xnor UO_1322 (O_1322,N_19891,N_19887);
nand UO_1323 (O_1323,N_19859,N_19960);
nand UO_1324 (O_1324,N_19932,N_19990);
and UO_1325 (O_1325,N_19908,N_19975);
or UO_1326 (O_1326,N_19806,N_19855);
nand UO_1327 (O_1327,N_19950,N_19825);
nor UO_1328 (O_1328,N_19909,N_19818);
or UO_1329 (O_1329,N_19901,N_19826);
nand UO_1330 (O_1330,N_19828,N_19976);
nor UO_1331 (O_1331,N_19978,N_19995);
or UO_1332 (O_1332,N_19994,N_19844);
nand UO_1333 (O_1333,N_19891,N_19903);
nand UO_1334 (O_1334,N_19803,N_19957);
and UO_1335 (O_1335,N_19929,N_19940);
xor UO_1336 (O_1336,N_19974,N_19890);
and UO_1337 (O_1337,N_19825,N_19971);
nor UO_1338 (O_1338,N_19873,N_19865);
nand UO_1339 (O_1339,N_19859,N_19923);
nand UO_1340 (O_1340,N_19916,N_19960);
nor UO_1341 (O_1341,N_19827,N_19871);
nor UO_1342 (O_1342,N_19830,N_19905);
nor UO_1343 (O_1343,N_19983,N_19923);
or UO_1344 (O_1344,N_19898,N_19979);
or UO_1345 (O_1345,N_19873,N_19958);
xor UO_1346 (O_1346,N_19919,N_19802);
and UO_1347 (O_1347,N_19911,N_19808);
and UO_1348 (O_1348,N_19995,N_19911);
and UO_1349 (O_1349,N_19980,N_19960);
nand UO_1350 (O_1350,N_19938,N_19905);
or UO_1351 (O_1351,N_19891,N_19838);
nor UO_1352 (O_1352,N_19843,N_19934);
xor UO_1353 (O_1353,N_19805,N_19813);
and UO_1354 (O_1354,N_19992,N_19884);
nand UO_1355 (O_1355,N_19867,N_19874);
nand UO_1356 (O_1356,N_19884,N_19980);
nand UO_1357 (O_1357,N_19966,N_19812);
or UO_1358 (O_1358,N_19853,N_19846);
nand UO_1359 (O_1359,N_19918,N_19866);
nand UO_1360 (O_1360,N_19986,N_19815);
nand UO_1361 (O_1361,N_19846,N_19838);
xor UO_1362 (O_1362,N_19944,N_19866);
nor UO_1363 (O_1363,N_19980,N_19908);
or UO_1364 (O_1364,N_19937,N_19967);
nor UO_1365 (O_1365,N_19856,N_19863);
or UO_1366 (O_1366,N_19931,N_19923);
xnor UO_1367 (O_1367,N_19985,N_19853);
nand UO_1368 (O_1368,N_19847,N_19923);
xnor UO_1369 (O_1369,N_19994,N_19909);
xnor UO_1370 (O_1370,N_19977,N_19888);
nand UO_1371 (O_1371,N_19965,N_19819);
xor UO_1372 (O_1372,N_19909,N_19958);
xnor UO_1373 (O_1373,N_19809,N_19854);
xor UO_1374 (O_1374,N_19843,N_19965);
nand UO_1375 (O_1375,N_19913,N_19837);
xor UO_1376 (O_1376,N_19963,N_19854);
nand UO_1377 (O_1377,N_19896,N_19831);
nor UO_1378 (O_1378,N_19810,N_19948);
and UO_1379 (O_1379,N_19905,N_19893);
nor UO_1380 (O_1380,N_19871,N_19986);
nor UO_1381 (O_1381,N_19994,N_19967);
nor UO_1382 (O_1382,N_19865,N_19957);
nand UO_1383 (O_1383,N_19948,N_19960);
nand UO_1384 (O_1384,N_19828,N_19805);
nand UO_1385 (O_1385,N_19920,N_19905);
xnor UO_1386 (O_1386,N_19823,N_19869);
or UO_1387 (O_1387,N_19992,N_19968);
nor UO_1388 (O_1388,N_19903,N_19940);
and UO_1389 (O_1389,N_19934,N_19901);
nor UO_1390 (O_1390,N_19868,N_19834);
and UO_1391 (O_1391,N_19895,N_19969);
or UO_1392 (O_1392,N_19817,N_19872);
nor UO_1393 (O_1393,N_19911,N_19809);
nor UO_1394 (O_1394,N_19957,N_19910);
xnor UO_1395 (O_1395,N_19956,N_19817);
nor UO_1396 (O_1396,N_19887,N_19982);
and UO_1397 (O_1397,N_19972,N_19924);
nor UO_1398 (O_1398,N_19985,N_19874);
and UO_1399 (O_1399,N_19938,N_19963);
or UO_1400 (O_1400,N_19959,N_19950);
or UO_1401 (O_1401,N_19949,N_19862);
or UO_1402 (O_1402,N_19912,N_19807);
nor UO_1403 (O_1403,N_19952,N_19842);
and UO_1404 (O_1404,N_19984,N_19814);
nand UO_1405 (O_1405,N_19987,N_19942);
xor UO_1406 (O_1406,N_19869,N_19825);
nand UO_1407 (O_1407,N_19813,N_19943);
xnor UO_1408 (O_1408,N_19817,N_19986);
or UO_1409 (O_1409,N_19811,N_19907);
nor UO_1410 (O_1410,N_19986,N_19974);
and UO_1411 (O_1411,N_19935,N_19813);
nand UO_1412 (O_1412,N_19968,N_19849);
nand UO_1413 (O_1413,N_19803,N_19961);
xnor UO_1414 (O_1414,N_19829,N_19995);
xnor UO_1415 (O_1415,N_19907,N_19850);
xnor UO_1416 (O_1416,N_19899,N_19923);
xor UO_1417 (O_1417,N_19814,N_19853);
nand UO_1418 (O_1418,N_19835,N_19817);
xor UO_1419 (O_1419,N_19822,N_19825);
or UO_1420 (O_1420,N_19813,N_19972);
and UO_1421 (O_1421,N_19951,N_19835);
xnor UO_1422 (O_1422,N_19807,N_19925);
or UO_1423 (O_1423,N_19977,N_19889);
or UO_1424 (O_1424,N_19958,N_19892);
or UO_1425 (O_1425,N_19838,N_19935);
nor UO_1426 (O_1426,N_19945,N_19826);
nor UO_1427 (O_1427,N_19895,N_19968);
nand UO_1428 (O_1428,N_19928,N_19978);
xnor UO_1429 (O_1429,N_19819,N_19834);
nor UO_1430 (O_1430,N_19981,N_19948);
nand UO_1431 (O_1431,N_19957,N_19967);
xnor UO_1432 (O_1432,N_19810,N_19942);
or UO_1433 (O_1433,N_19940,N_19961);
xor UO_1434 (O_1434,N_19843,N_19950);
nor UO_1435 (O_1435,N_19998,N_19877);
nand UO_1436 (O_1436,N_19913,N_19866);
xor UO_1437 (O_1437,N_19852,N_19963);
and UO_1438 (O_1438,N_19887,N_19820);
or UO_1439 (O_1439,N_19809,N_19868);
and UO_1440 (O_1440,N_19827,N_19973);
nor UO_1441 (O_1441,N_19916,N_19851);
nand UO_1442 (O_1442,N_19964,N_19873);
and UO_1443 (O_1443,N_19842,N_19820);
and UO_1444 (O_1444,N_19962,N_19869);
and UO_1445 (O_1445,N_19997,N_19917);
or UO_1446 (O_1446,N_19815,N_19971);
nor UO_1447 (O_1447,N_19966,N_19981);
nand UO_1448 (O_1448,N_19900,N_19877);
or UO_1449 (O_1449,N_19858,N_19960);
and UO_1450 (O_1450,N_19908,N_19946);
or UO_1451 (O_1451,N_19986,N_19882);
nand UO_1452 (O_1452,N_19837,N_19827);
or UO_1453 (O_1453,N_19980,N_19888);
nand UO_1454 (O_1454,N_19843,N_19838);
and UO_1455 (O_1455,N_19902,N_19952);
xnor UO_1456 (O_1456,N_19817,N_19926);
xnor UO_1457 (O_1457,N_19903,N_19946);
xor UO_1458 (O_1458,N_19894,N_19941);
or UO_1459 (O_1459,N_19976,N_19863);
and UO_1460 (O_1460,N_19897,N_19892);
xnor UO_1461 (O_1461,N_19884,N_19926);
or UO_1462 (O_1462,N_19829,N_19877);
xnor UO_1463 (O_1463,N_19931,N_19804);
nand UO_1464 (O_1464,N_19923,N_19997);
xor UO_1465 (O_1465,N_19988,N_19825);
nor UO_1466 (O_1466,N_19936,N_19863);
xnor UO_1467 (O_1467,N_19805,N_19829);
and UO_1468 (O_1468,N_19801,N_19991);
nor UO_1469 (O_1469,N_19899,N_19982);
or UO_1470 (O_1470,N_19840,N_19948);
nor UO_1471 (O_1471,N_19832,N_19993);
nor UO_1472 (O_1472,N_19993,N_19920);
or UO_1473 (O_1473,N_19884,N_19835);
and UO_1474 (O_1474,N_19969,N_19913);
or UO_1475 (O_1475,N_19843,N_19947);
nor UO_1476 (O_1476,N_19875,N_19901);
nand UO_1477 (O_1477,N_19999,N_19898);
or UO_1478 (O_1478,N_19863,N_19965);
xnor UO_1479 (O_1479,N_19932,N_19973);
nor UO_1480 (O_1480,N_19896,N_19968);
nor UO_1481 (O_1481,N_19984,N_19904);
nor UO_1482 (O_1482,N_19935,N_19956);
xor UO_1483 (O_1483,N_19816,N_19961);
and UO_1484 (O_1484,N_19967,N_19902);
nor UO_1485 (O_1485,N_19866,N_19928);
or UO_1486 (O_1486,N_19803,N_19804);
nor UO_1487 (O_1487,N_19827,N_19815);
nand UO_1488 (O_1488,N_19826,N_19958);
nor UO_1489 (O_1489,N_19814,N_19921);
nand UO_1490 (O_1490,N_19816,N_19905);
nand UO_1491 (O_1491,N_19980,N_19904);
xnor UO_1492 (O_1492,N_19880,N_19973);
or UO_1493 (O_1493,N_19823,N_19856);
or UO_1494 (O_1494,N_19979,N_19803);
xnor UO_1495 (O_1495,N_19876,N_19911);
and UO_1496 (O_1496,N_19981,N_19959);
nand UO_1497 (O_1497,N_19931,N_19870);
nor UO_1498 (O_1498,N_19980,N_19868);
xnor UO_1499 (O_1499,N_19956,N_19910);
nand UO_1500 (O_1500,N_19941,N_19897);
and UO_1501 (O_1501,N_19819,N_19961);
xnor UO_1502 (O_1502,N_19868,N_19894);
nor UO_1503 (O_1503,N_19977,N_19999);
nor UO_1504 (O_1504,N_19868,N_19905);
or UO_1505 (O_1505,N_19841,N_19995);
nor UO_1506 (O_1506,N_19986,N_19822);
and UO_1507 (O_1507,N_19810,N_19889);
nor UO_1508 (O_1508,N_19887,N_19938);
xor UO_1509 (O_1509,N_19867,N_19912);
nor UO_1510 (O_1510,N_19895,N_19896);
nor UO_1511 (O_1511,N_19951,N_19824);
nor UO_1512 (O_1512,N_19884,N_19901);
xor UO_1513 (O_1513,N_19819,N_19960);
and UO_1514 (O_1514,N_19913,N_19806);
and UO_1515 (O_1515,N_19935,N_19981);
or UO_1516 (O_1516,N_19821,N_19869);
and UO_1517 (O_1517,N_19963,N_19989);
or UO_1518 (O_1518,N_19809,N_19838);
xnor UO_1519 (O_1519,N_19955,N_19809);
xor UO_1520 (O_1520,N_19847,N_19897);
nor UO_1521 (O_1521,N_19834,N_19924);
nor UO_1522 (O_1522,N_19879,N_19814);
and UO_1523 (O_1523,N_19862,N_19842);
nor UO_1524 (O_1524,N_19989,N_19809);
xor UO_1525 (O_1525,N_19935,N_19884);
nand UO_1526 (O_1526,N_19850,N_19916);
nor UO_1527 (O_1527,N_19925,N_19948);
xnor UO_1528 (O_1528,N_19956,N_19858);
and UO_1529 (O_1529,N_19868,N_19915);
nor UO_1530 (O_1530,N_19908,N_19851);
or UO_1531 (O_1531,N_19875,N_19804);
or UO_1532 (O_1532,N_19859,N_19974);
and UO_1533 (O_1533,N_19890,N_19802);
and UO_1534 (O_1534,N_19915,N_19935);
and UO_1535 (O_1535,N_19998,N_19977);
and UO_1536 (O_1536,N_19955,N_19877);
and UO_1537 (O_1537,N_19881,N_19910);
nand UO_1538 (O_1538,N_19883,N_19809);
xnor UO_1539 (O_1539,N_19804,N_19883);
xor UO_1540 (O_1540,N_19908,N_19819);
nor UO_1541 (O_1541,N_19825,N_19897);
nor UO_1542 (O_1542,N_19933,N_19929);
or UO_1543 (O_1543,N_19963,N_19808);
xnor UO_1544 (O_1544,N_19875,N_19964);
xor UO_1545 (O_1545,N_19939,N_19905);
or UO_1546 (O_1546,N_19869,N_19948);
nor UO_1547 (O_1547,N_19820,N_19901);
or UO_1548 (O_1548,N_19864,N_19971);
nor UO_1549 (O_1549,N_19804,N_19865);
nor UO_1550 (O_1550,N_19927,N_19824);
nand UO_1551 (O_1551,N_19905,N_19937);
or UO_1552 (O_1552,N_19936,N_19824);
nor UO_1553 (O_1553,N_19908,N_19916);
nor UO_1554 (O_1554,N_19965,N_19807);
and UO_1555 (O_1555,N_19894,N_19895);
or UO_1556 (O_1556,N_19902,N_19895);
xor UO_1557 (O_1557,N_19977,N_19978);
and UO_1558 (O_1558,N_19973,N_19925);
nand UO_1559 (O_1559,N_19884,N_19943);
and UO_1560 (O_1560,N_19959,N_19922);
nor UO_1561 (O_1561,N_19950,N_19868);
or UO_1562 (O_1562,N_19843,N_19848);
and UO_1563 (O_1563,N_19808,N_19980);
nor UO_1564 (O_1564,N_19895,N_19994);
nor UO_1565 (O_1565,N_19911,N_19847);
and UO_1566 (O_1566,N_19905,N_19991);
nor UO_1567 (O_1567,N_19908,N_19900);
xnor UO_1568 (O_1568,N_19821,N_19927);
xor UO_1569 (O_1569,N_19901,N_19807);
xnor UO_1570 (O_1570,N_19910,N_19962);
nand UO_1571 (O_1571,N_19932,N_19887);
nor UO_1572 (O_1572,N_19992,N_19975);
nand UO_1573 (O_1573,N_19839,N_19992);
nor UO_1574 (O_1574,N_19921,N_19941);
and UO_1575 (O_1575,N_19957,N_19815);
nor UO_1576 (O_1576,N_19988,N_19898);
or UO_1577 (O_1577,N_19808,N_19890);
nand UO_1578 (O_1578,N_19889,N_19909);
or UO_1579 (O_1579,N_19984,N_19967);
and UO_1580 (O_1580,N_19888,N_19870);
or UO_1581 (O_1581,N_19908,N_19952);
and UO_1582 (O_1582,N_19975,N_19885);
xnor UO_1583 (O_1583,N_19998,N_19852);
or UO_1584 (O_1584,N_19972,N_19818);
nor UO_1585 (O_1585,N_19920,N_19954);
and UO_1586 (O_1586,N_19810,N_19892);
or UO_1587 (O_1587,N_19944,N_19819);
or UO_1588 (O_1588,N_19969,N_19924);
nand UO_1589 (O_1589,N_19821,N_19804);
nor UO_1590 (O_1590,N_19944,N_19899);
xor UO_1591 (O_1591,N_19850,N_19844);
xor UO_1592 (O_1592,N_19842,N_19980);
and UO_1593 (O_1593,N_19836,N_19984);
nand UO_1594 (O_1594,N_19919,N_19923);
nand UO_1595 (O_1595,N_19988,N_19910);
nand UO_1596 (O_1596,N_19912,N_19973);
and UO_1597 (O_1597,N_19958,N_19951);
xor UO_1598 (O_1598,N_19978,N_19933);
xor UO_1599 (O_1599,N_19899,N_19894);
xnor UO_1600 (O_1600,N_19885,N_19870);
or UO_1601 (O_1601,N_19973,N_19826);
nor UO_1602 (O_1602,N_19846,N_19899);
nand UO_1603 (O_1603,N_19890,N_19839);
xnor UO_1604 (O_1604,N_19938,N_19897);
nor UO_1605 (O_1605,N_19858,N_19892);
xnor UO_1606 (O_1606,N_19922,N_19966);
xor UO_1607 (O_1607,N_19902,N_19813);
xor UO_1608 (O_1608,N_19916,N_19849);
xor UO_1609 (O_1609,N_19971,N_19871);
xnor UO_1610 (O_1610,N_19895,N_19958);
and UO_1611 (O_1611,N_19913,N_19998);
nor UO_1612 (O_1612,N_19889,N_19951);
and UO_1613 (O_1613,N_19846,N_19938);
nand UO_1614 (O_1614,N_19992,N_19891);
or UO_1615 (O_1615,N_19849,N_19908);
and UO_1616 (O_1616,N_19995,N_19876);
nor UO_1617 (O_1617,N_19947,N_19806);
or UO_1618 (O_1618,N_19883,N_19912);
nand UO_1619 (O_1619,N_19896,N_19947);
or UO_1620 (O_1620,N_19908,N_19974);
or UO_1621 (O_1621,N_19915,N_19991);
nor UO_1622 (O_1622,N_19852,N_19870);
and UO_1623 (O_1623,N_19905,N_19865);
and UO_1624 (O_1624,N_19837,N_19859);
or UO_1625 (O_1625,N_19910,N_19941);
or UO_1626 (O_1626,N_19984,N_19860);
xor UO_1627 (O_1627,N_19884,N_19819);
nand UO_1628 (O_1628,N_19902,N_19921);
xnor UO_1629 (O_1629,N_19834,N_19926);
nand UO_1630 (O_1630,N_19858,N_19860);
nand UO_1631 (O_1631,N_19913,N_19966);
or UO_1632 (O_1632,N_19956,N_19946);
or UO_1633 (O_1633,N_19872,N_19932);
nand UO_1634 (O_1634,N_19843,N_19907);
nand UO_1635 (O_1635,N_19924,N_19896);
or UO_1636 (O_1636,N_19824,N_19924);
nand UO_1637 (O_1637,N_19975,N_19973);
xor UO_1638 (O_1638,N_19974,N_19867);
or UO_1639 (O_1639,N_19963,N_19860);
xor UO_1640 (O_1640,N_19817,N_19917);
nor UO_1641 (O_1641,N_19851,N_19828);
or UO_1642 (O_1642,N_19842,N_19880);
nand UO_1643 (O_1643,N_19951,N_19942);
or UO_1644 (O_1644,N_19819,N_19824);
nand UO_1645 (O_1645,N_19882,N_19910);
xor UO_1646 (O_1646,N_19857,N_19808);
or UO_1647 (O_1647,N_19819,N_19913);
nand UO_1648 (O_1648,N_19876,N_19809);
nor UO_1649 (O_1649,N_19899,N_19863);
xnor UO_1650 (O_1650,N_19957,N_19952);
or UO_1651 (O_1651,N_19827,N_19890);
or UO_1652 (O_1652,N_19957,N_19810);
nand UO_1653 (O_1653,N_19807,N_19854);
and UO_1654 (O_1654,N_19884,N_19811);
or UO_1655 (O_1655,N_19822,N_19834);
nand UO_1656 (O_1656,N_19964,N_19806);
and UO_1657 (O_1657,N_19987,N_19908);
xnor UO_1658 (O_1658,N_19981,N_19830);
nor UO_1659 (O_1659,N_19945,N_19935);
xor UO_1660 (O_1660,N_19833,N_19969);
nor UO_1661 (O_1661,N_19913,N_19896);
or UO_1662 (O_1662,N_19857,N_19938);
or UO_1663 (O_1663,N_19817,N_19837);
xnor UO_1664 (O_1664,N_19975,N_19934);
xor UO_1665 (O_1665,N_19927,N_19851);
nand UO_1666 (O_1666,N_19843,N_19879);
nand UO_1667 (O_1667,N_19915,N_19992);
and UO_1668 (O_1668,N_19949,N_19917);
nor UO_1669 (O_1669,N_19982,N_19855);
nor UO_1670 (O_1670,N_19922,N_19946);
nand UO_1671 (O_1671,N_19817,N_19800);
xor UO_1672 (O_1672,N_19938,N_19866);
or UO_1673 (O_1673,N_19939,N_19975);
xor UO_1674 (O_1674,N_19913,N_19957);
or UO_1675 (O_1675,N_19924,N_19802);
xnor UO_1676 (O_1676,N_19892,N_19974);
xor UO_1677 (O_1677,N_19899,N_19996);
nand UO_1678 (O_1678,N_19875,N_19918);
xor UO_1679 (O_1679,N_19884,N_19928);
nor UO_1680 (O_1680,N_19922,N_19816);
and UO_1681 (O_1681,N_19896,N_19956);
and UO_1682 (O_1682,N_19874,N_19884);
or UO_1683 (O_1683,N_19994,N_19904);
or UO_1684 (O_1684,N_19955,N_19897);
xor UO_1685 (O_1685,N_19956,N_19836);
nor UO_1686 (O_1686,N_19965,N_19921);
and UO_1687 (O_1687,N_19849,N_19822);
and UO_1688 (O_1688,N_19845,N_19818);
or UO_1689 (O_1689,N_19815,N_19949);
nand UO_1690 (O_1690,N_19863,N_19864);
or UO_1691 (O_1691,N_19825,N_19860);
and UO_1692 (O_1692,N_19877,N_19963);
or UO_1693 (O_1693,N_19869,N_19979);
nand UO_1694 (O_1694,N_19954,N_19982);
or UO_1695 (O_1695,N_19814,N_19802);
nand UO_1696 (O_1696,N_19818,N_19833);
and UO_1697 (O_1697,N_19968,N_19825);
or UO_1698 (O_1698,N_19901,N_19938);
nor UO_1699 (O_1699,N_19988,N_19824);
and UO_1700 (O_1700,N_19904,N_19915);
and UO_1701 (O_1701,N_19864,N_19867);
nor UO_1702 (O_1702,N_19901,N_19813);
nor UO_1703 (O_1703,N_19989,N_19973);
xnor UO_1704 (O_1704,N_19950,N_19864);
xor UO_1705 (O_1705,N_19907,N_19832);
nor UO_1706 (O_1706,N_19965,N_19839);
nor UO_1707 (O_1707,N_19912,N_19946);
or UO_1708 (O_1708,N_19904,N_19886);
nand UO_1709 (O_1709,N_19966,N_19931);
xor UO_1710 (O_1710,N_19996,N_19867);
or UO_1711 (O_1711,N_19929,N_19956);
or UO_1712 (O_1712,N_19948,N_19880);
nand UO_1713 (O_1713,N_19876,N_19825);
xor UO_1714 (O_1714,N_19829,N_19879);
nand UO_1715 (O_1715,N_19971,N_19865);
xnor UO_1716 (O_1716,N_19913,N_19975);
xor UO_1717 (O_1717,N_19989,N_19895);
nor UO_1718 (O_1718,N_19805,N_19933);
nand UO_1719 (O_1719,N_19863,N_19957);
nor UO_1720 (O_1720,N_19926,N_19907);
or UO_1721 (O_1721,N_19983,N_19858);
or UO_1722 (O_1722,N_19957,N_19921);
nor UO_1723 (O_1723,N_19914,N_19916);
and UO_1724 (O_1724,N_19890,N_19962);
xnor UO_1725 (O_1725,N_19837,N_19890);
and UO_1726 (O_1726,N_19818,N_19877);
and UO_1727 (O_1727,N_19979,N_19835);
nor UO_1728 (O_1728,N_19902,N_19841);
nand UO_1729 (O_1729,N_19961,N_19937);
xor UO_1730 (O_1730,N_19883,N_19992);
xnor UO_1731 (O_1731,N_19941,N_19998);
nor UO_1732 (O_1732,N_19935,N_19959);
nand UO_1733 (O_1733,N_19936,N_19889);
xnor UO_1734 (O_1734,N_19924,N_19910);
xnor UO_1735 (O_1735,N_19997,N_19913);
nor UO_1736 (O_1736,N_19984,N_19882);
and UO_1737 (O_1737,N_19966,N_19977);
and UO_1738 (O_1738,N_19993,N_19855);
and UO_1739 (O_1739,N_19862,N_19934);
or UO_1740 (O_1740,N_19926,N_19881);
and UO_1741 (O_1741,N_19958,N_19827);
nand UO_1742 (O_1742,N_19892,N_19942);
nor UO_1743 (O_1743,N_19938,N_19825);
and UO_1744 (O_1744,N_19961,N_19971);
nor UO_1745 (O_1745,N_19976,N_19854);
and UO_1746 (O_1746,N_19848,N_19943);
xor UO_1747 (O_1747,N_19845,N_19904);
nand UO_1748 (O_1748,N_19923,N_19975);
and UO_1749 (O_1749,N_19930,N_19967);
nor UO_1750 (O_1750,N_19906,N_19912);
or UO_1751 (O_1751,N_19911,N_19958);
and UO_1752 (O_1752,N_19903,N_19907);
and UO_1753 (O_1753,N_19959,N_19825);
nand UO_1754 (O_1754,N_19945,N_19980);
and UO_1755 (O_1755,N_19832,N_19984);
or UO_1756 (O_1756,N_19822,N_19912);
xnor UO_1757 (O_1757,N_19880,N_19859);
and UO_1758 (O_1758,N_19896,N_19855);
nand UO_1759 (O_1759,N_19954,N_19887);
nor UO_1760 (O_1760,N_19958,N_19923);
nor UO_1761 (O_1761,N_19975,N_19802);
nor UO_1762 (O_1762,N_19836,N_19832);
nand UO_1763 (O_1763,N_19906,N_19890);
nor UO_1764 (O_1764,N_19899,N_19999);
nor UO_1765 (O_1765,N_19895,N_19948);
nor UO_1766 (O_1766,N_19993,N_19843);
xnor UO_1767 (O_1767,N_19912,N_19938);
xnor UO_1768 (O_1768,N_19890,N_19899);
xnor UO_1769 (O_1769,N_19925,N_19861);
nand UO_1770 (O_1770,N_19977,N_19988);
xor UO_1771 (O_1771,N_19836,N_19856);
and UO_1772 (O_1772,N_19916,N_19874);
or UO_1773 (O_1773,N_19904,N_19849);
or UO_1774 (O_1774,N_19990,N_19969);
or UO_1775 (O_1775,N_19882,N_19905);
xor UO_1776 (O_1776,N_19849,N_19976);
nand UO_1777 (O_1777,N_19945,N_19974);
nor UO_1778 (O_1778,N_19983,N_19877);
nor UO_1779 (O_1779,N_19982,N_19809);
xor UO_1780 (O_1780,N_19845,N_19945);
and UO_1781 (O_1781,N_19998,N_19823);
nor UO_1782 (O_1782,N_19915,N_19964);
xnor UO_1783 (O_1783,N_19877,N_19931);
or UO_1784 (O_1784,N_19901,N_19992);
nor UO_1785 (O_1785,N_19909,N_19918);
or UO_1786 (O_1786,N_19865,N_19958);
nor UO_1787 (O_1787,N_19917,N_19857);
xor UO_1788 (O_1788,N_19989,N_19897);
nand UO_1789 (O_1789,N_19985,N_19820);
nor UO_1790 (O_1790,N_19909,N_19830);
or UO_1791 (O_1791,N_19825,N_19879);
nor UO_1792 (O_1792,N_19803,N_19901);
and UO_1793 (O_1793,N_19985,N_19813);
or UO_1794 (O_1794,N_19904,N_19966);
xor UO_1795 (O_1795,N_19891,N_19986);
nor UO_1796 (O_1796,N_19857,N_19921);
xnor UO_1797 (O_1797,N_19810,N_19875);
xnor UO_1798 (O_1798,N_19945,N_19966);
nor UO_1799 (O_1799,N_19816,N_19897);
or UO_1800 (O_1800,N_19931,N_19906);
nand UO_1801 (O_1801,N_19977,N_19894);
or UO_1802 (O_1802,N_19869,N_19964);
nor UO_1803 (O_1803,N_19943,N_19999);
and UO_1804 (O_1804,N_19839,N_19896);
xnor UO_1805 (O_1805,N_19802,N_19858);
xor UO_1806 (O_1806,N_19802,N_19888);
nor UO_1807 (O_1807,N_19931,N_19800);
nor UO_1808 (O_1808,N_19906,N_19873);
nor UO_1809 (O_1809,N_19858,N_19813);
xor UO_1810 (O_1810,N_19955,N_19999);
xnor UO_1811 (O_1811,N_19931,N_19991);
nand UO_1812 (O_1812,N_19875,N_19856);
or UO_1813 (O_1813,N_19921,N_19981);
and UO_1814 (O_1814,N_19901,N_19898);
xnor UO_1815 (O_1815,N_19854,N_19988);
nand UO_1816 (O_1816,N_19994,N_19955);
nor UO_1817 (O_1817,N_19821,N_19863);
nor UO_1818 (O_1818,N_19952,N_19810);
and UO_1819 (O_1819,N_19904,N_19931);
nand UO_1820 (O_1820,N_19860,N_19946);
xor UO_1821 (O_1821,N_19859,N_19907);
xor UO_1822 (O_1822,N_19937,N_19959);
xnor UO_1823 (O_1823,N_19957,N_19985);
nand UO_1824 (O_1824,N_19803,N_19832);
and UO_1825 (O_1825,N_19851,N_19984);
or UO_1826 (O_1826,N_19830,N_19972);
or UO_1827 (O_1827,N_19984,N_19820);
and UO_1828 (O_1828,N_19892,N_19989);
or UO_1829 (O_1829,N_19949,N_19855);
nand UO_1830 (O_1830,N_19994,N_19963);
nand UO_1831 (O_1831,N_19972,N_19863);
xnor UO_1832 (O_1832,N_19950,N_19870);
nor UO_1833 (O_1833,N_19930,N_19841);
and UO_1834 (O_1834,N_19918,N_19869);
xor UO_1835 (O_1835,N_19850,N_19861);
and UO_1836 (O_1836,N_19934,N_19814);
xnor UO_1837 (O_1837,N_19887,N_19854);
nor UO_1838 (O_1838,N_19899,N_19861);
nor UO_1839 (O_1839,N_19995,N_19964);
xnor UO_1840 (O_1840,N_19963,N_19956);
and UO_1841 (O_1841,N_19852,N_19888);
xor UO_1842 (O_1842,N_19874,N_19931);
and UO_1843 (O_1843,N_19901,N_19802);
or UO_1844 (O_1844,N_19837,N_19902);
xnor UO_1845 (O_1845,N_19845,N_19875);
and UO_1846 (O_1846,N_19946,N_19818);
xor UO_1847 (O_1847,N_19867,N_19894);
xnor UO_1848 (O_1848,N_19891,N_19820);
nand UO_1849 (O_1849,N_19922,N_19822);
nand UO_1850 (O_1850,N_19860,N_19896);
xnor UO_1851 (O_1851,N_19830,N_19919);
xor UO_1852 (O_1852,N_19909,N_19933);
nor UO_1853 (O_1853,N_19853,N_19823);
xor UO_1854 (O_1854,N_19880,N_19818);
xor UO_1855 (O_1855,N_19827,N_19845);
and UO_1856 (O_1856,N_19836,N_19996);
and UO_1857 (O_1857,N_19820,N_19941);
xor UO_1858 (O_1858,N_19961,N_19896);
nor UO_1859 (O_1859,N_19984,N_19924);
nand UO_1860 (O_1860,N_19952,N_19899);
nand UO_1861 (O_1861,N_19913,N_19994);
nor UO_1862 (O_1862,N_19852,N_19967);
nand UO_1863 (O_1863,N_19831,N_19836);
or UO_1864 (O_1864,N_19812,N_19855);
xnor UO_1865 (O_1865,N_19920,N_19844);
xnor UO_1866 (O_1866,N_19944,N_19992);
xor UO_1867 (O_1867,N_19864,N_19892);
and UO_1868 (O_1868,N_19934,N_19867);
nand UO_1869 (O_1869,N_19830,N_19862);
nor UO_1870 (O_1870,N_19855,N_19801);
xnor UO_1871 (O_1871,N_19803,N_19971);
nor UO_1872 (O_1872,N_19844,N_19926);
xor UO_1873 (O_1873,N_19967,N_19966);
or UO_1874 (O_1874,N_19817,N_19830);
and UO_1875 (O_1875,N_19973,N_19889);
nor UO_1876 (O_1876,N_19842,N_19853);
nand UO_1877 (O_1877,N_19838,N_19967);
or UO_1878 (O_1878,N_19816,N_19834);
or UO_1879 (O_1879,N_19925,N_19987);
xnor UO_1880 (O_1880,N_19821,N_19862);
or UO_1881 (O_1881,N_19901,N_19841);
and UO_1882 (O_1882,N_19893,N_19957);
or UO_1883 (O_1883,N_19946,N_19837);
xnor UO_1884 (O_1884,N_19992,N_19856);
or UO_1885 (O_1885,N_19868,N_19946);
xor UO_1886 (O_1886,N_19865,N_19986);
nand UO_1887 (O_1887,N_19923,N_19905);
or UO_1888 (O_1888,N_19819,N_19962);
nand UO_1889 (O_1889,N_19886,N_19887);
nor UO_1890 (O_1890,N_19995,N_19881);
and UO_1891 (O_1891,N_19886,N_19860);
or UO_1892 (O_1892,N_19988,N_19944);
and UO_1893 (O_1893,N_19969,N_19916);
and UO_1894 (O_1894,N_19810,N_19834);
nand UO_1895 (O_1895,N_19883,N_19939);
and UO_1896 (O_1896,N_19814,N_19933);
or UO_1897 (O_1897,N_19809,N_19977);
and UO_1898 (O_1898,N_19814,N_19926);
nor UO_1899 (O_1899,N_19804,N_19854);
or UO_1900 (O_1900,N_19845,N_19931);
or UO_1901 (O_1901,N_19865,N_19859);
nand UO_1902 (O_1902,N_19895,N_19878);
nor UO_1903 (O_1903,N_19895,N_19800);
and UO_1904 (O_1904,N_19932,N_19807);
or UO_1905 (O_1905,N_19844,N_19993);
or UO_1906 (O_1906,N_19919,N_19856);
or UO_1907 (O_1907,N_19809,N_19879);
xor UO_1908 (O_1908,N_19872,N_19825);
or UO_1909 (O_1909,N_19978,N_19908);
and UO_1910 (O_1910,N_19929,N_19903);
nor UO_1911 (O_1911,N_19946,N_19827);
nand UO_1912 (O_1912,N_19830,N_19958);
and UO_1913 (O_1913,N_19906,N_19959);
nand UO_1914 (O_1914,N_19977,N_19924);
xor UO_1915 (O_1915,N_19973,N_19815);
nand UO_1916 (O_1916,N_19919,N_19818);
or UO_1917 (O_1917,N_19864,N_19872);
and UO_1918 (O_1918,N_19877,N_19879);
nand UO_1919 (O_1919,N_19971,N_19855);
nand UO_1920 (O_1920,N_19802,N_19884);
nor UO_1921 (O_1921,N_19926,N_19975);
or UO_1922 (O_1922,N_19919,N_19820);
and UO_1923 (O_1923,N_19966,N_19800);
xnor UO_1924 (O_1924,N_19990,N_19804);
nor UO_1925 (O_1925,N_19911,N_19813);
nor UO_1926 (O_1926,N_19918,N_19858);
or UO_1927 (O_1927,N_19936,N_19975);
nor UO_1928 (O_1928,N_19921,N_19861);
nand UO_1929 (O_1929,N_19987,N_19807);
or UO_1930 (O_1930,N_19989,N_19943);
nor UO_1931 (O_1931,N_19939,N_19979);
nor UO_1932 (O_1932,N_19961,N_19853);
nand UO_1933 (O_1933,N_19988,N_19920);
nand UO_1934 (O_1934,N_19969,N_19874);
xnor UO_1935 (O_1935,N_19907,N_19983);
nor UO_1936 (O_1936,N_19814,N_19999);
nand UO_1937 (O_1937,N_19831,N_19829);
nor UO_1938 (O_1938,N_19834,N_19800);
nor UO_1939 (O_1939,N_19840,N_19808);
or UO_1940 (O_1940,N_19884,N_19872);
and UO_1941 (O_1941,N_19917,N_19893);
nand UO_1942 (O_1942,N_19864,N_19805);
or UO_1943 (O_1943,N_19950,N_19972);
nor UO_1944 (O_1944,N_19801,N_19918);
xnor UO_1945 (O_1945,N_19809,N_19938);
nor UO_1946 (O_1946,N_19818,N_19838);
and UO_1947 (O_1947,N_19912,N_19978);
or UO_1948 (O_1948,N_19889,N_19966);
and UO_1949 (O_1949,N_19971,N_19957);
nor UO_1950 (O_1950,N_19935,N_19926);
nor UO_1951 (O_1951,N_19806,N_19844);
xnor UO_1952 (O_1952,N_19993,N_19910);
nand UO_1953 (O_1953,N_19807,N_19945);
xnor UO_1954 (O_1954,N_19895,N_19880);
and UO_1955 (O_1955,N_19943,N_19852);
xnor UO_1956 (O_1956,N_19913,N_19826);
nor UO_1957 (O_1957,N_19837,N_19970);
nand UO_1958 (O_1958,N_19878,N_19802);
nand UO_1959 (O_1959,N_19876,N_19957);
and UO_1960 (O_1960,N_19873,N_19859);
and UO_1961 (O_1961,N_19974,N_19899);
and UO_1962 (O_1962,N_19849,N_19943);
or UO_1963 (O_1963,N_19939,N_19894);
nor UO_1964 (O_1964,N_19846,N_19801);
nor UO_1965 (O_1965,N_19815,N_19923);
nand UO_1966 (O_1966,N_19833,N_19952);
xor UO_1967 (O_1967,N_19879,N_19891);
nor UO_1968 (O_1968,N_19848,N_19879);
and UO_1969 (O_1969,N_19885,N_19883);
xnor UO_1970 (O_1970,N_19976,N_19862);
xor UO_1971 (O_1971,N_19915,N_19861);
nand UO_1972 (O_1972,N_19849,N_19828);
xor UO_1973 (O_1973,N_19848,N_19962);
nand UO_1974 (O_1974,N_19876,N_19823);
nor UO_1975 (O_1975,N_19847,N_19890);
and UO_1976 (O_1976,N_19856,N_19932);
nand UO_1977 (O_1977,N_19875,N_19849);
and UO_1978 (O_1978,N_19815,N_19848);
and UO_1979 (O_1979,N_19881,N_19930);
nand UO_1980 (O_1980,N_19895,N_19962);
xnor UO_1981 (O_1981,N_19811,N_19904);
and UO_1982 (O_1982,N_19949,N_19942);
xor UO_1983 (O_1983,N_19815,N_19817);
nor UO_1984 (O_1984,N_19986,N_19953);
nand UO_1985 (O_1985,N_19945,N_19840);
and UO_1986 (O_1986,N_19813,N_19976);
and UO_1987 (O_1987,N_19896,N_19898);
or UO_1988 (O_1988,N_19973,N_19858);
xnor UO_1989 (O_1989,N_19854,N_19962);
or UO_1990 (O_1990,N_19894,N_19888);
nand UO_1991 (O_1991,N_19894,N_19833);
xnor UO_1992 (O_1992,N_19934,N_19985);
nand UO_1993 (O_1993,N_19959,N_19946);
and UO_1994 (O_1994,N_19858,N_19948);
and UO_1995 (O_1995,N_19835,N_19988);
xor UO_1996 (O_1996,N_19961,N_19899);
nor UO_1997 (O_1997,N_19939,N_19832);
or UO_1998 (O_1998,N_19825,N_19980);
nor UO_1999 (O_1999,N_19817,N_19853);
nand UO_2000 (O_2000,N_19859,N_19883);
and UO_2001 (O_2001,N_19859,N_19958);
or UO_2002 (O_2002,N_19929,N_19920);
nand UO_2003 (O_2003,N_19919,N_19983);
nor UO_2004 (O_2004,N_19857,N_19836);
or UO_2005 (O_2005,N_19834,N_19869);
or UO_2006 (O_2006,N_19931,N_19895);
nor UO_2007 (O_2007,N_19836,N_19992);
xnor UO_2008 (O_2008,N_19934,N_19805);
nand UO_2009 (O_2009,N_19805,N_19891);
or UO_2010 (O_2010,N_19951,N_19955);
nor UO_2011 (O_2011,N_19887,N_19812);
nor UO_2012 (O_2012,N_19885,N_19876);
and UO_2013 (O_2013,N_19887,N_19811);
or UO_2014 (O_2014,N_19856,N_19834);
nand UO_2015 (O_2015,N_19990,N_19943);
nor UO_2016 (O_2016,N_19934,N_19970);
nand UO_2017 (O_2017,N_19809,N_19899);
or UO_2018 (O_2018,N_19900,N_19959);
or UO_2019 (O_2019,N_19995,N_19827);
or UO_2020 (O_2020,N_19897,N_19823);
and UO_2021 (O_2021,N_19976,N_19884);
nand UO_2022 (O_2022,N_19828,N_19803);
nor UO_2023 (O_2023,N_19839,N_19994);
nor UO_2024 (O_2024,N_19906,N_19933);
and UO_2025 (O_2025,N_19929,N_19880);
xnor UO_2026 (O_2026,N_19828,N_19902);
and UO_2027 (O_2027,N_19826,N_19892);
nand UO_2028 (O_2028,N_19896,N_19912);
and UO_2029 (O_2029,N_19933,N_19965);
xor UO_2030 (O_2030,N_19964,N_19937);
or UO_2031 (O_2031,N_19917,N_19957);
nand UO_2032 (O_2032,N_19829,N_19957);
or UO_2033 (O_2033,N_19978,N_19849);
nand UO_2034 (O_2034,N_19884,N_19868);
or UO_2035 (O_2035,N_19848,N_19956);
and UO_2036 (O_2036,N_19945,N_19877);
nor UO_2037 (O_2037,N_19960,N_19833);
or UO_2038 (O_2038,N_19928,N_19837);
or UO_2039 (O_2039,N_19855,N_19889);
or UO_2040 (O_2040,N_19994,N_19896);
and UO_2041 (O_2041,N_19982,N_19910);
or UO_2042 (O_2042,N_19921,N_19884);
nor UO_2043 (O_2043,N_19904,N_19995);
xnor UO_2044 (O_2044,N_19830,N_19858);
nand UO_2045 (O_2045,N_19924,N_19825);
nor UO_2046 (O_2046,N_19957,N_19844);
nand UO_2047 (O_2047,N_19965,N_19831);
and UO_2048 (O_2048,N_19905,N_19800);
nor UO_2049 (O_2049,N_19802,N_19874);
nand UO_2050 (O_2050,N_19991,N_19862);
xor UO_2051 (O_2051,N_19846,N_19901);
or UO_2052 (O_2052,N_19957,N_19834);
xor UO_2053 (O_2053,N_19977,N_19910);
nor UO_2054 (O_2054,N_19907,N_19817);
or UO_2055 (O_2055,N_19860,N_19996);
xnor UO_2056 (O_2056,N_19883,N_19938);
xnor UO_2057 (O_2057,N_19932,N_19934);
nand UO_2058 (O_2058,N_19819,N_19852);
nor UO_2059 (O_2059,N_19946,N_19865);
and UO_2060 (O_2060,N_19995,N_19848);
nor UO_2061 (O_2061,N_19873,N_19951);
nor UO_2062 (O_2062,N_19866,N_19950);
nand UO_2063 (O_2063,N_19851,N_19914);
or UO_2064 (O_2064,N_19801,N_19997);
or UO_2065 (O_2065,N_19888,N_19970);
or UO_2066 (O_2066,N_19878,N_19914);
xor UO_2067 (O_2067,N_19921,N_19894);
nor UO_2068 (O_2068,N_19800,N_19876);
nand UO_2069 (O_2069,N_19935,N_19932);
nand UO_2070 (O_2070,N_19960,N_19882);
and UO_2071 (O_2071,N_19852,N_19896);
and UO_2072 (O_2072,N_19937,N_19864);
xnor UO_2073 (O_2073,N_19845,N_19893);
or UO_2074 (O_2074,N_19938,N_19922);
and UO_2075 (O_2075,N_19873,N_19971);
nand UO_2076 (O_2076,N_19975,N_19842);
or UO_2077 (O_2077,N_19896,N_19970);
or UO_2078 (O_2078,N_19921,N_19980);
nor UO_2079 (O_2079,N_19994,N_19993);
xor UO_2080 (O_2080,N_19806,N_19890);
nor UO_2081 (O_2081,N_19857,N_19926);
nand UO_2082 (O_2082,N_19840,N_19829);
xor UO_2083 (O_2083,N_19885,N_19857);
or UO_2084 (O_2084,N_19964,N_19802);
and UO_2085 (O_2085,N_19958,N_19974);
xor UO_2086 (O_2086,N_19851,N_19859);
xnor UO_2087 (O_2087,N_19939,N_19956);
or UO_2088 (O_2088,N_19981,N_19983);
or UO_2089 (O_2089,N_19931,N_19850);
nor UO_2090 (O_2090,N_19804,N_19992);
or UO_2091 (O_2091,N_19840,N_19862);
or UO_2092 (O_2092,N_19926,N_19968);
and UO_2093 (O_2093,N_19951,N_19833);
or UO_2094 (O_2094,N_19804,N_19962);
or UO_2095 (O_2095,N_19870,N_19877);
and UO_2096 (O_2096,N_19940,N_19942);
or UO_2097 (O_2097,N_19855,N_19805);
nor UO_2098 (O_2098,N_19836,N_19932);
nor UO_2099 (O_2099,N_19877,N_19872);
nor UO_2100 (O_2100,N_19917,N_19894);
xnor UO_2101 (O_2101,N_19962,N_19862);
nor UO_2102 (O_2102,N_19870,N_19835);
and UO_2103 (O_2103,N_19876,N_19971);
nor UO_2104 (O_2104,N_19982,N_19864);
nand UO_2105 (O_2105,N_19929,N_19917);
nand UO_2106 (O_2106,N_19942,N_19803);
and UO_2107 (O_2107,N_19908,N_19998);
nor UO_2108 (O_2108,N_19903,N_19875);
or UO_2109 (O_2109,N_19841,N_19906);
and UO_2110 (O_2110,N_19993,N_19973);
nor UO_2111 (O_2111,N_19819,N_19879);
xnor UO_2112 (O_2112,N_19944,N_19955);
xnor UO_2113 (O_2113,N_19841,N_19907);
nand UO_2114 (O_2114,N_19882,N_19810);
and UO_2115 (O_2115,N_19978,N_19876);
xnor UO_2116 (O_2116,N_19907,N_19971);
nand UO_2117 (O_2117,N_19992,N_19889);
and UO_2118 (O_2118,N_19990,N_19974);
nor UO_2119 (O_2119,N_19946,N_19899);
nor UO_2120 (O_2120,N_19876,N_19986);
nor UO_2121 (O_2121,N_19933,N_19871);
nand UO_2122 (O_2122,N_19958,N_19952);
and UO_2123 (O_2123,N_19885,N_19887);
and UO_2124 (O_2124,N_19901,N_19987);
nand UO_2125 (O_2125,N_19975,N_19822);
or UO_2126 (O_2126,N_19887,N_19880);
nor UO_2127 (O_2127,N_19894,N_19843);
and UO_2128 (O_2128,N_19883,N_19881);
and UO_2129 (O_2129,N_19858,N_19922);
xnor UO_2130 (O_2130,N_19850,N_19817);
and UO_2131 (O_2131,N_19864,N_19855);
and UO_2132 (O_2132,N_19873,N_19816);
nand UO_2133 (O_2133,N_19840,N_19990);
nor UO_2134 (O_2134,N_19938,N_19836);
nand UO_2135 (O_2135,N_19869,N_19929);
or UO_2136 (O_2136,N_19965,N_19844);
and UO_2137 (O_2137,N_19854,N_19926);
nand UO_2138 (O_2138,N_19823,N_19934);
xor UO_2139 (O_2139,N_19955,N_19880);
or UO_2140 (O_2140,N_19997,N_19883);
and UO_2141 (O_2141,N_19977,N_19938);
xor UO_2142 (O_2142,N_19873,N_19999);
or UO_2143 (O_2143,N_19926,N_19951);
and UO_2144 (O_2144,N_19855,N_19863);
xnor UO_2145 (O_2145,N_19810,N_19933);
xor UO_2146 (O_2146,N_19903,N_19956);
and UO_2147 (O_2147,N_19921,N_19803);
xor UO_2148 (O_2148,N_19997,N_19951);
xor UO_2149 (O_2149,N_19853,N_19810);
and UO_2150 (O_2150,N_19970,N_19998);
xor UO_2151 (O_2151,N_19999,N_19838);
nand UO_2152 (O_2152,N_19847,N_19875);
or UO_2153 (O_2153,N_19892,N_19913);
nand UO_2154 (O_2154,N_19854,N_19930);
and UO_2155 (O_2155,N_19846,N_19849);
or UO_2156 (O_2156,N_19900,N_19910);
nand UO_2157 (O_2157,N_19982,N_19953);
or UO_2158 (O_2158,N_19821,N_19966);
nand UO_2159 (O_2159,N_19815,N_19953);
nor UO_2160 (O_2160,N_19830,N_19852);
or UO_2161 (O_2161,N_19858,N_19977);
xnor UO_2162 (O_2162,N_19865,N_19825);
nor UO_2163 (O_2163,N_19928,N_19940);
and UO_2164 (O_2164,N_19832,N_19914);
and UO_2165 (O_2165,N_19803,N_19899);
nand UO_2166 (O_2166,N_19826,N_19891);
xnor UO_2167 (O_2167,N_19991,N_19937);
nor UO_2168 (O_2168,N_19912,N_19988);
and UO_2169 (O_2169,N_19944,N_19860);
or UO_2170 (O_2170,N_19895,N_19859);
nor UO_2171 (O_2171,N_19916,N_19947);
or UO_2172 (O_2172,N_19835,N_19887);
xor UO_2173 (O_2173,N_19925,N_19940);
nand UO_2174 (O_2174,N_19867,N_19930);
nor UO_2175 (O_2175,N_19862,N_19847);
or UO_2176 (O_2176,N_19805,N_19989);
nand UO_2177 (O_2177,N_19899,N_19878);
or UO_2178 (O_2178,N_19927,N_19925);
xnor UO_2179 (O_2179,N_19913,N_19944);
nand UO_2180 (O_2180,N_19833,N_19881);
nand UO_2181 (O_2181,N_19923,N_19929);
nand UO_2182 (O_2182,N_19918,N_19833);
xnor UO_2183 (O_2183,N_19935,N_19864);
nand UO_2184 (O_2184,N_19900,N_19885);
xnor UO_2185 (O_2185,N_19926,N_19829);
or UO_2186 (O_2186,N_19906,N_19987);
xnor UO_2187 (O_2187,N_19848,N_19964);
nand UO_2188 (O_2188,N_19957,N_19911);
nor UO_2189 (O_2189,N_19824,N_19800);
and UO_2190 (O_2190,N_19869,N_19971);
and UO_2191 (O_2191,N_19806,N_19979);
xor UO_2192 (O_2192,N_19848,N_19910);
xor UO_2193 (O_2193,N_19943,N_19912);
nand UO_2194 (O_2194,N_19901,N_19835);
xnor UO_2195 (O_2195,N_19947,N_19882);
nand UO_2196 (O_2196,N_19964,N_19871);
nand UO_2197 (O_2197,N_19921,N_19843);
and UO_2198 (O_2198,N_19914,N_19975);
xor UO_2199 (O_2199,N_19989,N_19816);
and UO_2200 (O_2200,N_19960,N_19800);
and UO_2201 (O_2201,N_19994,N_19877);
nand UO_2202 (O_2202,N_19958,N_19870);
nand UO_2203 (O_2203,N_19954,N_19991);
nand UO_2204 (O_2204,N_19974,N_19825);
nor UO_2205 (O_2205,N_19917,N_19998);
or UO_2206 (O_2206,N_19906,N_19826);
and UO_2207 (O_2207,N_19899,N_19893);
nand UO_2208 (O_2208,N_19807,N_19942);
nand UO_2209 (O_2209,N_19874,N_19906);
nor UO_2210 (O_2210,N_19829,N_19875);
nor UO_2211 (O_2211,N_19995,N_19950);
nand UO_2212 (O_2212,N_19879,N_19880);
or UO_2213 (O_2213,N_19912,N_19957);
nor UO_2214 (O_2214,N_19969,N_19842);
or UO_2215 (O_2215,N_19800,N_19841);
xnor UO_2216 (O_2216,N_19854,N_19996);
and UO_2217 (O_2217,N_19988,N_19919);
xnor UO_2218 (O_2218,N_19877,N_19860);
or UO_2219 (O_2219,N_19920,N_19865);
and UO_2220 (O_2220,N_19822,N_19978);
xor UO_2221 (O_2221,N_19986,N_19866);
xnor UO_2222 (O_2222,N_19970,N_19921);
or UO_2223 (O_2223,N_19825,N_19854);
xnor UO_2224 (O_2224,N_19850,N_19976);
or UO_2225 (O_2225,N_19818,N_19982);
nor UO_2226 (O_2226,N_19885,N_19865);
xor UO_2227 (O_2227,N_19957,N_19974);
nor UO_2228 (O_2228,N_19991,N_19904);
xor UO_2229 (O_2229,N_19926,N_19800);
nor UO_2230 (O_2230,N_19895,N_19813);
and UO_2231 (O_2231,N_19990,N_19852);
xnor UO_2232 (O_2232,N_19803,N_19844);
nor UO_2233 (O_2233,N_19850,N_19912);
and UO_2234 (O_2234,N_19827,N_19907);
or UO_2235 (O_2235,N_19990,N_19845);
xor UO_2236 (O_2236,N_19847,N_19942);
and UO_2237 (O_2237,N_19859,N_19825);
nand UO_2238 (O_2238,N_19943,N_19901);
nor UO_2239 (O_2239,N_19900,N_19860);
nor UO_2240 (O_2240,N_19887,N_19852);
nand UO_2241 (O_2241,N_19872,N_19919);
and UO_2242 (O_2242,N_19996,N_19989);
or UO_2243 (O_2243,N_19999,N_19915);
xnor UO_2244 (O_2244,N_19961,N_19834);
xnor UO_2245 (O_2245,N_19847,N_19827);
and UO_2246 (O_2246,N_19888,N_19951);
nand UO_2247 (O_2247,N_19826,N_19801);
nand UO_2248 (O_2248,N_19963,N_19907);
xor UO_2249 (O_2249,N_19917,N_19844);
xnor UO_2250 (O_2250,N_19922,N_19884);
and UO_2251 (O_2251,N_19850,N_19990);
xor UO_2252 (O_2252,N_19872,N_19826);
xnor UO_2253 (O_2253,N_19938,N_19860);
xor UO_2254 (O_2254,N_19926,N_19909);
nand UO_2255 (O_2255,N_19895,N_19952);
and UO_2256 (O_2256,N_19950,N_19997);
nand UO_2257 (O_2257,N_19919,N_19897);
and UO_2258 (O_2258,N_19990,N_19813);
or UO_2259 (O_2259,N_19855,N_19847);
xor UO_2260 (O_2260,N_19927,N_19806);
and UO_2261 (O_2261,N_19900,N_19962);
xor UO_2262 (O_2262,N_19934,N_19809);
nor UO_2263 (O_2263,N_19966,N_19871);
xnor UO_2264 (O_2264,N_19996,N_19965);
or UO_2265 (O_2265,N_19936,N_19872);
and UO_2266 (O_2266,N_19960,N_19845);
xnor UO_2267 (O_2267,N_19953,N_19859);
or UO_2268 (O_2268,N_19913,N_19824);
and UO_2269 (O_2269,N_19855,N_19929);
nor UO_2270 (O_2270,N_19946,N_19976);
and UO_2271 (O_2271,N_19897,N_19835);
nand UO_2272 (O_2272,N_19996,N_19962);
nor UO_2273 (O_2273,N_19927,N_19853);
or UO_2274 (O_2274,N_19899,N_19912);
or UO_2275 (O_2275,N_19979,N_19845);
or UO_2276 (O_2276,N_19821,N_19896);
and UO_2277 (O_2277,N_19963,N_19855);
nand UO_2278 (O_2278,N_19993,N_19811);
xor UO_2279 (O_2279,N_19830,N_19865);
or UO_2280 (O_2280,N_19936,N_19868);
xnor UO_2281 (O_2281,N_19966,N_19959);
xnor UO_2282 (O_2282,N_19880,N_19935);
or UO_2283 (O_2283,N_19876,N_19952);
and UO_2284 (O_2284,N_19990,N_19926);
xor UO_2285 (O_2285,N_19956,N_19967);
xnor UO_2286 (O_2286,N_19980,N_19840);
nand UO_2287 (O_2287,N_19918,N_19871);
or UO_2288 (O_2288,N_19906,N_19848);
or UO_2289 (O_2289,N_19869,N_19936);
or UO_2290 (O_2290,N_19957,N_19989);
and UO_2291 (O_2291,N_19881,N_19982);
xor UO_2292 (O_2292,N_19949,N_19857);
nor UO_2293 (O_2293,N_19868,N_19964);
xor UO_2294 (O_2294,N_19828,N_19826);
xor UO_2295 (O_2295,N_19905,N_19808);
and UO_2296 (O_2296,N_19819,N_19820);
nand UO_2297 (O_2297,N_19864,N_19887);
xor UO_2298 (O_2298,N_19885,N_19810);
nor UO_2299 (O_2299,N_19825,N_19894);
nand UO_2300 (O_2300,N_19898,N_19997);
or UO_2301 (O_2301,N_19980,N_19999);
and UO_2302 (O_2302,N_19863,N_19950);
xor UO_2303 (O_2303,N_19988,N_19976);
nor UO_2304 (O_2304,N_19988,N_19841);
nand UO_2305 (O_2305,N_19807,N_19956);
xor UO_2306 (O_2306,N_19963,N_19955);
and UO_2307 (O_2307,N_19879,N_19944);
and UO_2308 (O_2308,N_19991,N_19907);
and UO_2309 (O_2309,N_19942,N_19998);
and UO_2310 (O_2310,N_19832,N_19823);
or UO_2311 (O_2311,N_19924,N_19876);
nand UO_2312 (O_2312,N_19977,N_19909);
and UO_2313 (O_2313,N_19823,N_19936);
and UO_2314 (O_2314,N_19973,N_19832);
nand UO_2315 (O_2315,N_19926,N_19896);
nand UO_2316 (O_2316,N_19878,N_19815);
and UO_2317 (O_2317,N_19937,N_19934);
nor UO_2318 (O_2318,N_19859,N_19850);
nor UO_2319 (O_2319,N_19839,N_19988);
nor UO_2320 (O_2320,N_19953,N_19917);
xnor UO_2321 (O_2321,N_19847,N_19921);
nor UO_2322 (O_2322,N_19830,N_19802);
or UO_2323 (O_2323,N_19821,N_19984);
or UO_2324 (O_2324,N_19940,N_19872);
and UO_2325 (O_2325,N_19931,N_19892);
and UO_2326 (O_2326,N_19814,N_19950);
nor UO_2327 (O_2327,N_19977,N_19831);
nand UO_2328 (O_2328,N_19875,N_19967);
nor UO_2329 (O_2329,N_19807,N_19825);
nand UO_2330 (O_2330,N_19872,N_19937);
nand UO_2331 (O_2331,N_19831,N_19987);
xnor UO_2332 (O_2332,N_19895,N_19854);
xor UO_2333 (O_2333,N_19967,N_19914);
nand UO_2334 (O_2334,N_19995,N_19859);
or UO_2335 (O_2335,N_19899,N_19935);
xor UO_2336 (O_2336,N_19939,N_19853);
and UO_2337 (O_2337,N_19814,N_19968);
or UO_2338 (O_2338,N_19847,N_19948);
nor UO_2339 (O_2339,N_19915,N_19844);
and UO_2340 (O_2340,N_19886,N_19952);
and UO_2341 (O_2341,N_19804,N_19963);
nand UO_2342 (O_2342,N_19962,N_19849);
nand UO_2343 (O_2343,N_19997,N_19822);
nand UO_2344 (O_2344,N_19908,N_19979);
xnor UO_2345 (O_2345,N_19909,N_19879);
or UO_2346 (O_2346,N_19979,N_19865);
and UO_2347 (O_2347,N_19963,N_19949);
or UO_2348 (O_2348,N_19815,N_19869);
nor UO_2349 (O_2349,N_19926,N_19985);
xor UO_2350 (O_2350,N_19957,N_19955);
or UO_2351 (O_2351,N_19990,N_19982);
nor UO_2352 (O_2352,N_19968,N_19821);
nand UO_2353 (O_2353,N_19965,N_19947);
xor UO_2354 (O_2354,N_19943,N_19966);
xnor UO_2355 (O_2355,N_19966,N_19845);
xor UO_2356 (O_2356,N_19921,N_19855);
xor UO_2357 (O_2357,N_19947,N_19929);
or UO_2358 (O_2358,N_19864,N_19927);
nor UO_2359 (O_2359,N_19929,N_19978);
nand UO_2360 (O_2360,N_19991,N_19977);
or UO_2361 (O_2361,N_19819,N_19836);
or UO_2362 (O_2362,N_19950,N_19909);
nand UO_2363 (O_2363,N_19981,N_19949);
xnor UO_2364 (O_2364,N_19942,N_19868);
nor UO_2365 (O_2365,N_19825,N_19896);
nor UO_2366 (O_2366,N_19932,N_19926);
nand UO_2367 (O_2367,N_19977,N_19933);
nor UO_2368 (O_2368,N_19868,N_19826);
or UO_2369 (O_2369,N_19840,N_19846);
nand UO_2370 (O_2370,N_19840,N_19981);
nand UO_2371 (O_2371,N_19926,N_19838);
xnor UO_2372 (O_2372,N_19848,N_19938);
and UO_2373 (O_2373,N_19816,N_19864);
and UO_2374 (O_2374,N_19853,N_19801);
nand UO_2375 (O_2375,N_19880,N_19945);
and UO_2376 (O_2376,N_19978,N_19966);
nand UO_2377 (O_2377,N_19802,N_19826);
nand UO_2378 (O_2378,N_19928,N_19930);
nor UO_2379 (O_2379,N_19909,N_19897);
nor UO_2380 (O_2380,N_19881,N_19820);
nand UO_2381 (O_2381,N_19878,N_19979);
nor UO_2382 (O_2382,N_19859,N_19830);
or UO_2383 (O_2383,N_19847,N_19899);
nor UO_2384 (O_2384,N_19988,N_19867);
nand UO_2385 (O_2385,N_19868,N_19932);
or UO_2386 (O_2386,N_19824,N_19994);
and UO_2387 (O_2387,N_19810,N_19877);
nor UO_2388 (O_2388,N_19909,N_19947);
xor UO_2389 (O_2389,N_19935,N_19876);
nor UO_2390 (O_2390,N_19879,N_19803);
nor UO_2391 (O_2391,N_19894,N_19942);
or UO_2392 (O_2392,N_19923,N_19906);
or UO_2393 (O_2393,N_19836,N_19885);
nand UO_2394 (O_2394,N_19854,N_19967);
nand UO_2395 (O_2395,N_19846,N_19834);
nand UO_2396 (O_2396,N_19911,N_19838);
nor UO_2397 (O_2397,N_19940,N_19889);
nor UO_2398 (O_2398,N_19804,N_19827);
or UO_2399 (O_2399,N_19882,N_19868);
nand UO_2400 (O_2400,N_19895,N_19924);
xor UO_2401 (O_2401,N_19852,N_19921);
nand UO_2402 (O_2402,N_19987,N_19891);
xnor UO_2403 (O_2403,N_19810,N_19829);
nor UO_2404 (O_2404,N_19888,N_19918);
nor UO_2405 (O_2405,N_19864,N_19888);
nand UO_2406 (O_2406,N_19970,N_19822);
xnor UO_2407 (O_2407,N_19938,N_19965);
nor UO_2408 (O_2408,N_19953,N_19900);
and UO_2409 (O_2409,N_19854,N_19980);
nor UO_2410 (O_2410,N_19925,N_19936);
xnor UO_2411 (O_2411,N_19961,N_19955);
and UO_2412 (O_2412,N_19917,N_19882);
xor UO_2413 (O_2413,N_19810,N_19870);
and UO_2414 (O_2414,N_19891,N_19997);
xor UO_2415 (O_2415,N_19966,N_19851);
nor UO_2416 (O_2416,N_19833,N_19937);
nand UO_2417 (O_2417,N_19857,N_19892);
and UO_2418 (O_2418,N_19876,N_19812);
and UO_2419 (O_2419,N_19977,N_19996);
and UO_2420 (O_2420,N_19929,N_19976);
or UO_2421 (O_2421,N_19935,N_19834);
nand UO_2422 (O_2422,N_19840,N_19932);
xnor UO_2423 (O_2423,N_19868,N_19837);
nor UO_2424 (O_2424,N_19871,N_19917);
or UO_2425 (O_2425,N_19865,N_19925);
nor UO_2426 (O_2426,N_19832,N_19964);
xor UO_2427 (O_2427,N_19912,N_19966);
and UO_2428 (O_2428,N_19896,N_19967);
and UO_2429 (O_2429,N_19895,N_19890);
and UO_2430 (O_2430,N_19936,N_19943);
nand UO_2431 (O_2431,N_19962,N_19816);
or UO_2432 (O_2432,N_19876,N_19811);
nor UO_2433 (O_2433,N_19993,N_19804);
nand UO_2434 (O_2434,N_19869,N_19922);
and UO_2435 (O_2435,N_19976,N_19865);
nor UO_2436 (O_2436,N_19843,N_19928);
xor UO_2437 (O_2437,N_19879,N_19912);
xnor UO_2438 (O_2438,N_19840,N_19974);
nand UO_2439 (O_2439,N_19860,N_19948);
xor UO_2440 (O_2440,N_19871,N_19927);
and UO_2441 (O_2441,N_19996,N_19909);
and UO_2442 (O_2442,N_19849,N_19871);
and UO_2443 (O_2443,N_19995,N_19992);
nand UO_2444 (O_2444,N_19909,N_19842);
or UO_2445 (O_2445,N_19848,N_19866);
and UO_2446 (O_2446,N_19880,N_19871);
and UO_2447 (O_2447,N_19813,N_19834);
and UO_2448 (O_2448,N_19872,N_19930);
nor UO_2449 (O_2449,N_19969,N_19851);
nand UO_2450 (O_2450,N_19961,N_19931);
and UO_2451 (O_2451,N_19912,N_19876);
nor UO_2452 (O_2452,N_19840,N_19816);
xor UO_2453 (O_2453,N_19949,N_19878);
and UO_2454 (O_2454,N_19903,N_19823);
nor UO_2455 (O_2455,N_19851,N_19972);
nor UO_2456 (O_2456,N_19897,N_19834);
xnor UO_2457 (O_2457,N_19877,N_19887);
or UO_2458 (O_2458,N_19873,N_19822);
nor UO_2459 (O_2459,N_19985,N_19869);
nor UO_2460 (O_2460,N_19847,N_19846);
and UO_2461 (O_2461,N_19867,N_19965);
nand UO_2462 (O_2462,N_19818,N_19852);
xor UO_2463 (O_2463,N_19831,N_19879);
nor UO_2464 (O_2464,N_19988,N_19901);
xnor UO_2465 (O_2465,N_19863,N_19955);
xor UO_2466 (O_2466,N_19971,N_19892);
xor UO_2467 (O_2467,N_19891,N_19963);
xnor UO_2468 (O_2468,N_19904,N_19986);
nand UO_2469 (O_2469,N_19817,N_19910);
and UO_2470 (O_2470,N_19987,N_19993);
nand UO_2471 (O_2471,N_19819,N_19947);
and UO_2472 (O_2472,N_19988,N_19884);
and UO_2473 (O_2473,N_19908,N_19896);
and UO_2474 (O_2474,N_19826,N_19979);
and UO_2475 (O_2475,N_19827,N_19977);
or UO_2476 (O_2476,N_19917,N_19936);
or UO_2477 (O_2477,N_19892,N_19844);
xnor UO_2478 (O_2478,N_19857,N_19904);
xnor UO_2479 (O_2479,N_19966,N_19886);
and UO_2480 (O_2480,N_19889,N_19924);
nor UO_2481 (O_2481,N_19878,N_19935);
or UO_2482 (O_2482,N_19817,N_19840);
nand UO_2483 (O_2483,N_19848,N_19981);
xor UO_2484 (O_2484,N_19962,N_19992);
and UO_2485 (O_2485,N_19993,N_19980);
or UO_2486 (O_2486,N_19835,N_19905);
or UO_2487 (O_2487,N_19838,N_19987);
and UO_2488 (O_2488,N_19857,N_19815);
xnor UO_2489 (O_2489,N_19916,N_19919);
and UO_2490 (O_2490,N_19890,N_19949);
and UO_2491 (O_2491,N_19850,N_19918);
nor UO_2492 (O_2492,N_19800,N_19903);
xnor UO_2493 (O_2493,N_19801,N_19989);
nor UO_2494 (O_2494,N_19923,N_19804);
and UO_2495 (O_2495,N_19915,N_19857);
or UO_2496 (O_2496,N_19888,N_19964);
and UO_2497 (O_2497,N_19875,N_19897);
xor UO_2498 (O_2498,N_19973,N_19845);
xnor UO_2499 (O_2499,N_19847,N_19842);
endmodule