module basic_750_5000_1000_25_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xor U0 (N_0,In_571,In_121);
xor U1 (N_1,In_404,In_274);
and U2 (N_2,In_272,In_537);
xnor U3 (N_3,In_97,In_314);
and U4 (N_4,In_6,In_592);
or U5 (N_5,In_625,In_99);
nand U6 (N_6,In_207,In_224);
and U7 (N_7,In_688,In_645);
nand U8 (N_8,In_8,In_171);
nor U9 (N_9,In_353,In_640);
xnor U10 (N_10,In_409,In_647);
nor U11 (N_11,In_101,In_489);
nand U12 (N_12,In_576,In_7);
nand U13 (N_13,In_710,In_604);
nor U14 (N_14,In_355,In_259);
or U15 (N_15,In_295,In_23);
nand U16 (N_16,In_313,In_133);
nand U17 (N_17,In_87,In_330);
xor U18 (N_18,In_550,In_75);
nand U19 (N_19,In_651,In_648);
and U20 (N_20,In_174,In_247);
nor U21 (N_21,In_299,In_316);
nor U22 (N_22,In_568,In_368);
and U23 (N_23,In_459,In_211);
nor U24 (N_24,In_672,In_40);
nor U25 (N_25,In_292,In_414);
and U26 (N_26,In_466,In_472);
xor U27 (N_27,In_311,In_159);
nand U28 (N_28,In_193,In_469);
xnor U29 (N_29,In_579,In_72);
and U30 (N_30,In_38,In_398);
nor U31 (N_31,In_257,In_666);
nor U32 (N_32,In_690,In_115);
xnor U33 (N_33,In_59,In_30);
and U34 (N_34,In_83,In_183);
nor U35 (N_35,In_417,In_57);
and U36 (N_36,In_531,In_153);
nor U37 (N_37,In_574,In_51);
nand U38 (N_38,In_650,In_399);
or U39 (N_39,In_315,In_561);
xnor U40 (N_40,In_407,In_79);
or U41 (N_41,In_745,In_552);
nand U42 (N_42,In_608,In_77);
xnor U43 (N_43,In_149,In_678);
nor U44 (N_44,In_29,In_103);
and U45 (N_45,In_162,In_278);
and U46 (N_46,In_463,In_366);
nand U47 (N_47,In_662,In_435);
xor U48 (N_48,In_208,In_518);
xor U49 (N_49,In_492,In_364);
nand U50 (N_50,In_328,In_416);
and U51 (N_51,In_529,In_725);
nand U52 (N_52,In_200,In_467);
xor U53 (N_53,In_124,In_433);
nand U54 (N_54,In_670,In_406);
and U55 (N_55,In_660,In_252);
nand U56 (N_56,In_178,In_334);
nand U57 (N_57,In_700,In_239);
or U58 (N_58,In_285,In_607);
nand U59 (N_59,In_521,In_391);
and U60 (N_60,In_719,In_545);
xor U61 (N_61,In_743,In_535);
nor U62 (N_62,In_323,In_383);
nand U63 (N_63,In_369,In_542);
and U64 (N_64,In_481,In_464);
xor U65 (N_65,In_623,In_122);
nor U66 (N_66,In_677,In_73);
xor U67 (N_67,In_715,In_611);
or U68 (N_68,In_210,In_628);
or U69 (N_69,In_515,In_215);
nor U70 (N_70,In_260,In_653);
nand U71 (N_71,In_388,In_28);
and U72 (N_72,In_746,In_89);
xor U73 (N_73,In_284,In_184);
nand U74 (N_74,In_289,In_452);
or U75 (N_75,In_712,In_303);
nor U76 (N_76,In_168,In_254);
nand U77 (N_77,In_534,In_696);
or U78 (N_78,In_199,In_723);
xor U79 (N_79,In_620,In_67);
nor U80 (N_80,In_27,In_468);
or U81 (N_81,In_375,In_4);
and U82 (N_82,In_60,In_170);
or U83 (N_83,In_18,In_10);
xnor U84 (N_84,In_641,In_716);
xor U85 (N_85,In_395,In_680);
nand U86 (N_86,In_93,In_714);
nor U87 (N_87,In_127,In_350);
xnor U88 (N_88,In_708,In_646);
nand U89 (N_89,In_68,In_737);
xor U90 (N_90,In_504,In_474);
nor U91 (N_91,In_727,In_172);
xor U92 (N_92,In_243,In_455);
xor U93 (N_93,In_594,In_674);
xnor U94 (N_94,In_340,In_639);
and U95 (N_95,In_359,In_325);
or U96 (N_96,In_621,In_373);
and U97 (N_97,In_160,In_175);
xnor U98 (N_98,In_108,In_381);
or U99 (N_99,In_687,In_502);
nand U100 (N_100,In_161,In_735);
or U101 (N_101,In_186,In_182);
or U102 (N_102,In_437,In_196);
nand U103 (N_103,In_302,In_638);
nor U104 (N_104,In_42,In_513);
nand U105 (N_105,In_562,In_533);
nand U106 (N_106,In_32,In_412);
or U107 (N_107,In_610,In_74);
nand U108 (N_108,In_496,In_480);
nor U109 (N_109,In_730,In_573);
nand U110 (N_110,In_280,In_589);
nor U111 (N_111,In_382,In_487);
and U112 (N_112,In_556,In_229);
or U113 (N_113,In_304,In_113);
xor U114 (N_114,In_308,In_98);
nand U115 (N_115,In_107,In_403);
and U116 (N_116,In_460,In_490);
nand U117 (N_117,In_692,In_205);
and U118 (N_118,In_82,In_749);
or U119 (N_119,In_636,In_413);
nor U120 (N_120,In_577,In_116);
and U121 (N_121,In_269,In_479);
or U122 (N_122,In_270,In_441);
and U123 (N_123,In_50,In_477);
xor U124 (N_124,In_614,In_606);
nor U125 (N_125,In_34,In_493);
xor U126 (N_126,In_389,In_250);
nor U127 (N_127,In_671,In_519);
nand U128 (N_128,In_164,In_400);
nor U129 (N_129,In_232,In_258);
nand U130 (N_130,In_219,In_106);
and U131 (N_131,In_551,In_432);
nand U132 (N_132,In_351,In_158);
and U133 (N_133,In_682,In_405);
nor U134 (N_134,In_26,In_118);
and U135 (N_135,In_586,In_283);
and U136 (N_136,In_294,In_429);
and U137 (N_137,In_190,In_36);
nor U138 (N_138,In_420,In_94);
xor U139 (N_139,In_661,In_197);
or U140 (N_140,In_377,In_557);
or U141 (N_141,In_447,In_233);
xor U142 (N_142,In_185,In_703);
and U143 (N_143,In_216,In_333);
nand U144 (N_144,In_145,In_191);
or U145 (N_145,In_267,In_155);
xor U146 (N_146,In_522,In_341);
or U147 (N_147,In_483,In_442);
and U148 (N_148,In_20,In_618);
nor U149 (N_149,In_578,In_335);
nand U150 (N_150,In_686,In_736);
and U151 (N_151,In_90,In_33);
nand U152 (N_152,In_498,In_704);
and U153 (N_153,In_506,In_721);
xnor U154 (N_154,In_629,In_613);
or U155 (N_155,In_236,In_540);
or U156 (N_156,In_387,In_129);
and U157 (N_157,In_582,In_624);
or U158 (N_158,In_227,In_600);
nand U159 (N_159,In_201,In_43);
xor U160 (N_160,In_591,In_206);
xor U161 (N_161,In_598,In_450);
or U162 (N_162,In_748,In_202);
or U163 (N_163,In_512,In_142);
nand U164 (N_164,In_223,In_478);
xor U165 (N_165,In_378,In_62);
and U166 (N_166,In_742,In_738);
xnor U167 (N_167,In_689,In_148);
nor U168 (N_168,In_81,In_151);
or U169 (N_169,In_726,In_597);
or U170 (N_170,In_626,In_635);
and U171 (N_171,In_198,In_44);
xnor U172 (N_172,In_279,In_297);
nor U173 (N_173,In_532,In_39);
xor U174 (N_174,In_156,In_695);
and U175 (N_175,In_194,In_110);
nand U176 (N_176,In_656,In_14);
or U177 (N_177,In_318,In_706);
or U178 (N_178,In_265,In_136);
and U179 (N_179,In_235,In_543);
xor U180 (N_180,In_553,In_658);
xnor U181 (N_181,In_343,In_560);
or U182 (N_182,In_443,In_189);
xor U183 (N_183,In_61,In_286);
nor U184 (N_184,In_84,In_218);
or U185 (N_185,In_192,In_601);
xor U186 (N_186,In_271,In_609);
and U187 (N_187,In_525,In_80);
or U188 (N_188,In_634,In_664);
or U189 (N_189,In_428,In_566);
or U190 (N_190,In_209,In_451);
and U191 (N_191,In_546,In_312);
nand U192 (N_192,In_360,In_222);
and U193 (N_193,In_22,In_665);
nand U194 (N_194,In_49,In_587);
nand U195 (N_195,In_177,In_66);
xnor U196 (N_196,In_332,In_602);
nand U197 (N_197,In_427,In_123);
or U198 (N_198,In_140,In_394);
nor U199 (N_199,In_713,In_71);
xor U200 (N_200,N_35,In_390);
and U201 (N_201,In_273,In_415);
nand U202 (N_202,N_7,In_337);
and U203 (N_203,N_172,In_449);
nor U204 (N_204,In_212,N_118);
and U205 (N_205,In_230,N_174);
or U206 (N_206,In_54,In_539);
or U207 (N_207,N_180,N_98);
xnor U208 (N_208,In_627,N_58);
or U209 (N_209,N_97,In_17);
xnor U210 (N_210,In_245,In_347);
xnor U211 (N_211,N_190,In_64);
nand U212 (N_212,In_76,In_471);
nand U213 (N_213,N_166,In_514);
nor U214 (N_214,In_747,In_702);
nor U215 (N_215,In_263,In_261);
nor U216 (N_216,N_159,N_39);
and U217 (N_217,In_583,In_13);
nand U218 (N_218,N_20,N_186);
or U219 (N_219,In_221,In_495);
nor U220 (N_220,In_491,In_130);
xor U221 (N_221,N_95,In_457);
and U222 (N_222,In_691,In_86);
nor U223 (N_223,N_109,In_2);
and U224 (N_224,N_163,In_264);
nand U225 (N_225,N_79,N_158);
nor U226 (N_226,N_47,N_89);
or U227 (N_227,In_281,In_376);
xor U228 (N_228,In_401,N_153);
and U229 (N_229,In_731,In_329);
nand U230 (N_230,In_709,In_154);
nor U231 (N_231,In_338,In_371);
or U232 (N_232,In_152,In_605);
or U233 (N_233,N_162,N_178);
nor U234 (N_234,In_448,N_192);
nor U235 (N_235,In_570,In_507);
nor U236 (N_236,In_585,In_675);
and U237 (N_237,In_317,N_120);
and U238 (N_238,In_249,N_113);
xor U239 (N_239,In_262,In_511);
nor U240 (N_240,In_56,N_161);
or U241 (N_241,N_15,In_203);
and U242 (N_242,N_144,N_188);
and U243 (N_243,In_430,In_616);
or U244 (N_244,In_138,In_440);
nor U245 (N_245,In_47,In_549);
nand U246 (N_246,In_520,In_526);
nor U247 (N_247,In_226,In_425);
nand U248 (N_248,In_436,N_104);
and U249 (N_249,N_30,In_321);
nand U250 (N_250,In_575,N_36);
nor U251 (N_251,In_244,In_593);
or U252 (N_252,In_679,N_173);
xor U253 (N_253,In_422,In_374);
nor U254 (N_254,N_199,In_728);
and U255 (N_255,In_352,In_372);
or U256 (N_256,N_164,In_698);
nor U257 (N_257,In_55,In_473);
and U258 (N_258,In_741,N_94);
xor U259 (N_259,In_176,In_402);
xor U260 (N_260,In_91,In_501);
nand U261 (N_261,In_434,N_156);
nand U262 (N_262,N_177,N_119);
xnor U263 (N_263,N_195,In_188);
or U264 (N_264,N_88,In_676);
or U265 (N_265,N_73,N_14);
nand U266 (N_266,N_17,N_55);
xor U267 (N_267,In_70,N_29);
xnor U268 (N_268,In_125,In_141);
nand U269 (N_269,In_45,N_129);
nand U270 (N_270,N_126,In_5);
nor U271 (N_271,In_275,N_184);
xnor U272 (N_272,N_13,In_309);
nor U273 (N_273,In_657,In_41);
and U274 (N_274,N_171,N_110);
nor U275 (N_275,In_655,In_733);
nand U276 (N_276,N_136,In_348);
and U277 (N_277,N_147,In_165);
and U278 (N_278,N_21,In_724);
or U279 (N_279,N_187,In_65);
or U280 (N_280,In_612,In_524);
nand U281 (N_281,N_107,In_109);
and U282 (N_282,N_42,N_2);
or U283 (N_283,In_718,N_194);
and U284 (N_284,In_580,In_117);
and U285 (N_285,N_93,In_287);
xnor U286 (N_286,In_555,In_362);
or U287 (N_287,In_169,In_370);
nand U288 (N_288,In_240,N_152);
nor U289 (N_289,N_141,N_138);
and U290 (N_290,N_167,In_642);
nor U291 (N_291,N_53,In_411);
or U292 (N_292,In_242,N_92);
and U293 (N_293,In_96,In_357);
xnor U294 (N_294,In_3,In_143);
and U295 (N_295,N_198,N_0);
nand U296 (N_296,In_187,N_31);
nand U297 (N_297,In_517,In_69);
and U298 (N_298,In_541,N_179);
and U299 (N_299,N_101,N_61);
nand U300 (N_300,N_66,In_644);
or U301 (N_301,In_392,N_19);
xor U302 (N_302,N_165,In_462);
xor U303 (N_303,N_40,In_538);
nor U304 (N_304,N_140,N_1);
or U305 (N_305,N_197,In_126);
or U306 (N_306,In_363,In_681);
nor U307 (N_307,N_123,In_131);
and U308 (N_308,In_722,In_418);
and U309 (N_309,In_166,In_484);
and U310 (N_310,N_18,N_6);
xnor U311 (N_311,N_157,In_509);
or U312 (N_312,In_46,In_697);
or U313 (N_313,In_547,In_669);
nor U314 (N_314,In_684,In_488);
or U315 (N_315,N_127,N_38);
nor U316 (N_316,In_445,N_25);
nand U317 (N_317,N_43,In_423);
nand U318 (N_318,In_85,In_421);
and U319 (N_319,In_617,N_5);
or U320 (N_320,In_16,In_282);
nor U321 (N_321,N_82,N_134);
nor U322 (N_322,In_503,N_23);
and U323 (N_323,In_63,In_288);
nand U324 (N_324,In_290,In_354);
and U325 (N_325,In_386,N_191);
or U326 (N_326,N_90,In_426);
and U327 (N_327,In_58,In_581);
and U328 (N_328,In_564,In_25);
nor U329 (N_329,In_24,N_28);
xnor U330 (N_330,N_34,N_106);
nor U331 (N_331,N_57,In_1);
nand U332 (N_332,N_128,In_384);
or U333 (N_333,In_204,In_11);
nand U334 (N_334,N_76,In_572);
nand U335 (N_335,In_12,In_147);
and U336 (N_336,N_63,In_307);
and U337 (N_337,N_83,N_105);
and U338 (N_338,In_508,N_114);
nor U339 (N_339,N_41,In_365);
nor U340 (N_340,N_149,In_19);
nand U341 (N_341,N_50,N_11);
nand U342 (N_342,In_319,In_228);
xnor U343 (N_343,In_663,In_567);
xnor U344 (N_344,In_652,N_148);
nor U345 (N_345,In_300,N_8);
or U346 (N_346,N_112,In_461);
nor U347 (N_347,In_132,In_163);
and U348 (N_348,N_3,In_699);
nand U349 (N_349,In_707,In_277);
xnor U350 (N_350,In_37,N_87);
or U351 (N_351,In_558,In_266);
nor U352 (N_352,N_130,N_146);
nand U353 (N_353,N_108,N_48);
xnor U354 (N_354,In_569,In_523);
nor U355 (N_355,In_444,In_327);
or U356 (N_356,In_633,N_56);
and U357 (N_357,N_60,In_120);
xor U358 (N_358,In_114,In_234);
xnor U359 (N_359,In_298,In_320);
nor U360 (N_360,In_322,N_67);
nor U361 (N_361,In_146,In_554);
nor U362 (N_362,In_424,In_213);
or U363 (N_363,In_637,In_454);
xnor U364 (N_364,In_499,N_99);
nor U365 (N_365,In_324,N_24);
and U366 (N_366,In_528,In_536);
or U367 (N_367,N_52,N_181);
xor U368 (N_368,N_12,In_482);
nand U369 (N_369,In_476,In_310);
or U370 (N_370,In_214,In_134);
nand U371 (N_371,N_68,In_379);
nor U372 (N_372,In_599,N_49);
or U373 (N_373,N_71,N_132);
or U374 (N_374,N_117,In_485);
nor U375 (N_375,In_565,In_15);
nand U376 (N_376,In_631,In_0);
nand U377 (N_377,In_102,In_361);
nand U378 (N_378,In_701,In_128);
and U379 (N_379,N_81,N_135);
or U380 (N_380,In_431,In_397);
nand U381 (N_381,In_668,In_144);
nand U382 (N_382,In_268,N_26);
nor U383 (N_383,In_596,In_622);
nand U384 (N_384,N_182,In_683);
and U385 (N_385,N_70,In_276);
or U386 (N_386,N_46,In_475);
nand U387 (N_387,N_189,N_77);
nand U388 (N_388,In_225,In_35);
nand U389 (N_389,In_251,In_88);
or U390 (N_390,N_151,In_135);
nor U391 (N_391,N_193,In_667);
xnor U392 (N_392,In_603,N_80);
and U393 (N_393,In_632,In_659);
nand U394 (N_394,In_385,In_438);
nand U395 (N_395,N_154,In_21);
nor U396 (N_396,In_705,In_588);
and U397 (N_397,In_173,N_84);
xnor U398 (N_398,In_104,In_356);
nand U399 (N_399,N_155,In_179);
nand U400 (N_400,In_527,N_100);
and U401 (N_401,N_319,N_311);
nor U402 (N_402,N_247,In_367);
and U403 (N_403,N_228,In_544);
nand U404 (N_404,N_354,N_203);
and U405 (N_405,N_332,N_250);
nand U406 (N_406,N_216,N_237);
or U407 (N_407,N_321,In_326);
nor U408 (N_408,N_348,In_220);
or U409 (N_409,N_196,N_150);
nand U410 (N_410,N_304,N_208);
nand U411 (N_411,In_630,N_238);
nor U412 (N_412,N_252,In_720);
or U413 (N_413,In_729,N_373);
or U414 (N_414,In_139,N_330);
nor U415 (N_415,N_242,In_711);
and U416 (N_416,N_255,In_342);
xnor U417 (N_417,In_654,N_78);
nor U418 (N_418,In_410,N_139);
xor U419 (N_419,In_439,N_277);
nor U420 (N_420,N_241,In_739);
nand U421 (N_421,N_270,N_392);
or U422 (N_422,In_446,N_398);
nand U423 (N_423,In_643,N_303);
and U424 (N_424,N_266,In_548);
or U425 (N_425,N_305,In_181);
and U426 (N_426,N_33,N_337);
xnor U427 (N_427,N_335,N_372);
and U428 (N_428,N_291,N_368);
nor U429 (N_429,N_142,N_221);
nor U430 (N_430,N_251,N_176);
or U431 (N_431,N_381,N_296);
or U432 (N_432,N_357,In_119);
nor U433 (N_433,N_394,N_268);
nor U434 (N_434,N_318,N_295);
and U435 (N_435,N_168,In_231);
or U436 (N_436,N_125,N_299);
nand U437 (N_437,N_334,N_386);
and U438 (N_438,N_314,N_286);
nand U439 (N_439,N_280,N_384);
or U440 (N_440,N_271,N_293);
nand U441 (N_441,N_320,N_387);
or U442 (N_442,N_379,In_217);
nand U443 (N_443,N_333,In_336);
or U444 (N_444,N_22,N_160);
or U445 (N_445,N_103,N_102);
or U446 (N_446,N_133,In_293);
or U447 (N_447,N_262,N_374);
and U448 (N_448,In_345,In_157);
nand U449 (N_449,N_325,N_269);
nand U450 (N_450,N_265,In_419);
and U451 (N_451,In_255,N_301);
xnor U452 (N_452,N_360,In_331);
and U453 (N_453,N_388,In_497);
or U454 (N_454,In_465,In_53);
nand U455 (N_455,N_390,N_353);
nand U456 (N_456,In_380,N_239);
nand U457 (N_457,N_204,In_31);
xor U458 (N_458,N_382,N_326);
xor U459 (N_459,N_16,In_590);
nor U460 (N_460,N_232,N_312);
or U461 (N_461,N_145,In_516);
or U462 (N_462,N_246,In_408);
or U463 (N_463,In_246,N_383);
nand U464 (N_464,N_331,N_10);
nand U465 (N_465,N_340,N_343);
nor U466 (N_466,N_115,N_116);
nor U467 (N_467,N_391,In_559);
and U468 (N_468,In_344,In_393);
and U469 (N_469,N_341,N_276);
and U470 (N_470,N_205,In_619);
nand U471 (N_471,In_744,In_180);
nor U472 (N_472,N_185,N_74);
nand U473 (N_473,In_456,In_693);
nor U474 (N_474,N_356,N_310);
nand U475 (N_475,In_734,N_292);
nor U476 (N_476,N_338,In_563);
nor U477 (N_477,N_207,N_236);
and U478 (N_478,In_649,N_219);
or U479 (N_479,In_238,N_290);
or U480 (N_480,N_389,N_377);
nand U481 (N_481,N_249,In_346);
nand U482 (N_482,In_732,N_288);
nor U483 (N_483,N_69,N_218);
or U484 (N_484,N_283,N_327);
nand U485 (N_485,N_344,N_258);
or U486 (N_486,In_453,N_206);
nand U487 (N_487,In_500,In_150);
xnor U488 (N_488,In_694,N_91);
xor U489 (N_489,N_350,N_297);
nand U490 (N_490,In_112,N_395);
nor U491 (N_491,In_105,In_595);
nand U492 (N_492,In_9,N_300);
and U493 (N_493,In_673,N_231);
and U494 (N_494,In_717,N_349);
xnor U495 (N_495,In_167,N_336);
and U496 (N_496,N_220,N_169);
and U497 (N_497,N_201,N_342);
or U498 (N_498,N_267,N_234);
and U499 (N_499,N_111,In_248);
xor U500 (N_500,N_279,N_346);
nor U501 (N_501,N_351,In_78);
xor U502 (N_502,N_72,N_235);
and U503 (N_503,N_62,In_306);
xor U504 (N_504,In_241,N_322);
xor U505 (N_505,In_494,N_352);
nand U506 (N_506,N_263,N_370);
and U507 (N_507,N_274,N_363);
and U508 (N_508,N_254,In_195);
nand U509 (N_509,N_278,N_75);
xnor U510 (N_510,N_212,N_358);
and U511 (N_511,N_309,N_380);
or U512 (N_512,N_44,N_272);
nand U513 (N_513,N_85,N_323);
nand U514 (N_514,In_111,N_217);
nor U515 (N_515,N_9,N_329);
nand U516 (N_516,N_260,N_65);
nand U517 (N_517,N_256,In_615);
and U518 (N_518,N_170,N_308);
or U519 (N_519,N_361,N_243);
nor U520 (N_520,In_237,N_122);
nand U521 (N_521,In_92,In_305);
xnor U522 (N_522,N_264,N_244);
and U523 (N_523,N_51,N_328);
nand U524 (N_524,N_27,N_366);
or U525 (N_525,N_284,In_253);
or U526 (N_526,N_143,N_306);
or U527 (N_527,N_124,In_740);
nor U528 (N_528,In_358,N_365);
or U529 (N_529,N_285,N_289);
and U530 (N_530,N_226,N_302);
or U531 (N_531,N_183,N_287);
nor U532 (N_532,N_59,N_345);
xnor U533 (N_533,N_227,N_281);
nand U534 (N_534,N_282,N_175);
xor U535 (N_535,In_296,N_248);
and U536 (N_536,N_121,In_95);
nand U537 (N_537,In_685,In_256);
or U538 (N_538,N_298,N_257);
nor U539 (N_539,In_349,N_64);
or U540 (N_540,N_362,N_369);
and U541 (N_541,N_376,N_261);
nor U542 (N_542,N_316,N_131);
nand U543 (N_543,N_202,N_45);
and U544 (N_544,N_215,In_505);
nand U545 (N_545,N_367,N_224);
or U546 (N_546,N_324,In_530);
nor U547 (N_547,N_294,N_211);
and U548 (N_548,N_229,N_225);
nand U549 (N_549,N_54,In_396);
or U550 (N_550,N_214,In_291);
and U551 (N_551,N_359,In_301);
and U552 (N_552,N_86,N_230);
xnor U553 (N_553,N_259,N_223);
and U554 (N_554,N_96,N_378);
nand U555 (N_555,N_273,N_339);
and U556 (N_556,N_313,N_200);
nor U557 (N_557,In_48,In_510);
nor U558 (N_558,N_222,N_37);
xnor U559 (N_559,N_385,In_458);
nor U560 (N_560,N_245,N_397);
nor U561 (N_561,N_253,N_355);
nand U562 (N_562,In_486,N_233);
and U563 (N_563,N_213,In_52);
or U564 (N_564,N_371,In_470);
nor U565 (N_565,N_375,N_307);
nand U566 (N_566,In_584,N_275);
nor U567 (N_567,In_100,N_399);
nand U568 (N_568,N_137,N_209);
nand U569 (N_569,N_210,N_32);
nor U570 (N_570,N_240,In_137);
or U571 (N_571,N_396,N_315);
nand U572 (N_572,N_393,In_339);
nand U573 (N_573,N_347,N_4);
or U574 (N_574,N_317,N_364);
and U575 (N_575,In_654,In_253);
nand U576 (N_576,N_16,N_251);
nand U577 (N_577,N_237,N_103);
and U578 (N_578,N_237,N_245);
nor U579 (N_579,In_595,In_739);
or U580 (N_580,N_150,N_255);
or U581 (N_581,N_185,N_286);
and U582 (N_582,N_169,N_255);
nor U583 (N_583,In_95,N_45);
and U584 (N_584,N_217,In_505);
and U585 (N_585,In_419,In_694);
nand U586 (N_586,In_349,N_196);
or U587 (N_587,In_339,N_355);
nand U588 (N_588,N_325,N_296);
or U589 (N_589,N_168,N_296);
xnor U590 (N_590,N_347,N_316);
nor U591 (N_591,N_388,N_390);
nand U592 (N_592,N_321,N_295);
or U593 (N_593,N_299,In_53);
or U594 (N_594,N_337,N_275);
or U595 (N_595,N_388,N_383);
nand U596 (N_596,N_208,In_255);
xnor U597 (N_597,N_203,N_272);
or U598 (N_598,N_350,In_231);
nand U599 (N_599,In_137,N_226);
nand U600 (N_600,N_542,N_589);
xnor U601 (N_601,N_574,N_406);
nand U602 (N_602,N_492,N_517);
nand U603 (N_603,N_428,N_535);
nand U604 (N_604,N_532,N_412);
and U605 (N_605,N_422,N_426);
or U606 (N_606,N_560,N_482);
nor U607 (N_607,N_416,N_480);
and U608 (N_608,N_464,N_553);
nand U609 (N_609,N_497,N_414);
and U610 (N_610,N_448,N_457);
nor U611 (N_611,N_570,N_483);
xnor U612 (N_612,N_521,N_586);
nand U613 (N_613,N_523,N_544);
xor U614 (N_614,N_546,N_400);
xor U615 (N_615,N_593,N_530);
and U616 (N_616,N_502,N_456);
and U617 (N_617,N_442,N_498);
nor U618 (N_618,N_520,N_467);
nand U619 (N_619,N_518,N_441);
xor U620 (N_620,N_562,N_539);
or U621 (N_621,N_564,N_487);
nor U622 (N_622,N_450,N_488);
or U623 (N_623,N_580,N_431);
nand U624 (N_624,N_433,N_410);
nor U625 (N_625,N_451,N_404);
nand U626 (N_626,N_460,N_411);
or U627 (N_627,N_522,N_413);
or U628 (N_628,N_478,N_587);
and U629 (N_629,N_514,N_573);
and U630 (N_630,N_515,N_435);
nor U631 (N_631,N_545,N_582);
nor U632 (N_632,N_525,N_407);
nor U633 (N_633,N_496,N_561);
xnor U634 (N_634,N_434,N_531);
and U635 (N_635,N_436,N_556);
nand U636 (N_636,N_503,N_405);
and U637 (N_637,N_500,N_432);
or U638 (N_638,N_446,N_519);
xor U639 (N_639,N_491,N_481);
xor U640 (N_640,N_534,N_507);
nor U641 (N_641,N_470,N_566);
nor U642 (N_642,N_490,N_438);
xnor U643 (N_643,N_477,N_588);
xnor U644 (N_644,N_552,N_453);
nor U645 (N_645,N_569,N_445);
and U646 (N_646,N_462,N_415);
xor U647 (N_647,N_575,N_468);
nor U648 (N_648,N_557,N_501);
nor U649 (N_649,N_479,N_455);
nand U650 (N_650,N_548,N_463);
nor U651 (N_651,N_471,N_537);
nor U652 (N_652,N_461,N_430);
nor U653 (N_653,N_590,N_549);
xnor U654 (N_654,N_579,N_576);
or U655 (N_655,N_506,N_536);
and U656 (N_656,N_594,N_452);
nor U657 (N_657,N_499,N_485);
or U658 (N_658,N_505,N_540);
and U659 (N_659,N_538,N_528);
nor U660 (N_660,N_559,N_401);
or U661 (N_661,N_550,N_489);
xnor U662 (N_662,N_444,N_554);
or U663 (N_663,N_565,N_476);
xor U664 (N_664,N_458,N_425);
or U665 (N_665,N_427,N_584);
xor U666 (N_666,N_526,N_578);
or U667 (N_667,N_585,N_598);
xor U668 (N_668,N_403,N_543);
and U669 (N_669,N_474,N_509);
or U670 (N_670,N_583,N_597);
nand U671 (N_671,N_402,N_555);
xnor U672 (N_672,N_475,N_420);
and U673 (N_673,N_591,N_409);
nand U674 (N_674,N_473,N_443);
and U675 (N_675,N_429,N_437);
nor U676 (N_676,N_454,N_533);
or U677 (N_677,N_440,N_558);
and U678 (N_678,N_465,N_596);
nor U679 (N_679,N_504,N_486);
or U680 (N_680,N_469,N_581);
nor U681 (N_681,N_577,N_508);
and U682 (N_682,N_527,N_516);
nand U683 (N_683,N_511,N_595);
xor U684 (N_684,N_408,N_493);
and U685 (N_685,N_417,N_421);
and U686 (N_686,N_571,N_419);
or U687 (N_687,N_568,N_484);
nand U688 (N_688,N_466,N_449);
nand U689 (N_689,N_424,N_472);
or U690 (N_690,N_529,N_459);
nand U691 (N_691,N_572,N_423);
or U692 (N_692,N_447,N_592);
xor U693 (N_693,N_547,N_599);
xor U694 (N_694,N_541,N_567);
nand U695 (N_695,N_495,N_510);
and U696 (N_696,N_513,N_512);
nor U697 (N_697,N_563,N_439);
and U698 (N_698,N_524,N_418);
nand U699 (N_699,N_551,N_494);
xor U700 (N_700,N_561,N_415);
xor U701 (N_701,N_457,N_569);
and U702 (N_702,N_492,N_580);
nand U703 (N_703,N_480,N_452);
xor U704 (N_704,N_534,N_463);
xnor U705 (N_705,N_473,N_591);
and U706 (N_706,N_406,N_581);
nand U707 (N_707,N_484,N_597);
or U708 (N_708,N_480,N_437);
or U709 (N_709,N_447,N_546);
or U710 (N_710,N_531,N_478);
and U711 (N_711,N_565,N_464);
xor U712 (N_712,N_470,N_409);
nor U713 (N_713,N_490,N_439);
xor U714 (N_714,N_597,N_442);
or U715 (N_715,N_538,N_470);
and U716 (N_716,N_466,N_599);
xnor U717 (N_717,N_417,N_436);
nor U718 (N_718,N_552,N_508);
nand U719 (N_719,N_580,N_545);
or U720 (N_720,N_461,N_544);
nand U721 (N_721,N_586,N_427);
or U722 (N_722,N_464,N_568);
and U723 (N_723,N_492,N_432);
or U724 (N_724,N_529,N_460);
and U725 (N_725,N_511,N_598);
xor U726 (N_726,N_508,N_463);
and U727 (N_727,N_459,N_428);
nand U728 (N_728,N_484,N_474);
nor U729 (N_729,N_513,N_486);
nand U730 (N_730,N_409,N_481);
nand U731 (N_731,N_493,N_481);
and U732 (N_732,N_516,N_478);
and U733 (N_733,N_510,N_526);
and U734 (N_734,N_496,N_430);
and U735 (N_735,N_521,N_519);
and U736 (N_736,N_406,N_441);
nand U737 (N_737,N_535,N_435);
and U738 (N_738,N_586,N_488);
or U739 (N_739,N_550,N_574);
and U740 (N_740,N_429,N_539);
nand U741 (N_741,N_542,N_550);
or U742 (N_742,N_439,N_555);
nor U743 (N_743,N_510,N_473);
and U744 (N_744,N_583,N_564);
or U745 (N_745,N_499,N_462);
nand U746 (N_746,N_502,N_473);
nor U747 (N_747,N_559,N_430);
nor U748 (N_748,N_516,N_532);
nor U749 (N_749,N_557,N_515);
or U750 (N_750,N_531,N_442);
xor U751 (N_751,N_432,N_525);
or U752 (N_752,N_414,N_444);
nor U753 (N_753,N_590,N_419);
xor U754 (N_754,N_428,N_487);
nand U755 (N_755,N_573,N_566);
xor U756 (N_756,N_438,N_515);
xnor U757 (N_757,N_467,N_454);
nor U758 (N_758,N_521,N_468);
or U759 (N_759,N_536,N_551);
xnor U760 (N_760,N_535,N_581);
xnor U761 (N_761,N_547,N_591);
xor U762 (N_762,N_449,N_480);
nand U763 (N_763,N_561,N_504);
nand U764 (N_764,N_580,N_504);
and U765 (N_765,N_476,N_418);
or U766 (N_766,N_584,N_519);
or U767 (N_767,N_466,N_409);
nand U768 (N_768,N_550,N_484);
xnor U769 (N_769,N_582,N_566);
or U770 (N_770,N_458,N_566);
xnor U771 (N_771,N_455,N_559);
nand U772 (N_772,N_580,N_488);
or U773 (N_773,N_508,N_512);
nor U774 (N_774,N_508,N_581);
nand U775 (N_775,N_563,N_438);
and U776 (N_776,N_475,N_482);
and U777 (N_777,N_570,N_597);
or U778 (N_778,N_447,N_439);
xnor U779 (N_779,N_467,N_524);
nand U780 (N_780,N_515,N_447);
nand U781 (N_781,N_499,N_580);
and U782 (N_782,N_586,N_596);
and U783 (N_783,N_494,N_417);
or U784 (N_784,N_593,N_504);
and U785 (N_785,N_403,N_445);
nand U786 (N_786,N_464,N_448);
or U787 (N_787,N_465,N_425);
and U788 (N_788,N_415,N_441);
or U789 (N_789,N_575,N_464);
nor U790 (N_790,N_506,N_490);
and U791 (N_791,N_454,N_580);
nand U792 (N_792,N_579,N_470);
nand U793 (N_793,N_563,N_464);
nor U794 (N_794,N_564,N_445);
and U795 (N_795,N_533,N_552);
xor U796 (N_796,N_546,N_415);
or U797 (N_797,N_551,N_528);
nand U798 (N_798,N_429,N_402);
or U799 (N_799,N_410,N_566);
or U800 (N_800,N_764,N_608);
nor U801 (N_801,N_716,N_770);
nor U802 (N_802,N_742,N_769);
nand U803 (N_803,N_664,N_730);
nor U804 (N_804,N_658,N_725);
and U805 (N_805,N_699,N_708);
and U806 (N_806,N_724,N_617);
nand U807 (N_807,N_729,N_672);
or U808 (N_808,N_726,N_743);
xnor U809 (N_809,N_633,N_788);
xnor U810 (N_810,N_652,N_747);
xor U811 (N_811,N_762,N_607);
xor U812 (N_812,N_787,N_686);
nand U813 (N_813,N_645,N_719);
xnor U814 (N_814,N_697,N_755);
xnor U815 (N_815,N_626,N_684);
xnor U816 (N_816,N_701,N_659);
or U817 (N_817,N_622,N_741);
nor U818 (N_818,N_717,N_750);
or U819 (N_819,N_761,N_651);
and U820 (N_820,N_648,N_620);
and U821 (N_821,N_738,N_649);
xnor U822 (N_822,N_694,N_792);
xor U823 (N_823,N_783,N_692);
nand U824 (N_824,N_777,N_793);
or U825 (N_825,N_687,N_759);
or U826 (N_826,N_654,N_707);
xor U827 (N_827,N_675,N_722);
and U828 (N_828,N_682,N_778);
nor U829 (N_829,N_776,N_765);
and U830 (N_830,N_720,N_737);
xnor U831 (N_831,N_732,N_683);
nor U832 (N_832,N_733,N_670);
xnor U833 (N_833,N_657,N_632);
xnor U834 (N_834,N_621,N_727);
or U835 (N_835,N_736,N_754);
and U836 (N_836,N_756,N_735);
xor U837 (N_837,N_774,N_685);
or U838 (N_838,N_693,N_690);
and U839 (N_839,N_642,N_640);
and U840 (N_840,N_680,N_606);
nand U841 (N_841,N_695,N_782);
nor U842 (N_842,N_627,N_638);
nor U843 (N_843,N_799,N_634);
xor U844 (N_844,N_705,N_748);
nor U845 (N_845,N_772,N_602);
nor U846 (N_846,N_603,N_669);
xnor U847 (N_847,N_610,N_731);
nor U848 (N_848,N_624,N_676);
and U849 (N_849,N_618,N_631);
xor U850 (N_850,N_797,N_698);
nor U851 (N_851,N_714,N_791);
nor U852 (N_852,N_785,N_775);
or U853 (N_853,N_665,N_666);
nand U854 (N_854,N_794,N_641);
and U855 (N_855,N_789,N_655);
and U856 (N_856,N_679,N_700);
nand U857 (N_857,N_712,N_619);
nor U858 (N_858,N_681,N_758);
or U859 (N_859,N_790,N_625);
or U860 (N_860,N_779,N_798);
nand U861 (N_861,N_723,N_744);
nand U862 (N_862,N_612,N_611);
and U863 (N_863,N_673,N_745);
nand U864 (N_864,N_767,N_711);
nor U865 (N_865,N_639,N_615);
or U866 (N_866,N_771,N_663);
nand U867 (N_867,N_616,N_739);
nand U868 (N_868,N_601,N_749);
or U869 (N_869,N_662,N_757);
or U870 (N_870,N_629,N_702);
and U871 (N_871,N_796,N_709);
and U872 (N_872,N_751,N_656);
nand U873 (N_873,N_704,N_746);
xnor U874 (N_874,N_734,N_691);
xnor U875 (N_875,N_678,N_766);
and U876 (N_876,N_643,N_760);
nand U877 (N_877,N_613,N_706);
or U878 (N_878,N_688,N_674);
nor U879 (N_879,N_650,N_668);
nand U880 (N_880,N_646,N_773);
and U881 (N_881,N_715,N_628);
and U882 (N_882,N_635,N_637);
xnor U883 (N_883,N_713,N_740);
nand U884 (N_884,N_710,N_677);
nand U885 (N_885,N_786,N_689);
or U886 (N_886,N_636,N_623);
xnor U887 (N_887,N_660,N_703);
nand U888 (N_888,N_605,N_752);
or U889 (N_889,N_667,N_718);
nor U890 (N_890,N_661,N_768);
xor U891 (N_891,N_728,N_600);
and U892 (N_892,N_630,N_753);
nand U893 (N_893,N_795,N_784);
nand U894 (N_894,N_721,N_644);
xnor U895 (N_895,N_671,N_781);
or U896 (N_896,N_696,N_604);
nor U897 (N_897,N_763,N_614);
nand U898 (N_898,N_609,N_647);
nand U899 (N_899,N_780,N_653);
or U900 (N_900,N_602,N_716);
xor U901 (N_901,N_687,N_757);
and U902 (N_902,N_771,N_676);
or U903 (N_903,N_629,N_751);
and U904 (N_904,N_727,N_639);
nand U905 (N_905,N_633,N_682);
or U906 (N_906,N_600,N_786);
nand U907 (N_907,N_759,N_778);
xor U908 (N_908,N_755,N_678);
or U909 (N_909,N_761,N_714);
and U910 (N_910,N_713,N_704);
xor U911 (N_911,N_622,N_605);
or U912 (N_912,N_619,N_644);
xnor U913 (N_913,N_767,N_606);
xor U914 (N_914,N_625,N_674);
and U915 (N_915,N_671,N_660);
nand U916 (N_916,N_704,N_675);
and U917 (N_917,N_680,N_629);
nand U918 (N_918,N_764,N_701);
or U919 (N_919,N_730,N_635);
or U920 (N_920,N_604,N_621);
and U921 (N_921,N_748,N_627);
nor U922 (N_922,N_604,N_725);
and U923 (N_923,N_706,N_644);
and U924 (N_924,N_663,N_709);
or U925 (N_925,N_639,N_779);
xnor U926 (N_926,N_626,N_677);
xor U927 (N_927,N_634,N_722);
and U928 (N_928,N_600,N_726);
xnor U929 (N_929,N_621,N_755);
nor U930 (N_930,N_645,N_682);
xnor U931 (N_931,N_787,N_794);
nand U932 (N_932,N_656,N_729);
or U933 (N_933,N_606,N_683);
nand U934 (N_934,N_615,N_628);
and U935 (N_935,N_665,N_703);
or U936 (N_936,N_704,N_618);
nand U937 (N_937,N_654,N_611);
nand U938 (N_938,N_642,N_763);
nand U939 (N_939,N_683,N_725);
xor U940 (N_940,N_699,N_628);
xor U941 (N_941,N_778,N_627);
nand U942 (N_942,N_623,N_685);
nor U943 (N_943,N_655,N_753);
xor U944 (N_944,N_779,N_664);
nor U945 (N_945,N_714,N_726);
nand U946 (N_946,N_664,N_687);
nor U947 (N_947,N_699,N_652);
xnor U948 (N_948,N_741,N_677);
nor U949 (N_949,N_673,N_684);
nand U950 (N_950,N_790,N_779);
nand U951 (N_951,N_752,N_603);
nor U952 (N_952,N_799,N_710);
xnor U953 (N_953,N_663,N_778);
or U954 (N_954,N_718,N_760);
nand U955 (N_955,N_614,N_625);
xor U956 (N_956,N_790,N_739);
or U957 (N_957,N_626,N_609);
or U958 (N_958,N_735,N_774);
nor U959 (N_959,N_698,N_731);
nand U960 (N_960,N_772,N_776);
nand U961 (N_961,N_617,N_745);
nor U962 (N_962,N_669,N_670);
and U963 (N_963,N_778,N_746);
xnor U964 (N_964,N_756,N_694);
or U965 (N_965,N_666,N_729);
nand U966 (N_966,N_642,N_754);
xnor U967 (N_967,N_602,N_780);
nor U968 (N_968,N_660,N_707);
nand U969 (N_969,N_692,N_732);
or U970 (N_970,N_652,N_637);
and U971 (N_971,N_654,N_747);
nand U972 (N_972,N_604,N_671);
xor U973 (N_973,N_614,N_623);
xor U974 (N_974,N_604,N_609);
nor U975 (N_975,N_796,N_700);
and U976 (N_976,N_649,N_747);
nor U977 (N_977,N_612,N_720);
xnor U978 (N_978,N_703,N_720);
nor U979 (N_979,N_765,N_791);
or U980 (N_980,N_660,N_686);
nand U981 (N_981,N_680,N_642);
and U982 (N_982,N_694,N_678);
nand U983 (N_983,N_649,N_795);
or U984 (N_984,N_612,N_758);
nand U985 (N_985,N_776,N_713);
or U986 (N_986,N_622,N_781);
nor U987 (N_987,N_669,N_700);
or U988 (N_988,N_771,N_781);
nand U989 (N_989,N_754,N_751);
and U990 (N_990,N_653,N_702);
nand U991 (N_991,N_756,N_622);
or U992 (N_992,N_605,N_685);
nor U993 (N_993,N_617,N_783);
and U994 (N_994,N_642,N_663);
and U995 (N_995,N_742,N_639);
nor U996 (N_996,N_684,N_794);
nand U997 (N_997,N_676,N_699);
or U998 (N_998,N_722,N_776);
or U999 (N_999,N_738,N_794);
or U1000 (N_1000,N_961,N_980);
or U1001 (N_1001,N_854,N_890);
nor U1002 (N_1002,N_814,N_923);
and U1003 (N_1003,N_835,N_971);
nand U1004 (N_1004,N_896,N_869);
and U1005 (N_1005,N_800,N_990);
nand U1006 (N_1006,N_924,N_902);
and U1007 (N_1007,N_852,N_839);
or U1008 (N_1008,N_843,N_982);
xnor U1009 (N_1009,N_930,N_859);
nand U1010 (N_1010,N_891,N_948);
nand U1011 (N_1011,N_880,N_874);
nor U1012 (N_1012,N_818,N_806);
or U1013 (N_1013,N_953,N_870);
and U1014 (N_1014,N_824,N_809);
and U1015 (N_1015,N_978,N_884);
and U1016 (N_1016,N_872,N_855);
and U1017 (N_1017,N_932,N_865);
nand U1018 (N_1018,N_974,N_899);
or U1019 (N_1019,N_907,N_949);
nor U1020 (N_1020,N_937,N_986);
xor U1021 (N_1021,N_813,N_850);
nand U1022 (N_1022,N_952,N_936);
and U1023 (N_1023,N_917,N_901);
nor U1024 (N_1024,N_941,N_878);
and U1025 (N_1025,N_885,N_864);
nor U1026 (N_1026,N_807,N_987);
nor U1027 (N_1027,N_945,N_996);
nand U1028 (N_1028,N_916,N_886);
nor U1029 (N_1029,N_808,N_900);
and U1030 (N_1030,N_960,N_823);
xnor U1031 (N_1031,N_810,N_938);
xor U1032 (N_1032,N_903,N_909);
nor U1033 (N_1033,N_956,N_889);
and U1034 (N_1034,N_993,N_841);
nor U1035 (N_1035,N_848,N_828);
and U1036 (N_1036,N_820,N_867);
or U1037 (N_1037,N_860,N_853);
or U1038 (N_1038,N_959,N_910);
and U1039 (N_1039,N_933,N_888);
nor U1040 (N_1040,N_929,N_887);
and U1041 (N_1041,N_825,N_955);
and U1042 (N_1042,N_877,N_829);
nand U1043 (N_1043,N_881,N_898);
and U1044 (N_1044,N_897,N_816);
and U1045 (N_1045,N_995,N_983);
nand U1046 (N_1046,N_926,N_908);
xnor U1047 (N_1047,N_866,N_946);
or U1048 (N_1048,N_992,N_973);
xnor U1049 (N_1049,N_939,N_943);
or U1050 (N_1050,N_944,N_957);
xnor U1051 (N_1051,N_803,N_914);
and U1052 (N_1052,N_912,N_970);
nor U1053 (N_1053,N_940,N_984);
nor U1054 (N_1054,N_882,N_951);
nand U1055 (N_1055,N_994,N_858);
nand U1056 (N_1056,N_845,N_827);
xnor U1057 (N_1057,N_977,N_892);
nand U1058 (N_1058,N_964,N_906);
or U1059 (N_1059,N_849,N_817);
nor U1060 (N_1060,N_947,N_851);
or U1061 (N_1061,N_921,N_991);
nand U1062 (N_1062,N_805,N_833);
or U1063 (N_1063,N_904,N_861);
nand U1064 (N_1064,N_975,N_966);
or U1065 (N_1065,N_918,N_837);
and U1066 (N_1066,N_875,N_963);
nand U1067 (N_1067,N_811,N_804);
xor U1068 (N_1068,N_831,N_913);
nor U1069 (N_1069,N_801,N_979);
and U1070 (N_1070,N_962,N_942);
nand U1071 (N_1071,N_838,N_997);
nor U1072 (N_1072,N_931,N_830);
and U1073 (N_1073,N_883,N_895);
xnor U1074 (N_1074,N_998,N_863);
xor U1075 (N_1075,N_935,N_972);
nand U1076 (N_1076,N_812,N_976);
xnor U1077 (N_1077,N_868,N_844);
nand U1078 (N_1078,N_919,N_950);
xnor U1079 (N_1079,N_989,N_846);
xnor U1080 (N_1080,N_842,N_922);
and U1081 (N_1081,N_840,N_894);
xnor U1082 (N_1082,N_915,N_965);
or U1083 (N_1083,N_819,N_847);
or U1084 (N_1084,N_815,N_985);
nand U1085 (N_1085,N_857,N_832);
nor U1086 (N_1086,N_834,N_822);
nor U1087 (N_1087,N_969,N_958);
or U1088 (N_1088,N_836,N_920);
nor U1089 (N_1089,N_999,N_934);
nor U1090 (N_1090,N_927,N_928);
nor U1091 (N_1091,N_856,N_826);
or U1092 (N_1092,N_911,N_988);
xnor U1093 (N_1093,N_821,N_981);
and U1094 (N_1094,N_862,N_879);
nor U1095 (N_1095,N_876,N_905);
nand U1096 (N_1096,N_967,N_968);
nor U1097 (N_1097,N_893,N_871);
xor U1098 (N_1098,N_873,N_925);
xor U1099 (N_1099,N_802,N_954);
nor U1100 (N_1100,N_846,N_991);
and U1101 (N_1101,N_833,N_927);
and U1102 (N_1102,N_900,N_997);
nor U1103 (N_1103,N_906,N_896);
nand U1104 (N_1104,N_914,N_937);
nor U1105 (N_1105,N_876,N_930);
or U1106 (N_1106,N_995,N_810);
and U1107 (N_1107,N_876,N_824);
and U1108 (N_1108,N_966,N_904);
and U1109 (N_1109,N_902,N_968);
nand U1110 (N_1110,N_942,N_937);
nor U1111 (N_1111,N_874,N_996);
or U1112 (N_1112,N_863,N_874);
nand U1113 (N_1113,N_803,N_895);
or U1114 (N_1114,N_970,N_887);
xnor U1115 (N_1115,N_832,N_821);
nor U1116 (N_1116,N_922,N_846);
xor U1117 (N_1117,N_884,N_972);
nor U1118 (N_1118,N_833,N_884);
xor U1119 (N_1119,N_900,N_922);
nand U1120 (N_1120,N_966,N_909);
or U1121 (N_1121,N_952,N_879);
and U1122 (N_1122,N_993,N_857);
or U1123 (N_1123,N_966,N_944);
nor U1124 (N_1124,N_919,N_932);
or U1125 (N_1125,N_809,N_901);
xnor U1126 (N_1126,N_879,N_802);
xor U1127 (N_1127,N_902,N_812);
or U1128 (N_1128,N_876,N_911);
or U1129 (N_1129,N_919,N_941);
nor U1130 (N_1130,N_972,N_810);
and U1131 (N_1131,N_983,N_988);
nand U1132 (N_1132,N_957,N_878);
nand U1133 (N_1133,N_984,N_915);
nand U1134 (N_1134,N_979,N_934);
and U1135 (N_1135,N_871,N_846);
xor U1136 (N_1136,N_947,N_862);
nor U1137 (N_1137,N_864,N_860);
or U1138 (N_1138,N_977,N_910);
and U1139 (N_1139,N_916,N_847);
xnor U1140 (N_1140,N_832,N_906);
or U1141 (N_1141,N_923,N_836);
nand U1142 (N_1142,N_928,N_966);
nand U1143 (N_1143,N_969,N_820);
and U1144 (N_1144,N_815,N_957);
or U1145 (N_1145,N_812,N_977);
nor U1146 (N_1146,N_871,N_982);
and U1147 (N_1147,N_853,N_885);
xnor U1148 (N_1148,N_909,N_857);
and U1149 (N_1149,N_876,N_836);
nand U1150 (N_1150,N_974,N_823);
xnor U1151 (N_1151,N_801,N_812);
and U1152 (N_1152,N_878,N_888);
xor U1153 (N_1153,N_970,N_836);
nand U1154 (N_1154,N_930,N_879);
xor U1155 (N_1155,N_931,N_947);
and U1156 (N_1156,N_912,N_824);
nor U1157 (N_1157,N_804,N_960);
or U1158 (N_1158,N_842,N_831);
nand U1159 (N_1159,N_933,N_932);
or U1160 (N_1160,N_985,N_954);
or U1161 (N_1161,N_869,N_958);
nand U1162 (N_1162,N_808,N_963);
nor U1163 (N_1163,N_924,N_921);
xnor U1164 (N_1164,N_939,N_969);
and U1165 (N_1165,N_932,N_970);
and U1166 (N_1166,N_957,N_866);
or U1167 (N_1167,N_980,N_987);
or U1168 (N_1168,N_927,N_803);
or U1169 (N_1169,N_854,N_868);
xnor U1170 (N_1170,N_942,N_801);
nand U1171 (N_1171,N_984,N_858);
and U1172 (N_1172,N_836,N_834);
nor U1173 (N_1173,N_930,N_972);
nand U1174 (N_1174,N_992,N_985);
xor U1175 (N_1175,N_964,N_991);
and U1176 (N_1176,N_807,N_959);
or U1177 (N_1177,N_996,N_891);
nor U1178 (N_1178,N_924,N_896);
nand U1179 (N_1179,N_972,N_952);
xnor U1180 (N_1180,N_947,N_913);
or U1181 (N_1181,N_980,N_862);
and U1182 (N_1182,N_990,N_858);
or U1183 (N_1183,N_946,N_819);
or U1184 (N_1184,N_813,N_834);
or U1185 (N_1185,N_969,N_968);
or U1186 (N_1186,N_984,N_834);
nor U1187 (N_1187,N_884,N_832);
xor U1188 (N_1188,N_991,N_975);
or U1189 (N_1189,N_955,N_808);
nand U1190 (N_1190,N_926,N_922);
and U1191 (N_1191,N_829,N_889);
xnor U1192 (N_1192,N_875,N_970);
xnor U1193 (N_1193,N_839,N_855);
or U1194 (N_1194,N_831,N_845);
nor U1195 (N_1195,N_836,N_965);
nor U1196 (N_1196,N_961,N_817);
and U1197 (N_1197,N_819,N_916);
nor U1198 (N_1198,N_867,N_895);
or U1199 (N_1199,N_854,N_849);
nand U1200 (N_1200,N_1146,N_1032);
and U1201 (N_1201,N_1067,N_1093);
xor U1202 (N_1202,N_1052,N_1091);
or U1203 (N_1203,N_1018,N_1153);
and U1204 (N_1204,N_1169,N_1098);
or U1205 (N_1205,N_1001,N_1117);
nand U1206 (N_1206,N_1081,N_1128);
and U1207 (N_1207,N_1180,N_1078);
or U1208 (N_1208,N_1171,N_1121);
and U1209 (N_1209,N_1134,N_1050);
and U1210 (N_1210,N_1163,N_1111);
nor U1211 (N_1211,N_1149,N_1004);
nor U1212 (N_1212,N_1104,N_1123);
and U1213 (N_1213,N_1119,N_1063);
or U1214 (N_1214,N_1009,N_1089);
nand U1215 (N_1215,N_1110,N_1065);
nor U1216 (N_1216,N_1054,N_1141);
nand U1217 (N_1217,N_1184,N_1190);
or U1218 (N_1218,N_1040,N_1122);
xnor U1219 (N_1219,N_1112,N_1099);
and U1220 (N_1220,N_1088,N_1186);
and U1221 (N_1221,N_1114,N_1011);
or U1222 (N_1222,N_1116,N_1154);
xor U1223 (N_1223,N_1115,N_1191);
and U1224 (N_1224,N_1107,N_1138);
and U1225 (N_1225,N_1025,N_1181);
nor U1226 (N_1226,N_1042,N_1103);
nand U1227 (N_1227,N_1195,N_1158);
nand U1228 (N_1228,N_1064,N_1113);
xnor U1229 (N_1229,N_1159,N_1148);
xor U1230 (N_1230,N_1048,N_1027);
xor U1231 (N_1231,N_1192,N_1179);
or U1232 (N_1232,N_1071,N_1196);
and U1233 (N_1233,N_1022,N_1079);
nand U1234 (N_1234,N_1125,N_1068);
nand U1235 (N_1235,N_1132,N_1036);
and U1236 (N_1236,N_1030,N_1076);
and U1237 (N_1237,N_1057,N_1150);
or U1238 (N_1238,N_1177,N_1198);
nand U1239 (N_1239,N_1126,N_1096);
xor U1240 (N_1240,N_1189,N_1167);
nor U1241 (N_1241,N_1188,N_1014);
nor U1242 (N_1242,N_1162,N_1173);
nand U1243 (N_1243,N_1017,N_1072);
and U1244 (N_1244,N_1194,N_1049);
and U1245 (N_1245,N_1174,N_1140);
nor U1246 (N_1246,N_1170,N_1015);
nor U1247 (N_1247,N_1039,N_1199);
xnor U1248 (N_1248,N_1092,N_1124);
xnor U1249 (N_1249,N_1016,N_1108);
nand U1250 (N_1250,N_1130,N_1183);
or U1251 (N_1251,N_1164,N_1034);
or U1252 (N_1252,N_1035,N_1145);
or U1253 (N_1253,N_1106,N_1021);
nor U1254 (N_1254,N_1005,N_1053);
xnor U1255 (N_1255,N_1043,N_1031);
or U1256 (N_1256,N_1129,N_1058);
nor U1257 (N_1257,N_1139,N_1070);
xor U1258 (N_1258,N_1037,N_1143);
nand U1259 (N_1259,N_1097,N_1008);
and U1260 (N_1260,N_1012,N_1073);
nor U1261 (N_1261,N_1080,N_1029);
and U1262 (N_1262,N_1055,N_1010);
or U1263 (N_1263,N_1155,N_1087);
or U1264 (N_1264,N_1028,N_1193);
nand U1265 (N_1265,N_1044,N_1136);
xnor U1266 (N_1266,N_1175,N_1045);
nand U1267 (N_1267,N_1061,N_1095);
nand U1268 (N_1268,N_1056,N_1075);
nor U1269 (N_1269,N_1182,N_1133);
nand U1270 (N_1270,N_1038,N_1041);
xnor U1271 (N_1271,N_1176,N_1074);
xor U1272 (N_1272,N_1156,N_1168);
nor U1273 (N_1273,N_1102,N_1127);
xor U1274 (N_1274,N_1051,N_1152);
and U1275 (N_1275,N_1135,N_1178);
nand U1276 (N_1276,N_1185,N_1142);
nand U1277 (N_1277,N_1019,N_1100);
nor U1278 (N_1278,N_1131,N_1109);
or U1279 (N_1279,N_1082,N_1033);
nand U1280 (N_1280,N_1062,N_1060);
or U1281 (N_1281,N_1144,N_1084);
nand U1282 (N_1282,N_1105,N_1000);
nor U1283 (N_1283,N_1069,N_1003);
and U1284 (N_1284,N_1059,N_1187);
nor U1285 (N_1285,N_1118,N_1006);
and U1286 (N_1286,N_1086,N_1090);
nor U1287 (N_1287,N_1047,N_1077);
or U1288 (N_1288,N_1160,N_1013);
nor U1289 (N_1289,N_1066,N_1101);
xor U1290 (N_1290,N_1083,N_1197);
xnor U1291 (N_1291,N_1147,N_1085);
and U1292 (N_1292,N_1157,N_1166);
or U1293 (N_1293,N_1094,N_1002);
nor U1294 (N_1294,N_1046,N_1172);
nor U1295 (N_1295,N_1120,N_1165);
xor U1296 (N_1296,N_1024,N_1020);
nor U1297 (N_1297,N_1026,N_1137);
xnor U1298 (N_1298,N_1023,N_1007);
or U1299 (N_1299,N_1161,N_1151);
nor U1300 (N_1300,N_1008,N_1015);
nand U1301 (N_1301,N_1023,N_1134);
xnor U1302 (N_1302,N_1004,N_1070);
or U1303 (N_1303,N_1001,N_1146);
and U1304 (N_1304,N_1177,N_1039);
xor U1305 (N_1305,N_1025,N_1142);
or U1306 (N_1306,N_1075,N_1153);
or U1307 (N_1307,N_1195,N_1086);
nand U1308 (N_1308,N_1088,N_1170);
or U1309 (N_1309,N_1181,N_1030);
and U1310 (N_1310,N_1018,N_1077);
xor U1311 (N_1311,N_1048,N_1012);
and U1312 (N_1312,N_1028,N_1088);
xor U1313 (N_1313,N_1097,N_1018);
or U1314 (N_1314,N_1127,N_1041);
and U1315 (N_1315,N_1193,N_1055);
xnor U1316 (N_1316,N_1197,N_1170);
nand U1317 (N_1317,N_1172,N_1159);
xor U1318 (N_1318,N_1127,N_1089);
and U1319 (N_1319,N_1000,N_1197);
nor U1320 (N_1320,N_1195,N_1137);
xor U1321 (N_1321,N_1166,N_1117);
xor U1322 (N_1322,N_1102,N_1170);
nor U1323 (N_1323,N_1049,N_1173);
xnor U1324 (N_1324,N_1152,N_1043);
xor U1325 (N_1325,N_1116,N_1016);
nor U1326 (N_1326,N_1104,N_1183);
or U1327 (N_1327,N_1043,N_1104);
and U1328 (N_1328,N_1173,N_1005);
or U1329 (N_1329,N_1072,N_1065);
nor U1330 (N_1330,N_1140,N_1064);
and U1331 (N_1331,N_1159,N_1150);
or U1332 (N_1332,N_1104,N_1170);
and U1333 (N_1333,N_1167,N_1040);
nand U1334 (N_1334,N_1124,N_1050);
or U1335 (N_1335,N_1063,N_1010);
nand U1336 (N_1336,N_1146,N_1149);
or U1337 (N_1337,N_1038,N_1096);
nor U1338 (N_1338,N_1023,N_1093);
and U1339 (N_1339,N_1067,N_1057);
xor U1340 (N_1340,N_1044,N_1098);
nor U1341 (N_1341,N_1036,N_1086);
and U1342 (N_1342,N_1133,N_1007);
nand U1343 (N_1343,N_1073,N_1150);
nand U1344 (N_1344,N_1014,N_1117);
nand U1345 (N_1345,N_1007,N_1140);
nor U1346 (N_1346,N_1042,N_1047);
nor U1347 (N_1347,N_1185,N_1052);
nand U1348 (N_1348,N_1110,N_1040);
or U1349 (N_1349,N_1118,N_1122);
xor U1350 (N_1350,N_1040,N_1022);
xor U1351 (N_1351,N_1129,N_1172);
or U1352 (N_1352,N_1117,N_1192);
nand U1353 (N_1353,N_1152,N_1052);
nand U1354 (N_1354,N_1083,N_1043);
xor U1355 (N_1355,N_1179,N_1003);
xnor U1356 (N_1356,N_1159,N_1136);
xnor U1357 (N_1357,N_1156,N_1189);
or U1358 (N_1358,N_1037,N_1112);
or U1359 (N_1359,N_1027,N_1034);
and U1360 (N_1360,N_1137,N_1054);
or U1361 (N_1361,N_1179,N_1056);
nand U1362 (N_1362,N_1086,N_1098);
xor U1363 (N_1363,N_1077,N_1190);
nor U1364 (N_1364,N_1049,N_1096);
nand U1365 (N_1365,N_1173,N_1086);
and U1366 (N_1366,N_1117,N_1062);
and U1367 (N_1367,N_1007,N_1044);
nor U1368 (N_1368,N_1008,N_1099);
nand U1369 (N_1369,N_1150,N_1124);
nand U1370 (N_1370,N_1108,N_1120);
nor U1371 (N_1371,N_1034,N_1009);
nor U1372 (N_1372,N_1183,N_1181);
nor U1373 (N_1373,N_1010,N_1175);
and U1374 (N_1374,N_1149,N_1109);
or U1375 (N_1375,N_1175,N_1020);
or U1376 (N_1376,N_1120,N_1008);
and U1377 (N_1377,N_1142,N_1155);
nand U1378 (N_1378,N_1162,N_1077);
nand U1379 (N_1379,N_1110,N_1026);
or U1380 (N_1380,N_1175,N_1113);
and U1381 (N_1381,N_1051,N_1054);
nand U1382 (N_1382,N_1130,N_1005);
or U1383 (N_1383,N_1173,N_1199);
nand U1384 (N_1384,N_1058,N_1013);
nor U1385 (N_1385,N_1057,N_1030);
or U1386 (N_1386,N_1118,N_1127);
nand U1387 (N_1387,N_1078,N_1041);
and U1388 (N_1388,N_1041,N_1176);
nor U1389 (N_1389,N_1097,N_1145);
and U1390 (N_1390,N_1188,N_1169);
and U1391 (N_1391,N_1134,N_1084);
xnor U1392 (N_1392,N_1035,N_1168);
or U1393 (N_1393,N_1062,N_1154);
nor U1394 (N_1394,N_1031,N_1145);
nand U1395 (N_1395,N_1003,N_1009);
xor U1396 (N_1396,N_1013,N_1176);
nor U1397 (N_1397,N_1187,N_1031);
and U1398 (N_1398,N_1042,N_1086);
xnor U1399 (N_1399,N_1121,N_1024);
or U1400 (N_1400,N_1281,N_1204);
and U1401 (N_1401,N_1262,N_1258);
nand U1402 (N_1402,N_1337,N_1219);
nor U1403 (N_1403,N_1313,N_1330);
nor U1404 (N_1404,N_1344,N_1268);
nor U1405 (N_1405,N_1238,N_1240);
and U1406 (N_1406,N_1282,N_1208);
or U1407 (N_1407,N_1353,N_1247);
nor U1408 (N_1408,N_1320,N_1211);
xor U1409 (N_1409,N_1273,N_1260);
nand U1410 (N_1410,N_1371,N_1249);
or U1411 (N_1411,N_1373,N_1386);
xor U1412 (N_1412,N_1316,N_1291);
or U1413 (N_1413,N_1216,N_1251);
and U1414 (N_1414,N_1221,N_1252);
xor U1415 (N_1415,N_1305,N_1369);
nand U1416 (N_1416,N_1376,N_1379);
nor U1417 (N_1417,N_1389,N_1237);
xnor U1418 (N_1418,N_1399,N_1235);
and U1419 (N_1419,N_1390,N_1383);
nor U1420 (N_1420,N_1334,N_1246);
or U1421 (N_1421,N_1375,N_1349);
and U1422 (N_1422,N_1277,N_1362);
or U1423 (N_1423,N_1385,N_1239);
nor U1424 (N_1424,N_1271,N_1321);
xnor U1425 (N_1425,N_1367,N_1307);
or U1426 (N_1426,N_1299,N_1267);
and U1427 (N_1427,N_1265,N_1361);
nand U1428 (N_1428,N_1276,N_1377);
xor U1429 (N_1429,N_1359,N_1311);
xnor U1430 (N_1430,N_1236,N_1279);
nor U1431 (N_1431,N_1205,N_1290);
nand U1432 (N_1432,N_1333,N_1241);
xor U1433 (N_1433,N_1336,N_1210);
and U1434 (N_1434,N_1254,N_1278);
nor U1435 (N_1435,N_1222,N_1341);
xnor U1436 (N_1436,N_1326,N_1253);
xor U1437 (N_1437,N_1209,N_1374);
xor U1438 (N_1438,N_1391,N_1248);
and U1439 (N_1439,N_1229,N_1308);
nand U1440 (N_1440,N_1306,N_1275);
nand U1441 (N_1441,N_1263,N_1225);
and U1442 (N_1442,N_1200,N_1244);
xnor U1443 (N_1443,N_1280,N_1212);
and U1444 (N_1444,N_1342,N_1346);
or U1445 (N_1445,N_1380,N_1310);
or U1446 (N_1446,N_1269,N_1365);
and U1447 (N_1447,N_1231,N_1207);
or U1448 (N_1448,N_1245,N_1259);
xnor U1449 (N_1449,N_1398,N_1360);
or U1450 (N_1450,N_1256,N_1312);
nor U1451 (N_1451,N_1227,N_1345);
nand U1452 (N_1452,N_1397,N_1234);
and U1453 (N_1453,N_1315,N_1351);
nor U1454 (N_1454,N_1348,N_1220);
nor U1455 (N_1455,N_1352,N_1395);
or U1456 (N_1456,N_1270,N_1230);
and U1457 (N_1457,N_1301,N_1224);
nand U1458 (N_1458,N_1382,N_1228);
nor U1459 (N_1459,N_1203,N_1257);
or U1460 (N_1460,N_1293,N_1296);
or U1461 (N_1461,N_1322,N_1366);
xnor U1462 (N_1462,N_1232,N_1288);
xnor U1463 (N_1463,N_1294,N_1388);
and U1464 (N_1464,N_1350,N_1226);
or U1465 (N_1465,N_1242,N_1327);
nand U1466 (N_1466,N_1370,N_1261);
and U1467 (N_1467,N_1319,N_1378);
nand U1468 (N_1468,N_1392,N_1300);
nand U1469 (N_1469,N_1338,N_1340);
nor U1470 (N_1470,N_1297,N_1202);
and U1471 (N_1471,N_1214,N_1303);
or U1472 (N_1472,N_1201,N_1285);
nand U1473 (N_1473,N_1272,N_1335);
nor U1474 (N_1474,N_1358,N_1217);
or U1475 (N_1475,N_1381,N_1304);
nor U1476 (N_1476,N_1283,N_1324);
and U1477 (N_1477,N_1266,N_1309);
nor U1478 (N_1478,N_1368,N_1331);
xor U1479 (N_1479,N_1325,N_1287);
or U1480 (N_1480,N_1223,N_1289);
nor U1481 (N_1481,N_1292,N_1355);
or U1482 (N_1482,N_1393,N_1332);
or U1483 (N_1483,N_1356,N_1364);
nand U1484 (N_1484,N_1243,N_1357);
and U1485 (N_1485,N_1396,N_1218);
and U1486 (N_1486,N_1329,N_1274);
and U1487 (N_1487,N_1284,N_1215);
and U1488 (N_1488,N_1264,N_1233);
nor U1489 (N_1489,N_1286,N_1328);
nand U1490 (N_1490,N_1347,N_1372);
and U1491 (N_1491,N_1384,N_1298);
and U1492 (N_1492,N_1302,N_1363);
or U1493 (N_1493,N_1387,N_1354);
nor U1494 (N_1494,N_1295,N_1255);
xnor U1495 (N_1495,N_1250,N_1339);
and U1496 (N_1496,N_1317,N_1318);
nand U1497 (N_1497,N_1394,N_1343);
xnor U1498 (N_1498,N_1314,N_1323);
and U1499 (N_1499,N_1206,N_1213);
and U1500 (N_1500,N_1371,N_1298);
nor U1501 (N_1501,N_1286,N_1331);
or U1502 (N_1502,N_1360,N_1309);
nand U1503 (N_1503,N_1297,N_1366);
nor U1504 (N_1504,N_1208,N_1257);
or U1505 (N_1505,N_1325,N_1326);
and U1506 (N_1506,N_1256,N_1351);
nor U1507 (N_1507,N_1254,N_1335);
nor U1508 (N_1508,N_1376,N_1302);
and U1509 (N_1509,N_1219,N_1289);
xor U1510 (N_1510,N_1369,N_1296);
nand U1511 (N_1511,N_1349,N_1324);
nand U1512 (N_1512,N_1239,N_1209);
nor U1513 (N_1513,N_1303,N_1348);
nor U1514 (N_1514,N_1201,N_1347);
xnor U1515 (N_1515,N_1390,N_1396);
nor U1516 (N_1516,N_1242,N_1379);
nor U1517 (N_1517,N_1375,N_1389);
and U1518 (N_1518,N_1329,N_1261);
nand U1519 (N_1519,N_1287,N_1269);
nor U1520 (N_1520,N_1342,N_1394);
nand U1521 (N_1521,N_1315,N_1258);
nor U1522 (N_1522,N_1232,N_1397);
and U1523 (N_1523,N_1326,N_1221);
nor U1524 (N_1524,N_1233,N_1376);
or U1525 (N_1525,N_1246,N_1277);
or U1526 (N_1526,N_1277,N_1339);
and U1527 (N_1527,N_1336,N_1317);
and U1528 (N_1528,N_1220,N_1218);
nand U1529 (N_1529,N_1362,N_1315);
nor U1530 (N_1530,N_1222,N_1205);
and U1531 (N_1531,N_1386,N_1337);
and U1532 (N_1532,N_1333,N_1374);
or U1533 (N_1533,N_1208,N_1286);
and U1534 (N_1534,N_1266,N_1229);
and U1535 (N_1535,N_1246,N_1368);
nand U1536 (N_1536,N_1228,N_1376);
nand U1537 (N_1537,N_1361,N_1253);
or U1538 (N_1538,N_1388,N_1231);
or U1539 (N_1539,N_1311,N_1276);
nor U1540 (N_1540,N_1272,N_1229);
nand U1541 (N_1541,N_1282,N_1319);
xnor U1542 (N_1542,N_1263,N_1224);
or U1543 (N_1543,N_1329,N_1387);
nor U1544 (N_1544,N_1220,N_1317);
and U1545 (N_1545,N_1229,N_1399);
nor U1546 (N_1546,N_1325,N_1379);
nand U1547 (N_1547,N_1347,N_1376);
or U1548 (N_1548,N_1352,N_1369);
nand U1549 (N_1549,N_1371,N_1239);
nand U1550 (N_1550,N_1340,N_1364);
xnor U1551 (N_1551,N_1267,N_1264);
nor U1552 (N_1552,N_1265,N_1215);
xor U1553 (N_1553,N_1259,N_1274);
xor U1554 (N_1554,N_1308,N_1396);
xnor U1555 (N_1555,N_1254,N_1325);
and U1556 (N_1556,N_1265,N_1208);
xnor U1557 (N_1557,N_1342,N_1371);
xor U1558 (N_1558,N_1361,N_1351);
or U1559 (N_1559,N_1375,N_1372);
xnor U1560 (N_1560,N_1304,N_1255);
nand U1561 (N_1561,N_1291,N_1228);
nand U1562 (N_1562,N_1201,N_1359);
or U1563 (N_1563,N_1333,N_1349);
and U1564 (N_1564,N_1363,N_1314);
nand U1565 (N_1565,N_1391,N_1395);
nor U1566 (N_1566,N_1390,N_1337);
and U1567 (N_1567,N_1227,N_1205);
and U1568 (N_1568,N_1386,N_1247);
nand U1569 (N_1569,N_1317,N_1313);
nor U1570 (N_1570,N_1297,N_1323);
nor U1571 (N_1571,N_1306,N_1395);
and U1572 (N_1572,N_1339,N_1321);
xor U1573 (N_1573,N_1352,N_1299);
xnor U1574 (N_1574,N_1368,N_1388);
and U1575 (N_1575,N_1256,N_1271);
or U1576 (N_1576,N_1347,N_1203);
or U1577 (N_1577,N_1271,N_1349);
and U1578 (N_1578,N_1250,N_1208);
or U1579 (N_1579,N_1244,N_1327);
xnor U1580 (N_1580,N_1355,N_1344);
nand U1581 (N_1581,N_1399,N_1307);
or U1582 (N_1582,N_1311,N_1233);
or U1583 (N_1583,N_1294,N_1398);
or U1584 (N_1584,N_1206,N_1376);
nor U1585 (N_1585,N_1334,N_1376);
nor U1586 (N_1586,N_1230,N_1316);
nand U1587 (N_1587,N_1366,N_1228);
xnor U1588 (N_1588,N_1292,N_1340);
nand U1589 (N_1589,N_1206,N_1382);
xor U1590 (N_1590,N_1332,N_1381);
and U1591 (N_1591,N_1394,N_1372);
nand U1592 (N_1592,N_1296,N_1349);
xnor U1593 (N_1593,N_1363,N_1326);
xnor U1594 (N_1594,N_1398,N_1367);
nor U1595 (N_1595,N_1391,N_1331);
nand U1596 (N_1596,N_1233,N_1302);
or U1597 (N_1597,N_1225,N_1345);
nor U1598 (N_1598,N_1368,N_1376);
or U1599 (N_1599,N_1299,N_1220);
and U1600 (N_1600,N_1590,N_1593);
nor U1601 (N_1601,N_1488,N_1573);
or U1602 (N_1602,N_1454,N_1476);
and U1603 (N_1603,N_1427,N_1560);
nand U1604 (N_1604,N_1457,N_1438);
or U1605 (N_1605,N_1518,N_1465);
xnor U1606 (N_1606,N_1406,N_1545);
or U1607 (N_1607,N_1410,N_1579);
nand U1608 (N_1608,N_1564,N_1402);
and U1609 (N_1609,N_1522,N_1539);
nor U1610 (N_1610,N_1581,N_1565);
and U1611 (N_1611,N_1469,N_1534);
nor U1612 (N_1612,N_1591,N_1481);
xnor U1613 (N_1613,N_1559,N_1415);
and U1614 (N_1614,N_1589,N_1507);
and U1615 (N_1615,N_1436,N_1434);
xor U1616 (N_1616,N_1414,N_1475);
nor U1617 (N_1617,N_1555,N_1541);
or U1618 (N_1618,N_1503,N_1405);
nor U1619 (N_1619,N_1568,N_1480);
nand U1620 (N_1620,N_1485,N_1474);
nor U1621 (N_1621,N_1597,N_1484);
nand U1622 (N_1622,N_1528,N_1420);
nor U1623 (N_1623,N_1463,N_1566);
xnor U1624 (N_1624,N_1458,N_1426);
or U1625 (N_1625,N_1595,N_1441);
and U1626 (N_1626,N_1431,N_1435);
xnor U1627 (N_1627,N_1504,N_1538);
and U1628 (N_1628,N_1482,N_1586);
xnor U1629 (N_1629,N_1417,N_1571);
xnor U1630 (N_1630,N_1547,N_1491);
xnor U1631 (N_1631,N_1498,N_1536);
and U1632 (N_1632,N_1502,N_1452);
nor U1633 (N_1633,N_1506,N_1442);
xnor U1634 (N_1634,N_1432,N_1455);
nor U1635 (N_1635,N_1527,N_1461);
xor U1636 (N_1636,N_1466,N_1421);
or U1637 (N_1637,N_1584,N_1514);
and U1638 (N_1638,N_1487,N_1412);
or U1639 (N_1639,N_1445,N_1429);
and U1640 (N_1640,N_1479,N_1513);
xor U1641 (N_1641,N_1501,N_1575);
xnor U1642 (N_1642,N_1599,N_1540);
or U1643 (N_1643,N_1400,N_1592);
or U1644 (N_1644,N_1567,N_1462);
or U1645 (N_1645,N_1447,N_1515);
and U1646 (N_1646,N_1508,N_1556);
nand U1647 (N_1647,N_1499,N_1428);
or U1648 (N_1648,N_1489,N_1585);
and U1649 (N_1649,N_1470,N_1587);
xor U1650 (N_1650,N_1443,N_1510);
nor U1651 (N_1651,N_1562,N_1509);
or U1652 (N_1652,N_1530,N_1588);
xnor U1653 (N_1653,N_1561,N_1425);
nor U1654 (N_1654,N_1492,N_1576);
or U1655 (N_1655,N_1598,N_1486);
and U1656 (N_1656,N_1582,N_1450);
nand U1657 (N_1657,N_1424,N_1549);
or U1658 (N_1658,N_1456,N_1558);
nor U1659 (N_1659,N_1516,N_1451);
or U1660 (N_1660,N_1529,N_1460);
xor U1661 (N_1661,N_1537,N_1533);
nand U1662 (N_1662,N_1594,N_1483);
nand U1663 (N_1663,N_1403,N_1563);
xnor U1664 (N_1664,N_1531,N_1446);
nand U1665 (N_1665,N_1496,N_1437);
nand U1666 (N_1666,N_1557,N_1543);
nor U1667 (N_1667,N_1577,N_1583);
xor U1668 (N_1668,N_1439,N_1548);
nand U1669 (N_1669,N_1574,N_1521);
or U1670 (N_1670,N_1493,N_1411);
nor U1671 (N_1671,N_1526,N_1550);
nand U1672 (N_1672,N_1430,N_1532);
or U1673 (N_1673,N_1497,N_1542);
and U1674 (N_1674,N_1449,N_1433);
and U1675 (N_1675,N_1495,N_1490);
and U1676 (N_1676,N_1517,N_1546);
or U1677 (N_1677,N_1448,N_1535);
nor U1678 (N_1678,N_1409,N_1578);
nor U1679 (N_1679,N_1404,N_1570);
and U1680 (N_1680,N_1471,N_1416);
xor U1681 (N_1681,N_1596,N_1418);
and U1682 (N_1682,N_1552,N_1569);
nor U1683 (N_1683,N_1444,N_1401);
or U1684 (N_1684,N_1467,N_1464);
xnor U1685 (N_1685,N_1477,N_1505);
nor U1686 (N_1686,N_1512,N_1544);
nand U1687 (N_1687,N_1572,N_1494);
or U1688 (N_1688,N_1524,N_1413);
nand U1689 (N_1689,N_1468,N_1459);
xor U1690 (N_1690,N_1500,N_1472);
nor U1691 (N_1691,N_1440,N_1419);
xnor U1692 (N_1692,N_1580,N_1553);
nor U1693 (N_1693,N_1525,N_1478);
and U1694 (N_1694,N_1519,N_1511);
nor U1695 (N_1695,N_1407,N_1453);
and U1696 (N_1696,N_1423,N_1523);
nor U1697 (N_1697,N_1520,N_1408);
or U1698 (N_1698,N_1473,N_1422);
and U1699 (N_1699,N_1554,N_1551);
or U1700 (N_1700,N_1591,N_1445);
nand U1701 (N_1701,N_1523,N_1584);
xnor U1702 (N_1702,N_1472,N_1497);
or U1703 (N_1703,N_1428,N_1454);
nand U1704 (N_1704,N_1426,N_1430);
nor U1705 (N_1705,N_1547,N_1418);
nand U1706 (N_1706,N_1544,N_1539);
and U1707 (N_1707,N_1567,N_1453);
and U1708 (N_1708,N_1405,N_1555);
and U1709 (N_1709,N_1595,N_1538);
nor U1710 (N_1710,N_1448,N_1598);
nand U1711 (N_1711,N_1532,N_1473);
xnor U1712 (N_1712,N_1598,N_1542);
xor U1713 (N_1713,N_1483,N_1569);
and U1714 (N_1714,N_1534,N_1594);
and U1715 (N_1715,N_1529,N_1535);
or U1716 (N_1716,N_1599,N_1503);
or U1717 (N_1717,N_1567,N_1583);
and U1718 (N_1718,N_1537,N_1421);
nand U1719 (N_1719,N_1538,N_1428);
xor U1720 (N_1720,N_1572,N_1538);
xnor U1721 (N_1721,N_1456,N_1549);
or U1722 (N_1722,N_1433,N_1568);
nor U1723 (N_1723,N_1545,N_1403);
nand U1724 (N_1724,N_1466,N_1498);
and U1725 (N_1725,N_1484,N_1517);
or U1726 (N_1726,N_1598,N_1427);
or U1727 (N_1727,N_1428,N_1501);
and U1728 (N_1728,N_1571,N_1558);
nor U1729 (N_1729,N_1511,N_1589);
and U1730 (N_1730,N_1461,N_1454);
or U1731 (N_1731,N_1595,N_1439);
or U1732 (N_1732,N_1400,N_1496);
nand U1733 (N_1733,N_1491,N_1568);
nand U1734 (N_1734,N_1420,N_1406);
nor U1735 (N_1735,N_1499,N_1514);
and U1736 (N_1736,N_1496,N_1558);
nor U1737 (N_1737,N_1527,N_1583);
nand U1738 (N_1738,N_1529,N_1556);
nand U1739 (N_1739,N_1427,N_1562);
nand U1740 (N_1740,N_1450,N_1491);
nor U1741 (N_1741,N_1587,N_1424);
nor U1742 (N_1742,N_1416,N_1539);
or U1743 (N_1743,N_1581,N_1579);
xnor U1744 (N_1744,N_1527,N_1561);
and U1745 (N_1745,N_1438,N_1509);
xor U1746 (N_1746,N_1404,N_1432);
or U1747 (N_1747,N_1539,N_1500);
nand U1748 (N_1748,N_1502,N_1562);
nor U1749 (N_1749,N_1485,N_1480);
and U1750 (N_1750,N_1589,N_1504);
nor U1751 (N_1751,N_1472,N_1428);
and U1752 (N_1752,N_1467,N_1566);
xnor U1753 (N_1753,N_1592,N_1556);
nand U1754 (N_1754,N_1453,N_1506);
or U1755 (N_1755,N_1558,N_1523);
or U1756 (N_1756,N_1419,N_1561);
nor U1757 (N_1757,N_1486,N_1491);
xnor U1758 (N_1758,N_1474,N_1472);
or U1759 (N_1759,N_1468,N_1529);
or U1760 (N_1760,N_1404,N_1564);
nand U1761 (N_1761,N_1446,N_1577);
and U1762 (N_1762,N_1406,N_1433);
nor U1763 (N_1763,N_1408,N_1563);
nand U1764 (N_1764,N_1458,N_1557);
nand U1765 (N_1765,N_1420,N_1513);
nor U1766 (N_1766,N_1439,N_1544);
and U1767 (N_1767,N_1503,N_1551);
xor U1768 (N_1768,N_1496,N_1453);
nand U1769 (N_1769,N_1475,N_1492);
and U1770 (N_1770,N_1472,N_1519);
nand U1771 (N_1771,N_1447,N_1596);
xnor U1772 (N_1772,N_1439,N_1562);
nor U1773 (N_1773,N_1419,N_1447);
nand U1774 (N_1774,N_1488,N_1578);
nand U1775 (N_1775,N_1553,N_1502);
nand U1776 (N_1776,N_1513,N_1579);
or U1777 (N_1777,N_1404,N_1434);
or U1778 (N_1778,N_1478,N_1581);
nor U1779 (N_1779,N_1512,N_1469);
nor U1780 (N_1780,N_1488,N_1501);
nor U1781 (N_1781,N_1557,N_1517);
xnor U1782 (N_1782,N_1487,N_1461);
nor U1783 (N_1783,N_1435,N_1467);
xnor U1784 (N_1784,N_1540,N_1564);
and U1785 (N_1785,N_1482,N_1467);
and U1786 (N_1786,N_1428,N_1434);
or U1787 (N_1787,N_1509,N_1573);
and U1788 (N_1788,N_1589,N_1436);
nand U1789 (N_1789,N_1475,N_1458);
and U1790 (N_1790,N_1591,N_1563);
nand U1791 (N_1791,N_1456,N_1412);
xnor U1792 (N_1792,N_1537,N_1591);
nor U1793 (N_1793,N_1447,N_1437);
or U1794 (N_1794,N_1449,N_1504);
nand U1795 (N_1795,N_1489,N_1505);
nor U1796 (N_1796,N_1552,N_1585);
xor U1797 (N_1797,N_1491,N_1519);
and U1798 (N_1798,N_1527,N_1501);
and U1799 (N_1799,N_1482,N_1462);
xnor U1800 (N_1800,N_1739,N_1693);
or U1801 (N_1801,N_1763,N_1720);
and U1802 (N_1802,N_1680,N_1627);
nor U1803 (N_1803,N_1766,N_1715);
xor U1804 (N_1804,N_1690,N_1607);
xor U1805 (N_1805,N_1610,N_1683);
and U1806 (N_1806,N_1788,N_1730);
nor U1807 (N_1807,N_1787,N_1692);
or U1808 (N_1808,N_1604,N_1784);
nand U1809 (N_1809,N_1716,N_1746);
nor U1810 (N_1810,N_1799,N_1762);
or U1811 (N_1811,N_1660,N_1719);
nand U1812 (N_1812,N_1758,N_1780);
xor U1813 (N_1813,N_1662,N_1779);
nand U1814 (N_1814,N_1653,N_1707);
xnor U1815 (N_1815,N_1616,N_1712);
or U1816 (N_1816,N_1760,N_1732);
nor U1817 (N_1817,N_1733,N_1635);
nor U1818 (N_1818,N_1731,N_1659);
nand U1819 (N_1819,N_1626,N_1698);
and U1820 (N_1820,N_1602,N_1646);
or U1821 (N_1821,N_1709,N_1771);
xor U1822 (N_1822,N_1710,N_1679);
nand U1823 (N_1823,N_1668,N_1754);
nor U1824 (N_1824,N_1657,N_1767);
and U1825 (N_1825,N_1783,N_1703);
nor U1826 (N_1826,N_1777,N_1745);
nor U1827 (N_1827,N_1724,N_1792);
nand U1828 (N_1828,N_1634,N_1648);
and U1829 (N_1829,N_1644,N_1773);
nor U1830 (N_1830,N_1614,N_1751);
nor U1831 (N_1831,N_1617,N_1681);
or U1832 (N_1832,N_1649,N_1661);
nand U1833 (N_1833,N_1785,N_1664);
and U1834 (N_1834,N_1714,N_1631);
and U1835 (N_1835,N_1689,N_1738);
nor U1836 (N_1836,N_1636,N_1797);
and U1837 (N_1837,N_1743,N_1633);
xor U1838 (N_1838,N_1639,N_1619);
xnor U1839 (N_1839,N_1670,N_1624);
nand U1840 (N_1840,N_1629,N_1700);
nand U1841 (N_1841,N_1694,N_1685);
xor U1842 (N_1842,N_1713,N_1729);
xor U1843 (N_1843,N_1711,N_1620);
nor U1844 (N_1844,N_1755,N_1641);
and U1845 (N_1845,N_1750,N_1618);
nor U1846 (N_1846,N_1782,N_1786);
xnor U1847 (N_1847,N_1674,N_1774);
nor U1848 (N_1848,N_1687,N_1625);
or U1849 (N_1849,N_1789,N_1726);
nor U1850 (N_1850,N_1621,N_1667);
nand U1851 (N_1851,N_1748,N_1752);
nand U1852 (N_1852,N_1706,N_1795);
and U1853 (N_1853,N_1672,N_1798);
nand U1854 (N_1854,N_1628,N_1718);
nor U1855 (N_1855,N_1622,N_1701);
xnor U1856 (N_1856,N_1736,N_1638);
nor U1857 (N_1857,N_1695,N_1765);
or U1858 (N_1858,N_1728,N_1704);
and U1859 (N_1859,N_1769,N_1640);
nand U1860 (N_1860,N_1725,N_1735);
xnor U1861 (N_1861,N_1761,N_1702);
and U1862 (N_1862,N_1645,N_1605);
nor U1863 (N_1863,N_1772,N_1722);
nor U1864 (N_1864,N_1642,N_1663);
xor U1865 (N_1865,N_1699,N_1630);
and U1866 (N_1866,N_1609,N_1790);
and U1867 (N_1867,N_1654,N_1611);
or U1868 (N_1868,N_1776,N_1734);
nor U1869 (N_1869,N_1775,N_1647);
nor U1870 (N_1870,N_1697,N_1656);
xnor U1871 (N_1871,N_1673,N_1666);
nand U1872 (N_1872,N_1793,N_1669);
xnor U1873 (N_1873,N_1612,N_1705);
xor U1874 (N_1874,N_1603,N_1658);
xnor U1875 (N_1875,N_1768,N_1791);
nor U1876 (N_1876,N_1675,N_1623);
nor U1877 (N_1877,N_1613,N_1688);
or U1878 (N_1878,N_1781,N_1671);
nand U1879 (N_1879,N_1637,N_1615);
nor U1880 (N_1880,N_1655,N_1606);
nor U1881 (N_1881,N_1665,N_1756);
xnor U1882 (N_1882,N_1749,N_1682);
xor U1883 (N_1883,N_1759,N_1796);
nor U1884 (N_1884,N_1770,N_1632);
and U1885 (N_1885,N_1643,N_1696);
nor U1886 (N_1886,N_1757,N_1686);
nand U1887 (N_1887,N_1778,N_1741);
xnor U1888 (N_1888,N_1652,N_1684);
or U1889 (N_1889,N_1600,N_1747);
or U1890 (N_1890,N_1678,N_1676);
nand U1891 (N_1891,N_1601,N_1744);
or U1892 (N_1892,N_1794,N_1764);
xnor U1893 (N_1893,N_1737,N_1717);
and U1894 (N_1894,N_1608,N_1651);
nor U1895 (N_1895,N_1740,N_1721);
xor U1896 (N_1896,N_1723,N_1742);
nor U1897 (N_1897,N_1727,N_1650);
nor U1898 (N_1898,N_1708,N_1677);
and U1899 (N_1899,N_1691,N_1753);
nand U1900 (N_1900,N_1622,N_1639);
nand U1901 (N_1901,N_1601,N_1777);
nor U1902 (N_1902,N_1697,N_1769);
or U1903 (N_1903,N_1756,N_1694);
nand U1904 (N_1904,N_1663,N_1601);
xor U1905 (N_1905,N_1681,N_1700);
or U1906 (N_1906,N_1605,N_1704);
xnor U1907 (N_1907,N_1720,N_1783);
or U1908 (N_1908,N_1688,N_1615);
xor U1909 (N_1909,N_1725,N_1624);
nor U1910 (N_1910,N_1645,N_1756);
or U1911 (N_1911,N_1744,N_1647);
nor U1912 (N_1912,N_1616,N_1741);
xnor U1913 (N_1913,N_1681,N_1657);
nand U1914 (N_1914,N_1717,N_1773);
nor U1915 (N_1915,N_1702,N_1719);
xnor U1916 (N_1916,N_1624,N_1632);
or U1917 (N_1917,N_1791,N_1718);
nand U1918 (N_1918,N_1787,N_1737);
nor U1919 (N_1919,N_1621,N_1717);
nand U1920 (N_1920,N_1758,N_1607);
or U1921 (N_1921,N_1726,N_1763);
nand U1922 (N_1922,N_1705,N_1726);
or U1923 (N_1923,N_1761,N_1604);
or U1924 (N_1924,N_1681,N_1650);
and U1925 (N_1925,N_1691,N_1687);
nand U1926 (N_1926,N_1783,N_1734);
or U1927 (N_1927,N_1674,N_1657);
and U1928 (N_1928,N_1611,N_1790);
nand U1929 (N_1929,N_1707,N_1758);
and U1930 (N_1930,N_1758,N_1682);
and U1931 (N_1931,N_1792,N_1612);
and U1932 (N_1932,N_1619,N_1701);
xnor U1933 (N_1933,N_1797,N_1688);
and U1934 (N_1934,N_1656,N_1717);
or U1935 (N_1935,N_1636,N_1724);
and U1936 (N_1936,N_1663,N_1643);
nand U1937 (N_1937,N_1746,N_1736);
or U1938 (N_1938,N_1762,N_1752);
xnor U1939 (N_1939,N_1771,N_1772);
or U1940 (N_1940,N_1741,N_1628);
nor U1941 (N_1941,N_1775,N_1610);
nand U1942 (N_1942,N_1605,N_1673);
nand U1943 (N_1943,N_1756,N_1621);
nand U1944 (N_1944,N_1627,N_1778);
or U1945 (N_1945,N_1680,N_1771);
and U1946 (N_1946,N_1765,N_1749);
nor U1947 (N_1947,N_1631,N_1775);
nor U1948 (N_1948,N_1725,N_1713);
nand U1949 (N_1949,N_1785,N_1688);
nand U1950 (N_1950,N_1690,N_1770);
and U1951 (N_1951,N_1676,N_1756);
and U1952 (N_1952,N_1650,N_1619);
nand U1953 (N_1953,N_1690,N_1673);
xor U1954 (N_1954,N_1703,N_1728);
nor U1955 (N_1955,N_1766,N_1669);
or U1956 (N_1956,N_1752,N_1696);
nand U1957 (N_1957,N_1617,N_1770);
xor U1958 (N_1958,N_1784,N_1648);
xor U1959 (N_1959,N_1688,N_1746);
xnor U1960 (N_1960,N_1788,N_1600);
or U1961 (N_1961,N_1618,N_1666);
and U1962 (N_1962,N_1666,N_1611);
xor U1963 (N_1963,N_1685,N_1627);
nor U1964 (N_1964,N_1705,N_1782);
xnor U1965 (N_1965,N_1731,N_1674);
xor U1966 (N_1966,N_1685,N_1622);
xnor U1967 (N_1967,N_1645,N_1795);
nand U1968 (N_1968,N_1680,N_1713);
nor U1969 (N_1969,N_1673,N_1642);
nor U1970 (N_1970,N_1608,N_1756);
nor U1971 (N_1971,N_1612,N_1787);
xor U1972 (N_1972,N_1655,N_1645);
and U1973 (N_1973,N_1650,N_1759);
nor U1974 (N_1974,N_1650,N_1798);
xor U1975 (N_1975,N_1730,N_1648);
xnor U1976 (N_1976,N_1765,N_1794);
xor U1977 (N_1977,N_1653,N_1629);
nor U1978 (N_1978,N_1719,N_1664);
nor U1979 (N_1979,N_1648,N_1772);
and U1980 (N_1980,N_1647,N_1724);
xor U1981 (N_1981,N_1702,N_1713);
nor U1982 (N_1982,N_1606,N_1788);
nor U1983 (N_1983,N_1735,N_1740);
or U1984 (N_1984,N_1733,N_1729);
nand U1985 (N_1985,N_1792,N_1618);
or U1986 (N_1986,N_1684,N_1731);
and U1987 (N_1987,N_1776,N_1626);
or U1988 (N_1988,N_1649,N_1782);
nand U1989 (N_1989,N_1647,N_1624);
nand U1990 (N_1990,N_1694,N_1677);
xor U1991 (N_1991,N_1751,N_1673);
xnor U1992 (N_1992,N_1626,N_1772);
or U1993 (N_1993,N_1737,N_1675);
xor U1994 (N_1994,N_1696,N_1756);
xnor U1995 (N_1995,N_1775,N_1693);
and U1996 (N_1996,N_1635,N_1737);
or U1997 (N_1997,N_1671,N_1702);
and U1998 (N_1998,N_1673,N_1740);
and U1999 (N_1999,N_1701,N_1659);
xnor U2000 (N_2000,N_1980,N_1901);
xnor U2001 (N_2001,N_1930,N_1881);
xor U2002 (N_2002,N_1906,N_1806);
and U2003 (N_2003,N_1941,N_1863);
nor U2004 (N_2004,N_1955,N_1878);
and U2005 (N_2005,N_1846,N_1935);
or U2006 (N_2006,N_1999,N_1943);
nor U2007 (N_2007,N_1920,N_1956);
nor U2008 (N_2008,N_1982,N_1889);
nand U2009 (N_2009,N_1815,N_1986);
nor U2010 (N_2010,N_1812,N_1991);
nand U2011 (N_2011,N_1963,N_1954);
nand U2012 (N_2012,N_1953,N_1841);
and U2013 (N_2013,N_1844,N_1974);
nor U2014 (N_2014,N_1870,N_1938);
nand U2015 (N_2015,N_1854,N_1940);
nand U2016 (N_2016,N_1979,N_1874);
nor U2017 (N_2017,N_1958,N_1823);
nor U2018 (N_2018,N_1957,N_1811);
and U2019 (N_2019,N_1871,N_1971);
or U2020 (N_2020,N_1989,N_1837);
nor U2021 (N_2021,N_1879,N_1966);
nor U2022 (N_2022,N_1895,N_1990);
nor U2023 (N_2023,N_1910,N_1832);
and U2024 (N_2024,N_1808,N_1807);
or U2025 (N_2025,N_1978,N_1964);
nand U2026 (N_2026,N_1973,N_1861);
or U2027 (N_2027,N_1976,N_1907);
nand U2028 (N_2028,N_1801,N_1876);
or U2029 (N_2029,N_1865,N_1884);
nor U2030 (N_2030,N_1872,N_1850);
nand U2031 (N_2031,N_1947,N_1987);
and U2032 (N_2032,N_1800,N_1908);
nand U2033 (N_2033,N_1857,N_1917);
and U2034 (N_2034,N_1927,N_1993);
nor U2035 (N_2035,N_1899,N_1968);
xor U2036 (N_2036,N_1926,N_1890);
and U2037 (N_2037,N_1931,N_1869);
or U2038 (N_2038,N_1802,N_1977);
nor U2039 (N_2039,N_1952,N_1833);
and U2040 (N_2040,N_1834,N_1849);
or U2041 (N_2041,N_1921,N_1919);
or U2042 (N_2042,N_1824,N_1996);
nand U2043 (N_2043,N_1803,N_1859);
and U2044 (N_2044,N_1992,N_1894);
xor U2045 (N_2045,N_1867,N_1972);
nor U2046 (N_2046,N_1825,N_1836);
and U2047 (N_2047,N_1818,N_1918);
nand U2048 (N_2048,N_1961,N_1914);
nand U2049 (N_2049,N_1924,N_1985);
or U2050 (N_2050,N_1860,N_1877);
and U2051 (N_2051,N_1840,N_1932);
nor U2052 (N_2052,N_1885,N_1853);
nor U2053 (N_2053,N_1928,N_1967);
nor U2054 (N_2054,N_1903,N_1862);
nor U2055 (N_2055,N_1835,N_1909);
nand U2056 (N_2056,N_1898,N_1913);
xnor U2057 (N_2057,N_1923,N_1880);
and U2058 (N_2058,N_1933,N_1905);
nand U2059 (N_2059,N_1827,N_1998);
or U2060 (N_2060,N_1962,N_1892);
nor U2061 (N_2061,N_1843,N_1883);
or U2062 (N_2062,N_1951,N_1830);
or U2063 (N_2063,N_1934,N_1822);
or U2064 (N_2064,N_1842,N_1904);
nor U2065 (N_2065,N_1916,N_1944);
or U2066 (N_2066,N_1831,N_1929);
or U2067 (N_2067,N_1851,N_1886);
nor U2068 (N_2068,N_1981,N_1997);
xnor U2069 (N_2069,N_1939,N_1839);
xnor U2070 (N_2070,N_1847,N_1949);
nand U2071 (N_2071,N_1922,N_1821);
or U2072 (N_2072,N_1950,N_1925);
nor U2073 (N_2073,N_1994,N_1809);
and U2074 (N_2074,N_1845,N_1817);
nand U2075 (N_2075,N_1866,N_1893);
and U2076 (N_2076,N_1826,N_1942);
or U2077 (N_2077,N_1975,N_1902);
nor U2078 (N_2078,N_1984,N_1810);
nor U2079 (N_2079,N_1887,N_1896);
or U2080 (N_2080,N_1988,N_1816);
or U2081 (N_2081,N_1858,N_1970);
xor U2082 (N_2082,N_1969,N_1873);
xor U2083 (N_2083,N_1864,N_1915);
xnor U2084 (N_2084,N_1888,N_1882);
nand U2085 (N_2085,N_1855,N_1848);
or U2086 (N_2086,N_1805,N_1937);
and U2087 (N_2087,N_1960,N_1936);
nand U2088 (N_2088,N_1852,N_1983);
xnor U2089 (N_2089,N_1911,N_1868);
or U2090 (N_2090,N_1829,N_1959);
and U2091 (N_2091,N_1804,N_1813);
nor U2092 (N_2092,N_1891,N_1820);
nand U2093 (N_2093,N_1828,N_1838);
nand U2094 (N_2094,N_1945,N_1965);
nor U2095 (N_2095,N_1900,N_1946);
nand U2096 (N_2096,N_1814,N_1819);
xor U2097 (N_2097,N_1948,N_1875);
or U2098 (N_2098,N_1856,N_1995);
nor U2099 (N_2099,N_1912,N_1897);
nor U2100 (N_2100,N_1906,N_1960);
or U2101 (N_2101,N_1953,N_1910);
nor U2102 (N_2102,N_1919,N_1948);
nand U2103 (N_2103,N_1932,N_1910);
nand U2104 (N_2104,N_1958,N_1972);
nand U2105 (N_2105,N_1934,N_1843);
nor U2106 (N_2106,N_1851,N_1997);
nor U2107 (N_2107,N_1985,N_1806);
xor U2108 (N_2108,N_1926,N_1892);
and U2109 (N_2109,N_1855,N_1912);
nor U2110 (N_2110,N_1973,N_1845);
or U2111 (N_2111,N_1950,N_1853);
nor U2112 (N_2112,N_1876,N_1817);
and U2113 (N_2113,N_1918,N_1993);
or U2114 (N_2114,N_1929,N_1813);
or U2115 (N_2115,N_1956,N_1918);
nand U2116 (N_2116,N_1873,N_1835);
or U2117 (N_2117,N_1947,N_1925);
xor U2118 (N_2118,N_1823,N_1860);
and U2119 (N_2119,N_1958,N_1998);
nand U2120 (N_2120,N_1927,N_1810);
nand U2121 (N_2121,N_1953,N_1913);
or U2122 (N_2122,N_1953,N_1808);
nand U2123 (N_2123,N_1885,N_1845);
or U2124 (N_2124,N_1841,N_1852);
and U2125 (N_2125,N_1831,N_1971);
nor U2126 (N_2126,N_1811,N_1950);
nand U2127 (N_2127,N_1911,N_1999);
xnor U2128 (N_2128,N_1810,N_1968);
nand U2129 (N_2129,N_1991,N_1971);
nor U2130 (N_2130,N_1874,N_1940);
xor U2131 (N_2131,N_1954,N_1829);
and U2132 (N_2132,N_1905,N_1848);
nor U2133 (N_2133,N_1903,N_1870);
xor U2134 (N_2134,N_1881,N_1934);
xor U2135 (N_2135,N_1877,N_1807);
nor U2136 (N_2136,N_1969,N_1974);
or U2137 (N_2137,N_1974,N_1909);
and U2138 (N_2138,N_1810,N_1941);
and U2139 (N_2139,N_1846,N_1877);
and U2140 (N_2140,N_1966,N_1907);
nand U2141 (N_2141,N_1972,N_1804);
nand U2142 (N_2142,N_1857,N_1956);
or U2143 (N_2143,N_1940,N_1867);
and U2144 (N_2144,N_1875,N_1946);
or U2145 (N_2145,N_1987,N_1998);
and U2146 (N_2146,N_1938,N_1923);
or U2147 (N_2147,N_1841,N_1981);
and U2148 (N_2148,N_1808,N_1913);
or U2149 (N_2149,N_1827,N_1958);
and U2150 (N_2150,N_1930,N_1942);
nor U2151 (N_2151,N_1918,N_1991);
xor U2152 (N_2152,N_1931,N_1920);
or U2153 (N_2153,N_1850,N_1975);
or U2154 (N_2154,N_1809,N_1986);
nor U2155 (N_2155,N_1928,N_1997);
nor U2156 (N_2156,N_1871,N_1852);
or U2157 (N_2157,N_1859,N_1990);
and U2158 (N_2158,N_1895,N_1837);
nor U2159 (N_2159,N_1802,N_1980);
xnor U2160 (N_2160,N_1960,N_1860);
xnor U2161 (N_2161,N_1924,N_1809);
or U2162 (N_2162,N_1874,N_1869);
nand U2163 (N_2163,N_1856,N_1913);
nand U2164 (N_2164,N_1980,N_1924);
nor U2165 (N_2165,N_1806,N_1831);
xor U2166 (N_2166,N_1932,N_1936);
nor U2167 (N_2167,N_1817,N_1800);
xnor U2168 (N_2168,N_1840,N_1969);
nand U2169 (N_2169,N_1897,N_1922);
nor U2170 (N_2170,N_1993,N_1921);
nand U2171 (N_2171,N_1804,N_1978);
nor U2172 (N_2172,N_1918,N_1871);
nand U2173 (N_2173,N_1889,N_1916);
and U2174 (N_2174,N_1994,N_1895);
xnor U2175 (N_2175,N_1851,N_1805);
or U2176 (N_2176,N_1817,N_1840);
or U2177 (N_2177,N_1985,N_1934);
xnor U2178 (N_2178,N_1948,N_1857);
nor U2179 (N_2179,N_1826,N_1852);
or U2180 (N_2180,N_1974,N_1845);
or U2181 (N_2181,N_1841,N_1932);
nor U2182 (N_2182,N_1933,N_1957);
nand U2183 (N_2183,N_1935,N_1866);
and U2184 (N_2184,N_1941,N_1948);
xor U2185 (N_2185,N_1878,N_1836);
or U2186 (N_2186,N_1968,N_1977);
or U2187 (N_2187,N_1845,N_1910);
and U2188 (N_2188,N_1899,N_1853);
nand U2189 (N_2189,N_1911,N_1806);
and U2190 (N_2190,N_1971,N_1929);
or U2191 (N_2191,N_1998,N_1817);
nand U2192 (N_2192,N_1887,N_1914);
nor U2193 (N_2193,N_1895,N_1929);
xor U2194 (N_2194,N_1828,N_1946);
xnor U2195 (N_2195,N_1969,N_1806);
or U2196 (N_2196,N_1926,N_1827);
nand U2197 (N_2197,N_1882,N_1954);
or U2198 (N_2198,N_1852,N_1811);
nand U2199 (N_2199,N_1993,N_1889);
xor U2200 (N_2200,N_2110,N_2172);
nor U2201 (N_2201,N_2116,N_2169);
nand U2202 (N_2202,N_2179,N_2111);
xnor U2203 (N_2203,N_2056,N_2166);
nor U2204 (N_2204,N_2152,N_2019);
nand U2205 (N_2205,N_2188,N_2085);
nor U2206 (N_2206,N_2144,N_2108);
and U2207 (N_2207,N_2138,N_2105);
xor U2208 (N_2208,N_2196,N_2071);
or U2209 (N_2209,N_2027,N_2190);
nand U2210 (N_2210,N_2078,N_2147);
and U2211 (N_2211,N_2069,N_2174);
nand U2212 (N_2212,N_2070,N_2009);
xor U2213 (N_2213,N_2053,N_2163);
and U2214 (N_2214,N_2058,N_2016);
and U2215 (N_2215,N_2049,N_2041);
nor U2216 (N_2216,N_2162,N_2185);
nand U2217 (N_2217,N_2164,N_2018);
or U2218 (N_2218,N_2098,N_2124);
xor U2219 (N_2219,N_2060,N_2126);
xnor U2220 (N_2220,N_2125,N_2195);
xnor U2221 (N_2221,N_2052,N_2021);
xor U2222 (N_2222,N_2134,N_2079);
or U2223 (N_2223,N_2097,N_2023);
nand U2224 (N_2224,N_2064,N_2033);
and U2225 (N_2225,N_2047,N_2072);
xor U2226 (N_2226,N_2150,N_2132);
or U2227 (N_2227,N_2136,N_2106);
or U2228 (N_2228,N_2039,N_2182);
or U2229 (N_2229,N_2165,N_2030);
and U2230 (N_2230,N_2008,N_2156);
nor U2231 (N_2231,N_2117,N_2092);
xnor U2232 (N_2232,N_2113,N_2029);
nor U2233 (N_2233,N_2006,N_2084);
nor U2234 (N_2234,N_2095,N_2109);
nand U2235 (N_2235,N_2044,N_2123);
and U2236 (N_2236,N_2114,N_2187);
or U2237 (N_2237,N_2131,N_2103);
and U2238 (N_2238,N_2067,N_2139);
or U2239 (N_2239,N_2112,N_2192);
or U2240 (N_2240,N_2082,N_2051);
nand U2241 (N_2241,N_2014,N_2062);
nand U2242 (N_2242,N_2099,N_2080);
nor U2243 (N_2243,N_2007,N_2042);
and U2244 (N_2244,N_2118,N_2028);
nor U2245 (N_2245,N_2149,N_2170);
and U2246 (N_2246,N_2040,N_2083);
and U2247 (N_2247,N_2148,N_2004);
xor U2248 (N_2248,N_2005,N_2096);
and U2249 (N_2249,N_2199,N_2075);
and U2250 (N_2250,N_2153,N_2177);
and U2251 (N_2251,N_2000,N_2063);
nand U2252 (N_2252,N_2141,N_2151);
xnor U2253 (N_2253,N_2121,N_2173);
nand U2254 (N_2254,N_2193,N_2038);
or U2255 (N_2255,N_2159,N_2130);
nor U2256 (N_2256,N_2128,N_2100);
xnor U2257 (N_2257,N_2020,N_2076);
or U2258 (N_2258,N_2175,N_2065);
nor U2259 (N_2259,N_2054,N_2093);
nand U2260 (N_2260,N_2102,N_2012);
nand U2261 (N_2261,N_2154,N_2167);
and U2262 (N_2262,N_2145,N_2013);
or U2263 (N_2263,N_2101,N_2010);
or U2264 (N_2264,N_2186,N_2129);
xor U2265 (N_2265,N_2094,N_2168);
nand U2266 (N_2266,N_2183,N_2017);
or U2267 (N_2267,N_2061,N_2036);
nand U2268 (N_2268,N_2035,N_2180);
or U2269 (N_2269,N_2157,N_2155);
nor U2270 (N_2270,N_2178,N_2050);
or U2271 (N_2271,N_2088,N_2087);
xnor U2272 (N_2272,N_2073,N_2001);
nor U2273 (N_2273,N_2043,N_2197);
or U2274 (N_2274,N_2086,N_2057);
nand U2275 (N_2275,N_2081,N_2025);
xnor U2276 (N_2276,N_2037,N_2107);
nor U2277 (N_2277,N_2055,N_2122);
and U2278 (N_2278,N_2135,N_2158);
nand U2279 (N_2279,N_2003,N_2189);
or U2280 (N_2280,N_2104,N_2059);
xnor U2281 (N_2281,N_2160,N_2045);
xor U2282 (N_2282,N_2133,N_2022);
nor U2283 (N_2283,N_2194,N_2191);
nand U2284 (N_2284,N_2140,N_2026);
or U2285 (N_2285,N_2142,N_2143);
or U2286 (N_2286,N_2066,N_2015);
xnor U2287 (N_2287,N_2046,N_2048);
and U2288 (N_2288,N_2198,N_2068);
nand U2289 (N_2289,N_2032,N_2031);
nand U2290 (N_2290,N_2137,N_2024);
or U2291 (N_2291,N_2171,N_2091);
nor U2292 (N_2292,N_2089,N_2090);
and U2293 (N_2293,N_2161,N_2002);
and U2294 (N_2294,N_2146,N_2120);
or U2295 (N_2295,N_2127,N_2074);
nor U2296 (N_2296,N_2011,N_2034);
nor U2297 (N_2297,N_2119,N_2077);
and U2298 (N_2298,N_2176,N_2115);
xnor U2299 (N_2299,N_2184,N_2181);
or U2300 (N_2300,N_2193,N_2008);
xnor U2301 (N_2301,N_2052,N_2136);
or U2302 (N_2302,N_2152,N_2085);
nor U2303 (N_2303,N_2165,N_2180);
nand U2304 (N_2304,N_2097,N_2190);
xor U2305 (N_2305,N_2174,N_2188);
nand U2306 (N_2306,N_2042,N_2064);
nor U2307 (N_2307,N_2014,N_2164);
and U2308 (N_2308,N_2126,N_2074);
nand U2309 (N_2309,N_2129,N_2021);
nor U2310 (N_2310,N_2135,N_2103);
or U2311 (N_2311,N_2001,N_2048);
xnor U2312 (N_2312,N_2078,N_2094);
nand U2313 (N_2313,N_2190,N_2070);
or U2314 (N_2314,N_2046,N_2040);
nor U2315 (N_2315,N_2083,N_2014);
nor U2316 (N_2316,N_2058,N_2093);
and U2317 (N_2317,N_2064,N_2131);
xnor U2318 (N_2318,N_2070,N_2194);
xor U2319 (N_2319,N_2079,N_2025);
or U2320 (N_2320,N_2114,N_2048);
xnor U2321 (N_2321,N_2163,N_2083);
or U2322 (N_2322,N_2137,N_2051);
xnor U2323 (N_2323,N_2142,N_2195);
xor U2324 (N_2324,N_2002,N_2170);
nor U2325 (N_2325,N_2076,N_2048);
nand U2326 (N_2326,N_2119,N_2161);
or U2327 (N_2327,N_2011,N_2125);
or U2328 (N_2328,N_2035,N_2123);
and U2329 (N_2329,N_2056,N_2069);
and U2330 (N_2330,N_2043,N_2112);
and U2331 (N_2331,N_2077,N_2127);
nor U2332 (N_2332,N_2047,N_2070);
xor U2333 (N_2333,N_2129,N_2190);
xnor U2334 (N_2334,N_2165,N_2021);
nand U2335 (N_2335,N_2116,N_2096);
xnor U2336 (N_2336,N_2176,N_2016);
xnor U2337 (N_2337,N_2177,N_2012);
nand U2338 (N_2338,N_2049,N_2031);
and U2339 (N_2339,N_2098,N_2040);
or U2340 (N_2340,N_2103,N_2077);
or U2341 (N_2341,N_2153,N_2159);
nor U2342 (N_2342,N_2103,N_2044);
xor U2343 (N_2343,N_2118,N_2199);
nand U2344 (N_2344,N_2039,N_2018);
nand U2345 (N_2345,N_2128,N_2027);
xnor U2346 (N_2346,N_2154,N_2001);
nor U2347 (N_2347,N_2081,N_2154);
nand U2348 (N_2348,N_2003,N_2052);
xor U2349 (N_2349,N_2136,N_2123);
nand U2350 (N_2350,N_2020,N_2000);
nand U2351 (N_2351,N_2151,N_2196);
nand U2352 (N_2352,N_2120,N_2016);
nor U2353 (N_2353,N_2196,N_2029);
nand U2354 (N_2354,N_2167,N_2176);
nor U2355 (N_2355,N_2070,N_2046);
xnor U2356 (N_2356,N_2134,N_2004);
nand U2357 (N_2357,N_2174,N_2097);
or U2358 (N_2358,N_2160,N_2129);
and U2359 (N_2359,N_2076,N_2127);
or U2360 (N_2360,N_2101,N_2061);
nand U2361 (N_2361,N_2070,N_2163);
and U2362 (N_2362,N_2068,N_2142);
xor U2363 (N_2363,N_2091,N_2051);
or U2364 (N_2364,N_2185,N_2056);
xnor U2365 (N_2365,N_2188,N_2064);
or U2366 (N_2366,N_2050,N_2193);
or U2367 (N_2367,N_2106,N_2096);
nor U2368 (N_2368,N_2173,N_2048);
nor U2369 (N_2369,N_2101,N_2175);
nor U2370 (N_2370,N_2115,N_2031);
and U2371 (N_2371,N_2078,N_2124);
nor U2372 (N_2372,N_2164,N_2126);
xor U2373 (N_2373,N_2173,N_2092);
or U2374 (N_2374,N_2047,N_2042);
nor U2375 (N_2375,N_2169,N_2161);
or U2376 (N_2376,N_2179,N_2148);
and U2377 (N_2377,N_2074,N_2034);
nor U2378 (N_2378,N_2100,N_2155);
xnor U2379 (N_2379,N_2141,N_2037);
or U2380 (N_2380,N_2171,N_2048);
or U2381 (N_2381,N_2012,N_2001);
and U2382 (N_2382,N_2138,N_2167);
nand U2383 (N_2383,N_2042,N_2170);
xor U2384 (N_2384,N_2089,N_2114);
nor U2385 (N_2385,N_2160,N_2094);
nand U2386 (N_2386,N_2140,N_2178);
nor U2387 (N_2387,N_2043,N_2005);
and U2388 (N_2388,N_2100,N_2042);
nor U2389 (N_2389,N_2182,N_2151);
or U2390 (N_2390,N_2041,N_2003);
nor U2391 (N_2391,N_2138,N_2034);
xor U2392 (N_2392,N_2032,N_2052);
xor U2393 (N_2393,N_2173,N_2106);
xnor U2394 (N_2394,N_2005,N_2155);
xnor U2395 (N_2395,N_2184,N_2022);
nor U2396 (N_2396,N_2178,N_2126);
or U2397 (N_2397,N_2035,N_2058);
or U2398 (N_2398,N_2072,N_2025);
nand U2399 (N_2399,N_2163,N_2094);
xor U2400 (N_2400,N_2289,N_2212);
xnor U2401 (N_2401,N_2380,N_2230);
and U2402 (N_2402,N_2321,N_2329);
and U2403 (N_2403,N_2214,N_2353);
and U2404 (N_2404,N_2290,N_2254);
nor U2405 (N_2405,N_2315,N_2285);
xor U2406 (N_2406,N_2213,N_2222);
nand U2407 (N_2407,N_2372,N_2236);
nand U2408 (N_2408,N_2203,N_2271);
nand U2409 (N_2409,N_2324,N_2238);
nand U2410 (N_2410,N_2202,N_2361);
and U2411 (N_2411,N_2211,N_2266);
nor U2412 (N_2412,N_2355,N_2338);
or U2413 (N_2413,N_2277,N_2249);
or U2414 (N_2414,N_2345,N_2358);
and U2415 (N_2415,N_2336,N_2375);
or U2416 (N_2416,N_2239,N_2330);
nor U2417 (N_2417,N_2267,N_2326);
nand U2418 (N_2418,N_2245,N_2346);
nor U2419 (N_2419,N_2291,N_2250);
and U2420 (N_2420,N_2357,N_2246);
or U2421 (N_2421,N_2244,N_2260);
xor U2422 (N_2422,N_2282,N_2354);
xor U2423 (N_2423,N_2365,N_2226);
or U2424 (N_2424,N_2343,N_2264);
and U2425 (N_2425,N_2297,N_2397);
nand U2426 (N_2426,N_2287,N_2347);
xor U2427 (N_2427,N_2229,N_2310);
and U2428 (N_2428,N_2320,N_2257);
xor U2429 (N_2429,N_2322,N_2369);
nor U2430 (N_2430,N_2387,N_2356);
or U2431 (N_2431,N_2327,N_2206);
or U2432 (N_2432,N_2348,N_2296);
xor U2433 (N_2433,N_2390,N_2304);
and U2434 (N_2434,N_2272,N_2314);
nor U2435 (N_2435,N_2234,N_2233);
and U2436 (N_2436,N_2363,N_2335);
xnor U2437 (N_2437,N_2374,N_2333);
xnor U2438 (N_2438,N_2395,N_2303);
or U2439 (N_2439,N_2224,N_2216);
and U2440 (N_2440,N_2286,N_2370);
or U2441 (N_2441,N_2298,N_2378);
or U2442 (N_2442,N_2283,N_2237);
or U2443 (N_2443,N_2388,N_2399);
nand U2444 (N_2444,N_2377,N_2259);
and U2445 (N_2445,N_2342,N_2398);
and U2446 (N_2446,N_2302,N_2367);
or U2447 (N_2447,N_2208,N_2268);
xor U2448 (N_2448,N_2219,N_2349);
xnor U2449 (N_2449,N_2243,N_2337);
and U2450 (N_2450,N_2306,N_2325);
nor U2451 (N_2451,N_2209,N_2385);
xor U2452 (N_2452,N_2247,N_2223);
nor U2453 (N_2453,N_2341,N_2352);
nand U2454 (N_2454,N_2318,N_2396);
or U2455 (N_2455,N_2201,N_2328);
xnor U2456 (N_2456,N_2274,N_2218);
nor U2457 (N_2457,N_2275,N_2340);
nor U2458 (N_2458,N_2235,N_2221);
and U2459 (N_2459,N_2384,N_2232);
nand U2460 (N_2460,N_2359,N_2200);
nand U2461 (N_2461,N_2261,N_2255);
or U2462 (N_2462,N_2292,N_2299);
and U2463 (N_2463,N_2251,N_2263);
xnor U2464 (N_2464,N_2293,N_2210);
nand U2465 (N_2465,N_2205,N_2204);
or U2466 (N_2466,N_2227,N_2301);
nor U2467 (N_2467,N_2316,N_2373);
nor U2468 (N_2468,N_2344,N_2256);
nand U2469 (N_2469,N_2313,N_2331);
xnor U2470 (N_2470,N_2265,N_2288);
nor U2471 (N_2471,N_2312,N_2295);
or U2472 (N_2472,N_2383,N_2269);
and U2473 (N_2473,N_2394,N_2240);
or U2474 (N_2474,N_2280,N_2225);
nand U2475 (N_2475,N_2248,N_2332);
or U2476 (N_2476,N_2284,N_2381);
or U2477 (N_2477,N_2317,N_2270);
and U2478 (N_2478,N_2339,N_2351);
nor U2479 (N_2479,N_2308,N_2276);
and U2480 (N_2480,N_2262,N_2220);
or U2481 (N_2481,N_2207,N_2391);
xnor U2482 (N_2482,N_2215,N_2311);
and U2483 (N_2483,N_2379,N_2376);
nand U2484 (N_2484,N_2334,N_2371);
nand U2485 (N_2485,N_2393,N_2253);
xnor U2486 (N_2486,N_2392,N_2319);
nand U2487 (N_2487,N_2307,N_2389);
nor U2488 (N_2488,N_2273,N_2386);
xnor U2489 (N_2489,N_2309,N_2382);
and U2490 (N_2490,N_2300,N_2252);
and U2491 (N_2491,N_2323,N_2360);
nand U2492 (N_2492,N_2228,N_2258);
nand U2493 (N_2493,N_2305,N_2241);
nor U2494 (N_2494,N_2278,N_2281);
nor U2495 (N_2495,N_2366,N_2294);
or U2496 (N_2496,N_2362,N_2242);
or U2497 (N_2497,N_2368,N_2364);
xnor U2498 (N_2498,N_2350,N_2279);
nand U2499 (N_2499,N_2231,N_2217);
nand U2500 (N_2500,N_2363,N_2398);
or U2501 (N_2501,N_2348,N_2379);
nand U2502 (N_2502,N_2270,N_2210);
nor U2503 (N_2503,N_2248,N_2245);
and U2504 (N_2504,N_2210,N_2221);
nand U2505 (N_2505,N_2359,N_2362);
xor U2506 (N_2506,N_2249,N_2341);
or U2507 (N_2507,N_2337,N_2240);
or U2508 (N_2508,N_2279,N_2329);
xor U2509 (N_2509,N_2259,N_2242);
xor U2510 (N_2510,N_2307,N_2285);
xnor U2511 (N_2511,N_2269,N_2237);
xor U2512 (N_2512,N_2317,N_2211);
nand U2513 (N_2513,N_2249,N_2345);
or U2514 (N_2514,N_2238,N_2355);
nor U2515 (N_2515,N_2344,N_2386);
xnor U2516 (N_2516,N_2350,N_2272);
or U2517 (N_2517,N_2246,N_2324);
nand U2518 (N_2518,N_2326,N_2312);
nand U2519 (N_2519,N_2307,N_2315);
xor U2520 (N_2520,N_2378,N_2269);
xnor U2521 (N_2521,N_2385,N_2288);
nor U2522 (N_2522,N_2284,N_2364);
or U2523 (N_2523,N_2304,N_2318);
and U2524 (N_2524,N_2212,N_2318);
nor U2525 (N_2525,N_2318,N_2328);
or U2526 (N_2526,N_2220,N_2243);
xnor U2527 (N_2527,N_2331,N_2343);
nor U2528 (N_2528,N_2217,N_2308);
and U2529 (N_2529,N_2362,N_2215);
and U2530 (N_2530,N_2347,N_2235);
or U2531 (N_2531,N_2219,N_2251);
nor U2532 (N_2532,N_2273,N_2321);
or U2533 (N_2533,N_2252,N_2353);
nor U2534 (N_2534,N_2366,N_2339);
and U2535 (N_2535,N_2318,N_2374);
xor U2536 (N_2536,N_2245,N_2220);
and U2537 (N_2537,N_2286,N_2202);
xnor U2538 (N_2538,N_2311,N_2272);
nor U2539 (N_2539,N_2352,N_2335);
xor U2540 (N_2540,N_2303,N_2351);
or U2541 (N_2541,N_2239,N_2254);
xnor U2542 (N_2542,N_2250,N_2322);
nand U2543 (N_2543,N_2242,N_2207);
and U2544 (N_2544,N_2208,N_2356);
nand U2545 (N_2545,N_2346,N_2209);
nor U2546 (N_2546,N_2325,N_2230);
and U2547 (N_2547,N_2308,N_2287);
xor U2548 (N_2548,N_2248,N_2255);
xor U2549 (N_2549,N_2262,N_2304);
or U2550 (N_2550,N_2224,N_2312);
nand U2551 (N_2551,N_2241,N_2319);
xor U2552 (N_2552,N_2238,N_2389);
nor U2553 (N_2553,N_2216,N_2296);
or U2554 (N_2554,N_2219,N_2335);
and U2555 (N_2555,N_2335,N_2337);
nor U2556 (N_2556,N_2201,N_2232);
nor U2557 (N_2557,N_2343,N_2200);
or U2558 (N_2558,N_2358,N_2262);
nand U2559 (N_2559,N_2204,N_2224);
and U2560 (N_2560,N_2320,N_2345);
nand U2561 (N_2561,N_2363,N_2255);
nor U2562 (N_2562,N_2342,N_2317);
xor U2563 (N_2563,N_2255,N_2399);
nand U2564 (N_2564,N_2230,N_2283);
or U2565 (N_2565,N_2265,N_2327);
xnor U2566 (N_2566,N_2395,N_2293);
and U2567 (N_2567,N_2238,N_2348);
xnor U2568 (N_2568,N_2201,N_2353);
and U2569 (N_2569,N_2394,N_2297);
and U2570 (N_2570,N_2227,N_2376);
nand U2571 (N_2571,N_2265,N_2273);
nand U2572 (N_2572,N_2241,N_2310);
or U2573 (N_2573,N_2353,N_2259);
or U2574 (N_2574,N_2209,N_2338);
or U2575 (N_2575,N_2393,N_2243);
or U2576 (N_2576,N_2376,N_2205);
and U2577 (N_2577,N_2269,N_2262);
nor U2578 (N_2578,N_2238,N_2266);
nand U2579 (N_2579,N_2269,N_2204);
xnor U2580 (N_2580,N_2354,N_2209);
nor U2581 (N_2581,N_2207,N_2368);
nor U2582 (N_2582,N_2253,N_2250);
or U2583 (N_2583,N_2350,N_2231);
or U2584 (N_2584,N_2232,N_2364);
or U2585 (N_2585,N_2344,N_2228);
nor U2586 (N_2586,N_2393,N_2201);
or U2587 (N_2587,N_2276,N_2275);
nor U2588 (N_2588,N_2206,N_2205);
nand U2589 (N_2589,N_2246,N_2369);
and U2590 (N_2590,N_2210,N_2334);
or U2591 (N_2591,N_2328,N_2233);
and U2592 (N_2592,N_2365,N_2324);
nand U2593 (N_2593,N_2352,N_2302);
nor U2594 (N_2594,N_2246,N_2223);
or U2595 (N_2595,N_2202,N_2222);
and U2596 (N_2596,N_2248,N_2228);
nand U2597 (N_2597,N_2259,N_2306);
nand U2598 (N_2598,N_2349,N_2252);
or U2599 (N_2599,N_2299,N_2242);
nor U2600 (N_2600,N_2505,N_2454);
nor U2601 (N_2601,N_2567,N_2522);
xor U2602 (N_2602,N_2450,N_2595);
or U2603 (N_2603,N_2401,N_2512);
nand U2604 (N_2604,N_2417,N_2467);
or U2605 (N_2605,N_2459,N_2564);
nand U2606 (N_2606,N_2566,N_2481);
nand U2607 (N_2607,N_2476,N_2406);
nor U2608 (N_2608,N_2561,N_2463);
nor U2609 (N_2609,N_2432,N_2426);
nand U2610 (N_2610,N_2445,N_2488);
and U2611 (N_2611,N_2557,N_2420);
nand U2612 (N_2612,N_2437,N_2591);
nor U2613 (N_2613,N_2455,N_2461);
nor U2614 (N_2614,N_2542,N_2535);
and U2615 (N_2615,N_2416,N_2465);
nor U2616 (N_2616,N_2599,N_2438);
xor U2617 (N_2617,N_2515,N_2593);
nor U2618 (N_2618,N_2530,N_2583);
xnor U2619 (N_2619,N_2543,N_2533);
nor U2620 (N_2620,N_2596,N_2453);
nor U2621 (N_2621,N_2590,N_2474);
and U2622 (N_2622,N_2485,N_2460);
and U2623 (N_2623,N_2419,N_2525);
or U2624 (N_2624,N_2569,N_2477);
xnor U2625 (N_2625,N_2410,N_2486);
xnor U2626 (N_2626,N_2579,N_2422);
xnor U2627 (N_2627,N_2504,N_2584);
nand U2628 (N_2628,N_2578,N_2544);
nand U2629 (N_2629,N_2571,N_2430);
nor U2630 (N_2630,N_2497,N_2421);
and U2631 (N_2631,N_2527,N_2451);
nand U2632 (N_2632,N_2570,N_2506);
nand U2633 (N_2633,N_2447,N_2491);
and U2634 (N_2634,N_2439,N_2499);
and U2635 (N_2635,N_2409,N_2514);
and U2636 (N_2636,N_2517,N_2449);
and U2637 (N_2637,N_2518,N_2553);
xnor U2638 (N_2638,N_2594,N_2452);
xnor U2639 (N_2639,N_2494,N_2493);
and U2640 (N_2640,N_2427,N_2457);
nand U2641 (N_2641,N_2425,N_2592);
and U2642 (N_2642,N_2540,N_2536);
nand U2643 (N_2643,N_2479,N_2573);
nand U2644 (N_2644,N_2577,N_2532);
nand U2645 (N_2645,N_2576,N_2586);
or U2646 (N_2646,N_2433,N_2423);
nor U2647 (N_2647,N_2428,N_2496);
nand U2648 (N_2648,N_2434,N_2404);
nor U2649 (N_2649,N_2466,N_2547);
xor U2650 (N_2650,N_2513,N_2495);
xnor U2651 (N_2651,N_2511,N_2519);
or U2652 (N_2652,N_2526,N_2405);
or U2653 (N_2653,N_2501,N_2458);
or U2654 (N_2654,N_2407,N_2524);
and U2655 (N_2655,N_2550,N_2443);
nor U2656 (N_2656,N_2538,N_2444);
and U2657 (N_2657,N_2531,N_2554);
nor U2658 (N_2658,N_2468,N_2548);
xnor U2659 (N_2659,N_2555,N_2442);
nand U2660 (N_2660,N_2509,N_2503);
nand U2661 (N_2661,N_2559,N_2572);
nand U2662 (N_2662,N_2429,N_2478);
or U2663 (N_2663,N_2558,N_2541);
nor U2664 (N_2664,N_2470,N_2588);
nor U2665 (N_2665,N_2574,N_2539);
nand U2666 (N_2666,N_2487,N_2440);
nand U2667 (N_2667,N_2523,N_2563);
and U2668 (N_2668,N_2411,N_2402);
xor U2669 (N_2669,N_2471,N_2424);
nand U2670 (N_2670,N_2446,N_2472);
nor U2671 (N_2671,N_2545,N_2483);
xor U2672 (N_2672,N_2502,N_2489);
nor U2673 (N_2673,N_2598,N_2520);
xnor U2674 (N_2674,N_2562,N_2537);
or U2675 (N_2675,N_2510,N_2498);
xnor U2676 (N_2676,N_2435,N_2412);
and U2677 (N_2677,N_2415,N_2441);
xnor U2678 (N_2678,N_2534,N_2546);
or U2679 (N_2679,N_2462,N_2500);
or U2680 (N_2680,N_2551,N_2580);
and U2681 (N_2681,N_2581,N_2565);
nor U2682 (N_2682,N_2587,N_2431);
xnor U2683 (N_2683,N_2568,N_2589);
or U2684 (N_2684,N_2480,N_2484);
nand U2685 (N_2685,N_2597,N_2464);
or U2686 (N_2686,N_2490,N_2418);
and U2687 (N_2687,N_2414,N_2528);
or U2688 (N_2688,N_2400,N_2582);
or U2689 (N_2689,N_2507,N_2448);
nand U2690 (N_2690,N_2436,N_2482);
nand U2691 (N_2691,N_2475,N_2575);
nor U2692 (N_2692,N_2552,N_2529);
nor U2693 (N_2693,N_2549,N_2521);
nand U2694 (N_2694,N_2469,N_2473);
and U2695 (N_2695,N_2556,N_2408);
and U2696 (N_2696,N_2585,N_2413);
xnor U2697 (N_2697,N_2492,N_2456);
nor U2698 (N_2698,N_2508,N_2403);
xnor U2699 (N_2699,N_2516,N_2560);
nand U2700 (N_2700,N_2543,N_2439);
nor U2701 (N_2701,N_2408,N_2479);
nor U2702 (N_2702,N_2589,N_2565);
nor U2703 (N_2703,N_2466,N_2568);
and U2704 (N_2704,N_2402,N_2425);
and U2705 (N_2705,N_2498,N_2419);
or U2706 (N_2706,N_2418,N_2481);
and U2707 (N_2707,N_2516,N_2558);
nor U2708 (N_2708,N_2514,N_2574);
and U2709 (N_2709,N_2430,N_2569);
nor U2710 (N_2710,N_2538,N_2593);
nand U2711 (N_2711,N_2537,N_2400);
nand U2712 (N_2712,N_2495,N_2482);
nand U2713 (N_2713,N_2467,N_2452);
and U2714 (N_2714,N_2552,N_2534);
nand U2715 (N_2715,N_2544,N_2401);
nand U2716 (N_2716,N_2553,N_2527);
and U2717 (N_2717,N_2565,N_2504);
nand U2718 (N_2718,N_2490,N_2468);
nand U2719 (N_2719,N_2517,N_2541);
nand U2720 (N_2720,N_2419,N_2510);
xor U2721 (N_2721,N_2530,N_2560);
xnor U2722 (N_2722,N_2469,N_2569);
or U2723 (N_2723,N_2453,N_2464);
nor U2724 (N_2724,N_2474,N_2539);
and U2725 (N_2725,N_2518,N_2449);
or U2726 (N_2726,N_2590,N_2406);
nand U2727 (N_2727,N_2537,N_2446);
or U2728 (N_2728,N_2562,N_2435);
nor U2729 (N_2729,N_2598,N_2466);
nand U2730 (N_2730,N_2403,N_2528);
and U2731 (N_2731,N_2463,N_2527);
or U2732 (N_2732,N_2412,N_2477);
nor U2733 (N_2733,N_2561,N_2598);
xor U2734 (N_2734,N_2401,N_2511);
or U2735 (N_2735,N_2408,N_2462);
nand U2736 (N_2736,N_2578,N_2412);
or U2737 (N_2737,N_2446,N_2479);
nor U2738 (N_2738,N_2406,N_2510);
xor U2739 (N_2739,N_2538,N_2407);
xnor U2740 (N_2740,N_2527,N_2404);
nor U2741 (N_2741,N_2479,N_2471);
nand U2742 (N_2742,N_2590,N_2475);
nand U2743 (N_2743,N_2469,N_2557);
and U2744 (N_2744,N_2596,N_2506);
or U2745 (N_2745,N_2541,N_2512);
and U2746 (N_2746,N_2520,N_2449);
or U2747 (N_2747,N_2448,N_2537);
nor U2748 (N_2748,N_2401,N_2482);
and U2749 (N_2749,N_2485,N_2534);
xor U2750 (N_2750,N_2578,N_2594);
and U2751 (N_2751,N_2498,N_2426);
and U2752 (N_2752,N_2575,N_2583);
or U2753 (N_2753,N_2474,N_2580);
nor U2754 (N_2754,N_2453,N_2426);
and U2755 (N_2755,N_2450,N_2588);
nor U2756 (N_2756,N_2559,N_2440);
xnor U2757 (N_2757,N_2472,N_2541);
and U2758 (N_2758,N_2407,N_2445);
or U2759 (N_2759,N_2509,N_2454);
nor U2760 (N_2760,N_2408,N_2573);
nor U2761 (N_2761,N_2442,N_2492);
or U2762 (N_2762,N_2518,N_2547);
xnor U2763 (N_2763,N_2460,N_2521);
xor U2764 (N_2764,N_2431,N_2434);
and U2765 (N_2765,N_2426,N_2402);
and U2766 (N_2766,N_2420,N_2491);
nor U2767 (N_2767,N_2422,N_2582);
nand U2768 (N_2768,N_2560,N_2504);
nand U2769 (N_2769,N_2431,N_2504);
nor U2770 (N_2770,N_2510,N_2435);
xor U2771 (N_2771,N_2458,N_2549);
nor U2772 (N_2772,N_2502,N_2562);
nor U2773 (N_2773,N_2576,N_2518);
nand U2774 (N_2774,N_2404,N_2489);
or U2775 (N_2775,N_2500,N_2551);
or U2776 (N_2776,N_2444,N_2584);
or U2777 (N_2777,N_2580,N_2410);
or U2778 (N_2778,N_2590,N_2583);
nand U2779 (N_2779,N_2547,N_2418);
and U2780 (N_2780,N_2522,N_2505);
nor U2781 (N_2781,N_2541,N_2492);
nand U2782 (N_2782,N_2546,N_2515);
nand U2783 (N_2783,N_2426,N_2563);
xor U2784 (N_2784,N_2442,N_2589);
xnor U2785 (N_2785,N_2480,N_2500);
and U2786 (N_2786,N_2550,N_2510);
xor U2787 (N_2787,N_2411,N_2472);
and U2788 (N_2788,N_2559,N_2436);
xor U2789 (N_2789,N_2432,N_2574);
or U2790 (N_2790,N_2489,N_2484);
and U2791 (N_2791,N_2585,N_2495);
and U2792 (N_2792,N_2444,N_2546);
nor U2793 (N_2793,N_2414,N_2523);
or U2794 (N_2794,N_2486,N_2456);
nand U2795 (N_2795,N_2579,N_2465);
nor U2796 (N_2796,N_2427,N_2467);
nand U2797 (N_2797,N_2457,N_2499);
xor U2798 (N_2798,N_2511,N_2569);
or U2799 (N_2799,N_2584,N_2535);
nor U2800 (N_2800,N_2611,N_2636);
xnor U2801 (N_2801,N_2685,N_2624);
nand U2802 (N_2802,N_2601,N_2607);
xnor U2803 (N_2803,N_2658,N_2621);
or U2804 (N_2804,N_2723,N_2672);
and U2805 (N_2805,N_2620,N_2654);
nand U2806 (N_2806,N_2604,N_2681);
and U2807 (N_2807,N_2757,N_2650);
nor U2808 (N_2808,N_2762,N_2710);
nand U2809 (N_2809,N_2702,N_2662);
nor U2810 (N_2810,N_2722,N_2663);
and U2811 (N_2811,N_2694,N_2619);
or U2812 (N_2812,N_2706,N_2708);
nand U2813 (N_2813,N_2673,N_2798);
and U2814 (N_2814,N_2632,N_2637);
xor U2815 (N_2815,N_2605,N_2652);
or U2816 (N_2816,N_2678,N_2661);
xor U2817 (N_2817,N_2765,N_2742);
and U2818 (N_2818,N_2760,N_2704);
or U2819 (N_2819,N_2638,N_2764);
and U2820 (N_2820,N_2730,N_2697);
nand U2821 (N_2821,N_2747,N_2627);
or U2822 (N_2822,N_2689,N_2631);
and U2823 (N_2823,N_2660,N_2781);
xnor U2824 (N_2824,N_2616,N_2776);
or U2825 (N_2825,N_2749,N_2759);
and U2826 (N_2826,N_2609,N_2698);
and U2827 (N_2827,N_2664,N_2614);
xor U2828 (N_2828,N_2795,N_2653);
nor U2829 (N_2829,N_2770,N_2761);
nor U2830 (N_2830,N_2771,N_2623);
and U2831 (N_2831,N_2714,N_2777);
nor U2832 (N_2832,N_2726,N_2671);
nand U2833 (N_2833,N_2645,N_2602);
nand U2834 (N_2834,N_2766,N_2792);
nand U2835 (N_2835,N_2717,N_2625);
nor U2836 (N_2836,N_2745,N_2754);
nand U2837 (N_2837,N_2600,N_2768);
xor U2838 (N_2838,N_2750,N_2680);
and U2839 (N_2839,N_2786,N_2669);
and U2840 (N_2840,N_2629,N_2720);
nand U2841 (N_2841,N_2780,N_2646);
xor U2842 (N_2842,N_2793,N_2705);
and U2843 (N_2843,N_2736,N_2783);
and U2844 (N_2844,N_2670,N_2691);
or U2845 (N_2845,N_2612,N_2622);
xnor U2846 (N_2846,N_2740,N_2721);
nor U2847 (N_2847,N_2679,N_2751);
and U2848 (N_2848,N_2718,N_2642);
and U2849 (N_2849,N_2731,N_2635);
xor U2850 (N_2850,N_2606,N_2744);
nor U2851 (N_2851,N_2756,N_2692);
nand U2852 (N_2852,N_2758,N_2613);
nor U2853 (N_2853,N_2639,N_2787);
nand U2854 (N_2854,N_2659,N_2739);
and U2855 (N_2855,N_2729,N_2769);
xnor U2856 (N_2856,N_2633,N_2666);
or U2857 (N_2857,N_2703,N_2668);
nand U2858 (N_2858,N_2674,N_2615);
nand U2859 (N_2859,N_2647,N_2667);
xnor U2860 (N_2860,N_2763,N_2693);
nor U2861 (N_2861,N_2640,N_2695);
nor U2862 (N_2862,N_2700,N_2699);
or U2863 (N_2863,N_2779,N_2755);
or U2864 (N_2864,N_2711,N_2772);
and U2865 (N_2865,N_2648,N_2684);
and U2866 (N_2866,N_2649,N_2790);
nand U2867 (N_2867,N_2728,N_2709);
and U2868 (N_2868,N_2683,N_2785);
nand U2869 (N_2869,N_2707,N_2724);
xnor U2870 (N_2870,N_2686,N_2712);
and U2871 (N_2871,N_2799,N_2796);
and U2872 (N_2872,N_2676,N_2687);
nor U2873 (N_2873,N_2748,N_2746);
xor U2874 (N_2874,N_2719,N_2789);
nor U2875 (N_2875,N_2634,N_2696);
xnor U2876 (N_2876,N_2741,N_2767);
xor U2877 (N_2877,N_2733,N_2690);
xnor U2878 (N_2878,N_2784,N_2628);
nand U2879 (N_2879,N_2738,N_2713);
and U2880 (N_2880,N_2665,N_2752);
xor U2881 (N_2881,N_2773,N_2655);
nor U2882 (N_2882,N_2753,N_2618);
nor U2883 (N_2883,N_2774,N_2657);
nand U2884 (N_2884,N_2617,N_2608);
and U2885 (N_2885,N_2610,N_2716);
xor U2886 (N_2886,N_2644,N_2715);
xor U2887 (N_2887,N_2701,N_2682);
nor U2888 (N_2888,N_2732,N_2788);
and U2889 (N_2889,N_2734,N_2775);
xor U2890 (N_2890,N_2603,N_2743);
or U2891 (N_2891,N_2677,N_2778);
nand U2892 (N_2892,N_2675,N_2735);
nand U2893 (N_2893,N_2630,N_2791);
or U2894 (N_2894,N_2656,N_2797);
nor U2895 (N_2895,N_2651,N_2626);
nor U2896 (N_2896,N_2643,N_2782);
nor U2897 (N_2897,N_2725,N_2794);
xnor U2898 (N_2898,N_2641,N_2737);
xnor U2899 (N_2899,N_2727,N_2688);
xnor U2900 (N_2900,N_2679,N_2749);
nand U2901 (N_2901,N_2612,N_2609);
nor U2902 (N_2902,N_2623,N_2681);
nand U2903 (N_2903,N_2677,N_2767);
or U2904 (N_2904,N_2724,N_2663);
nor U2905 (N_2905,N_2785,N_2638);
nor U2906 (N_2906,N_2657,N_2744);
and U2907 (N_2907,N_2703,N_2684);
xnor U2908 (N_2908,N_2791,N_2744);
or U2909 (N_2909,N_2704,N_2795);
xnor U2910 (N_2910,N_2656,N_2717);
or U2911 (N_2911,N_2777,N_2682);
xnor U2912 (N_2912,N_2725,N_2724);
nor U2913 (N_2913,N_2692,N_2733);
and U2914 (N_2914,N_2634,N_2743);
nand U2915 (N_2915,N_2760,N_2677);
xnor U2916 (N_2916,N_2608,N_2653);
nand U2917 (N_2917,N_2718,N_2612);
and U2918 (N_2918,N_2635,N_2663);
xnor U2919 (N_2919,N_2736,N_2746);
and U2920 (N_2920,N_2686,N_2655);
nor U2921 (N_2921,N_2611,N_2665);
or U2922 (N_2922,N_2640,N_2731);
nand U2923 (N_2923,N_2784,N_2611);
nand U2924 (N_2924,N_2763,N_2658);
and U2925 (N_2925,N_2775,N_2631);
nand U2926 (N_2926,N_2671,N_2730);
or U2927 (N_2927,N_2613,N_2768);
or U2928 (N_2928,N_2730,N_2716);
or U2929 (N_2929,N_2757,N_2714);
or U2930 (N_2930,N_2656,N_2621);
nor U2931 (N_2931,N_2644,N_2712);
nand U2932 (N_2932,N_2789,N_2663);
xor U2933 (N_2933,N_2777,N_2638);
nand U2934 (N_2934,N_2730,N_2710);
xnor U2935 (N_2935,N_2708,N_2769);
or U2936 (N_2936,N_2742,N_2753);
nand U2937 (N_2937,N_2641,N_2741);
xor U2938 (N_2938,N_2759,N_2636);
and U2939 (N_2939,N_2764,N_2644);
or U2940 (N_2940,N_2601,N_2735);
nand U2941 (N_2941,N_2663,N_2709);
nor U2942 (N_2942,N_2789,N_2721);
xnor U2943 (N_2943,N_2602,N_2704);
xor U2944 (N_2944,N_2643,N_2640);
nand U2945 (N_2945,N_2615,N_2656);
nand U2946 (N_2946,N_2688,N_2662);
nand U2947 (N_2947,N_2603,N_2669);
and U2948 (N_2948,N_2787,N_2693);
and U2949 (N_2949,N_2735,N_2783);
nand U2950 (N_2950,N_2795,N_2640);
xnor U2951 (N_2951,N_2700,N_2677);
xnor U2952 (N_2952,N_2693,N_2625);
nand U2953 (N_2953,N_2606,N_2799);
nor U2954 (N_2954,N_2791,N_2745);
nand U2955 (N_2955,N_2791,N_2657);
and U2956 (N_2956,N_2741,N_2613);
nor U2957 (N_2957,N_2666,N_2740);
nor U2958 (N_2958,N_2645,N_2708);
xor U2959 (N_2959,N_2722,N_2685);
xnor U2960 (N_2960,N_2719,N_2763);
and U2961 (N_2961,N_2648,N_2685);
xnor U2962 (N_2962,N_2735,N_2792);
xor U2963 (N_2963,N_2703,N_2618);
or U2964 (N_2964,N_2634,N_2622);
nor U2965 (N_2965,N_2645,N_2631);
nor U2966 (N_2966,N_2649,N_2761);
and U2967 (N_2967,N_2635,N_2607);
and U2968 (N_2968,N_2618,N_2719);
xor U2969 (N_2969,N_2713,N_2769);
or U2970 (N_2970,N_2703,N_2665);
nand U2971 (N_2971,N_2744,N_2603);
xor U2972 (N_2972,N_2631,N_2755);
nand U2973 (N_2973,N_2635,N_2701);
xor U2974 (N_2974,N_2669,N_2694);
and U2975 (N_2975,N_2748,N_2656);
or U2976 (N_2976,N_2672,N_2603);
xor U2977 (N_2977,N_2662,N_2698);
or U2978 (N_2978,N_2720,N_2767);
or U2979 (N_2979,N_2673,N_2614);
and U2980 (N_2980,N_2745,N_2711);
nor U2981 (N_2981,N_2714,N_2616);
nor U2982 (N_2982,N_2757,N_2646);
and U2983 (N_2983,N_2738,N_2700);
xor U2984 (N_2984,N_2659,N_2668);
and U2985 (N_2985,N_2685,N_2687);
and U2986 (N_2986,N_2666,N_2678);
xor U2987 (N_2987,N_2796,N_2705);
xnor U2988 (N_2988,N_2731,N_2762);
and U2989 (N_2989,N_2780,N_2698);
or U2990 (N_2990,N_2789,N_2737);
nor U2991 (N_2991,N_2740,N_2778);
xor U2992 (N_2992,N_2717,N_2701);
xor U2993 (N_2993,N_2611,N_2750);
xnor U2994 (N_2994,N_2668,N_2724);
nand U2995 (N_2995,N_2696,N_2705);
nand U2996 (N_2996,N_2791,N_2620);
and U2997 (N_2997,N_2701,N_2698);
xor U2998 (N_2998,N_2759,N_2786);
nor U2999 (N_2999,N_2745,N_2603);
or U3000 (N_3000,N_2838,N_2912);
or U3001 (N_3001,N_2996,N_2911);
nand U3002 (N_3002,N_2950,N_2953);
or U3003 (N_3003,N_2801,N_2968);
nor U3004 (N_3004,N_2827,N_2805);
xor U3005 (N_3005,N_2837,N_2949);
nor U3006 (N_3006,N_2800,N_2978);
xor U3007 (N_3007,N_2807,N_2867);
xor U3008 (N_3008,N_2990,N_2983);
and U3009 (N_3009,N_2901,N_2850);
or U3010 (N_3010,N_2900,N_2834);
or U3011 (N_3011,N_2859,N_2981);
nand U3012 (N_3012,N_2813,N_2829);
nor U3013 (N_3013,N_2848,N_2874);
or U3014 (N_3014,N_2977,N_2988);
and U3015 (N_3015,N_2864,N_2931);
nor U3016 (N_3016,N_2811,N_2934);
or U3017 (N_3017,N_2964,N_2921);
nor U3018 (N_3018,N_2866,N_2865);
and U3019 (N_3019,N_2963,N_2979);
xor U3020 (N_3020,N_2843,N_2833);
or U3021 (N_3021,N_2962,N_2836);
and U3022 (N_3022,N_2839,N_2965);
xnor U3023 (N_3023,N_2902,N_2857);
xor U3024 (N_3024,N_2817,N_2909);
nand U3025 (N_3025,N_2890,N_2942);
or U3026 (N_3026,N_2893,N_2876);
or U3027 (N_3027,N_2885,N_2819);
nor U3028 (N_3028,N_2828,N_2926);
and U3029 (N_3029,N_2928,N_2967);
nor U3030 (N_3030,N_2896,N_2815);
or U3031 (N_3031,N_2980,N_2997);
and U3032 (N_3032,N_2913,N_2892);
nor U3033 (N_3033,N_2869,N_2899);
xnor U3034 (N_3034,N_2898,N_2835);
nor U3035 (N_3035,N_2861,N_2881);
xnor U3036 (N_3036,N_2841,N_2952);
or U3037 (N_3037,N_2930,N_2916);
or U3038 (N_3038,N_2948,N_2907);
xor U3039 (N_3039,N_2856,N_2989);
or U3040 (N_3040,N_2944,N_2973);
nand U3041 (N_3041,N_2905,N_2895);
nor U3042 (N_3042,N_2941,N_2947);
xnor U3043 (N_3043,N_2825,N_2936);
and U3044 (N_3044,N_2946,N_2940);
xor U3045 (N_3045,N_2812,N_2903);
nand U3046 (N_3046,N_2814,N_2802);
nand U3047 (N_3047,N_2976,N_2927);
xnor U3048 (N_3048,N_2938,N_2974);
or U3049 (N_3049,N_2832,N_2993);
nor U3050 (N_3050,N_2932,N_2826);
and U3051 (N_3051,N_2957,N_2924);
xnor U3052 (N_3052,N_2886,N_2919);
nor U3053 (N_3053,N_2831,N_2958);
or U3054 (N_3054,N_2917,N_2860);
nand U3055 (N_3055,N_2822,N_2808);
nor U3056 (N_3056,N_2880,N_2803);
xor U3057 (N_3057,N_2854,N_2945);
xor U3058 (N_3058,N_2966,N_2875);
nand U3059 (N_3059,N_2969,N_2956);
and U3060 (N_3060,N_2972,N_2852);
or U3061 (N_3061,N_2960,N_2820);
nand U3062 (N_3062,N_2862,N_2821);
nand U3063 (N_3063,N_2824,N_2830);
nand U3064 (N_3064,N_2954,N_2918);
and U3065 (N_3065,N_2987,N_2884);
nand U3066 (N_3066,N_2994,N_2809);
or U3067 (N_3067,N_2925,N_2951);
nor U3068 (N_3068,N_2998,N_2889);
or U3069 (N_3069,N_2975,N_2970);
nand U3070 (N_3070,N_2894,N_2806);
or U3071 (N_3071,N_2882,N_2816);
xor U3072 (N_3072,N_2986,N_2877);
nand U3073 (N_3073,N_2863,N_2840);
or U3074 (N_3074,N_2904,N_2914);
or U3075 (N_3075,N_2851,N_2937);
and U3076 (N_3076,N_2823,N_2935);
nand U3077 (N_3077,N_2878,N_2995);
and U3078 (N_3078,N_2871,N_2910);
or U3079 (N_3079,N_2915,N_2872);
nor U3080 (N_3080,N_2906,N_2804);
and U3081 (N_3081,N_2923,N_2853);
and U3082 (N_3082,N_2984,N_2845);
or U3083 (N_3083,N_2846,N_2929);
or U3084 (N_3084,N_2943,N_2920);
nor U3085 (N_3085,N_2922,N_2810);
xnor U3086 (N_3086,N_2992,N_2891);
nand U3087 (N_3087,N_2842,N_2933);
xnor U3088 (N_3088,N_2858,N_2847);
nand U3089 (N_3089,N_2870,N_2897);
nor U3090 (N_3090,N_2879,N_2982);
or U3091 (N_3091,N_2999,N_2985);
nand U3092 (N_3092,N_2868,N_2955);
nor U3093 (N_3093,N_2888,N_2818);
nor U3094 (N_3094,N_2887,N_2883);
and U3095 (N_3095,N_2971,N_2959);
nand U3096 (N_3096,N_2939,N_2844);
nand U3097 (N_3097,N_2849,N_2961);
nor U3098 (N_3098,N_2873,N_2908);
xnor U3099 (N_3099,N_2855,N_2991);
nand U3100 (N_3100,N_2992,N_2943);
nand U3101 (N_3101,N_2990,N_2866);
nor U3102 (N_3102,N_2846,N_2992);
and U3103 (N_3103,N_2802,N_2933);
or U3104 (N_3104,N_2828,N_2908);
xnor U3105 (N_3105,N_2859,N_2878);
nand U3106 (N_3106,N_2915,N_2810);
nor U3107 (N_3107,N_2815,N_2963);
xnor U3108 (N_3108,N_2968,N_2848);
nor U3109 (N_3109,N_2870,N_2893);
nand U3110 (N_3110,N_2990,N_2805);
and U3111 (N_3111,N_2883,N_2982);
nand U3112 (N_3112,N_2962,N_2817);
or U3113 (N_3113,N_2825,N_2869);
and U3114 (N_3114,N_2880,N_2967);
xor U3115 (N_3115,N_2806,N_2815);
nor U3116 (N_3116,N_2955,N_2858);
xnor U3117 (N_3117,N_2817,N_2955);
xor U3118 (N_3118,N_2865,N_2988);
or U3119 (N_3119,N_2979,N_2887);
xnor U3120 (N_3120,N_2932,N_2805);
nor U3121 (N_3121,N_2958,N_2816);
or U3122 (N_3122,N_2919,N_2848);
and U3123 (N_3123,N_2983,N_2916);
nand U3124 (N_3124,N_2946,N_2941);
or U3125 (N_3125,N_2976,N_2960);
nor U3126 (N_3126,N_2926,N_2865);
nand U3127 (N_3127,N_2867,N_2819);
nor U3128 (N_3128,N_2923,N_2999);
nor U3129 (N_3129,N_2933,N_2983);
nor U3130 (N_3130,N_2931,N_2904);
nor U3131 (N_3131,N_2849,N_2876);
nor U3132 (N_3132,N_2989,N_2945);
nand U3133 (N_3133,N_2834,N_2839);
and U3134 (N_3134,N_2829,N_2856);
nor U3135 (N_3135,N_2970,N_2861);
nor U3136 (N_3136,N_2881,N_2962);
xnor U3137 (N_3137,N_2836,N_2804);
nor U3138 (N_3138,N_2836,N_2882);
xnor U3139 (N_3139,N_2808,N_2946);
nand U3140 (N_3140,N_2800,N_2811);
or U3141 (N_3141,N_2804,N_2848);
or U3142 (N_3142,N_2861,N_2831);
xnor U3143 (N_3143,N_2949,N_2810);
and U3144 (N_3144,N_2885,N_2849);
xnor U3145 (N_3145,N_2967,N_2996);
nand U3146 (N_3146,N_2859,N_2852);
xnor U3147 (N_3147,N_2921,N_2857);
nand U3148 (N_3148,N_2929,N_2879);
xnor U3149 (N_3149,N_2855,N_2973);
nand U3150 (N_3150,N_2897,N_2867);
or U3151 (N_3151,N_2890,N_2815);
and U3152 (N_3152,N_2813,N_2858);
nor U3153 (N_3153,N_2818,N_2902);
nand U3154 (N_3154,N_2886,N_2892);
or U3155 (N_3155,N_2940,N_2877);
xor U3156 (N_3156,N_2833,N_2984);
nor U3157 (N_3157,N_2903,N_2932);
nand U3158 (N_3158,N_2856,N_2802);
or U3159 (N_3159,N_2833,N_2909);
and U3160 (N_3160,N_2867,N_2811);
nand U3161 (N_3161,N_2989,N_2909);
nand U3162 (N_3162,N_2944,N_2849);
and U3163 (N_3163,N_2965,N_2804);
nand U3164 (N_3164,N_2986,N_2906);
nand U3165 (N_3165,N_2805,N_2945);
or U3166 (N_3166,N_2979,N_2806);
xor U3167 (N_3167,N_2968,N_2826);
nor U3168 (N_3168,N_2923,N_2930);
and U3169 (N_3169,N_2851,N_2889);
nand U3170 (N_3170,N_2920,N_2975);
nand U3171 (N_3171,N_2885,N_2938);
xnor U3172 (N_3172,N_2864,N_2965);
xnor U3173 (N_3173,N_2916,N_2832);
and U3174 (N_3174,N_2820,N_2883);
nand U3175 (N_3175,N_2855,N_2947);
nand U3176 (N_3176,N_2862,N_2869);
xor U3177 (N_3177,N_2849,N_2863);
and U3178 (N_3178,N_2831,N_2989);
or U3179 (N_3179,N_2819,N_2843);
or U3180 (N_3180,N_2876,N_2998);
xnor U3181 (N_3181,N_2817,N_2809);
and U3182 (N_3182,N_2865,N_2861);
nor U3183 (N_3183,N_2997,N_2964);
nor U3184 (N_3184,N_2990,N_2975);
xor U3185 (N_3185,N_2850,N_2812);
and U3186 (N_3186,N_2834,N_2877);
nand U3187 (N_3187,N_2815,N_2999);
xnor U3188 (N_3188,N_2900,N_2986);
nand U3189 (N_3189,N_2909,N_2937);
nand U3190 (N_3190,N_2952,N_2879);
and U3191 (N_3191,N_2938,N_2836);
or U3192 (N_3192,N_2916,N_2933);
xor U3193 (N_3193,N_2919,N_2959);
nor U3194 (N_3194,N_2837,N_2896);
and U3195 (N_3195,N_2877,N_2970);
or U3196 (N_3196,N_2849,N_2865);
xor U3197 (N_3197,N_2892,N_2987);
and U3198 (N_3198,N_2991,N_2845);
xor U3199 (N_3199,N_2988,N_2853);
nand U3200 (N_3200,N_3032,N_3055);
nor U3201 (N_3201,N_3090,N_3084);
xnor U3202 (N_3202,N_3120,N_3148);
nor U3203 (N_3203,N_3106,N_3174);
nor U3204 (N_3204,N_3069,N_3087);
nand U3205 (N_3205,N_3089,N_3104);
xnor U3206 (N_3206,N_3024,N_3199);
nand U3207 (N_3207,N_3077,N_3165);
or U3208 (N_3208,N_3196,N_3149);
nand U3209 (N_3209,N_3125,N_3096);
or U3210 (N_3210,N_3137,N_3117);
xnor U3211 (N_3211,N_3029,N_3160);
nor U3212 (N_3212,N_3133,N_3092);
nor U3213 (N_3213,N_3008,N_3152);
nand U3214 (N_3214,N_3060,N_3080);
or U3215 (N_3215,N_3019,N_3054);
nand U3216 (N_3216,N_3094,N_3138);
nor U3217 (N_3217,N_3097,N_3088);
or U3218 (N_3218,N_3131,N_3041);
xnor U3219 (N_3219,N_3095,N_3052);
and U3220 (N_3220,N_3048,N_3122);
or U3221 (N_3221,N_3134,N_3187);
and U3222 (N_3222,N_3033,N_3103);
and U3223 (N_3223,N_3079,N_3176);
nor U3224 (N_3224,N_3059,N_3034);
or U3225 (N_3225,N_3167,N_3166);
and U3226 (N_3226,N_3171,N_3023);
xnor U3227 (N_3227,N_3040,N_3028);
and U3228 (N_3228,N_3169,N_3192);
nand U3229 (N_3229,N_3156,N_3082);
nor U3230 (N_3230,N_3045,N_3142);
and U3231 (N_3231,N_3065,N_3011);
nand U3232 (N_3232,N_3015,N_3100);
nor U3233 (N_3233,N_3067,N_3083);
or U3234 (N_3234,N_3189,N_3136);
or U3235 (N_3235,N_3107,N_3158);
nor U3236 (N_3236,N_3168,N_3042);
xnor U3237 (N_3237,N_3190,N_3074);
nor U3238 (N_3238,N_3001,N_3162);
or U3239 (N_3239,N_3066,N_3078);
xor U3240 (N_3240,N_3073,N_3068);
nand U3241 (N_3241,N_3075,N_3180);
and U3242 (N_3242,N_3076,N_3184);
and U3243 (N_3243,N_3007,N_3081);
nor U3244 (N_3244,N_3173,N_3056);
and U3245 (N_3245,N_3113,N_3179);
nor U3246 (N_3246,N_3026,N_3153);
nand U3247 (N_3247,N_3004,N_3126);
nor U3248 (N_3248,N_3058,N_3013);
and U3249 (N_3249,N_3036,N_3195);
nor U3250 (N_3250,N_3016,N_3177);
and U3251 (N_3251,N_3038,N_3050);
xnor U3252 (N_3252,N_3157,N_3147);
and U3253 (N_3253,N_3099,N_3186);
and U3254 (N_3254,N_3151,N_3030);
or U3255 (N_3255,N_3150,N_3010);
nor U3256 (N_3256,N_3020,N_3051);
nand U3257 (N_3257,N_3039,N_3098);
nand U3258 (N_3258,N_3123,N_3044);
nand U3259 (N_3259,N_3127,N_3183);
or U3260 (N_3260,N_3110,N_3116);
nor U3261 (N_3261,N_3049,N_3062);
and U3262 (N_3262,N_3071,N_3053);
nand U3263 (N_3263,N_3035,N_3182);
and U3264 (N_3264,N_3021,N_3057);
and U3265 (N_3265,N_3188,N_3197);
or U3266 (N_3266,N_3121,N_3018);
and U3267 (N_3267,N_3119,N_3118);
xnor U3268 (N_3268,N_3002,N_3114);
xnor U3269 (N_3269,N_3014,N_3086);
and U3270 (N_3270,N_3129,N_3159);
nor U3271 (N_3271,N_3006,N_3144);
nor U3272 (N_3272,N_3009,N_3145);
xnor U3273 (N_3273,N_3108,N_3064);
or U3274 (N_3274,N_3164,N_3141);
and U3275 (N_3275,N_3025,N_3130);
or U3276 (N_3276,N_3155,N_3198);
nand U3277 (N_3277,N_3178,N_3161);
and U3278 (N_3278,N_3191,N_3132);
nor U3279 (N_3279,N_3193,N_3109);
nor U3280 (N_3280,N_3135,N_3163);
xnor U3281 (N_3281,N_3146,N_3063);
nor U3282 (N_3282,N_3194,N_3061);
nand U3283 (N_3283,N_3017,N_3031);
nor U3284 (N_3284,N_3139,N_3027);
and U3285 (N_3285,N_3000,N_3005);
or U3286 (N_3286,N_3093,N_3085);
and U3287 (N_3287,N_3043,N_3143);
xnor U3288 (N_3288,N_3105,N_3175);
nand U3289 (N_3289,N_3003,N_3012);
nand U3290 (N_3290,N_3124,N_3037);
or U3291 (N_3291,N_3112,N_3072);
or U3292 (N_3292,N_3172,N_3046);
nor U3293 (N_3293,N_3115,N_3022);
and U3294 (N_3294,N_3181,N_3070);
and U3295 (N_3295,N_3102,N_3047);
or U3296 (N_3296,N_3154,N_3091);
or U3297 (N_3297,N_3101,N_3185);
xnor U3298 (N_3298,N_3111,N_3128);
or U3299 (N_3299,N_3140,N_3170);
nor U3300 (N_3300,N_3134,N_3196);
xnor U3301 (N_3301,N_3126,N_3139);
nand U3302 (N_3302,N_3124,N_3105);
or U3303 (N_3303,N_3163,N_3158);
xnor U3304 (N_3304,N_3052,N_3073);
nor U3305 (N_3305,N_3074,N_3186);
nor U3306 (N_3306,N_3103,N_3060);
nor U3307 (N_3307,N_3192,N_3054);
and U3308 (N_3308,N_3193,N_3118);
or U3309 (N_3309,N_3086,N_3169);
nand U3310 (N_3310,N_3197,N_3163);
or U3311 (N_3311,N_3171,N_3181);
xnor U3312 (N_3312,N_3094,N_3199);
xnor U3313 (N_3313,N_3095,N_3188);
xor U3314 (N_3314,N_3011,N_3102);
nand U3315 (N_3315,N_3104,N_3027);
or U3316 (N_3316,N_3082,N_3155);
nand U3317 (N_3317,N_3161,N_3159);
nor U3318 (N_3318,N_3093,N_3034);
xor U3319 (N_3319,N_3167,N_3180);
nor U3320 (N_3320,N_3071,N_3135);
nand U3321 (N_3321,N_3120,N_3035);
xnor U3322 (N_3322,N_3121,N_3111);
nor U3323 (N_3323,N_3034,N_3134);
xor U3324 (N_3324,N_3011,N_3116);
or U3325 (N_3325,N_3029,N_3011);
xor U3326 (N_3326,N_3063,N_3109);
and U3327 (N_3327,N_3149,N_3199);
or U3328 (N_3328,N_3159,N_3127);
and U3329 (N_3329,N_3081,N_3061);
nand U3330 (N_3330,N_3125,N_3089);
nor U3331 (N_3331,N_3108,N_3132);
xor U3332 (N_3332,N_3109,N_3017);
xnor U3333 (N_3333,N_3017,N_3026);
and U3334 (N_3334,N_3190,N_3135);
xnor U3335 (N_3335,N_3117,N_3024);
or U3336 (N_3336,N_3086,N_3027);
nand U3337 (N_3337,N_3113,N_3101);
xor U3338 (N_3338,N_3085,N_3148);
xor U3339 (N_3339,N_3082,N_3153);
xnor U3340 (N_3340,N_3042,N_3111);
and U3341 (N_3341,N_3101,N_3096);
or U3342 (N_3342,N_3159,N_3148);
and U3343 (N_3343,N_3187,N_3127);
xor U3344 (N_3344,N_3121,N_3157);
and U3345 (N_3345,N_3102,N_3032);
and U3346 (N_3346,N_3044,N_3134);
or U3347 (N_3347,N_3076,N_3009);
or U3348 (N_3348,N_3189,N_3041);
xor U3349 (N_3349,N_3020,N_3112);
and U3350 (N_3350,N_3159,N_3126);
and U3351 (N_3351,N_3020,N_3157);
nor U3352 (N_3352,N_3160,N_3079);
or U3353 (N_3353,N_3146,N_3060);
and U3354 (N_3354,N_3190,N_3157);
and U3355 (N_3355,N_3173,N_3034);
nand U3356 (N_3356,N_3113,N_3138);
nor U3357 (N_3357,N_3008,N_3013);
or U3358 (N_3358,N_3176,N_3151);
nand U3359 (N_3359,N_3041,N_3032);
and U3360 (N_3360,N_3018,N_3152);
nand U3361 (N_3361,N_3014,N_3192);
or U3362 (N_3362,N_3128,N_3022);
or U3363 (N_3363,N_3075,N_3051);
xnor U3364 (N_3364,N_3033,N_3049);
xor U3365 (N_3365,N_3038,N_3059);
xnor U3366 (N_3366,N_3039,N_3049);
nor U3367 (N_3367,N_3057,N_3185);
and U3368 (N_3368,N_3026,N_3041);
nand U3369 (N_3369,N_3132,N_3129);
nand U3370 (N_3370,N_3143,N_3189);
xnor U3371 (N_3371,N_3070,N_3145);
and U3372 (N_3372,N_3144,N_3019);
or U3373 (N_3373,N_3150,N_3132);
xor U3374 (N_3374,N_3136,N_3170);
nor U3375 (N_3375,N_3192,N_3089);
xor U3376 (N_3376,N_3095,N_3036);
nor U3377 (N_3377,N_3004,N_3085);
or U3378 (N_3378,N_3147,N_3050);
nor U3379 (N_3379,N_3151,N_3047);
nand U3380 (N_3380,N_3090,N_3128);
and U3381 (N_3381,N_3043,N_3158);
nor U3382 (N_3382,N_3028,N_3023);
xnor U3383 (N_3383,N_3016,N_3018);
and U3384 (N_3384,N_3062,N_3125);
or U3385 (N_3385,N_3084,N_3039);
and U3386 (N_3386,N_3029,N_3199);
nand U3387 (N_3387,N_3101,N_3168);
nand U3388 (N_3388,N_3152,N_3061);
or U3389 (N_3389,N_3068,N_3074);
xor U3390 (N_3390,N_3137,N_3161);
and U3391 (N_3391,N_3055,N_3139);
nor U3392 (N_3392,N_3192,N_3179);
nand U3393 (N_3393,N_3119,N_3189);
nor U3394 (N_3394,N_3049,N_3125);
or U3395 (N_3395,N_3037,N_3116);
and U3396 (N_3396,N_3048,N_3069);
and U3397 (N_3397,N_3108,N_3028);
xnor U3398 (N_3398,N_3105,N_3123);
nor U3399 (N_3399,N_3036,N_3056);
nor U3400 (N_3400,N_3361,N_3328);
or U3401 (N_3401,N_3362,N_3381);
or U3402 (N_3402,N_3283,N_3336);
nor U3403 (N_3403,N_3372,N_3228);
and U3404 (N_3404,N_3212,N_3257);
and U3405 (N_3405,N_3256,N_3326);
nand U3406 (N_3406,N_3255,N_3285);
nand U3407 (N_3407,N_3376,N_3341);
xnor U3408 (N_3408,N_3277,N_3245);
or U3409 (N_3409,N_3281,N_3315);
nor U3410 (N_3410,N_3343,N_3317);
or U3411 (N_3411,N_3339,N_3370);
nand U3412 (N_3412,N_3221,N_3349);
nor U3413 (N_3413,N_3288,N_3269);
nor U3414 (N_3414,N_3322,N_3214);
nand U3415 (N_3415,N_3387,N_3286);
or U3416 (N_3416,N_3330,N_3350);
xnor U3417 (N_3417,N_3394,N_3296);
or U3418 (N_3418,N_3204,N_3272);
or U3419 (N_3419,N_3385,N_3319);
xor U3420 (N_3420,N_3201,N_3226);
or U3421 (N_3421,N_3227,N_3267);
xor U3422 (N_3422,N_3359,N_3300);
or U3423 (N_3423,N_3305,N_3251);
nand U3424 (N_3424,N_3247,N_3383);
nand U3425 (N_3425,N_3232,N_3364);
nand U3426 (N_3426,N_3241,N_3211);
and U3427 (N_3427,N_3301,N_3260);
and U3428 (N_3428,N_3252,N_3268);
or U3429 (N_3429,N_3363,N_3275);
or U3430 (N_3430,N_3235,N_3389);
xor U3431 (N_3431,N_3205,N_3324);
or U3432 (N_3432,N_3332,N_3248);
and U3433 (N_3433,N_3230,N_3384);
and U3434 (N_3434,N_3331,N_3207);
xnor U3435 (N_3435,N_3292,N_3274);
nor U3436 (N_3436,N_3264,N_3223);
nand U3437 (N_3437,N_3271,N_3365);
and U3438 (N_3438,N_3311,N_3282);
xnor U3439 (N_3439,N_3346,N_3279);
nor U3440 (N_3440,N_3342,N_3373);
nor U3441 (N_3441,N_3391,N_3357);
nor U3442 (N_3442,N_3378,N_3367);
or U3443 (N_3443,N_3392,N_3234);
nand U3444 (N_3444,N_3360,N_3289);
nor U3445 (N_3445,N_3395,N_3345);
nand U3446 (N_3446,N_3219,N_3368);
xnor U3447 (N_3447,N_3351,N_3276);
xor U3448 (N_3448,N_3278,N_3229);
nand U3449 (N_3449,N_3356,N_3240);
xnor U3450 (N_3450,N_3294,N_3329);
and U3451 (N_3451,N_3273,N_3318);
or U3452 (N_3452,N_3284,N_3388);
nor U3453 (N_3453,N_3390,N_3246);
or U3454 (N_3454,N_3263,N_3323);
nor U3455 (N_3455,N_3344,N_3254);
and U3456 (N_3456,N_3242,N_3215);
xor U3457 (N_3457,N_3220,N_3354);
nand U3458 (N_3458,N_3216,N_3217);
nor U3459 (N_3459,N_3386,N_3369);
nor U3460 (N_3460,N_3222,N_3313);
and U3461 (N_3461,N_3398,N_3335);
or U3462 (N_3462,N_3209,N_3358);
or U3463 (N_3463,N_3262,N_3314);
or U3464 (N_3464,N_3287,N_3377);
nand U3465 (N_3465,N_3347,N_3352);
xor U3466 (N_3466,N_3213,N_3338);
nand U3467 (N_3467,N_3397,N_3308);
or U3468 (N_3468,N_3253,N_3303);
nand U3469 (N_3469,N_3224,N_3366);
and U3470 (N_3470,N_3225,N_3316);
or U3471 (N_3471,N_3348,N_3320);
or U3472 (N_3472,N_3304,N_3243);
or U3473 (N_3473,N_3250,N_3295);
nor U3474 (N_3474,N_3293,N_3393);
and U3475 (N_3475,N_3297,N_3299);
nor U3476 (N_3476,N_3333,N_3327);
xor U3477 (N_3477,N_3265,N_3249);
nand U3478 (N_3478,N_3298,N_3306);
and U3479 (N_3479,N_3290,N_3259);
or U3480 (N_3480,N_3379,N_3355);
or U3481 (N_3481,N_3337,N_3380);
nand U3482 (N_3482,N_3309,N_3202);
or U3483 (N_3483,N_3237,N_3210);
and U3484 (N_3484,N_3334,N_3382);
and U3485 (N_3485,N_3340,N_3321);
nand U3486 (N_3486,N_3371,N_3233);
nand U3487 (N_3487,N_3261,N_3353);
nor U3488 (N_3488,N_3325,N_3231);
nor U3489 (N_3489,N_3270,N_3208);
nand U3490 (N_3490,N_3291,N_3312);
nor U3491 (N_3491,N_3396,N_3218);
xnor U3492 (N_3492,N_3399,N_3244);
nor U3493 (N_3493,N_3310,N_3374);
and U3494 (N_3494,N_3200,N_3203);
nand U3495 (N_3495,N_3307,N_3238);
or U3496 (N_3496,N_3236,N_3206);
and U3497 (N_3497,N_3239,N_3302);
and U3498 (N_3498,N_3266,N_3258);
and U3499 (N_3499,N_3375,N_3280);
nand U3500 (N_3500,N_3352,N_3267);
nand U3501 (N_3501,N_3379,N_3305);
nor U3502 (N_3502,N_3265,N_3358);
xnor U3503 (N_3503,N_3395,N_3230);
or U3504 (N_3504,N_3241,N_3202);
xnor U3505 (N_3505,N_3396,N_3235);
nand U3506 (N_3506,N_3230,N_3223);
or U3507 (N_3507,N_3237,N_3225);
and U3508 (N_3508,N_3301,N_3300);
nor U3509 (N_3509,N_3222,N_3245);
nor U3510 (N_3510,N_3295,N_3273);
xor U3511 (N_3511,N_3311,N_3357);
xor U3512 (N_3512,N_3229,N_3344);
nand U3513 (N_3513,N_3255,N_3223);
nand U3514 (N_3514,N_3316,N_3246);
nand U3515 (N_3515,N_3356,N_3276);
or U3516 (N_3516,N_3256,N_3345);
xnor U3517 (N_3517,N_3280,N_3321);
or U3518 (N_3518,N_3243,N_3207);
and U3519 (N_3519,N_3364,N_3240);
or U3520 (N_3520,N_3356,N_3331);
or U3521 (N_3521,N_3260,N_3203);
xnor U3522 (N_3522,N_3230,N_3213);
and U3523 (N_3523,N_3383,N_3256);
nor U3524 (N_3524,N_3286,N_3260);
xor U3525 (N_3525,N_3272,N_3352);
nor U3526 (N_3526,N_3336,N_3255);
xnor U3527 (N_3527,N_3222,N_3286);
or U3528 (N_3528,N_3359,N_3233);
and U3529 (N_3529,N_3390,N_3204);
nand U3530 (N_3530,N_3361,N_3222);
nor U3531 (N_3531,N_3294,N_3264);
nor U3532 (N_3532,N_3281,N_3391);
xor U3533 (N_3533,N_3282,N_3276);
nand U3534 (N_3534,N_3283,N_3319);
nand U3535 (N_3535,N_3291,N_3346);
and U3536 (N_3536,N_3340,N_3262);
xnor U3537 (N_3537,N_3263,N_3288);
nand U3538 (N_3538,N_3210,N_3273);
xor U3539 (N_3539,N_3275,N_3358);
or U3540 (N_3540,N_3221,N_3305);
xor U3541 (N_3541,N_3280,N_3322);
xnor U3542 (N_3542,N_3229,N_3374);
and U3543 (N_3543,N_3259,N_3398);
nand U3544 (N_3544,N_3284,N_3237);
or U3545 (N_3545,N_3236,N_3354);
nor U3546 (N_3546,N_3223,N_3372);
xor U3547 (N_3547,N_3277,N_3365);
nand U3548 (N_3548,N_3298,N_3294);
and U3549 (N_3549,N_3212,N_3344);
and U3550 (N_3550,N_3377,N_3301);
xnor U3551 (N_3551,N_3223,N_3388);
and U3552 (N_3552,N_3311,N_3235);
or U3553 (N_3553,N_3262,N_3331);
or U3554 (N_3554,N_3250,N_3384);
xnor U3555 (N_3555,N_3234,N_3312);
xnor U3556 (N_3556,N_3356,N_3255);
or U3557 (N_3557,N_3312,N_3252);
or U3558 (N_3558,N_3236,N_3269);
xor U3559 (N_3559,N_3249,N_3272);
nand U3560 (N_3560,N_3234,N_3246);
or U3561 (N_3561,N_3273,N_3320);
or U3562 (N_3562,N_3267,N_3317);
and U3563 (N_3563,N_3388,N_3256);
nand U3564 (N_3564,N_3391,N_3237);
nor U3565 (N_3565,N_3315,N_3259);
or U3566 (N_3566,N_3366,N_3387);
nand U3567 (N_3567,N_3396,N_3371);
or U3568 (N_3568,N_3251,N_3394);
nand U3569 (N_3569,N_3262,N_3389);
and U3570 (N_3570,N_3355,N_3358);
xor U3571 (N_3571,N_3365,N_3228);
nor U3572 (N_3572,N_3247,N_3374);
nand U3573 (N_3573,N_3270,N_3286);
and U3574 (N_3574,N_3211,N_3289);
nor U3575 (N_3575,N_3285,N_3378);
and U3576 (N_3576,N_3230,N_3337);
xor U3577 (N_3577,N_3289,N_3249);
or U3578 (N_3578,N_3314,N_3392);
nand U3579 (N_3579,N_3300,N_3311);
and U3580 (N_3580,N_3361,N_3295);
nand U3581 (N_3581,N_3393,N_3349);
nand U3582 (N_3582,N_3247,N_3306);
and U3583 (N_3583,N_3386,N_3364);
nor U3584 (N_3584,N_3251,N_3286);
nor U3585 (N_3585,N_3323,N_3273);
nand U3586 (N_3586,N_3390,N_3321);
nor U3587 (N_3587,N_3293,N_3271);
nand U3588 (N_3588,N_3253,N_3326);
or U3589 (N_3589,N_3338,N_3346);
nor U3590 (N_3590,N_3302,N_3383);
or U3591 (N_3591,N_3379,N_3294);
xor U3592 (N_3592,N_3260,N_3249);
xor U3593 (N_3593,N_3385,N_3322);
and U3594 (N_3594,N_3356,N_3368);
nor U3595 (N_3595,N_3215,N_3284);
or U3596 (N_3596,N_3269,N_3243);
nand U3597 (N_3597,N_3342,N_3275);
and U3598 (N_3598,N_3349,N_3367);
xnor U3599 (N_3599,N_3367,N_3255);
nand U3600 (N_3600,N_3510,N_3578);
and U3601 (N_3601,N_3404,N_3539);
nor U3602 (N_3602,N_3563,N_3569);
or U3603 (N_3603,N_3464,N_3587);
xnor U3604 (N_3604,N_3504,N_3544);
nand U3605 (N_3605,N_3523,N_3541);
nand U3606 (N_3606,N_3502,N_3490);
and U3607 (N_3607,N_3420,N_3434);
nand U3608 (N_3608,N_3535,N_3422);
or U3609 (N_3609,N_3497,N_3531);
xnor U3610 (N_3610,N_3577,N_3586);
or U3611 (N_3611,N_3468,N_3459);
nand U3612 (N_3612,N_3414,N_3552);
xor U3613 (N_3613,N_3448,N_3551);
or U3614 (N_3614,N_3425,N_3482);
and U3615 (N_3615,N_3528,N_3565);
xor U3616 (N_3616,N_3471,N_3534);
nand U3617 (N_3617,N_3419,N_3584);
and U3618 (N_3618,N_3516,N_3579);
xor U3619 (N_3619,N_3407,N_3598);
nand U3620 (N_3620,N_3415,N_3472);
xor U3621 (N_3621,N_3431,N_3596);
nand U3622 (N_3622,N_3462,N_3485);
or U3623 (N_3623,N_3483,N_3487);
and U3624 (N_3624,N_3580,N_3532);
or U3625 (N_3625,N_3517,N_3403);
xor U3626 (N_3626,N_3488,N_3410);
xor U3627 (N_3627,N_3426,N_3424);
nor U3628 (N_3628,N_3455,N_3494);
nor U3629 (N_3629,N_3433,N_3540);
xnor U3630 (N_3630,N_3521,N_3545);
nor U3631 (N_3631,N_3416,N_3476);
nor U3632 (N_3632,N_3595,N_3511);
or U3633 (N_3633,N_3445,N_3499);
xnor U3634 (N_3634,N_3439,N_3553);
nor U3635 (N_3635,N_3430,N_3457);
nand U3636 (N_3636,N_3489,N_3571);
nand U3637 (N_3637,N_3465,N_3546);
nor U3638 (N_3638,N_3458,N_3493);
and U3639 (N_3639,N_3581,N_3543);
and U3640 (N_3640,N_3484,N_3442);
nand U3641 (N_3641,N_3550,N_3437);
nand U3642 (N_3642,N_3583,N_3573);
nor U3643 (N_3643,N_3466,N_3594);
or U3644 (N_3644,N_3500,N_3556);
and U3645 (N_3645,N_3401,N_3507);
nand U3646 (N_3646,N_3402,N_3412);
and U3647 (N_3647,N_3557,N_3505);
nor U3648 (N_3648,N_3460,N_3486);
or U3649 (N_3649,N_3428,N_3559);
xnor U3650 (N_3650,N_3512,N_3526);
nor U3651 (N_3651,N_3548,N_3436);
and U3652 (N_3652,N_3566,N_3574);
or U3653 (N_3653,N_3525,N_3506);
and U3654 (N_3654,N_3496,N_3441);
and U3655 (N_3655,N_3452,N_3474);
or U3656 (N_3656,N_3406,N_3570);
nor U3657 (N_3657,N_3519,N_3467);
nand U3658 (N_3658,N_3405,N_3447);
nor U3659 (N_3659,N_3492,N_3520);
and U3660 (N_3660,N_3562,N_3530);
nand U3661 (N_3661,N_3537,N_3588);
and U3662 (N_3662,N_3427,N_3440);
nor U3663 (N_3663,N_3429,N_3538);
xnor U3664 (N_3664,N_3478,N_3590);
nand U3665 (N_3665,N_3443,N_3582);
nand U3666 (N_3666,N_3451,N_3515);
xnor U3667 (N_3667,N_3423,N_3514);
xor U3668 (N_3668,N_3524,N_3438);
or U3669 (N_3669,N_3585,N_3498);
and U3670 (N_3670,N_3572,N_3555);
nand U3671 (N_3671,N_3454,N_3513);
nand U3672 (N_3672,N_3473,N_3592);
nor U3673 (N_3673,N_3432,N_3593);
nand U3674 (N_3674,N_3475,N_3446);
xnor U3675 (N_3675,N_3547,N_3413);
and U3676 (N_3676,N_3461,N_3560);
nor U3677 (N_3677,N_3576,N_3564);
and U3678 (N_3678,N_3495,N_3463);
or U3679 (N_3679,N_3503,N_3518);
and U3680 (N_3680,N_3456,N_3409);
or U3681 (N_3681,N_3568,N_3527);
xor U3682 (N_3682,N_3529,N_3533);
xnor U3683 (N_3683,N_3480,N_3417);
and U3684 (N_3684,N_3554,N_3558);
xnor U3685 (N_3685,N_3536,N_3589);
xnor U3686 (N_3686,N_3470,N_3522);
nor U3687 (N_3687,N_3509,N_3599);
xnor U3688 (N_3688,N_3450,N_3591);
nand U3689 (N_3689,N_3411,N_3418);
nand U3690 (N_3690,N_3408,N_3501);
xor U3691 (N_3691,N_3575,N_3597);
nor U3692 (N_3692,N_3477,N_3542);
nand U3693 (N_3693,N_3481,N_3567);
nor U3694 (N_3694,N_3561,N_3400);
nand U3695 (N_3695,N_3449,N_3508);
xnor U3696 (N_3696,N_3479,N_3444);
or U3697 (N_3697,N_3421,N_3469);
nand U3698 (N_3698,N_3435,N_3453);
xnor U3699 (N_3699,N_3491,N_3549);
and U3700 (N_3700,N_3523,N_3475);
nand U3701 (N_3701,N_3524,N_3492);
or U3702 (N_3702,N_3409,N_3557);
and U3703 (N_3703,N_3435,N_3442);
or U3704 (N_3704,N_3441,N_3449);
and U3705 (N_3705,N_3422,N_3403);
nand U3706 (N_3706,N_3517,N_3427);
or U3707 (N_3707,N_3536,N_3414);
or U3708 (N_3708,N_3557,N_3428);
and U3709 (N_3709,N_3585,N_3570);
or U3710 (N_3710,N_3435,N_3455);
xor U3711 (N_3711,N_3596,N_3455);
nor U3712 (N_3712,N_3563,N_3579);
nor U3713 (N_3713,N_3459,N_3579);
nor U3714 (N_3714,N_3492,N_3597);
xor U3715 (N_3715,N_3544,N_3507);
xnor U3716 (N_3716,N_3517,N_3523);
nor U3717 (N_3717,N_3445,N_3400);
or U3718 (N_3718,N_3408,N_3476);
or U3719 (N_3719,N_3427,N_3430);
xnor U3720 (N_3720,N_3530,N_3418);
and U3721 (N_3721,N_3564,N_3479);
xnor U3722 (N_3722,N_3508,N_3435);
nor U3723 (N_3723,N_3456,N_3416);
or U3724 (N_3724,N_3572,N_3590);
and U3725 (N_3725,N_3423,N_3461);
xnor U3726 (N_3726,N_3538,N_3408);
xor U3727 (N_3727,N_3505,N_3513);
xnor U3728 (N_3728,N_3503,N_3496);
and U3729 (N_3729,N_3549,N_3483);
or U3730 (N_3730,N_3415,N_3405);
xnor U3731 (N_3731,N_3508,N_3509);
nor U3732 (N_3732,N_3538,N_3437);
xnor U3733 (N_3733,N_3421,N_3500);
or U3734 (N_3734,N_3505,N_3554);
xnor U3735 (N_3735,N_3573,N_3590);
nand U3736 (N_3736,N_3554,N_3408);
and U3737 (N_3737,N_3537,N_3565);
and U3738 (N_3738,N_3456,N_3432);
nor U3739 (N_3739,N_3437,N_3551);
nand U3740 (N_3740,N_3456,N_3414);
or U3741 (N_3741,N_3407,N_3541);
xor U3742 (N_3742,N_3473,N_3482);
nor U3743 (N_3743,N_3550,N_3435);
nand U3744 (N_3744,N_3574,N_3597);
nor U3745 (N_3745,N_3543,N_3528);
nand U3746 (N_3746,N_3441,N_3544);
and U3747 (N_3747,N_3402,N_3428);
nand U3748 (N_3748,N_3546,N_3537);
nor U3749 (N_3749,N_3479,N_3518);
or U3750 (N_3750,N_3423,N_3477);
xor U3751 (N_3751,N_3556,N_3440);
nand U3752 (N_3752,N_3462,N_3489);
and U3753 (N_3753,N_3521,N_3501);
xnor U3754 (N_3754,N_3468,N_3462);
or U3755 (N_3755,N_3533,N_3403);
or U3756 (N_3756,N_3470,N_3537);
or U3757 (N_3757,N_3560,N_3591);
and U3758 (N_3758,N_3445,N_3512);
and U3759 (N_3759,N_3497,N_3585);
nand U3760 (N_3760,N_3599,N_3435);
nor U3761 (N_3761,N_3485,N_3544);
or U3762 (N_3762,N_3441,N_3550);
or U3763 (N_3763,N_3523,N_3400);
nor U3764 (N_3764,N_3506,N_3591);
nor U3765 (N_3765,N_3574,N_3493);
xnor U3766 (N_3766,N_3545,N_3518);
or U3767 (N_3767,N_3471,N_3517);
nor U3768 (N_3768,N_3463,N_3479);
xor U3769 (N_3769,N_3568,N_3596);
nor U3770 (N_3770,N_3572,N_3576);
or U3771 (N_3771,N_3435,N_3552);
nand U3772 (N_3772,N_3521,N_3417);
nand U3773 (N_3773,N_3490,N_3453);
nand U3774 (N_3774,N_3590,N_3531);
nor U3775 (N_3775,N_3582,N_3581);
xnor U3776 (N_3776,N_3489,N_3481);
or U3777 (N_3777,N_3576,N_3493);
and U3778 (N_3778,N_3493,N_3419);
and U3779 (N_3779,N_3569,N_3522);
nand U3780 (N_3780,N_3524,N_3564);
or U3781 (N_3781,N_3552,N_3485);
or U3782 (N_3782,N_3482,N_3514);
or U3783 (N_3783,N_3537,N_3428);
nand U3784 (N_3784,N_3573,N_3422);
nand U3785 (N_3785,N_3516,N_3569);
nand U3786 (N_3786,N_3450,N_3472);
nand U3787 (N_3787,N_3425,N_3474);
xor U3788 (N_3788,N_3412,N_3477);
nor U3789 (N_3789,N_3446,N_3432);
and U3790 (N_3790,N_3464,N_3574);
nand U3791 (N_3791,N_3415,N_3593);
or U3792 (N_3792,N_3527,N_3468);
and U3793 (N_3793,N_3485,N_3422);
nand U3794 (N_3794,N_3553,N_3451);
nand U3795 (N_3795,N_3510,N_3434);
xor U3796 (N_3796,N_3591,N_3443);
nand U3797 (N_3797,N_3592,N_3420);
xnor U3798 (N_3798,N_3598,N_3432);
nor U3799 (N_3799,N_3545,N_3452);
or U3800 (N_3800,N_3794,N_3763);
and U3801 (N_3801,N_3739,N_3664);
nand U3802 (N_3802,N_3657,N_3781);
nand U3803 (N_3803,N_3643,N_3661);
nor U3804 (N_3804,N_3637,N_3716);
or U3805 (N_3805,N_3782,N_3662);
xnor U3806 (N_3806,N_3628,N_3747);
xnor U3807 (N_3807,N_3754,N_3721);
nor U3808 (N_3808,N_3713,N_3722);
and U3809 (N_3809,N_3609,N_3789);
xor U3810 (N_3810,N_3627,N_3697);
and U3811 (N_3811,N_3613,N_3792);
nand U3812 (N_3812,N_3788,N_3607);
xor U3813 (N_3813,N_3751,N_3614);
nor U3814 (N_3814,N_3731,N_3787);
xnor U3815 (N_3815,N_3785,N_3652);
xnor U3816 (N_3816,N_3798,N_3619);
and U3817 (N_3817,N_3645,N_3725);
and U3818 (N_3818,N_3603,N_3714);
and U3819 (N_3819,N_3755,N_3704);
and U3820 (N_3820,N_3771,N_3605);
and U3821 (N_3821,N_3633,N_3689);
xor U3822 (N_3822,N_3703,N_3783);
nand U3823 (N_3823,N_3799,N_3653);
nor U3824 (N_3824,N_3711,N_3659);
and U3825 (N_3825,N_3629,N_3730);
and U3826 (N_3826,N_3702,N_3793);
or U3827 (N_3827,N_3700,N_3655);
nand U3828 (N_3828,N_3620,N_3675);
xnor U3829 (N_3829,N_3669,N_3682);
xor U3830 (N_3830,N_3687,N_3737);
nor U3831 (N_3831,N_3705,N_3776);
nor U3832 (N_3832,N_3647,N_3724);
xnor U3833 (N_3833,N_3760,N_3750);
or U3834 (N_3834,N_3604,N_3624);
or U3835 (N_3835,N_3774,N_3630);
or U3836 (N_3836,N_3756,N_3676);
xor U3837 (N_3837,N_3727,N_3708);
nand U3838 (N_3838,N_3753,N_3752);
nand U3839 (N_3839,N_3728,N_3671);
or U3840 (N_3840,N_3601,N_3644);
xor U3841 (N_3841,N_3690,N_3767);
or U3842 (N_3842,N_3608,N_3717);
nand U3843 (N_3843,N_3648,N_3762);
nor U3844 (N_3844,N_3636,N_3660);
nand U3845 (N_3845,N_3635,N_3735);
nand U3846 (N_3846,N_3765,N_3759);
and U3847 (N_3847,N_3694,N_3695);
and U3848 (N_3848,N_3748,N_3723);
or U3849 (N_3849,N_3606,N_3769);
and U3850 (N_3850,N_3761,N_3612);
and U3851 (N_3851,N_3663,N_3733);
and U3852 (N_3852,N_3784,N_3670);
nand U3853 (N_3853,N_3691,N_3631);
xor U3854 (N_3854,N_3642,N_3678);
nand U3855 (N_3855,N_3600,N_3649);
or U3856 (N_3856,N_3623,N_3651);
nor U3857 (N_3857,N_3621,N_3681);
nor U3858 (N_3858,N_3720,N_3715);
nor U3859 (N_3859,N_3791,N_3786);
or U3860 (N_3860,N_3683,N_3706);
xor U3861 (N_3861,N_3618,N_3790);
nor U3862 (N_3862,N_3743,N_3672);
or U3863 (N_3863,N_3656,N_3658);
nor U3864 (N_3864,N_3738,N_3732);
and U3865 (N_3865,N_3746,N_3638);
nor U3866 (N_3866,N_3734,N_3712);
xnor U3867 (N_3867,N_3742,N_3780);
nand U3868 (N_3868,N_3654,N_3797);
and U3869 (N_3869,N_3772,N_3709);
xnor U3870 (N_3870,N_3680,N_3667);
nor U3871 (N_3871,N_3736,N_3778);
nand U3872 (N_3872,N_3749,N_3779);
xnor U3873 (N_3873,N_3679,N_3745);
nand U3874 (N_3874,N_3611,N_3701);
or U3875 (N_3875,N_3622,N_3646);
or U3876 (N_3876,N_3718,N_3685);
nor U3877 (N_3877,N_3764,N_3773);
nor U3878 (N_3878,N_3770,N_3796);
or U3879 (N_3879,N_3674,N_3777);
or U3880 (N_3880,N_3699,N_3615);
xor U3881 (N_3881,N_3684,N_3626);
xor U3882 (N_3882,N_3666,N_3696);
or U3883 (N_3883,N_3610,N_3625);
or U3884 (N_3884,N_3693,N_3650);
and U3885 (N_3885,N_3719,N_3665);
or U3886 (N_3886,N_3686,N_3757);
nor U3887 (N_3887,N_3616,N_3775);
xor U3888 (N_3888,N_3640,N_3688);
and U3889 (N_3889,N_3677,N_3795);
and U3890 (N_3890,N_3768,N_3729);
nor U3891 (N_3891,N_3641,N_3673);
nand U3892 (N_3892,N_3766,N_3692);
xor U3893 (N_3893,N_3698,N_3710);
nor U3894 (N_3894,N_3707,N_3602);
or U3895 (N_3895,N_3632,N_3668);
or U3896 (N_3896,N_3639,N_3634);
nand U3897 (N_3897,N_3740,N_3617);
or U3898 (N_3898,N_3758,N_3744);
and U3899 (N_3899,N_3741,N_3726);
and U3900 (N_3900,N_3743,N_3620);
nand U3901 (N_3901,N_3780,N_3644);
and U3902 (N_3902,N_3712,N_3713);
or U3903 (N_3903,N_3729,N_3750);
nand U3904 (N_3904,N_3618,N_3623);
and U3905 (N_3905,N_3699,N_3713);
nand U3906 (N_3906,N_3680,N_3764);
nor U3907 (N_3907,N_3701,N_3735);
xnor U3908 (N_3908,N_3666,N_3687);
xnor U3909 (N_3909,N_3766,N_3695);
xnor U3910 (N_3910,N_3766,N_3606);
or U3911 (N_3911,N_3790,N_3739);
nand U3912 (N_3912,N_3745,N_3647);
xnor U3913 (N_3913,N_3710,N_3677);
nor U3914 (N_3914,N_3695,N_3602);
or U3915 (N_3915,N_3713,N_3613);
and U3916 (N_3916,N_3721,N_3621);
or U3917 (N_3917,N_3745,N_3648);
xnor U3918 (N_3918,N_3728,N_3778);
nor U3919 (N_3919,N_3799,N_3627);
and U3920 (N_3920,N_3648,N_3657);
and U3921 (N_3921,N_3605,N_3675);
and U3922 (N_3922,N_3628,N_3741);
xor U3923 (N_3923,N_3652,N_3775);
nor U3924 (N_3924,N_3717,N_3730);
and U3925 (N_3925,N_3666,N_3750);
xor U3926 (N_3926,N_3717,N_3701);
nand U3927 (N_3927,N_3713,N_3730);
and U3928 (N_3928,N_3735,N_3641);
nand U3929 (N_3929,N_3621,N_3730);
nor U3930 (N_3930,N_3764,N_3668);
nor U3931 (N_3931,N_3688,N_3609);
and U3932 (N_3932,N_3677,N_3757);
and U3933 (N_3933,N_3730,N_3668);
or U3934 (N_3934,N_3707,N_3658);
xor U3935 (N_3935,N_3781,N_3626);
and U3936 (N_3936,N_3786,N_3641);
xnor U3937 (N_3937,N_3763,N_3691);
nand U3938 (N_3938,N_3708,N_3633);
xnor U3939 (N_3939,N_3698,N_3697);
xnor U3940 (N_3940,N_3602,N_3671);
or U3941 (N_3941,N_3784,N_3680);
nor U3942 (N_3942,N_3638,N_3712);
or U3943 (N_3943,N_3665,N_3704);
or U3944 (N_3944,N_3744,N_3619);
xnor U3945 (N_3945,N_3628,N_3777);
or U3946 (N_3946,N_3793,N_3602);
nand U3947 (N_3947,N_3700,N_3718);
or U3948 (N_3948,N_3651,N_3606);
nor U3949 (N_3949,N_3602,N_3636);
nor U3950 (N_3950,N_3729,N_3695);
nand U3951 (N_3951,N_3626,N_3790);
nor U3952 (N_3952,N_3616,N_3742);
and U3953 (N_3953,N_3733,N_3755);
or U3954 (N_3954,N_3763,N_3721);
xnor U3955 (N_3955,N_3618,N_3763);
and U3956 (N_3956,N_3659,N_3759);
xor U3957 (N_3957,N_3736,N_3665);
nand U3958 (N_3958,N_3720,N_3744);
or U3959 (N_3959,N_3623,N_3773);
and U3960 (N_3960,N_3607,N_3734);
nor U3961 (N_3961,N_3701,N_3718);
and U3962 (N_3962,N_3615,N_3648);
or U3963 (N_3963,N_3766,N_3649);
nand U3964 (N_3964,N_3709,N_3614);
xor U3965 (N_3965,N_3617,N_3786);
or U3966 (N_3966,N_3718,N_3620);
nor U3967 (N_3967,N_3651,N_3668);
xnor U3968 (N_3968,N_3762,N_3725);
nand U3969 (N_3969,N_3603,N_3638);
or U3970 (N_3970,N_3755,N_3762);
and U3971 (N_3971,N_3736,N_3686);
xnor U3972 (N_3972,N_3799,N_3791);
nand U3973 (N_3973,N_3692,N_3655);
or U3974 (N_3974,N_3653,N_3685);
nor U3975 (N_3975,N_3656,N_3790);
xnor U3976 (N_3976,N_3773,N_3688);
nor U3977 (N_3977,N_3662,N_3676);
nand U3978 (N_3978,N_3781,N_3748);
or U3979 (N_3979,N_3764,N_3600);
nor U3980 (N_3980,N_3644,N_3729);
nor U3981 (N_3981,N_3648,N_3726);
and U3982 (N_3982,N_3602,N_3784);
or U3983 (N_3983,N_3794,N_3629);
nor U3984 (N_3984,N_3623,N_3729);
nor U3985 (N_3985,N_3672,N_3611);
and U3986 (N_3986,N_3627,N_3606);
or U3987 (N_3987,N_3737,N_3698);
or U3988 (N_3988,N_3730,N_3678);
nor U3989 (N_3989,N_3720,N_3611);
and U3990 (N_3990,N_3714,N_3679);
and U3991 (N_3991,N_3717,N_3790);
nand U3992 (N_3992,N_3717,N_3757);
and U3993 (N_3993,N_3715,N_3649);
or U3994 (N_3994,N_3726,N_3699);
or U3995 (N_3995,N_3678,N_3747);
nand U3996 (N_3996,N_3647,N_3706);
and U3997 (N_3997,N_3750,N_3743);
nand U3998 (N_3998,N_3681,N_3769);
xor U3999 (N_3999,N_3607,N_3708);
nor U4000 (N_4000,N_3876,N_3920);
nand U4001 (N_4001,N_3861,N_3870);
and U4002 (N_4002,N_3814,N_3896);
nor U4003 (N_4003,N_3985,N_3924);
nor U4004 (N_4004,N_3986,N_3815);
or U4005 (N_4005,N_3973,N_3913);
xor U4006 (N_4006,N_3840,N_3884);
and U4007 (N_4007,N_3858,N_3944);
and U4008 (N_4008,N_3965,N_3975);
and U4009 (N_4009,N_3830,N_3904);
nand U4010 (N_4010,N_3889,N_3871);
nand U4011 (N_4011,N_3996,N_3885);
nor U4012 (N_4012,N_3992,N_3969);
nand U4013 (N_4013,N_3911,N_3857);
and U4014 (N_4014,N_3988,N_3955);
and U4015 (N_4015,N_3806,N_3898);
nand U4016 (N_4016,N_3917,N_3802);
and U4017 (N_4017,N_3964,N_3923);
xor U4018 (N_4018,N_3895,N_3853);
nand U4019 (N_4019,N_3843,N_3834);
or U4020 (N_4020,N_3966,N_3852);
nor U4021 (N_4021,N_3831,N_3872);
xor U4022 (N_4022,N_3844,N_3998);
and U4023 (N_4023,N_3826,N_3954);
or U4024 (N_4024,N_3932,N_3842);
nor U4025 (N_4025,N_3981,N_3801);
xor U4026 (N_4026,N_3945,N_3820);
nand U4027 (N_4027,N_3883,N_3971);
and U4028 (N_4028,N_3894,N_3899);
xnor U4029 (N_4029,N_3990,N_3929);
and U4030 (N_4030,N_3846,N_3869);
xor U4031 (N_4031,N_3963,N_3914);
or U4032 (N_4032,N_3850,N_3949);
xnor U4033 (N_4033,N_3999,N_3823);
xor U4034 (N_4034,N_3978,N_3866);
and U4035 (N_4035,N_3951,N_3931);
and U4036 (N_4036,N_3824,N_3910);
and U4037 (N_4037,N_3811,N_3926);
or U4038 (N_4038,N_3908,N_3817);
xor U4039 (N_4039,N_3822,N_3841);
nand U4040 (N_4040,N_3982,N_3912);
xor U4041 (N_4041,N_3859,N_3995);
and U4042 (N_4042,N_3836,N_3915);
xnor U4043 (N_4043,N_3886,N_3902);
nor U4044 (N_4044,N_3854,N_3979);
or U4045 (N_4045,N_3942,N_3862);
xor U4046 (N_4046,N_3903,N_3930);
xor U4047 (N_4047,N_3891,N_3922);
xnor U4048 (N_4048,N_3934,N_3882);
or U4049 (N_4049,N_3860,N_3878);
nor U4050 (N_4050,N_3959,N_3827);
or U4051 (N_4051,N_3909,N_3893);
nand U4052 (N_4052,N_3984,N_3938);
nand U4053 (N_4053,N_3993,N_3851);
or U4054 (N_4054,N_3818,N_3863);
nand U4055 (N_4055,N_3936,N_3808);
and U4056 (N_4056,N_3807,N_3897);
nor U4057 (N_4057,N_3901,N_3928);
nor U4058 (N_4058,N_3812,N_3989);
nand U4059 (N_4059,N_3968,N_3875);
nor U4060 (N_4060,N_3868,N_3848);
xnor U4061 (N_4061,N_3948,N_3877);
nor U4062 (N_4062,N_3892,N_3864);
nor U4063 (N_4063,N_3977,N_3916);
and U4064 (N_4064,N_3974,N_3907);
and U4065 (N_4065,N_3810,N_3967);
and U4066 (N_4066,N_3970,N_3925);
and U4067 (N_4067,N_3941,N_3813);
or U4068 (N_4068,N_3957,N_3900);
and U4069 (N_4069,N_3953,N_3919);
and U4070 (N_4070,N_3879,N_3888);
or U4071 (N_4071,N_3956,N_3839);
and U4072 (N_4072,N_3927,N_3890);
nand U4073 (N_4073,N_3994,N_3983);
and U4074 (N_4074,N_3825,N_3943);
and U4075 (N_4075,N_3873,N_3952);
nand U4076 (N_4076,N_3947,N_3935);
xor U4077 (N_4077,N_3991,N_3906);
xor U4078 (N_4078,N_3865,N_3921);
or U4079 (N_4079,N_3855,N_3980);
xor U4080 (N_4080,N_3962,N_3805);
and U4081 (N_4081,N_3958,N_3880);
nand U4082 (N_4082,N_3939,N_3918);
nor U4083 (N_4083,N_3804,N_3881);
nor U4084 (N_4084,N_3946,N_3856);
xor U4085 (N_4085,N_3960,N_3835);
nand U4086 (N_4086,N_3933,N_3937);
and U4087 (N_4087,N_3837,N_3816);
nor U4088 (N_4088,N_3950,N_3976);
and U4089 (N_4089,N_3809,N_3972);
nand U4090 (N_4090,N_3819,N_3905);
nand U4091 (N_4091,N_3803,N_3961);
and U4092 (N_4092,N_3987,N_3874);
or U4093 (N_4093,N_3849,N_3940);
or U4094 (N_4094,N_3832,N_3800);
and U4095 (N_4095,N_3828,N_3821);
nand U4096 (N_4096,N_3887,N_3997);
nor U4097 (N_4097,N_3845,N_3867);
and U4098 (N_4098,N_3833,N_3847);
or U4099 (N_4099,N_3829,N_3838);
and U4100 (N_4100,N_3871,N_3858);
and U4101 (N_4101,N_3886,N_3830);
or U4102 (N_4102,N_3837,N_3933);
and U4103 (N_4103,N_3811,N_3829);
and U4104 (N_4104,N_3945,N_3872);
nor U4105 (N_4105,N_3954,N_3956);
and U4106 (N_4106,N_3816,N_3998);
and U4107 (N_4107,N_3969,N_3844);
xor U4108 (N_4108,N_3928,N_3833);
or U4109 (N_4109,N_3933,N_3850);
and U4110 (N_4110,N_3987,N_3960);
and U4111 (N_4111,N_3985,N_3967);
or U4112 (N_4112,N_3823,N_3826);
and U4113 (N_4113,N_3855,N_3823);
nor U4114 (N_4114,N_3918,N_3934);
nand U4115 (N_4115,N_3923,N_3807);
nand U4116 (N_4116,N_3934,N_3822);
nand U4117 (N_4117,N_3874,N_3941);
or U4118 (N_4118,N_3837,N_3917);
and U4119 (N_4119,N_3824,N_3812);
and U4120 (N_4120,N_3880,N_3928);
nor U4121 (N_4121,N_3894,N_3968);
xnor U4122 (N_4122,N_3981,N_3867);
nand U4123 (N_4123,N_3869,N_3994);
nand U4124 (N_4124,N_3806,N_3999);
nand U4125 (N_4125,N_3918,N_3870);
nor U4126 (N_4126,N_3873,N_3980);
nand U4127 (N_4127,N_3974,N_3806);
nand U4128 (N_4128,N_3839,N_3806);
xnor U4129 (N_4129,N_3968,N_3896);
and U4130 (N_4130,N_3846,N_3818);
nor U4131 (N_4131,N_3936,N_3872);
or U4132 (N_4132,N_3919,N_3875);
nand U4133 (N_4133,N_3913,N_3814);
nand U4134 (N_4134,N_3946,N_3993);
nand U4135 (N_4135,N_3932,N_3885);
xnor U4136 (N_4136,N_3921,N_3958);
or U4137 (N_4137,N_3925,N_3932);
or U4138 (N_4138,N_3871,N_3854);
and U4139 (N_4139,N_3973,N_3938);
and U4140 (N_4140,N_3977,N_3878);
xnor U4141 (N_4141,N_3933,N_3897);
nand U4142 (N_4142,N_3903,N_3853);
or U4143 (N_4143,N_3938,N_3842);
xnor U4144 (N_4144,N_3810,N_3977);
or U4145 (N_4145,N_3801,N_3866);
xnor U4146 (N_4146,N_3807,N_3823);
or U4147 (N_4147,N_3834,N_3951);
xnor U4148 (N_4148,N_3863,N_3973);
nand U4149 (N_4149,N_3965,N_3905);
and U4150 (N_4150,N_3905,N_3884);
xor U4151 (N_4151,N_3909,N_3825);
or U4152 (N_4152,N_3877,N_3896);
nor U4153 (N_4153,N_3848,N_3832);
and U4154 (N_4154,N_3982,N_3981);
xnor U4155 (N_4155,N_3840,N_3912);
xnor U4156 (N_4156,N_3855,N_3973);
or U4157 (N_4157,N_3833,N_3933);
nand U4158 (N_4158,N_3862,N_3907);
or U4159 (N_4159,N_3807,N_3892);
nor U4160 (N_4160,N_3868,N_3893);
or U4161 (N_4161,N_3907,N_3965);
nand U4162 (N_4162,N_3814,N_3824);
xor U4163 (N_4163,N_3962,N_3814);
or U4164 (N_4164,N_3958,N_3970);
xor U4165 (N_4165,N_3826,N_3987);
nand U4166 (N_4166,N_3935,N_3927);
xor U4167 (N_4167,N_3830,N_3991);
nor U4168 (N_4168,N_3862,N_3922);
and U4169 (N_4169,N_3939,N_3920);
and U4170 (N_4170,N_3882,N_3983);
or U4171 (N_4171,N_3967,N_3938);
nor U4172 (N_4172,N_3875,N_3928);
and U4173 (N_4173,N_3897,N_3829);
xnor U4174 (N_4174,N_3865,N_3829);
or U4175 (N_4175,N_3905,N_3999);
xnor U4176 (N_4176,N_3882,N_3924);
xor U4177 (N_4177,N_3806,N_3844);
nor U4178 (N_4178,N_3915,N_3875);
or U4179 (N_4179,N_3860,N_3911);
nand U4180 (N_4180,N_3988,N_3805);
and U4181 (N_4181,N_3852,N_3932);
nand U4182 (N_4182,N_3948,N_3990);
nor U4183 (N_4183,N_3962,N_3893);
nand U4184 (N_4184,N_3860,N_3953);
nor U4185 (N_4185,N_3938,N_3885);
nand U4186 (N_4186,N_3944,N_3936);
xnor U4187 (N_4187,N_3812,N_3902);
nand U4188 (N_4188,N_3869,N_3808);
nor U4189 (N_4189,N_3820,N_3983);
nand U4190 (N_4190,N_3922,N_3957);
nand U4191 (N_4191,N_3842,N_3837);
nand U4192 (N_4192,N_3818,N_3972);
nor U4193 (N_4193,N_3807,N_3874);
nand U4194 (N_4194,N_3866,N_3914);
and U4195 (N_4195,N_3906,N_3860);
nor U4196 (N_4196,N_3884,N_3830);
nand U4197 (N_4197,N_3968,N_3980);
nand U4198 (N_4198,N_3886,N_3816);
and U4199 (N_4199,N_3898,N_3909);
and U4200 (N_4200,N_4140,N_4100);
nor U4201 (N_4201,N_4044,N_4060);
xnor U4202 (N_4202,N_4025,N_4030);
nor U4203 (N_4203,N_4127,N_4155);
xor U4204 (N_4204,N_4034,N_4046);
or U4205 (N_4205,N_4033,N_4063);
or U4206 (N_4206,N_4028,N_4106);
nor U4207 (N_4207,N_4168,N_4075);
or U4208 (N_4208,N_4066,N_4018);
and U4209 (N_4209,N_4058,N_4142);
nor U4210 (N_4210,N_4143,N_4072);
nand U4211 (N_4211,N_4111,N_4029);
nand U4212 (N_4212,N_4012,N_4045);
or U4213 (N_4213,N_4015,N_4067);
or U4214 (N_4214,N_4107,N_4059);
or U4215 (N_4215,N_4164,N_4102);
xnor U4216 (N_4216,N_4192,N_4162);
or U4217 (N_4217,N_4176,N_4190);
nor U4218 (N_4218,N_4126,N_4198);
nor U4219 (N_4219,N_4175,N_4180);
nand U4220 (N_4220,N_4091,N_4119);
nand U4221 (N_4221,N_4146,N_4123);
nand U4222 (N_4222,N_4195,N_4170);
or U4223 (N_4223,N_4035,N_4154);
xnor U4224 (N_4224,N_4006,N_4010);
nor U4225 (N_4225,N_4054,N_4014);
nand U4226 (N_4226,N_4134,N_4169);
xor U4227 (N_4227,N_4062,N_4113);
nor U4228 (N_4228,N_4101,N_4189);
and U4229 (N_4229,N_4158,N_4160);
nor U4230 (N_4230,N_4116,N_4019);
nor U4231 (N_4231,N_4112,N_4009);
and U4232 (N_4232,N_4088,N_4089);
or U4233 (N_4233,N_4026,N_4157);
nand U4234 (N_4234,N_4159,N_4078);
or U4235 (N_4235,N_4007,N_4120);
and U4236 (N_4236,N_4086,N_4039);
and U4237 (N_4237,N_4103,N_4055);
or U4238 (N_4238,N_4027,N_4031);
or U4239 (N_4239,N_4183,N_4108);
nor U4240 (N_4240,N_4130,N_4191);
or U4241 (N_4241,N_4016,N_4070);
nand U4242 (N_4242,N_4095,N_4185);
xor U4243 (N_4243,N_4093,N_4109);
and U4244 (N_4244,N_4133,N_4068);
and U4245 (N_4245,N_4177,N_4043);
nor U4246 (N_4246,N_4197,N_4051);
or U4247 (N_4247,N_4135,N_4056);
xor U4248 (N_4248,N_4121,N_4129);
and U4249 (N_4249,N_4124,N_4136);
nand U4250 (N_4250,N_4047,N_4079);
nand U4251 (N_4251,N_4053,N_4057);
and U4252 (N_4252,N_4132,N_4110);
or U4253 (N_4253,N_4000,N_4049);
or U4254 (N_4254,N_4005,N_4147);
nand U4255 (N_4255,N_4090,N_4115);
nand U4256 (N_4256,N_4167,N_4117);
xnor U4257 (N_4257,N_4036,N_4144);
or U4258 (N_4258,N_4024,N_4118);
and U4259 (N_4259,N_4153,N_4064);
nand U4260 (N_4260,N_4184,N_4181);
nor U4261 (N_4261,N_4122,N_4131);
nor U4262 (N_4262,N_4125,N_4004);
nor U4263 (N_4263,N_4077,N_4148);
or U4264 (N_4264,N_4071,N_4069);
or U4265 (N_4265,N_4179,N_4186);
xor U4266 (N_4266,N_4073,N_4032);
xnor U4267 (N_4267,N_4194,N_4038);
nand U4268 (N_4268,N_4161,N_4023);
or U4269 (N_4269,N_4096,N_4137);
nor U4270 (N_4270,N_4080,N_4040);
nand U4271 (N_4271,N_4017,N_4022);
xor U4272 (N_4272,N_4082,N_4138);
nand U4273 (N_4273,N_4002,N_4196);
nand U4274 (N_4274,N_4052,N_4182);
nor U4275 (N_4275,N_4152,N_4061);
nand U4276 (N_4276,N_4074,N_4065);
nor U4277 (N_4277,N_4188,N_4174);
and U4278 (N_4278,N_4084,N_4081);
nor U4279 (N_4279,N_4163,N_4139);
xor U4280 (N_4280,N_4105,N_4001);
nand U4281 (N_4281,N_4149,N_4150);
nor U4282 (N_4282,N_4041,N_4156);
or U4283 (N_4283,N_4011,N_4172);
nand U4284 (N_4284,N_4141,N_4128);
or U4285 (N_4285,N_4099,N_4173);
or U4286 (N_4286,N_4166,N_4165);
or U4287 (N_4287,N_4104,N_4021);
and U4288 (N_4288,N_4050,N_4042);
or U4289 (N_4289,N_4087,N_4097);
nand U4290 (N_4290,N_4114,N_4094);
nand U4291 (N_4291,N_4092,N_4178);
xnor U4292 (N_4292,N_4008,N_4013);
nor U4293 (N_4293,N_4076,N_4145);
nor U4294 (N_4294,N_4199,N_4037);
and U4295 (N_4295,N_4098,N_4083);
nor U4296 (N_4296,N_4003,N_4187);
nand U4297 (N_4297,N_4151,N_4085);
nor U4298 (N_4298,N_4020,N_4171);
and U4299 (N_4299,N_4193,N_4048);
nand U4300 (N_4300,N_4172,N_4122);
nand U4301 (N_4301,N_4096,N_4017);
nor U4302 (N_4302,N_4053,N_4192);
nand U4303 (N_4303,N_4110,N_4116);
nand U4304 (N_4304,N_4100,N_4191);
nor U4305 (N_4305,N_4130,N_4029);
and U4306 (N_4306,N_4055,N_4007);
or U4307 (N_4307,N_4048,N_4197);
or U4308 (N_4308,N_4027,N_4171);
nor U4309 (N_4309,N_4114,N_4104);
nand U4310 (N_4310,N_4039,N_4115);
or U4311 (N_4311,N_4037,N_4071);
and U4312 (N_4312,N_4109,N_4139);
nor U4313 (N_4313,N_4104,N_4164);
nor U4314 (N_4314,N_4098,N_4189);
and U4315 (N_4315,N_4124,N_4083);
nor U4316 (N_4316,N_4141,N_4011);
nand U4317 (N_4317,N_4165,N_4022);
or U4318 (N_4318,N_4105,N_4041);
nand U4319 (N_4319,N_4052,N_4146);
or U4320 (N_4320,N_4008,N_4102);
nand U4321 (N_4321,N_4072,N_4063);
or U4322 (N_4322,N_4106,N_4134);
and U4323 (N_4323,N_4144,N_4070);
nor U4324 (N_4324,N_4063,N_4094);
or U4325 (N_4325,N_4113,N_4079);
nand U4326 (N_4326,N_4009,N_4055);
nand U4327 (N_4327,N_4026,N_4138);
nand U4328 (N_4328,N_4006,N_4199);
nor U4329 (N_4329,N_4100,N_4097);
xor U4330 (N_4330,N_4143,N_4122);
xor U4331 (N_4331,N_4149,N_4160);
or U4332 (N_4332,N_4145,N_4114);
nor U4333 (N_4333,N_4029,N_4092);
nand U4334 (N_4334,N_4011,N_4026);
xnor U4335 (N_4335,N_4077,N_4079);
nor U4336 (N_4336,N_4127,N_4198);
and U4337 (N_4337,N_4192,N_4050);
and U4338 (N_4338,N_4170,N_4073);
and U4339 (N_4339,N_4140,N_4171);
xor U4340 (N_4340,N_4128,N_4185);
nand U4341 (N_4341,N_4070,N_4103);
and U4342 (N_4342,N_4108,N_4123);
nand U4343 (N_4343,N_4143,N_4168);
nor U4344 (N_4344,N_4167,N_4186);
and U4345 (N_4345,N_4002,N_4006);
xnor U4346 (N_4346,N_4053,N_4044);
or U4347 (N_4347,N_4047,N_4010);
xor U4348 (N_4348,N_4144,N_4182);
and U4349 (N_4349,N_4144,N_4138);
nand U4350 (N_4350,N_4028,N_4006);
nand U4351 (N_4351,N_4156,N_4057);
nand U4352 (N_4352,N_4024,N_4115);
nand U4353 (N_4353,N_4170,N_4005);
nor U4354 (N_4354,N_4192,N_4123);
or U4355 (N_4355,N_4045,N_4069);
or U4356 (N_4356,N_4002,N_4123);
and U4357 (N_4357,N_4177,N_4090);
and U4358 (N_4358,N_4088,N_4099);
nand U4359 (N_4359,N_4029,N_4146);
and U4360 (N_4360,N_4113,N_4082);
nor U4361 (N_4361,N_4067,N_4193);
or U4362 (N_4362,N_4091,N_4114);
or U4363 (N_4363,N_4150,N_4138);
nand U4364 (N_4364,N_4026,N_4196);
or U4365 (N_4365,N_4060,N_4038);
xnor U4366 (N_4366,N_4090,N_4184);
nor U4367 (N_4367,N_4089,N_4077);
and U4368 (N_4368,N_4003,N_4011);
and U4369 (N_4369,N_4126,N_4049);
nor U4370 (N_4370,N_4108,N_4004);
nor U4371 (N_4371,N_4027,N_4053);
nor U4372 (N_4372,N_4027,N_4047);
nand U4373 (N_4373,N_4019,N_4100);
and U4374 (N_4374,N_4036,N_4073);
nand U4375 (N_4375,N_4021,N_4005);
and U4376 (N_4376,N_4035,N_4088);
nor U4377 (N_4377,N_4073,N_4035);
nor U4378 (N_4378,N_4135,N_4178);
xor U4379 (N_4379,N_4028,N_4036);
and U4380 (N_4380,N_4002,N_4115);
nor U4381 (N_4381,N_4085,N_4070);
nand U4382 (N_4382,N_4149,N_4084);
xnor U4383 (N_4383,N_4094,N_4033);
and U4384 (N_4384,N_4176,N_4083);
nor U4385 (N_4385,N_4067,N_4102);
xor U4386 (N_4386,N_4139,N_4154);
and U4387 (N_4387,N_4045,N_4146);
or U4388 (N_4388,N_4025,N_4184);
or U4389 (N_4389,N_4137,N_4091);
xor U4390 (N_4390,N_4072,N_4137);
nor U4391 (N_4391,N_4190,N_4033);
nor U4392 (N_4392,N_4072,N_4003);
xor U4393 (N_4393,N_4180,N_4093);
nor U4394 (N_4394,N_4108,N_4026);
nand U4395 (N_4395,N_4040,N_4068);
nand U4396 (N_4396,N_4025,N_4087);
nand U4397 (N_4397,N_4074,N_4183);
or U4398 (N_4398,N_4140,N_4152);
xor U4399 (N_4399,N_4181,N_4057);
and U4400 (N_4400,N_4383,N_4399);
or U4401 (N_4401,N_4361,N_4259);
and U4402 (N_4402,N_4376,N_4203);
xnor U4403 (N_4403,N_4229,N_4318);
or U4404 (N_4404,N_4336,N_4366);
nand U4405 (N_4405,N_4202,N_4211);
xor U4406 (N_4406,N_4220,N_4377);
nor U4407 (N_4407,N_4360,N_4291);
nand U4408 (N_4408,N_4289,N_4260);
and U4409 (N_4409,N_4236,N_4321);
or U4410 (N_4410,N_4276,N_4355);
xnor U4411 (N_4411,N_4219,N_4392);
or U4412 (N_4412,N_4348,N_4325);
xnor U4413 (N_4413,N_4396,N_4225);
or U4414 (N_4414,N_4226,N_4232);
and U4415 (N_4415,N_4333,N_4313);
and U4416 (N_4416,N_4239,N_4300);
and U4417 (N_4417,N_4204,N_4246);
nor U4418 (N_4418,N_4372,N_4322);
or U4419 (N_4419,N_4307,N_4279);
nor U4420 (N_4420,N_4359,N_4310);
nor U4421 (N_4421,N_4234,N_4273);
nand U4422 (N_4422,N_4367,N_4268);
nor U4423 (N_4423,N_4212,N_4323);
nand U4424 (N_4424,N_4255,N_4341);
or U4425 (N_4425,N_4337,N_4274);
and U4426 (N_4426,N_4314,N_4262);
nand U4427 (N_4427,N_4209,N_4328);
and U4428 (N_4428,N_4356,N_4213);
nand U4429 (N_4429,N_4252,N_4292);
nand U4430 (N_4430,N_4309,N_4240);
nor U4431 (N_4431,N_4388,N_4261);
nor U4432 (N_4432,N_4216,N_4210);
and U4433 (N_4433,N_4285,N_4277);
nand U4434 (N_4434,N_4271,N_4208);
xnor U4435 (N_4435,N_4218,N_4228);
and U4436 (N_4436,N_4231,N_4339);
and U4437 (N_4437,N_4223,N_4242);
xnor U4438 (N_4438,N_4342,N_4389);
nor U4439 (N_4439,N_4296,N_4230);
nor U4440 (N_4440,N_4283,N_4397);
or U4441 (N_4441,N_4326,N_4329);
xor U4442 (N_4442,N_4264,N_4272);
nor U4443 (N_4443,N_4354,N_4373);
xor U4444 (N_4444,N_4308,N_4381);
nor U4445 (N_4445,N_4254,N_4221);
xnor U4446 (N_4446,N_4269,N_4374);
nor U4447 (N_4447,N_4335,N_4351);
nand U4448 (N_4448,N_4304,N_4334);
nor U4449 (N_4449,N_4306,N_4350);
xor U4450 (N_4450,N_4345,N_4298);
nor U4451 (N_4451,N_4244,N_4340);
and U4452 (N_4452,N_4214,N_4281);
nand U4453 (N_4453,N_4352,N_4257);
nor U4454 (N_4454,N_4235,N_4245);
or U4455 (N_4455,N_4327,N_4284);
nand U4456 (N_4456,N_4275,N_4349);
or U4457 (N_4457,N_4287,N_4302);
and U4458 (N_4458,N_4294,N_4398);
xnor U4459 (N_4459,N_4247,N_4295);
and U4460 (N_4460,N_4293,N_4286);
xor U4461 (N_4461,N_4280,N_4370);
xor U4462 (N_4462,N_4251,N_4332);
or U4463 (N_4463,N_4394,N_4317);
or U4464 (N_4464,N_4200,N_4311);
and U4465 (N_4465,N_4353,N_4201);
or U4466 (N_4466,N_4324,N_4331);
or U4467 (N_4467,N_4303,N_4364);
xnor U4468 (N_4468,N_4344,N_4362);
and U4469 (N_4469,N_4206,N_4258);
xor U4470 (N_4470,N_4301,N_4267);
nand U4471 (N_4471,N_4358,N_4363);
xnor U4472 (N_4472,N_4316,N_4346);
nor U4473 (N_4473,N_4343,N_4369);
or U4474 (N_4474,N_4215,N_4266);
xor U4475 (N_4475,N_4393,N_4238);
xor U4476 (N_4476,N_4385,N_4305);
and U4477 (N_4477,N_4379,N_4384);
and U4478 (N_4478,N_4391,N_4256);
nor U4479 (N_4479,N_4222,N_4382);
xnor U4480 (N_4480,N_4338,N_4288);
xnor U4481 (N_4481,N_4319,N_4375);
and U4482 (N_4482,N_4250,N_4320);
or U4483 (N_4483,N_4270,N_4368);
nand U4484 (N_4484,N_4227,N_4249);
nand U4485 (N_4485,N_4387,N_4371);
or U4486 (N_4486,N_4312,N_4207);
or U4487 (N_4487,N_4330,N_4365);
and U4488 (N_4488,N_4205,N_4253);
nand U4489 (N_4489,N_4297,N_4357);
nand U4490 (N_4490,N_4217,N_4395);
nor U4491 (N_4491,N_4386,N_4233);
nand U4492 (N_4492,N_4380,N_4390);
nor U4493 (N_4493,N_4315,N_4237);
or U4494 (N_4494,N_4378,N_4265);
nor U4495 (N_4495,N_4263,N_4299);
xnor U4496 (N_4496,N_4243,N_4224);
nor U4497 (N_4497,N_4290,N_4347);
and U4498 (N_4498,N_4278,N_4241);
nor U4499 (N_4499,N_4248,N_4282);
nand U4500 (N_4500,N_4220,N_4351);
xnor U4501 (N_4501,N_4364,N_4339);
nor U4502 (N_4502,N_4314,N_4214);
and U4503 (N_4503,N_4389,N_4328);
xnor U4504 (N_4504,N_4363,N_4329);
xnor U4505 (N_4505,N_4200,N_4263);
or U4506 (N_4506,N_4268,N_4205);
and U4507 (N_4507,N_4345,N_4337);
and U4508 (N_4508,N_4324,N_4325);
nor U4509 (N_4509,N_4375,N_4233);
nor U4510 (N_4510,N_4246,N_4387);
and U4511 (N_4511,N_4240,N_4290);
nand U4512 (N_4512,N_4321,N_4288);
nand U4513 (N_4513,N_4331,N_4261);
xnor U4514 (N_4514,N_4350,N_4340);
nand U4515 (N_4515,N_4378,N_4211);
xnor U4516 (N_4516,N_4291,N_4359);
nor U4517 (N_4517,N_4294,N_4256);
nor U4518 (N_4518,N_4271,N_4280);
nand U4519 (N_4519,N_4235,N_4210);
nand U4520 (N_4520,N_4336,N_4324);
and U4521 (N_4521,N_4348,N_4397);
nand U4522 (N_4522,N_4307,N_4235);
nor U4523 (N_4523,N_4237,N_4373);
nand U4524 (N_4524,N_4232,N_4282);
nor U4525 (N_4525,N_4292,N_4350);
nand U4526 (N_4526,N_4332,N_4237);
nand U4527 (N_4527,N_4375,N_4291);
nand U4528 (N_4528,N_4215,N_4362);
xor U4529 (N_4529,N_4297,N_4300);
nor U4530 (N_4530,N_4299,N_4260);
or U4531 (N_4531,N_4283,N_4338);
nand U4532 (N_4532,N_4330,N_4329);
and U4533 (N_4533,N_4329,N_4247);
or U4534 (N_4534,N_4226,N_4274);
nand U4535 (N_4535,N_4389,N_4312);
xnor U4536 (N_4536,N_4343,N_4384);
nor U4537 (N_4537,N_4367,N_4328);
or U4538 (N_4538,N_4245,N_4231);
or U4539 (N_4539,N_4234,N_4390);
or U4540 (N_4540,N_4333,N_4218);
xor U4541 (N_4541,N_4281,N_4212);
nor U4542 (N_4542,N_4357,N_4329);
xor U4543 (N_4543,N_4298,N_4220);
xor U4544 (N_4544,N_4297,N_4299);
nand U4545 (N_4545,N_4369,N_4222);
nor U4546 (N_4546,N_4220,N_4384);
or U4547 (N_4547,N_4358,N_4255);
nor U4548 (N_4548,N_4284,N_4258);
or U4549 (N_4549,N_4204,N_4373);
nor U4550 (N_4550,N_4378,N_4360);
nor U4551 (N_4551,N_4327,N_4200);
and U4552 (N_4552,N_4309,N_4359);
nand U4553 (N_4553,N_4314,N_4379);
and U4554 (N_4554,N_4291,N_4383);
and U4555 (N_4555,N_4331,N_4382);
or U4556 (N_4556,N_4282,N_4287);
or U4557 (N_4557,N_4240,N_4361);
nand U4558 (N_4558,N_4269,N_4219);
nand U4559 (N_4559,N_4244,N_4374);
nor U4560 (N_4560,N_4291,N_4218);
nand U4561 (N_4561,N_4355,N_4349);
xor U4562 (N_4562,N_4206,N_4319);
nand U4563 (N_4563,N_4293,N_4204);
xnor U4564 (N_4564,N_4311,N_4319);
nand U4565 (N_4565,N_4348,N_4363);
xnor U4566 (N_4566,N_4214,N_4225);
nand U4567 (N_4567,N_4370,N_4393);
nor U4568 (N_4568,N_4325,N_4372);
nand U4569 (N_4569,N_4335,N_4391);
nor U4570 (N_4570,N_4365,N_4394);
nand U4571 (N_4571,N_4366,N_4312);
and U4572 (N_4572,N_4358,N_4261);
nand U4573 (N_4573,N_4293,N_4395);
nand U4574 (N_4574,N_4377,N_4258);
or U4575 (N_4575,N_4292,N_4365);
and U4576 (N_4576,N_4367,N_4336);
xor U4577 (N_4577,N_4293,N_4209);
xor U4578 (N_4578,N_4212,N_4370);
xor U4579 (N_4579,N_4269,N_4275);
xnor U4580 (N_4580,N_4288,N_4336);
xor U4581 (N_4581,N_4355,N_4250);
nor U4582 (N_4582,N_4361,N_4366);
nand U4583 (N_4583,N_4269,N_4308);
xnor U4584 (N_4584,N_4318,N_4321);
or U4585 (N_4585,N_4363,N_4251);
nand U4586 (N_4586,N_4347,N_4316);
and U4587 (N_4587,N_4254,N_4327);
nor U4588 (N_4588,N_4352,N_4212);
nor U4589 (N_4589,N_4326,N_4256);
and U4590 (N_4590,N_4308,N_4275);
xnor U4591 (N_4591,N_4275,N_4287);
nand U4592 (N_4592,N_4369,N_4316);
xor U4593 (N_4593,N_4234,N_4269);
or U4594 (N_4594,N_4245,N_4302);
and U4595 (N_4595,N_4322,N_4379);
and U4596 (N_4596,N_4237,N_4370);
and U4597 (N_4597,N_4359,N_4380);
xnor U4598 (N_4598,N_4295,N_4246);
or U4599 (N_4599,N_4288,N_4340);
and U4600 (N_4600,N_4518,N_4446);
nand U4601 (N_4601,N_4526,N_4503);
or U4602 (N_4602,N_4595,N_4598);
and U4603 (N_4603,N_4570,N_4542);
or U4604 (N_4604,N_4596,N_4591);
xor U4605 (N_4605,N_4530,N_4495);
nand U4606 (N_4606,N_4492,N_4505);
and U4607 (N_4607,N_4471,N_4525);
and U4608 (N_4608,N_4478,N_4462);
and U4609 (N_4609,N_4594,N_4425);
or U4610 (N_4610,N_4479,N_4476);
nand U4611 (N_4611,N_4507,N_4403);
and U4612 (N_4612,N_4430,N_4539);
nand U4613 (N_4613,N_4447,N_4597);
nor U4614 (N_4614,N_4407,N_4512);
or U4615 (N_4615,N_4535,N_4514);
or U4616 (N_4616,N_4494,N_4435);
nor U4617 (N_4617,N_4441,N_4470);
nor U4618 (N_4618,N_4577,N_4592);
and U4619 (N_4619,N_4451,N_4418);
or U4620 (N_4620,N_4419,N_4454);
and U4621 (N_4621,N_4496,N_4438);
xnor U4622 (N_4622,N_4431,N_4500);
or U4623 (N_4623,N_4448,N_4485);
nand U4624 (N_4624,N_4458,N_4456);
nand U4625 (N_4625,N_4569,N_4566);
or U4626 (N_4626,N_4581,N_4547);
and U4627 (N_4627,N_4587,N_4422);
nor U4628 (N_4628,N_4499,N_4497);
xnor U4629 (N_4629,N_4410,N_4538);
nor U4630 (N_4630,N_4585,N_4416);
xnor U4631 (N_4631,N_4589,N_4506);
nor U4632 (N_4632,N_4540,N_4423);
or U4633 (N_4633,N_4437,N_4558);
xor U4634 (N_4634,N_4408,N_4473);
nor U4635 (N_4635,N_4546,N_4417);
nor U4636 (N_4636,N_4405,N_4459);
or U4637 (N_4637,N_4467,N_4561);
xnor U4638 (N_4638,N_4564,N_4582);
nor U4639 (N_4639,N_4529,N_4532);
nor U4640 (N_4640,N_4412,N_4434);
and U4641 (N_4641,N_4554,N_4468);
xnor U4642 (N_4642,N_4536,N_4552);
nor U4643 (N_4643,N_4583,N_4520);
xor U4644 (N_4644,N_4426,N_4450);
or U4645 (N_4645,N_4534,N_4504);
nor U4646 (N_4646,N_4574,N_4599);
or U4647 (N_4647,N_4519,N_4556);
nand U4648 (N_4648,N_4511,N_4593);
and U4649 (N_4649,N_4449,N_4572);
xor U4650 (N_4650,N_4527,N_4560);
nand U4651 (N_4651,N_4442,N_4464);
nor U4652 (N_4652,N_4444,N_4439);
or U4653 (N_4653,N_4414,N_4409);
or U4654 (N_4654,N_4513,N_4579);
and U4655 (N_4655,N_4477,N_4573);
and U4656 (N_4656,N_4401,N_4490);
xnor U4657 (N_4657,N_4484,N_4411);
nor U4658 (N_4658,N_4548,N_4567);
nand U4659 (N_4659,N_4455,N_4420);
and U4660 (N_4660,N_4432,N_4491);
xnor U4661 (N_4661,N_4565,N_4559);
xor U4662 (N_4662,N_4509,N_4400);
xor U4663 (N_4663,N_4580,N_4588);
nand U4664 (N_4664,N_4537,N_4481);
nor U4665 (N_4665,N_4404,N_4533);
and U4666 (N_4666,N_4555,N_4571);
xor U4667 (N_4667,N_4475,N_4487);
nand U4668 (N_4668,N_4590,N_4493);
nor U4669 (N_4669,N_4550,N_4543);
or U4670 (N_4670,N_4578,N_4469);
or U4671 (N_4671,N_4452,N_4482);
and U4672 (N_4672,N_4413,N_4551);
nor U4673 (N_4673,N_4510,N_4415);
or U4674 (N_4674,N_4428,N_4460);
xnor U4675 (N_4675,N_4429,N_4562);
xor U4676 (N_4676,N_4576,N_4465);
nand U4677 (N_4677,N_4402,N_4501);
or U4678 (N_4678,N_4463,N_4515);
nand U4679 (N_4679,N_4440,N_4457);
or U4680 (N_4680,N_4483,N_4472);
xor U4681 (N_4681,N_4433,N_4524);
xor U4682 (N_4682,N_4563,N_4466);
and U4683 (N_4683,N_4406,N_4474);
xnor U4684 (N_4684,N_4461,N_4445);
or U4685 (N_4685,N_4522,N_4528);
xor U4686 (N_4686,N_4427,N_4523);
nor U4687 (N_4687,N_4586,N_4531);
and U4688 (N_4688,N_4488,N_4553);
and U4689 (N_4689,N_4424,N_4421);
xnor U4690 (N_4690,N_4541,N_4545);
nand U4691 (N_4691,N_4549,N_4443);
xor U4692 (N_4692,N_4557,N_4489);
xnor U4693 (N_4693,N_4508,N_4486);
xnor U4694 (N_4694,N_4521,N_4568);
nor U4695 (N_4695,N_4498,N_4516);
xor U4696 (N_4696,N_4502,N_4453);
or U4697 (N_4697,N_4517,N_4480);
xor U4698 (N_4698,N_4436,N_4584);
nor U4699 (N_4699,N_4544,N_4575);
nand U4700 (N_4700,N_4439,N_4462);
or U4701 (N_4701,N_4447,N_4405);
nand U4702 (N_4702,N_4539,N_4535);
and U4703 (N_4703,N_4582,N_4569);
nand U4704 (N_4704,N_4417,N_4572);
nand U4705 (N_4705,N_4544,N_4588);
nor U4706 (N_4706,N_4499,N_4568);
nor U4707 (N_4707,N_4429,N_4582);
xnor U4708 (N_4708,N_4595,N_4524);
nor U4709 (N_4709,N_4425,N_4595);
or U4710 (N_4710,N_4548,N_4511);
xnor U4711 (N_4711,N_4420,N_4544);
nand U4712 (N_4712,N_4508,N_4580);
nor U4713 (N_4713,N_4527,N_4578);
or U4714 (N_4714,N_4469,N_4580);
xor U4715 (N_4715,N_4495,N_4499);
and U4716 (N_4716,N_4415,N_4470);
xnor U4717 (N_4717,N_4512,N_4465);
xnor U4718 (N_4718,N_4555,N_4446);
or U4719 (N_4719,N_4599,N_4417);
or U4720 (N_4720,N_4426,N_4579);
nand U4721 (N_4721,N_4568,N_4567);
xor U4722 (N_4722,N_4478,N_4535);
or U4723 (N_4723,N_4520,N_4558);
and U4724 (N_4724,N_4447,N_4440);
nand U4725 (N_4725,N_4489,N_4592);
nor U4726 (N_4726,N_4458,N_4423);
and U4727 (N_4727,N_4494,N_4545);
or U4728 (N_4728,N_4423,N_4538);
xor U4729 (N_4729,N_4514,N_4463);
xor U4730 (N_4730,N_4432,N_4435);
and U4731 (N_4731,N_4474,N_4582);
and U4732 (N_4732,N_4442,N_4466);
or U4733 (N_4733,N_4587,N_4538);
or U4734 (N_4734,N_4422,N_4487);
or U4735 (N_4735,N_4456,N_4508);
xnor U4736 (N_4736,N_4556,N_4522);
xnor U4737 (N_4737,N_4596,N_4580);
and U4738 (N_4738,N_4434,N_4415);
or U4739 (N_4739,N_4444,N_4540);
and U4740 (N_4740,N_4530,N_4434);
nand U4741 (N_4741,N_4552,N_4527);
and U4742 (N_4742,N_4491,N_4583);
and U4743 (N_4743,N_4545,N_4538);
nand U4744 (N_4744,N_4416,N_4400);
xor U4745 (N_4745,N_4561,N_4576);
nand U4746 (N_4746,N_4500,N_4429);
nand U4747 (N_4747,N_4595,N_4552);
nand U4748 (N_4748,N_4473,N_4495);
nand U4749 (N_4749,N_4521,N_4451);
and U4750 (N_4750,N_4543,N_4460);
nand U4751 (N_4751,N_4459,N_4524);
nand U4752 (N_4752,N_4433,N_4441);
and U4753 (N_4753,N_4486,N_4480);
nor U4754 (N_4754,N_4539,N_4449);
and U4755 (N_4755,N_4527,N_4522);
or U4756 (N_4756,N_4514,N_4533);
xnor U4757 (N_4757,N_4580,N_4552);
or U4758 (N_4758,N_4560,N_4401);
or U4759 (N_4759,N_4593,N_4514);
or U4760 (N_4760,N_4423,N_4454);
nand U4761 (N_4761,N_4536,N_4534);
nor U4762 (N_4762,N_4469,N_4582);
xor U4763 (N_4763,N_4406,N_4482);
xnor U4764 (N_4764,N_4554,N_4493);
and U4765 (N_4765,N_4553,N_4566);
or U4766 (N_4766,N_4514,N_4404);
nand U4767 (N_4767,N_4454,N_4549);
nor U4768 (N_4768,N_4560,N_4593);
nor U4769 (N_4769,N_4558,N_4574);
xnor U4770 (N_4770,N_4485,N_4451);
nand U4771 (N_4771,N_4589,N_4530);
xnor U4772 (N_4772,N_4592,N_4546);
nor U4773 (N_4773,N_4512,N_4472);
xor U4774 (N_4774,N_4570,N_4410);
nor U4775 (N_4775,N_4549,N_4464);
and U4776 (N_4776,N_4498,N_4576);
nand U4777 (N_4777,N_4576,N_4573);
nand U4778 (N_4778,N_4590,N_4505);
and U4779 (N_4779,N_4470,N_4536);
nor U4780 (N_4780,N_4538,N_4567);
nand U4781 (N_4781,N_4548,N_4427);
or U4782 (N_4782,N_4552,N_4576);
nor U4783 (N_4783,N_4470,N_4565);
nor U4784 (N_4784,N_4500,N_4562);
or U4785 (N_4785,N_4461,N_4562);
xor U4786 (N_4786,N_4484,N_4483);
nor U4787 (N_4787,N_4525,N_4548);
xnor U4788 (N_4788,N_4413,N_4542);
and U4789 (N_4789,N_4577,N_4447);
or U4790 (N_4790,N_4596,N_4459);
or U4791 (N_4791,N_4455,N_4425);
and U4792 (N_4792,N_4450,N_4435);
and U4793 (N_4793,N_4456,N_4463);
nor U4794 (N_4794,N_4456,N_4400);
nand U4795 (N_4795,N_4448,N_4535);
xor U4796 (N_4796,N_4485,N_4426);
or U4797 (N_4797,N_4493,N_4524);
and U4798 (N_4798,N_4551,N_4484);
xor U4799 (N_4799,N_4564,N_4563);
or U4800 (N_4800,N_4626,N_4651);
xnor U4801 (N_4801,N_4666,N_4757);
nor U4802 (N_4802,N_4774,N_4676);
nand U4803 (N_4803,N_4617,N_4613);
or U4804 (N_4804,N_4646,N_4788);
and U4805 (N_4805,N_4687,N_4760);
xor U4806 (N_4806,N_4686,N_4604);
xnor U4807 (N_4807,N_4717,N_4710);
nor U4808 (N_4808,N_4649,N_4732);
and U4809 (N_4809,N_4729,N_4795);
nor U4810 (N_4810,N_4691,N_4727);
xor U4811 (N_4811,N_4678,N_4681);
and U4812 (N_4812,N_4643,N_4719);
nand U4813 (N_4813,N_4690,N_4754);
or U4814 (N_4814,N_4654,N_4749);
nand U4815 (N_4815,N_4724,N_4636);
nand U4816 (N_4816,N_4665,N_4793);
and U4817 (N_4817,N_4694,N_4752);
nand U4818 (N_4818,N_4737,N_4645);
xnor U4819 (N_4819,N_4782,N_4722);
nand U4820 (N_4820,N_4794,N_4735);
nand U4821 (N_4821,N_4620,N_4769);
or U4822 (N_4822,N_4607,N_4638);
or U4823 (N_4823,N_4775,N_4743);
or U4824 (N_4824,N_4639,N_4618);
and U4825 (N_4825,N_4712,N_4787);
and U4826 (N_4826,N_4693,N_4670);
or U4827 (N_4827,N_4742,N_4781);
or U4828 (N_4828,N_4606,N_4672);
nand U4829 (N_4829,N_4635,N_4704);
xor U4830 (N_4830,N_4658,N_4718);
and U4831 (N_4831,N_4758,N_4616);
nand U4832 (N_4832,N_4792,N_4627);
nand U4833 (N_4833,N_4675,N_4648);
and U4834 (N_4834,N_4716,N_4730);
xor U4835 (N_4835,N_4789,N_4707);
and U4836 (N_4836,N_4685,N_4667);
and U4837 (N_4837,N_4623,N_4725);
or U4838 (N_4838,N_4631,N_4714);
xor U4839 (N_4839,N_4709,N_4771);
xor U4840 (N_4840,N_4711,N_4747);
xor U4841 (N_4841,N_4736,N_4673);
or U4842 (N_4842,N_4728,N_4761);
nand U4843 (N_4843,N_4799,N_4652);
xnor U4844 (N_4844,N_4679,N_4700);
nand U4845 (N_4845,N_4664,N_4759);
xnor U4846 (N_4846,N_4680,N_4695);
xnor U4847 (N_4847,N_4756,N_4653);
xor U4848 (N_4848,N_4772,N_4706);
xnor U4849 (N_4849,N_4753,N_4777);
nor U4850 (N_4850,N_4798,N_4605);
nand U4851 (N_4851,N_4750,N_4696);
xnor U4852 (N_4852,N_4768,N_4647);
nor U4853 (N_4853,N_4739,N_4703);
nand U4854 (N_4854,N_4790,N_4660);
nand U4855 (N_4855,N_4601,N_4628);
nand U4856 (N_4856,N_4726,N_4655);
or U4857 (N_4857,N_4796,N_4765);
and U4858 (N_4858,N_4698,N_4755);
xnor U4859 (N_4859,N_4662,N_4766);
and U4860 (N_4860,N_4671,N_4634);
and U4861 (N_4861,N_4740,N_4744);
xnor U4862 (N_4862,N_4784,N_4723);
xnor U4863 (N_4863,N_4783,N_4708);
or U4864 (N_4864,N_4734,N_4689);
or U4865 (N_4865,N_4612,N_4640);
or U4866 (N_4866,N_4731,N_4763);
nor U4867 (N_4867,N_4773,N_4659);
and U4868 (N_4868,N_4770,N_4746);
or U4869 (N_4869,N_4713,N_4776);
xor U4870 (N_4870,N_4797,N_4786);
xor U4871 (N_4871,N_4745,N_4622);
and U4872 (N_4872,N_4669,N_4668);
or U4873 (N_4873,N_4656,N_4600);
xor U4874 (N_4874,N_4619,N_4684);
or U4875 (N_4875,N_4630,N_4741);
nor U4876 (N_4876,N_4692,N_4641);
or U4877 (N_4877,N_4702,N_4762);
nor U4878 (N_4878,N_4682,N_4611);
or U4879 (N_4879,N_4699,N_4779);
xnor U4880 (N_4880,N_4602,N_4608);
nor U4881 (N_4881,N_4632,N_4624);
or U4882 (N_4882,N_4701,N_4642);
nand U4883 (N_4883,N_4764,N_4720);
or U4884 (N_4884,N_4683,N_4688);
nand U4885 (N_4885,N_4633,N_4610);
nor U4886 (N_4886,N_4637,N_4791);
and U4887 (N_4887,N_4738,N_4674);
nand U4888 (N_4888,N_4621,N_4625);
xnor U4889 (N_4889,N_4650,N_4629);
nand U4890 (N_4890,N_4644,N_4778);
nor U4891 (N_4891,N_4715,N_4748);
nor U4892 (N_4892,N_4603,N_4697);
nand U4893 (N_4893,N_4785,N_4614);
and U4894 (N_4894,N_4657,N_4677);
nor U4895 (N_4895,N_4705,N_4721);
xnor U4896 (N_4896,N_4663,N_4615);
nand U4897 (N_4897,N_4733,N_4661);
nand U4898 (N_4898,N_4609,N_4767);
xnor U4899 (N_4899,N_4780,N_4751);
and U4900 (N_4900,N_4721,N_4636);
or U4901 (N_4901,N_4695,N_4609);
and U4902 (N_4902,N_4706,N_4699);
xor U4903 (N_4903,N_4617,N_4639);
nor U4904 (N_4904,N_4744,N_4787);
nand U4905 (N_4905,N_4729,N_4683);
nand U4906 (N_4906,N_4734,N_4666);
or U4907 (N_4907,N_4703,N_4610);
and U4908 (N_4908,N_4671,N_4713);
nor U4909 (N_4909,N_4655,N_4737);
nor U4910 (N_4910,N_4784,N_4638);
and U4911 (N_4911,N_4645,N_4700);
nor U4912 (N_4912,N_4765,N_4617);
and U4913 (N_4913,N_4679,N_4693);
nor U4914 (N_4914,N_4631,N_4780);
xnor U4915 (N_4915,N_4696,N_4740);
nor U4916 (N_4916,N_4739,N_4775);
nand U4917 (N_4917,N_4715,N_4743);
nand U4918 (N_4918,N_4766,N_4790);
and U4919 (N_4919,N_4765,N_4606);
and U4920 (N_4920,N_4743,N_4799);
nand U4921 (N_4921,N_4658,N_4685);
or U4922 (N_4922,N_4736,N_4764);
and U4923 (N_4923,N_4600,N_4601);
nor U4924 (N_4924,N_4682,N_4718);
and U4925 (N_4925,N_4684,N_4630);
and U4926 (N_4926,N_4684,N_4681);
nor U4927 (N_4927,N_4715,N_4710);
or U4928 (N_4928,N_4729,N_4601);
and U4929 (N_4929,N_4720,N_4688);
and U4930 (N_4930,N_4647,N_4705);
or U4931 (N_4931,N_4652,N_4788);
or U4932 (N_4932,N_4715,N_4620);
or U4933 (N_4933,N_4683,N_4768);
nand U4934 (N_4934,N_4745,N_4659);
and U4935 (N_4935,N_4714,N_4635);
and U4936 (N_4936,N_4706,N_4610);
nor U4937 (N_4937,N_4634,N_4731);
or U4938 (N_4938,N_4685,N_4644);
nor U4939 (N_4939,N_4615,N_4657);
nor U4940 (N_4940,N_4705,N_4642);
nor U4941 (N_4941,N_4777,N_4649);
xor U4942 (N_4942,N_4629,N_4739);
nand U4943 (N_4943,N_4656,N_4679);
or U4944 (N_4944,N_4759,N_4721);
xnor U4945 (N_4945,N_4646,N_4631);
or U4946 (N_4946,N_4666,N_4615);
or U4947 (N_4947,N_4674,N_4748);
or U4948 (N_4948,N_4790,N_4683);
xor U4949 (N_4949,N_4651,N_4750);
xor U4950 (N_4950,N_4704,N_4776);
nand U4951 (N_4951,N_4754,N_4614);
nand U4952 (N_4952,N_4750,N_4719);
xor U4953 (N_4953,N_4781,N_4614);
nand U4954 (N_4954,N_4746,N_4655);
nor U4955 (N_4955,N_4635,N_4766);
nand U4956 (N_4956,N_4630,N_4705);
and U4957 (N_4957,N_4771,N_4671);
xnor U4958 (N_4958,N_4773,N_4660);
or U4959 (N_4959,N_4741,N_4687);
nor U4960 (N_4960,N_4718,N_4661);
nand U4961 (N_4961,N_4742,N_4740);
nor U4962 (N_4962,N_4754,N_4677);
and U4963 (N_4963,N_4640,N_4695);
nor U4964 (N_4964,N_4684,N_4712);
and U4965 (N_4965,N_4785,N_4704);
or U4966 (N_4966,N_4637,N_4619);
xnor U4967 (N_4967,N_4766,N_4665);
xor U4968 (N_4968,N_4672,N_4662);
nand U4969 (N_4969,N_4647,N_4657);
nand U4970 (N_4970,N_4629,N_4740);
nor U4971 (N_4971,N_4767,N_4638);
nor U4972 (N_4972,N_4685,N_4689);
and U4973 (N_4973,N_4650,N_4685);
and U4974 (N_4974,N_4646,N_4660);
nor U4975 (N_4975,N_4760,N_4656);
nand U4976 (N_4976,N_4683,N_4677);
nor U4977 (N_4977,N_4646,N_4685);
xor U4978 (N_4978,N_4768,N_4697);
or U4979 (N_4979,N_4631,N_4789);
xor U4980 (N_4980,N_4719,N_4745);
nand U4981 (N_4981,N_4785,N_4798);
nand U4982 (N_4982,N_4638,N_4775);
or U4983 (N_4983,N_4656,N_4635);
and U4984 (N_4984,N_4736,N_4781);
nand U4985 (N_4985,N_4762,N_4780);
nor U4986 (N_4986,N_4686,N_4682);
nor U4987 (N_4987,N_4748,N_4708);
nand U4988 (N_4988,N_4790,N_4788);
or U4989 (N_4989,N_4704,N_4629);
nor U4990 (N_4990,N_4707,N_4788);
xor U4991 (N_4991,N_4659,N_4724);
or U4992 (N_4992,N_4789,N_4649);
or U4993 (N_4993,N_4711,N_4725);
nand U4994 (N_4994,N_4799,N_4786);
and U4995 (N_4995,N_4729,N_4784);
xnor U4996 (N_4996,N_4657,N_4603);
nand U4997 (N_4997,N_4611,N_4699);
nor U4998 (N_4998,N_4744,N_4619);
xor U4999 (N_4999,N_4648,N_4628);
and UO_0 (O_0,N_4827,N_4980);
nor UO_1 (O_1,N_4888,N_4837);
nand UO_2 (O_2,N_4857,N_4983);
nand UO_3 (O_3,N_4999,N_4886);
and UO_4 (O_4,N_4903,N_4877);
or UO_5 (O_5,N_4961,N_4951);
xor UO_6 (O_6,N_4977,N_4802);
and UO_7 (O_7,N_4950,N_4893);
xor UO_8 (O_8,N_4883,N_4973);
and UO_9 (O_9,N_4940,N_4800);
and UO_10 (O_10,N_4807,N_4863);
xnor UO_11 (O_11,N_4957,N_4833);
nand UO_12 (O_12,N_4892,N_4904);
and UO_13 (O_13,N_4933,N_4869);
nand UO_14 (O_14,N_4941,N_4835);
and UO_15 (O_15,N_4874,N_4810);
or UO_16 (O_16,N_4806,N_4954);
or UO_17 (O_17,N_4936,N_4910);
nor UO_18 (O_18,N_4914,N_4852);
xnor UO_19 (O_19,N_4953,N_4830);
and UO_20 (O_20,N_4998,N_4817);
xnor UO_21 (O_21,N_4839,N_4938);
and UO_22 (O_22,N_4952,N_4944);
nand UO_23 (O_23,N_4885,N_4978);
or UO_24 (O_24,N_4974,N_4841);
nand UO_25 (O_25,N_4905,N_4862);
or UO_26 (O_26,N_4822,N_4889);
xor UO_27 (O_27,N_4934,N_4887);
nand UO_28 (O_28,N_4947,N_4923);
nand UO_29 (O_29,N_4894,N_4884);
xnor UO_30 (O_30,N_4860,N_4897);
nand UO_31 (O_31,N_4815,N_4819);
and UO_32 (O_32,N_4891,N_4908);
and UO_33 (O_33,N_4962,N_4967);
nand UO_34 (O_34,N_4823,N_4868);
and UO_35 (O_35,N_4937,N_4928);
nand UO_36 (O_36,N_4917,N_4955);
nand UO_37 (O_37,N_4930,N_4964);
or UO_38 (O_38,N_4963,N_4945);
xor UO_39 (O_39,N_4927,N_4882);
or UO_40 (O_40,N_4804,N_4926);
and UO_41 (O_41,N_4913,N_4820);
or UO_42 (O_42,N_4932,N_4909);
or UO_43 (O_43,N_4831,N_4821);
and UO_44 (O_44,N_4811,N_4829);
xor UO_45 (O_45,N_4872,N_4971);
xnor UO_46 (O_46,N_4994,N_4968);
nand UO_47 (O_47,N_4946,N_4834);
or UO_48 (O_48,N_4881,N_4920);
and UO_49 (O_49,N_4854,N_4912);
nand UO_50 (O_50,N_4879,N_4981);
xor UO_51 (O_51,N_4838,N_4918);
xor UO_52 (O_52,N_4921,N_4939);
nor UO_53 (O_53,N_4986,N_4808);
nor UO_54 (O_54,N_4942,N_4846);
xor UO_55 (O_55,N_4958,N_4989);
nor UO_56 (O_56,N_4825,N_4890);
nand UO_57 (O_57,N_4925,N_4842);
xnor UO_58 (O_58,N_4997,N_4924);
nor UO_59 (O_59,N_4898,N_4972);
xnor UO_60 (O_60,N_4818,N_4844);
and UO_61 (O_61,N_4959,N_4824);
or UO_62 (O_62,N_4993,N_4960);
and UO_63 (O_63,N_4840,N_4803);
nor UO_64 (O_64,N_4876,N_4979);
and UO_65 (O_65,N_4864,N_4956);
or UO_66 (O_66,N_4809,N_4965);
and UO_67 (O_67,N_4856,N_4985);
nand UO_68 (O_68,N_4943,N_4853);
xnor UO_69 (O_69,N_4875,N_4901);
xnor UO_70 (O_70,N_4988,N_4896);
nand UO_71 (O_71,N_4919,N_4902);
or UO_72 (O_72,N_4915,N_4849);
xor UO_73 (O_73,N_4870,N_4812);
or UO_74 (O_74,N_4848,N_4899);
or UO_75 (O_75,N_4975,N_4966);
or UO_76 (O_76,N_4929,N_4949);
xor UO_77 (O_77,N_4995,N_4832);
xor UO_78 (O_78,N_4935,N_4805);
and UO_79 (O_79,N_4992,N_4865);
nand UO_80 (O_80,N_4991,N_4866);
and UO_81 (O_81,N_4801,N_4814);
xnor UO_82 (O_82,N_4878,N_4987);
nand UO_83 (O_83,N_4907,N_4931);
xor UO_84 (O_84,N_4916,N_4996);
or UO_85 (O_85,N_4922,N_4948);
nand UO_86 (O_86,N_4826,N_4906);
nand UO_87 (O_87,N_4984,N_4873);
nand UO_88 (O_88,N_4990,N_4847);
nand UO_89 (O_89,N_4976,N_4867);
and UO_90 (O_90,N_4836,N_4843);
nand UO_91 (O_91,N_4861,N_4880);
and UO_92 (O_92,N_4970,N_4828);
xor UO_93 (O_93,N_4850,N_4813);
or UO_94 (O_94,N_4859,N_4900);
nor UO_95 (O_95,N_4845,N_4858);
and UO_96 (O_96,N_4871,N_4855);
or UO_97 (O_97,N_4969,N_4911);
and UO_98 (O_98,N_4816,N_4982);
xor UO_99 (O_99,N_4895,N_4851);
nor UO_100 (O_100,N_4938,N_4972);
and UO_101 (O_101,N_4924,N_4971);
nor UO_102 (O_102,N_4838,N_4955);
nor UO_103 (O_103,N_4973,N_4813);
nor UO_104 (O_104,N_4844,N_4992);
xor UO_105 (O_105,N_4895,N_4876);
or UO_106 (O_106,N_4953,N_4866);
and UO_107 (O_107,N_4963,N_4956);
or UO_108 (O_108,N_4857,N_4969);
nand UO_109 (O_109,N_4879,N_4896);
nand UO_110 (O_110,N_4823,N_4944);
nand UO_111 (O_111,N_4910,N_4985);
or UO_112 (O_112,N_4854,N_4863);
xor UO_113 (O_113,N_4963,N_4893);
and UO_114 (O_114,N_4907,N_4812);
xor UO_115 (O_115,N_4827,N_4941);
xor UO_116 (O_116,N_4897,N_4927);
nor UO_117 (O_117,N_4887,N_4804);
nand UO_118 (O_118,N_4807,N_4834);
nand UO_119 (O_119,N_4879,N_4812);
or UO_120 (O_120,N_4847,N_4857);
nor UO_121 (O_121,N_4913,N_4814);
or UO_122 (O_122,N_4894,N_4901);
nand UO_123 (O_123,N_4999,N_4994);
nand UO_124 (O_124,N_4910,N_4876);
and UO_125 (O_125,N_4998,N_4951);
xor UO_126 (O_126,N_4935,N_4874);
or UO_127 (O_127,N_4920,N_4949);
xor UO_128 (O_128,N_4802,N_4903);
xnor UO_129 (O_129,N_4914,N_4829);
nor UO_130 (O_130,N_4969,N_4946);
xnor UO_131 (O_131,N_4806,N_4973);
or UO_132 (O_132,N_4940,N_4943);
nand UO_133 (O_133,N_4890,N_4989);
nand UO_134 (O_134,N_4835,N_4884);
nand UO_135 (O_135,N_4802,N_4899);
or UO_136 (O_136,N_4967,N_4845);
xor UO_137 (O_137,N_4806,N_4941);
nand UO_138 (O_138,N_4938,N_4964);
or UO_139 (O_139,N_4808,N_4946);
or UO_140 (O_140,N_4904,N_4894);
nand UO_141 (O_141,N_4815,N_4989);
xnor UO_142 (O_142,N_4923,N_4969);
xor UO_143 (O_143,N_4973,N_4833);
xor UO_144 (O_144,N_4817,N_4811);
nand UO_145 (O_145,N_4825,N_4943);
and UO_146 (O_146,N_4822,N_4827);
nor UO_147 (O_147,N_4921,N_4884);
nand UO_148 (O_148,N_4832,N_4870);
or UO_149 (O_149,N_4878,N_4953);
or UO_150 (O_150,N_4929,N_4914);
nor UO_151 (O_151,N_4830,N_4984);
nand UO_152 (O_152,N_4845,N_4884);
nand UO_153 (O_153,N_4862,N_4849);
nand UO_154 (O_154,N_4918,N_4858);
and UO_155 (O_155,N_4813,N_4863);
nand UO_156 (O_156,N_4832,N_4852);
or UO_157 (O_157,N_4802,N_4817);
nor UO_158 (O_158,N_4846,N_4943);
nor UO_159 (O_159,N_4911,N_4866);
and UO_160 (O_160,N_4931,N_4942);
and UO_161 (O_161,N_4827,N_4947);
or UO_162 (O_162,N_4974,N_4881);
nor UO_163 (O_163,N_4884,N_4841);
nor UO_164 (O_164,N_4959,N_4905);
and UO_165 (O_165,N_4846,N_4849);
nand UO_166 (O_166,N_4994,N_4911);
or UO_167 (O_167,N_4909,N_4995);
nor UO_168 (O_168,N_4923,N_4997);
nand UO_169 (O_169,N_4842,N_4803);
or UO_170 (O_170,N_4850,N_4824);
nor UO_171 (O_171,N_4950,N_4843);
nor UO_172 (O_172,N_4921,N_4898);
or UO_173 (O_173,N_4813,N_4890);
or UO_174 (O_174,N_4886,N_4862);
or UO_175 (O_175,N_4894,N_4983);
xnor UO_176 (O_176,N_4975,N_4839);
nor UO_177 (O_177,N_4879,N_4986);
xnor UO_178 (O_178,N_4974,N_4925);
nor UO_179 (O_179,N_4955,N_4834);
or UO_180 (O_180,N_4920,N_4929);
xnor UO_181 (O_181,N_4951,N_4905);
nand UO_182 (O_182,N_4819,N_4947);
nor UO_183 (O_183,N_4828,N_4920);
nor UO_184 (O_184,N_4956,N_4903);
and UO_185 (O_185,N_4861,N_4955);
xnor UO_186 (O_186,N_4986,N_4927);
xor UO_187 (O_187,N_4807,N_4821);
or UO_188 (O_188,N_4985,N_4803);
xnor UO_189 (O_189,N_4961,N_4812);
and UO_190 (O_190,N_4973,N_4945);
and UO_191 (O_191,N_4808,N_4824);
or UO_192 (O_192,N_4863,N_4867);
or UO_193 (O_193,N_4940,N_4832);
and UO_194 (O_194,N_4824,N_4868);
nor UO_195 (O_195,N_4960,N_4866);
and UO_196 (O_196,N_4834,N_4803);
and UO_197 (O_197,N_4861,N_4892);
nor UO_198 (O_198,N_4945,N_4915);
nand UO_199 (O_199,N_4993,N_4979);
or UO_200 (O_200,N_4889,N_4840);
or UO_201 (O_201,N_4951,N_4931);
xor UO_202 (O_202,N_4817,N_4840);
nor UO_203 (O_203,N_4989,N_4922);
or UO_204 (O_204,N_4958,N_4854);
and UO_205 (O_205,N_4847,N_4886);
or UO_206 (O_206,N_4916,N_4920);
xnor UO_207 (O_207,N_4934,N_4800);
xor UO_208 (O_208,N_4811,N_4918);
nand UO_209 (O_209,N_4850,N_4832);
and UO_210 (O_210,N_4873,N_4904);
xor UO_211 (O_211,N_4953,N_4918);
and UO_212 (O_212,N_4808,N_4945);
and UO_213 (O_213,N_4838,N_4875);
xor UO_214 (O_214,N_4836,N_4908);
or UO_215 (O_215,N_4888,N_4947);
xnor UO_216 (O_216,N_4966,N_4896);
nand UO_217 (O_217,N_4938,N_4824);
or UO_218 (O_218,N_4856,N_4954);
and UO_219 (O_219,N_4872,N_4961);
nand UO_220 (O_220,N_4924,N_4825);
and UO_221 (O_221,N_4983,N_4811);
nor UO_222 (O_222,N_4909,N_4805);
xor UO_223 (O_223,N_4831,N_4946);
and UO_224 (O_224,N_4993,N_4890);
or UO_225 (O_225,N_4831,N_4912);
xor UO_226 (O_226,N_4867,N_4801);
or UO_227 (O_227,N_4968,N_4816);
or UO_228 (O_228,N_4808,N_4982);
xor UO_229 (O_229,N_4806,N_4917);
and UO_230 (O_230,N_4913,N_4968);
nor UO_231 (O_231,N_4923,N_4820);
and UO_232 (O_232,N_4824,N_4915);
xnor UO_233 (O_233,N_4848,N_4963);
and UO_234 (O_234,N_4857,N_4827);
or UO_235 (O_235,N_4815,N_4895);
and UO_236 (O_236,N_4896,N_4921);
and UO_237 (O_237,N_4819,N_4948);
nor UO_238 (O_238,N_4901,N_4827);
nor UO_239 (O_239,N_4869,N_4968);
nor UO_240 (O_240,N_4963,N_4964);
or UO_241 (O_241,N_4842,N_4997);
xor UO_242 (O_242,N_4934,N_4998);
or UO_243 (O_243,N_4990,N_4991);
nor UO_244 (O_244,N_4816,N_4997);
or UO_245 (O_245,N_4867,N_4902);
nor UO_246 (O_246,N_4859,N_4960);
or UO_247 (O_247,N_4954,N_4961);
nor UO_248 (O_248,N_4996,N_4888);
and UO_249 (O_249,N_4990,N_4870);
xnor UO_250 (O_250,N_4940,N_4855);
and UO_251 (O_251,N_4949,N_4851);
or UO_252 (O_252,N_4864,N_4871);
nor UO_253 (O_253,N_4878,N_4875);
nand UO_254 (O_254,N_4811,N_4854);
and UO_255 (O_255,N_4856,N_4871);
nand UO_256 (O_256,N_4809,N_4909);
nor UO_257 (O_257,N_4970,N_4801);
nor UO_258 (O_258,N_4917,N_4949);
nor UO_259 (O_259,N_4918,N_4994);
nand UO_260 (O_260,N_4956,N_4883);
and UO_261 (O_261,N_4995,N_4828);
nand UO_262 (O_262,N_4840,N_4849);
or UO_263 (O_263,N_4983,N_4887);
or UO_264 (O_264,N_4854,N_4993);
or UO_265 (O_265,N_4804,N_4840);
or UO_266 (O_266,N_4935,N_4856);
xor UO_267 (O_267,N_4838,N_4872);
nor UO_268 (O_268,N_4941,N_4805);
or UO_269 (O_269,N_4878,N_4881);
nor UO_270 (O_270,N_4952,N_4945);
and UO_271 (O_271,N_4929,N_4885);
and UO_272 (O_272,N_4935,N_4984);
or UO_273 (O_273,N_4816,N_4908);
nand UO_274 (O_274,N_4946,N_4838);
xnor UO_275 (O_275,N_4905,N_4808);
xnor UO_276 (O_276,N_4902,N_4863);
or UO_277 (O_277,N_4976,N_4950);
nor UO_278 (O_278,N_4905,N_4848);
and UO_279 (O_279,N_4867,N_4982);
nor UO_280 (O_280,N_4922,N_4923);
and UO_281 (O_281,N_4929,N_4911);
nand UO_282 (O_282,N_4913,N_4815);
and UO_283 (O_283,N_4993,N_4909);
nor UO_284 (O_284,N_4830,N_4856);
nor UO_285 (O_285,N_4879,N_4878);
and UO_286 (O_286,N_4882,N_4819);
nand UO_287 (O_287,N_4902,N_4943);
and UO_288 (O_288,N_4906,N_4996);
or UO_289 (O_289,N_4829,N_4817);
nand UO_290 (O_290,N_4827,N_4992);
nand UO_291 (O_291,N_4826,N_4834);
nand UO_292 (O_292,N_4876,N_4854);
nand UO_293 (O_293,N_4975,N_4875);
xor UO_294 (O_294,N_4999,N_4945);
nor UO_295 (O_295,N_4969,N_4950);
or UO_296 (O_296,N_4914,N_4990);
nor UO_297 (O_297,N_4938,N_4891);
nor UO_298 (O_298,N_4910,N_4930);
or UO_299 (O_299,N_4967,N_4985);
or UO_300 (O_300,N_4951,N_4872);
nor UO_301 (O_301,N_4936,N_4871);
xor UO_302 (O_302,N_4976,N_4943);
nor UO_303 (O_303,N_4963,N_4993);
xor UO_304 (O_304,N_4846,N_4828);
xnor UO_305 (O_305,N_4978,N_4872);
nor UO_306 (O_306,N_4921,N_4809);
nand UO_307 (O_307,N_4801,N_4994);
and UO_308 (O_308,N_4994,N_4946);
or UO_309 (O_309,N_4818,N_4839);
nand UO_310 (O_310,N_4802,N_4934);
or UO_311 (O_311,N_4892,N_4883);
or UO_312 (O_312,N_4807,N_4992);
and UO_313 (O_313,N_4918,N_4934);
and UO_314 (O_314,N_4920,N_4811);
nor UO_315 (O_315,N_4847,N_4914);
or UO_316 (O_316,N_4873,N_4881);
and UO_317 (O_317,N_4845,N_4848);
xor UO_318 (O_318,N_4880,N_4957);
and UO_319 (O_319,N_4988,N_4807);
nor UO_320 (O_320,N_4849,N_4925);
xor UO_321 (O_321,N_4800,N_4858);
nand UO_322 (O_322,N_4838,N_4904);
xnor UO_323 (O_323,N_4926,N_4810);
and UO_324 (O_324,N_4968,N_4862);
nand UO_325 (O_325,N_4888,N_4906);
nor UO_326 (O_326,N_4924,N_4886);
and UO_327 (O_327,N_4873,N_4890);
nand UO_328 (O_328,N_4805,N_4931);
nor UO_329 (O_329,N_4985,N_4954);
xnor UO_330 (O_330,N_4936,N_4903);
and UO_331 (O_331,N_4957,N_4976);
nor UO_332 (O_332,N_4834,N_4940);
nor UO_333 (O_333,N_4872,N_4989);
or UO_334 (O_334,N_4867,N_4893);
and UO_335 (O_335,N_4975,N_4870);
or UO_336 (O_336,N_4875,N_4919);
nand UO_337 (O_337,N_4849,N_4850);
nor UO_338 (O_338,N_4987,N_4937);
and UO_339 (O_339,N_4851,N_4947);
nor UO_340 (O_340,N_4961,N_4887);
or UO_341 (O_341,N_4914,N_4885);
or UO_342 (O_342,N_4901,N_4848);
and UO_343 (O_343,N_4978,N_4969);
nand UO_344 (O_344,N_4830,N_4902);
xor UO_345 (O_345,N_4804,N_4965);
nor UO_346 (O_346,N_4802,N_4902);
or UO_347 (O_347,N_4918,N_4917);
nand UO_348 (O_348,N_4978,N_4800);
nor UO_349 (O_349,N_4814,N_4832);
and UO_350 (O_350,N_4909,N_4858);
nand UO_351 (O_351,N_4971,N_4822);
and UO_352 (O_352,N_4849,N_4897);
xnor UO_353 (O_353,N_4985,N_4971);
xor UO_354 (O_354,N_4989,N_4939);
or UO_355 (O_355,N_4953,N_4962);
nor UO_356 (O_356,N_4830,N_4929);
and UO_357 (O_357,N_4931,N_4976);
nor UO_358 (O_358,N_4891,N_4996);
nand UO_359 (O_359,N_4894,N_4838);
and UO_360 (O_360,N_4928,N_4816);
and UO_361 (O_361,N_4884,N_4977);
nor UO_362 (O_362,N_4937,N_4865);
nor UO_363 (O_363,N_4996,N_4847);
and UO_364 (O_364,N_4885,N_4834);
and UO_365 (O_365,N_4959,N_4814);
xor UO_366 (O_366,N_4822,N_4819);
nand UO_367 (O_367,N_4977,N_4953);
nand UO_368 (O_368,N_4981,N_4825);
nor UO_369 (O_369,N_4825,N_4845);
and UO_370 (O_370,N_4889,N_4811);
or UO_371 (O_371,N_4964,N_4974);
and UO_372 (O_372,N_4972,N_4868);
or UO_373 (O_373,N_4962,N_4985);
nand UO_374 (O_374,N_4829,N_4836);
or UO_375 (O_375,N_4967,N_4850);
xor UO_376 (O_376,N_4953,N_4932);
xnor UO_377 (O_377,N_4885,N_4980);
nor UO_378 (O_378,N_4944,N_4956);
or UO_379 (O_379,N_4923,N_4952);
or UO_380 (O_380,N_4927,N_4922);
xor UO_381 (O_381,N_4872,N_4824);
and UO_382 (O_382,N_4982,N_4873);
nand UO_383 (O_383,N_4965,N_4860);
nor UO_384 (O_384,N_4844,N_4926);
nand UO_385 (O_385,N_4911,N_4874);
or UO_386 (O_386,N_4845,N_4965);
or UO_387 (O_387,N_4970,N_4818);
xnor UO_388 (O_388,N_4961,N_4861);
and UO_389 (O_389,N_4874,N_4895);
nand UO_390 (O_390,N_4991,N_4822);
or UO_391 (O_391,N_4940,N_4856);
or UO_392 (O_392,N_4875,N_4841);
and UO_393 (O_393,N_4912,N_4932);
nand UO_394 (O_394,N_4900,N_4986);
nor UO_395 (O_395,N_4981,N_4813);
nand UO_396 (O_396,N_4977,N_4880);
nand UO_397 (O_397,N_4969,N_4917);
and UO_398 (O_398,N_4908,N_4955);
nor UO_399 (O_399,N_4848,N_4980);
xor UO_400 (O_400,N_4960,N_4940);
xor UO_401 (O_401,N_4884,N_4866);
nor UO_402 (O_402,N_4865,N_4934);
xor UO_403 (O_403,N_4965,N_4949);
nand UO_404 (O_404,N_4875,N_4936);
and UO_405 (O_405,N_4892,N_4944);
xor UO_406 (O_406,N_4968,N_4807);
nor UO_407 (O_407,N_4989,N_4845);
or UO_408 (O_408,N_4964,N_4818);
or UO_409 (O_409,N_4920,N_4823);
nand UO_410 (O_410,N_4888,N_4859);
nor UO_411 (O_411,N_4824,N_4922);
or UO_412 (O_412,N_4807,N_4967);
nand UO_413 (O_413,N_4834,N_4816);
nand UO_414 (O_414,N_4869,N_4948);
or UO_415 (O_415,N_4816,N_4994);
nor UO_416 (O_416,N_4935,N_4944);
nor UO_417 (O_417,N_4908,N_4839);
nand UO_418 (O_418,N_4947,N_4809);
xnor UO_419 (O_419,N_4849,N_4917);
or UO_420 (O_420,N_4966,N_4972);
nand UO_421 (O_421,N_4800,N_4908);
and UO_422 (O_422,N_4857,N_4884);
and UO_423 (O_423,N_4957,N_4816);
nand UO_424 (O_424,N_4952,N_4814);
or UO_425 (O_425,N_4833,N_4975);
nor UO_426 (O_426,N_4808,N_4918);
or UO_427 (O_427,N_4860,N_4904);
and UO_428 (O_428,N_4872,N_4863);
nand UO_429 (O_429,N_4917,N_4972);
nand UO_430 (O_430,N_4808,N_4863);
nor UO_431 (O_431,N_4821,N_4916);
nor UO_432 (O_432,N_4863,N_4843);
nor UO_433 (O_433,N_4835,N_4902);
and UO_434 (O_434,N_4928,N_4921);
and UO_435 (O_435,N_4818,N_4923);
and UO_436 (O_436,N_4993,N_4828);
xor UO_437 (O_437,N_4907,N_4925);
or UO_438 (O_438,N_4814,N_4843);
xor UO_439 (O_439,N_4928,N_4957);
nand UO_440 (O_440,N_4986,N_4813);
or UO_441 (O_441,N_4909,N_4848);
and UO_442 (O_442,N_4889,N_4932);
nand UO_443 (O_443,N_4835,N_4873);
or UO_444 (O_444,N_4866,N_4904);
or UO_445 (O_445,N_4885,N_4953);
nand UO_446 (O_446,N_4982,N_4958);
nor UO_447 (O_447,N_4940,N_4941);
nor UO_448 (O_448,N_4898,N_4802);
nor UO_449 (O_449,N_4826,N_4874);
and UO_450 (O_450,N_4969,N_4896);
xor UO_451 (O_451,N_4837,N_4999);
nor UO_452 (O_452,N_4825,N_4866);
and UO_453 (O_453,N_4927,N_4952);
xor UO_454 (O_454,N_4834,N_4837);
nor UO_455 (O_455,N_4981,N_4973);
nand UO_456 (O_456,N_4848,N_4987);
xnor UO_457 (O_457,N_4891,N_4932);
nor UO_458 (O_458,N_4957,N_4912);
nand UO_459 (O_459,N_4981,N_4803);
nor UO_460 (O_460,N_4914,N_4864);
nor UO_461 (O_461,N_4857,N_4837);
xor UO_462 (O_462,N_4914,N_4935);
xor UO_463 (O_463,N_4874,N_4846);
nand UO_464 (O_464,N_4962,N_4838);
nor UO_465 (O_465,N_4924,N_4807);
xor UO_466 (O_466,N_4903,N_4828);
and UO_467 (O_467,N_4991,N_4835);
nor UO_468 (O_468,N_4959,N_4819);
nand UO_469 (O_469,N_4974,N_4981);
or UO_470 (O_470,N_4986,N_4892);
or UO_471 (O_471,N_4834,N_4932);
nor UO_472 (O_472,N_4808,N_4900);
and UO_473 (O_473,N_4985,N_4886);
xnor UO_474 (O_474,N_4947,N_4802);
and UO_475 (O_475,N_4834,N_4809);
xor UO_476 (O_476,N_4874,N_4948);
or UO_477 (O_477,N_4936,N_4941);
nand UO_478 (O_478,N_4873,N_4854);
or UO_479 (O_479,N_4983,N_4830);
and UO_480 (O_480,N_4825,N_4907);
nor UO_481 (O_481,N_4939,N_4823);
nor UO_482 (O_482,N_4870,N_4878);
and UO_483 (O_483,N_4934,N_4959);
or UO_484 (O_484,N_4947,N_4903);
nand UO_485 (O_485,N_4883,N_4819);
xnor UO_486 (O_486,N_4943,N_4953);
nor UO_487 (O_487,N_4933,N_4810);
and UO_488 (O_488,N_4818,N_4889);
nor UO_489 (O_489,N_4911,N_4963);
nor UO_490 (O_490,N_4895,N_4835);
and UO_491 (O_491,N_4884,N_4997);
nand UO_492 (O_492,N_4951,N_4987);
nand UO_493 (O_493,N_4924,N_4898);
nand UO_494 (O_494,N_4888,N_4867);
xor UO_495 (O_495,N_4994,N_4856);
and UO_496 (O_496,N_4931,N_4978);
nor UO_497 (O_497,N_4917,N_4898);
nand UO_498 (O_498,N_4965,N_4888);
or UO_499 (O_499,N_4838,N_4936);
xnor UO_500 (O_500,N_4918,N_4841);
and UO_501 (O_501,N_4959,N_4841);
nand UO_502 (O_502,N_4801,N_4872);
and UO_503 (O_503,N_4993,N_4830);
nand UO_504 (O_504,N_4901,N_4979);
and UO_505 (O_505,N_4936,N_4925);
and UO_506 (O_506,N_4934,N_4933);
and UO_507 (O_507,N_4833,N_4807);
and UO_508 (O_508,N_4966,N_4962);
and UO_509 (O_509,N_4985,N_4852);
or UO_510 (O_510,N_4982,N_4914);
nor UO_511 (O_511,N_4970,N_4966);
xor UO_512 (O_512,N_4883,N_4995);
and UO_513 (O_513,N_4886,N_4940);
nand UO_514 (O_514,N_4874,N_4873);
nor UO_515 (O_515,N_4810,N_4953);
nand UO_516 (O_516,N_4809,N_4940);
or UO_517 (O_517,N_4979,N_4848);
nand UO_518 (O_518,N_4818,N_4830);
xor UO_519 (O_519,N_4840,N_4801);
and UO_520 (O_520,N_4837,N_4848);
or UO_521 (O_521,N_4923,N_4946);
xor UO_522 (O_522,N_4846,N_4819);
nor UO_523 (O_523,N_4970,N_4981);
nor UO_524 (O_524,N_4944,N_4820);
xnor UO_525 (O_525,N_4891,N_4870);
xnor UO_526 (O_526,N_4817,N_4939);
or UO_527 (O_527,N_4955,N_4940);
nand UO_528 (O_528,N_4807,N_4969);
or UO_529 (O_529,N_4890,N_4978);
and UO_530 (O_530,N_4830,N_4924);
and UO_531 (O_531,N_4986,N_4945);
nor UO_532 (O_532,N_4810,N_4969);
nor UO_533 (O_533,N_4976,N_4948);
or UO_534 (O_534,N_4805,N_4811);
and UO_535 (O_535,N_4972,N_4875);
nor UO_536 (O_536,N_4831,N_4872);
and UO_537 (O_537,N_4919,N_4969);
nor UO_538 (O_538,N_4895,N_4930);
and UO_539 (O_539,N_4875,N_4935);
nand UO_540 (O_540,N_4972,N_4925);
xnor UO_541 (O_541,N_4825,N_4892);
xnor UO_542 (O_542,N_4936,N_4977);
nand UO_543 (O_543,N_4901,N_4851);
nand UO_544 (O_544,N_4926,N_4869);
nand UO_545 (O_545,N_4895,N_4887);
xor UO_546 (O_546,N_4932,N_4968);
or UO_547 (O_547,N_4995,N_4962);
and UO_548 (O_548,N_4994,N_4803);
xor UO_549 (O_549,N_4857,N_4936);
xnor UO_550 (O_550,N_4871,N_4898);
and UO_551 (O_551,N_4860,N_4912);
nor UO_552 (O_552,N_4901,N_4959);
or UO_553 (O_553,N_4814,N_4888);
and UO_554 (O_554,N_4853,N_4922);
nor UO_555 (O_555,N_4899,N_4832);
nand UO_556 (O_556,N_4837,N_4987);
nor UO_557 (O_557,N_4838,N_4844);
and UO_558 (O_558,N_4929,N_4859);
nand UO_559 (O_559,N_4965,N_4867);
and UO_560 (O_560,N_4940,N_4894);
nor UO_561 (O_561,N_4914,N_4804);
nand UO_562 (O_562,N_4935,N_4831);
xor UO_563 (O_563,N_4974,N_4896);
xnor UO_564 (O_564,N_4953,N_4814);
or UO_565 (O_565,N_4994,N_4916);
nor UO_566 (O_566,N_4961,N_4911);
xor UO_567 (O_567,N_4968,N_4964);
nand UO_568 (O_568,N_4921,N_4871);
and UO_569 (O_569,N_4961,N_4955);
and UO_570 (O_570,N_4902,N_4871);
xor UO_571 (O_571,N_4858,N_4934);
and UO_572 (O_572,N_4841,N_4881);
nor UO_573 (O_573,N_4824,N_4855);
and UO_574 (O_574,N_4877,N_4860);
or UO_575 (O_575,N_4814,N_4974);
or UO_576 (O_576,N_4920,N_4865);
xor UO_577 (O_577,N_4827,N_4916);
or UO_578 (O_578,N_4801,N_4903);
nand UO_579 (O_579,N_4916,N_4977);
xor UO_580 (O_580,N_4849,N_4883);
nor UO_581 (O_581,N_4991,N_4969);
nor UO_582 (O_582,N_4901,N_4925);
and UO_583 (O_583,N_4960,N_4969);
or UO_584 (O_584,N_4873,N_4845);
nor UO_585 (O_585,N_4827,N_4838);
xnor UO_586 (O_586,N_4967,N_4895);
or UO_587 (O_587,N_4986,N_4855);
nand UO_588 (O_588,N_4958,N_4977);
and UO_589 (O_589,N_4887,N_4914);
and UO_590 (O_590,N_4884,N_4937);
xor UO_591 (O_591,N_4845,N_4988);
nand UO_592 (O_592,N_4840,N_4882);
or UO_593 (O_593,N_4984,N_4867);
xnor UO_594 (O_594,N_4903,N_4852);
nor UO_595 (O_595,N_4921,N_4979);
nand UO_596 (O_596,N_4922,N_4951);
xor UO_597 (O_597,N_4801,N_4893);
and UO_598 (O_598,N_4852,N_4883);
and UO_599 (O_599,N_4982,N_4898);
or UO_600 (O_600,N_4852,N_4887);
xor UO_601 (O_601,N_4941,N_4834);
and UO_602 (O_602,N_4984,N_4944);
or UO_603 (O_603,N_4889,N_4843);
and UO_604 (O_604,N_4920,N_4951);
nand UO_605 (O_605,N_4919,N_4845);
nand UO_606 (O_606,N_4985,N_4824);
xnor UO_607 (O_607,N_4943,N_4882);
nand UO_608 (O_608,N_4975,N_4891);
xor UO_609 (O_609,N_4951,N_4812);
nor UO_610 (O_610,N_4882,N_4835);
or UO_611 (O_611,N_4861,N_4922);
nand UO_612 (O_612,N_4847,N_4904);
or UO_613 (O_613,N_4928,N_4832);
and UO_614 (O_614,N_4976,N_4937);
nor UO_615 (O_615,N_4822,N_4928);
or UO_616 (O_616,N_4834,N_4943);
nor UO_617 (O_617,N_4821,N_4999);
nand UO_618 (O_618,N_4839,N_4911);
or UO_619 (O_619,N_4814,N_4899);
or UO_620 (O_620,N_4877,N_4986);
xor UO_621 (O_621,N_4826,N_4888);
nor UO_622 (O_622,N_4824,N_4862);
and UO_623 (O_623,N_4826,N_4868);
nor UO_624 (O_624,N_4821,N_4966);
and UO_625 (O_625,N_4990,N_4982);
or UO_626 (O_626,N_4831,N_4972);
and UO_627 (O_627,N_4944,N_4839);
nand UO_628 (O_628,N_4893,N_4928);
and UO_629 (O_629,N_4827,N_4826);
xor UO_630 (O_630,N_4849,N_4842);
and UO_631 (O_631,N_4967,N_4983);
nand UO_632 (O_632,N_4874,N_4967);
xor UO_633 (O_633,N_4905,N_4889);
nand UO_634 (O_634,N_4900,N_4969);
xnor UO_635 (O_635,N_4900,N_4911);
or UO_636 (O_636,N_4931,N_4955);
xor UO_637 (O_637,N_4950,N_4815);
nand UO_638 (O_638,N_4845,N_4979);
xnor UO_639 (O_639,N_4945,N_4858);
and UO_640 (O_640,N_4850,N_4953);
nor UO_641 (O_641,N_4993,N_4895);
xnor UO_642 (O_642,N_4822,N_4813);
and UO_643 (O_643,N_4997,N_4975);
or UO_644 (O_644,N_4815,N_4881);
or UO_645 (O_645,N_4998,N_4959);
and UO_646 (O_646,N_4840,N_4910);
nor UO_647 (O_647,N_4863,N_4820);
xnor UO_648 (O_648,N_4809,N_4830);
or UO_649 (O_649,N_4994,N_4895);
or UO_650 (O_650,N_4881,N_4890);
or UO_651 (O_651,N_4893,N_4932);
nand UO_652 (O_652,N_4827,N_4831);
or UO_653 (O_653,N_4898,N_4970);
or UO_654 (O_654,N_4967,N_4963);
and UO_655 (O_655,N_4819,N_4810);
xor UO_656 (O_656,N_4867,N_4862);
and UO_657 (O_657,N_4942,N_4802);
nand UO_658 (O_658,N_4836,N_4831);
xnor UO_659 (O_659,N_4912,N_4834);
or UO_660 (O_660,N_4990,N_4800);
nor UO_661 (O_661,N_4878,N_4800);
xnor UO_662 (O_662,N_4916,N_4897);
or UO_663 (O_663,N_4816,N_4870);
xnor UO_664 (O_664,N_4901,N_4828);
or UO_665 (O_665,N_4854,N_4991);
xor UO_666 (O_666,N_4997,N_4831);
nor UO_667 (O_667,N_4932,N_4942);
or UO_668 (O_668,N_4897,N_4911);
and UO_669 (O_669,N_4849,N_4959);
nor UO_670 (O_670,N_4815,N_4985);
or UO_671 (O_671,N_4935,N_4977);
xnor UO_672 (O_672,N_4974,N_4803);
nor UO_673 (O_673,N_4990,N_4976);
xnor UO_674 (O_674,N_4925,N_4876);
nor UO_675 (O_675,N_4818,N_4854);
and UO_676 (O_676,N_4830,N_4966);
or UO_677 (O_677,N_4895,N_4836);
nor UO_678 (O_678,N_4983,N_4951);
xor UO_679 (O_679,N_4953,N_4976);
or UO_680 (O_680,N_4856,N_4805);
nand UO_681 (O_681,N_4939,N_4804);
xnor UO_682 (O_682,N_4960,N_4868);
nor UO_683 (O_683,N_4811,N_4934);
xnor UO_684 (O_684,N_4960,N_4973);
and UO_685 (O_685,N_4933,N_4896);
or UO_686 (O_686,N_4837,N_4995);
nor UO_687 (O_687,N_4907,N_4823);
or UO_688 (O_688,N_4895,N_4850);
nor UO_689 (O_689,N_4899,N_4864);
nor UO_690 (O_690,N_4938,N_4803);
or UO_691 (O_691,N_4978,N_4873);
or UO_692 (O_692,N_4964,N_4950);
nor UO_693 (O_693,N_4928,N_4828);
and UO_694 (O_694,N_4985,N_4855);
xor UO_695 (O_695,N_4802,N_4864);
or UO_696 (O_696,N_4958,N_4839);
and UO_697 (O_697,N_4862,N_4828);
and UO_698 (O_698,N_4948,N_4824);
or UO_699 (O_699,N_4992,N_4984);
nor UO_700 (O_700,N_4889,N_4912);
nor UO_701 (O_701,N_4996,N_4871);
or UO_702 (O_702,N_4952,N_4951);
nand UO_703 (O_703,N_4962,N_4981);
nor UO_704 (O_704,N_4873,N_4914);
nor UO_705 (O_705,N_4879,N_4907);
nor UO_706 (O_706,N_4885,N_4908);
nor UO_707 (O_707,N_4876,N_4883);
nand UO_708 (O_708,N_4958,N_4889);
and UO_709 (O_709,N_4804,N_4815);
nand UO_710 (O_710,N_4869,N_4984);
and UO_711 (O_711,N_4864,N_4921);
or UO_712 (O_712,N_4862,N_4900);
nor UO_713 (O_713,N_4839,N_4986);
and UO_714 (O_714,N_4860,N_4906);
nor UO_715 (O_715,N_4996,N_4821);
nor UO_716 (O_716,N_4814,N_4940);
or UO_717 (O_717,N_4963,N_4894);
or UO_718 (O_718,N_4903,N_4803);
xnor UO_719 (O_719,N_4989,N_4905);
nor UO_720 (O_720,N_4934,N_4835);
and UO_721 (O_721,N_4956,N_4829);
nand UO_722 (O_722,N_4898,N_4938);
or UO_723 (O_723,N_4979,N_4893);
and UO_724 (O_724,N_4821,N_4875);
xnor UO_725 (O_725,N_4835,N_4900);
nand UO_726 (O_726,N_4859,N_4850);
or UO_727 (O_727,N_4999,N_4846);
nand UO_728 (O_728,N_4895,N_4824);
or UO_729 (O_729,N_4810,N_4862);
nor UO_730 (O_730,N_4901,N_4801);
and UO_731 (O_731,N_4864,N_4941);
xor UO_732 (O_732,N_4939,N_4814);
nand UO_733 (O_733,N_4909,N_4970);
xnor UO_734 (O_734,N_4831,N_4898);
or UO_735 (O_735,N_4961,N_4827);
nand UO_736 (O_736,N_4958,N_4907);
nor UO_737 (O_737,N_4888,N_4989);
or UO_738 (O_738,N_4852,N_4938);
or UO_739 (O_739,N_4935,N_4863);
or UO_740 (O_740,N_4813,N_4878);
nor UO_741 (O_741,N_4924,N_4938);
and UO_742 (O_742,N_4961,N_4834);
nor UO_743 (O_743,N_4967,N_4961);
nand UO_744 (O_744,N_4950,N_4840);
nand UO_745 (O_745,N_4869,N_4805);
or UO_746 (O_746,N_4955,N_4993);
and UO_747 (O_747,N_4951,N_4879);
or UO_748 (O_748,N_4877,N_4912);
nand UO_749 (O_749,N_4848,N_4950);
and UO_750 (O_750,N_4893,N_4991);
or UO_751 (O_751,N_4819,N_4830);
or UO_752 (O_752,N_4839,N_4928);
and UO_753 (O_753,N_4950,N_4932);
and UO_754 (O_754,N_4986,N_4841);
nand UO_755 (O_755,N_4852,N_4919);
nor UO_756 (O_756,N_4970,N_4831);
or UO_757 (O_757,N_4863,N_4801);
nand UO_758 (O_758,N_4990,N_4986);
or UO_759 (O_759,N_4901,N_4915);
xor UO_760 (O_760,N_4925,N_4999);
and UO_761 (O_761,N_4968,N_4991);
nor UO_762 (O_762,N_4932,N_4904);
and UO_763 (O_763,N_4912,N_4906);
nand UO_764 (O_764,N_4804,N_4856);
and UO_765 (O_765,N_4882,N_4836);
or UO_766 (O_766,N_4839,N_4953);
nand UO_767 (O_767,N_4807,N_4962);
nand UO_768 (O_768,N_4954,N_4992);
and UO_769 (O_769,N_4991,N_4882);
nor UO_770 (O_770,N_4868,N_4860);
nand UO_771 (O_771,N_4892,N_4932);
nand UO_772 (O_772,N_4802,N_4858);
and UO_773 (O_773,N_4963,N_4881);
nand UO_774 (O_774,N_4972,N_4950);
nor UO_775 (O_775,N_4855,N_4829);
nor UO_776 (O_776,N_4970,N_4821);
nor UO_777 (O_777,N_4906,N_4833);
xor UO_778 (O_778,N_4985,N_4951);
or UO_779 (O_779,N_4858,N_4963);
and UO_780 (O_780,N_4850,N_4947);
or UO_781 (O_781,N_4995,N_4834);
nor UO_782 (O_782,N_4902,N_4989);
or UO_783 (O_783,N_4956,N_4974);
nand UO_784 (O_784,N_4980,N_4892);
or UO_785 (O_785,N_4838,N_4840);
xor UO_786 (O_786,N_4863,N_4829);
and UO_787 (O_787,N_4885,N_4840);
and UO_788 (O_788,N_4912,N_4856);
nor UO_789 (O_789,N_4982,N_4957);
and UO_790 (O_790,N_4923,N_4848);
nand UO_791 (O_791,N_4965,N_4982);
or UO_792 (O_792,N_4850,N_4980);
or UO_793 (O_793,N_4925,N_4802);
and UO_794 (O_794,N_4967,N_4871);
xor UO_795 (O_795,N_4818,N_4819);
or UO_796 (O_796,N_4971,N_4840);
or UO_797 (O_797,N_4833,N_4921);
xnor UO_798 (O_798,N_4805,N_4999);
nor UO_799 (O_799,N_4965,N_4961);
or UO_800 (O_800,N_4886,N_4893);
xor UO_801 (O_801,N_4920,N_4973);
nor UO_802 (O_802,N_4940,N_4860);
nor UO_803 (O_803,N_4834,N_4841);
xor UO_804 (O_804,N_4969,N_4916);
nand UO_805 (O_805,N_4824,N_4888);
or UO_806 (O_806,N_4900,N_4881);
or UO_807 (O_807,N_4932,N_4951);
and UO_808 (O_808,N_4965,N_4821);
xnor UO_809 (O_809,N_4935,N_4876);
and UO_810 (O_810,N_4948,N_4890);
and UO_811 (O_811,N_4978,N_4833);
or UO_812 (O_812,N_4852,N_4817);
and UO_813 (O_813,N_4820,N_4806);
or UO_814 (O_814,N_4831,N_4941);
nor UO_815 (O_815,N_4835,N_4852);
or UO_816 (O_816,N_4940,N_4861);
nor UO_817 (O_817,N_4828,N_4932);
nand UO_818 (O_818,N_4993,N_4880);
nor UO_819 (O_819,N_4910,N_4955);
and UO_820 (O_820,N_4814,N_4835);
nor UO_821 (O_821,N_4860,N_4803);
xor UO_822 (O_822,N_4855,N_4889);
nor UO_823 (O_823,N_4821,N_4937);
nor UO_824 (O_824,N_4974,N_4866);
and UO_825 (O_825,N_4838,N_4958);
or UO_826 (O_826,N_4917,N_4968);
or UO_827 (O_827,N_4935,N_4922);
or UO_828 (O_828,N_4940,N_4991);
and UO_829 (O_829,N_4865,N_4949);
nand UO_830 (O_830,N_4881,N_4847);
and UO_831 (O_831,N_4813,N_4883);
nor UO_832 (O_832,N_4820,N_4813);
and UO_833 (O_833,N_4883,N_4924);
or UO_834 (O_834,N_4897,N_4839);
and UO_835 (O_835,N_4951,N_4910);
nor UO_836 (O_836,N_4801,N_4813);
nand UO_837 (O_837,N_4802,N_4895);
xnor UO_838 (O_838,N_4913,N_4905);
and UO_839 (O_839,N_4940,N_4885);
or UO_840 (O_840,N_4891,N_4944);
xnor UO_841 (O_841,N_4932,N_4914);
nor UO_842 (O_842,N_4851,N_4969);
or UO_843 (O_843,N_4889,N_4888);
and UO_844 (O_844,N_4995,N_4983);
nor UO_845 (O_845,N_4827,N_4861);
and UO_846 (O_846,N_4881,N_4883);
nor UO_847 (O_847,N_4897,N_4913);
nor UO_848 (O_848,N_4909,N_4859);
nor UO_849 (O_849,N_4816,N_4826);
nand UO_850 (O_850,N_4949,N_4872);
nor UO_851 (O_851,N_4934,N_4891);
nor UO_852 (O_852,N_4995,N_4933);
or UO_853 (O_853,N_4809,N_4821);
and UO_854 (O_854,N_4870,N_4946);
nor UO_855 (O_855,N_4929,N_4996);
xnor UO_856 (O_856,N_4837,N_4818);
or UO_857 (O_857,N_4822,N_4962);
xnor UO_858 (O_858,N_4990,N_4856);
nor UO_859 (O_859,N_4970,N_4995);
and UO_860 (O_860,N_4827,N_4897);
xnor UO_861 (O_861,N_4942,N_4857);
xnor UO_862 (O_862,N_4813,N_4959);
nor UO_863 (O_863,N_4933,N_4898);
nand UO_864 (O_864,N_4838,N_4888);
xnor UO_865 (O_865,N_4820,N_4987);
xnor UO_866 (O_866,N_4882,N_4994);
or UO_867 (O_867,N_4954,N_4999);
nand UO_868 (O_868,N_4965,N_4919);
xnor UO_869 (O_869,N_4846,N_4939);
xor UO_870 (O_870,N_4975,N_4926);
nand UO_871 (O_871,N_4983,N_4973);
nor UO_872 (O_872,N_4933,N_4808);
nor UO_873 (O_873,N_4860,N_4988);
nand UO_874 (O_874,N_4991,N_4942);
xor UO_875 (O_875,N_4829,N_4864);
nor UO_876 (O_876,N_4991,N_4839);
and UO_877 (O_877,N_4948,N_4891);
nand UO_878 (O_878,N_4983,N_4809);
and UO_879 (O_879,N_4840,N_4911);
xor UO_880 (O_880,N_4853,N_4939);
or UO_881 (O_881,N_4805,N_4888);
nor UO_882 (O_882,N_4809,N_4972);
or UO_883 (O_883,N_4928,N_4851);
nand UO_884 (O_884,N_4910,N_4836);
and UO_885 (O_885,N_4858,N_4953);
and UO_886 (O_886,N_4900,N_4960);
xor UO_887 (O_887,N_4822,N_4864);
and UO_888 (O_888,N_4966,N_4818);
xor UO_889 (O_889,N_4880,N_4922);
xnor UO_890 (O_890,N_4816,N_4907);
xnor UO_891 (O_891,N_4826,N_4803);
nor UO_892 (O_892,N_4843,N_4895);
nor UO_893 (O_893,N_4999,N_4972);
and UO_894 (O_894,N_4992,N_4961);
nor UO_895 (O_895,N_4878,N_4912);
or UO_896 (O_896,N_4882,N_4875);
nor UO_897 (O_897,N_4999,N_4966);
nor UO_898 (O_898,N_4837,N_4852);
xor UO_899 (O_899,N_4824,N_4836);
or UO_900 (O_900,N_4951,N_4949);
nand UO_901 (O_901,N_4953,N_4845);
xor UO_902 (O_902,N_4964,N_4922);
and UO_903 (O_903,N_4995,N_4898);
xor UO_904 (O_904,N_4883,N_4903);
xnor UO_905 (O_905,N_4946,N_4859);
and UO_906 (O_906,N_4841,N_4988);
or UO_907 (O_907,N_4946,N_4914);
nor UO_908 (O_908,N_4834,N_4865);
and UO_909 (O_909,N_4944,N_4863);
nand UO_910 (O_910,N_4839,N_4902);
or UO_911 (O_911,N_4833,N_4981);
nand UO_912 (O_912,N_4851,N_4939);
or UO_913 (O_913,N_4914,N_4863);
nand UO_914 (O_914,N_4973,N_4943);
or UO_915 (O_915,N_4856,N_4820);
and UO_916 (O_916,N_4998,N_4881);
and UO_917 (O_917,N_4808,N_4892);
and UO_918 (O_918,N_4978,N_4910);
xnor UO_919 (O_919,N_4887,N_4904);
nand UO_920 (O_920,N_4802,N_4933);
or UO_921 (O_921,N_4976,N_4877);
xor UO_922 (O_922,N_4940,N_4916);
or UO_923 (O_923,N_4895,N_4944);
and UO_924 (O_924,N_4822,N_4908);
and UO_925 (O_925,N_4859,N_4819);
xnor UO_926 (O_926,N_4991,N_4842);
or UO_927 (O_927,N_4868,N_4891);
xor UO_928 (O_928,N_4958,N_4971);
nor UO_929 (O_929,N_4977,N_4822);
or UO_930 (O_930,N_4832,N_4920);
nand UO_931 (O_931,N_4810,N_4966);
nand UO_932 (O_932,N_4932,N_4818);
and UO_933 (O_933,N_4999,N_4965);
nor UO_934 (O_934,N_4825,N_4913);
nand UO_935 (O_935,N_4807,N_4885);
nand UO_936 (O_936,N_4838,N_4997);
and UO_937 (O_937,N_4948,N_4900);
or UO_938 (O_938,N_4997,N_4925);
xnor UO_939 (O_939,N_4960,N_4832);
nand UO_940 (O_940,N_4865,N_4923);
nand UO_941 (O_941,N_4966,N_4816);
xnor UO_942 (O_942,N_4941,N_4921);
nor UO_943 (O_943,N_4900,N_4997);
xnor UO_944 (O_944,N_4826,N_4936);
nor UO_945 (O_945,N_4906,N_4894);
nand UO_946 (O_946,N_4994,N_4944);
nand UO_947 (O_947,N_4907,N_4880);
and UO_948 (O_948,N_4932,N_4902);
xor UO_949 (O_949,N_4975,N_4980);
nor UO_950 (O_950,N_4938,N_4979);
xor UO_951 (O_951,N_4996,N_4904);
and UO_952 (O_952,N_4896,N_4963);
nor UO_953 (O_953,N_4966,N_4964);
xor UO_954 (O_954,N_4972,N_4835);
nor UO_955 (O_955,N_4989,N_4973);
nor UO_956 (O_956,N_4924,N_4834);
or UO_957 (O_957,N_4829,N_4860);
nor UO_958 (O_958,N_4922,N_4889);
or UO_959 (O_959,N_4894,N_4808);
nand UO_960 (O_960,N_4802,N_4844);
or UO_961 (O_961,N_4974,N_4859);
xnor UO_962 (O_962,N_4937,N_4855);
nor UO_963 (O_963,N_4959,N_4809);
nor UO_964 (O_964,N_4887,N_4889);
or UO_965 (O_965,N_4986,N_4880);
and UO_966 (O_966,N_4987,N_4935);
and UO_967 (O_967,N_4846,N_4873);
nor UO_968 (O_968,N_4929,N_4833);
xor UO_969 (O_969,N_4862,N_4856);
xor UO_970 (O_970,N_4946,N_4879);
nor UO_971 (O_971,N_4939,N_4985);
nand UO_972 (O_972,N_4855,N_4813);
xnor UO_973 (O_973,N_4933,N_4844);
xor UO_974 (O_974,N_4973,N_4864);
or UO_975 (O_975,N_4963,N_4900);
and UO_976 (O_976,N_4927,N_4848);
and UO_977 (O_977,N_4864,N_4845);
nor UO_978 (O_978,N_4806,N_4828);
nor UO_979 (O_979,N_4894,N_4964);
and UO_980 (O_980,N_4832,N_4839);
and UO_981 (O_981,N_4844,N_4908);
nand UO_982 (O_982,N_4905,N_4892);
or UO_983 (O_983,N_4926,N_4910);
and UO_984 (O_984,N_4852,N_4987);
xnor UO_985 (O_985,N_4831,N_4999);
and UO_986 (O_986,N_4912,N_4893);
or UO_987 (O_987,N_4937,N_4852);
xor UO_988 (O_988,N_4820,N_4945);
and UO_989 (O_989,N_4901,N_4809);
and UO_990 (O_990,N_4895,N_4902);
and UO_991 (O_991,N_4991,N_4890);
nor UO_992 (O_992,N_4917,N_4802);
nand UO_993 (O_993,N_4800,N_4917);
and UO_994 (O_994,N_4969,N_4951);
or UO_995 (O_995,N_4990,N_4854);
xnor UO_996 (O_996,N_4954,N_4979);
xnor UO_997 (O_997,N_4811,N_4863);
and UO_998 (O_998,N_4995,N_4951);
or UO_999 (O_999,N_4950,N_4819);
endmodule