module basic_1000_10000_1500_5_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_846,In_784);
nand U1 (N_1,In_217,In_964);
xor U2 (N_2,In_622,In_441);
and U3 (N_3,In_838,In_799);
or U4 (N_4,In_228,In_718);
or U5 (N_5,In_797,In_35);
nor U6 (N_6,In_956,In_743);
xor U7 (N_7,In_316,In_648);
and U8 (N_8,In_330,In_485);
xor U9 (N_9,In_963,In_407);
xnor U10 (N_10,In_56,In_917);
or U11 (N_11,In_844,In_971);
nand U12 (N_12,In_147,In_763);
and U13 (N_13,In_238,In_195);
or U14 (N_14,In_438,In_654);
xor U15 (N_15,In_570,In_786);
xnor U16 (N_16,In_978,In_153);
or U17 (N_17,In_841,In_290);
or U18 (N_18,In_873,In_31);
nor U19 (N_19,In_976,In_883);
and U20 (N_20,In_564,In_588);
nor U21 (N_21,In_89,In_311);
nor U22 (N_22,In_600,In_794);
xor U23 (N_23,In_855,In_853);
xor U24 (N_24,In_875,In_33);
nand U25 (N_25,In_867,In_244);
nand U26 (N_26,In_504,In_440);
xnor U27 (N_27,In_674,In_443);
xnor U28 (N_28,In_966,In_858);
or U29 (N_29,In_691,In_833);
xor U30 (N_30,In_327,In_542);
xor U31 (N_31,In_302,In_211);
xor U32 (N_32,In_519,In_744);
nor U33 (N_33,In_126,In_641);
xor U34 (N_34,In_116,In_493);
xnor U35 (N_35,In_948,In_909);
xor U36 (N_36,In_977,In_901);
xor U37 (N_37,In_673,In_307);
nor U38 (N_38,In_111,In_986);
xor U39 (N_39,In_732,In_262);
nor U40 (N_40,In_52,In_605);
and U41 (N_41,In_677,In_466);
or U42 (N_42,In_907,In_606);
and U43 (N_43,In_240,In_706);
xnor U44 (N_44,In_649,In_834);
nand U45 (N_45,In_903,In_27);
nor U46 (N_46,In_83,In_599);
xor U47 (N_47,In_702,In_364);
nor U48 (N_48,In_406,In_630);
nor U49 (N_49,In_765,In_224);
nor U50 (N_50,In_480,In_270);
and U51 (N_51,In_3,In_132);
xnor U52 (N_52,In_420,In_719);
xor U53 (N_53,In_814,In_950);
nor U54 (N_54,In_124,In_617);
nand U55 (N_55,In_879,In_453);
nand U56 (N_56,In_513,In_386);
and U57 (N_57,In_762,In_435);
nand U58 (N_58,In_292,In_468);
and U59 (N_59,In_467,In_220);
nand U60 (N_60,In_698,In_457);
or U61 (N_61,In_81,In_106);
and U62 (N_62,In_87,In_8);
nor U63 (N_63,In_996,In_144);
and U64 (N_64,In_852,In_534);
or U65 (N_65,In_297,In_676);
or U66 (N_66,In_395,In_821);
nor U67 (N_67,In_491,In_614);
nand U68 (N_68,In_573,In_989);
xnor U69 (N_69,In_824,In_768);
nand U70 (N_70,In_358,In_965);
nor U71 (N_71,In_304,In_496);
nand U72 (N_72,In_260,In_105);
xnor U73 (N_73,In_612,In_635);
nand U74 (N_74,In_384,In_162);
or U75 (N_75,In_701,In_456);
and U76 (N_76,In_350,In_816);
or U77 (N_77,In_526,In_792);
nor U78 (N_78,In_382,In_968);
or U79 (N_79,In_227,In_766);
nand U80 (N_80,In_159,In_334);
nor U81 (N_81,In_157,In_323);
xnor U82 (N_82,In_957,In_512);
xor U83 (N_83,In_587,In_708);
nor U84 (N_84,In_865,In_626);
or U85 (N_85,In_695,In_775);
and U86 (N_86,In_773,In_121);
nand U87 (N_87,In_138,In_923);
or U88 (N_88,In_390,In_114);
and U89 (N_89,In_403,In_325);
nor U90 (N_90,In_442,In_843);
xnor U91 (N_91,In_990,In_926);
nor U92 (N_92,In_608,In_548);
nand U93 (N_93,In_284,In_886);
nor U94 (N_94,In_688,In_394);
nor U95 (N_95,In_857,In_300);
or U96 (N_96,In_51,In_280);
nand U97 (N_97,In_409,In_528);
nand U98 (N_98,In_631,In_679);
or U99 (N_99,In_954,In_835);
or U100 (N_100,In_722,In_259);
nor U101 (N_101,In_748,In_827);
or U102 (N_102,In_992,In_177);
or U103 (N_103,In_267,In_585);
nor U104 (N_104,In_417,In_984);
xnor U105 (N_105,In_357,In_269);
and U106 (N_106,In_46,In_815);
and U107 (N_107,In_699,In_642);
or U108 (N_108,In_200,In_789);
and U109 (N_109,In_139,In_283);
and U110 (N_110,In_632,In_680);
nand U111 (N_111,In_532,In_595);
xor U112 (N_112,In_980,In_724);
nand U113 (N_113,In_7,In_991);
nor U114 (N_114,In_837,In_825);
nor U115 (N_115,In_484,In_222);
and U116 (N_116,In_309,In_374);
nor U117 (N_117,In_900,In_940);
xnor U118 (N_118,In_308,In_94);
or U119 (N_119,In_876,In_783);
and U120 (N_120,In_850,In_800);
or U121 (N_121,In_749,In_319);
nand U122 (N_122,In_158,In_385);
or U123 (N_123,In_524,In_434);
xor U124 (N_124,In_932,In_776);
nor U125 (N_125,In_801,In_717);
or U126 (N_126,In_6,In_100);
nor U127 (N_127,In_970,In_165);
nand U128 (N_128,In_771,In_554);
nor U129 (N_129,In_296,In_368);
xnor U130 (N_130,In_348,In_671);
or U131 (N_131,In_757,In_263);
or U132 (N_132,In_933,In_753);
and U133 (N_133,In_819,In_919);
nand U134 (N_134,In_565,In_329);
and U135 (N_135,In_870,In_198);
or U136 (N_136,In_878,In_34);
and U137 (N_137,In_1,In_667);
and U138 (N_138,In_143,In_333);
and U139 (N_139,In_337,In_481);
nand U140 (N_140,In_232,In_508);
xnor U141 (N_141,In_133,In_666);
xor U142 (N_142,In_258,In_298);
nor U143 (N_143,In_320,In_877);
nand U144 (N_144,In_938,In_944);
and U145 (N_145,In_725,In_507);
or U146 (N_146,In_633,In_469);
nand U147 (N_147,In_988,In_99);
nor U148 (N_148,In_890,In_772);
and U149 (N_149,In_119,In_328);
nand U150 (N_150,In_285,In_710);
and U151 (N_151,In_301,In_663);
and U152 (N_152,In_709,In_860);
and U153 (N_153,In_346,In_571);
and U154 (N_154,In_317,In_893);
or U155 (N_155,In_108,In_445);
xor U156 (N_156,In_233,In_125);
or U157 (N_157,In_859,In_498);
or U158 (N_158,In_49,In_416);
nor U159 (N_159,In_60,In_922);
or U160 (N_160,In_908,In_905);
nor U161 (N_161,In_408,In_70);
and U162 (N_162,In_643,In_546);
xor U163 (N_163,In_539,In_74);
or U164 (N_164,In_619,In_823);
and U165 (N_165,In_525,In_896);
and U166 (N_166,In_345,In_73);
xor U167 (N_167,In_175,In_229);
xnor U168 (N_168,In_482,In_904);
and U169 (N_169,In_577,In_711);
or U170 (N_170,In_609,In_354);
xor U171 (N_171,In_785,In_192);
nand U172 (N_172,In_418,In_254);
or U173 (N_173,In_646,In_377);
or U174 (N_174,In_523,In_979);
nand U175 (N_175,In_665,In_104);
xnor U176 (N_176,In_912,In_118);
nand U177 (N_177,In_898,In_93);
nor U178 (N_178,In_193,In_471);
xnor U179 (N_179,In_312,In_90);
xor U180 (N_180,In_848,In_840);
or U181 (N_181,In_14,In_172);
and U182 (N_182,In_576,In_624);
or U183 (N_183,In_194,In_117);
or U184 (N_184,In_553,In_266);
and U185 (N_185,In_109,In_826);
or U186 (N_186,In_128,In_537);
nor U187 (N_187,In_129,In_552);
nand U188 (N_188,In_378,In_758);
or U189 (N_189,In_560,In_282);
and U190 (N_190,In_914,In_340);
xnor U191 (N_191,In_683,In_734);
nor U192 (N_192,In_77,In_943);
and U193 (N_193,In_804,In_874);
xnor U194 (N_194,In_461,In_592);
or U195 (N_195,In_343,In_568);
or U196 (N_196,In_656,In_313);
xor U197 (N_197,In_974,In_444);
nor U198 (N_198,In_97,In_563);
nor U199 (N_199,In_154,In_847);
or U200 (N_200,In_293,In_221);
and U201 (N_201,In_741,In_218);
xor U202 (N_202,In_934,In_255);
and U203 (N_203,In_809,In_366);
nor U204 (N_204,In_64,In_433);
nor U205 (N_205,In_767,In_413);
or U206 (N_206,In_169,In_715);
and U207 (N_207,In_180,In_399);
xnor U208 (N_208,In_72,In_419);
nand U209 (N_209,In_245,In_616);
and U210 (N_210,In_851,In_289);
or U211 (N_211,In_644,In_306);
or U212 (N_212,In_22,In_726);
and U213 (N_213,In_55,In_183);
and U214 (N_214,In_729,In_291);
nand U215 (N_215,In_370,In_149);
and U216 (N_216,In_120,In_98);
and U217 (N_217,In_470,In_995);
and U218 (N_218,In_361,In_286);
xor U219 (N_219,In_806,In_69);
xor U220 (N_220,In_854,In_798);
xor U221 (N_221,In_376,In_618);
or U222 (N_222,In_2,In_54);
nor U223 (N_223,In_892,In_557);
and U224 (N_224,In_716,In_359);
xnor U225 (N_225,In_705,In_235);
nor U226 (N_226,In_728,In_25);
nand U227 (N_227,In_130,In_778);
and U228 (N_228,In_520,In_547);
and U229 (N_229,In_448,In_272);
xor U230 (N_230,In_911,In_439);
xnor U231 (N_231,In_845,In_521);
or U232 (N_232,In_182,In_566);
nor U233 (N_233,In_655,In_59);
and U234 (N_234,In_20,In_856);
xnor U235 (N_235,In_223,In_381);
and U236 (N_236,In_92,In_492);
and U237 (N_237,In_899,In_431);
xnor U238 (N_238,In_582,In_488);
or U239 (N_239,In_536,In_246);
nand U240 (N_240,In_13,In_723);
and U241 (N_241,In_603,In_700);
and U242 (N_242,In_322,In_959);
or U243 (N_243,In_953,In_146);
or U244 (N_244,In_43,In_915);
nor U245 (N_245,In_829,In_682);
or U246 (N_246,In_897,In_115);
xnor U247 (N_247,In_16,In_199);
nor U248 (N_248,In_602,In_868);
and U249 (N_249,In_181,In_730);
xor U250 (N_250,In_985,In_424);
or U251 (N_251,In_812,In_342);
xnor U252 (N_252,In_459,In_86);
or U253 (N_253,In_91,In_264);
nand U254 (N_254,In_610,In_315);
or U255 (N_255,In_279,In_380);
or U256 (N_256,In_805,In_48);
or U257 (N_257,In_131,In_414);
and U258 (N_258,In_392,In_339);
and U259 (N_259,In_662,In_379);
and U260 (N_260,In_372,In_754);
nand U261 (N_261,In_37,In_449);
and U262 (N_262,In_880,In_972);
and U263 (N_263,In_347,In_551);
or U264 (N_264,In_212,In_982);
nor U265 (N_265,In_249,In_415);
xnor U266 (N_266,In_822,In_659);
nand U267 (N_267,In_692,In_428);
nand U268 (N_268,In_63,In_363);
or U269 (N_269,In_405,In_866);
and U270 (N_270,In_353,In_733);
and U271 (N_271,In_447,In_38);
nand U272 (N_272,In_894,In_696);
nor U273 (N_273,In_593,In_787);
nor U274 (N_274,In_769,In_951);
nand U275 (N_275,In_882,In_47);
and U276 (N_276,In_261,In_518);
nand U277 (N_277,In_425,In_881);
and U278 (N_278,In_678,In_672);
or U279 (N_279,In_236,In_774);
nor U280 (N_280,In_556,In_973);
or U281 (N_281,In_360,In_849);
xor U282 (N_282,In_650,In_9);
and U283 (N_283,In_697,In_490);
xor U284 (N_284,In_755,In_681);
and U285 (N_285,In_895,In_574);
nor U286 (N_286,In_205,In_945);
nand U287 (N_287,In_949,In_225);
or U288 (N_288,In_615,In_994);
and U289 (N_289,In_113,In_450);
nand U290 (N_290,In_863,In_651);
nand U291 (N_291,In_53,In_216);
xor U292 (N_292,In_44,In_476);
nand U293 (N_293,In_828,In_201);
nand U294 (N_294,In_522,In_179);
or U295 (N_295,In_527,In_503);
and U296 (N_296,In_26,In_421);
or U297 (N_297,In_742,In_188);
or U298 (N_298,In_367,In_36);
or U299 (N_299,In_497,In_740);
nor U300 (N_300,In_242,In_167);
nor U301 (N_301,In_176,In_10);
nor U302 (N_302,In_777,In_214);
xnor U303 (N_303,In_462,In_918);
nor U304 (N_304,In_684,In_924);
xor U305 (N_305,In_640,In_84);
or U306 (N_306,In_4,In_685);
nand U307 (N_307,In_253,In_18);
xnor U308 (N_308,In_460,In_930);
and U309 (N_309,In_952,In_668);
and U310 (N_310,In_714,In_861);
nand U311 (N_311,In_356,In_23);
nor U312 (N_312,In_430,In_647);
xnor U313 (N_313,In_135,In_543);
nand U314 (N_314,In_318,In_190);
and U315 (N_315,In_920,In_278);
xnor U316 (N_316,In_652,In_598);
xor U317 (N_317,In_475,In_997);
or U318 (N_318,In_590,In_219);
and U319 (N_319,In_436,In_506);
or U320 (N_320,In_910,In_514);
nor U321 (N_321,In_184,In_540);
nor U322 (N_322,In_398,In_30);
xor U323 (N_323,In_40,In_887);
nor U324 (N_324,In_832,In_362);
nor U325 (N_325,In_21,In_657);
nor U326 (N_326,In_810,In_538);
or U327 (N_327,In_45,In_530);
nor U328 (N_328,In_210,In_830);
and U329 (N_329,In_299,In_243);
or U330 (N_330,In_487,In_738);
nor U331 (N_331,In_955,In_281);
or U332 (N_332,In_929,In_401);
and U333 (N_333,In_969,In_693);
xnor U334 (N_334,In_795,In_226);
nor U335 (N_335,In_5,In_545);
nand U336 (N_336,In_256,In_151);
xnor U337 (N_337,In_597,In_474);
or U338 (N_338,In_101,In_141);
nor U339 (N_339,In_727,In_426);
and U340 (N_340,In_842,In_687);
nor U341 (N_341,In_669,In_75);
nand U342 (N_342,In_721,In_276);
or U343 (N_343,In_931,In_925);
nor U344 (N_344,In_134,In_621);
and U345 (N_345,In_287,In_41);
and U346 (N_346,In_661,In_817);
xor U347 (N_347,In_96,In_884);
nor U348 (N_348,In_501,In_209);
and U349 (N_349,In_203,In_704);
xor U350 (N_350,In_889,In_639);
and U351 (N_351,In_446,In_752);
nor U352 (N_352,In_637,In_625);
nor U353 (N_353,In_250,In_464);
or U354 (N_354,In_562,In_839);
or U355 (N_355,In_782,In_248);
and U356 (N_356,In_387,In_591);
and U357 (N_357,In_24,In_185);
nor U358 (N_358,In_103,In_349);
nor U359 (N_359,In_981,In_234);
or U360 (N_360,In_230,In_790);
xor U361 (N_361,In_735,In_636);
nor U362 (N_362,In_375,In_578);
or U363 (N_363,In_288,In_906);
or U364 (N_364,In_383,In_80);
nand U365 (N_365,In_294,In_252);
and U366 (N_366,In_561,In_472);
nand U367 (N_367,In_458,In_916);
nand U368 (N_368,In_544,In_788);
xor U369 (N_369,In_831,In_432);
nor U370 (N_370,In_336,In_935);
or U371 (N_371,In_170,In_739);
nand U372 (N_372,In_921,In_65);
and U373 (N_373,In_509,In_66);
and U374 (N_374,In_888,In_601);
nor U375 (N_375,In_196,In_869);
nand U376 (N_376,In_596,In_477);
nand U377 (N_377,In_770,In_197);
nor U378 (N_378,In_690,In_510);
nor U379 (N_379,In_483,In_107);
and U380 (N_380,In_611,In_168);
xor U381 (N_381,In_712,In_215);
xnor U382 (N_382,In_529,In_17);
or U383 (N_383,In_781,In_579);
nand U384 (N_384,In_265,In_303);
and U385 (N_385,In_555,In_620);
and U386 (N_386,In_32,In_331);
xor U387 (N_387,In_764,In_166);
or U388 (N_388,In_173,In_533);
nand U389 (N_389,In_422,In_397);
nand U390 (N_390,In_628,In_670);
and U391 (N_391,In_231,In_452);
nand U392 (N_392,In_891,In_112);
or U393 (N_393,In_946,In_463);
and U394 (N_394,In_156,In_737);
nor U395 (N_395,In_499,In_796);
nor U396 (N_396,In_204,In_171);
and U397 (N_397,In_206,In_29);
nand U398 (N_398,In_960,In_102);
and U399 (N_399,In_213,In_164);
nor U400 (N_400,In_404,In_505);
or U401 (N_401,In_85,In_275);
xor U402 (N_402,In_19,In_836);
or U403 (N_403,In_584,In_324);
and U404 (N_404,In_567,In_396);
or U405 (N_405,In_277,In_928);
or U406 (N_406,In_658,In_79);
nor U407 (N_407,In_50,In_335);
xor U408 (N_408,In_885,In_241);
nor U409 (N_409,In_427,In_160);
and U410 (N_410,In_402,In_607);
or U411 (N_411,In_140,In_237);
xnor U412 (N_412,In_594,In_987);
xor U413 (N_413,In_412,In_746);
or U414 (N_414,In_604,In_186);
and U415 (N_415,In_163,In_793);
or U416 (N_416,In_207,In_295);
and U417 (N_417,In_67,In_486);
and U418 (N_418,In_78,In_627);
or U419 (N_419,In_756,In_110);
nand U420 (N_420,In_760,In_638);
nor U421 (N_421,In_583,In_150);
nor U422 (N_422,In_489,In_411);
xor U423 (N_423,In_962,In_549);
nand U424 (N_424,In_88,In_811);
and U425 (N_425,In_541,In_818);
and U426 (N_426,In_0,In_454);
xnor U427 (N_427,In_208,In_967);
nor U428 (N_428,In_473,In_451);
nor U429 (N_429,In_558,In_759);
nand U430 (N_430,In_613,In_983);
or U431 (N_431,In_62,In_780);
nor U432 (N_432,In_58,In_707);
nand U433 (N_433,In_586,In_161);
nand U434 (N_434,In_122,In_393);
nor U435 (N_435,In_502,In_391);
nor U436 (N_436,In_268,In_127);
nor U437 (N_437,In_15,In_515);
xnor U438 (N_438,In_57,In_731);
or U439 (N_439,In_189,In_429);
nor U440 (N_440,In_257,In_572);
nand U441 (N_441,In_629,In_12);
or U442 (N_442,In_191,In_747);
nand U443 (N_443,In_751,In_388);
nand U444 (N_444,In_437,In_95);
or U445 (N_445,In_148,In_961);
or U446 (N_446,In_511,In_937);
xnor U447 (N_447,In_137,In_251);
xnor U448 (N_448,In_145,In_271);
nand U449 (N_449,In_465,In_713);
nor U450 (N_450,In_802,In_239);
and U451 (N_451,In_305,In_569);
or U452 (N_452,In_371,In_479);
xnor U453 (N_453,In_664,In_580);
nor U454 (N_454,In_675,In_936);
nand U455 (N_455,In_820,In_338);
or U456 (N_456,In_39,In_689);
nor U457 (N_457,In_273,In_142);
nor U458 (N_458,In_750,In_939);
nor U459 (N_459,In_581,In_589);
xor U460 (N_460,In_634,In_351);
nand U461 (N_461,In_28,In_314);
nand U462 (N_462,In_500,In_202);
nand U463 (N_463,In_535,In_178);
and U464 (N_464,In_61,In_947);
and U465 (N_465,In_975,In_373);
and U466 (N_466,In_645,In_400);
nand U467 (N_467,In_913,In_745);
nor U468 (N_468,In_247,In_761);
nor U469 (N_469,In_862,In_82);
or U470 (N_470,In_155,In_187);
or U471 (N_471,In_410,In_872);
or U472 (N_472,In_71,In_495);
xnor U473 (N_473,In_365,In_369);
nand U474 (N_474,In_152,In_927);
and U475 (N_475,In_326,In_321);
nand U476 (N_476,In_344,In_864);
or U477 (N_477,In_123,In_341);
nand U478 (N_478,In_998,In_807);
and U479 (N_479,In_653,In_791);
xnor U480 (N_480,In_389,In_531);
nand U481 (N_481,In_686,In_310);
nand U482 (N_482,In_455,In_68);
xnor U483 (N_483,In_136,In_736);
nand U484 (N_484,In_42,In_779);
nor U485 (N_485,In_871,In_274);
xnor U486 (N_486,In_550,In_494);
and U487 (N_487,In_516,In_941);
and U488 (N_488,In_623,In_174);
and U489 (N_489,In_902,In_423);
nor U490 (N_490,In_808,In_703);
xnor U491 (N_491,In_720,In_11);
xnor U492 (N_492,In_993,In_813);
xnor U493 (N_493,In_76,In_332);
or U494 (N_494,In_355,In_559);
xnor U495 (N_495,In_942,In_958);
nor U496 (N_496,In_352,In_803);
nand U497 (N_497,In_999,In_660);
and U498 (N_498,In_478,In_575);
or U499 (N_499,In_517,In_694);
nand U500 (N_500,In_147,In_314);
xnor U501 (N_501,In_80,In_547);
nor U502 (N_502,In_148,In_657);
xnor U503 (N_503,In_535,In_774);
or U504 (N_504,In_923,In_879);
xnor U505 (N_505,In_336,In_397);
or U506 (N_506,In_468,In_371);
or U507 (N_507,In_435,In_922);
nor U508 (N_508,In_747,In_759);
nand U509 (N_509,In_537,In_664);
and U510 (N_510,In_809,In_874);
nand U511 (N_511,In_643,In_372);
or U512 (N_512,In_665,In_801);
nand U513 (N_513,In_530,In_234);
and U514 (N_514,In_8,In_486);
and U515 (N_515,In_176,In_29);
and U516 (N_516,In_705,In_366);
and U517 (N_517,In_864,In_105);
nand U518 (N_518,In_261,In_668);
nand U519 (N_519,In_853,In_34);
xor U520 (N_520,In_49,In_957);
nand U521 (N_521,In_882,In_524);
nand U522 (N_522,In_418,In_838);
nor U523 (N_523,In_585,In_72);
xnor U524 (N_524,In_369,In_995);
nor U525 (N_525,In_394,In_92);
nor U526 (N_526,In_847,In_176);
nor U527 (N_527,In_885,In_126);
nand U528 (N_528,In_619,In_424);
nand U529 (N_529,In_803,In_112);
nand U530 (N_530,In_585,In_936);
nor U531 (N_531,In_938,In_428);
and U532 (N_532,In_474,In_936);
and U533 (N_533,In_723,In_260);
and U534 (N_534,In_53,In_968);
nor U535 (N_535,In_463,In_108);
nor U536 (N_536,In_572,In_210);
nor U537 (N_537,In_237,In_733);
or U538 (N_538,In_310,In_145);
and U539 (N_539,In_865,In_307);
nor U540 (N_540,In_965,In_930);
and U541 (N_541,In_567,In_554);
and U542 (N_542,In_351,In_376);
xor U543 (N_543,In_806,In_566);
and U544 (N_544,In_161,In_641);
and U545 (N_545,In_785,In_368);
nand U546 (N_546,In_551,In_448);
and U547 (N_547,In_558,In_236);
or U548 (N_548,In_481,In_845);
xnor U549 (N_549,In_423,In_387);
or U550 (N_550,In_358,In_426);
or U551 (N_551,In_333,In_816);
xor U552 (N_552,In_359,In_399);
and U553 (N_553,In_142,In_51);
nor U554 (N_554,In_853,In_630);
nor U555 (N_555,In_988,In_91);
xnor U556 (N_556,In_282,In_157);
nor U557 (N_557,In_842,In_765);
or U558 (N_558,In_95,In_390);
and U559 (N_559,In_537,In_84);
nand U560 (N_560,In_93,In_772);
or U561 (N_561,In_71,In_975);
nor U562 (N_562,In_321,In_113);
or U563 (N_563,In_578,In_920);
nor U564 (N_564,In_763,In_917);
and U565 (N_565,In_348,In_379);
or U566 (N_566,In_826,In_623);
nor U567 (N_567,In_194,In_418);
and U568 (N_568,In_925,In_825);
or U569 (N_569,In_971,In_739);
and U570 (N_570,In_274,In_843);
xor U571 (N_571,In_805,In_794);
nand U572 (N_572,In_495,In_589);
and U573 (N_573,In_298,In_648);
and U574 (N_574,In_707,In_638);
nor U575 (N_575,In_299,In_113);
xor U576 (N_576,In_717,In_547);
xor U577 (N_577,In_75,In_512);
and U578 (N_578,In_526,In_176);
or U579 (N_579,In_591,In_431);
nor U580 (N_580,In_232,In_715);
nand U581 (N_581,In_731,In_302);
and U582 (N_582,In_118,In_490);
or U583 (N_583,In_801,In_583);
or U584 (N_584,In_484,In_147);
nand U585 (N_585,In_855,In_498);
or U586 (N_586,In_32,In_212);
or U587 (N_587,In_564,In_576);
nor U588 (N_588,In_280,In_9);
or U589 (N_589,In_986,In_257);
nand U590 (N_590,In_733,In_962);
xnor U591 (N_591,In_528,In_236);
or U592 (N_592,In_409,In_332);
nand U593 (N_593,In_624,In_300);
or U594 (N_594,In_730,In_260);
or U595 (N_595,In_389,In_399);
or U596 (N_596,In_860,In_374);
and U597 (N_597,In_979,In_711);
and U598 (N_598,In_86,In_376);
nand U599 (N_599,In_985,In_18);
xor U600 (N_600,In_745,In_35);
nor U601 (N_601,In_687,In_59);
xnor U602 (N_602,In_116,In_525);
xnor U603 (N_603,In_569,In_189);
or U604 (N_604,In_673,In_857);
and U605 (N_605,In_482,In_440);
or U606 (N_606,In_390,In_301);
and U607 (N_607,In_383,In_106);
nor U608 (N_608,In_300,In_728);
and U609 (N_609,In_562,In_642);
nor U610 (N_610,In_249,In_40);
or U611 (N_611,In_539,In_208);
nand U612 (N_612,In_609,In_981);
nand U613 (N_613,In_808,In_123);
xor U614 (N_614,In_369,In_63);
nand U615 (N_615,In_313,In_290);
nor U616 (N_616,In_521,In_348);
nor U617 (N_617,In_59,In_492);
and U618 (N_618,In_876,In_772);
xor U619 (N_619,In_362,In_879);
nand U620 (N_620,In_874,In_883);
xor U621 (N_621,In_118,In_732);
nor U622 (N_622,In_5,In_145);
and U623 (N_623,In_736,In_56);
and U624 (N_624,In_245,In_241);
xnor U625 (N_625,In_202,In_640);
or U626 (N_626,In_664,In_423);
or U627 (N_627,In_186,In_119);
and U628 (N_628,In_384,In_698);
and U629 (N_629,In_981,In_371);
xor U630 (N_630,In_315,In_401);
nand U631 (N_631,In_100,In_354);
nor U632 (N_632,In_893,In_344);
or U633 (N_633,In_754,In_70);
or U634 (N_634,In_591,In_567);
or U635 (N_635,In_594,In_920);
nor U636 (N_636,In_951,In_808);
and U637 (N_637,In_528,In_192);
or U638 (N_638,In_578,In_616);
nor U639 (N_639,In_182,In_811);
xor U640 (N_640,In_727,In_369);
xnor U641 (N_641,In_264,In_155);
nand U642 (N_642,In_618,In_87);
nand U643 (N_643,In_999,In_411);
nand U644 (N_644,In_824,In_51);
and U645 (N_645,In_162,In_477);
and U646 (N_646,In_882,In_595);
nor U647 (N_647,In_329,In_582);
or U648 (N_648,In_759,In_446);
nand U649 (N_649,In_753,In_790);
nand U650 (N_650,In_994,In_816);
nor U651 (N_651,In_394,In_553);
and U652 (N_652,In_566,In_630);
and U653 (N_653,In_785,In_605);
nor U654 (N_654,In_955,In_908);
xnor U655 (N_655,In_996,In_183);
and U656 (N_656,In_617,In_387);
nand U657 (N_657,In_77,In_155);
xnor U658 (N_658,In_165,In_625);
nor U659 (N_659,In_351,In_367);
nor U660 (N_660,In_41,In_637);
xnor U661 (N_661,In_238,In_691);
nand U662 (N_662,In_843,In_634);
xor U663 (N_663,In_607,In_530);
and U664 (N_664,In_324,In_610);
nor U665 (N_665,In_59,In_500);
xor U666 (N_666,In_346,In_216);
nor U667 (N_667,In_678,In_249);
or U668 (N_668,In_23,In_997);
xor U669 (N_669,In_223,In_822);
nor U670 (N_670,In_792,In_833);
or U671 (N_671,In_650,In_646);
or U672 (N_672,In_189,In_347);
nand U673 (N_673,In_326,In_643);
nand U674 (N_674,In_677,In_732);
nand U675 (N_675,In_915,In_557);
or U676 (N_676,In_823,In_383);
xor U677 (N_677,In_843,In_516);
xor U678 (N_678,In_970,In_450);
or U679 (N_679,In_26,In_155);
nor U680 (N_680,In_893,In_403);
xor U681 (N_681,In_883,In_104);
xnor U682 (N_682,In_948,In_729);
xor U683 (N_683,In_622,In_531);
and U684 (N_684,In_81,In_218);
nor U685 (N_685,In_996,In_47);
or U686 (N_686,In_633,In_141);
or U687 (N_687,In_571,In_69);
and U688 (N_688,In_127,In_515);
nor U689 (N_689,In_976,In_687);
and U690 (N_690,In_562,In_604);
and U691 (N_691,In_900,In_975);
nor U692 (N_692,In_393,In_457);
or U693 (N_693,In_57,In_942);
xor U694 (N_694,In_513,In_918);
nor U695 (N_695,In_761,In_385);
or U696 (N_696,In_106,In_361);
and U697 (N_697,In_641,In_962);
xnor U698 (N_698,In_208,In_894);
or U699 (N_699,In_578,In_610);
xor U700 (N_700,In_661,In_181);
and U701 (N_701,In_230,In_548);
nand U702 (N_702,In_482,In_417);
or U703 (N_703,In_927,In_470);
nand U704 (N_704,In_138,In_179);
nand U705 (N_705,In_644,In_566);
nand U706 (N_706,In_925,In_194);
xnor U707 (N_707,In_189,In_350);
or U708 (N_708,In_890,In_153);
xnor U709 (N_709,In_540,In_854);
nor U710 (N_710,In_257,In_721);
and U711 (N_711,In_288,In_493);
nor U712 (N_712,In_832,In_904);
xnor U713 (N_713,In_540,In_382);
nand U714 (N_714,In_255,In_309);
or U715 (N_715,In_83,In_17);
or U716 (N_716,In_9,In_250);
xnor U717 (N_717,In_336,In_342);
nor U718 (N_718,In_139,In_985);
xor U719 (N_719,In_293,In_884);
xor U720 (N_720,In_335,In_254);
xor U721 (N_721,In_460,In_814);
xor U722 (N_722,In_632,In_812);
and U723 (N_723,In_300,In_589);
nand U724 (N_724,In_349,In_983);
and U725 (N_725,In_245,In_715);
and U726 (N_726,In_82,In_36);
and U727 (N_727,In_92,In_647);
and U728 (N_728,In_79,In_717);
nor U729 (N_729,In_886,In_452);
nor U730 (N_730,In_485,In_722);
nand U731 (N_731,In_640,In_742);
nand U732 (N_732,In_426,In_790);
nand U733 (N_733,In_635,In_964);
nor U734 (N_734,In_767,In_254);
nand U735 (N_735,In_717,In_780);
nand U736 (N_736,In_119,In_23);
and U737 (N_737,In_631,In_371);
xor U738 (N_738,In_718,In_449);
nor U739 (N_739,In_749,In_776);
nor U740 (N_740,In_154,In_231);
xor U741 (N_741,In_114,In_703);
nand U742 (N_742,In_478,In_6);
xor U743 (N_743,In_874,In_944);
nor U744 (N_744,In_125,In_548);
nor U745 (N_745,In_39,In_787);
nand U746 (N_746,In_711,In_92);
nor U747 (N_747,In_527,In_60);
nor U748 (N_748,In_386,In_918);
nand U749 (N_749,In_560,In_375);
or U750 (N_750,In_558,In_900);
xor U751 (N_751,In_857,In_982);
or U752 (N_752,In_41,In_253);
nand U753 (N_753,In_939,In_763);
or U754 (N_754,In_842,In_811);
and U755 (N_755,In_915,In_146);
nor U756 (N_756,In_242,In_647);
nor U757 (N_757,In_285,In_496);
xnor U758 (N_758,In_736,In_626);
nor U759 (N_759,In_529,In_948);
or U760 (N_760,In_625,In_216);
nand U761 (N_761,In_351,In_953);
xor U762 (N_762,In_875,In_377);
or U763 (N_763,In_605,In_104);
nor U764 (N_764,In_393,In_207);
and U765 (N_765,In_346,In_749);
nor U766 (N_766,In_179,In_296);
nand U767 (N_767,In_231,In_728);
or U768 (N_768,In_885,In_542);
xnor U769 (N_769,In_794,In_484);
and U770 (N_770,In_632,In_606);
xor U771 (N_771,In_636,In_644);
nand U772 (N_772,In_860,In_980);
or U773 (N_773,In_175,In_194);
nand U774 (N_774,In_469,In_199);
or U775 (N_775,In_99,In_750);
xnor U776 (N_776,In_901,In_325);
nor U777 (N_777,In_653,In_28);
or U778 (N_778,In_845,In_664);
nor U779 (N_779,In_793,In_720);
or U780 (N_780,In_224,In_422);
xor U781 (N_781,In_244,In_764);
or U782 (N_782,In_853,In_449);
xnor U783 (N_783,In_342,In_960);
nand U784 (N_784,In_478,In_422);
nand U785 (N_785,In_628,In_263);
nand U786 (N_786,In_627,In_450);
nand U787 (N_787,In_591,In_170);
and U788 (N_788,In_696,In_788);
and U789 (N_789,In_674,In_768);
xor U790 (N_790,In_204,In_858);
or U791 (N_791,In_121,In_379);
and U792 (N_792,In_488,In_382);
or U793 (N_793,In_242,In_727);
and U794 (N_794,In_388,In_490);
xnor U795 (N_795,In_823,In_250);
nand U796 (N_796,In_956,In_922);
or U797 (N_797,In_136,In_179);
nand U798 (N_798,In_512,In_676);
xor U799 (N_799,In_236,In_708);
xnor U800 (N_800,In_888,In_80);
xnor U801 (N_801,In_398,In_519);
and U802 (N_802,In_258,In_713);
and U803 (N_803,In_578,In_17);
nor U804 (N_804,In_604,In_579);
or U805 (N_805,In_795,In_558);
or U806 (N_806,In_593,In_771);
xor U807 (N_807,In_705,In_762);
nand U808 (N_808,In_726,In_592);
nor U809 (N_809,In_109,In_981);
nor U810 (N_810,In_139,In_973);
xor U811 (N_811,In_999,In_343);
nand U812 (N_812,In_874,In_556);
and U813 (N_813,In_790,In_337);
xor U814 (N_814,In_870,In_582);
nor U815 (N_815,In_428,In_353);
xor U816 (N_816,In_327,In_323);
nor U817 (N_817,In_238,In_899);
xor U818 (N_818,In_111,In_175);
nor U819 (N_819,In_30,In_315);
or U820 (N_820,In_886,In_547);
nor U821 (N_821,In_754,In_417);
nand U822 (N_822,In_364,In_39);
or U823 (N_823,In_512,In_680);
xnor U824 (N_824,In_481,In_223);
nor U825 (N_825,In_438,In_890);
or U826 (N_826,In_850,In_464);
xnor U827 (N_827,In_745,In_68);
nand U828 (N_828,In_122,In_386);
nand U829 (N_829,In_572,In_380);
xor U830 (N_830,In_406,In_211);
or U831 (N_831,In_622,In_522);
or U832 (N_832,In_317,In_319);
nand U833 (N_833,In_107,In_276);
nand U834 (N_834,In_426,In_219);
and U835 (N_835,In_891,In_547);
or U836 (N_836,In_139,In_724);
xor U837 (N_837,In_314,In_693);
or U838 (N_838,In_755,In_239);
nor U839 (N_839,In_984,In_575);
nand U840 (N_840,In_836,In_583);
nand U841 (N_841,In_901,In_590);
nand U842 (N_842,In_84,In_950);
xnor U843 (N_843,In_141,In_31);
or U844 (N_844,In_437,In_616);
xnor U845 (N_845,In_826,In_823);
nand U846 (N_846,In_568,In_207);
nor U847 (N_847,In_6,In_989);
xnor U848 (N_848,In_343,In_938);
nor U849 (N_849,In_548,In_378);
xnor U850 (N_850,In_69,In_768);
nor U851 (N_851,In_73,In_334);
or U852 (N_852,In_499,In_154);
or U853 (N_853,In_842,In_940);
and U854 (N_854,In_998,In_216);
or U855 (N_855,In_673,In_668);
or U856 (N_856,In_271,In_207);
nor U857 (N_857,In_708,In_335);
or U858 (N_858,In_966,In_683);
xor U859 (N_859,In_859,In_231);
xor U860 (N_860,In_618,In_693);
nor U861 (N_861,In_406,In_262);
and U862 (N_862,In_235,In_586);
and U863 (N_863,In_452,In_614);
nor U864 (N_864,In_182,In_235);
xnor U865 (N_865,In_964,In_859);
nand U866 (N_866,In_657,In_925);
and U867 (N_867,In_206,In_857);
xnor U868 (N_868,In_464,In_304);
xor U869 (N_869,In_624,In_429);
and U870 (N_870,In_922,In_217);
nand U871 (N_871,In_108,In_793);
nor U872 (N_872,In_682,In_134);
nand U873 (N_873,In_458,In_162);
nor U874 (N_874,In_907,In_496);
and U875 (N_875,In_901,In_493);
xor U876 (N_876,In_928,In_522);
xnor U877 (N_877,In_557,In_74);
nor U878 (N_878,In_789,In_610);
or U879 (N_879,In_353,In_361);
nand U880 (N_880,In_153,In_830);
and U881 (N_881,In_862,In_815);
and U882 (N_882,In_501,In_372);
or U883 (N_883,In_723,In_870);
nor U884 (N_884,In_845,In_823);
and U885 (N_885,In_275,In_578);
or U886 (N_886,In_738,In_914);
nand U887 (N_887,In_811,In_215);
and U888 (N_888,In_649,In_177);
or U889 (N_889,In_946,In_370);
xnor U890 (N_890,In_126,In_79);
nor U891 (N_891,In_877,In_244);
nand U892 (N_892,In_829,In_985);
and U893 (N_893,In_566,In_49);
xnor U894 (N_894,In_11,In_731);
nand U895 (N_895,In_654,In_535);
nor U896 (N_896,In_278,In_390);
xnor U897 (N_897,In_952,In_620);
nor U898 (N_898,In_352,In_660);
nand U899 (N_899,In_866,In_58);
nor U900 (N_900,In_291,In_294);
xnor U901 (N_901,In_329,In_869);
nor U902 (N_902,In_470,In_563);
nand U903 (N_903,In_639,In_124);
nor U904 (N_904,In_23,In_773);
or U905 (N_905,In_377,In_771);
nor U906 (N_906,In_727,In_661);
nor U907 (N_907,In_608,In_959);
nand U908 (N_908,In_246,In_530);
xor U909 (N_909,In_557,In_285);
nand U910 (N_910,In_808,In_974);
nand U911 (N_911,In_333,In_176);
nor U912 (N_912,In_491,In_259);
or U913 (N_913,In_482,In_387);
xor U914 (N_914,In_899,In_493);
xnor U915 (N_915,In_729,In_609);
or U916 (N_916,In_950,In_524);
nor U917 (N_917,In_923,In_590);
and U918 (N_918,In_41,In_361);
or U919 (N_919,In_933,In_956);
nand U920 (N_920,In_120,In_871);
xor U921 (N_921,In_193,In_743);
xnor U922 (N_922,In_614,In_346);
or U923 (N_923,In_522,In_584);
xor U924 (N_924,In_971,In_411);
nor U925 (N_925,In_3,In_367);
nor U926 (N_926,In_109,In_679);
nor U927 (N_927,In_976,In_97);
nor U928 (N_928,In_715,In_428);
nor U929 (N_929,In_941,In_437);
xor U930 (N_930,In_945,In_130);
nor U931 (N_931,In_879,In_438);
nand U932 (N_932,In_421,In_239);
or U933 (N_933,In_552,In_976);
or U934 (N_934,In_475,In_367);
xor U935 (N_935,In_26,In_839);
or U936 (N_936,In_518,In_842);
or U937 (N_937,In_127,In_5);
and U938 (N_938,In_647,In_766);
nor U939 (N_939,In_141,In_438);
nor U940 (N_940,In_273,In_665);
xor U941 (N_941,In_698,In_235);
or U942 (N_942,In_813,In_171);
nor U943 (N_943,In_27,In_83);
xnor U944 (N_944,In_908,In_19);
xor U945 (N_945,In_248,In_261);
xnor U946 (N_946,In_960,In_195);
nand U947 (N_947,In_274,In_322);
nor U948 (N_948,In_437,In_971);
nand U949 (N_949,In_715,In_339);
nor U950 (N_950,In_968,In_301);
nand U951 (N_951,In_87,In_31);
xnor U952 (N_952,In_280,In_343);
and U953 (N_953,In_652,In_34);
and U954 (N_954,In_531,In_760);
and U955 (N_955,In_31,In_165);
and U956 (N_956,In_603,In_402);
and U957 (N_957,In_166,In_529);
or U958 (N_958,In_961,In_879);
nor U959 (N_959,In_730,In_768);
nand U960 (N_960,In_812,In_360);
and U961 (N_961,In_102,In_925);
xnor U962 (N_962,In_170,In_101);
or U963 (N_963,In_510,In_237);
and U964 (N_964,In_680,In_320);
or U965 (N_965,In_710,In_945);
or U966 (N_966,In_869,In_490);
xor U967 (N_967,In_448,In_967);
nand U968 (N_968,In_412,In_963);
nor U969 (N_969,In_772,In_55);
xor U970 (N_970,In_144,In_386);
xnor U971 (N_971,In_888,In_884);
nand U972 (N_972,In_839,In_360);
xor U973 (N_973,In_248,In_950);
nor U974 (N_974,In_490,In_456);
and U975 (N_975,In_63,In_636);
xnor U976 (N_976,In_927,In_452);
xor U977 (N_977,In_242,In_657);
nor U978 (N_978,In_987,In_382);
xnor U979 (N_979,In_115,In_173);
and U980 (N_980,In_417,In_940);
and U981 (N_981,In_186,In_796);
xnor U982 (N_982,In_878,In_577);
or U983 (N_983,In_138,In_714);
nor U984 (N_984,In_238,In_637);
or U985 (N_985,In_403,In_260);
nor U986 (N_986,In_21,In_827);
and U987 (N_987,In_718,In_719);
nand U988 (N_988,In_202,In_723);
nand U989 (N_989,In_567,In_463);
xnor U990 (N_990,In_347,In_908);
or U991 (N_991,In_408,In_284);
or U992 (N_992,In_889,In_781);
nand U993 (N_993,In_317,In_392);
and U994 (N_994,In_390,In_99);
or U995 (N_995,In_862,In_382);
and U996 (N_996,In_681,In_652);
or U997 (N_997,In_54,In_235);
and U998 (N_998,In_922,In_112);
and U999 (N_999,In_342,In_373);
nand U1000 (N_1000,In_824,In_686);
xor U1001 (N_1001,In_950,In_460);
or U1002 (N_1002,In_643,In_685);
nor U1003 (N_1003,In_788,In_937);
or U1004 (N_1004,In_592,In_7);
and U1005 (N_1005,In_93,In_184);
nand U1006 (N_1006,In_690,In_561);
and U1007 (N_1007,In_423,In_382);
and U1008 (N_1008,In_469,In_264);
nand U1009 (N_1009,In_731,In_480);
and U1010 (N_1010,In_205,In_154);
nor U1011 (N_1011,In_844,In_982);
and U1012 (N_1012,In_485,In_120);
or U1013 (N_1013,In_175,In_841);
nand U1014 (N_1014,In_162,In_600);
nor U1015 (N_1015,In_276,In_982);
nor U1016 (N_1016,In_674,In_25);
nand U1017 (N_1017,In_557,In_523);
and U1018 (N_1018,In_634,In_750);
and U1019 (N_1019,In_771,In_78);
nand U1020 (N_1020,In_103,In_656);
nand U1021 (N_1021,In_114,In_14);
xnor U1022 (N_1022,In_133,In_40);
nand U1023 (N_1023,In_48,In_724);
xnor U1024 (N_1024,In_152,In_473);
or U1025 (N_1025,In_435,In_651);
nand U1026 (N_1026,In_339,In_698);
and U1027 (N_1027,In_45,In_896);
nor U1028 (N_1028,In_133,In_67);
nand U1029 (N_1029,In_660,In_582);
and U1030 (N_1030,In_886,In_907);
or U1031 (N_1031,In_768,In_341);
or U1032 (N_1032,In_171,In_703);
nor U1033 (N_1033,In_180,In_75);
nor U1034 (N_1034,In_936,In_981);
and U1035 (N_1035,In_90,In_701);
or U1036 (N_1036,In_252,In_325);
nor U1037 (N_1037,In_853,In_713);
nor U1038 (N_1038,In_995,In_266);
and U1039 (N_1039,In_122,In_943);
and U1040 (N_1040,In_164,In_155);
or U1041 (N_1041,In_70,In_240);
xor U1042 (N_1042,In_131,In_760);
and U1043 (N_1043,In_414,In_158);
and U1044 (N_1044,In_955,In_340);
nand U1045 (N_1045,In_140,In_869);
or U1046 (N_1046,In_55,In_222);
xor U1047 (N_1047,In_615,In_123);
nand U1048 (N_1048,In_718,In_791);
nand U1049 (N_1049,In_629,In_318);
or U1050 (N_1050,In_167,In_115);
or U1051 (N_1051,In_321,In_14);
and U1052 (N_1052,In_708,In_638);
xor U1053 (N_1053,In_290,In_708);
xnor U1054 (N_1054,In_769,In_281);
nand U1055 (N_1055,In_88,In_831);
xnor U1056 (N_1056,In_451,In_304);
nor U1057 (N_1057,In_498,In_765);
or U1058 (N_1058,In_644,In_907);
nor U1059 (N_1059,In_103,In_618);
nand U1060 (N_1060,In_657,In_225);
nand U1061 (N_1061,In_219,In_943);
nand U1062 (N_1062,In_43,In_527);
nand U1063 (N_1063,In_441,In_612);
nand U1064 (N_1064,In_53,In_989);
xnor U1065 (N_1065,In_501,In_306);
xor U1066 (N_1066,In_396,In_512);
or U1067 (N_1067,In_162,In_807);
xnor U1068 (N_1068,In_271,In_938);
nand U1069 (N_1069,In_778,In_769);
nor U1070 (N_1070,In_241,In_660);
and U1071 (N_1071,In_113,In_95);
nor U1072 (N_1072,In_217,In_564);
xnor U1073 (N_1073,In_34,In_703);
or U1074 (N_1074,In_77,In_100);
or U1075 (N_1075,In_419,In_862);
xnor U1076 (N_1076,In_752,In_400);
and U1077 (N_1077,In_516,In_145);
xor U1078 (N_1078,In_788,In_672);
and U1079 (N_1079,In_653,In_95);
nand U1080 (N_1080,In_88,In_614);
xnor U1081 (N_1081,In_819,In_820);
nor U1082 (N_1082,In_115,In_782);
nand U1083 (N_1083,In_138,In_519);
or U1084 (N_1084,In_641,In_296);
nor U1085 (N_1085,In_203,In_832);
and U1086 (N_1086,In_746,In_880);
xor U1087 (N_1087,In_166,In_234);
and U1088 (N_1088,In_843,In_63);
nor U1089 (N_1089,In_847,In_812);
nor U1090 (N_1090,In_464,In_285);
and U1091 (N_1091,In_705,In_656);
nand U1092 (N_1092,In_329,In_597);
and U1093 (N_1093,In_856,In_165);
nor U1094 (N_1094,In_461,In_776);
nand U1095 (N_1095,In_231,In_865);
nor U1096 (N_1096,In_344,In_922);
xor U1097 (N_1097,In_10,In_49);
or U1098 (N_1098,In_300,In_4);
nand U1099 (N_1099,In_355,In_224);
nand U1100 (N_1100,In_833,In_800);
xor U1101 (N_1101,In_622,In_692);
or U1102 (N_1102,In_786,In_909);
or U1103 (N_1103,In_38,In_131);
nand U1104 (N_1104,In_966,In_701);
or U1105 (N_1105,In_954,In_744);
nand U1106 (N_1106,In_176,In_362);
and U1107 (N_1107,In_61,In_682);
nand U1108 (N_1108,In_760,In_554);
nor U1109 (N_1109,In_574,In_618);
nor U1110 (N_1110,In_138,In_195);
xnor U1111 (N_1111,In_76,In_857);
nor U1112 (N_1112,In_167,In_792);
or U1113 (N_1113,In_781,In_994);
nand U1114 (N_1114,In_198,In_279);
or U1115 (N_1115,In_690,In_224);
nand U1116 (N_1116,In_964,In_992);
nand U1117 (N_1117,In_46,In_967);
nand U1118 (N_1118,In_71,In_293);
and U1119 (N_1119,In_847,In_755);
xor U1120 (N_1120,In_736,In_909);
or U1121 (N_1121,In_449,In_638);
and U1122 (N_1122,In_553,In_814);
xor U1123 (N_1123,In_399,In_392);
and U1124 (N_1124,In_674,In_761);
or U1125 (N_1125,In_769,In_95);
nand U1126 (N_1126,In_754,In_744);
or U1127 (N_1127,In_818,In_380);
nand U1128 (N_1128,In_777,In_392);
and U1129 (N_1129,In_644,In_315);
xor U1130 (N_1130,In_763,In_860);
or U1131 (N_1131,In_762,In_510);
nor U1132 (N_1132,In_6,In_440);
nor U1133 (N_1133,In_413,In_886);
or U1134 (N_1134,In_70,In_470);
nand U1135 (N_1135,In_801,In_198);
nand U1136 (N_1136,In_177,In_935);
and U1137 (N_1137,In_674,In_571);
xor U1138 (N_1138,In_447,In_327);
or U1139 (N_1139,In_251,In_670);
nor U1140 (N_1140,In_625,In_2);
xor U1141 (N_1141,In_471,In_713);
nor U1142 (N_1142,In_762,In_103);
nor U1143 (N_1143,In_861,In_500);
nor U1144 (N_1144,In_407,In_898);
or U1145 (N_1145,In_421,In_976);
or U1146 (N_1146,In_14,In_212);
or U1147 (N_1147,In_856,In_215);
or U1148 (N_1148,In_464,In_798);
or U1149 (N_1149,In_58,In_80);
and U1150 (N_1150,In_785,In_6);
xor U1151 (N_1151,In_855,In_227);
or U1152 (N_1152,In_943,In_632);
or U1153 (N_1153,In_986,In_455);
nand U1154 (N_1154,In_248,In_191);
nand U1155 (N_1155,In_173,In_659);
xnor U1156 (N_1156,In_566,In_610);
nor U1157 (N_1157,In_481,In_112);
or U1158 (N_1158,In_221,In_387);
xnor U1159 (N_1159,In_836,In_714);
nand U1160 (N_1160,In_940,In_32);
nor U1161 (N_1161,In_738,In_21);
nor U1162 (N_1162,In_387,In_486);
and U1163 (N_1163,In_267,In_574);
or U1164 (N_1164,In_493,In_73);
xnor U1165 (N_1165,In_196,In_876);
or U1166 (N_1166,In_422,In_179);
nor U1167 (N_1167,In_806,In_339);
nor U1168 (N_1168,In_611,In_913);
nor U1169 (N_1169,In_53,In_896);
nor U1170 (N_1170,In_499,In_995);
or U1171 (N_1171,In_627,In_333);
and U1172 (N_1172,In_126,In_350);
or U1173 (N_1173,In_345,In_777);
nand U1174 (N_1174,In_384,In_860);
nor U1175 (N_1175,In_9,In_109);
nand U1176 (N_1176,In_837,In_466);
nor U1177 (N_1177,In_713,In_574);
or U1178 (N_1178,In_122,In_319);
nand U1179 (N_1179,In_331,In_436);
nand U1180 (N_1180,In_655,In_520);
xor U1181 (N_1181,In_774,In_813);
nor U1182 (N_1182,In_104,In_507);
nor U1183 (N_1183,In_535,In_585);
nor U1184 (N_1184,In_612,In_345);
xor U1185 (N_1185,In_51,In_56);
xnor U1186 (N_1186,In_984,In_656);
xnor U1187 (N_1187,In_219,In_211);
or U1188 (N_1188,In_534,In_972);
or U1189 (N_1189,In_607,In_17);
nor U1190 (N_1190,In_852,In_770);
or U1191 (N_1191,In_262,In_637);
nand U1192 (N_1192,In_234,In_581);
nand U1193 (N_1193,In_284,In_999);
or U1194 (N_1194,In_106,In_561);
nand U1195 (N_1195,In_824,In_933);
nor U1196 (N_1196,In_419,In_386);
nor U1197 (N_1197,In_410,In_548);
or U1198 (N_1198,In_759,In_407);
nor U1199 (N_1199,In_755,In_612);
xor U1200 (N_1200,In_489,In_943);
nor U1201 (N_1201,In_184,In_186);
and U1202 (N_1202,In_765,In_299);
xor U1203 (N_1203,In_379,In_761);
or U1204 (N_1204,In_511,In_73);
nand U1205 (N_1205,In_332,In_836);
and U1206 (N_1206,In_61,In_827);
and U1207 (N_1207,In_538,In_191);
xnor U1208 (N_1208,In_797,In_31);
nand U1209 (N_1209,In_999,In_725);
and U1210 (N_1210,In_588,In_108);
and U1211 (N_1211,In_250,In_870);
nand U1212 (N_1212,In_316,In_588);
xor U1213 (N_1213,In_770,In_192);
and U1214 (N_1214,In_322,In_890);
xnor U1215 (N_1215,In_68,In_829);
or U1216 (N_1216,In_523,In_466);
nor U1217 (N_1217,In_280,In_594);
nand U1218 (N_1218,In_714,In_367);
nor U1219 (N_1219,In_70,In_411);
xnor U1220 (N_1220,In_834,In_382);
xnor U1221 (N_1221,In_679,In_54);
nor U1222 (N_1222,In_782,In_747);
nor U1223 (N_1223,In_985,In_657);
and U1224 (N_1224,In_167,In_275);
xnor U1225 (N_1225,In_102,In_896);
nor U1226 (N_1226,In_257,In_158);
nand U1227 (N_1227,In_351,In_799);
nand U1228 (N_1228,In_846,In_608);
or U1229 (N_1229,In_310,In_277);
or U1230 (N_1230,In_953,In_21);
or U1231 (N_1231,In_677,In_187);
xnor U1232 (N_1232,In_962,In_726);
nand U1233 (N_1233,In_895,In_681);
or U1234 (N_1234,In_754,In_265);
or U1235 (N_1235,In_460,In_31);
nor U1236 (N_1236,In_477,In_390);
nand U1237 (N_1237,In_55,In_734);
nand U1238 (N_1238,In_805,In_415);
and U1239 (N_1239,In_224,In_416);
nor U1240 (N_1240,In_871,In_737);
nor U1241 (N_1241,In_413,In_338);
or U1242 (N_1242,In_175,In_456);
and U1243 (N_1243,In_285,In_315);
xnor U1244 (N_1244,In_867,In_967);
nand U1245 (N_1245,In_234,In_230);
xor U1246 (N_1246,In_233,In_803);
nand U1247 (N_1247,In_203,In_372);
nand U1248 (N_1248,In_510,In_47);
nor U1249 (N_1249,In_520,In_412);
or U1250 (N_1250,In_679,In_391);
or U1251 (N_1251,In_616,In_159);
nand U1252 (N_1252,In_788,In_384);
xnor U1253 (N_1253,In_997,In_663);
or U1254 (N_1254,In_189,In_55);
and U1255 (N_1255,In_312,In_206);
xor U1256 (N_1256,In_231,In_709);
xor U1257 (N_1257,In_609,In_307);
or U1258 (N_1258,In_76,In_623);
nand U1259 (N_1259,In_510,In_351);
or U1260 (N_1260,In_586,In_889);
nor U1261 (N_1261,In_815,In_385);
nand U1262 (N_1262,In_445,In_685);
nand U1263 (N_1263,In_942,In_207);
or U1264 (N_1264,In_868,In_644);
nand U1265 (N_1265,In_517,In_578);
nor U1266 (N_1266,In_896,In_12);
or U1267 (N_1267,In_417,In_600);
and U1268 (N_1268,In_762,In_487);
nand U1269 (N_1269,In_789,In_485);
xor U1270 (N_1270,In_906,In_102);
xnor U1271 (N_1271,In_356,In_298);
or U1272 (N_1272,In_269,In_389);
xor U1273 (N_1273,In_148,In_506);
and U1274 (N_1274,In_139,In_117);
nor U1275 (N_1275,In_993,In_258);
nand U1276 (N_1276,In_188,In_289);
and U1277 (N_1277,In_27,In_979);
or U1278 (N_1278,In_411,In_509);
or U1279 (N_1279,In_809,In_852);
xnor U1280 (N_1280,In_93,In_489);
xor U1281 (N_1281,In_677,In_399);
xor U1282 (N_1282,In_718,In_198);
nor U1283 (N_1283,In_812,In_837);
xor U1284 (N_1284,In_666,In_360);
and U1285 (N_1285,In_369,In_480);
xor U1286 (N_1286,In_292,In_412);
and U1287 (N_1287,In_321,In_492);
nand U1288 (N_1288,In_331,In_247);
or U1289 (N_1289,In_479,In_212);
xnor U1290 (N_1290,In_837,In_728);
or U1291 (N_1291,In_125,In_186);
or U1292 (N_1292,In_278,In_72);
nor U1293 (N_1293,In_939,In_646);
nor U1294 (N_1294,In_73,In_848);
nor U1295 (N_1295,In_939,In_290);
nand U1296 (N_1296,In_369,In_393);
or U1297 (N_1297,In_332,In_495);
nand U1298 (N_1298,In_319,In_813);
or U1299 (N_1299,In_244,In_440);
or U1300 (N_1300,In_97,In_510);
xnor U1301 (N_1301,In_857,In_587);
nand U1302 (N_1302,In_112,In_872);
nand U1303 (N_1303,In_496,In_616);
nor U1304 (N_1304,In_392,In_728);
xor U1305 (N_1305,In_407,In_584);
or U1306 (N_1306,In_941,In_521);
or U1307 (N_1307,In_1,In_411);
and U1308 (N_1308,In_466,In_227);
and U1309 (N_1309,In_769,In_687);
xnor U1310 (N_1310,In_320,In_26);
and U1311 (N_1311,In_917,In_885);
xor U1312 (N_1312,In_311,In_390);
nor U1313 (N_1313,In_903,In_721);
or U1314 (N_1314,In_128,In_846);
xnor U1315 (N_1315,In_54,In_754);
nor U1316 (N_1316,In_638,In_109);
and U1317 (N_1317,In_19,In_180);
or U1318 (N_1318,In_259,In_910);
nand U1319 (N_1319,In_716,In_513);
or U1320 (N_1320,In_998,In_982);
nand U1321 (N_1321,In_171,In_538);
nor U1322 (N_1322,In_9,In_332);
nor U1323 (N_1323,In_517,In_282);
and U1324 (N_1324,In_601,In_835);
nand U1325 (N_1325,In_129,In_176);
and U1326 (N_1326,In_287,In_40);
nand U1327 (N_1327,In_193,In_348);
xnor U1328 (N_1328,In_482,In_939);
xor U1329 (N_1329,In_113,In_126);
xnor U1330 (N_1330,In_649,In_234);
and U1331 (N_1331,In_12,In_945);
and U1332 (N_1332,In_538,In_565);
nand U1333 (N_1333,In_627,In_703);
xnor U1334 (N_1334,In_61,In_346);
and U1335 (N_1335,In_655,In_400);
nor U1336 (N_1336,In_163,In_346);
nor U1337 (N_1337,In_468,In_37);
xor U1338 (N_1338,In_648,In_868);
nor U1339 (N_1339,In_46,In_897);
and U1340 (N_1340,In_488,In_541);
nor U1341 (N_1341,In_488,In_592);
nand U1342 (N_1342,In_799,In_958);
nand U1343 (N_1343,In_21,In_878);
or U1344 (N_1344,In_433,In_720);
nand U1345 (N_1345,In_617,In_467);
or U1346 (N_1346,In_191,In_696);
nor U1347 (N_1347,In_576,In_223);
nand U1348 (N_1348,In_883,In_137);
and U1349 (N_1349,In_196,In_294);
nand U1350 (N_1350,In_547,In_104);
xnor U1351 (N_1351,In_280,In_74);
nor U1352 (N_1352,In_398,In_265);
nor U1353 (N_1353,In_569,In_664);
or U1354 (N_1354,In_111,In_585);
nand U1355 (N_1355,In_241,In_502);
xnor U1356 (N_1356,In_710,In_557);
or U1357 (N_1357,In_836,In_94);
or U1358 (N_1358,In_706,In_865);
nor U1359 (N_1359,In_926,In_329);
xor U1360 (N_1360,In_337,In_319);
or U1361 (N_1361,In_148,In_6);
and U1362 (N_1362,In_360,In_755);
and U1363 (N_1363,In_612,In_451);
nor U1364 (N_1364,In_851,In_135);
xnor U1365 (N_1365,In_470,In_438);
xnor U1366 (N_1366,In_797,In_434);
and U1367 (N_1367,In_844,In_300);
nor U1368 (N_1368,In_938,In_808);
or U1369 (N_1369,In_656,In_427);
or U1370 (N_1370,In_836,In_454);
nand U1371 (N_1371,In_793,In_522);
and U1372 (N_1372,In_9,In_496);
or U1373 (N_1373,In_658,In_911);
or U1374 (N_1374,In_595,In_719);
nor U1375 (N_1375,In_196,In_0);
xor U1376 (N_1376,In_541,In_329);
or U1377 (N_1377,In_153,In_284);
nor U1378 (N_1378,In_556,In_875);
xnor U1379 (N_1379,In_309,In_59);
nor U1380 (N_1380,In_144,In_39);
nor U1381 (N_1381,In_35,In_670);
nand U1382 (N_1382,In_867,In_399);
nand U1383 (N_1383,In_154,In_658);
nor U1384 (N_1384,In_616,In_448);
nor U1385 (N_1385,In_10,In_576);
nor U1386 (N_1386,In_556,In_127);
xor U1387 (N_1387,In_278,In_823);
xor U1388 (N_1388,In_878,In_674);
nand U1389 (N_1389,In_779,In_274);
or U1390 (N_1390,In_974,In_263);
and U1391 (N_1391,In_319,In_58);
nor U1392 (N_1392,In_188,In_10);
nor U1393 (N_1393,In_131,In_53);
xor U1394 (N_1394,In_579,In_889);
or U1395 (N_1395,In_942,In_614);
nor U1396 (N_1396,In_708,In_438);
or U1397 (N_1397,In_188,In_244);
or U1398 (N_1398,In_872,In_334);
nor U1399 (N_1399,In_959,In_419);
nand U1400 (N_1400,In_93,In_565);
nand U1401 (N_1401,In_258,In_577);
or U1402 (N_1402,In_395,In_577);
nor U1403 (N_1403,In_476,In_64);
nand U1404 (N_1404,In_90,In_353);
nor U1405 (N_1405,In_959,In_541);
nor U1406 (N_1406,In_649,In_509);
and U1407 (N_1407,In_424,In_860);
xnor U1408 (N_1408,In_706,In_888);
nand U1409 (N_1409,In_841,In_652);
xnor U1410 (N_1410,In_546,In_298);
or U1411 (N_1411,In_646,In_825);
nor U1412 (N_1412,In_938,In_936);
or U1413 (N_1413,In_326,In_734);
or U1414 (N_1414,In_37,In_102);
nand U1415 (N_1415,In_870,In_358);
and U1416 (N_1416,In_170,In_717);
nor U1417 (N_1417,In_695,In_602);
or U1418 (N_1418,In_359,In_373);
and U1419 (N_1419,In_639,In_499);
xor U1420 (N_1420,In_860,In_482);
and U1421 (N_1421,In_336,In_369);
nor U1422 (N_1422,In_535,In_324);
or U1423 (N_1423,In_40,In_418);
nand U1424 (N_1424,In_233,In_973);
nand U1425 (N_1425,In_495,In_875);
nand U1426 (N_1426,In_340,In_79);
nand U1427 (N_1427,In_477,In_353);
nor U1428 (N_1428,In_462,In_335);
nand U1429 (N_1429,In_887,In_498);
nand U1430 (N_1430,In_335,In_250);
or U1431 (N_1431,In_152,In_998);
nor U1432 (N_1432,In_759,In_779);
nor U1433 (N_1433,In_103,In_406);
nor U1434 (N_1434,In_669,In_520);
and U1435 (N_1435,In_580,In_759);
nor U1436 (N_1436,In_710,In_931);
nand U1437 (N_1437,In_102,In_490);
xor U1438 (N_1438,In_314,In_500);
xnor U1439 (N_1439,In_258,In_73);
nand U1440 (N_1440,In_480,In_964);
or U1441 (N_1441,In_854,In_85);
or U1442 (N_1442,In_525,In_426);
or U1443 (N_1443,In_824,In_237);
and U1444 (N_1444,In_798,In_598);
and U1445 (N_1445,In_512,In_893);
and U1446 (N_1446,In_391,In_505);
nor U1447 (N_1447,In_881,In_53);
or U1448 (N_1448,In_200,In_267);
or U1449 (N_1449,In_869,In_32);
nand U1450 (N_1450,In_769,In_804);
nor U1451 (N_1451,In_513,In_879);
or U1452 (N_1452,In_299,In_626);
nor U1453 (N_1453,In_370,In_389);
and U1454 (N_1454,In_627,In_880);
nor U1455 (N_1455,In_523,In_344);
nor U1456 (N_1456,In_992,In_172);
and U1457 (N_1457,In_223,In_990);
nand U1458 (N_1458,In_229,In_31);
or U1459 (N_1459,In_118,In_77);
or U1460 (N_1460,In_365,In_215);
nand U1461 (N_1461,In_209,In_792);
nor U1462 (N_1462,In_814,In_611);
and U1463 (N_1463,In_694,In_870);
and U1464 (N_1464,In_47,In_429);
xor U1465 (N_1465,In_605,In_930);
nand U1466 (N_1466,In_153,In_947);
or U1467 (N_1467,In_742,In_112);
or U1468 (N_1468,In_195,In_190);
xnor U1469 (N_1469,In_152,In_976);
xor U1470 (N_1470,In_447,In_222);
nand U1471 (N_1471,In_371,In_175);
and U1472 (N_1472,In_894,In_262);
nor U1473 (N_1473,In_52,In_430);
nand U1474 (N_1474,In_198,In_947);
nand U1475 (N_1475,In_320,In_948);
or U1476 (N_1476,In_92,In_55);
xnor U1477 (N_1477,In_719,In_689);
nand U1478 (N_1478,In_836,In_95);
xnor U1479 (N_1479,In_162,In_252);
and U1480 (N_1480,In_2,In_816);
nand U1481 (N_1481,In_634,In_987);
and U1482 (N_1482,In_379,In_67);
xor U1483 (N_1483,In_448,In_326);
xnor U1484 (N_1484,In_845,In_440);
xnor U1485 (N_1485,In_903,In_939);
nand U1486 (N_1486,In_185,In_486);
and U1487 (N_1487,In_296,In_338);
and U1488 (N_1488,In_380,In_484);
nand U1489 (N_1489,In_637,In_343);
and U1490 (N_1490,In_133,In_216);
nand U1491 (N_1491,In_994,In_761);
and U1492 (N_1492,In_671,In_309);
or U1493 (N_1493,In_868,In_280);
xor U1494 (N_1494,In_918,In_143);
xor U1495 (N_1495,In_990,In_158);
nand U1496 (N_1496,In_286,In_862);
or U1497 (N_1497,In_507,In_311);
nand U1498 (N_1498,In_585,In_315);
xnor U1499 (N_1499,In_77,In_827);
or U1500 (N_1500,In_302,In_355);
nand U1501 (N_1501,In_922,In_792);
nor U1502 (N_1502,In_644,In_413);
xnor U1503 (N_1503,In_716,In_250);
nor U1504 (N_1504,In_633,In_321);
nor U1505 (N_1505,In_483,In_799);
and U1506 (N_1506,In_660,In_273);
or U1507 (N_1507,In_146,In_567);
nand U1508 (N_1508,In_41,In_790);
or U1509 (N_1509,In_975,In_625);
or U1510 (N_1510,In_599,In_976);
nand U1511 (N_1511,In_302,In_551);
or U1512 (N_1512,In_380,In_79);
and U1513 (N_1513,In_893,In_933);
nand U1514 (N_1514,In_761,In_91);
or U1515 (N_1515,In_35,In_765);
or U1516 (N_1516,In_947,In_86);
and U1517 (N_1517,In_673,In_107);
and U1518 (N_1518,In_405,In_708);
nand U1519 (N_1519,In_587,In_854);
xor U1520 (N_1520,In_504,In_263);
nand U1521 (N_1521,In_147,In_161);
nor U1522 (N_1522,In_701,In_782);
xor U1523 (N_1523,In_165,In_580);
nor U1524 (N_1524,In_47,In_585);
nand U1525 (N_1525,In_996,In_735);
nor U1526 (N_1526,In_995,In_38);
xor U1527 (N_1527,In_35,In_237);
xor U1528 (N_1528,In_487,In_315);
and U1529 (N_1529,In_768,In_844);
and U1530 (N_1530,In_704,In_48);
xor U1531 (N_1531,In_275,In_928);
nor U1532 (N_1532,In_848,In_628);
or U1533 (N_1533,In_696,In_553);
nor U1534 (N_1534,In_442,In_306);
nor U1535 (N_1535,In_875,In_937);
and U1536 (N_1536,In_274,In_958);
or U1537 (N_1537,In_283,In_985);
nor U1538 (N_1538,In_160,In_835);
and U1539 (N_1539,In_640,In_823);
nor U1540 (N_1540,In_912,In_796);
nand U1541 (N_1541,In_655,In_121);
xnor U1542 (N_1542,In_320,In_373);
and U1543 (N_1543,In_935,In_799);
nor U1544 (N_1544,In_957,In_160);
xnor U1545 (N_1545,In_620,In_21);
or U1546 (N_1546,In_975,In_8);
or U1547 (N_1547,In_897,In_889);
nand U1548 (N_1548,In_747,In_709);
and U1549 (N_1549,In_341,In_840);
or U1550 (N_1550,In_727,In_755);
or U1551 (N_1551,In_730,In_174);
xnor U1552 (N_1552,In_865,In_818);
xor U1553 (N_1553,In_30,In_676);
or U1554 (N_1554,In_679,In_266);
nand U1555 (N_1555,In_720,In_728);
or U1556 (N_1556,In_752,In_36);
xnor U1557 (N_1557,In_699,In_307);
xor U1558 (N_1558,In_613,In_185);
nand U1559 (N_1559,In_144,In_857);
nand U1560 (N_1560,In_467,In_687);
or U1561 (N_1561,In_81,In_610);
nand U1562 (N_1562,In_702,In_730);
or U1563 (N_1563,In_303,In_242);
or U1564 (N_1564,In_600,In_977);
nand U1565 (N_1565,In_989,In_203);
nor U1566 (N_1566,In_140,In_959);
xnor U1567 (N_1567,In_579,In_697);
or U1568 (N_1568,In_671,In_448);
and U1569 (N_1569,In_314,In_184);
nor U1570 (N_1570,In_682,In_653);
and U1571 (N_1571,In_409,In_393);
nor U1572 (N_1572,In_738,In_156);
and U1573 (N_1573,In_333,In_993);
xor U1574 (N_1574,In_160,In_198);
nor U1575 (N_1575,In_956,In_600);
nand U1576 (N_1576,In_972,In_742);
nor U1577 (N_1577,In_206,In_78);
nand U1578 (N_1578,In_314,In_458);
nor U1579 (N_1579,In_520,In_391);
or U1580 (N_1580,In_640,In_678);
nand U1581 (N_1581,In_902,In_977);
and U1582 (N_1582,In_531,In_384);
or U1583 (N_1583,In_382,In_895);
nand U1584 (N_1584,In_639,In_168);
or U1585 (N_1585,In_23,In_521);
or U1586 (N_1586,In_385,In_225);
and U1587 (N_1587,In_117,In_606);
and U1588 (N_1588,In_81,In_873);
nor U1589 (N_1589,In_349,In_55);
or U1590 (N_1590,In_234,In_241);
and U1591 (N_1591,In_112,In_656);
nor U1592 (N_1592,In_590,In_531);
and U1593 (N_1593,In_104,In_168);
nor U1594 (N_1594,In_243,In_981);
and U1595 (N_1595,In_902,In_31);
nand U1596 (N_1596,In_229,In_429);
nand U1597 (N_1597,In_976,In_907);
nor U1598 (N_1598,In_275,In_24);
and U1599 (N_1599,In_353,In_233);
xor U1600 (N_1600,In_356,In_556);
or U1601 (N_1601,In_110,In_59);
or U1602 (N_1602,In_266,In_733);
nand U1603 (N_1603,In_594,In_362);
nor U1604 (N_1604,In_300,In_316);
nor U1605 (N_1605,In_915,In_879);
nor U1606 (N_1606,In_473,In_354);
or U1607 (N_1607,In_754,In_358);
nand U1608 (N_1608,In_73,In_95);
xor U1609 (N_1609,In_586,In_754);
nand U1610 (N_1610,In_787,In_373);
nor U1611 (N_1611,In_357,In_532);
and U1612 (N_1612,In_217,In_982);
nor U1613 (N_1613,In_946,In_944);
nand U1614 (N_1614,In_905,In_853);
and U1615 (N_1615,In_236,In_788);
xnor U1616 (N_1616,In_540,In_71);
nand U1617 (N_1617,In_392,In_911);
xor U1618 (N_1618,In_323,In_915);
and U1619 (N_1619,In_520,In_501);
nand U1620 (N_1620,In_308,In_431);
and U1621 (N_1621,In_432,In_166);
or U1622 (N_1622,In_652,In_764);
or U1623 (N_1623,In_643,In_633);
nand U1624 (N_1624,In_878,In_709);
nand U1625 (N_1625,In_717,In_6);
xnor U1626 (N_1626,In_51,In_82);
and U1627 (N_1627,In_295,In_62);
nor U1628 (N_1628,In_144,In_361);
or U1629 (N_1629,In_858,In_519);
nor U1630 (N_1630,In_871,In_92);
nor U1631 (N_1631,In_232,In_268);
or U1632 (N_1632,In_59,In_398);
or U1633 (N_1633,In_468,In_288);
nor U1634 (N_1634,In_585,In_704);
nor U1635 (N_1635,In_40,In_35);
nor U1636 (N_1636,In_581,In_597);
nor U1637 (N_1637,In_796,In_864);
xnor U1638 (N_1638,In_9,In_412);
or U1639 (N_1639,In_661,In_793);
nor U1640 (N_1640,In_430,In_333);
or U1641 (N_1641,In_776,In_213);
nand U1642 (N_1642,In_812,In_943);
nor U1643 (N_1643,In_594,In_24);
nand U1644 (N_1644,In_632,In_935);
nand U1645 (N_1645,In_496,In_826);
xnor U1646 (N_1646,In_501,In_875);
and U1647 (N_1647,In_986,In_766);
and U1648 (N_1648,In_311,In_990);
nand U1649 (N_1649,In_503,In_239);
or U1650 (N_1650,In_343,In_668);
nand U1651 (N_1651,In_81,In_979);
and U1652 (N_1652,In_391,In_237);
or U1653 (N_1653,In_365,In_171);
xnor U1654 (N_1654,In_282,In_554);
nand U1655 (N_1655,In_239,In_450);
and U1656 (N_1656,In_279,In_396);
nor U1657 (N_1657,In_400,In_299);
and U1658 (N_1658,In_703,In_96);
or U1659 (N_1659,In_724,In_367);
xor U1660 (N_1660,In_589,In_189);
nor U1661 (N_1661,In_574,In_517);
nor U1662 (N_1662,In_54,In_393);
or U1663 (N_1663,In_207,In_767);
and U1664 (N_1664,In_349,In_15);
nand U1665 (N_1665,In_486,In_812);
nand U1666 (N_1666,In_236,In_155);
nand U1667 (N_1667,In_873,In_153);
nor U1668 (N_1668,In_137,In_651);
or U1669 (N_1669,In_496,In_725);
nand U1670 (N_1670,In_22,In_899);
nor U1671 (N_1671,In_83,In_858);
or U1672 (N_1672,In_883,In_800);
or U1673 (N_1673,In_219,In_637);
nor U1674 (N_1674,In_728,In_278);
and U1675 (N_1675,In_74,In_21);
and U1676 (N_1676,In_509,In_655);
and U1677 (N_1677,In_659,In_619);
or U1678 (N_1678,In_18,In_434);
nor U1679 (N_1679,In_806,In_559);
nor U1680 (N_1680,In_258,In_529);
and U1681 (N_1681,In_487,In_376);
nand U1682 (N_1682,In_21,In_512);
xor U1683 (N_1683,In_400,In_608);
nor U1684 (N_1684,In_464,In_486);
and U1685 (N_1685,In_971,In_628);
xnor U1686 (N_1686,In_688,In_530);
or U1687 (N_1687,In_824,In_121);
and U1688 (N_1688,In_503,In_720);
or U1689 (N_1689,In_728,In_117);
and U1690 (N_1690,In_880,In_147);
nor U1691 (N_1691,In_176,In_47);
and U1692 (N_1692,In_815,In_10);
xor U1693 (N_1693,In_580,In_476);
xor U1694 (N_1694,In_849,In_283);
or U1695 (N_1695,In_950,In_580);
nand U1696 (N_1696,In_357,In_948);
nor U1697 (N_1697,In_588,In_722);
xor U1698 (N_1698,In_889,In_823);
and U1699 (N_1699,In_571,In_393);
or U1700 (N_1700,In_154,In_373);
xnor U1701 (N_1701,In_694,In_603);
nand U1702 (N_1702,In_438,In_246);
nor U1703 (N_1703,In_663,In_434);
nand U1704 (N_1704,In_667,In_43);
nor U1705 (N_1705,In_295,In_676);
xor U1706 (N_1706,In_927,In_512);
or U1707 (N_1707,In_987,In_128);
nor U1708 (N_1708,In_897,In_240);
and U1709 (N_1709,In_774,In_451);
and U1710 (N_1710,In_184,In_526);
and U1711 (N_1711,In_846,In_786);
xnor U1712 (N_1712,In_951,In_447);
and U1713 (N_1713,In_766,In_18);
xnor U1714 (N_1714,In_24,In_616);
nor U1715 (N_1715,In_867,In_9);
nand U1716 (N_1716,In_942,In_3);
xor U1717 (N_1717,In_231,In_756);
and U1718 (N_1718,In_322,In_861);
nand U1719 (N_1719,In_629,In_144);
and U1720 (N_1720,In_187,In_337);
nor U1721 (N_1721,In_695,In_530);
and U1722 (N_1722,In_360,In_389);
or U1723 (N_1723,In_238,In_25);
xor U1724 (N_1724,In_91,In_659);
and U1725 (N_1725,In_59,In_245);
and U1726 (N_1726,In_765,In_286);
xor U1727 (N_1727,In_586,In_411);
nor U1728 (N_1728,In_876,In_684);
nor U1729 (N_1729,In_684,In_43);
xor U1730 (N_1730,In_714,In_416);
xnor U1731 (N_1731,In_376,In_591);
nor U1732 (N_1732,In_63,In_288);
nand U1733 (N_1733,In_456,In_690);
or U1734 (N_1734,In_880,In_762);
nand U1735 (N_1735,In_188,In_917);
nor U1736 (N_1736,In_47,In_944);
and U1737 (N_1737,In_126,In_828);
xor U1738 (N_1738,In_995,In_982);
and U1739 (N_1739,In_667,In_147);
or U1740 (N_1740,In_368,In_482);
xnor U1741 (N_1741,In_48,In_968);
xnor U1742 (N_1742,In_434,In_776);
nand U1743 (N_1743,In_276,In_13);
nor U1744 (N_1744,In_500,In_896);
xor U1745 (N_1745,In_173,In_727);
xor U1746 (N_1746,In_651,In_462);
nand U1747 (N_1747,In_670,In_913);
and U1748 (N_1748,In_251,In_855);
nor U1749 (N_1749,In_452,In_172);
or U1750 (N_1750,In_767,In_362);
xnor U1751 (N_1751,In_143,In_565);
and U1752 (N_1752,In_419,In_590);
nand U1753 (N_1753,In_898,In_914);
nand U1754 (N_1754,In_700,In_464);
or U1755 (N_1755,In_848,In_351);
xor U1756 (N_1756,In_753,In_663);
nor U1757 (N_1757,In_554,In_827);
xnor U1758 (N_1758,In_586,In_139);
and U1759 (N_1759,In_328,In_630);
xnor U1760 (N_1760,In_40,In_268);
nor U1761 (N_1761,In_693,In_424);
nand U1762 (N_1762,In_462,In_644);
nor U1763 (N_1763,In_214,In_615);
nand U1764 (N_1764,In_795,In_802);
xor U1765 (N_1765,In_555,In_262);
and U1766 (N_1766,In_540,In_615);
xor U1767 (N_1767,In_29,In_917);
and U1768 (N_1768,In_176,In_105);
nor U1769 (N_1769,In_176,In_502);
nand U1770 (N_1770,In_936,In_733);
or U1771 (N_1771,In_948,In_288);
and U1772 (N_1772,In_654,In_423);
xnor U1773 (N_1773,In_705,In_581);
nand U1774 (N_1774,In_126,In_467);
xnor U1775 (N_1775,In_905,In_337);
nor U1776 (N_1776,In_510,In_689);
and U1777 (N_1777,In_354,In_677);
xnor U1778 (N_1778,In_635,In_926);
and U1779 (N_1779,In_545,In_119);
xnor U1780 (N_1780,In_902,In_350);
nor U1781 (N_1781,In_161,In_682);
nand U1782 (N_1782,In_911,In_367);
or U1783 (N_1783,In_893,In_197);
or U1784 (N_1784,In_281,In_849);
and U1785 (N_1785,In_801,In_223);
or U1786 (N_1786,In_111,In_199);
or U1787 (N_1787,In_999,In_493);
or U1788 (N_1788,In_803,In_887);
nor U1789 (N_1789,In_403,In_46);
or U1790 (N_1790,In_298,In_402);
and U1791 (N_1791,In_308,In_948);
or U1792 (N_1792,In_316,In_243);
nor U1793 (N_1793,In_15,In_970);
or U1794 (N_1794,In_293,In_358);
xor U1795 (N_1795,In_509,In_880);
nand U1796 (N_1796,In_346,In_807);
nor U1797 (N_1797,In_888,In_151);
nor U1798 (N_1798,In_241,In_667);
nor U1799 (N_1799,In_362,In_769);
nor U1800 (N_1800,In_20,In_431);
or U1801 (N_1801,In_0,In_77);
or U1802 (N_1802,In_208,In_634);
nor U1803 (N_1803,In_672,In_292);
nand U1804 (N_1804,In_577,In_441);
or U1805 (N_1805,In_271,In_691);
nand U1806 (N_1806,In_500,In_14);
nor U1807 (N_1807,In_636,In_718);
nand U1808 (N_1808,In_419,In_650);
nand U1809 (N_1809,In_976,In_10);
or U1810 (N_1810,In_526,In_497);
nand U1811 (N_1811,In_366,In_43);
xnor U1812 (N_1812,In_620,In_551);
xor U1813 (N_1813,In_139,In_845);
nand U1814 (N_1814,In_906,In_713);
and U1815 (N_1815,In_118,In_254);
or U1816 (N_1816,In_709,In_493);
or U1817 (N_1817,In_432,In_624);
xor U1818 (N_1818,In_486,In_291);
xor U1819 (N_1819,In_503,In_798);
and U1820 (N_1820,In_53,In_560);
nand U1821 (N_1821,In_907,In_293);
xor U1822 (N_1822,In_798,In_563);
nand U1823 (N_1823,In_161,In_150);
nand U1824 (N_1824,In_56,In_685);
nand U1825 (N_1825,In_286,In_735);
xnor U1826 (N_1826,In_642,In_994);
xor U1827 (N_1827,In_514,In_668);
nand U1828 (N_1828,In_975,In_978);
nor U1829 (N_1829,In_684,In_214);
and U1830 (N_1830,In_914,In_582);
and U1831 (N_1831,In_471,In_451);
nand U1832 (N_1832,In_161,In_605);
xnor U1833 (N_1833,In_838,In_664);
nand U1834 (N_1834,In_251,In_554);
xor U1835 (N_1835,In_722,In_836);
xor U1836 (N_1836,In_210,In_378);
xor U1837 (N_1837,In_669,In_25);
nand U1838 (N_1838,In_695,In_517);
xor U1839 (N_1839,In_770,In_418);
and U1840 (N_1840,In_290,In_509);
xnor U1841 (N_1841,In_857,In_682);
nand U1842 (N_1842,In_114,In_107);
xor U1843 (N_1843,In_171,In_4);
or U1844 (N_1844,In_892,In_96);
xnor U1845 (N_1845,In_681,In_397);
and U1846 (N_1846,In_756,In_768);
xnor U1847 (N_1847,In_663,In_584);
nor U1848 (N_1848,In_957,In_785);
nand U1849 (N_1849,In_415,In_868);
nand U1850 (N_1850,In_193,In_215);
or U1851 (N_1851,In_854,In_350);
nor U1852 (N_1852,In_28,In_820);
nand U1853 (N_1853,In_796,In_26);
or U1854 (N_1854,In_754,In_888);
or U1855 (N_1855,In_20,In_105);
nor U1856 (N_1856,In_133,In_590);
nor U1857 (N_1857,In_448,In_463);
and U1858 (N_1858,In_3,In_934);
nor U1859 (N_1859,In_100,In_984);
or U1860 (N_1860,In_331,In_46);
and U1861 (N_1861,In_846,In_193);
nor U1862 (N_1862,In_969,In_837);
nor U1863 (N_1863,In_459,In_511);
nand U1864 (N_1864,In_439,In_495);
nand U1865 (N_1865,In_961,In_334);
and U1866 (N_1866,In_731,In_738);
or U1867 (N_1867,In_420,In_267);
xor U1868 (N_1868,In_263,In_408);
xor U1869 (N_1869,In_828,In_124);
and U1870 (N_1870,In_824,In_82);
xor U1871 (N_1871,In_937,In_632);
nand U1872 (N_1872,In_571,In_867);
nand U1873 (N_1873,In_861,In_831);
or U1874 (N_1874,In_961,In_448);
nand U1875 (N_1875,In_558,In_515);
or U1876 (N_1876,In_551,In_495);
nor U1877 (N_1877,In_790,In_687);
nand U1878 (N_1878,In_990,In_823);
and U1879 (N_1879,In_268,In_782);
or U1880 (N_1880,In_304,In_560);
and U1881 (N_1881,In_248,In_96);
nor U1882 (N_1882,In_989,In_336);
nor U1883 (N_1883,In_494,In_596);
nor U1884 (N_1884,In_318,In_333);
nand U1885 (N_1885,In_186,In_115);
or U1886 (N_1886,In_519,In_645);
nor U1887 (N_1887,In_65,In_52);
xor U1888 (N_1888,In_727,In_143);
xor U1889 (N_1889,In_937,In_886);
nor U1890 (N_1890,In_224,In_667);
or U1891 (N_1891,In_928,In_169);
nand U1892 (N_1892,In_996,In_980);
and U1893 (N_1893,In_687,In_920);
nor U1894 (N_1894,In_458,In_390);
nand U1895 (N_1895,In_7,In_581);
xor U1896 (N_1896,In_665,In_838);
xnor U1897 (N_1897,In_662,In_425);
xnor U1898 (N_1898,In_854,In_765);
or U1899 (N_1899,In_251,In_847);
or U1900 (N_1900,In_390,In_647);
xnor U1901 (N_1901,In_518,In_252);
and U1902 (N_1902,In_359,In_763);
or U1903 (N_1903,In_878,In_605);
xnor U1904 (N_1904,In_131,In_699);
xnor U1905 (N_1905,In_856,In_708);
xor U1906 (N_1906,In_466,In_756);
xnor U1907 (N_1907,In_609,In_102);
and U1908 (N_1908,In_55,In_219);
and U1909 (N_1909,In_344,In_623);
nor U1910 (N_1910,In_75,In_678);
or U1911 (N_1911,In_831,In_234);
nor U1912 (N_1912,In_330,In_471);
or U1913 (N_1913,In_410,In_827);
and U1914 (N_1914,In_804,In_244);
nand U1915 (N_1915,In_472,In_427);
or U1916 (N_1916,In_262,In_835);
nor U1917 (N_1917,In_722,In_126);
or U1918 (N_1918,In_847,In_690);
nand U1919 (N_1919,In_236,In_931);
nand U1920 (N_1920,In_931,In_816);
nand U1921 (N_1921,In_114,In_865);
xnor U1922 (N_1922,In_576,In_665);
xnor U1923 (N_1923,In_572,In_147);
xor U1924 (N_1924,In_333,In_512);
nor U1925 (N_1925,In_820,In_446);
nor U1926 (N_1926,In_615,In_377);
or U1927 (N_1927,In_130,In_890);
and U1928 (N_1928,In_828,In_640);
xor U1929 (N_1929,In_257,In_610);
nand U1930 (N_1930,In_295,In_396);
nand U1931 (N_1931,In_352,In_840);
nand U1932 (N_1932,In_388,In_814);
or U1933 (N_1933,In_739,In_882);
xnor U1934 (N_1934,In_246,In_457);
and U1935 (N_1935,In_565,In_405);
and U1936 (N_1936,In_399,In_539);
xor U1937 (N_1937,In_991,In_367);
or U1938 (N_1938,In_609,In_507);
xnor U1939 (N_1939,In_220,In_394);
xnor U1940 (N_1940,In_553,In_743);
xnor U1941 (N_1941,In_184,In_937);
xnor U1942 (N_1942,In_913,In_192);
xnor U1943 (N_1943,In_416,In_934);
nor U1944 (N_1944,In_726,In_783);
or U1945 (N_1945,In_707,In_295);
xnor U1946 (N_1946,In_411,In_310);
xor U1947 (N_1947,In_328,In_285);
or U1948 (N_1948,In_521,In_493);
or U1949 (N_1949,In_722,In_94);
nor U1950 (N_1950,In_945,In_220);
nand U1951 (N_1951,In_208,In_873);
nand U1952 (N_1952,In_812,In_96);
and U1953 (N_1953,In_80,In_566);
nand U1954 (N_1954,In_865,In_11);
or U1955 (N_1955,In_41,In_646);
xnor U1956 (N_1956,In_573,In_531);
nand U1957 (N_1957,In_340,In_262);
and U1958 (N_1958,In_42,In_694);
nor U1959 (N_1959,In_561,In_713);
xnor U1960 (N_1960,In_608,In_417);
nand U1961 (N_1961,In_461,In_11);
nor U1962 (N_1962,In_245,In_703);
or U1963 (N_1963,In_967,In_545);
or U1964 (N_1964,In_597,In_748);
and U1965 (N_1965,In_235,In_716);
or U1966 (N_1966,In_70,In_976);
and U1967 (N_1967,In_696,In_291);
or U1968 (N_1968,In_35,In_54);
and U1969 (N_1969,In_172,In_402);
nor U1970 (N_1970,In_283,In_48);
and U1971 (N_1971,In_961,In_884);
and U1972 (N_1972,In_928,In_35);
nor U1973 (N_1973,In_284,In_904);
nor U1974 (N_1974,In_140,In_686);
xnor U1975 (N_1975,In_715,In_243);
nor U1976 (N_1976,In_90,In_781);
nand U1977 (N_1977,In_821,In_537);
xnor U1978 (N_1978,In_11,In_568);
nor U1979 (N_1979,In_240,In_654);
or U1980 (N_1980,In_138,In_308);
and U1981 (N_1981,In_536,In_591);
nor U1982 (N_1982,In_81,In_98);
and U1983 (N_1983,In_278,In_356);
or U1984 (N_1984,In_847,In_235);
xor U1985 (N_1985,In_755,In_109);
xnor U1986 (N_1986,In_767,In_804);
and U1987 (N_1987,In_49,In_455);
or U1988 (N_1988,In_66,In_727);
or U1989 (N_1989,In_574,In_148);
nor U1990 (N_1990,In_42,In_678);
xnor U1991 (N_1991,In_163,In_572);
and U1992 (N_1992,In_87,In_842);
nor U1993 (N_1993,In_12,In_808);
and U1994 (N_1994,In_586,In_456);
xor U1995 (N_1995,In_491,In_78);
or U1996 (N_1996,In_607,In_779);
nor U1997 (N_1997,In_718,In_333);
nor U1998 (N_1998,In_906,In_920);
nor U1999 (N_1999,In_34,In_501);
and U2000 (N_2000,N_1557,N_1224);
nor U2001 (N_2001,N_1638,N_112);
nor U2002 (N_2002,N_1682,N_79);
nor U2003 (N_2003,N_242,N_1772);
nand U2004 (N_2004,N_585,N_1900);
or U2005 (N_2005,N_1724,N_1037);
xor U2006 (N_2006,N_455,N_1694);
nor U2007 (N_2007,N_1028,N_301);
nor U2008 (N_2008,N_215,N_724);
nor U2009 (N_2009,N_879,N_1891);
nor U2010 (N_2010,N_219,N_509);
nor U2011 (N_2011,N_1793,N_760);
xor U2012 (N_2012,N_306,N_676);
nand U2013 (N_2013,N_1725,N_1381);
xor U2014 (N_2014,N_627,N_479);
or U2015 (N_2015,N_273,N_1915);
or U2016 (N_2016,N_717,N_1610);
xnor U2017 (N_2017,N_1080,N_593);
xnor U2018 (N_2018,N_1306,N_737);
nor U2019 (N_2019,N_145,N_1388);
nand U2020 (N_2020,N_1147,N_1288);
nor U2021 (N_2021,N_116,N_1957);
nand U2022 (N_2022,N_17,N_1951);
xor U2023 (N_2023,N_784,N_200);
nor U2024 (N_2024,N_608,N_1966);
nand U2025 (N_2025,N_1971,N_1829);
nand U2026 (N_2026,N_247,N_1251);
or U2027 (N_2027,N_1707,N_682);
and U2028 (N_2028,N_844,N_1267);
xnor U2029 (N_2029,N_1249,N_349);
and U2030 (N_2030,N_113,N_1089);
and U2031 (N_2031,N_117,N_594);
nor U2032 (N_2032,N_141,N_334);
or U2033 (N_2033,N_8,N_262);
or U2034 (N_2034,N_119,N_933);
or U2035 (N_2035,N_581,N_507);
and U2036 (N_2036,N_1454,N_625);
nor U2037 (N_2037,N_487,N_263);
xnor U2038 (N_2038,N_723,N_1507);
nand U2039 (N_2039,N_123,N_900);
nor U2040 (N_2040,N_605,N_577);
and U2041 (N_2041,N_1247,N_1452);
or U2042 (N_2042,N_1355,N_87);
or U2043 (N_2043,N_224,N_328);
and U2044 (N_2044,N_1887,N_1161);
xnor U2045 (N_2045,N_1601,N_427);
nand U2046 (N_2046,N_418,N_482);
nor U2047 (N_2047,N_1589,N_1988);
nand U2048 (N_2048,N_1778,N_408);
nor U2049 (N_2049,N_1660,N_503);
xor U2050 (N_2050,N_1121,N_718);
nand U2051 (N_2051,N_1976,N_586);
nor U2052 (N_2052,N_189,N_1349);
xnor U2053 (N_2053,N_1266,N_1359);
and U2054 (N_2054,N_1204,N_284);
and U2055 (N_2055,N_1406,N_788);
nand U2056 (N_2056,N_310,N_1624);
or U2057 (N_2057,N_1869,N_1759);
nor U2058 (N_2058,N_557,N_1628);
nand U2059 (N_2059,N_777,N_1006);
or U2060 (N_2060,N_130,N_144);
xor U2061 (N_2061,N_673,N_1415);
or U2062 (N_2062,N_1835,N_97);
xor U2063 (N_2063,N_965,N_587);
xor U2064 (N_2064,N_748,N_1180);
or U2065 (N_2065,N_960,N_822);
nand U2066 (N_2066,N_1491,N_1334);
nand U2067 (N_2067,N_1100,N_190);
and U2068 (N_2068,N_1408,N_388);
xor U2069 (N_2069,N_1310,N_160);
or U2070 (N_2070,N_1220,N_640);
and U2071 (N_2071,N_1853,N_369);
or U2072 (N_2072,N_1146,N_149);
and U2073 (N_2073,N_1409,N_1139);
or U2074 (N_2074,N_83,N_691);
nand U2075 (N_2075,N_966,N_1559);
and U2076 (N_2076,N_1997,N_1656);
and U2077 (N_2077,N_1486,N_878);
and U2078 (N_2078,N_483,N_456);
and U2079 (N_2079,N_1546,N_931);
and U2080 (N_2080,N_704,N_1014);
nor U2081 (N_2081,N_1088,N_647);
nor U2082 (N_2082,N_1038,N_196);
xnor U2083 (N_2083,N_322,N_244);
nand U2084 (N_2084,N_1307,N_122);
and U2085 (N_2085,N_228,N_710);
nand U2086 (N_2086,N_610,N_615);
and U2087 (N_2087,N_1313,N_1308);
xnor U2088 (N_2088,N_1558,N_1376);
nand U2089 (N_2089,N_340,N_1646);
and U2090 (N_2090,N_1169,N_1556);
nor U2091 (N_2091,N_287,N_77);
nor U2092 (N_2092,N_1234,N_513);
nand U2093 (N_2093,N_600,N_1154);
nor U2094 (N_2094,N_510,N_296);
nor U2095 (N_2095,N_982,N_887);
xnor U2096 (N_2096,N_1398,N_693);
xor U2097 (N_2097,N_424,N_72);
nand U2098 (N_2098,N_414,N_1873);
or U2099 (N_2099,N_2,N_103);
xnor U2100 (N_2100,N_411,N_516);
xor U2101 (N_2101,N_431,N_1010);
or U2102 (N_2102,N_99,N_1843);
or U2103 (N_2103,N_1492,N_1751);
nand U2104 (N_2104,N_667,N_1296);
xor U2105 (N_2105,N_1049,N_1289);
nor U2106 (N_2106,N_1199,N_352);
or U2107 (N_2107,N_152,N_1292);
nand U2108 (N_2108,N_1612,N_311);
xnor U2109 (N_2109,N_867,N_641);
and U2110 (N_2110,N_781,N_1893);
nand U2111 (N_2111,N_1807,N_279);
and U2112 (N_2112,N_203,N_675);
nor U2113 (N_2113,N_1851,N_642);
or U2114 (N_2114,N_683,N_810);
xor U2115 (N_2115,N_70,N_1105);
nor U2116 (N_2116,N_801,N_1324);
xor U2117 (N_2117,N_134,N_670);
nand U2118 (N_2118,N_1577,N_1475);
nand U2119 (N_2119,N_156,N_1283);
xor U2120 (N_2120,N_106,N_1757);
nand U2121 (N_2121,N_1762,N_1440);
and U2122 (N_2122,N_237,N_750);
or U2123 (N_2123,N_502,N_1422);
xor U2124 (N_2124,N_841,N_1305);
and U2125 (N_2125,N_1539,N_857);
xor U2126 (N_2126,N_1630,N_297);
or U2127 (N_2127,N_623,N_29);
or U2128 (N_2128,N_533,N_899);
nand U2129 (N_2129,N_257,N_406);
nand U2130 (N_2130,N_1791,N_715);
nor U2131 (N_2131,N_1705,N_1077);
xnor U2132 (N_2132,N_1270,N_47);
nor U2133 (N_2133,N_1389,N_901);
xnor U2134 (N_2134,N_162,N_3);
nand U2135 (N_2135,N_882,N_959);
or U2136 (N_2136,N_1438,N_1788);
nand U2137 (N_2137,N_1,N_1547);
nor U2138 (N_2138,N_1836,N_873);
xnor U2139 (N_2139,N_752,N_800);
xor U2140 (N_2140,N_1832,N_762);
nand U2141 (N_2141,N_726,N_1644);
nor U2142 (N_2142,N_1719,N_823);
xor U2143 (N_2143,N_1698,N_1984);
and U2144 (N_2144,N_656,N_1321);
nor U2145 (N_2145,N_536,N_293);
xor U2146 (N_2146,N_1593,N_1095);
or U2147 (N_2147,N_778,N_572);
nor U2148 (N_2148,N_942,N_1463);
nor U2149 (N_2149,N_1050,N_551);
nor U2150 (N_2150,N_570,N_923);
or U2151 (N_2151,N_1250,N_1140);
or U2152 (N_2152,N_816,N_1684);
nor U2153 (N_2153,N_1320,N_1116);
or U2154 (N_2154,N_1258,N_926);
or U2155 (N_2155,N_735,N_688);
xnor U2156 (N_2156,N_542,N_288);
or U2157 (N_2157,N_1091,N_568);
or U2158 (N_2158,N_1239,N_904);
nor U2159 (N_2159,N_1040,N_1280);
nand U2160 (N_2160,N_884,N_1527);
or U2161 (N_2161,N_23,N_269);
or U2162 (N_2162,N_839,N_1399);
and U2163 (N_2163,N_1735,N_938);
xor U2164 (N_2164,N_876,N_1530);
or U2165 (N_2165,N_1651,N_378);
nand U2166 (N_2166,N_654,N_1622);
or U2167 (N_2167,N_1513,N_1036);
nand U2168 (N_2168,N_1924,N_681);
and U2169 (N_2169,N_1943,N_558);
or U2170 (N_2170,N_360,N_1072);
xnor U2171 (N_2171,N_11,N_469);
nor U2172 (N_2172,N_606,N_265);
or U2173 (N_2173,N_383,N_1695);
and U2174 (N_2174,N_1773,N_208);
nand U2175 (N_2175,N_1803,N_1103);
and U2176 (N_2176,N_1822,N_1002);
nor U2177 (N_2177,N_906,N_1564);
and U2178 (N_2178,N_394,N_961);
nand U2179 (N_2179,N_1143,N_711);
nor U2180 (N_2180,N_1493,N_1537);
nand U2181 (N_2181,N_1022,N_973);
nor U2182 (N_2182,N_381,N_1738);
xor U2183 (N_2183,N_1828,N_853);
xor U2184 (N_2184,N_1183,N_1244);
xor U2185 (N_2185,N_1108,N_604);
nor U2186 (N_2186,N_253,N_1590);
or U2187 (N_2187,N_1850,N_184);
or U2188 (N_2188,N_912,N_815);
or U2189 (N_2189,N_1386,N_1153);
and U2190 (N_2190,N_1083,N_1930);
xor U2191 (N_2191,N_1882,N_1472);
xor U2192 (N_2192,N_776,N_1366);
xor U2193 (N_2193,N_1343,N_147);
and U2194 (N_2194,N_1114,N_1134);
xor U2195 (N_2195,N_1563,N_695);
and U2196 (N_2196,N_1008,N_1649);
nor U2197 (N_2197,N_150,N_1098);
and U2198 (N_2198,N_1716,N_1060);
xnor U2199 (N_2199,N_1240,N_372);
nor U2200 (N_2200,N_477,N_1057);
nor U2201 (N_2201,N_896,N_1074);
nor U2202 (N_2202,N_1519,N_798);
xnor U2203 (N_2203,N_261,N_744);
xnor U2204 (N_2204,N_775,N_1795);
nor U2205 (N_2205,N_1506,N_539);
and U2206 (N_2206,N_802,N_1046);
and U2207 (N_2207,N_1858,N_575);
and U2208 (N_2208,N_1992,N_1554);
nand U2209 (N_2209,N_1065,N_1727);
and U2210 (N_2210,N_1344,N_1595);
xnor U2211 (N_2211,N_108,N_1841);
nor U2212 (N_2212,N_211,N_1647);
xor U2213 (N_2213,N_1721,N_1462);
xor U2214 (N_2214,N_927,N_580);
nor U2215 (N_2215,N_1973,N_1362);
and U2216 (N_2216,N_1207,N_1482);
xor U2217 (N_2217,N_1261,N_1185);
nand U2218 (N_2218,N_246,N_1588);
xor U2219 (N_2219,N_1063,N_1871);
and U2220 (N_2220,N_639,N_964);
xnor U2221 (N_2221,N_1503,N_620);
nand U2222 (N_2222,N_866,N_36);
nor U2223 (N_2223,N_1808,N_826);
and U2224 (N_2224,N_1238,N_94);
and U2225 (N_2225,N_102,N_1094);
nand U2226 (N_2226,N_733,N_561);
nor U2227 (N_2227,N_170,N_1713);
nand U2228 (N_2228,N_741,N_588);
nand U2229 (N_2229,N_1200,N_451);
and U2230 (N_2230,N_62,N_1823);
xor U2231 (N_2231,N_146,N_535);
and U2232 (N_2232,N_463,N_1096);
nor U2233 (N_2233,N_1416,N_720);
nand U2234 (N_2234,N_1410,N_183);
nor U2235 (N_2235,N_63,N_1332);
nand U2236 (N_2236,N_836,N_974);
nor U2237 (N_2237,N_1230,N_1173);
or U2238 (N_2238,N_793,N_1403);
nand U2239 (N_2239,N_1627,N_1617);
and U2240 (N_2240,N_435,N_1412);
and U2241 (N_2241,N_1863,N_848);
xnor U2242 (N_2242,N_674,N_1780);
xor U2243 (N_2243,N_1710,N_234);
nand U2244 (N_2244,N_1205,N_924);
and U2245 (N_2245,N_12,N_703);
or U2246 (N_2246,N_598,N_562);
xnor U2247 (N_2247,N_484,N_114);
and U2248 (N_2248,N_1168,N_1796);
nor U2249 (N_2249,N_366,N_191);
and U2250 (N_2250,N_1771,N_413);
or U2251 (N_2251,N_1608,N_607);
nor U2252 (N_2252,N_1110,N_543);
xnor U2253 (N_2253,N_1777,N_163);
and U2254 (N_2254,N_1404,N_1905);
nand U2255 (N_2255,N_528,N_1112);
and U2256 (N_2256,N_1192,N_1030);
and U2257 (N_2257,N_612,N_467);
nor U2258 (N_2258,N_1004,N_172);
and U2259 (N_2259,N_902,N_277);
nand U2260 (N_2260,N_345,N_1550);
nand U2261 (N_2261,N_1208,N_1446);
and U2262 (N_2262,N_9,N_1193);
nor U2263 (N_2263,N_852,N_1394);
nand U2264 (N_2264,N_1113,N_127);
nor U2265 (N_2265,N_1831,N_721);
or U2266 (N_2266,N_1418,N_1342);
or U2267 (N_2267,N_1323,N_1980);
and U2268 (N_2268,N_429,N_1212);
nand U2269 (N_2269,N_1825,N_259);
and U2270 (N_2270,N_664,N_506);
nor U2271 (N_2271,N_18,N_359);
or U2272 (N_2272,N_1625,N_1675);
nand U2273 (N_2273,N_1687,N_1963);
or U2274 (N_2274,N_1717,N_35);
xor U2275 (N_2275,N_448,N_1352);
and U2276 (N_2276,N_24,N_1782);
and U2277 (N_2277,N_473,N_390);
or U2278 (N_2278,N_1696,N_313);
and U2279 (N_2279,N_1340,N_375);
nor U2280 (N_2280,N_619,N_1521);
and U2281 (N_2281,N_85,N_790);
nand U2282 (N_2282,N_1549,N_1948);
and U2283 (N_2283,N_1137,N_417);
nand U2284 (N_2284,N_419,N_1718);
and U2285 (N_2285,N_895,N_1448);
or U2286 (N_2286,N_1812,N_1935);
nor U2287 (N_2287,N_1445,N_751);
nand U2288 (N_2288,N_1487,N_660);
nand U2289 (N_2289,N_1297,N_550);
nor U2290 (N_2290,N_1552,N_1026);
and U2291 (N_2291,N_314,N_139);
and U2292 (N_2292,N_474,N_1723);
xor U2293 (N_2293,N_519,N_338);
nor U2294 (N_2294,N_986,N_1701);
xnor U2295 (N_2295,N_104,N_1286);
xor U2296 (N_2296,N_115,N_480);
and U2297 (N_2297,N_1035,N_412);
or U2298 (N_2298,N_1439,N_1369);
or U2299 (N_2299,N_1998,N_553);
or U2300 (N_2300,N_1879,N_1889);
nor U2301 (N_2301,N_532,N_874);
and U2302 (N_2302,N_565,N_166);
and U2303 (N_2303,N_1155,N_967);
xor U2304 (N_2304,N_441,N_1184);
nor U2305 (N_2305,N_1740,N_1222);
xor U2306 (N_2306,N_227,N_754);
or U2307 (N_2307,N_1954,N_779);
xnor U2308 (N_2308,N_1587,N_426);
nand U2309 (N_2309,N_1163,N_285);
or U2310 (N_2310,N_1986,N_552);
nand U2311 (N_2311,N_643,N_522);
nand U2312 (N_2312,N_1485,N_730);
and U2313 (N_2313,N_814,N_1387);
or U2314 (N_2314,N_168,N_1523);
and U2315 (N_2315,N_1714,N_1581);
xor U2316 (N_2316,N_1372,N_651);
nor U2317 (N_2317,N_1385,N_1319);
xor U2318 (N_2318,N_124,N_1594);
xnor U2319 (N_2319,N_493,N_450);
nand U2320 (N_2320,N_997,N_105);
or U2321 (N_2321,N_290,N_1195);
nor U2322 (N_2322,N_1479,N_364);
and U2323 (N_2323,N_327,N_1237);
nand U2324 (N_2324,N_1805,N_555);
nand U2325 (N_2325,N_517,N_1532);
or U2326 (N_2326,N_1819,N_492);
or U2327 (N_2327,N_201,N_1081);
nand U2328 (N_2328,N_302,N_919);
and U2329 (N_2329,N_1309,N_1177);
and U2330 (N_2330,N_1464,N_278);
or U2331 (N_2331,N_729,N_1068);
or U2332 (N_2332,N_834,N_131);
or U2333 (N_2333,N_993,N_1353);
or U2334 (N_2334,N_109,N_1000);
xor U2335 (N_2335,N_1602,N_1728);
xor U2336 (N_2336,N_174,N_365);
nor U2337 (N_2337,N_1923,N_1910);
or U2338 (N_2338,N_1364,N_885);
nand U2339 (N_2339,N_1544,N_1637);
nand U2340 (N_2340,N_1400,N_348);
nor U2341 (N_2341,N_52,N_763);
or U2342 (N_2342,N_1395,N_100);
and U2343 (N_2343,N_657,N_849);
and U2344 (N_2344,N_1102,N_1356);
and U2345 (N_2345,N_1371,N_1241);
xor U2346 (N_2346,N_169,N_21);
nand U2347 (N_2347,N_1509,N_1766);
nor U2348 (N_2348,N_1806,N_1062);
nand U2349 (N_2349,N_1969,N_1736);
or U2350 (N_2350,N_1459,N_1281);
nor U2351 (N_2351,N_541,N_1571);
nand U2352 (N_2352,N_566,N_1929);
xnor U2353 (N_2353,N_403,N_1578);
or U2354 (N_2354,N_1045,N_745);
or U2355 (N_2355,N_446,N_1654);
xnor U2356 (N_2356,N_1449,N_333);
nand U2357 (N_2357,N_795,N_351);
or U2358 (N_2358,N_1614,N_303);
nand U2359 (N_2359,N_1333,N_1397);
and U2360 (N_2360,N_1926,N_1164);
nor U2361 (N_2361,N_1073,N_819);
and U2362 (N_2362,N_1011,N_1326);
and U2363 (N_2363,N_233,N_792);
and U2364 (N_2364,N_1517,N_680);
nor U2365 (N_2365,N_478,N_1754);
or U2366 (N_2366,N_1162,N_315);
xor U2367 (N_2367,N_205,N_860);
and U2368 (N_2368,N_405,N_61);
and U2369 (N_2369,N_292,N_787);
or U2370 (N_2370,N_336,N_1059);
xnor U2371 (N_2371,N_363,N_350);
and U2372 (N_2372,N_1260,N_121);
or U2373 (N_2373,N_1775,N_192);
xor U2374 (N_2374,N_1708,N_68);
nor U2375 (N_2375,N_1661,N_1864);
or U2376 (N_2376,N_387,N_1756);
and U2377 (N_2377,N_1936,N_355);
nand U2378 (N_2378,N_1681,N_433);
nor U2379 (N_2379,N_829,N_1555);
xor U2380 (N_2380,N_1282,N_5);
nand U2381 (N_2381,N_71,N_892);
nor U2382 (N_2382,N_84,N_1975);
or U2383 (N_2383,N_941,N_571);
nand U2384 (N_2384,N_1335,N_1460);
or U2385 (N_2385,N_438,N_952);
xor U2386 (N_2386,N_661,N_574);
and U2387 (N_2387,N_548,N_1079);
xor U2388 (N_2388,N_1693,N_1840);
nor U2389 (N_2389,N_700,N_110);
and U2390 (N_2390,N_264,N_1568);
nor U2391 (N_2391,N_1149,N_1592);
and U2392 (N_2392,N_443,N_225);
xor U2393 (N_2393,N_231,N_78);
nand U2394 (N_2394,N_797,N_195);
and U2395 (N_2395,N_1671,N_1938);
nand U2396 (N_2396,N_1987,N_13);
xnor U2397 (N_2397,N_384,N_44);
or U2398 (N_2398,N_389,N_218);
nor U2399 (N_2399,N_1417,N_136);
or U2400 (N_2400,N_1393,N_1316);
or U2401 (N_2401,N_569,N_1833);
nor U2402 (N_2402,N_1743,N_1846);
xnor U2403 (N_2403,N_436,N_1774);
xnor U2404 (N_2404,N_1023,N_1051);
or U2405 (N_2405,N_1582,N_1514);
xor U2406 (N_2406,N_258,N_687);
xor U2407 (N_2407,N_1277,N_1361);
nand U2408 (N_2408,N_236,N_1314);
xnor U2409 (N_2409,N_1243,N_1859);
xnor U2410 (N_2410,N_1787,N_1918);
xor U2411 (N_2411,N_101,N_1123);
nor U2412 (N_2412,N_805,N_1672);
xnor U2413 (N_2413,N_240,N_179);
nor U2414 (N_2414,N_1090,N_1890);
nand U2415 (N_2415,N_1540,N_1330);
or U2416 (N_2416,N_1156,N_56);
nand U2417 (N_2417,N_1674,N_1597);
or U2418 (N_2418,N_341,N_804);
and U2419 (N_2419,N_45,N_1176);
xor U2420 (N_2420,N_1685,N_402);
nand U2421 (N_2421,N_1515,N_1295);
nor U2422 (N_2422,N_1606,N_1444);
xnor U2423 (N_2423,N_850,N_1107);
or U2424 (N_2424,N_1378,N_530);
xor U2425 (N_2425,N_267,N_377);
nor U2426 (N_2426,N_1958,N_701);
nand U2427 (N_2427,N_1522,N_308);
nand U2428 (N_2428,N_1826,N_582);
nor U2429 (N_2429,N_1436,N_511);
nor U2430 (N_2430,N_1977,N_624);
nor U2431 (N_2431,N_1553,N_573);
nand U2432 (N_2432,N_996,N_1979);
nor U2433 (N_2433,N_252,N_346);
nor U2434 (N_2434,N_1086,N_789);
nor U2435 (N_2435,N_422,N_1560);
nand U2436 (N_2436,N_1383,N_1003);
and U2437 (N_2437,N_512,N_1465);
nand U2438 (N_2438,N_1603,N_880);
xor U2439 (N_2439,N_159,N_1894);
or U2440 (N_2440,N_368,N_132);
or U2441 (N_2441,N_157,N_1396);
xnor U2442 (N_2442,N_1466,N_1262);
xor U2443 (N_2443,N_1175,N_992);
or U2444 (N_2444,N_1734,N_1955);
nand U2445 (N_2445,N_663,N_957);
nand U2446 (N_2446,N_209,N_1903);
and U2447 (N_2447,N_1076,N_698);
xnor U2448 (N_2448,N_1048,N_1039);
nand U2449 (N_2449,N_1377,N_716);
and U2450 (N_2450,N_1531,N_975);
xnor U2451 (N_2451,N_524,N_1133);
xnor U2452 (N_2452,N_1217,N_1329);
nor U2453 (N_2453,N_1962,N_1689);
or U2454 (N_2454,N_692,N_1233);
nand U2455 (N_2455,N_1178,N_1151);
nand U2456 (N_2456,N_1663,N_1502);
xor U2457 (N_2457,N_1567,N_1252);
xnor U2458 (N_2458,N_1433,N_1336);
or U2459 (N_2459,N_515,N_1817);
and U2460 (N_2460,N_500,N_374);
xor U2461 (N_2461,N_1730,N_983);
and U2462 (N_2462,N_1348,N_538);
nor U2463 (N_2463,N_1995,N_28);
or U2464 (N_2464,N_499,N_821);
nor U2465 (N_2465,N_770,N_320);
xor U2466 (N_2466,N_415,N_537);
nor U2467 (N_2467,N_1937,N_19);
nor U2468 (N_2468,N_222,N_1024);
xor U2469 (N_2469,N_1054,N_330);
xor U2470 (N_2470,N_1990,N_1370);
or U2471 (N_2471,N_1119,N_1981);
xor U2472 (N_2472,N_1883,N_270);
xor U2473 (N_2473,N_1457,N_229);
xor U2474 (N_2474,N_1007,N_916);
and U2475 (N_2475,N_198,N_713);
nand U2476 (N_2476,N_1639,N_1363);
xnor U2477 (N_2477,N_1274,N_1005);
or U2478 (N_2478,N_397,N_1215);
and U2479 (N_2479,N_60,N_1665);
and U2480 (N_2480,N_846,N_1902);
and U2481 (N_2481,N_544,N_1913);
and U2482 (N_2482,N_707,N_1842);
nor U2483 (N_2483,N_917,N_92);
nor U2484 (N_2484,N_361,N_1055);
xor U2485 (N_2485,N_1033,N_1202);
nor U2486 (N_2486,N_1201,N_93);
nor U2487 (N_2487,N_1970,N_1471);
and U2488 (N_2488,N_595,N_1426);
nand U2489 (N_2489,N_324,N_120);
xnor U2490 (N_2490,N_1927,N_221);
and U2491 (N_2491,N_148,N_38);
xnor U2492 (N_2492,N_618,N_1392);
nand U2493 (N_2493,N_1510,N_171);
and U2494 (N_2494,N_1520,N_175);
nor U2495 (N_2495,N_1345,N_1844);
or U2496 (N_2496,N_1518,N_1700);
or U2497 (N_2497,N_1679,N_783);
xnor U2498 (N_2498,N_1253,N_937);
and U2499 (N_2499,N_317,N_658);
and U2500 (N_2500,N_809,N_1613);
nand U2501 (N_2501,N_165,N_653);
or U2502 (N_2502,N_972,N_1985);
xor U2503 (N_2503,N_1761,N_1809);
nor U2504 (N_2504,N_953,N_1901);
xor U2505 (N_2505,N_31,N_447);
or U2506 (N_2506,N_1401,N_1269);
or U2507 (N_2507,N_903,N_1331);
xor U2508 (N_2508,N_89,N_423);
nor U2509 (N_2509,N_865,N_1586);
and U2510 (N_2510,N_1830,N_339);
or U2511 (N_2511,N_602,N_1120);
or U2512 (N_2512,N_1061,N_905);
or U2513 (N_2513,N_1750,N_1141);
and U2514 (N_2514,N_1814,N_886);
xnor U2515 (N_2515,N_1203,N_1034);
or U2516 (N_2516,N_817,N_1816);
or U2517 (N_2517,N_485,N_765);
nand U2518 (N_2518,N_694,N_407);
nor U2519 (N_2519,N_603,N_847);
and U2520 (N_2520,N_1414,N_875);
nand U2521 (N_2521,N_1504,N_799);
and U2522 (N_2522,N_495,N_46);
nor U2523 (N_2523,N_1758,N_1657);
or U2524 (N_2524,N_1275,N_1895);
or U2525 (N_2525,N_769,N_75);
xor U2526 (N_2526,N_980,N_434);
or U2527 (N_2527,N_981,N_154);
nor U2528 (N_2528,N_1868,N_1596);
and U2529 (N_2529,N_1468,N_894);
nor U2530 (N_2530,N_1848,N_371);
or U2531 (N_2531,N_1167,N_476);
nand U2532 (N_2532,N_749,N_1481);
or U2533 (N_2533,N_457,N_1019);
nor U2534 (N_2534,N_742,N_1755);
nand U2535 (N_2535,N_1018,N_1256);
xor U2536 (N_2536,N_15,N_1093);
xor U2537 (N_2537,N_1747,N_1453);
nand U2538 (N_2538,N_1699,N_1294);
or U2539 (N_2539,N_1744,N_1499);
xnor U2540 (N_2540,N_1742,N_950);
or U2541 (N_2541,N_343,N_1232);
or U2542 (N_2542,N_1078,N_630);
and U2543 (N_2543,N_1402,N_858);
nor U2544 (N_2544,N_416,N_1856);
nor U2545 (N_2545,N_243,N_1538);
nand U2546 (N_2546,N_995,N_1786);
nand U2547 (N_2547,N_1609,N_877);
nor U2548 (N_2548,N_404,N_979);
nand U2549 (N_2549,N_1029,N_1179);
nor U2550 (N_2550,N_1291,N_1631);
nor U2551 (N_2551,N_260,N_1317);
and U2552 (N_2552,N_945,N_216);
nand U2553 (N_2553,N_794,N_1769);
nand U2554 (N_2554,N_1748,N_768);
xnor U2555 (N_2555,N_1692,N_684);
or U2556 (N_2556,N_1712,N_655);
and U2557 (N_2557,N_890,N_1318);
xor U2558 (N_2558,N_1337,N_1218);
nand U2559 (N_2559,N_1476,N_1271);
nand U2560 (N_2560,N_453,N_1870);
nand U2561 (N_2561,N_1585,N_910);
and U2562 (N_2562,N_353,N_820);
and U2563 (N_2563,N_1405,N_1824);
xor U2564 (N_2564,N_420,N_547);
xnor U2565 (N_2565,N_988,N_250);
and U2566 (N_2566,N_1432,N_758);
nand U2567 (N_2567,N_4,N_1373);
nor U2568 (N_2568,N_1382,N_940);
and U2569 (N_2569,N_1874,N_727);
xnor U2570 (N_2570,N_276,N_1273);
or U2571 (N_2571,N_576,N_140);
nand U2572 (N_2572,N_842,N_1961);
and U2573 (N_2573,N_1741,N_1122);
nor U2574 (N_2574,N_501,N_1983);
and U2575 (N_2575,N_1875,N_1784);
and U2576 (N_2576,N_34,N_1996);
or U2577 (N_2577,N_1508,N_197);
nand U2578 (N_2578,N_559,N_915);
and U2579 (N_2579,N_1354,N_67);
or U2580 (N_2580,N_678,N_1315);
or U2581 (N_2581,N_468,N_629);
and U2582 (N_2582,N_1191,N_459);
and U2583 (N_2583,N_958,N_1231);
and U2584 (N_2584,N_1745,N_771);
xnor U2585 (N_2585,N_425,N_1726);
or U2586 (N_2586,N_212,N_1174);
or U2587 (N_2587,N_773,N_1670);
and U2588 (N_2588,N_767,N_791);
or U2589 (N_2589,N_321,N_118);
and U2590 (N_2590,N_738,N_1683);
nand U2591 (N_2591,N_689,N_1953);
nand U2592 (N_2592,N_199,N_1126);
or U2593 (N_2593,N_531,N_828);
nor U2594 (N_2594,N_268,N_948);
and U2595 (N_2595,N_1346,N_883);
and U2596 (N_2596,N_1770,N_632);
or U2597 (N_2597,N_739,N_1876);
and U2598 (N_2598,N_617,N_1419);
xor U2599 (N_2599,N_1619,N_428);
nor U2600 (N_2600,N_440,N_757);
nand U2601 (N_2601,N_1171,N_1431);
or U2602 (N_2602,N_1912,N_1645);
nor U2603 (N_2603,N_1495,N_1196);
or U2604 (N_2604,N_888,N_1922);
or U2605 (N_2605,N_1666,N_1720);
xor U2606 (N_2606,N_1680,N_1686);
nor U2607 (N_2607,N_245,N_863);
nand U2608 (N_2608,N_1952,N_217);
or U2609 (N_2609,N_1576,N_1157);
nand U2610 (N_2610,N_1272,N_299);
and U2611 (N_2611,N_272,N_399);
nor U2612 (N_2612,N_1264,N_1043);
nor U2613 (N_2613,N_864,N_1959);
nor U2614 (N_2614,N_845,N_280);
or U2615 (N_2615,N_1357,N_833);
or U2616 (N_2616,N_1673,N_1633);
xor U2617 (N_2617,N_143,N_1827);
xnor U2618 (N_2618,N_1082,N_1991);
nand U2619 (N_2619,N_1925,N_914);
or U2620 (N_2620,N_999,N_786);
xnor U2621 (N_2621,N_1702,N_1434);
nand U2622 (N_2622,N_1430,N_1839);
and U2623 (N_2623,N_944,N_990);
or U2624 (N_2624,N_318,N_266);
nand U2625 (N_2625,N_392,N_1934);
and U2626 (N_2626,N_989,N_870);
nor U2627 (N_2627,N_907,N_1265);
xor U2628 (N_2628,N_1573,N_1852);
nand U2629 (N_2629,N_991,N_1776);
xor U2630 (N_2630,N_1993,N_1731);
and U2631 (N_2631,N_490,N_1792);
nor U2632 (N_2632,N_458,N_1384);
xnor U2633 (N_2633,N_1669,N_1904);
or U2634 (N_2634,N_719,N_57);
and U2635 (N_2635,N_1128,N_697);
and U2636 (N_2636,N_871,N_32);
and U2637 (N_2637,N_838,N_616);
nor U2638 (N_2638,N_400,N_951);
nor U2639 (N_2639,N_1569,N_64);
or U2640 (N_2640,N_30,N_669);
nand U2641 (N_2641,N_1437,N_69);
nor U2642 (N_2642,N_592,N_319);
nor U2643 (N_2643,N_725,N_1303);
or U2644 (N_2644,N_668,N_488);
or U2645 (N_2645,N_1411,N_129);
or U2646 (N_2646,N_1621,N_645);
and U2647 (N_2647,N_20,N_897);
xnor U2648 (N_2648,N_1798,N_452);
or U2649 (N_2649,N_1562,N_597);
or U2650 (N_2650,N_949,N_921);
and U2651 (N_2651,N_782,N_1311);
or U2652 (N_2652,N_1494,N_1668);
xor U2653 (N_2653,N_1284,N_382);
xor U2654 (N_2654,N_1643,N_50);
xor U2655 (N_2655,N_48,N_59);
and U2656 (N_2656,N_180,N_1015);
or U2657 (N_2657,N_1551,N_185);
nand U2658 (N_2658,N_549,N_679);
xnor U2659 (N_2659,N_1498,N_635);
or U2660 (N_2660,N_238,N_1629);
nand U2661 (N_2661,N_1170,N_51);
nor U2662 (N_2662,N_358,N_1351);
xor U2663 (N_2663,N_465,N_249);
and U2664 (N_2664,N_746,N_690);
or U2665 (N_2665,N_1259,N_994);
nor U2666 (N_2666,N_840,N_920);
xnor U2667 (N_2667,N_1941,N_1254);
and U2668 (N_2668,N_1339,N_1255);
nor U2669 (N_2669,N_743,N_373);
nor U2670 (N_2670,N_634,N_111);
nor U2671 (N_2671,N_55,N_628);
xnor U2672 (N_2672,N_96,N_1228);
nor U2673 (N_2673,N_74,N_1135);
and U2674 (N_2674,N_1982,N_1536);
or U2675 (N_2675,N_1867,N_283);
and U2676 (N_2676,N_564,N_445);
and U2677 (N_2677,N_1181,N_42);
nand U2678 (N_2678,N_193,N_1223);
and U2679 (N_2679,N_650,N_891);
nand U2680 (N_2680,N_1198,N_312);
or U2681 (N_2681,N_1676,N_126);
xor U2682 (N_2682,N_1391,N_1942);
xnor U2683 (N_2683,N_1042,N_971);
or U2684 (N_2684,N_755,N_295);
nand U2685 (N_2685,N_291,N_590);
nor U2686 (N_2686,N_1677,N_176);
or U2687 (N_2687,N_1579,N_1561);
or U2688 (N_2688,N_1505,N_728);
nor U2689 (N_2689,N_1021,N_955);
xnor U2690 (N_2690,N_843,N_1794);
nand U2691 (N_2691,N_893,N_128);
xor U2692 (N_2692,N_1130,N_911);
nand U2693 (N_2693,N_1467,N_1058);
nand U2694 (N_2694,N_856,N_1312);
xnor U2695 (N_2695,N_1999,N_984);
nand U2696 (N_2696,N_633,N_1804);
or U2697 (N_2697,N_646,N_379);
nand U2698 (N_2698,N_281,N_611);
nand U2699 (N_2699,N_722,N_1325);
nor U2700 (N_2700,N_922,N_1118);
xor U2701 (N_2701,N_386,N_354);
nor U2702 (N_2702,N_204,N_1944);
and U2703 (N_2703,N_342,N_1599);
nor U2704 (N_2704,N_1928,N_1659);
nand U2705 (N_2705,N_470,N_1545);
nor U2706 (N_2706,N_1235,N_309);
nor U2707 (N_2707,N_521,N_563);
or U2708 (N_2708,N_1768,N_1441);
xnor U2709 (N_2709,N_1811,N_925);
nor U2710 (N_2710,N_1580,N_780);
nor U2711 (N_2711,N_81,N_1972);
xnor U2712 (N_2712,N_1455,N_1447);
or U2713 (N_2713,N_376,N_316);
nand U2714 (N_2714,N_1800,N_579);
nand U2715 (N_2715,N_1960,N_58);
or U2716 (N_2716,N_98,N_1810);
xor U2717 (N_2717,N_1821,N_282);
nor U2718 (N_2718,N_1186,N_1572);
or U2719 (N_2719,N_529,N_1190);
nor U2720 (N_2720,N_7,N_1069);
or U2721 (N_2721,N_1092,N_1490);
nand U2722 (N_2722,N_25,N_1379);
or U2723 (N_2723,N_1634,N_88);
nand U2724 (N_2724,N_232,N_1642);
nor U2725 (N_2725,N_167,N_1257);
and U2726 (N_2726,N_1965,N_1380);
and U2727 (N_2727,N_1709,N_764);
nand U2728 (N_2728,N_1500,N_824);
or U2729 (N_2729,N_589,N_699);
xor U2730 (N_2730,N_1885,N_1583);
or U2731 (N_2731,N_1516,N_1390);
and U2732 (N_2732,N_1374,N_1801);
or U2733 (N_2733,N_1044,N_1548);
nand U2734 (N_2734,N_207,N_969);
nand U2735 (N_2735,N_248,N_626);
or U2736 (N_2736,N_1111,N_939);
or U2737 (N_2737,N_1025,N_1697);
nor U2738 (N_2738,N_648,N_39);
nand U2739 (N_2739,N_534,N_1921);
nand U2740 (N_2740,N_254,N_40);
or U2741 (N_2741,N_1299,N_1219);
xnor U2742 (N_2742,N_835,N_584);
xnor U2743 (N_2743,N_1528,N_1301);
and U2744 (N_2744,N_956,N_494);
nor U2745 (N_2745,N_963,N_1956);
nor U2746 (N_2746,N_430,N_1245);
xor U2747 (N_2747,N_659,N_489);
and U2748 (N_2748,N_1300,N_796);
and U2749 (N_2749,N_685,N_1862);
nand U2750 (N_2750,N_1884,N_66);
nand U2751 (N_2751,N_686,N_706);
xor U2752 (N_2752,N_1648,N_432);
xnor U2753 (N_2753,N_702,N_614);
xor U2754 (N_2754,N_1834,N_1620);
nand U2755 (N_2755,N_1435,N_491);
xor U2756 (N_2756,N_142,N_1211);
and U2757 (N_2757,N_1461,N_1933);
nand U2758 (N_2758,N_1964,N_1242);
or U2759 (N_2759,N_325,N_1375);
and U2760 (N_2760,N_1407,N_1166);
or U2761 (N_2761,N_1974,N_298);
nor U2762 (N_2762,N_830,N_380);
and U2763 (N_2763,N_1994,N_182);
and U2764 (N_2764,N_1968,N_396);
or U2765 (N_2765,N_462,N_596);
nand U2766 (N_2766,N_859,N_1932);
nor U2767 (N_2767,N_1636,N_1541);
xnor U2768 (N_2768,N_1989,N_672);
nand U2769 (N_2769,N_1125,N_1287);
xnor U2770 (N_2770,N_91,N_1001);
nor U2771 (N_2771,N_811,N_1752);
and U2772 (N_2772,N_1706,N_1279);
and U2773 (N_2773,N_1070,N_1268);
nand U2774 (N_2774,N_370,N_294);
and U2775 (N_2775,N_1189,N_213);
nand U2776 (N_2776,N_1652,N_1543);
xor U2777 (N_2777,N_1298,N_135);
xor U2778 (N_2778,N_1611,N_151);
xor U2779 (N_2779,N_471,N_1109);
and U2780 (N_2780,N_158,N_946);
xnor U2781 (N_2781,N_1838,N_1477);
or U2782 (N_2782,N_1899,N_497);
nor U2783 (N_2783,N_1946,N_567);
xor U2784 (N_2784,N_968,N_1715);
nand U2785 (N_2785,N_1136,N_1565);
nand U2786 (N_2786,N_1591,N_1064);
xor U2787 (N_2787,N_37,N_1575);
and U2788 (N_2788,N_1641,N_708);
and U2789 (N_2789,N_736,N_286);
nand U2790 (N_2790,N_766,N_357);
xnor U2791 (N_2791,N_1084,N_107);
nand U2792 (N_2792,N_1031,N_987);
nor U2793 (N_2793,N_1327,N_747);
or U2794 (N_2794,N_1420,N_421);
nor U2795 (N_2795,N_1152,N_918);
or U2796 (N_2796,N_181,N_464);
xnor U2797 (N_2797,N_1360,N_1845);
xnor U2798 (N_2798,N_344,N_1525);
or U2799 (N_2799,N_1097,N_638);
nand U2800 (N_2800,N_1818,N_409);
nor U2801 (N_2801,N_1443,N_1703);
nor U2802 (N_2802,N_1749,N_1138);
nor U2803 (N_2803,N_898,N_486);
and U2804 (N_2804,N_1512,N_1322);
xor U2805 (N_2805,N_1496,N_1947);
nand U2806 (N_2806,N_1896,N_1931);
or U2807 (N_2807,N_1584,N_1052);
nor U2808 (N_2808,N_546,N_1524);
nor U2809 (N_2809,N_1854,N_161);
or U2810 (N_2810,N_1878,N_230);
nand U2811 (N_2811,N_954,N_1967);
nand U2812 (N_2812,N_1469,N_86);
nor U2813 (N_2813,N_665,N_27);
nor U2814 (N_2814,N_1159,N_662);
xor U2815 (N_2815,N_1815,N_881);
and U2816 (N_2816,N_1188,N_932);
nor U2817 (N_2817,N_1898,N_304);
nand U2818 (N_2818,N_210,N_1328);
or U2819 (N_2819,N_454,N_1221);
nor U2820 (N_2820,N_300,N_1529);
or U2821 (N_2821,N_1012,N_812);
nor U2822 (N_2822,N_591,N_837);
xnor U2823 (N_2823,N_498,N_540);
and U2824 (N_2824,N_1635,N_1542);
nand U2825 (N_2825,N_1598,N_1802);
or U2826 (N_2826,N_1906,N_275);
or U2827 (N_2827,N_1013,N_1618);
and U2828 (N_2828,N_331,N_1450);
and U2829 (N_2829,N_1765,N_807);
and U2830 (N_2830,N_1763,N_1837);
and U2831 (N_2831,N_1767,N_1939);
nand U2832 (N_2832,N_740,N_256);
nand U2833 (N_2833,N_696,N_356);
and U2834 (N_2834,N_1760,N_395);
and U2835 (N_2835,N_43,N_1187);
xor U2836 (N_2836,N_761,N_1877);
xnor U2837 (N_2837,N_1746,N_1041);
xor U2838 (N_2838,N_803,N_731);
xnor U2839 (N_2839,N_337,N_978);
nand U2840 (N_2840,N_1914,N_1124);
or U2841 (N_2841,N_1131,N_1605);
and U2842 (N_2842,N_347,N_943);
nor U2843 (N_2843,N_1027,N_95);
nand U2844 (N_2844,N_1127,N_401);
nor U2845 (N_2845,N_391,N_861);
and U2846 (N_2846,N_22,N_1662);
xnor U2847 (N_2847,N_1276,N_1917);
nand U2848 (N_2848,N_1442,N_854);
nor U2849 (N_2849,N_1533,N_1789);
nand U2850 (N_2850,N_1148,N_1368);
nand U2851 (N_2851,N_1732,N_444);
and U2852 (N_2852,N_1071,N_554);
xnor U2853 (N_2853,N_1213,N_251);
and U2854 (N_2854,N_289,N_1470);
or U2855 (N_2855,N_214,N_1860);
xor U2856 (N_2856,N_934,N_1423);
and U2857 (N_2857,N_73,N_1632);
or U2858 (N_2858,N_908,N_518);
xnor U2859 (N_2859,N_813,N_774);
nor U2860 (N_2860,N_578,N_851);
and U2861 (N_2861,N_1478,N_523);
and U2862 (N_2862,N_1483,N_235);
nor U2863 (N_2863,N_1949,N_1160);
nor U2864 (N_2864,N_326,N_1145);
or U2865 (N_2865,N_1658,N_649);
and U2866 (N_2866,N_1501,N_560);
or U2867 (N_2867,N_1341,N_53);
nand U2868 (N_2868,N_1285,N_460);
and U2869 (N_2869,N_1691,N_1857);
or U2870 (N_2870,N_1350,N_1908);
or U2871 (N_2871,N_80,N_609);
or U2872 (N_2872,N_1626,N_1880);
nand U2873 (N_2873,N_1849,N_1047);
and U2874 (N_2874,N_241,N_1704);
xnor U2875 (N_2875,N_49,N_1129);
or U2876 (N_2876,N_1907,N_239);
nor U2877 (N_2877,N_1655,N_1429);
and U2878 (N_2878,N_827,N_335);
and U2879 (N_2879,N_188,N_976);
nand U2880 (N_2880,N_862,N_1729);
nand U2881 (N_2881,N_1497,N_307);
nand U2882 (N_2882,N_1872,N_164);
and U2883 (N_2883,N_636,N_65);
or U2884 (N_2884,N_601,N_1101);
xor U2885 (N_2885,N_505,N_466);
nor U2886 (N_2886,N_332,N_1067);
or U2887 (N_2887,N_1511,N_1892);
or U2888 (N_2888,N_613,N_520);
and U2889 (N_2889,N_1358,N_54);
xnor U2890 (N_2890,N_1484,N_439);
xnor U2891 (N_2891,N_1607,N_274);
and U2892 (N_2892,N_10,N_1066);
nor U2893 (N_2893,N_1790,N_527);
nand U2894 (N_2894,N_1117,N_1909);
xnor U2895 (N_2895,N_220,N_410);
nor U2896 (N_2896,N_714,N_1016);
nor U2897 (N_2897,N_753,N_226);
nor U2898 (N_2898,N_935,N_583);
nor U2899 (N_2899,N_475,N_153);
nor U2900 (N_2900,N_1690,N_666);
or U2901 (N_2901,N_772,N_1209);
nand U2902 (N_2902,N_872,N_998);
nor U2903 (N_2903,N_1210,N_1623);
xnor U2904 (N_2904,N_1293,N_186);
or U2905 (N_2905,N_1722,N_930);
nand U2906 (N_2906,N_1032,N_1640);
xor U2907 (N_2907,N_1087,N_271);
nand U2908 (N_2908,N_1056,N_1678);
or U2909 (N_2909,N_1182,N_599);
or U2910 (N_2910,N_1813,N_82);
xnor U2911 (N_2911,N_1534,N_329);
nor U2912 (N_2912,N_545,N_481);
and U2913 (N_2913,N_1451,N_831);
nand U2914 (N_2914,N_1115,N_177);
xor U2915 (N_2915,N_868,N_1009);
nand U2916 (N_2916,N_1797,N_1142);
or U2917 (N_2917,N_1488,N_1604);
xnor U2918 (N_2918,N_1474,N_705);
or U2919 (N_2919,N_1616,N_1785);
nand U2920 (N_2920,N_1950,N_173);
nor U2921 (N_2921,N_1978,N_1425);
nor U2922 (N_2922,N_1158,N_1473);
or U2923 (N_2923,N_6,N_90);
nand U2924 (N_2924,N_1480,N_0);
nor U2925 (N_2925,N_631,N_1144);
nand U2926 (N_2926,N_305,N_449);
xnor U2927 (N_2927,N_556,N_806);
xor U2928 (N_2928,N_622,N_393);
or U2929 (N_2929,N_1197,N_1886);
or U2930 (N_2930,N_1688,N_1132);
nand U2931 (N_2931,N_677,N_1172);
nor U2932 (N_2932,N_1302,N_442);
and U2933 (N_2933,N_732,N_1427);
nand U2934 (N_2934,N_508,N_1940);
or U2935 (N_2935,N_1206,N_1861);
or U2936 (N_2936,N_759,N_1456);
and U2937 (N_2937,N_437,N_644);
and U2938 (N_2938,N_756,N_1236);
xnor U2939 (N_2939,N_1570,N_1615);
nand U2940 (N_2940,N_1365,N_977);
nand U2941 (N_2941,N_818,N_14);
nor U2942 (N_2942,N_1600,N_514);
xnor U2943 (N_2943,N_1779,N_1263);
or U2944 (N_2944,N_1020,N_206);
nor U2945 (N_2945,N_1367,N_1150);
xor U2946 (N_2946,N_1526,N_1888);
and U2947 (N_2947,N_1711,N_1214);
and U2948 (N_2948,N_1347,N_1246);
nand U2949 (N_2949,N_1085,N_1855);
or U2950 (N_2950,N_889,N_1820);
or U2951 (N_2951,N_962,N_16);
nor U2952 (N_2952,N_1781,N_255);
xnor U2953 (N_2953,N_138,N_936);
nor U2954 (N_2954,N_1739,N_1650);
and U2955 (N_2955,N_504,N_928);
or U2956 (N_2956,N_1566,N_133);
xnor U2957 (N_2957,N_1304,N_1664);
nor U2958 (N_2958,N_1165,N_1017);
xor U2959 (N_2959,N_825,N_525);
nor U2960 (N_2960,N_1535,N_808);
xnor U2961 (N_2961,N_1428,N_1075);
xnor U2962 (N_2962,N_1053,N_832);
and U2963 (N_2963,N_472,N_1290);
xor U2964 (N_2964,N_137,N_1226);
or U2965 (N_2965,N_1424,N_947);
nand U2966 (N_2966,N_367,N_202);
or U2967 (N_2967,N_1653,N_1458);
or U2968 (N_2968,N_1753,N_909);
nand U2969 (N_2969,N_1667,N_496);
nor U2970 (N_2970,N_1421,N_1897);
nor U2971 (N_2971,N_1194,N_1881);
nor U2972 (N_2972,N_785,N_652);
nand U2973 (N_2973,N_1225,N_398);
nor U2974 (N_2974,N_1945,N_1229);
or U2975 (N_2975,N_734,N_1764);
or U2976 (N_2976,N_223,N_155);
xor U2977 (N_2977,N_621,N_385);
xnor U2978 (N_2978,N_1799,N_1413);
nor U2979 (N_2979,N_1574,N_33);
nand U2980 (N_2980,N_1104,N_187);
xnor U2981 (N_2981,N_712,N_1338);
xor U2982 (N_2982,N_1783,N_1919);
or U2983 (N_2983,N_855,N_1248);
or U2984 (N_2984,N_1099,N_526);
nand U2985 (N_2985,N_709,N_194);
and U2986 (N_2986,N_1847,N_985);
nand U2987 (N_2987,N_1911,N_323);
nor U2988 (N_2988,N_26,N_362);
or U2989 (N_2989,N_1489,N_869);
and U2990 (N_2990,N_929,N_1106);
nand U2991 (N_2991,N_1920,N_637);
xnor U2992 (N_2992,N_1733,N_461);
and U2993 (N_2993,N_671,N_1227);
xor U2994 (N_2994,N_178,N_1737);
and U2995 (N_2995,N_125,N_1216);
xor U2996 (N_2996,N_41,N_913);
and U2997 (N_2997,N_1865,N_970);
xnor U2998 (N_2998,N_1916,N_1278);
xnor U2999 (N_2999,N_1866,N_76);
nand U3000 (N_3000,N_1797,N_948);
and U3001 (N_3001,N_1205,N_514);
nor U3002 (N_3002,N_1306,N_732);
nor U3003 (N_3003,N_1284,N_1128);
nor U3004 (N_3004,N_1523,N_999);
xnor U3005 (N_3005,N_946,N_1329);
nand U3006 (N_3006,N_1653,N_94);
and U3007 (N_3007,N_1623,N_246);
nor U3008 (N_3008,N_1002,N_686);
or U3009 (N_3009,N_1376,N_1867);
nand U3010 (N_3010,N_188,N_1108);
or U3011 (N_3011,N_1193,N_1951);
nand U3012 (N_3012,N_1074,N_404);
xor U3013 (N_3013,N_1027,N_522);
xor U3014 (N_3014,N_1946,N_1758);
nand U3015 (N_3015,N_1608,N_1019);
nor U3016 (N_3016,N_1947,N_1190);
and U3017 (N_3017,N_1616,N_1516);
nand U3018 (N_3018,N_1923,N_1751);
nand U3019 (N_3019,N_305,N_1764);
xnor U3020 (N_3020,N_1893,N_1810);
nand U3021 (N_3021,N_1169,N_739);
nand U3022 (N_3022,N_1524,N_1759);
nor U3023 (N_3023,N_812,N_1735);
xnor U3024 (N_3024,N_1166,N_1446);
nand U3025 (N_3025,N_1097,N_1022);
and U3026 (N_3026,N_871,N_1933);
xnor U3027 (N_3027,N_1013,N_917);
and U3028 (N_3028,N_868,N_1293);
nand U3029 (N_3029,N_1459,N_1303);
xor U3030 (N_3030,N_1060,N_567);
xnor U3031 (N_3031,N_812,N_1373);
xor U3032 (N_3032,N_1391,N_95);
nor U3033 (N_3033,N_505,N_261);
and U3034 (N_3034,N_1321,N_334);
nor U3035 (N_3035,N_425,N_876);
or U3036 (N_3036,N_1995,N_373);
xnor U3037 (N_3037,N_473,N_1679);
nor U3038 (N_3038,N_1216,N_1468);
or U3039 (N_3039,N_1628,N_1409);
nor U3040 (N_3040,N_534,N_1404);
and U3041 (N_3041,N_1946,N_1812);
xor U3042 (N_3042,N_10,N_428);
and U3043 (N_3043,N_1002,N_1173);
or U3044 (N_3044,N_519,N_435);
or U3045 (N_3045,N_1716,N_864);
and U3046 (N_3046,N_1221,N_1464);
xnor U3047 (N_3047,N_1680,N_180);
nor U3048 (N_3048,N_1752,N_561);
and U3049 (N_3049,N_525,N_979);
nand U3050 (N_3050,N_1731,N_32);
nand U3051 (N_3051,N_1609,N_297);
xor U3052 (N_3052,N_61,N_2);
or U3053 (N_3053,N_1595,N_1133);
and U3054 (N_3054,N_1339,N_299);
nand U3055 (N_3055,N_1704,N_263);
or U3056 (N_3056,N_1777,N_1095);
nand U3057 (N_3057,N_1394,N_145);
or U3058 (N_3058,N_1299,N_173);
and U3059 (N_3059,N_677,N_1701);
nand U3060 (N_3060,N_1171,N_1582);
and U3061 (N_3061,N_121,N_1098);
nand U3062 (N_3062,N_851,N_1236);
xnor U3063 (N_3063,N_1285,N_1017);
nor U3064 (N_3064,N_28,N_1406);
nand U3065 (N_3065,N_1322,N_61);
nand U3066 (N_3066,N_635,N_1603);
and U3067 (N_3067,N_1003,N_1743);
xor U3068 (N_3068,N_1852,N_1922);
xnor U3069 (N_3069,N_387,N_713);
and U3070 (N_3070,N_1923,N_1007);
xor U3071 (N_3071,N_907,N_87);
nand U3072 (N_3072,N_825,N_1260);
xnor U3073 (N_3073,N_492,N_990);
nand U3074 (N_3074,N_442,N_1588);
or U3075 (N_3075,N_636,N_1869);
nand U3076 (N_3076,N_476,N_333);
nor U3077 (N_3077,N_634,N_433);
xnor U3078 (N_3078,N_469,N_1982);
nor U3079 (N_3079,N_1092,N_887);
or U3080 (N_3080,N_1903,N_788);
xor U3081 (N_3081,N_1163,N_905);
nand U3082 (N_3082,N_502,N_1987);
xor U3083 (N_3083,N_1591,N_96);
nand U3084 (N_3084,N_517,N_374);
or U3085 (N_3085,N_1780,N_1510);
nor U3086 (N_3086,N_317,N_1663);
and U3087 (N_3087,N_662,N_592);
nor U3088 (N_3088,N_1365,N_695);
nand U3089 (N_3089,N_961,N_1559);
or U3090 (N_3090,N_787,N_1711);
xnor U3091 (N_3091,N_655,N_752);
nand U3092 (N_3092,N_153,N_854);
nand U3093 (N_3093,N_682,N_766);
or U3094 (N_3094,N_661,N_1610);
nand U3095 (N_3095,N_1931,N_766);
and U3096 (N_3096,N_1380,N_707);
nand U3097 (N_3097,N_935,N_639);
nand U3098 (N_3098,N_193,N_113);
or U3099 (N_3099,N_1049,N_1982);
nand U3100 (N_3100,N_1324,N_1778);
and U3101 (N_3101,N_17,N_1785);
xor U3102 (N_3102,N_1748,N_928);
and U3103 (N_3103,N_1647,N_1809);
or U3104 (N_3104,N_452,N_927);
or U3105 (N_3105,N_873,N_1805);
and U3106 (N_3106,N_115,N_610);
nand U3107 (N_3107,N_1412,N_757);
nand U3108 (N_3108,N_1841,N_686);
or U3109 (N_3109,N_1310,N_1608);
nand U3110 (N_3110,N_92,N_495);
xor U3111 (N_3111,N_1283,N_1372);
nor U3112 (N_3112,N_1792,N_500);
xor U3113 (N_3113,N_1205,N_245);
nor U3114 (N_3114,N_1779,N_618);
or U3115 (N_3115,N_392,N_593);
or U3116 (N_3116,N_570,N_767);
xor U3117 (N_3117,N_1368,N_1039);
or U3118 (N_3118,N_367,N_1358);
nor U3119 (N_3119,N_970,N_1611);
nand U3120 (N_3120,N_1925,N_1163);
and U3121 (N_3121,N_1461,N_738);
xnor U3122 (N_3122,N_1230,N_157);
xnor U3123 (N_3123,N_1633,N_640);
and U3124 (N_3124,N_1777,N_849);
xor U3125 (N_3125,N_95,N_283);
or U3126 (N_3126,N_1384,N_482);
xor U3127 (N_3127,N_1230,N_1970);
and U3128 (N_3128,N_1859,N_1944);
and U3129 (N_3129,N_1495,N_1963);
and U3130 (N_3130,N_247,N_1681);
or U3131 (N_3131,N_1918,N_1817);
nor U3132 (N_3132,N_1839,N_313);
xor U3133 (N_3133,N_1905,N_1588);
or U3134 (N_3134,N_684,N_944);
nor U3135 (N_3135,N_1852,N_257);
and U3136 (N_3136,N_1972,N_1069);
or U3137 (N_3137,N_418,N_1668);
nor U3138 (N_3138,N_1610,N_185);
nand U3139 (N_3139,N_916,N_137);
xnor U3140 (N_3140,N_604,N_60);
nor U3141 (N_3141,N_663,N_111);
xor U3142 (N_3142,N_1807,N_1888);
xor U3143 (N_3143,N_612,N_921);
nand U3144 (N_3144,N_134,N_1145);
nor U3145 (N_3145,N_1635,N_551);
and U3146 (N_3146,N_914,N_138);
or U3147 (N_3147,N_1287,N_708);
and U3148 (N_3148,N_997,N_669);
nand U3149 (N_3149,N_851,N_786);
and U3150 (N_3150,N_917,N_1927);
nor U3151 (N_3151,N_222,N_1194);
nor U3152 (N_3152,N_1029,N_1938);
or U3153 (N_3153,N_1184,N_303);
nand U3154 (N_3154,N_964,N_1426);
xnor U3155 (N_3155,N_1824,N_1701);
nor U3156 (N_3156,N_1069,N_1093);
nor U3157 (N_3157,N_358,N_1520);
and U3158 (N_3158,N_1369,N_1473);
nand U3159 (N_3159,N_863,N_1880);
nand U3160 (N_3160,N_898,N_1107);
xor U3161 (N_3161,N_1790,N_972);
xor U3162 (N_3162,N_358,N_1304);
nor U3163 (N_3163,N_342,N_1030);
and U3164 (N_3164,N_276,N_868);
and U3165 (N_3165,N_567,N_1127);
xnor U3166 (N_3166,N_868,N_913);
nand U3167 (N_3167,N_1888,N_114);
or U3168 (N_3168,N_942,N_1947);
nand U3169 (N_3169,N_1041,N_1302);
and U3170 (N_3170,N_1347,N_1064);
xnor U3171 (N_3171,N_1289,N_1234);
nor U3172 (N_3172,N_225,N_1355);
nand U3173 (N_3173,N_1197,N_1401);
nor U3174 (N_3174,N_899,N_64);
or U3175 (N_3175,N_667,N_1627);
nor U3176 (N_3176,N_1684,N_343);
nor U3177 (N_3177,N_915,N_1251);
nand U3178 (N_3178,N_1021,N_1330);
xor U3179 (N_3179,N_534,N_668);
nand U3180 (N_3180,N_852,N_598);
nor U3181 (N_3181,N_865,N_581);
and U3182 (N_3182,N_300,N_567);
nor U3183 (N_3183,N_1357,N_1737);
xnor U3184 (N_3184,N_57,N_289);
and U3185 (N_3185,N_660,N_1399);
nand U3186 (N_3186,N_1501,N_1492);
or U3187 (N_3187,N_942,N_636);
nor U3188 (N_3188,N_1654,N_1115);
or U3189 (N_3189,N_145,N_1391);
nand U3190 (N_3190,N_70,N_347);
nand U3191 (N_3191,N_832,N_918);
or U3192 (N_3192,N_527,N_478);
nand U3193 (N_3193,N_1152,N_1709);
xor U3194 (N_3194,N_1092,N_1646);
xor U3195 (N_3195,N_267,N_701);
nor U3196 (N_3196,N_8,N_469);
nor U3197 (N_3197,N_904,N_178);
nor U3198 (N_3198,N_1912,N_470);
or U3199 (N_3199,N_491,N_1311);
nor U3200 (N_3200,N_751,N_179);
nor U3201 (N_3201,N_1229,N_1913);
or U3202 (N_3202,N_1343,N_837);
nor U3203 (N_3203,N_674,N_364);
or U3204 (N_3204,N_468,N_1405);
nand U3205 (N_3205,N_105,N_935);
xnor U3206 (N_3206,N_591,N_724);
nand U3207 (N_3207,N_1893,N_651);
or U3208 (N_3208,N_1437,N_1891);
nand U3209 (N_3209,N_1946,N_1256);
nand U3210 (N_3210,N_1066,N_1284);
or U3211 (N_3211,N_659,N_1854);
or U3212 (N_3212,N_453,N_1482);
xnor U3213 (N_3213,N_1801,N_358);
xor U3214 (N_3214,N_1247,N_1085);
nand U3215 (N_3215,N_249,N_741);
and U3216 (N_3216,N_1754,N_1482);
nand U3217 (N_3217,N_756,N_1393);
and U3218 (N_3218,N_225,N_1223);
nor U3219 (N_3219,N_1049,N_970);
or U3220 (N_3220,N_43,N_186);
nand U3221 (N_3221,N_1661,N_1928);
and U3222 (N_3222,N_1332,N_1738);
or U3223 (N_3223,N_908,N_8);
and U3224 (N_3224,N_506,N_605);
nand U3225 (N_3225,N_643,N_1518);
nor U3226 (N_3226,N_568,N_78);
and U3227 (N_3227,N_493,N_1568);
nand U3228 (N_3228,N_927,N_1197);
or U3229 (N_3229,N_1893,N_708);
nor U3230 (N_3230,N_724,N_1853);
and U3231 (N_3231,N_1432,N_435);
nor U3232 (N_3232,N_1264,N_750);
nand U3233 (N_3233,N_1965,N_1994);
nor U3234 (N_3234,N_1641,N_1340);
or U3235 (N_3235,N_69,N_350);
nand U3236 (N_3236,N_1169,N_1998);
xor U3237 (N_3237,N_417,N_1714);
xnor U3238 (N_3238,N_631,N_1178);
and U3239 (N_3239,N_807,N_1293);
or U3240 (N_3240,N_945,N_1693);
and U3241 (N_3241,N_66,N_540);
or U3242 (N_3242,N_1949,N_325);
and U3243 (N_3243,N_716,N_582);
xor U3244 (N_3244,N_588,N_660);
and U3245 (N_3245,N_1859,N_1872);
and U3246 (N_3246,N_537,N_723);
nor U3247 (N_3247,N_892,N_1380);
and U3248 (N_3248,N_967,N_1487);
nand U3249 (N_3249,N_1045,N_1981);
nand U3250 (N_3250,N_491,N_40);
and U3251 (N_3251,N_1042,N_902);
nand U3252 (N_3252,N_1856,N_263);
nand U3253 (N_3253,N_1912,N_1434);
nor U3254 (N_3254,N_246,N_757);
nor U3255 (N_3255,N_1395,N_338);
or U3256 (N_3256,N_938,N_1288);
xor U3257 (N_3257,N_41,N_386);
nand U3258 (N_3258,N_1692,N_747);
nor U3259 (N_3259,N_632,N_348);
xor U3260 (N_3260,N_1670,N_183);
nand U3261 (N_3261,N_1423,N_342);
or U3262 (N_3262,N_1396,N_1357);
or U3263 (N_3263,N_812,N_1142);
nand U3264 (N_3264,N_347,N_405);
nand U3265 (N_3265,N_35,N_1866);
nand U3266 (N_3266,N_1380,N_592);
nor U3267 (N_3267,N_389,N_1459);
and U3268 (N_3268,N_824,N_848);
and U3269 (N_3269,N_1951,N_810);
xor U3270 (N_3270,N_1673,N_784);
and U3271 (N_3271,N_152,N_337);
or U3272 (N_3272,N_15,N_372);
nor U3273 (N_3273,N_785,N_1099);
nor U3274 (N_3274,N_596,N_1284);
xnor U3275 (N_3275,N_154,N_1658);
xnor U3276 (N_3276,N_295,N_1417);
nor U3277 (N_3277,N_900,N_1408);
xor U3278 (N_3278,N_148,N_1878);
nor U3279 (N_3279,N_334,N_982);
and U3280 (N_3280,N_1010,N_1096);
xnor U3281 (N_3281,N_1833,N_832);
nand U3282 (N_3282,N_571,N_1218);
xnor U3283 (N_3283,N_1745,N_1916);
and U3284 (N_3284,N_1572,N_1781);
nor U3285 (N_3285,N_919,N_928);
and U3286 (N_3286,N_1062,N_527);
nor U3287 (N_3287,N_1211,N_1550);
or U3288 (N_3288,N_646,N_1717);
xnor U3289 (N_3289,N_1334,N_1735);
or U3290 (N_3290,N_1455,N_1133);
and U3291 (N_3291,N_1628,N_812);
xnor U3292 (N_3292,N_1916,N_1866);
and U3293 (N_3293,N_1535,N_1319);
and U3294 (N_3294,N_1306,N_1230);
nand U3295 (N_3295,N_650,N_964);
xor U3296 (N_3296,N_471,N_437);
nand U3297 (N_3297,N_1225,N_323);
and U3298 (N_3298,N_335,N_1517);
nor U3299 (N_3299,N_335,N_1316);
nand U3300 (N_3300,N_366,N_1961);
xor U3301 (N_3301,N_426,N_1490);
nand U3302 (N_3302,N_1157,N_1315);
or U3303 (N_3303,N_1950,N_1010);
and U3304 (N_3304,N_479,N_931);
or U3305 (N_3305,N_800,N_1121);
or U3306 (N_3306,N_1178,N_1722);
nand U3307 (N_3307,N_1994,N_1614);
nor U3308 (N_3308,N_676,N_1491);
nor U3309 (N_3309,N_411,N_1652);
and U3310 (N_3310,N_788,N_389);
and U3311 (N_3311,N_1650,N_1687);
or U3312 (N_3312,N_738,N_498);
xor U3313 (N_3313,N_1051,N_1867);
nand U3314 (N_3314,N_672,N_879);
nor U3315 (N_3315,N_685,N_220);
xor U3316 (N_3316,N_1753,N_1867);
xnor U3317 (N_3317,N_1951,N_862);
and U3318 (N_3318,N_1167,N_1803);
and U3319 (N_3319,N_1505,N_1554);
nand U3320 (N_3320,N_1065,N_528);
or U3321 (N_3321,N_261,N_126);
xor U3322 (N_3322,N_1710,N_310);
and U3323 (N_3323,N_803,N_289);
xnor U3324 (N_3324,N_205,N_395);
or U3325 (N_3325,N_595,N_1657);
nor U3326 (N_3326,N_1431,N_1821);
and U3327 (N_3327,N_347,N_272);
nand U3328 (N_3328,N_1699,N_1730);
xnor U3329 (N_3329,N_562,N_339);
xor U3330 (N_3330,N_703,N_1248);
nor U3331 (N_3331,N_1565,N_470);
nand U3332 (N_3332,N_906,N_1504);
nor U3333 (N_3333,N_1172,N_1940);
nor U3334 (N_3334,N_1920,N_1522);
nand U3335 (N_3335,N_142,N_994);
xor U3336 (N_3336,N_1743,N_1291);
nand U3337 (N_3337,N_1634,N_1796);
and U3338 (N_3338,N_1881,N_1023);
nand U3339 (N_3339,N_1831,N_25);
nor U3340 (N_3340,N_1542,N_1810);
nor U3341 (N_3341,N_1491,N_1617);
xnor U3342 (N_3342,N_489,N_1207);
nor U3343 (N_3343,N_456,N_51);
nor U3344 (N_3344,N_1141,N_699);
nor U3345 (N_3345,N_349,N_588);
nor U3346 (N_3346,N_968,N_1187);
or U3347 (N_3347,N_594,N_1508);
and U3348 (N_3348,N_1876,N_1161);
nor U3349 (N_3349,N_985,N_1405);
nor U3350 (N_3350,N_1752,N_1616);
nand U3351 (N_3351,N_181,N_1457);
or U3352 (N_3352,N_850,N_841);
xor U3353 (N_3353,N_1346,N_1473);
nor U3354 (N_3354,N_1935,N_1873);
nor U3355 (N_3355,N_1271,N_412);
xor U3356 (N_3356,N_484,N_1340);
and U3357 (N_3357,N_435,N_1544);
nand U3358 (N_3358,N_435,N_1776);
nand U3359 (N_3359,N_101,N_1796);
nand U3360 (N_3360,N_604,N_517);
and U3361 (N_3361,N_591,N_786);
nor U3362 (N_3362,N_1780,N_1264);
or U3363 (N_3363,N_1230,N_804);
nor U3364 (N_3364,N_1159,N_603);
xor U3365 (N_3365,N_1822,N_1270);
nand U3366 (N_3366,N_830,N_240);
nand U3367 (N_3367,N_273,N_433);
and U3368 (N_3368,N_1652,N_1298);
nand U3369 (N_3369,N_453,N_1181);
xor U3370 (N_3370,N_1861,N_205);
nand U3371 (N_3371,N_1248,N_897);
nand U3372 (N_3372,N_419,N_1565);
or U3373 (N_3373,N_1863,N_1737);
xor U3374 (N_3374,N_228,N_1677);
and U3375 (N_3375,N_366,N_532);
and U3376 (N_3376,N_1015,N_997);
xor U3377 (N_3377,N_1247,N_291);
xor U3378 (N_3378,N_1363,N_1116);
xor U3379 (N_3379,N_232,N_1948);
nand U3380 (N_3380,N_1317,N_1959);
nand U3381 (N_3381,N_9,N_985);
and U3382 (N_3382,N_1261,N_973);
nor U3383 (N_3383,N_795,N_1723);
and U3384 (N_3384,N_961,N_1955);
and U3385 (N_3385,N_157,N_1695);
nand U3386 (N_3386,N_724,N_1613);
nor U3387 (N_3387,N_1426,N_1622);
or U3388 (N_3388,N_883,N_1106);
xor U3389 (N_3389,N_957,N_972);
nor U3390 (N_3390,N_1411,N_1179);
nand U3391 (N_3391,N_1245,N_1174);
xor U3392 (N_3392,N_1059,N_1834);
xnor U3393 (N_3393,N_1747,N_1314);
nand U3394 (N_3394,N_1213,N_1116);
nor U3395 (N_3395,N_374,N_1208);
nor U3396 (N_3396,N_1149,N_1304);
and U3397 (N_3397,N_938,N_1412);
xnor U3398 (N_3398,N_332,N_640);
or U3399 (N_3399,N_826,N_1067);
nand U3400 (N_3400,N_215,N_1202);
xnor U3401 (N_3401,N_114,N_1983);
and U3402 (N_3402,N_1004,N_1965);
xor U3403 (N_3403,N_799,N_1879);
or U3404 (N_3404,N_1793,N_1029);
nand U3405 (N_3405,N_1826,N_1997);
nand U3406 (N_3406,N_873,N_727);
nand U3407 (N_3407,N_1481,N_1200);
and U3408 (N_3408,N_1004,N_885);
nor U3409 (N_3409,N_1773,N_406);
xnor U3410 (N_3410,N_1917,N_233);
xor U3411 (N_3411,N_522,N_188);
xnor U3412 (N_3412,N_253,N_887);
nand U3413 (N_3413,N_236,N_1293);
xor U3414 (N_3414,N_1221,N_1572);
or U3415 (N_3415,N_1234,N_115);
or U3416 (N_3416,N_1236,N_777);
and U3417 (N_3417,N_863,N_639);
or U3418 (N_3418,N_92,N_52);
xnor U3419 (N_3419,N_497,N_897);
nand U3420 (N_3420,N_1952,N_1327);
nor U3421 (N_3421,N_65,N_727);
nand U3422 (N_3422,N_1077,N_1261);
nor U3423 (N_3423,N_631,N_541);
nor U3424 (N_3424,N_1916,N_422);
nand U3425 (N_3425,N_82,N_927);
nand U3426 (N_3426,N_546,N_84);
or U3427 (N_3427,N_980,N_1744);
nand U3428 (N_3428,N_1405,N_285);
nor U3429 (N_3429,N_1121,N_309);
nand U3430 (N_3430,N_677,N_898);
and U3431 (N_3431,N_1592,N_566);
or U3432 (N_3432,N_732,N_906);
nor U3433 (N_3433,N_605,N_949);
xor U3434 (N_3434,N_450,N_567);
or U3435 (N_3435,N_580,N_1928);
nand U3436 (N_3436,N_1199,N_1669);
xnor U3437 (N_3437,N_176,N_1007);
xnor U3438 (N_3438,N_652,N_677);
and U3439 (N_3439,N_1453,N_1098);
or U3440 (N_3440,N_588,N_1584);
nand U3441 (N_3441,N_1559,N_1908);
nand U3442 (N_3442,N_8,N_1857);
xor U3443 (N_3443,N_748,N_689);
nor U3444 (N_3444,N_172,N_1414);
or U3445 (N_3445,N_690,N_159);
xor U3446 (N_3446,N_484,N_252);
nor U3447 (N_3447,N_1763,N_1553);
or U3448 (N_3448,N_955,N_272);
nor U3449 (N_3449,N_1206,N_1122);
xor U3450 (N_3450,N_1835,N_693);
nor U3451 (N_3451,N_1069,N_1084);
and U3452 (N_3452,N_1333,N_430);
or U3453 (N_3453,N_1362,N_1557);
nor U3454 (N_3454,N_1401,N_1460);
and U3455 (N_3455,N_223,N_607);
xnor U3456 (N_3456,N_1633,N_1447);
or U3457 (N_3457,N_1948,N_1671);
or U3458 (N_3458,N_470,N_1979);
nor U3459 (N_3459,N_387,N_632);
nor U3460 (N_3460,N_380,N_1008);
nand U3461 (N_3461,N_1119,N_1863);
or U3462 (N_3462,N_10,N_1138);
or U3463 (N_3463,N_766,N_392);
nand U3464 (N_3464,N_1719,N_812);
xor U3465 (N_3465,N_158,N_1318);
nand U3466 (N_3466,N_375,N_1267);
nand U3467 (N_3467,N_556,N_257);
nor U3468 (N_3468,N_54,N_1239);
or U3469 (N_3469,N_943,N_1310);
or U3470 (N_3470,N_1165,N_101);
nor U3471 (N_3471,N_1464,N_697);
or U3472 (N_3472,N_964,N_562);
and U3473 (N_3473,N_808,N_840);
and U3474 (N_3474,N_752,N_491);
nand U3475 (N_3475,N_1443,N_1638);
nor U3476 (N_3476,N_1319,N_819);
nand U3477 (N_3477,N_1749,N_388);
xnor U3478 (N_3478,N_315,N_1977);
xnor U3479 (N_3479,N_901,N_1540);
nand U3480 (N_3480,N_669,N_1960);
nand U3481 (N_3481,N_21,N_1413);
nand U3482 (N_3482,N_27,N_1268);
xor U3483 (N_3483,N_1161,N_1072);
nor U3484 (N_3484,N_1700,N_1692);
or U3485 (N_3485,N_1746,N_69);
and U3486 (N_3486,N_959,N_751);
or U3487 (N_3487,N_1824,N_141);
nand U3488 (N_3488,N_623,N_1387);
nand U3489 (N_3489,N_958,N_965);
or U3490 (N_3490,N_1976,N_129);
nand U3491 (N_3491,N_841,N_1086);
xnor U3492 (N_3492,N_321,N_368);
nor U3493 (N_3493,N_747,N_1630);
nor U3494 (N_3494,N_1569,N_1357);
nand U3495 (N_3495,N_142,N_601);
and U3496 (N_3496,N_1970,N_1165);
xor U3497 (N_3497,N_109,N_1044);
nand U3498 (N_3498,N_1788,N_93);
nor U3499 (N_3499,N_1518,N_533);
nor U3500 (N_3500,N_1526,N_290);
and U3501 (N_3501,N_621,N_830);
nor U3502 (N_3502,N_630,N_1700);
or U3503 (N_3503,N_1340,N_1499);
or U3504 (N_3504,N_266,N_731);
nor U3505 (N_3505,N_17,N_795);
nand U3506 (N_3506,N_1761,N_1959);
nor U3507 (N_3507,N_200,N_1749);
and U3508 (N_3508,N_1742,N_169);
or U3509 (N_3509,N_146,N_1522);
nor U3510 (N_3510,N_975,N_1087);
and U3511 (N_3511,N_16,N_1248);
nand U3512 (N_3512,N_100,N_379);
nand U3513 (N_3513,N_23,N_109);
nand U3514 (N_3514,N_1238,N_725);
nor U3515 (N_3515,N_1790,N_595);
xor U3516 (N_3516,N_1857,N_1019);
xor U3517 (N_3517,N_1499,N_779);
and U3518 (N_3518,N_1306,N_1057);
xor U3519 (N_3519,N_1090,N_1313);
and U3520 (N_3520,N_716,N_110);
xnor U3521 (N_3521,N_1776,N_303);
and U3522 (N_3522,N_1488,N_311);
or U3523 (N_3523,N_663,N_1236);
nor U3524 (N_3524,N_1591,N_1576);
nand U3525 (N_3525,N_461,N_1125);
or U3526 (N_3526,N_1140,N_157);
and U3527 (N_3527,N_632,N_1025);
or U3528 (N_3528,N_1939,N_398);
nor U3529 (N_3529,N_778,N_1749);
and U3530 (N_3530,N_1484,N_377);
nor U3531 (N_3531,N_393,N_985);
or U3532 (N_3532,N_1862,N_565);
nand U3533 (N_3533,N_163,N_1148);
or U3534 (N_3534,N_366,N_802);
and U3535 (N_3535,N_1909,N_277);
nor U3536 (N_3536,N_167,N_1607);
and U3537 (N_3537,N_532,N_1815);
and U3538 (N_3538,N_436,N_51);
or U3539 (N_3539,N_1154,N_45);
nand U3540 (N_3540,N_1439,N_1676);
nor U3541 (N_3541,N_740,N_1950);
and U3542 (N_3542,N_31,N_1732);
and U3543 (N_3543,N_660,N_1338);
and U3544 (N_3544,N_1773,N_784);
or U3545 (N_3545,N_1025,N_360);
and U3546 (N_3546,N_984,N_1516);
xnor U3547 (N_3547,N_1940,N_1326);
nor U3548 (N_3548,N_11,N_1847);
xnor U3549 (N_3549,N_438,N_732);
and U3550 (N_3550,N_1435,N_1068);
nand U3551 (N_3551,N_1266,N_1041);
nand U3552 (N_3552,N_1772,N_1706);
nor U3553 (N_3553,N_1263,N_360);
and U3554 (N_3554,N_514,N_1639);
and U3555 (N_3555,N_1010,N_397);
nand U3556 (N_3556,N_186,N_1661);
or U3557 (N_3557,N_114,N_1145);
nor U3558 (N_3558,N_1443,N_667);
and U3559 (N_3559,N_1410,N_390);
nand U3560 (N_3560,N_1258,N_401);
nand U3561 (N_3561,N_476,N_1237);
and U3562 (N_3562,N_712,N_802);
xor U3563 (N_3563,N_1783,N_761);
xnor U3564 (N_3564,N_757,N_771);
and U3565 (N_3565,N_171,N_266);
xor U3566 (N_3566,N_1610,N_1708);
or U3567 (N_3567,N_1445,N_1012);
nand U3568 (N_3568,N_1853,N_73);
xnor U3569 (N_3569,N_514,N_1034);
and U3570 (N_3570,N_39,N_595);
nand U3571 (N_3571,N_1847,N_1928);
xor U3572 (N_3572,N_935,N_1065);
and U3573 (N_3573,N_306,N_501);
nand U3574 (N_3574,N_1175,N_1515);
or U3575 (N_3575,N_21,N_1659);
and U3576 (N_3576,N_46,N_896);
xor U3577 (N_3577,N_557,N_1818);
and U3578 (N_3578,N_1685,N_535);
or U3579 (N_3579,N_163,N_37);
xnor U3580 (N_3580,N_778,N_1342);
xnor U3581 (N_3581,N_1792,N_1281);
xnor U3582 (N_3582,N_1353,N_1891);
xor U3583 (N_3583,N_1467,N_86);
xor U3584 (N_3584,N_1539,N_781);
and U3585 (N_3585,N_1783,N_199);
and U3586 (N_3586,N_1757,N_1091);
or U3587 (N_3587,N_1368,N_1583);
xor U3588 (N_3588,N_1326,N_55);
nand U3589 (N_3589,N_1837,N_1291);
nor U3590 (N_3590,N_861,N_1761);
nor U3591 (N_3591,N_1512,N_1645);
and U3592 (N_3592,N_611,N_942);
and U3593 (N_3593,N_1487,N_1777);
or U3594 (N_3594,N_1916,N_469);
and U3595 (N_3595,N_1487,N_653);
and U3596 (N_3596,N_1839,N_1375);
and U3597 (N_3597,N_4,N_962);
nand U3598 (N_3598,N_118,N_1345);
nand U3599 (N_3599,N_707,N_1268);
xnor U3600 (N_3600,N_1948,N_1844);
nand U3601 (N_3601,N_1105,N_1574);
or U3602 (N_3602,N_443,N_1812);
and U3603 (N_3603,N_1276,N_175);
and U3604 (N_3604,N_40,N_782);
xor U3605 (N_3605,N_1845,N_1116);
nand U3606 (N_3606,N_1897,N_728);
or U3607 (N_3607,N_1938,N_1971);
nor U3608 (N_3608,N_579,N_1476);
and U3609 (N_3609,N_1846,N_780);
xnor U3610 (N_3610,N_1032,N_778);
and U3611 (N_3611,N_1492,N_1916);
nor U3612 (N_3612,N_122,N_607);
and U3613 (N_3613,N_1278,N_730);
or U3614 (N_3614,N_1915,N_424);
nor U3615 (N_3615,N_1201,N_1032);
or U3616 (N_3616,N_1563,N_1295);
xor U3617 (N_3617,N_988,N_826);
or U3618 (N_3618,N_1274,N_765);
xor U3619 (N_3619,N_544,N_1870);
nand U3620 (N_3620,N_1338,N_1514);
nand U3621 (N_3621,N_1052,N_912);
xnor U3622 (N_3622,N_1103,N_572);
nand U3623 (N_3623,N_160,N_347);
xnor U3624 (N_3624,N_825,N_1246);
and U3625 (N_3625,N_700,N_803);
nand U3626 (N_3626,N_482,N_942);
and U3627 (N_3627,N_1678,N_1042);
xnor U3628 (N_3628,N_1034,N_1950);
xor U3629 (N_3629,N_406,N_378);
nor U3630 (N_3630,N_1090,N_1531);
and U3631 (N_3631,N_582,N_809);
nor U3632 (N_3632,N_1300,N_43);
xnor U3633 (N_3633,N_268,N_986);
nor U3634 (N_3634,N_183,N_820);
nand U3635 (N_3635,N_156,N_966);
xor U3636 (N_3636,N_1337,N_1500);
xor U3637 (N_3637,N_1364,N_1154);
nand U3638 (N_3638,N_1450,N_1416);
nand U3639 (N_3639,N_1229,N_1608);
and U3640 (N_3640,N_1584,N_398);
nor U3641 (N_3641,N_431,N_12);
or U3642 (N_3642,N_1478,N_1725);
and U3643 (N_3643,N_342,N_1734);
nor U3644 (N_3644,N_1089,N_353);
and U3645 (N_3645,N_74,N_435);
or U3646 (N_3646,N_1804,N_916);
xnor U3647 (N_3647,N_102,N_1066);
xnor U3648 (N_3648,N_1099,N_1513);
and U3649 (N_3649,N_160,N_1013);
or U3650 (N_3650,N_973,N_497);
xor U3651 (N_3651,N_867,N_900);
nor U3652 (N_3652,N_1070,N_439);
or U3653 (N_3653,N_640,N_916);
xor U3654 (N_3654,N_240,N_363);
and U3655 (N_3655,N_1725,N_948);
and U3656 (N_3656,N_629,N_1025);
and U3657 (N_3657,N_1170,N_1940);
nor U3658 (N_3658,N_1213,N_1946);
xor U3659 (N_3659,N_1147,N_1316);
nand U3660 (N_3660,N_442,N_803);
nand U3661 (N_3661,N_1107,N_1739);
xnor U3662 (N_3662,N_1400,N_1680);
xnor U3663 (N_3663,N_681,N_940);
nor U3664 (N_3664,N_905,N_1703);
and U3665 (N_3665,N_9,N_1377);
nand U3666 (N_3666,N_2,N_1676);
or U3667 (N_3667,N_695,N_1374);
nor U3668 (N_3668,N_412,N_1317);
xor U3669 (N_3669,N_87,N_691);
or U3670 (N_3670,N_819,N_1310);
and U3671 (N_3671,N_797,N_1699);
and U3672 (N_3672,N_1264,N_1245);
nand U3673 (N_3673,N_1415,N_1173);
and U3674 (N_3674,N_1643,N_1765);
xor U3675 (N_3675,N_766,N_733);
xor U3676 (N_3676,N_1808,N_1560);
or U3677 (N_3677,N_1270,N_473);
and U3678 (N_3678,N_897,N_816);
xor U3679 (N_3679,N_868,N_728);
xnor U3680 (N_3680,N_670,N_1997);
nor U3681 (N_3681,N_1169,N_405);
and U3682 (N_3682,N_349,N_1569);
nor U3683 (N_3683,N_1601,N_20);
nand U3684 (N_3684,N_1615,N_450);
nand U3685 (N_3685,N_557,N_962);
nand U3686 (N_3686,N_803,N_202);
xnor U3687 (N_3687,N_33,N_1942);
and U3688 (N_3688,N_1368,N_480);
nand U3689 (N_3689,N_765,N_635);
and U3690 (N_3690,N_1304,N_1378);
and U3691 (N_3691,N_1193,N_838);
and U3692 (N_3692,N_1023,N_198);
nor U3693 (N_3693,N_97,N_1675);
and U3694 (N_3694,N_1287,N_1255);
nor U3695 (N_3695,N_935,N_1792);
or U3696 (N_3696,N_71,N_359);
or U3697 (N_3697,N_801,N_1935);
or U3698 (N_3698,N_1508,N_728);
and U3699 (N_3699,N_452,N_1529);
and U3700 (N_3700,N_205,N_1453);
xnor U3701 (N_3701,N_1304,N_1609);
or U3702 (N_3702,N_1501,N_323);
xor U3703 (N_3703,N_1420,N_735);
nor U3704 (N_3704,N_987,N_1723);
and U3705 (N_3705,N_1770,N_1935);
nor U3706 (N_3706,N_65,N_1025);
xnor U3707 (N_3707,N_874,N_1670);
xnor U3708 (N_3708,N_254,N_704);
nor U3709 (N_3709,N_570,N_957);
xnor U3710 (N_3710,N_1226,N_741);
nand U3711 (N_3711,N_1340,N_1335);
xnor U3712 (N_3712,N_265,N_334);
or U3713 (N_3713,N_310,N_1052);
xnor U3714 (N_3714,N_1850,N_99);
nor U3715 (N_3715,N_1912,N_566);
xor U3716 (N_3716,N_1786,N_1222);
nand U3717 (N_3717,N_762,N_471);
or U3718 (N_3718,N_337,N_26);
xor U3719 (N_3719,N_663,N_631);
nand U3720 (N_3720,N_1103,N_167);
nand U3721 (N_3721,N_1312,N_1897);
and U3722 (N_3722,N_1169,N_1227);
xor U3723 (N_3723,N_498,N_1234);
or U3724 (N_3724,N_706,N_1730);
or U3725 (N_3725,N_1437,N_855);
or U3726 (N_3726,N_1161,N_1018);
nor U3727 (N_3727,N_1139,N_118);
xnor U3728 (N_3728,N_436,N_498);
and U3729 (N_3729,N_106,N_660);
nand U3730 (N_3730,N_1972,N_188);
nor U3731 (N_3731,N_708,N_1668);
nand U3732 (N_3732,N_190,N_74);
or U3733 (N_3733,N_625,N_882);
nand U3734 (N_3734,N_1636,N_1310);
or U3735 (N_3735,N_964,N_918);
nor U3736 (N_3736,N_1172,N_550);
nand U3737 (N_3737,N_1024,N_655);
nand U3738 (N_3738,N_1176,N_1507);
nand U3739 (N_3739,N_969,N_1434);
nand U3740 (N_3740,N_1169,N_113);
nor U3741 (N_3741,N_206,N_506);
nor U3742 (N_3742,N_1443,N_1412);
nand U3743 (N_3743,N_1866,N_34);
nand U3744 (N_3744,N_342,N_1646);
nor U3745 (N_3745,N_407,N_325);
nand U3746 (N_3746,N_1304,N_1528);
and U3747 (N_3747,N_1435,N_1288);
and U3748 (N_3748,N_1578,N_1686);
nand U3749 (N_3749,N_1564,N_490);
xor U3750 (N_3750,N_382,N_1683);
nor U3751 (N_3751,N_1186,N_1454);
nor U3752 (N_3752,N_281,N_1134);
nor U3753 (N_3753,N_965,N_1670);
and U3754 (N_3754,N_1111,N_1834);
xor U3755 (N_3755,N_697,N_727);
xor U3756 (N_3756,N_1805,N_1435);
or U3757 (N_3757,N_349,N_774);
nand U3758 (N_3758,N_972,N_498);
nand U3759 (N_3759,N_176,N_1027);
or U3760 (N_3760,N_1633,N_494);
nand U3761 (N_3761,N_333,N_1906);
and U3762 (N_3762,N_1505,N_1454);
nor U3763 (N_3763,N_878,N_1973);
nor U3764 (N_3764,N_371,N_1843);
nor U3765 (N_3765,N_1893,N_1428);
nor U3766 (N_3766,N_746,N_442);
nand U3767 (N_3767,N_663,N_17);
or U3768 (N_3768,N_1889,N_1498);
nand U3769 (N_3769,N_1328,N_686);
or U3770 (N_3770,N_1542,N_835);
nor U3771 (N_3771,N_799,N_27);
and U3772 (N_3772,N_379,N_495);
nor U3773 (N_3773,N_697,N_1858);
or U3774 (N_3774,N_970,N_901);
nor U3775 (N_3775,N_652,N_193);
nor U3776 (N_3776,N_305,N_922);
nor U3777 (N_3777,N_1683,N_982);
or U3778 (N_3778,N_723,N_45);
nand U3779 (N_3779,N_529,N_1954);
and U3780 (N_3780,N_1168,N_975);
xnor U3781 (N_3781,N_1438,N_544);
or U3782 (N_3782,N_1198,N_126);
or U3783 (N_3783,N_1935,N_193);
nor U3784 (N_3784,N_1380,N_1178);
or U3785 (N_3785,N_430,N_1633);
nand U3786 (N_3786,N_582,N_1038);
nand U3787 (N_3787,N_1859,N_56);
xor U3788 (N_3788,N_626,N_1335);
nor U3789 (N_3789,N_1545,N_1664);
and U3790 (N_3790,N_1025,N_47);
or U3791 (N_3791,N_1308,N_727);
or U3792 (N_3792,N_809,N_764);
xor U3793 (N_3793,N_969,N_925);
and U3794 (N_3794,N_963,N_1175);
xor U3795 (N_3795,N_1049,N_484);
and U3796 (N_3796,N_344,N_1439);
xor U3797 (N_3797,N_354,N_858);
and U3798 (N_3798,N_1432,N_1679);
or U3799 (N_3799,N_1428,N_1626);
nand U3800 (N_3800,N_1929,N_1585);
xor U3801 (N_3801,N_1005,N_967);
nor U3802 (N_3802,N_353,N_669);
nand U3803 (N_3803,N_538,N_1851);
nor U3804 (N_3804,N_4,N_1166);
nor U3805 (N_3805,N_1645,N_1290);
nor U3806 (N_3806,N_1890,N_1119);
and U3807 (N_3807,N_1776,N_178);
and U3808 (N_3808,N_1744,N_1514);
or U3809 (N_3809,N_1312,N_261);
xor U3810 (N_3810,N_25,N_1447);
xor U3811 (N_3811,N_492,N_503);
and U3812 (N_3812,N_236,N_1488);
or U3813 (N_3813,N_645,N_1215);
nand U3814 (N_3814,N_1336,N_753);
nand U3815 (N_3815,N_823,N_968);
nor U3816 (N_3816,N_72,N_639);
or U3817 (N_3817,N_291,N_146);
xnor U3818 (N_3818,N_219,N_1975);
and U3819 (N_3819,N_547,N_1950);
xor U3820 (N_3820,N_496,N_213);
and U3821 (N_3821,N_1283,N_538);
nand U3822 (N_3822,N_331,N_565);
and U3823 (N_3823,N_1310,N_1490);
or U3824 (N_3824,N_1938,N_1337);
nor U3825 (N_3825,N_1610,N_839);
nand U3826 (N_3826,N_1303,N_381);
or U3827 (N_3827,N_1000,N_847);
nor U3828 (N_3828,N_499,N_1651);
or U3829 (N_3829,N_1650,N_271);
xnor U3830 (N_3830,N_995,N_1235);
xnor U3831 (N_3831,N_1973,N_576);
xor U3832 (N_3832,N_227,N_1306);
nor U3833 (N_3833,N_468,N_1532);
nand U3834 (N_3834,N_1546,N_1251);
nand U3835 (N_3835,N_1849,N_893);
nor U3836 (N_3836,N_1402,N_890);
xnor U3837 (N_3837,N_318,N_183);
nor U3838 (N_3838,N_1643,N_794);
and U3839 (N_3839,N_1481,N_906);
nor U3840 (N_3840,N_1182,N_1433);
xor U3841 (N_3841,N_1350,N_646);
nand U3842 (N_3842,N_1735,N_971);
nor U3843 (N_3843,N_1238,N_1912);
nor U3844 (N_3844,N_516,N_990);
and U3845 (N_3845,N_255,N_787);
nor U3846 (N_3846,N_603,N_1990);
or U3847 (N_3847,N_1099,N_630);
xor U3848 (N_3848,N_1050,N_1647);
and U3849 (N_3849,N_604,N_1844);
nor U3850 (N_3850,N_1209,N_601);
nand U3851 (N_3851,N_388,N_1937);
xor U3852 (N_3852,N_629,N_735);
xnor U3853 (N_3853,N_436,N_1414);
and U3854 (N_3854,N_1076,N_133);
xnor U3855 (N_3855,N_1724,N_627);
xor U3856 (N_3856,N_1377,N_1611);
xor U3857 (N_3857,N_1280,N_1876);
nand U3858 (N_3858,N_1585,N_1435);
and U3859 (N_3859,N_143,N_1329);
nand U3860 (N_3860,N_1421,N_1509);
nand U3861 (N_3861,N_581,N_1938);
and U3862 (N_3862,N_950,N_83);
xnor U3863 (N_3863,N_1771,N_1735);
xnor U3864 (N_3864,N_503,N_1013);
nor U3865 (N_3865,N_1553,N_557);
nor U3866 (N_3866,N_1,N_464);
xnor U3867 (N_3867,N_238,N_1166);
and U3868 (N_3868,N_931,N_970);
xor U3869 (N_3869,N_949,N_1989);
nor U3870 (N_3870,N_1592,N_1120);
xnor U3871 (N_3871,N_1523,N_1236);
and U3872 (N_3872,N_1069,N_1956);
nand U3873 (N_3873,N_361,N_1105);
and U3874 (N_3874,N_233,N_1181);
nor U3875 (N_3875,N_1042,N_596);
nor U3876 (N_3876,N_845,N_47);
xor U3877 (N_3877,N_1112,N_777);
nand U3878 (N_3878,N_930,N_1199);
or U3879 (N_3879,N_548,N_1394);
and U3880 (N_3880,N_1992,N_98);
xnor U3881 (N_3881,N_1585,N_389);
nand U3882 (N_3882,N_1445,N_1614);
or U3883 (N_3883,N_1849,N_1680);
xor U3884 (N_3884,N_1262,N_1532);
xor U3885 (N_3885,N_1613,N_990);
and U3886 (N_3886,N_776,N_223);
nor U3887 (N_3887,N_507,N_1356);
nor U3888 (N_3888,N_719,N_1795);
xnor U3889 (N_3889,N_1755,N_388);
nor U3890 (N_3890,N_1784,N_1655);
nor U3891 (N_3891,N_732,N_798);
nor U3892 (N_3892,N_1879,N_1685);
xor U3893 (N_3893,N_1762,N_66);
nand U3894 (N_3894,N_1710,N_407);
or U3895 (N_3895,N_1926,N_1660);
nand U3896 (N_3896,N_969,N_272);
xor U3897 (N_3897,N_1188,N_1169);
or U3898 (N_3898,N_740,N_599);
nand U3899 (N_3899,N_1184,N_1827);
xor U3900 (N_3900,N_491,N_1541);
xor U3901 (N_3901,N_853,N_1911);
xnor U3902 (N_3902,N_1956,N_527);
nand U3903 (N_3903,N_562,N_951);
and U3904 (N_3904,N_104,N_1910);
nor U3905 (N_3905,N_1942,N_343);
nand U3906 (N_3906,N_826,N_1754);
nor U3907 (N_3907,N_1869,N_677);
xnor U3908 (N_3908,N_1039,N_347);
nand U3909 (N_3909,N_1411,N_1463);
xor U3910 (N_3910,N_694,N_1317);
or U3911 (N_3911,N_155,N_915);
nand U3912 (N_3912,N_1675,N_294);
xor U3913 (N_3913,N_904,N_1713);
nor U3914 (N_3914,N_411,N_1714);
nand U3915 (N_3915,N_437,N_594);
and U3916 (N_3916,N_228,N_703);
and U3917 (N_3917,N_295,N_734);
and U3918 (N_3918,N_1587,N_1938);
or U3919 (N_3919,N_1931,N_948);
nand U3920 (N_3920,N_381,N_823);
xnor U3921 (N_3921,N_567,N_1144);
and U3922 (N_3922,N_1680,N_744);
xor U3923 (N_3923,N_1534,N_272);
and U3924 (N_3924,N_1542,N_1740);
nor U3925 (N_3925,N_1396,N_951);
nor U3926 (N_3926,N_1043,N_590);
nand U3927 (N_3927,N_1177,N_625);
xor U3928 (N_3928,N_596,N_1560);
or U3929 (N_3929,N_1446,N_941);
or U3930 (N_3930,N_1591,N_1127);
nor U3931 (N_3931,N_1860,N_1550);
nand U3932 (N_3932,N_1089,N_381);
or U3933 (N_3933,N_1741,N_489);
nand U3934 (N_3934,N_984,N_1350);
or U3935 (N_3935,N_1913,N_1192);
nor U3936 (N_3936,N_501,N_1378);
nand U3937 (N_3937,N_1105,N_988);
xor U3938 (N_3938,N_94,N_292);
nor U3939 (N_3939,N_1085,N_286);
xnor U3940 (N_3940,N_1118,N_1523);
xor U3941 (N_3941,N_1001,N_380);
nor U3942 (N_3942,N_357,N_620);
nand U3943 (N_3943,N_1828,N_1426);
nand U3944 (N_3944,N_33,N_59);
nand U3945 (N_3945,N_1400,N_710);
xnor U3946 (N_3946,N_1784,N_1684);
nor U3947 (N_3947,N_917,N_1150);
nor U3948 (N_3948,N_78,N_1828);
nor U3949 (N_3949,N_121,N_1676);
or U3950 (N_3950,N_892,N_516);
nor U3951 (N_3951,N_1797,N_584);
or U3952 (N_3952,N_266,N_997);
and U3953 (N_3953,N_1235,N_440);
and U3954 (N_3954,N_796,N_1161);
or U3955 (N_3955,N_872,N_1332);
or U3956 (N_3956,N_885,N_1318);
or U3957 (N_3957,N_1326,N_1733);
or U3958 (N_3958,N_417,N_334);
and U3959 (N_3959,N_1171,N_1617);
nor U3960 (N_3960,N_1697,N_189);
and U3961 (N_3961,N_1377,N_77);
nand U3962 (N_3962,N_593,N_265);
nor U3963 (N_3963,N_801,N_879);
or U3964 (N_3964,N_1106,N_466);
nand U3965 (N_3965,N_806,N_992);
xor U3966 (N_3966,N_1282,N_1012);
nor U3967 (N_3967,N_232,N_286);
or U3968 (N_3968,N_1524,N_419);
xnor U3969 (N_3969,N_1791,N_1658);
and U3970 (N_3970,N_844,N_1803);
nand U3971 (N_3971,N_256,N_1185);
nor U3972 (N_3972,N_363,N_974);
nor U3973 (N_3973,N_1337,N_985);
nor U3974 (N_3974,N_742,N_387);
and U3975 (N_3975,N_1926,N_1068);
nor U3976 (N_3976,N_843,N_1571);
nand U3977 (N_3977,N_780,N_1150);
nand U3978 (N_3978,N_1178,N_1579);
nand U3979 (N_3979,N_833,N_1131);
or U3980 (N_3980,N_1748,N_567);
or U3981 (N_3981,N_1298,N_1768);
nand U3982 (N_3982,N_760,N_294);
nor U3983 (N_3983,N_1849,N_1904);
xnor U3984 (N_3984,N_1251,N_1839);
xnor U3985 (N_3985,N_961,N_385);
or U3986 (N_3986,N_1266,N_405);
or U3987 (N_3987,N_1617,N_500);
xor U3988 (N_3988,N_1243,N_1336);
or U3989 (N_3989,N_560,N_1336);
nor U3990 (N_3990,N_319,N_113);
nor U3991 (N_3991,N_1733,N_1859);
nor U3992 (N_3992,N_398,N_40);
and U3993 (N_3993,N_1884,N_103);
xnor U3994 (N_3994,N_359,N_1371);
nor U3995 (N_3995,N_861,N_1908);
xnor U3996 (N_3996,N_1387,N_1742);
and U3997 (N_3997,N_1698,N_1191);
xnor U3998 (N_3998,N_1826,N_940);
nor U3999 (N_3999,N_701,N_1310);
nor U4000 (N_4000,N_3956,N_2166);
nor U4001 (N_4001,N_3474,N_2525);
and U4002 (N_4002,N_2480,N_3331);
nor U4003 (N_4003,N_2468,N_3872);
and U4004 (N_4004,N_3566,N_3122);
and U4005 (N_4005,N_2200,N_3778);
and U4006 (N_4006,N_2712,N_3810);
xor U4007 (N_4007,N_2957,N_3791);
xor U4008 (N_4008,N_3747,N_2120);
and U4009 (N_4009,N_3623,N_2337);
xnor U4010 (N_4010,N_2176,N_3323);
and U4011 (N_4011,N_3946,N_3183);
or U4012 (N_4012,N_3075,N_3460);
nor U4013 (N_4013,N_2377,N_3168);
nor U4014 (N_4014,N_3807,N_3248);
xor U4015 (N_4015,N_2429,N_2992);
nor U4016 (N_4016,N_2580,N_2511);
nor U4017 (N_4017,N_3702,N_3327);
nor U4018 (N_4018,N_2475,N_3280);
or U4019 (N_4019,N_2763,N_3031);
xor U4020 (N_4020,N_3079,N_3803);
nor U4021 (N_4021,N_3435,N_2430);
or U4022 (N_4022,N_2056,N_2087);
or U4023 (N_4023,N_3339,N_3355);
nand U4024 (N_4024,N_2604,N_2899);
and U4025 (N_4025,N_3948,N_2673);
xor U4026 (N_4026,N_3684,N_3061);
and U4027 (N_4027,N_3171,N_3772);
nor U4028 (N_4028,N_2578,N_2660);
or U4029 (N_4029,N_2886,N_2224);
and U4030 (N_4030,N_2452,N_3907);
xnor U4031 (N_4031,N_2782,N_2259);
nand U4032 (N_4032,N_3799,N_3535);
nand U4033 (N_4033,N_2102,N_2421);
and U4034 (N_4034,N_3935,N_3486);
or U4035 (N_4035,N_2380,N_2513);
nand U4036 (N_4036,N_2690,N_3551);
or U4037 (N_4037,N_2705,N_3133);
and U4038 (N_4038,N_3856,N_2472);
nor U4039 (N_4039,N_2461,N_3688);
nor U4040 (N_4040,N_3932,N_2512);
or U4041 (N_4041,N_3001,N_3796);
nor U4042 (N_4042,N_2314,N_3552);
nor U4043 (N_4043,N_3913,N_2347);
nor U4044 (N_4044,N_2987,N_2010);
xnor U4045 (N_4045,N_3157,N_2562);
or U4046 (N_4046,N_3569,N_2964);
nand U4047 (N_4047,N_2264,N_2691);
nor U4048 (N_4048,N_3720,N_2518);
or U4049 (N_4049,N_2789,N_2440);
or U4050 (N_4050,N_3522,N_3729);
xor U4051 (N_4051,N_3274,N_3124);
xnor U4052 (N_4052,N_2876,N_3144);
nor U4053 (N_4053,N_3230,N_3180);
nor U4054 (N_4054,N_3104,N_3528);
xor U4055 (N_4055,N_3867,N_3563);
nor U4056 (N_4056,N_3637,N_3295);
nand U4057 (N_4057,N_2679,N_3651);
and U4058 (N_4058,N_2640,N_3457);
nor U4059 (N_4059,N_2397,N_3325);
and U4060 (N_4060,N_3193,N_2569);
and U4061 (N_4061,N_2136,N_3638);
nor U4062 (N_4062,N_3223,N_2859);
and U4063 (N_4063,N_2301,N_2055);
or U4064 (N_4064,N_2893,N_3483);
nor U4065 (N_4065,N_2069,N_2365);
nand U4066 (N_4066,N_3080,N_2875);
nor U4067 (N_4067,N_2497,N_3661);
nor U4068 (N_4068,N_3046,N_3806);
nand U4069 (N_4069,N_2422,N_2496);
nand U4070 (N_4070,N_3829,N_2607);
or U4071 (N_4071,N_3613,N_2208);
and U4072 (N_4072,N_2379,N_3618);
and U4073 (N_4073,N_2822,N_2624);
xnor U4074 (N_4074,N_2650,N_2283);
xor U4075 (N_4075,N_2130,N_2537);
and U4076 (N_4076,N_3653,N_2535);
nor U4077 (N_4077,N_3650,N_2097);
and U4078 (N_4078,N_2317,N_2672);
nand U4079 (N_4079,N_3070,N_2107);
nor U4080 (N_4080,N_3681,N_3523);
and U4081 (N_4081,N_3822,N_3469);
nand U4082 (N_4082,N_2682,N_3383);
or U4083 (N_4083,N_2318,N_3450);
xor U4084 (N_4084,N_2404,N_3812);
or U4085 (N_4085,N_2601,N_2326);
and U4086 (N_4086,N_3683,N_3699);
nand U4087 (N_4087,N_3313,N_2570);
nor U4088 (N_4088,N_3240,N_2958);
nand U4089 (N_4089,N_2443,N_2500);
nor U4090 (N_4090,N_2156,N_3800);
or U4091 (N_4091,N_3801,N_2129);
xnor U4092 (N_4092,N_3758,N_2841);
xor U4093 (N_4093,N_3804,N_3925);
nand U4094 (N_4094,N_3555,N_3453);
nand U4095 (N_4095,N_3781,N_3832);
or U4096 (N_4096,N_3814,N_3251);
nor U4097 (N_4097,N_2204,N_3979);
and U4098 (N_4098,N_3545,N_3089);
nand U4099 (N_4099,N_2192,N_2025);
or U4100 (N_4100,N_2171,N_2944);
nor U4101 (N_4101,N_3304,N_2199);
and U4102 (N_4102,N_2993,N_2148);
or U4103 (N_4103,N_2004,N_2113);
nand U4104 (N_4104,N_2868,N_3348);
xor U4105 (N_4105,N_2565,N_2117);
xor U4106 (N_4106,N_3685,N_2692);
or U4107 (N_4107,N_3918,N_2592);
or U4108 (N_4108,N_2213,N_3477);
or U4109 (N_4109,N_3950,N_2403);
nor U4110 (N_4110,N_3021,N_3336);
and U4111 (N_4111,N_2392,N_2072);
or U4112 (N_4112,N_2357,N_3252);
or U4113 (N_4113,N_3045,N_3838);
nand U4114 (N_4114,N_3238,N_2433);
and U4115 (N_4115,N_3367,N_3161);
xnor U4116 (N_4116,N_3073,N_2411);
xnor U4117 (N_4117,N_2487,N_2424);
xnor U4118 (N_4118,N_2641,N_3817);
and U4119 (N_4119,N_3578,N_3627);
nand U4120 (N_4120,N_2294,N_2118);
xnor U4121 (N_4121,N_2867,N_2054);
and U4122 (N_4122,N_2310,N_2917);
or U4123 (N_4123,N_3141,N_2967);
nand U4124 (N_4124,N_3105,N_2343);
or U4125 (N_4125,N_2855,N_3287);
or U4126 (N_4126,N_2796,N_3657);
and U4127 (N_4127,N_2367,N_2638);
and U4128 (N_4128,N_2378,N_2460);
nand U4129 (N_4129,N_2559,N_3983);
nand U4130 (N_4130,N_3060,N_3356);
nor U4131 (N_4131,N_2646,N_2664);
and U4132 (N_4132,N_2193,N_2390);
and U4133 (N_4133,N_2329,N_3573);
xnor U4134 (N_4134,N_3710,N_3150);
and U4135 (N_4135,N_3920,N_3534);
or U4136 (N_4136,N_2866,N_3874);
and U4137 (N_4137,N_3707,N_2888);
nand U4138 (N_4138,N_2990,N_3004);
or U4139 (N_4139,N_3784,N_2544);
nand U4140 (N_4140,N_2962,N_2619);
nor U4141 (N_4141,N_3322,N_2162);
xnor U4142 (N_4142,N_3694,N_3571);
and U4143 (N_4143,N_2889,N_2585);
or U4144 (N_4144,N_3062,N_2246);
xor U4145 (N_4145,N_2319,N_3895);
or U4146 (N_4146,N_2582,N_2252);
nand U4147 (N_4147,N_2504,N_2188);
nor U4148 (N_4148,N_2140,N_2805);
and U4149 (N_4149,N_3439,N_2980);
and U4150 (N_4150,N_2564,N_3236);
xor U4151 (N_4151,N_2432,N_2187);
nand U4152 (N_4152,N_3420,N_3362);
nand U4153 (N_4153,N_3825,N_3713);
nand U4154 (N_4154,N_2738,N_3186);
nand U4155 (N_4155,N_2829,N_2265);
nor U4156 (N_4156,N_2082,N_2158);
or U4157 (N_4157,N_3283,N_2852);
or U4158 (N_4158,N_2297,N_3628);
or U4159 (N_4159,N_2960,N_2495);
and U4160 (N_4160,N_2744,N_3057);
and U4161 (N_4161,N_2183,N_2799);
nor U4162 (N_4162,N_2230,N_2747);
or U4163 (N_4163,N_2393,N_2776);
xor U4164 (N_4164,N_3140,N_3445);
nor U4165 (N_4165,N_3776,N_3992);
nand U4166 (N_4166,N_3278,N_2579);
xnor U4167 (N_4167,N_3518,N_3320);
and U4168 (N_4168,N_2645,N_2567);
or U4169 (N_4169,N_3083,N_2181);
nor U4170 (N_4170,N_3584,N_2292);
nand U4171 (N_4171,N_2320,N_3887);
or U4172 (N_4172,N_3225,N_3691);
or U4173 (N_4173,N_3763,N_3098);
or U4174 (N_4174,N_2689,N_3388);
xor U4175 (N_4175,N_3466,N_3052);
or U4176 (N_4176,N_2023,N_3754);
and U4177 (N_4177,N_3939,N_3705);
and U4178 (N_4178,N_3868,N_3769);
nand U4179 (N_4179,N_2736,N_3904);
nor U4180 (N_4180,N_2872,N_2700);
nand U4181 (N_4181,N_2746,N_3660);
nor U4182 (N_4182,N_2651,N_2434);
or U4183 (N_4183,N_2869,N_2172);
and U4184 (N_4184,N_3241,N_2989);
and U4185 (N_4185,N_3484,N_3505);
xnor U4186 (N_4186,N_3481,N_2066);
or U4187 (N_4187,N_2322,N_2669);
or U4188 (N_4188,N_2469,N_2795);
nor U4189 (N_4189,N_3167,N_2356);
or U4190 (N_4190,N_3464,N_2416);
nor U4191 (N_4191,N_2820,N_3659);
nand U4192 (N_4192,N_3063,N_3254);
nor U4193 (N_4193,N_2814,N_2998);
and U4194 (N_4194,N_3853,N_3300);
nand U4195 (N_4195,N_2413,N_2626);
or U4196 (N_4196,N_2808,N_2031);
xor U4197 (N_4197,N_3368,N_2146);
nand U4198 (N_4198,N_3081,N_2182);
nand U4199 (N_4199,N_3988,N_2750);
xnor U4200 (N_4200,N_3843,N_3415);
nor U4201 (N_4201,N_3123,N_2800);
nand U4202 (N_4202,N_3517,N_2375);
nand U4203 (N_4203,N_2126,N_3841);
xor U4204 (N_4204,N_2846,N_3148);
xor U4205 (N_4205,N_2105,N_2685);
nor U4206 (N_4206,N_3974,N_2289);
nor U4207 (N_4207,N_3390,N_3839);
nor U4208 (N_4208,N_2906,N_3159);
xor U4209 (N_4209,N_2395,N_3125);
nor U4210 (N_4210,N_2211,N_3101);
or U4211 (N_4211,N_2662,N_2271);
nand U4212 (N_4212,N_2787,N_3110);
nand U4213 (N_4213,N_3218,N_3883);
nand U4214 (N_4214,N_2458,N_3201);
and U4215 (N_4215,N_2353,N_3302);
xnor U4216 (N_4216,N_2332,N_2725);
and U4217 (N_4217,N_2788,N_3471);
or U4218 (N_4218,N_3858,N_3396);
nor U4219 (N_4219,N_2272,N_2729);
nand U4220 (N_4220,N_2355,N_3876);
and U4221 (N_4221,N_2951,N_3384);
nand U4222 (N_4222,N_2721,N_3014);
or U4223 (N_4223,N_2389,N_2410);
or U4224 (N_4224,N_3177,N_2697);
and U4225 (N_4225,N_2280,N_2642);
xnor U4226 (N_4226,N_3908,N_2704);
nor U4227 (N_4227,N_2342,N_3343);
and U4228 (N_4228,N_3862,N_3020);
and U4229 (N_4229,N_2111,N_2760);
or U4230 (N_4230,N_3345,N_2479);
or U4231 (N_4231,N_3968,N_3402);
nand U4232 (N_4232,N_2802,N_2086);
nor U4233 (N_4233,N_3850,N_2046);
and U4234 (N_4234,N_3109,N_3427);
xnor U4235 (N_4235,N_2236,N_2901);
or U4236 (N_4236,N_2401,N_2929);
or U4237 (N_4237,N_2628,N_2359);
nor U4238 (N_4238,N_2436,N_2765);
and U4239 (N_4239,N_3590,N_3941);
nand U4240 (N_4240,N_3130,N_2457);
or U4241 (N_4241,N_3202,N_2762);
xnor U4242 (N_4242,N_3069,N_2915);
nand U4243 (N_4243,N_2175,N_2683);
and U4244 (N_4244,N_3996,N_3525);
and U4245 (N_4245,N_3745,N_2939);
or U4246 (N_4246,N_2470,N_3126);
nand U4247 (N_4247,N_3565,N_3050);
and U4248 (N_4248,N_2414,N_3680);
nand U4249 (N_4249,N_2234,N_2935);
or U4250 (N_4250,N_3370,N_2291);
or U4251 (N_4251,N_3949,N_2445);
and U4252 (N_4252,N_3764,N_2128);
nor U4253 (N_4253,N_2005,N_2474);
nand U4254 (N_4254,N_3991,N_3044);
nor U4255 (N_4255,N_3154,N_3833);
and U4256 (N_4256,N_3330,N_3798);
or U4257 (N_4257,N_3733,N_3693);
and U4258 (N_4258,N_3042,N_3896);
and U4259 (N_4259,N_2834,N_2110);
xor U4260 (N_4260,N_2828,N_3993);
nor U4261 (N_4261,N_2016,N_2144);
xnor U4262 (N_4262,N_3615,N_3443);
and U4263 (N_4263,N_2139,N_3496);
nor U4264 (N_4264,N_3553,N_2299);
xor U4265 (N_4265,N_2221,N_3340);
or U4266 (N_4266,N_2084,N_3478);
xnor U4267 (N_4267,N_2620,N_3587);
and U4268 (N_4268,N_2801,N_3369);
and U4269 (N_4269,N_3977,N_3994);
nand U4270 (N_4270,N_3100,N_2473);
nand U4271 (N_4271,N_2398,N_2756);
nand U4272 (N_4272,N_3506,N_2486);
nor U4273 (N_4273,N_3281,N_3138);
nor U4274 (N_4274,N_3601,N_3092);
nand U4275 (N_4275,N_2058,N_3631);
xor U4276 (N_4276,N_2463,N_3306);
nand U4277 (N_4277,N_3146,N_3787);
xnor U4278 (N_4278,N_3214,N_2415);
nor U4279 (N_4279,N_3107,N_3371);
nand U4280 (N_4280,N_3735,N_2608);
nand U4281 (N_4281,N_2370,N_2880);
or U4282 (N_4282,N_3134,N_3873);
xor U4283 (N_4283,N_2373,N_3570);
or U4284 (N_4284,N_3115,N_2573);
and U4285 (N_4285,N_2405,N_2354);
nand U4286 (N_4286,N_3239,N_2268);
xnor U4287 (N_4287,N_2654,N_2761);
or U4288 (N_4288,N_2777,N_3824);
nand U4289 (N_4289,N_2083,N_3498);
nor U4290 (N_4290,N_3774,N_2062);
nor U4291 (N_4291,N_3392,N_3197);
xnor U4292 (N_4292,N_2686,N_2919);
nand U4293 (N_4293,N_3231,N_2052);
or U4294 (N_4294,N_2165,N_3645);
xnor U4295 (N_4295,N_2783,N_3562);
or U4296 (N_4296,N_2591,N_2648);
or U4297 (N_4297,N_3624,N_3863);
nor U4298 (N_4298,N_3931,N_2109);
nand U4299 (N_4299,N_3507,N_3112);
nor U4300 (N_4300,N_2767,N_2595);
or U4301 (N_4301,N_3748,N_2447);
and U4302 (N_4302,N_3921,N_2719);
xor U4303 (N_4303,N_3775,N_2657);
nor U4304 (N_4304,N_3458,N_2138);
and U4305 (N_4305,N_2132,N_2784);
nor U4306 (N_4306,N_3164,N_3906);
and U4307 (N_4307,N_3970,N_3654);
and U4308 (N_4308,N_3255,N_3944);
nor U4309 (N_4309,N_2349,N_3350);
xor U4310 (N_4310,N_2668,N_3023);
nor U4311 (N_4311,N_2041,N_2770);
nand U4312 (N_4312,N_2376,N_3451);
or U4313 (N_4313,N_3119,N_3972);
nor U4314 (N_4314,N_3997,N_3398);
nor U4315 (N_4315,N_2890,N_3761);
nor U4316 (N_4316,N_2164,N_3744);
and U4317 (N_4317,N_3952,N_2293);
nand U4318 (N_4318,N_3830,N_3890);
or U4319 (N_4319,N_3664,N_2262);
nand U4320 (N_4320,N_2364,N_2593);
nor U4321 (N_4321,N_2185,N_2602);
nand U4322 (N_4322,N_2816,N_3773);
xor U4323 (N_4323,N_3632,N_3059);
and U4324 (N_4324,N_2617,N_2209);
or U4325 (N_4325,N_3634,N_2837);
nor U4326 (N_4326,N_2091,N_3916);
and U4327 (N_4327,N_2178,N_2904);
xnor U4328 (N_4328,N_2918,N_3985);
nand U4329 (N_4329,N_3513,N_2625);
or U4330 (N_4330,N_2838,N_3291);
xnor U4331 (N_4331,N_2644,N_2286);
or U4332 (N_4332,N_3099,N_3431);
nor U4333 (N_4333,N_2194,N_2121);
xnor U4334 (N_4334,N_2873,N_2926);
nor U4335 (N_4335,N_3329,N_3759);
xnor U4336 (N_4336,N_3208,N_3786);
or U4337 (N_4337,N_2674,N_2002);
nand U4338 (N_4338,N_3421,N_2240);
xor U4339 (N_4339,N_3642,N_2634);
xor U4340 (N_4340,N_2726,N_3011);
and U4341 (N_4341,N_3746,N_3558);
xor U4342 (N_4342,N_2335,N_2968);
or U4343 (N_4343,N_2649,N_2001);
and U4344 (N_4344,N_3256,N_2145);
xnor U4345 (N_4345,N_3797,N_3554);
nand U4346 (N_4346,N_3725,N_2163);
xor U4347 (N_4347,N_3078,N_3181);
xor U4348 (N_4348,N_2698,N_2881);
and U4349 (N_4349,N_2437,N_2551);
and U4350 (N_4350,N_3065,N_3263);
or U4351 (N_4351,N_2557,N_2276);
xor U4352 (N_4352,N_3228,N_3588);
or U4353 (N_4353,N_2597,N_3428);
nand U4354 (N_4354,N_3179,N_3296);
xnor U4355 (N_4355,N_3527,N_3891);
xor U4356 (N_4356,N_2363,N_2231);
nand U4357 (N_4357,N_3819,N_2790);
nand U4358 (N_4358,N_3538,N_3844);
xnor U4359 (N_4359,N_3607,N_2854);
or U4360 (N_4360,N_3393,N_2879);
xnor U4361 (N_4361,N_3465,N_2722);
and U4362 (N_4362,N_3273,N_3782);
xnor U4363 (N_4363,N_2774,N_2387);
nand U4364 (N_4364,N_2715,N_3847);
nand U4365 (N_4365,N_2532,N_3185);
nand U4366 (N_4366,N_2833,N_3227);
nor U4367 (N_4367,N_2924,N_2089);
nor U4368 (N_4368,N_2142,N_3012);
nand U4369 (N_4369,N_2362,N_3963);
or U4370 (N_4370,N_3813,N_3840);
xnor U4371 (N_4371,N_3630,N_2298);
xnor U4372 (N_4372,N_2008,N_2530);
xnor U4373 (N_4373,N_2941,N_2227);
nor U4374 (N_4374,N_3793,N_2134);
nand U4375 (N_4375,N_2516,N_3409);
nand U4376 (N_4376,N_2863,N_3462);
and U4377 (N_4377,N_2603,N_2985);
or U4378 (N_4378,N_3172,N_3203);
xnor U4379 (N_4379,N_2125,N_2666);
or U4380 (N_4380,N_3372,N_2542);
xnor U4381 (N_4381,N_3220,N_3307);
or U4382 (N_4382,N_2212,N_3404);
or U4383 (N_4383,N_3815,N_2823);
or U4384 (N_4384,N_2499,N_3491);
and U4385 (N_4385,N_2489,N_3332);
or U4386 (N_4386,N_2523,N_2366);
or U4387 (N_4387,N_2971,N_3837);
and U4388 (N_4388,N_3173,N_3411);
nand U4389 (N_4389,N_3497,N_3901);
and U4390 (N_4390,N_3299,N_2707);
and U4391 (N_4391,N_2334,N_2214);
xnor U4392 (N_4392,N_2610,N_3048);
nor U4393 (N_4393,N_3442,N_2826);
nor U4394 (N_4394,N_2279,N_3893);
and U4395 (N_4395,N_2151,N_2711);
and U4396 (N_4396,N_2201,N_3543);
or U4397 (N_4397,N_2870,N_2179);
or U4398 (N_4398,N_3947,N_2892);
nor U4399 (N_4399,N_3902,N_3679);
xnor U4400 (N_4400,N_3335,N_2534);
nand U4401 (N_4401,N_3738,N_2940);
and U4402 (N_4402,N_3068,N_3721);
nor U4403 (N_4403,N_2174,N_3995);
nand U4404 (N_4404,N_2247,N_2581);
and U4405 (N_4405,N_3594,N_2543);
or U4406 (N_4406,N_2333,N_2587);
or U4407 (N_4407,N_2385,N_2028);
nand U4408 (N_4408,N_2563,N_2312);
or U4409 (N_4409,N_2029,N_3221);
nand U4410 (N_4410,N_3536,N_3544);
or U4411 (N_4411,N_2775,N_2999);
xor U4412 (N_4412,N_3303,N_3834);
nor U4413 (N_4413,N_3091,N_3399);
xnor U4414 (N_4414,N_2572,N_3516);
nand U4415 (N_4415,N_2652,N_2583);
xnor U4416 (N_4416,N_3285,N_3889);
and U4417 (N_4417,N_3811,N_2850);
and U4418 (N_4418,N_3174,N_3673);
nand U4419 (N_4419,N_2481,N_3722);
nor U4420 (N_4420,N_2517,N_2160);
xor U4421 (N_4421,N_3187,N_2408);
and U4422 (N_4422,N_2346,N_2241);
or U4423 (N_4423,N_3524,N_2059);
nor U4424 (N_4424,N_2561,N_2060);
nand U4425 (N_4425,N_3262,N_2013);
or U4426 (N_4426,N_2428,N_3264);
or U4427 (N_4427,N_3253,N_2900);
and U4428 (N_4428,N_3156,N_2623);
xor U4429 (N_4429,N_2643,N_3490);
and U4430 (N_4430,N_3040,N_3526);
xnor U4431 (N_4431,N_3200,N_2465);
and U4432 (N_4432,N_3789,N_2157);
or U4433 (N_4433,N_2556,N_2042);
nand U4434 (N_4434,N_3196,N_3696);
xor U4435 (N_4435,N_3576,N_2456);
and U4436 (N_4436,N_2027,N_3266);
or U4437 (N_4437,N_2155,N_2785);
or U4438 (N_4438,N_3492,N_2615);
or U4439 (N_4439,N_3047,N_2442);
or U4440 (N_4440,N_3606,N_2663);
xor U4441 (N_4441,N_3321,N_3459);
and U4442 (N_4442,N_2313,N_3053);
xnor U4443 (N_4443,N_3515,N_2249);
nand U4444 (N_4444,N_2665,N_2217);
xor U4445 (N_4445,N_2032,N_3940);
and U4446 (N_4446,N_3717,N_2521);
nor U4447 (N_4447,N_2418,N_3475);
nor U4448 (N_4448,N_3877,N_3358);
and U4449 (N_4449,N_2520,N_3127);
xnor U4450 (N_4450,N_3347,N_2019);
xnor U4451 (N_4451,N_2596,N_3644);
or U4452 (N_4452,N_3919,N_3363);
nand U4453 (N_4453,N_2051,N_2753);
and U4454 (N_4454,N_3743,N_2325);
nand U4455 (N_4455,N_2441,N_2483);
or U4456 (N_4456,N_2969,N_3885);
xor U4457 (N_4457,N_3512,N_3851);
nand U4458 (N_4458,N_2494,N_3360);
or U4459 (N_4459,N_3301,N_3088);
xor U4460 (N_4460,N_2858,N_2159);
xor U4461 (N_4461,N_3217,N_3547);
nor U4462 (N_4462,N_2963,N_3394);
xnor U4463 (N_4463,N_2733,N_3387);
xor U4464 (N_4464,N_3911,N_2553);
nand U4465 (N_4465,N_2505,N_3767);
or U4466 (N_4466,N_2186,N_3749);
nand U4467 (N_4467,N_3500,N_2050);
and U4468 (N_4468,N_2598,N_2701);
nor U4469 (N_4469,N_3783,N_2409);
xor U4470 (N_4470,N_2764,N_3636);
nor U4471 (N_4471,N_2577,N_2073);
and U4472 (N_4472,N_2267,N_3027);
or U4473 (N_4473,N_3085,N_3831);
and U4474 (N_4474,N_3731,N_3842);
nor U4475 (N_4475,N_3647,N_2937);
or U4476 (N_4476,N_2621,N_3113);
nor U4477 (N_4477,N_3448,N_3412);
and U4478 (N_4478,N_3090,N_3604);
nor U4479 (N_4479,N_2629,N_2566);
nand U4480 (N_4480,N_3884,N_3617);
or U4481 (N_4481,N_2902,N_2720);
xor U4482 (N_4482,N_2636,N_3675);
nand U4483 (N_4483,N_3656,N_3629);
or U4484 (N_4484,N_2527,N_3407);
xnor U4485 (N_4485,N_2897,N_2541);
nor U4486 (N_4486,N_2400,N_2104);
xnor U4487 (N_4487,N_2862,N_3310);
nand U4488 (N_4488,N_3998,N_2426);
and U4489 (N_4489,N_2751,N_3521);
xor U4490 (N_4490,N_3700,N_2694);
xor U4491 (N_4491,N_3821,N_3087);
xor U4492 (N_4492,N_2316,N_3926);
or U4493 (N_4493,N_3456,N_3597);
or U4494 (N_4494,N_3750,N_2269);
and U4495 (N_4495,N_3211,N_3184);
or U4496 (N_4496,N_2678,N_2945);
nor U4497 (N_4497,N_3976,N_3805);
or U4498 (N_4498,N_2954,N_3724);
nand U4499 (N_4499,N_3029,N_3910);
nand U4500 (N_4500,N_2284,N_2925);
nor U4501 (N_4501,N_3595,N_2718);
and U4502 (N_4502,N_3564,N_2498);
nand U4503 (N_4503,N_3643,N_2835);
and U4504 (N_4504,N_3086,N_2003);
nand U4505 (N_4505,N_2514,N_3753);
nor U4506 (N_4506,N_3620,N_3698);
or U4507 (N_4507,N_3441,N_3641);
xnor U4508 (N_4508,N_3583,N_2381);
or U4509 (N_4509,N_2821,N_3788);
nor U4510 (N_4510,N_3007,N_3894);
and U4511 (N_4511,N_3377,N_3690);
nand U4512 (N_4512,N_3957,N_2079);
xnor U4513 (N_4513,N_3210,N_3317);
or U4514 (N_4514,N_2519,N_3792);
xnor U4515 (N_4515,N_2180,N_3603);
nor U4516 (N_4516,N_3019,N_2482);
nor U4517 (N_4517,N_3132,N_3734);
nor U4518 (N_4518,N_3485,N_2396);
and U4519 (N_4519,N_2955,N_3959);
and U4520 (N_4520,N_2388,N_2898);
xnor U4521 (N_4521,N_2256,N_2454);
and U4522 (N_4522,N_3324,N_2490);
or U4523 (N_4523,N_3880,N_2716);
and U4524 (N_4524,N_3349,N_2907);
xnor U4525 (N_4525,N_2861,N_3927);
or U4526 (N_4526,N_2484,N_2748);
xnor U4527 (N_4527,N_3116,N_2938);
and U4528 (N_4528,N_3229,N_2270);
xnor U4529 (N_4529,N_2245,N_2806);
nand U4530 (N_4530,N_3933,N_2933);
nor U4531 (N_4531,N_2832,N_2606);
xor U4532 (N_4532,N_2986,N_3082);
xor U4533 (N_4533,N_2994,N_3226);
xnor U4534 (N_4534,N_3692,N_3808);
and U4535 (N_4535,N_3243,N_3076);
xor U4536 (N_4536,N_3344,N_3102);
xor U4537 (N_4537,N_3556,N_2037);
xor U4538 (N_4538,N_2916,N_3289);
or U4539 (N_4539,N_3000,N_2143);
or U4540 (N_4540,N_3723,N_2884);
xor U4541 (N_4541,N_3446,N_2202);
xor U4542 (N_4542,N_3479,N_3726);
nor U4543 (N_4543,N_3034,N_3577);
or U4544 (N_4544,N_2419,N_2189);
and U4545 (N_4545,N_3426,N_2786);
xnor U4546 (N_4546,N_2827,N_2550);
nand U4547 (N_4547,N_3865,N_3209);
and U4548 (N_4548,N_2708,N_2950);
nor U4549 (N_4549,N_2818,N_3592);
nor U4550 (N_4550,N_2450,N_2809);
nor U4551 (N_4551,N_2399,N_3117);
nor U4552 (N_4552,N_2444,N_2402);
xor U4553 (N_4553,N_3279,N_3857);
xor U4554 (N_4554,N_3328,N_2030);
nor U4555 (N_4555,N_3909,N_3149);
xnor U4556 (N_4556,N_3869,N_2681);
nand U4557 (N_4557,N_2740,N_2865);
xor U4558 (N_4558,N_2943,N_2344);
nand U4559 (N_4559,N_3669,N_2492);
nor U4560 (N_4560,N_2242,N_3771);
and U4561 (N_4561,N_2759,N_3682);
xor U4562 (N_4562,N_2632,N_2119);
nor U4563 (N_4563,N_3438,N_2921);
or U4564 (N_4564,N_3151,N_2571);
or U4565 (N_4565,N_3128,N_2699);
nand U4566 (N_4566,N_2195,N_3224);
and U4567 (N_4567,N_3338,N_3938);
xor U4568 (N_4568,N_2425,N_2198);
xor U4569 (N_4569,N_2435,N_3548);
xnor U4570 (N_4570,N_2020,N_3013);
and U4571 (N_4571,N_2693,N_3039);
nand U4572 (N_4572,N_2406,N_3129);
or U4573 (N_4573,N_2842,N_3520);
and U4574 (N_4574,N_2257,N_2609);
nand U4575 (N_4575,N_2732,N_2339);
nand U4576 (N_4576,N_2772,N_2154);
nand U4577 (N_4577,N_2077,N_3987);
and U4578 (N_4578,N_3695,N_3504);
xor U4579 (N_4579,N_2009,N_2305);
nand U4580 (N_4580,N_3309,N_3945);
and U4581 (N_4581,N_3250,N_2948);
xor U4582 (N_4582,N_2647,N_2982);
xnor U4583 (N_4583,N_3864,N_2350);
nand U4584 (N_4584,N_3602,N_3621);
and U4585 (N_4585,N_2878,N_3716);
nand U4586 (N_4586,N_3975,N_3242);
nor U4587 (N_4587,N_3581,N_3882);
nor U4588 (N_4588,N_3008,N_3414);
nand U4589 (N_4589,N_2124,N_2067);
nor U4590 (N_4590,N_3511,N_3598);
and U4591 (N_4591,N_3395,N_3108);
xnor U4592 (N_4592,N_3403,N_3574);
and U4593 (N_4593,N_3752,N_2309);
nand U4594 (N_4594,N_3888,N_3121);
and U4595 (N_4595,N_3028,N_3249);
or U4596 (N_4596,N_2035,N_2047);
and U4597 (N_4597,N_2049,N_2560);
nor U4598 (N_4598,N_3493,N_3600);
xnor U4599 (N_4599,N_3071,N_2244);
xor U4600 (N_4600,N_3828,N_2033);
xnor U4601 (N_4601,N_3417,N_3142);
and U4602 (N_4602,N_2768,N_3903);
xnor U4603 (N_4603,N_3378,N_3286);
nor U4604 (N_4604,N_2627,N_2090);
or U4605 (N_4605,N_3914,N_2478);
and U4606 (N_4606,N_3591,N_3826);
or U4607 (N_4607,N_3560,N_3986);
nand U4608 (N_4608,N_2341,N_2285);
and U4609 (N_4609,N_2044,N_3561);
and U4610 (N_4610,N_3319,N_3364);
xnor U4611 (N_4611,N_2459,N_2321);
or U4612 (N_4612,N_2345,N_3646);
or U4613 (N_4613,N_2228,N_2477);
nand U4614 (N_4614,N_2684,N_2758);
nor U4615 (N_4615,N_3870,N_3686);
and U4616 (N_4616,N_2065,N_2766);
and U4617 (N_4617,N_3163,N_3018);
or U4618 (N_4618,N_2196,N_3147);
or U4619 (N_4619,N_2169,N_2757);
or U4620 (N_4620,N_2824,N_3418);
and U4621 (N_4621,N_3715,N_2503);
xor U4622 (N_4622,N_2966,N_3670);
nor U4623 (N_4623,N_2446,N_2448);
or U4624 (N_4624,N_3709,N_3971);
or U4625 (N_4625,N_3640,N_3990);
and U4626 (N_4626,N_2351,N_2161);
nor U4627 (N_4627,N_3015,N_2811);
or U4628 (N_4628,N_3182,N_2914);
and U4629 (N_4629,N_2840,N_2730);
and U4630 (N_4630,N_2754,N_2100);
or U4631 (N_4631,N_3097,N_3703);
nand U4632 (N_4632,N_3381,N_3405);
nand U4633 (N_4633,N_3244,N_3294);
nand U4634 (N_4634,N_2427,N_3756);
nand U4635 (N_4635,N_2895,N_3917);
nor U4636 (N_4636,N_2501,N_2290);
or U4637 (N_4637,N_2778,N_3589);
nor U4638 (N_4638,N_2466,N_3290);
and U4639 (N_4639,N_3003,N_3848);
or U4640 (N_4640,N_3265,N_2614);
nand U4641 (N_4641,N_3429,N_3480);
nand U4642 (N_4642,N_2896,N_2203);
nor U4643 (N_4643,N_3373,N_2015);
and U4644 (N_4644,N_2825,N_2857);
or U4645 (N_4645,N_2912,N_2702);
or U4646 (N_4646,N_3234,N_3433);
nand U4647 (N_4647,N_2300,N_3260);
nor U4648 (N_4648,N_3488,N_3658);
nand U4649 (N_4649,N_2887,N_3540);
or U4650 (N_4650,N_3905,N_2755);
and U4651 (N_4651,N_2845,N_3035);
nor U4652 (N_4652,N_3024,N_3768);
nor U4653 (N_4653,N_2622,N_3755);
nand U4654 (N_4654,N_2853,N_2239);
and U4655 (N_4655,N_2836,N_3030);
or U4656 (N_4656,N_2605,N_2152);
nor U4657 (N_4657,N_3158,N_3989);
and U4658 (N_4658,N_3687,N_3470);
nor U4659 (N_4659,N_2979,N_2656);
nor U4660 (N_4660,N_2703,N_3314);
or U4661 (N_4661,N_3472,N_3131);
or U4662 (N_4662,N_2803,N_3619);
nor U4663 (N_4663,N_2210,N_3084);
or U4664 (N_4664,N_3790,N_2324);
nand U4665 (N_4665,N_2141,N_2168);
nand U4666 (N_4666,N_2696,N_3166);
or U4667 (N_4667,N_2507,N_3191);
nor U4668 (N_4668,N_2653,N_2229);
and U4669 (N_4669,N_2115,N_2536);
nand U4670 (N_4670,N_3096,N_3232);
xor U4671 (N_4671,N_3155,N_3845);
nand U4672 (N_4672,N_2812,N_2540);
xor U4673 (N_4673,N_2070,N_2936);
or U4674 (N_4674,N_3452,N_3106);
nor U4675 (N_4675,N_3354,N_2981);
nand U4676 (N_4676,N_3635,N_3333);
nor U4677 (N_4677,N_3579,N_3192);
and U4678 (N_4678,N_3677,N_2423);
nand U4679 (N_4679,N_3284,N_2233);
or U4680 (N_4680,N_3365,N_3499);
xor U4681 (N_4681,N_3633,N_3982);
nand U4682 (N_4682,N_2771,N_2659);
and U4683 (N_4683,N_2903,N_2476);
and U4684 (N_4684,N_3568,N_3002);
xnor U4685 (N_4685,N_2531,N_2661);
xnor U4686 (N_4686,N_2819,N_2123);
nor U4687 (N_4687,N_3671,N_2191);
or U4688 (N_4688,N_3235,N_2057);
and U4689 (N_4689,N_2630,N_2991);
and U4690 (N_4690,N_2095,N_3765);
xor U4691 (N_4691,N_3835,N_2338);
and U4692 (N_4692,N_3397,N_3258);
xor U4693 (N_4693,N_2167,N_2555);
nand U4694 (N_4694,N_2101,N_2589);
and U4695 (N_4695,N_3430,N_2099);
nor U4696 (N_4696,N_3999,N_3648);
or U4697 (N_4697,N_2374,N_3962);
nor U4698 (N_4698,N_2737,N_3190);
or U4699 (N_4699,N_2149,N_3550);
xor U4700 (N_4700,N_2509,N_2677);
nand U4701 (N_4701,N_3213,N_2358);
and U4702 (N_4702,N_3467,N_2014);
nor U4703 (N_4703,N_3929,N_2080);
nor U4704 (N_4704,N_2680,N_3881);
and U4705 (N_4705,N_3559,N_3608);
nor U4706 (N_4706,N_2538,N_2885);
nor U4707 (N_4707,N_2844,N_3215);
nor U4708 (N_4708,N_3697,N_2548);
xnor U4709 (N_4709,N_2048,N_3233);
or U4710 (N_4710,N_2773,N_3032);
and U4711 (N_4711,N_2064,N_2170);
and U4712 (N_4712,N_3170,N_2219);
or U4713 (N_4713,N_2849,N_2956);
xor U4714 (N_4714,N_2909,N_2611);
or U4715 (N_4715,N_3305,N_3585);
and U4716 (N_4716,N_2830,N_2391);
and U4717 (N_4717,N_2250,N_3964);
nor U4718 (N_4718,N_3337,N_2586);
nand U4719 (N_4719,N_3878,N_2094);
xor U4720 (N_4720,N_2769,N_2734);
xnor U4721 (N_4721,N_2372,N_3346);
or U4722 (N_4722,N_2713,N_3366);
and U4723 (N_4723,N_2038,N_3351);
or U4724 (N_4724,N_2368,N_3416);
nand U4725 (N_4725,N_2965,N_2092);
nand U4726 (N_4726,N_3610,N_2599);
nand U4727 (N_4727,N_3978,N_3860);
xnor U4728 (N_4728,N_3064,N_2116);
and U4729 (N_4729,N_2988,N_2184);
nand U4730 (N_4730,N_2612,N_2552);
and U4731 (N_4731,N_2533,N_3267);
and U4732 (N_4732,N_3385,N_3708);
nor U4733 (N_4733,N_2687,N_2745);
and U4734 (N_4734,N_2891,N_2190);
and U4735 (N_4735,N_2340,N_2243);
nand U4736 (N_4736,N_3923,N_3718);
or U4737 (N_4737,N_2576,N_3609);
or U4738 (N_4738,N_3852,N_3794);
xnor U4739 (N_4739,N_2780,N_3777);
or U4740 (N_4740,N_2045,N_3341);
or U4741 (N_4741,N_2848,N_3432);
and U4742 (N_4742,N_3719,N_2462);
or U4743 (N_4743,N_3593,N_3586);
nand U4744 (N_4744,N_3961,N_3074);
or U4745 (N_4745,N_2328,N_3143);
xnor U4746 (N_4746,N_2277,N_3423);
or U4747 (N_4747,N_3827,N_2282);
nand U4748 (N_4748,N_3386,N_3943);
or U4749 (N_4749,N_3195,N_3169);
nor U4750 (N_4750,N_3572,N_3139);
nand U4751 (N_4751,N_2017,N_2515);
nand U4752 (N_4752,N_2075,N_2088);
or U4753 (N_4753,N_2361,N_2254);
nand U4754 (N_4754,N_2177,N_3549);
and U4755 (N_4755,N_2281,N_3958);
nor U4756 (N_4756,N_2575,N_2308);
xnor U4757 (N_4757,N_2464,N_2584);
and U4758 (N_4758,N_2931,N_2360);
and U4759 (N_4759,N_2467,N_3809);
xnor U4760 (N_4760,N_3176,N_2336);
nor U4761 (N_4761,N_2547,N_2860);
nor U4762 (N_4762,N_2871,N_2510);
and U4763 (N_4763,N_3739,N_3652);
nand U4764 (N_4764,N_2797,N_3136);
nor U4765 (N_4765,N_3625,N_3912);
xor U4766 (N_4766,N_3072,N_2471);
nand U4767 (N_4767,N_2947,N_3514);
nand U4768 (N_4768,N_3503,N_2932);
nor U4769 (N_4769,N_3437,N_3400);
or U4770 (N_4770,N_3567,N_2928);
and U4771 (N_4771,N_2637,N_3376);
nand U4772 (N_4772,N_3879,N_3737);
nor U4773 (N_4773,N_2851,N_3454);
nor U4774 (N_4774,N_3198,N_2558);
nor U4775 (N_4775,N_2804,N_3969);
xnor U4776 (N_4776,N_3120,N_2792);
nand U4777 (N_4777,N_3033,N_3118);
nor U4778 (N_4778,N_3312,N_2173);
or U4779 (N_4779,N_3145,N_2554);
or U4780 (N_4780,N_2911,N_2923);
and U4781 (N_4781,N_3361,N_3605);
nand U4782 (N_4782,N_2295,N_2074);
nor U4783 (N_4783,N_3689,N_3436);
or U4784 (N_4784,N_2147,N_3668);
and U4785 (N_4785,N_3067,N_2946);
nand U4786 (N_4786,N_3599,N_3316);
xor U4787 (N_4787,N_2910,N_3836);
and U4788 (N_4788,N_3795,N_2631);
xor U4789 (N_4789,N_2417,N_3509);
xnor U4790 (N_4790,N_3359,N_2237);
nor U4791 (N_4791,N_2394,N_3741);
and U4792 (N_4792,N_2743,N_2007);
nand U4793 (N_4793,N_3596,N_2949);
and U4794 (N_4794,N_3770,N_3859);
or U4795 (N_4795,N_3531,N_3502);
xor U4796 (N_4796,N_3093,N_3382);
nor U4797 (N_4797,N_3616,N_3022);
nand U4798 (N_4798,N_2710,N_3965);
xor U4799 (N_4799,N_2995,N_3178);
nand U4800 (N_4800,N_2613,N_3425);
nand U4801 (N_4801,N_3461,N_3055);
xor U4802 (N_4802,N_3308,N_3025);
xor U4803 (N_4803,N_3137,N_3855);
nor U4804 (N_4804,N_3899,N_2369);
nand U4805 (N_4805,N_3557,N_3056);
and U4806 (N_4806,N_3016,N_2024);
xor U4807 (N_4807,N_2455,N_2220);
and U4808 (N_4808,N_2506,N_2348);
nand U4809 (N_4809,N_3297,N_2098);
or U4810 (N_4810,N_3751,N_3058);
nand U4811 (N_4811,N_3942,N_2667);
nand U4812 (N_4812,N_3247,N_3712);
or U4813 (N_4813,N_2108,N_2275);
or U4814 (N_4814,N_2920,N_3222);
or U4815 (N_4815,N_3216,N_3487);
or U4816 (N_4816,N_3886,N_2063);
nor U4817 (N_4817,N_3199,N_3846);
and U4818 (N_4818,N_3934,N_2794);
or U4819 (N_4819,N_3440,N_3017);
xor U4820 (N_4820,N_3212,N_3111);
and U4821 (N_4821,N_3189,N_2026);
and U4822 (N_4822,N_2085,N_3206);
and U4823 (N_4823,N_3413,N_3326);
nor U4824 (N_4824,N_2529,N_2232);
or U4825 (N_4825,N_3419,N_3779);
and U4826 (N_4826,N_2122,N_3672);
or U4827 (N_4827,N_3861,N_3482);
xor U4828 (N_4828,N_3802,N_3374);
nand U4829 (N_4829,N_2791,N_2330);
xnor U4830 (N_4830,N_2675,N_3288);
nand U4831 (N_4831,N_3219,N_3009);
nor U4832 (N_4832,N_3928,N_3532);
xnor U4833 (N_4833,N_2724,N_3649);
xor U4834 (N_4834,N_3051,N_2485);
nand U4835 (N_4835,N_3875,N_2831);
nor U4836 (N_4836,N_2205,N_3094);
nor U4837 (N_4837,N_3275,N_2930);
or U4838 (N_4838,N_3135,N_2635);
xnor U4839 (N_4839,N_2216,N_3406);
or U4840 (N_4840,N_3951,N_3389);
nand U4841 (N_4841,N_2522,N_3152);
nand U4842 (N_4842,N_3489,N_2451);
nor U4843 (N_4843,N_2894,N_2287);
or U4844 (N_4844,N_2488,N_2081);
xor U4845 (N_4845,N_2749,N_2114);
nor U4846 (N_4846,N_3542,N_3205);
and U4847 (N_4847,N_3293,N_3298);
xor U4848 (N_4848,N_3257,N_2071);
xor U4849 (N_4849,N_3501,N_3037);
nand U4850 (N_4850,N_3006,N_3866);
nand U4851 (N_4851,N_3237,N_2847);
nand U4852 (N_4852,N_2260,N_3704);
nor U4853 (N_4853,N_2526,N_2491);
and U4854 (N_4854,N_2225,N_3292);
xnor U4855 (N_4855,N_2741,N_2153);
nor U4856 (N_4856,N_2793,N_2779);
nand U4857 (N_4857,N_2752,N_3849);
nand U4858 (N_4858,N_3529,N_3449);
xor U4859 (N_4859,N_2382,N_3967);
xnor U4860 (N_4860,N_3900,N_3936);
nor U4861 (N_4861,N_2453,N_3473);
and U4862 (N_4862,N_2302,N_3973);
and U4863 (N_4863,N_2574,N_3662);
and U4864 (N_4864,N_2307,N_2043);
xor U4865 (N_4865,N_2882,N_2974);
xor U4866 (N_4866,N_2096,N_2323);
nor U4867 (N_4867,N_3049,N_3114);
or U4868 (N_4868,N_2695,N_2133);
and U4869 (N_4869,N_3038,N_2728);
and U4870 (N_4870,N_3468,N_2983);
xnor U4871 (N_4871,N_2905,N_2877);
and U4872 (N_4872,N_2658,N_3732);
and U4873 (N_4873,N_3207,N_3315);
nand U4874 (N_4874,N_2714,N_2807);
and U4875 (N_4875,N_2618,N_3915);
or U4876 (N_4876,N_2103,N_3980);
or U4877 (N_4877,N_2197,N_3495);
or U4878 (N_4878,N_3391,N_3476);
nand U4879 (N_4879,N_2843,N_2296);
xnor U4880 (N_4880,N_2545,N_2034);
nand U4881 (N_4881,N_3245,N_3674);
xnor U4882 (N_4882,N_3892,N_3447);
xnor U4883 (N_4883,N_2018,N_3353);
or U4884 (N_4884,N_3954,N_3714);
and U4885 (N_4885,N_3095,N_2616);
nand U4886 (N_4886,N_2978,N_2288);
nor U4887 (N_4887,N_3153,N_3960);
xor U4888 (N_4888,N_2493,N_2011);
or U4889 (N_4889,N_3357,N_2093);
xor U4890 (N_4890,N_2952,N_3667);
or U4891 (N_4891,N_3269,N_3930);
and U4892 (N_4892,N_3730,N_3165);
or U4893 (N_4893,N_2438,N_3678);
and U4894 (N_4894,N_2539,N_3742);
xnor U4895 (N_4895,N_2384,N_2273);
nand U4896 (N_4896,N_2331,N_3103);
nor U4897 (N_4897,N_2053,N_3924);
nand U4898 (N_4898,N_3727,N_3276);
or U4899 (N_4899,N_3043,N_3766);
nand U4900 (N_4900,N_3077,N_3401);
nor U4901 (N_4901,N_3160,N_3270);
or U4902 (N_4902,N_3816,N_3582);
nand U4903 (N_4903,N_2977,N_3041);
nor U4904 (N_4904,N_2839,N_3380);
and U4905 (N_4905,N_3663,N_2727);
nand U4906 (N_4906,N_3711,N_2731);
xor U4907 (N_4907,N_3444,N_3410);
and U4908 (N_4908,N_2996,N_2135);
nor U4909 (N_4909,N_2006,N_3010);
xor U4910 (N_4910,N_3268,N_2261);
and U4911 (N_4911,N_2106,N_2528);
nor U4912 (N_4912,N_2655,N_3530);
xor U4913 (N_4913,N_3575,N_3434);
nand U4914 (N_4914,N_2970,N_2263);
xor U4915 (N_4915,N_2251,N_2972);
or U4916 (N_4916,N_2973,N_2386);
nand U4917 (N_4917,N_3282,N_3854);
nor U4918 (N_4918,N_2439,N_2315);
xor U4919 (N_4919,N_3546,N_2546);
nor U4920 (N_4920,N_2304,N_3626);
and U4921 (N_4921,N_2913,N_2352);
xor U4922 (N_4922,N_3318,N_2218);
xor U4923 (N_4923,N_2311,N_2255);
xnor U4924 (N_4924,N_3736,N_3066);
xnor U4925 (N_4925,N_3762,N_3162);
nor U4926 (N_4926,N_2961,N_3455);
and U4927 (N_4927,N_3981,N_3005);
or U4928 (N_4928,N_2039,N_2639);
nor U4929 (N_4929,N_3655,N_3272);
or U4930 (N_4930,N_2371,N_3334);
and U4931 (N_4931,N_3054,N_3823);
nand U4932 (N_4932,N_3780,N_3508);
nand U4933 (N_4933,N_2112,N_2934);
nor U4934 (N_4934,N_3175,N_2590);
xnor U4935 (N_4935,N_3757,N_3204);
nand U4936 (N_4936,N_2883,N_3580);
and U4937 (N_4937,N_3510,N_3352);
and U4938 (N_4938,N_3966,N_2984);
and U4939 (N_4939,N_2040,N_2676);
and U4940 (N_4940,N_2131,N_3666);
or U4941 (N_4941,N_2068,N_3955);
nor U4942 (N_4942,N_2671,N_2420);
and U4943 (N_4943,N_2150,N_2226);
or U4944 (N_4944,N_2588,N_3871);
or U4945 (N_4945,N_2908,N_2327);
nor U4946 (N_4946,N_2449,N_2407);
nand U4947 (N_4947,N_3706,N_3953);
and U4948 (N_4948,N_3984,N_2303);
nand U4949 (N_4949,N_2781,N_2021);
nor U4950 (N_4950,N_2953,N_3541);
nor U4951 (N_4951,N_2235,N_2022);
nor U4952 (N_4952,N_2306,N_2856);
and U4953 (N_4953,N_2959,N_3271);
or U4954 (N_4954,N_2253,N_3676);
nor U4955 (N_4955,N_2709,N_2600);
nand U4956 (N_4956,N_2215,N_3494);
nor U4957 (N_4957,N_2670,N_3246);
and U4958 (N_4958,N_3026,N_2078);
or U4959 (N_4959,N_3375,N_2266);
nand U4960 (N_4960,N_3740,N_3611);
or U4961 (N_4961,N_2431,N_2723);
nand U4962 (N_4962,N_2568,N_3622);
or U4963 (N_4963,N_2207,N_2508);
or U4964 (N_4964,N_2258,N_2742);
nand U4965 (N_4965,N_3036,N_3785);
nand U4966 (N_4966,N_2549,N_3639);
and U4967 (N_4967,N_2739,N_3311);
and U4968 (N_4968,N_3728,N_3519);
nor U4969 (N_4969,N_2633,N_3422);
nand U4970 (N_4970,N_3537,N_2036);
and U4971 (N_4971,N_2206,N_3261);
or U4972 (N_4972,N_2238,N_2976);
xor U4973 (N_4973,N_3424,N_2874);
and U4974 (N_4974,N_2383,N_2706);
and U4975 (N_4975,N_2813,N_2717);
xnor U4976 (N_4976,N_2688,N_3937);
xnor U4977 (N_4977,N_2274,N_3922);
nand U4978 (N_4978,N_2815,N_2594);
xnor U4979 (N_4979,N_3665,N_2922);
or U4980 (N_4980,N_3614,N_2798);
or U4981 (N_4981,N_2502,N_2000);
nor U4982 (N_4982,N_3277,N_2223);
xor U4983 (N_4983,N_3818,N_3463);
or U4984 (N_4984,N_2817,N_2412);
nor U4985 (N_4985,N_2942,N_3760);
xor U4986 (N_4986,N_2524,N_2248);
xor U4987 (N_4987,N_2222,N_2864);
or U4988 (N_4988,N_2927,N_3898);
nand U4989 (N_4989,N_2975,N_2997);
or U4990 (N_4990,N_3897,N_3259);
nor U4991 (N_4991,N_3342,N_2061);
nand U4992 (N_4992,N_2076,N_3408);
nor U4993 (N_4993,N_2012,N_2278);
and U4994 (N_4994,N_3194,N_3612);
nand U4995 (N_4995,N_2127,N_2735);
nand U4996 (N_4996,N_2810,N_3533);
or U4997 (N_4997,N_3379,N_3701);
nor U4998 (N_4998,N_3820,N_3188);
and U4999 (N_4999,N_2137,N_3539);
or U5000 (N_5000,N_2810,N_3017);
and U5001 (N_5001,N_3608,N_3813);
xnor U5002 (N_5002,N_2279,N_2094);
or U5003 (N_5003,N_2296,N_2691);
xor U5004 (N_5004,N_2993,N_3362);
nand U5005 (N_5005,N_2645,N_3939);
or U5006 (N_5006,N_2534,N_3965);
or U5007 (N_5007,N_2006,N_3784);
and U5008 (N_5008,N_2404,N_3087);
nor U5009 (N_5009,N_3167,N_2096);
nand U5010 (N_5010,N_2213,N_3949);
nand U5011 (N_5011,N_2188,N_3924);
xor U5012 (N_5012,N_2093,N_3569);
nand U5013 (N_5013,N_2389,N_3942);
nand U5014 (N_5014,N_3236,N_2475);
nand U5015 (N_5015,N_3286,N_3499);
and U5016 (N_5016,N_3397,N_2620);
or U5017 (N_5017,N_2866,N_2658);
nand U5018 (N_5018,N_3843,N_3916);
or U5019 (N_5019,N_3044,N_3661);
or U5020 (N_5020,N_3794,N_2376);
xnor U5021 (N_5021,N_3624,N_3591);
or U5022 (N_5022,N_3754,N_3359);
or U5023 (N_5023,N_2872,N_2895);
nand U5024 (N_5024,N_3029,N_3941);
and U5025 (N_5025,N_2012,N_3280);
nand U5026 (N_5026,N_2832,N_3953);
and U5027 (N_5027,N_2118,N_2009);
nand U5028 (N_5028,N_2051,N_3669);
xor U5029 (N_5029,N_2255,N_2062);
xor U5030 (N_5030,N_2916,N_3554);
or U5031 (N_5031,N_2175,N_2325);
or U5032 (N_5032,N_3437,N_2557);
and U5033 (N_5033,N_3019,N_3491);
xnor U5034 (N_5034,N_3109,N_3987);
xor U5035 (N_5035,N_3418,N_2491);
nand U5036 (N_5036,N_3872,N_3184);
nor U5037 (N_5037,N_2199,N_3543);
and U5038 (N_5038,N_3342,N_3126);
nor U5039 (N_5039,N_3565,N_2221);
or U5040 (N_5040,N_2727,N_2876);
nor U5041 (N_5041,N_3026,N_3223);
or U5042 (N_5042,N_3307,N_2691);
xnor U5043 (N_5043,N_2760,N_3207);
nand U5044 (N_5044,N_3750,N_3497);
xor U5045 (N_5045,N_2431,N_2699);
and U5046 (N_5046,N_2938,N_2321);
and U5047 (N_5047,N_3115,N_2838);
nand U5048 (N_5048,N_3439,N_2908);
and U5049 (N_5049,N_3003,N_3362);
xnor U5050 (N_5050,N_3194,N_3505);
nor U5051 (N_5051,N_3710,N_2868);
or U5052 (N_5052,N_3838,N_3350);
or U5053 (N_5053,N_3500,N_2662);
nand U5054 (N_5054,N_3905,N_2924);
nand U5055 (N_5055,N_2456,N_3189);
nor U5056 (N_5056,N_3188,N_3339);
xor U5057 (N_5057,N_3538,N_3666);
nand U5058 (N_5058,N_3951,N_2642);
and U5059 (N_5059,N_2893,N_3075);
nand U5060 (N_5060,N_3961,N_2184);
nand U5061 (N_5061,N_3969,N_2540);
and U5062 (N_5062,N_2552,N_3807);
nand U5063 (N_5063,N_3015,N_3414);
nand U5064 (N_5064,N_3630,N_3873);
nand U5065 (N_5065,N_3031,N_3975);
nand U5066 (N_5066,N_3980,N_3587);
nor U5067 (N_5067,N_3365,N_3991);
nand U5068 (N_5068,N_3310,N_2754);
and U5069 (N_5069,N_3144,N_3396);
xor U5070 (N_5070,N_3274,N_2134);
and U5071 (N_5071,N_2245,N_3005);
nand U5072 (N_5072,N_2368,N_3355);
or U5073 (N_5073,N_2012,N_3428);
nor U5074 (N_5074,N_2249,N_3477);
or U5075 (N_5075,N_3978,N_2486);
and U5076 (N_5076,N_2865,N_2091);
and U5077 (N_5077,N_2887,N_3896);
xor U5078 (N_5078,N_3784,N_3541);
and U5079 (N_5079,N_3288,N_3436);
and U5080 (N_5080,N_3876,N_2176);
nand U5081 (N_5081,N_2817,N_2975);
and U5082 (N_5082,N_2405,N_3802);
and U5083 (N_5083,N_2510,N_2355);
and U5084 (N_5084,N_2642,N_2872);
xor U5085 (N_5085,N_2262,N_3191);
or U5086 (N_5086,N_3798,N_2599);
nand U5087 (N_5087,N_2093,N_2081);
or U5088 (N_5088,N_3194,N_2727);
nand U5089 (N_5089,N_3677,N_3316);
nand U5090 (N_5090,N_3186,N_2489);
xnor U5091 (N_5091,N_2515,N_2344);
nor U5092 (N_5092,N_2993,N_2509);
or U5093 (N_5093,N_3684,N_2910);
nor U5094 (N_5094,N_2235,N_3908);
nand U5095 (N_5095,N_2310,N_2658);
and U5096 (N_5096,N_2837,N_3788);
xor U5097 (N_5097,N_3740,N_3533);
nor U5098 (N_5098,N_2839,N_2049);
nand U5099 (N_5099,N_2885,N_2955);
xor U5100 (N_5100,N_3494,N_3755);
and U5101 (N_5101,N_2764,N_2426);
nor U5102 (N_5102,N_2064,N_2819);
and U5103 (N_5103,N_2783,N_2354);
and U5104 (N_5104,N_2318,N_3507);
or U5105 (N_5105,N_2395,N_3210);
or U5106 (N_5106,N_3736,N_3713);
or U5107 (N_5107,N_3632,N_3893);
or U5108 (N_5108,N_3746,N_2162);
or U5109 (N_5109,N_2313,N_3197);
nand U5110 (N_5110,N_3004,N_3844);
xor U5111 (N_5111,N_3854,N_2015);
or U5112 (N_5112,N_2607,N_3482);
nand U5113 (N_5113,N_2906,N_2571);
nand U5114 (N_5114,N_2677,N_3139);
and U5115 (N_5115,N_2137,N_3596);
nor U5116 (N_5116,N_2889,N_2239);
xor U5117 (N_5117,N_2157,N_3420);
xor U5118 (N_5118,N_2226,N_2037);
or U5119 (N_5119,N_2222,N_2560);
and U5120 (N_5120,N_3394,N_3393);
and U5121 (N_5121,N_2885,N_3625);
or U5122 (N_5122,N_2515,N_3507);
and U5123 (N_5123,N_2293,N_3694);
nor U5124 (N_5124,N_2364,N_3448);
and U5125 (N_5125,N_3019,N_3105);
xnor U5126 (N_5126,N_3328,N_3442);
nand U5127 (N_5127,N_2506,N_2163);
xor U5128 (N_5128,N_3488,N_2898);
xor U5129 (N_5129,N_2803,N_2144);
and U5130 (N_5130,N_2298,N_3740);
nand U5131 (N_5131,N_3459,N_3373);
nor U5132 (N_5132,N_3118,N_3920);
xor U5133 (N_5133,N_3927,N_2334);
nand U5134 (N_5134,N_3384,N_2979);
nor U5135 (N_5135,N_2557,N_3345);
nand U5136 (N_5136,N_2088,N_2748);
nor U5137 (N_5137,N_2548,N_2712);
and U5138 (N_5138,N_3451,N_2098);
xor U5139 (N_5139,N_3855,N_3274);
or U5140 (N_5140,N_3826,N_3232);
nand U5141 (N_5141,N_3698,N_3583);
nor U5142 (N_5142,N_3332,N_3248);
and U5143 (N_5143,N_2350,N_2745);
and U5144 (N_5144,N_2918,N_3529);
and U5145 (N_5145,N_3836,N_3684);
and U5146 (N_5146,N_3088,N_2454);
nand U5147 (N_5147,N_2322,N_2419);
nor U5148 (N_5148,N_2945,N_3943);
or U5149 (N_5149,N_2225,N_3800);
and U5150 (N_5150,N_2523,N_2539);
or U5151 (N_5151,N_3801,N_2952);
nand U5152 (N_5152,N_3012,N_3525);
and U5153 (N_5153,N_3682,N_3611);
and U5154 (N_5154,N_2769,N_3934);
xor U5155 (N_5155,N_2140,N_2230);
nand U5156 (N_5156,N_3481,N_3794);
or U5157 (N_5157,N_2327,N_2906);
nand U5158 (N_5158,N_2646,N_2910);
and U5159 (N_5159,N_2214,N_3458);
xnor U5160 (N_5160,N_3765,N_2561);
and U5161 (N_5161,N_3776,N_2986);
nor U5162 (N_5162,N_3533,N_3638);
and U5163 (N_5163,N_3965,N_2366);
nor U5164 (N_5164,N_2771,N_3885);
nand U5165 (N_5165,N_2950,N_3223);
xor U5166 (N_5166,N_3593,N_2084);
xnor U5167 (N_5167,N_2741,N_2539);
nor U5168 (N_5168,N_2672,N_2165);
nor U5169 (N_5169,N_3791,N_3596);
nor U5170 (N_5170,N_3856,N_2710);
and U5171 (N_5171,N_3566,N_2632);
xor U5172 (N_5172,N_2009,N_3527);
or U5173 (N_5173,N_2758,N_2988);
and U5174 (N_5174,N_2611,N_3619);
xor U5175 (N_5175,N_3145,N_2465);
xnor U5176 (N_5176,N_3855,N_3438);
xor U5177 (N_5177,N_2330,N_2273);
and U5178 (N_5178,N_3122,N_3491);
or U5179 (N_5179,N_3902,N_2672);
and U5180 (N_5180,N_2378,N_2918);
nand U5181 (N_5181,N_3102,N_3623);
nand U5182 (N_5182,N_2046,N_3251);
or U5183 (N_5183,N_3813,N_3452);
or U5184 (N_5184,N_3486,N_2964);
xnor U5185 (N_5185,N_3793,N_2520);
xor U5186 (N_5186,N_3755,N_3797);
and U5187 (N_5187,N_2081,N_3456);
nor U5188 (N_5188,N_2454,N_2025);
and U5189 (N_5189,N_3501,N_2367);
or U5190 (N_5190,N_3053,N_2880);
or U5191 (N_5191,N_3910,N_2520);
xnor U5192 (N_5192,N_3573,N_3447);
nand U5193 (N_5193,N_2965,N_2577);
xnor U5194 (N_5194,N_2279,N_3549);
xnor U5195 (N_5195,N_3817,N_2646);
nand U5196 (N_5196,N_2369,N_3220);
or U5197 (N_5197,N_3204,N_2295);
nand U5198 (N_5198,N_3004,N_2112);
nor U5199 (N_5199,N_3873,N_3742);
or U5200 (N_5200,N_3964,N_3325);
and U5201 (N_5201,N_2250,N_3818);
nand U5202 (N_5202,N_2505,N_2142);
and U5203 (N_5203,N_3129,N_3757);
nand U5204 (N_5204,N_3916,N_2549);
nor U5205 (N_5205,N_2189,N_3158);
and U5206 (N_5206,N_3390,N_2291);
nand U5207 (N_5207,N_3194,N_3882);
and U5208 (N_5208,N_3223,N_2366);
xnor U5209 (N_5209,N_3614,N_3784);
nor U5210 (N_5210,N_3359,N_3240);
and U5211 (N_5211,N_2922,N_2203);
xor U5212 (N_5212,N_2078,N_3229);
and U5213 (N_5213,N_2590,N_2118);
and U5214 (N_5214,N_2228,N_3853);
nor U5215 (N_5215,N_2648,N_3860);
and U5216 (N_5216,N_2445,N_2239);
nand U5217 (N_5217,N_2730,N_2583);
nor U5218 (N_5218,N_2814,N_3493);
and U5219 (N_5219,N_3387,N_2843);
or U5220 (N_5220,N_2633,N_2037);
and U5221 (N_5221,N_2935,N_2439);
nor U5222 (N_5222,N_3990,N_3662);
xnor U5223 (N_5223,N_3440,N_3537);
or U5224 (N_5224,N_2111,N_3065);
nor U5225 (N_5225,N_2463,N_3183);
nand U5226 (N_5226,N_3772,N_2730);
nand U5227 (N_5227,N_2623,N_3373);
nor U5228 (N_5228,N_2802,N_2120);
nor U5229 (N_5229,N_3707,N_3890);
nand U5230 (N_5230,N_3045,N_3748);
or U5231 (N_5231,N_3629,N_3199);
nor U5232 (N_5232,N_3039,N_3530);
nor U5233 (N_5233,N_2608,N_3368);
or U5234 (N_5234,N_3131,N_3224);
nand U5235 (N_5235,N_2666,N_2041);
and U5236 (N_5236,N_3060,N_2710);
nor U5237 (N_5237,N_3175,N_3177);
nand U5238 (N_5238,N_3317,N_3880);
xnor U5239 (N_5239,N_3211,N_2372);
xnor U5240 (N_5240,N_2863,N_3529);
or U5241 (N_5241,N_2641,N_3620);
or U5242 (N_5242,N_2410,N_2175);
and U5243 (N_5243,N_3646,N_2716);
and U5244 (N_5244,N_2405,N_2709);
nand U5245 (N_5245,N_3685,N_3385);
nor U5246 (N_5246,N_3710,N_2750);
nor U5247 (N_5247,N_2496,N_2626);
and U5248 (N_5248,N_3665,N_2979);
nor U5249 (N_5249,N_2757,N_2971);
nor U5250 (N_5250,N_3319,N_2204);
and U5251 (N_5251,N_2904,N_2947);
nand U5252 (N_5252,N_3993,N_2341);
nor U5253 (N_5253,N_2881,N_3409);
and U5254 (N_5254,N_2747,N_2528);
xnor U5255 (N_5255,N_2452,N_3771);
or U5256 (N_5256,N_3835,N_2218);
or U5257 (N_5257,N_2963,N_3388);
and U5258 (N_5258,N_2753,N_3045);
and U5259 (N_5259,N_3517,N_3753);
nand U5260 (N_5260,N_2493,N_3547);
xor U5261 (N_5261,N_2855,N_3320);
nand U5262 (N_5262,N_3397,N_3041);
nand U5263 (N_5263,N_2704,N_2910);
and U5264 (N_5264,N_3643,N_2008);
or U5265 (N_5265,N_3873,N_3510);
and U5266 (N_5266,N_3756,N_2404);
or U5267 (N_5267,N_2388,N_3449);
nand U5268 (N_5268,N_2324,N_3328);
and U5269 (N_5269,N_2715,N_2116);
or U5270 (N_5270,N_3761,N_3766);
xnor U5271 (N_5271,N_3034,N_2616);
and U5272 (N_5272,N_2814,N_2397);
xor U5273 (N_5273,N_3558,N_3218);
xnor U5274 (N_5274,N_3602,N_3915);
xnor U5275 (N_5275,N_3395,N_3533);
nor U5276 (N_5276,N_3269,N_2992);
or U5277 (N_5277,N_3523,N_3620);
nor U5278 (N_5278,N_3590,N_3073);
or U5279 (N_5279,N_3120,N_2904);
xor U5280 (N_5280,N_3914,N_2609);
nand U5281 (N_5281,N_2483,N_2000);
nand U5282 (N_5282,N_2117,N_3018);
nor U5283 (N_5283,N_3263,N_3678);
and U5284 (N_5284,N_2411,N_3343);
or U5285 (N_5285,N_3796,N_2045);
xor U5286 (N_5286,N_2808,N_3398);
or U5287 (N_5287,N_2115,N_3286);
and U5288 (N_5288,N_2442,N_2707);
nor U5289 (N_5289,N_2625,N_3952);
or U5290 (N_5290,N_3093,N_3006);
nor U5291 (N_5291,N_2608,N_2347);
nor U5292 (N_5292,N_2427,N_3013);
nand U5293 (N_5293,N_3232,N_2951);
nor U5294 (N_5294,N_2041,N_3462);
xnor U5295 (N_5295,N_2431,N_3381);
nor U5296 (N_5296,N_3746,N_3808);
or U5297 (N_5297,N_2111,N_2170);
xnor U5298 (N_5298,N_2239,N_3752);
nor U5299 (N_5299,N_2133,N_2417);
xnor U5300 (N_5300,N_2874,N_2154);
nand U5301 (N_5301,N_3797,N_3598);
or U5302 (N_5302,N_2761,N_2651);
or U5303 (N_5303,N_2983,N_2207);
xor U5304 (N_5304,N_3401,N_2558);
nor U5305 (N_5305,N_2108,N_2283);
nand U5306 (N_5306,N_2269,N_2315);
nand U5307 (N_5307,N_2020,N_3595);
or U5308 (N_5308,N_3181,N_3023);
xor U5309 (N_5309,N_2095,N_3232);
nor U5310 (N_5310,N_2483,N_3458);
xor U5311 (N_5311,N_2156,N_3105);
nand U5312 (N_5312,N_2580,N_2043);
and U5313 (N_5313,N_3533,N_3988);
and U5314 (N_5314,N_2061,N_2389);
nor U5315 (N_5315,N_2230,N_2163);
and U5316 (N_5316,N_2836,N_3051);
or U5317 (N_5317,N_3637,N_2869);
or U5318 (N_5318,N_3802,N_2039);
xnor U5319 (N_5319,N_3421,N_3061);
xor U5320 (N_5320,N_2280,N_2572);
or U5321 (N_5321,N_3772,N_3787);
or U5322 (N_5322,N_3312,N_3336);
or U5323 (N_5323,N_2047,N_3968);
or U5324 (N_5324,N_2265,N_3630);
xor U5325 (N_5325,N_2567,N_2621);
or U5326 (N_5326,N_3476,N_2871);
nor U5327 (N_5327,N_2872,N_3220);
nand U5328 (N_5328,N_2287,N_2465);
xnor U5329 (N_5329,N_2726,N_3276);
and U5330 (N_5330,N_2916,N_2870);
or U5331 (N_5331,N_2610,N_3026);
nor U5332 (N_5332,N_2946,N_2280);
and U5333 (N_5333,N_2233,N_3311);
and U5334 (N_5334,N_3423,N_2759);
nor U5335 (N_5335,N_3669,N_2404);
nand U5336 (N_5336,N_3046,N_3435);
or U5337 (N_5337,N_2304,N_2334);
and U5338 (N_5338,N_3685,N_3869);
or U5339 (N_5339,N_3990,N_3576);
or U5340 (N_5340,N_2298,N_3908);
and U5341 (N_5341,N_2232,N_3478);
and U5342 (N_5342,N_2300,N_2341);
xor U5343 (N_5343,N_2849,N_2720);
xor U5344 (N_5344,N_2064,N_3562);
nand U5345 (N_5345,N_2691,N_3717);
nor U5346 (N_5346,N_3045,N_2804);
nand U5347 (N_5347,N_3000,N_3282);
or U5348 (N_5348,N_2850,N_3699);
and U5349 (N_5349,N_3879,N_2369);
or U5350 (N_5350,N_3214,N_3472);
or U5351 (N_5351,N_3981,N_3245);
xnor U5352 (N_5352,N_3945,N_3652);
nor U5353 (N_5353,N_2767,N_3742);
or U5354 (N_5354,N_2375,N_2011);
xnor U5355 (N_5355,N_3406,N_2279);
nand U5356 (N_5356,N_2267,N_2577);
xor U5357 (N_5357,N_2658,N_3686);
xor U5358 (N_5358,N_2344,N_3553);
nor U5359 (N_5359,N_3336,N_2689);
nor U5360 (N_5360,N_2670,N_3140);
nor U5361 (N_5361,N_3462,N_2806);
and U5362 (N_5362,N_2084,N_2908);
or U5363 (N_5363,N_2778,N_3203);
or U5364 (N_5364,N_3387,N_2354);
nor U5365 (N_5365,N_2275,N_2367);
xor U5366 (N_5366,N_3396,N_2750);
xnor U5367 (N_5367,N_3399,N_2890);
or U5368 (N_5368,N_2139,N_2176);
and U5369 (N_5369,N_2023,N_3331);
nor U5370 (N_5370,N_2472,N_3159);
and U5371 (N_5371,N_3164,N_3750);
and U5372 (N_5372,N_2510,N_3856);
nand U5373 (N_5373,N_3246,N_3206);
xnor U5374 (N_5374,N_2830,N_3732);
and U5375 (N_5375,N_3373,N_3863);
nor U5376 (N_5376,N_2219,N_3200);
xor U5377 (N_5377,N_2622,N_2788);
xor U5378 (N_5378,N_2883,N_3927);
or U5379 (N_5379,N_2842,N_2896);
nor U5380 (N_5380,N_2568,N_3197);
nor U5381 (N_5381,N_2420,N_2288);
nand U5382 (N_5382,N_3508,N_2313);
xor U5383 (N_5383,N_3826,N_3929);
xnor U5384 (N_5384,N_3510,N_3394);
or U5385 (N_5385,N_2520,N_3631);
or U5386 (N_5386,N_2543,N_3635);
and U5387 (N_5387,N_3160,N_2645);
xnor U5388 (N_5388,N_2478,N_2676);
and U5389 (N_5389,N_3801,N_2537);
and U5390 (N_5390,N_3823,N_3173);
nor U5391 (N_5391,N_2511,N_3556);
nand U5392 (N_5392,N_2828,N_3127);
nor U5393 (N_5393,N_3175,N_2876);
nand U5394 (N_5394,N_3659,N_2046);
and U5395 (N_5395,N_2476,N_3999);
nor U5396 (N_5396,N_3804,N_2319);
or U5397 (N_5397,N_3852,N_2484);
or U5398 (N_5398,N_2605,N_3296);
nand U5399 (N_5399,N_2277,N_2163);
nor U5400 (N_5400,N_2283,N_3468);
xor U5401 (N_5401,N_2489,N_3191);
nor U5402 (N_5402,N_3326,N_3521);
nand U5403 (N_5403,N_2757,N_3476);
xor U5404 (N_5404,N_2291,N_3480);
nand U5405 (N_5405,N_2645,N_3265);
or U5406 (N_5406,N_2681,N_3961);
nand U5407 (N_5407,N_3068,N_3042);
xor U5408 (N_5408,N_2995,N_2797);
nand U5409 (N_5409,N_3211,N_2652);
and U5410 (N_5410,N_2806,N_2904);
xnor U5411 (N_5411,N_2099,N_2809);
nand U5412 (N_5412,N_2410,N_3353);
nand U5413 (N_5413,N_3261,N_2746);
nor U5414 (N_5414,N_2395,N_3722);
and U5415 (N_5415,N_2536,N_2715);
or U5416 (N_5416,N_3360,N_3194);
xor U5417 (N_5417,N_2731,N_2536);
nor U5418 (N_5418,N_2431,N_3472);
xnor U5419 (N_5419,N_2967,N_2995);
and U5420 (N_5420,N_3827,N_3650);
nor U5421 (N_5421,N_2991,N_2952);
xor U5422 (N_5422,N_3839,N_2937);
nor U5423 (N_5423,N_3287,N_3534);
and U5424 (N_5424,N_2202,N_3209);
nor U5425 (N_5425,N_3196,N_2886);
or U5426 (N_5426,N_3141,N_3831);
nor U5427 (N_5427,N_2384,N_3003);
or U5428 (N_5428,N_2046,N_2833);
nand U5429 (N_5429,N_3937,N_3142);
or U5430 (N_5430,N_3309,N_2567);
and U5431 (N_5431,N_3951,N_3977);
nand U5432 (N_5432,N_3740,N_3447);
nor U5433 (N_5433,N_2045,N_2808);
and U5434 (N_5434,N_3579,N_2144);
and U5435 (N_5435,N_3483,N_2962);
nand U5436 (N_5436,N_2423,N_2438);
nand U5437 (N_5437,N_3247,N_2816);
nor U5438 (N_5438,N_2599,N_2364);
nand U5439 (N_5439,N_2326,N_3895);
xor U5440 (N_5440,N_2774,N_2161);
nand U5441 (N_5441,N_3025,N_3279);
nor U5442 (N_5442,N_3363,N_3558);
xor U5443 (N_5443,N_2436,N_3482);
nor U5444 (N_5444,N_2333,N_3926);
xor U5445 (N_5445,N_3952,N_2177);
nand U5446 (N_5446,N_2184,N_3291);
and U5447 (N_5447,N_3266,N_2246);
nor U5448 (N_5448,N_3311,N_2216);
nor U5449 (N_5449,N_2848,N_2370);
and U5450 (N_5450,N_3166,N_2030);
or U5451 (N_5451,N_3876,N_2985);
and U5452 (N_5452,N_3770,N_2017);
or U5453 (N_5453,N_3242,N_3755);
xor U5454 (N_5454,N_2868,N_2354);
nor U5455 (N_5455,N_3866,N_3500);
nor U5456 (N_5456,N_2018,N_3778);
xnor U5457 (N_5457,N_2016,N_2811);
and U5458 (N_5458,N_3834,N_2621);
xor U5459 (N_5459,N_2841,N_3617);
and U5460 (N_5460,N_3069,N_2517);
or U5461 (N_5461,N_3623,N_3948);
xor U5462 (N_5462,N_2431,N_3141);
nand U5463 (N_5463,N_3686,N_3320);
nand U5464 (N_5464,N_2314,N_3224);
nor U5465 (N_5465,N_3325,N_3273);
nor U5466 (N_5466,N_2120,N_2314);
nand U5467 (N_5467,N_2128,N_2484);
xor U5468 (N_5468,N_3877,N_3617);
xnor U5469 (N_5469,N_2244,N_3653);
nand U5470 (N_5470,N_2821,N_3831);
nor U5471 (N_5471,N_3642,N_2328);
nor U5472 (N_5472,N_2082,N_3981);
or U5473 (N_5473,N_3743,N_2005);
xor U5474 (N_5474,N_2430,N_3089);
nor U5475 (N_5475,N_2155,N_2255);
or U5476 (N_5476,N_3474,N_3407);
and U5477 (N_5477,N_3146,N_2847);
nor U5478 (N_5478,N_3255,N_3092);
nor U5479 (N_5479,N_2180,N_2393);
xor U5480 (N_5480,N_3613,N_2143);
or U5481 (N_5481,N_3393,N_2943);
and U5482 (N_5482,N_3524,N_3360);
or U5483 (N_5483,N_2798,N_2899);
and U5484 (N_5484,N_3862,N_2653);
nor U5485 (N_5485,N_3713,N_2103);
or U5486 (N_5486,N_3161,N_2288);
nor U5487 (N_5487,N_3560,N_3124);
nand U5488 (N_5488,N_2254,N_2157);
nor U5489 (N_5489,N_2185,N_3139);
nand U5490 (N_5490,N_2783,N_2132);
nand U5491 (N_5491,N_3448,N_3562);
nand U5492 (N_5492,N_3491,N_3090);
nor U5493 (N_5493,N_2867,N_2321);
xnor U5494 (N_5494,N_2885,N_2261);
and U5495 (N_5495,N_2622,N_3859);
nor U5496 (N_5496,N_3729,N_3251);
nor U5497 (N_5497,N_3603,N_2204);
nand U5498 (N_5498,N_2353,N_2759);
or U5499 (N_5499,N_2036,N_2159);
and U5500 (N_5500,N_3968,N_3555);
xnor U5501 (N_5501,N_3259,N_3551);
or U5502 (N_5502,N_2207,N_3880);
xnor U5503 (N_5503,N_2676,N_3954);
nor U5504 (N_5504,N_2477,N_3847);
nor U5505 (N_5505,N_3267,N_2022);
nor U5506 (N_5506,N_3860,N_2277);
and U5507 (N_5507,N_2253,N_3728);
nand U5508 (N_5508,N_2208,N_2841);
xor U5509 (N_5509,N_3498,N_2374);
or U5510 (N_5510,N_2193,N_2609);
xnor U5511 (N_5511,N_3200,N_2625);
nor U5512 (N_5512,N_2836,N_3992);
xnor U5513 (N_5513,N_3824,N_2302);
xor U5514 (N_5514,N_2634,N_2435);
and U5515 (N_5515,N_3737,N_3421);
nand U5516 (N_5516,N_2021,N_2469);
nand U5517 (N_5517,N_3982,N_2697);
or U5518 (N_5518,N_2847,N_3864);
and U5519 (N_5519,N_2944,N_3465);
nand U5520 (N_5520,N_2875,N_3849);
xor U5521 (N_5521,N_3052,N_2220);
nor U5522 (N_5522,N_3024,N_3482);
xor U5523 (N_5523,N_2506,N_2530);
nand U5524 (N_5524,N_2198,N_2173);
xor U5525 (N_5525,N_3327,N_2241);
nor U5526 (N_5526,N_2355,N_3414);
nor U5527 (N_5527,N_2204,N_2069);
or U5528 (N_5528,N_3320,N_2165);
nand U5529 (N_5529,N_3512,N_2549);
xor U5530 (N_5530,N_2950,N_3117);
and U5531 (N_5531,N_3850,N_2072);
nand U5532 (N_5532,N_2782,N_3381);
nand U5533 (N_5533,N_2310,N_2592);
nand U5534 (N_5534,N_2569,N_2548);
or U5535 (N_5535,N_3571,N_2724);
and U5536 (N_5536,N_2937,N_2697);
nand U5537 (N_5537,N_3787,N_2133);
and U5538 (N_5538,N_3884,N_2244);
nor U5539 (N_5539,N_3626,N_3149);
nand U5540 (N_5540,N_3444,N_2844);
and U5541 (N_5541,N_2993,N_3292);
or U5542 (N_5542,N_2941,N_2884);
nor U5543 (N_5543,N_3902,N_3701);
and U5544 (N_5544,N_3191,N_3330);
xnor U5545 (N_5545,N_3751,N_3240);
and U5546 (N_5546,N_2256,N_2596);
and U5547 (N_5547,N_3334,N_2271);
or U5548 (N_5548,N_2418,N_3378);
or U5549 (N_5549,N_3885,N_3213);
xor U5550 (N_5550,N_2248,N_3783);
or U5551 (N_5551,N_2250,N_2644);
and U5552 (N_5552,N_3457,N_3116);
and U5553 (N_5553,N_2790,N_2851);
nor U5554 (N_5554,N_2276,N_2567);
and U5555 (N_5555,N_3380,N_2623);
xnor U5556 (N_5556,N_2477,N_2320);
nor U5557 (N_5557,N_3611,N_2895);
and U5558 (N_5558,N_2588,N_3127);
xor U5559 (N_5559,N_3144,N_2663);
xor U5560 (N_5560,N_2549,N_3893);
or U5561 (N_5561,N_2891,N_3470);
nand U5562 (N_5562,N_3390,N_3270);
nand U5563 (N_5563,N_3593,N_2388);
nor U5564 (N_5564,N_3255,N_2619);
or U5565 (N_5565,N_2684,N_3246);
and U5566 (N_5566,N_2653,N_2596);
nand U5567 (N_5567,N_2228,N_2041);
nand U5568 (N_5568,N_2157,N_3782);
or U5569 (N_5569,N_2936,N_3306);
and U5570 (N_5570,N_3416,N_2544);
nor U5571 (N_5571,N_2006,N_3478);
and U5572 (N_5572,N_2656,N_3227);
nor U5573 (N_5573,N_3868,N_2233);
or U5574 (N_5574,N_2462,N_3729);
or U5575 (N_5575,N_2707,N_3620);
nor U5576 (N_5576,N_2999,N_2096);
or U5577 (N_5577,N_2136,N_2273);
nor U5578 (N_5578,N_2733,N_3926);
xor U5579 (N_5579,N_2274,N_3091);
nand U5580 (N_5580,N_2900,N_3832);
nand U5581 (N_5581,N_2183,N_2791);
xor U5582 (N_5582,N_3073,N_3115);
or U5583 (N_5583,N_2333,N_3079);
nand U5584 (N_5584,N_3847,N_2294);
xnor U5585 (N_5585,N_3045,N_3255);
xnor U5586 (N_5586,N_3825,N_3387);
and U5587 (N_5587,N_2316,N_2264);
xnor U5588 (N_5588,N_2862,N_2635);
xor U5589 (N_5589,N_2098,N_3868);
nand U5590 (N_5590,N_3750,N_3360);
nor U5591 (N_5591,N_3792,N_3613);
xnor U5592 (N_5592,N_3685,N_3135);
nand U5593 (N_5593,N_2106,N_2639);
or U5594 (N_5594,N_2681,N_3298);
xnor U5595 (N_5595,N_3884,N_3535);
nor U5596 (N_5596,N_2441,N_2715);
and U5597 (N_5597,N_3651,N_2674);
and U5598 (N_5598,N_2621,N_3139);
nand U5599 (N_5599,N_2834,N_3701);
nor U5600 (N_5600,N_2736,N_3376);
nand U5601 (N_5601,N_2610,N_2068);
nand U5602 (N_5602,N_2864,N_3961);
nand U5603 (N_5603,N_2356,N_3634);
nor U5604 (N_5604,N_3389,N_3192);
xnor U5605 (N_5605,N_3390,N_2333);
and U5606 (N_5606,N_2985,N_3005);
nor U5607 (N_5607,N_2410,N_3746);
or U5608 (N_5608,N_2693,N_2718);
or U5609 (N_5609,N_2194,N_2144);
xor U5610 (N_5610,N_3604,N_2400);
nor U5611 (N_5611,N_3061,N_3436);
or U5612 (N_5612,N_3846,N_3590);
and U5613 (N_5613,N_3944,N_3453);
and U5614 (N_5614,N_2199,N_2121);
and U5615 (N_5615,N_3735,N_3280);
nor U5616 (N_5616,N_2853,N_2430);
or U5617 (N_5617,N_2393,N_3745);
nor U5618 (N_5618,N_3053,N_2430);
or U5619 (N_5619,N_3780,N_2667);
or U5620 (N_5620,N_3424,N_2691);
and U5621 (N_5621,N_2125,N_3433);
nor U5622 (N_5622,N_3930,N_3267);
or U5623 (N_5623,N_2501,N_2221);
xnor U5624 (N_5624,N_3246,N_2322);
nor U5625 (N_5625,N_3386,N_2437);
or U5626 (N_5626,N_3498,N_2128);
or U5627 (N_5627,N_3228,N_3432);
nand U5628 (N_5628,N_2977,N_3763);
nand U5629 (N_5629,N_3358,N_2958);
nor U5630 (N_5630,N_2345,N_3198);
nor U5631 (N_5631,N_3751,N_2006);
nand U5632 (N_5632,N_3977,N_2208);
xor U5633 (N_5633,N_3657,N_3199);
nor U5634 (N_5634,N_2682,N_2475);
nand U5635 (N_5635,N_2796,N_2923);
nand U5636 (N_5636,N_3223,N_2445);
xnor U5637 (N_5637,N_3495,N_3343);
nor U5638 (N_5638,N_3469,N_3049);
nor U5639 (N_5639,N_2666,N_3356);
xnor U5640 (N_5640,N_2169,N_3776);
or U5641 (N_5641,N_3413,N_2754);
nand U5642 (N_5642,N_3948,N_3896);
or U5643 (N_5643,N_3421,N_3926);
nand U5644 (N_5644,N_3882,N_3968);
nor U5645 (N_5645,N_2470,N_2057);
and U5646 (N_5646,N_2989,N_2927);
xor U5647 (N_5647,N_3194,N_3061);
or U5648 (N_5648,N_3424,N_2577);
nand U5649 (N_5649,N_2895,N_2316);
xnor U5650 (N_5650,N_2417,N_2569);
xnor U5651 (N_5651,N_2335,N_3432);
xnor U5652 (N_5652,N_2279,N_2445);
and U5653 (N_5653,N_3883,N_3916);
and U5654 (N_5654,N_3195,N_3290);
xor U5655 (N_5655,N_2151,N_3883);
nor U5656 (N_5656,N_2032,N_2798);
nand U5657 (N_5657,N_2168,N_2634);
and U5658 (N_5658,N_2524,N_2746);
nand U5659 (N_5659,N_3289,N_2258);
or U5660 (N_5660,N_3434,N_2867);
nand U5661 (N_5661,N_3521,N_3972);
nor U5662 (N_5662,N_3921,N_2482);
xor U5663 (N_5663,N_3424,N_2200);
nand U5664 (N_5664,N_2967,N_2366);
nand U5665 (N_5665,N_3225,N_2431);
or U5666 (N_5666,N_3874,N_2026);
nor U5667 (N_5667,N_3583,N_3071);
or U5668 (N_5668,N_3187,N_3226);
nor U5669 (N_5669,N_3140,N_2412);
nand U5670 (N_5670,N_3394,N_3538);
nand U5671 (N_5671,N_2739,N_2516);
nor U5672 (N_5672,N_3906,N_2933);
and U5673 (N_5673,N_3842,N_2911);
nor U5674 (N_5674,N_3364,N_3104);
and U5675 (N_5675,N_3956,N_2162);
and U5676 (N_5676,N_2090,N_3172);
xor U5677 (N_5677,N_2751,N_2843);
nand U5678 (N_5678,N_2260,N_3943);
or U5679 (N_5679,N_3320,N_2477);
nand U5680 (N_5680,N_3614,N_2373);
xnor U5681 (N_5681,N_2716,N_3143);
nor U5682 (N_5682,N_3480,N_3058);
nor U5683 (N_5683,N_3890,N_2491);
xnor U5684 (N_5684,N_3178,N_3535);
xor U5685 (N_5685,N_2852,N_2995);
nor U5686 (N_5686,N_3166,N_2595);
nor U5687 (N_5687,N_2607,N_3411);
and U5688 (N_5688,N_2258,N_3330);
or U5689 (N_5689,N_3155,N_3935);
nand U5690 (N_5690,N_2027,N_3463);
and U5691 (N_5691,N_2385,N_2175);
and U5692 (N_5692,N_3925,N_2347);
and U5693 (N_5693,N_2748,N_3099);
nand U5694 (N_5694,N_2553,N_3628);
and U5695 (N_5695,N_3243,N_2387);
and U5696 (N_5696,N_2087,N_2947);
nor U5697 (N_5697,N_2535,N_3056);
xnor U5698 (N_5698,N_2132,N_2641);
nor U5699 (N_5699,N_3091,N_3350);
xor U5700 (N_5700,N_2548,N_2563);
xnor U5701 (N_5701,N_3872,N_3770);
xor U5702 (N_5702,N_2631,N_3541);
or U5703 (N_5703,N_3769,N_3907);
or U5704 (N_5704,N_2346,N_2611);
or U5705 (N_5705,N_2215,N_2334);
and U5706 (N_5706,N_2258,N_2060);
and U5707 (N_5707,N_3673,N_2059);
xnor U5708 (N_5708,N_3442,N_2412);
and U5709 (N_5709,N_2223,N_2428);
nor U5710 (N_5710,N_3725,N_2678);
xor U5711 (N_5711,N_3500,N_3052);
and U5712 (N_5712,N_3762,N_2190);
or U5713 (N_5713,N_2493,N_3123);
nand U5714 (N_5714,N_3488,N_3701);
or U5715 (N_5715,N_3127,N_3210);
or U5716 (N_5716,N_3430,N_2229);
nor U5717 (N_5717,N_3063,N_2199);
nor U5718 (N_5718,N_2210,N_2054);
or U5719 (N_5719,N_2110,N_3440);
xnor U5720 (N_5720,N_2375,N_2440);
nand U5721 (N_5721,N_2179,N_3693);
xor U5722 (N_5722,N_3862,N_3408);
nand U5723 (N_5723,N_3231,N_3954);
and U5724 (N_5724,N_2906,N_3595);
xnor U5725 (N_5725,N_2058,N_2628);
or U5726 (N_5726,N_2707,N_3635);
nand U5727 (N_5727,N_3954,N_3194);
or U5728 (N_5728,N_2017,N_3541);
and U5729 (N_5729,N_3263,N_3253);
and U5730 (N_5730,N_3248,N_3541);
or U5731 (N_5731,N_3957,N_3261);
nor U5732 (N_5732,N_3236,N_2867);
nor U5733 (N_5733,N_2416,N_3916);
xor U5734 (N_5734,N_3779,N_2539);
or U5735 (N_5735,N_3072,N_3356);
nand U5736 (N_5736,N_3231,N_3323);
or U5737 (N_5737,N_3960,N_3314);
and U5738 (N_5738,N_3166,N_3690);
xor U5739 (N_5739,N_3476,N_3730);
xor U5740 (N_5740,N_3473,N_3860);
or U5741 (N_5741,N_2882,N_2920);
nor U5742 (N_5742,N_3990,N_3537);
or U5743 (N_5743,N_3014,N_3556);
nor U5744 (N_5744,N_2936,N_3451);
xnor U5745 (N_5745,N_3736,N_3409);
xor U5746 (N_5746,N_2308,N_3082);
nor U5747 (N_5747,N_3199,N_2735);
or U5748 (N_5748,N_3591,N_3019);
nand U5749 (N_5749,N_3573,N_3944);
and U5750 (N_5750,N_2845,N_2238);
nor U5751 (N_5751,N_3260,N_2707);
or U5752 (N_5752,N_3311,N_3963);
nor U5753 (N_5753,N_3086,N_2408);
and U5754 (N_5754,N_2956,N_3423);
nand U5755 (N_5755,N_3763,N_3357);
nor U5756 (N_5756,N_3939,N_3582);
and U5757 (N_5757,N_2872,N_3947);
xnor U5758 (N_5758,N_3591,N_3356);
xnor U5759 (N_5759,N_2967,N_3411);
nand U5760 (N_5760,N_3576,N_3641);
and U5761 (N_5761,N_3526,N_3754);
nor U5762 (N_5762,N_3792,N_3279);
xor U5763 (N_5763,N_2875,N_3646);
nor U5764 (N_5764,N_3592,N_2369);
or U5765 (N_5765,N_3477,N_3928);
xor U5766 (N_5766,N_2259,N_3687);
or U5767 (N_5767,N_2143,N_3389);
nor U5768 (N_5768,N_2120,N_2978);
nand U5769 (N_5769,N_3064,N_3560);
xor U5770 (N_5770,N_2879,N_2264);
nor U5771 (N_5771,N_3424,N_3718);
or U5772 (N_5772,N_3944,N_3884);
or U5773 (N_5773,N_3744,N_3039);
xnor U5774 (N_5774,N_2709,N_2821);
xnor U5775 (N_5775,N_3369,N_2484);
nor U5776 (N_5776,N_3877,N_3170);
and U5777 (N_5777,N_2750,N_2264);
xnor U5778 (N_5778,N_3633,N_3520);
xor U5779 (N_5779,N_3483,N_2323);
nor U5780 (N_5780,N_2998,N_3905);
and U5781 (N_5781,N_2561,N_3328);
nor U5782 (N_5782,N_3398,N_3112);
and U5783 (N_5783,N_2949,N_3924);
or U5784 (N_5784,N_2901,N_3814);
and U5785 (N_5785,N_3534,N_3667);
nor U5786 (N_5786,N_3616,N_3635);
nand U5787 (N_5787,N_2177,N_3350);
nand U5788 (N_5788,N_2646,N_2047);
or U5789 (N_5789,N_2715,N_2936);
xnor U5790 (N_5790,N_3024,N_2038);
or U5791 (N_5791,N_2209,N_3914);
nor U5792 (N_5792,N_3178,N_2373);
xor U5793 (N_5793,N_2468,N_2294);
and U5794 (N_5794,N_3310,N_3924);
nand U5795 (N_5795,N_2363,N_3730);
nand U5796 (N_5796,N_3593,N_3620);
xor U5797 (N_5797,N_3668,N_2272);
or U5798 (N_5798,N_2629,N_3048);
or U5799 (N_5799,N_3193,N_3090);
nand U5800 (N_5800,N_3532,N_3762);
xor U5801 (N_5801,N_3843,N_2218);
nand U5802 (N_5802,N_2075,N_2469);
nor U5803 (N_5803,N_3902,N_2644);
or U5804 (N_5804,N_2891,N_2994);
and U5805 (N_5805,N_2717,N_2263);
xnor U5806 (N_5806,N_2131,N_3549);
or U5807 (N_5807,N_3566,N_2857);
and U5808 (N_5808,N_2205,N_2157);
and U5809 (N_5809,N_3845,N_3926);
nor U5810 (N_5810,N_2815,N_2667);
xnor U5811 (N_5811,N_2362,N_2536);
nand U5812 (N_5812,N_2627,N_3443);
and U5813 (N_5813,N_3601,N_2257);
xor U5814 (N_5814,N_2409,N_3368);
or U5815 (N_5815,N_3431,N_2222);
and U5816 (N_5816,N_3042,N_2410);
xnor U5817 (N_5817,N_2455,N_3344);
nand U5818 (N_5818,N_2368,N_3326);
xnor U5819 (N_5819,N_3277,N_2607);
nand U5820 (N_5820,N_2119,N_2445);
nor U5821 (N_5821,N_2942,N_2240);
or U5822 (N_5822,N_2238,N_2182);
nor U5823 (N_5823,N_3924,N_2685);
nand U5824 (N_5824,N_2276,N_2003);
nand U5825 (N_5825,N_3996,N_3186);
or U5826 (N_5826,N_3408,N_2571);
or U5827 (N_5827,N_3861,N_2162);
nor U5828 (N_5828,N_2011,N_3337);
and U5829 (N_5829,N_3489,N_2165);
nand U5830 (N_5830,N_2928,N_3917);
nor U5831 (N_5831,N_2383,N_2396);
nor U5832 (N_5832,N_3205,N_3225);
and U5833 (N_5833,N_2181,N_2333);
and U5834 (N_5834,N_2939,N_2965);
and U5835 (N_5835,N_3534,N_2431);
and U5836 (N_5836,N_2027,N_2251);
nand U5837 (N_5837,N_2400,N_2148);
and U5838 (N_5838,N_3227,N_2299);
xor U5839 (N_5839,N_2360,N_2768);
nand U5840 (N_5840,N_2234,N_2212);
nand U5841 (N_5841,N_3181,N_2349);
xnor U5842 (N_5842,N_3835,N_2662);
or U5843 (N_5843,N_3773,N_2103);
and U5844 (N_5844,N_3966,N_2558);
xnor U5845 (N_5845,N_2912,N_2825);
nor U5846 (N_5846,N_2801,N_3006);
nand U5847 (N_5847,N_2307,N_2517);
nor U5848 (N_5848,N_3781,N_2769);
or U5849 (N_5849,N_3200,N_3672);
nand U5850 (N_5850,N_2835,N_2702);
nand U5851 (N_5851,N_2610,N_3243);
nand U5852 (N_5852,N_3618,N_3451);
and U5853 (N_5853,N_3290,N_2612);
nor U5854 (N_5854,N_3033,N_3945);
or U5855 (N_5855,N_3057,N_2108);
nand U5856 (N_5856,N_3623,N_3705);
nor U5857 (N_5857,N_3060,N_2471);
nand U5858 (N_5858,N_3651,N_3238);
nor U5859 (N_5859,N_2064,N_3097);
or U5860 (N_5860,N_3463,N_3433);
nor U5861 (N_5861,N_3929,N_2223);
nor U5862 (N_5862,N_2901,N_2702);
and U5863 (N_5863,N_3238,N_2242);
xor U5864 (N_5864,N_3503,N_2480);
or U5865 (N_5865,N_3447,N_3255);
and U5866 (N_5866,N_3351,N_2278);
or U5867 (N_5867,N_2367,N_2007);
nand U5868 (N_5868,N_2528,N_3206);
or U5869 (N_5869,N_2527,N_3637);
nor U5870 (N_5870,N_3677,N_2250);
and U5871 (N_5871,N_2464,N_3876);
xor U5872 (N_5872,N_3378,N_3618);
nand U5873 (N_5873,N_3733,N_3729);
and U5874 (N_5874,N_2243,N_3182);
nand U5875 (N_5875,N_3042,N_3033);
or U5876 (N_5876,N_2185,N_2153);
nand U5877 (N_5877,N_3850,N_3183);
and U5878 (N_5878,N_3316,N_2886);
nor U5879 (N_5879,N_2842,N_2282);
xor U5880 (N_5880,N_3221,N_3385);
nand U5881 (N_5881,N_2329,N_3292);
and U5882 (N_5882,N_2870,N_3240);
and U5883 (N_5883,N_3425,N_2497);
nor U5884 (N_5884,N_2633,N_3907);
nor U5885 (N_5885,N_2296,N_2229);
and U5886 (N_5886,N_2669,N_3402);
nand U5887 (N_5887,N_3375,N_2021);
nor U5888 (N_5888,N_2928,N_3868);
nand U5889 (N_5889,N_3851,N_3996);
and U5890 (N_5890,N_2201,N_2718);
nor U5891 (N_5891,N_2845,N_3526);
xnor U5892 (N_5892,N_2057,N_2990);
nand U5893 (N_5893,N_2013,N_3748);
and U5894 (N_5894,N_2381,N_2372);
nor U5895 (N_5895,N_2723,N_3794);
nor U5896 (N_5896,N_2108,N_3978);
nand U5897 (N_5897,N_2030,N_3739);
and U5898 (N_5898,N_3446,N_3513);
xor U5899 (N_5899,N_2265,N_3807);
and U5900 (N_5900,N_2924,N_2256);
or U5901 (N_5901,N_3998,N_2485);
xor U5902 (N_5902,N_3491,N_3220);
and U5903 (N_5903,N_2332,N_2605);
nor U5904 (N_5904,N_2786,N_2963);
or U5905 (N_5905,N_2838,N_3878);
nand U5906 (N_5906,N_2010,N_2875);
or U5907 (N_5907,N_2546,N_3266);
nand U5908 (N_5908,N_2129,N_2234);
xor U5909 (N_5909,N_2456,N_2346);
nand U5910 (N_5910,N_3610,N_3315);
xnor U5911 (N_5911,N_3067,N_3540);
or U5912 (N_5912,N_2007,N_2338);
xor U5913 (N_5913,N_2352,N_2035);
nor U5914 (N_5914,N_3095,N_2847);
or U5915 (N_5915,N_2298,N_2595);
nand U5916 (N_5916,N_3031,N_3186);
and U5917 (N_5917,N_2059,N_2593);
and U5918 (N_5918,N_3988,N_2026);
or U5919 (N_5919,N_2051,N_2634);
xnor U5920 (N_5920,N_3441,N_2267);
xor U5921 (N_5921,N_3969,N_2717);
nor U5922 (N_5922,N_3437,N_2530);
and U5923 (N_5923,N_2972,N_3944);
xor U5924 (N_5924,N_2610,N_2229);
nor U5925 (N_5925,N_3585,N_3932);
nor U5926 (N_5926,N_3226,N_2888);
or U5927 (N_5927,N_2034,N_3051);
nand U5928 (N_5928,N_3248,N_3713);
and U5929 (N_5929,N_2836,N_2317);
and U5930 (N_5930,N_3508,N_2804);
or U5931 (N_5931,N_3080,N_2753);
and U5932 (N_5932,N_3087,N_3579);
or U5933 (N_5933,N_3350,N_3441);
and U5934 (N_5934,N_3025,N_2889);
xnor U5935 (N_5935,N_2811,N_3854);
and U5936 (N_5936,N_2763,N_3997);
nand U5937 (N_5937,N_3048,N_2428);
or U5938 (N_5938,N_2800,N_3199);
or U5939 (N_5939,N_3663,N_3610);
nand U5940 (N_5940,N_2632,N_2692);
nand U5941 (N_5941,N_3029,N_2102);
xor U5942 (N_5942,N_2127,N_3550);
nand U5943 (N_5943,N_3858,N_3656);
or U5944 (N_5944,N_2120,N_2438);
and U5945 (N_5945,N_2637,N_3648);
nand U5946 (N_5946,N_2062,N_2136);
or U5947 (N_5947,N_3660,N_3311);
and U5948 (N_5948,N_3159,N_3519);
or U5949 (N_5949,N_3389,N_2165);
nand U5950 (N_5950,N_2447,N_3523);
or U5951 (N_5951,N_2555,N_2838);
nor U5952 (N_5952,N_2477,N_2527);
xor U5953 (N_5953,N_3006,N_3306);
and U5954 (N_5954,N_3351,N_3624);
nand U5955 (N_5955,N_2568,N_2914);
xnor U5956 (N_5956,N_3326,N_3350);
and U5957 (N_5957,N_3656,N_2320);
or U5958 (N_5958,N_2432,N_2692);
nor U5959 (N_5959,N_2679,N_3047);
xnor U5960 (N_5960,N_3424,N_3244);
and U5961 (N_5961,N_3340,N_3745);
nand U5962 (N_5962,N_2273,N_2272);
or U5963 (N_5963,N_2942,N_2419);
and U5964 (N_5964,N_2945,N_2552);
and U5965 (N_5965,N_3752,N_3978);
xnor U5966 (N_5966,N_2280,N_3146);
xnor U5967 (N_5967,N_2778,N_3618);
xnor U5968 (N_5968,N_3740,N_2268);
nand U5969 (N_5969,N_2535,N_2853);
or U5970 (N_5970,N_2083,N_3304);
xor U5971 (N_5971,N_2428,N_2588);
nand U5972 (N_5972,N_2242,N_3322);
xnor U5973 (N_5973,N_3080,N_3783);
nand U5974 (N_5974,N_2610,N_2046);
nor U5975 (N_5975,N_3627,N_3920);
or U5976 (N_5976,N_3116,N_2864);
nor U5977 (N_5977,N_3287,N_3578);
nor U5978 (N_5978,N_3809,N_2071);
and U5979 (N_5979,N_3382,N_3087);
nor U5980 (N_5980,N_3632,N_2614);
nand U5981 (N_5981,N_2819,N_3063);
nand U5982 (N_5982,N_3621,N_3652);
nand U5983 (N_5983,N_2226,N_2830);
or U5984 (N_5984,N_3102,N_2491);
and U5985 (N_5985,N_3697,N_2877);
nor U5986 (N_5986,N_3075,N_2691);
nand U5987 (N_5987,N_2784,N_3055);
nand U5988 (N_5988,N_3634,N_3557);
xor U5989 (N_5989,N_3881,N_2556);
or U5990 (N_5990,N_3149,N_3989);
xnor U5991 (N_5991,N_2342,N_3135);
or U5992 (N_5992,N_3774,N_3704);
and U5993 (N_5993,N_2216,N_2733);
nor U5994 (N_5994,N_2400,N_2343);
nand U5995 (N_5995,N_2570,N_3273);
nand U5996 (N_5996,N_3622,N_3893);
and U5997 (N_5997,N_3679,N_3231);
or U5998 (N_5998,N_3814,N_2393);
nand U5999 (N_5999,N_3771,N_3749);
or U6000 (N_6000,N_5598,N_4344);
nand U6001 (N_6001,N_4398,N_5852);
and U6002 (N_6002,N_5384,N_5758);
nand U6003 (N_6003,N_4973,N_4374);
or U6004 (N_6004,N_5222,N_4386);
and U6005 (N_6005,N_5670,N_5367);
xnor U6006 (N_6006,N_4888,N_5545);
nor U6007 (N_6007,N_4443,N_5233);
or U6008 (N_6008,N_4372,N_4106);
nor U6009 (N_6009,N_5812,N_5908);
and U6010 (N_6010,N_5606,N_5848);
nor U6011 (N_6011,N_4284,N_4307);
nor U6012 (N_6012,N_4606,N_5743);
nand U6013 (N_6013,N_4167,N_4590);
xor U6014 (N_6014,N_4485,N_5712);
xor U6015 (N_6015,N_4038,N_5491);
and U6016 (N_6016,N_4879,N_5085);
nor U6017 (N_6017,N_4423,N_5786);
nand U6018 (N_6018,N_5548,N_4325);
nand U6019 (N_6019,N_5292,N_4717);
xnor U6020 (N_6020,N_5637,N_4548);
or U6021 (N_6021,N_5087,N_5223);
nand U6022 (N_6022,N_5439,N_5977);
nor U6023 (N_6023,N_4122,N_4708);
nand U6024 (N_6024,N_4475,N_4225);
nand U6025 (N_6025,N_4319,N_5710);
or U6026 (N_6026,N_4088,N_5215);
nand U6027 (N_6027,N_4880,N_4781);
or U6028 (N_6028,N_5171,N_5132);
or U6029 (N_6029,N_4632,N_4745);
nor U6030 (N_6030,N_4896,N_4951);
xnor U6031 (N_6031,N_5892,N_4360);
or U6032 (N_6032,N_4193,N_4124);
and U6033 (N_6033,N_5399,N_5493);
or U6034 (N_6034,N_5285,N_5723);
nand U6035 (N_6035,N_5953,N_4634);
nor U6036 (N_6036,N_5414,N_4407);
nor U6037 (N_6037,N_4181,N_5949);
nand U6038 (N_6038,N_4388,N_4601);
or U6039 (N_6039,N_5027,N_4459);
and U6040 (N_6040,N_5785,N_5463);
or U6041 (N_6041,N_4927,N_5473);
nor U6042 (N_6042,N_4474,N_5058);
nand U6043 (N_6043,N_5377,N_4151);
and U6044 (N_6044,N_4988,N_5960);
nand U6045 (N_6045,N_4022,N_5555);
nor U6046 (N_6046,N_4529,N_4652);
or U6047 (N_6047,N_4435,N_5189);
xnor U6048 (N_6048,N_5693,N_5331);
and U6049 (N_6049,N_5921,N_4686);
nand U6050 (N_6050,N_5826,N_4065);
and U6051 (N_6051,N_5366,N_4889);
nand U6052 (N_6052,N_5795,N_4073);
nand U6053 (N_6053,N_5666,N_5247);
nor U6054 (N_6054,N_5181,N_5318);
nor U6055 (N_6055,N_5336,N_5602);
and U6056 (N_6056,N_4299,N_4539);
and U6057 (N_6057,N_5654,N_5824);
nand U6058 (N_6058,N_5457,N_5640);
or U6059 (N_6059,N_4148,N_4513);
xor U6060 (N_6060,N_4293,N_4046);
and U6061 (N_6061,N_4123,N_5748);
nor U6062 (N_6062,N_5459,N_5527);
nor U6063 (N_6063,N_4859,N_4204);
nor U6064 (N_6064,N_5154,N_5356);
xor U6065 (N_6065,N_5311,N_4570);
xnor U6066 (N_6066,N_5579,N_5387);
nor U6067 (N_6067,N_4010,N_5680);
or U6068 (N_6068,N_4800,N_4843);
and U6069 (N_6069,N_4137,N_5832);
or U6070 (N_6070,N_5220,N_5102);
and U6071 (N_6071,N_5009,N_4827);
or U6072 (N_6072,N_5252,N_5343);
and U6073 (N_6073,N_4092,N_4401);
or U6074 (N_6074,N_4807,N_5095);
and U6075 (N_6075,N_4466,N_4075);
nand U6076 (N_6076,N_5300,N_4791);
and U6077 (N_6077,N_5590,N_5264);
nor U6078 (N_6078,N_4817,N_4957);
nor U6079 (N_6079,N_4471,N_4554);
nor U6080 (N_6080,N_4308,N_5057);
nand U6081 (N_6081,N_5008,N_4503);
and U6082 (N_6082,N_5043,N_5665);
xor U6083 (N_6083,N_5747,N_5822);
and U6084 (N_6084,N_5973,N_5557);
and U6085 (N_6085,N_4077,N_4300);
or U6086 (N_6086,N_4079,N_5185);
xnor U6087 (N_6087,N_4239,N_5787);
xnor U6088 (N_6088,N_4107,N_5914);
nor U6089 (N_6089,N_5565,N_5141);
nor U6090 (N_6090,N_5597,N_4150);
or U6091 (N_6091,N_5583,N_5188);
nand U6092 (N_6092,N_5304,N_5989);
and U6093 (N_6093,N_5794,N_4187);
or U6094 (N_6094,N_4567,N_4014);
or U6095 (N_6095,N_4937,N_5775);
nor U6096 (N_6096,N_4602,N_4874);
xnor U6097 (N_6097,N_4694,N_5066);
nor U6098 (N_6098,N_4695,N_4909);
xnor U6099 (N_6099,N_5350,N_5465);
or U6100 (N_6100,N_4805,N_5175);
or U6101 (N_6101,N_4858,N_5005);
xnor U6102 (N_6102,N_5742,N_4796);
nor U6103 (N_6103,N_5445,N_5307);
xor U6104 (N_6104,N_4061,N_4960);
xor U6105 (N_6105,N_5950,N_4517);
nand U6106 (N_6106,N_5599,N_5289);
nor U6107 (N_6107,N_4507,N_4778);
nor U6108 (N_6108,N_4354,N_5418);
nor U6109 (N_6109,N_4774,N_5561);
or U6110 (N_6110,N_4835,N_5642);
xnor U6111 (N_6111,N_4076,N_4623);
or U6112 (N_6112,N_5047,N_4478);
nor U6113 (N_6113,N_5969,N_4387);
and U6114 (N_6114,N_5090,N_4560);
or U6115 (N_6115,N_4921,N_5684);
or U6116 (N_6116,N_4954,N_4565);
or U6117 (N_6117,N_4406,N_4950);
xnor U6118 (N_6118,N_4631,N_4058);
and U6119 (N_6119,N_5803,N_5297);
or U6120 (N_6120,N_5814,N_5338);
and U6121 (N_6121,N_4460,N_4506);
and U6122 (N_6122,N_5923,N_5487);
and U6123 (N_6123,N_5653,N_4218);
nor U6124 (N_6124,N_5157,N_4613);
and U6125 (N_6125,N_5481,N_4649);
nor U6126 (N_6126,N_4380,N_5595);
or U6127 (N_6127,N_5616,N_4655);
xor U6128 (N_6128,N_4233,N_5326);
nand U6129 (N_6129,N_5046,N_4078);
nand U6130 (N_6130,N_4002,N_4057);
nor U6131 (N_6131,N_5959,N_4765);
nand U6132 (N_6132,N_5104,N_5455);
xnor U6133 (N_6133,N_4861,N_4208);
and U6134 (N_6134,N_5919,N_4168);
nor U6135 (N_6135,N_4256,N_5070);
xnor U6136 (N_6136,N_4108,N_5206);
or U6137 (N_6137,N_4165,N_4339);
and U6138 (N_6138,N_5735,N_5869);
nand U6139 (N_6139,N_5641,N_5627);
xnor U6140 (N_6140,N_5408,N_4039);
nand U6141 (N_6141,N_4531,N_5855);
nand U6142 (N_6142,N_4666,N_4821);
xor U6143 (N_6143,N_4100,N_4579);
and U6144 (N_6144,N_4047,N_4183);
nor U6145 (N_6145,N_5987,N_5249);
nand U6146 (N_6146,N_5886,N_5131);
nor U6147 (N_6147,N_5781,N_5495);
and U6148 (N_6148,N_5127,N_5450);
and U6149 (N_6149,N_5738,N_5081);
nor U6150 (N_6150,N_5879,N_5155);
xor U6151 (N_6151,N_5346,N_5715);
nand U6152 (N_6152,N_4793,N_5514);
or U6153 (N_6153,N_5248,N_5353);
and U6154 (N_6154,N_4628,N_4509);
xor U6155 (N_6155,N_5902,N_5239);
xor U6156 (N_6156,N_4847,N_5807);
or U6157 (N_6157,N_5327,N_4510);
xnor U6158 (N_6158,N_4671,N_5759);
nor U6159 (N_6159,N_4312,N_5357);
and U6160 (N_6160,N_5745,N_5065);
and U6161 (N_6161,N_4865,N_5394);
xor U6162 (N_6162,N_5900,N_4878);
xor U6163 (N_6163,N_4673,N_4170);
and U6164 (N_6164,N_5881,N_5701);
nand U6165 (N_6165,N_5925,N_5490);
or U6166 (N_6166,N_4001,N_5773);
or U6167 (N_6167,N_4958,N_4886);
xor U6168 (N_6168,N_4274,N_4820);
nor U6169 (N_6169,N_5934,N_4259);
and U6170 (N_6170,N_5867,N_4241);
nor U6171 (N_6171,N_4715,N_5093);
or U6172 (N_6172,N_4409,N_4779);
nor U6173 (N_6173,N_4953,N_5101);
and U6174 (N_6174,N_5591,N_5898);
nand U6175 (N_6175,N_5732,N_5604);
nand U6176 (N_6176,N_4003,N_5859);
nand U6177 (N_6177,N_4147,N_4253);
nand U6178 (N_6178,N_5204,N_5755);
and U6179 (N_6179,N_5731,N_5038);
or U6180 (N_6180,N_4236,N_4157);
or U6181 (N_6181,N_5099,N_4521);
or U6182 (N_6182,N_4213,N_5880);
nor U6183 (N_6183,N_5507,N_5592);
nand U6184 (N_6184,N_5619,N_5303);
and U6185 (N_6185,N_4610,N_4191);
and U6186 (N_6186,N_4426,N_5720);
or U6187 (N_6187,N_4452,N_5169);
xor U6188 (N_6188,N_4670,N_4752);
and U6189 (N_6189,N_4195,N_4205);
and U6190 (N_6190,N_5910,N_5431);
nand U6191 (N_6191,N_5333,N_5655);
nor U6192 (N_6192,N_4904,N_5737);
nor U6193 (N_6193,N_5402,N_4557);
and U6194 (N_6194,N_4334,N_4172);
or U6195 (N_6195,N_5846,N_4357);
nand U6196 (N_6196,N_4371,N_4592);
nor U6197 (N_6197,N_4782,N_5649);
nand U6198 (N_6198,N_4598,N_5757);
xnor U6199 (N_6199,N_5623,N_5480);
nor U6200 (N_6200,N_4023,N_4365);
nor U6201 (N_6201,N_5505,N_5632);
or U6202 (N_6202,N_5643,N_5179);
nand U6203 (N_6203,N_4021,N_5834);
nand U6204 (N_6204,N_4737,N_5161);
nor U6205 (N_6205,N_5504,N_4411);
or U6206 (N_6206,N_4007,N_5906);
nor U6207 (N_6207,N_4445,N_4441);
or U6208 (N_6208,N_5412,N_5518);
and U6209 (N_6209,N_4599,N_5612);
nand U6210 (N_6210,N_5443,N_5589);
and U6211 (N_6211,N_5714,N_4709);
xor U6212 (N_6212,N_4101,N_5875);
or U6213 (N_6213,N_5593,N_4081);
xor U6214 (N_6214,N_4650,N_4134);
xor U6215 (N_6215,N_4373,N_4989);
nand U6216 (N_6216,N_5603,N_4250);
xor U6217 (N_6217,N_4713,N_4784);
or U6218 (N_6218,N_5993,N_4449);
or U6219 (N_6219,N_5177,N_4786);
and U6220 (N_6220,N_4635,N_5837);
xor U6221 (N_6221,N_5767,N_4564);
xor U6222 (N_6222,N_5485,N_4875);
xor U6223 (N_6223,N_4056,N_5139);
xnor U6224 (N_6224,N_5678,N_4285);
or U6225 (N_6225,N_4468,N_4015);
nor U6226 (N_6226,N_4050,N_4918);
and U6227 (N_6227,N_5531,N_4384);
nor U6228 (N_6228,N_5411,N_5254);
xnor U6229 (N_6229,N_4645,N_4550);
nand U6230 (N_6230,N_5113,N_5424);
xnor U6231 (N_6231,N_5585,N_4389);
nand U6232 (N_6232,N_4359,N_5309);
xor U6233 (N_6233,N_5976,N_5268);
and U6234 (N_6234,N_4866,N_5250);
or U6235 (N_6235,N_4586,N_4219);
nand U6236 (N_6236,N_4646,N_5920);
nor U6237 (N_6237,N_5392,N_4524);
and U6238 (N_6238,N_4029,N_4366);
and U6239 (N_6239,N_5668,N_4229);
and U6240 (N_6240,N_5274,N_5153);
and U6241 (N_6241,N_5075,N_4254);
or U6242 (N_6242,N_4566,N_4526);
nand U6243 (N_6243,N_5174,N_4622);
and U6244 (N_6244,N_5282,N_5429);
nand U6245 (N_6245,N_4146,N_4493);
nor U6246 (N_6246,N_5526,N_4145);
xor U6247 (N_6247,N_5051,N_4910);
nand U6248 (N_6248,N_5551,N_4026);
xnor U6249 (N_6249,N_4757,N_5744);
or U6250 (N_6250,N_5776,N_4573);
nor U6251 (N_6251,N_4541,N_4447);
or U6252 (N_6252,N_4690,N_4643);
nand U6253 (N_6253,N_5705,N_5946);
nor U6254 (N_6254,N_5314,N_5486);
nor U6255 (N_6255,N_5516,N_5479);
and U6256 (N_6256,N_4260,N_4223);
xor U6257 (N_6257,N_4094,N_5582);
and U6258 (N_6258,N_5352,N_5797);
nand U6259 (N_6259,N_4965,N_4648);
and U6260 (N_6260,N_4802,N_4928);
or U6261 (N_6261,N_4346,N_5286);
and U6262 (N_6262,N_5349,N_5226);
and U6263 (N_6263,N_4956,N_4248);
xnor U6264 (N_6264,N_4916,N_5928);
or U6265 (N_6265,N_4900,N_4385);
and U6266 (N_6266,N_5629,N_4399);
and U6267 (N_6267,N_4846,N_4390);
nor U6268 (N_6268,N_5260,N_4131);
nand U6269 (N_6269,N_4818,N_4055);
nor U6270 (N_6270,N_4221,N_5947);
or U6271 (N_6271,N_4922,N_5792);
nand U6272 (N_6272,N_4551,N_4759);
and U6273 (N_6273,N_5584,N_5194);
xor U6274 (N_6274,N_4328,N_5446);
nand U6275 (N_6275,N_4948,N_4587);
xor U6276 (N_6276,N_4016,N_4139);
and U6277 (N_6277,N_5427,N_5793);
and U6278 (N_6278,N_5615,N_5419);
nand U6279 (N_6279,N_5508,N_5148);
nor U6280 (N_6280,N_4701,N_4505);
and U6281 (N_6281,N_4605,N_4841);
and U6282 (N_6282,N_4895,N_5217);
or U6283 (N_6283,N_4281,N_5689);
nor U6284 (N_6284,N_5676,N_4637);
or U6285 (N_6285,N_4495,N_4196);
or U6286 (N_6286,N_4615,N_5151);
or U6287 (N_6287,N_4331,N_4060);
and U6288 (N_6288,N_5108,N_4395);
or U6289 (N_6289,N_4450,N_4104);
and U6290 (N_6290,N_5765,N_4391);
and U6291 (N_6291,N_4885,N_5319);
nand U6292 (N_6292,N_4159,N_4314);
xnor U6293 (N_6293,N_5277,N_4642);
xnor U6294 (N_6294,N_4271,N_5860);
nand U6295 (N_6295,N_4591,N_5556);
xnor U6296 (N_6296,N_5497,N_4034);
and U6297 (N_6297,N_5853,N_4549);
nand U6298 (N_6298,N_4589,N_5238);
nor U6299 (N_6299,N_5897,N_4762);
nand U6300 (N_6300,N_5760,N_4864);
nand U6301 (N_6301,N_4349,N_5883);
and U6302 (N_6302,N_4947,N_5625);
nor U6303 (N_6303,N_5240,N_4045);
nand U6304 (N_6304,N_5305,N_5064);
xor U6305 (N_6305,N_4404,N_4982);
or U6306 (N_6306,N_5230,N_4035);
nor U6307 (N_6307,N_4053,N_5729);
or U6308 (N_6308,N_4934,N_4898);
nand U6309 (N_6309,N_5173,N_4358);
nor U6310 (N_6310,N_5076,N_4899);
xor U6311 (N_6311,N_4659,N_5752);
nand U6312 (N_6312,N_4534,N_5060);
xor U6313 (N_6313,N_5638,N_4091);
nor U6314 (N_6314,N_4264,N_5961);
nor U6315 (N_6315,N_5052,N_5607);
nor U6316 (N_6316,N_5498,N_5287);
xnor U6317 (N_6317,N_5972,N_5894);
nand U6318 (N_6318,N_4863,N_5661);
or U6319 (N_6319,N_4877,N_5614);
and U6320 (N_6320,N_5187,N_4189);
nand U6321 (N_6321,N_4267,N_4336);
nor U6322 (N_6322,N_5454,N_5214);
and U6323 (N_6323,N_4066,N_5513);
or U6324 (N_6324,N_4665,N_5954);
nand U6325 (N_6325,N_5610,N_4929);
or U6326 (N_6326,N_5725,N_4719);
nand U6327 (N_6327,N_5422,N_4356);
nor U6328 (N_6328,N_4532,N_4855);
nand U6329 (N_6329,N_4318,N_5779);
xor U6330 (N_6330,N_5466,N_5523);
and U6331 (N_6331,N_5324,N_4559);
or U6332 (N_6332,N_5764,N_4674);
nor U6333 (N_6333,N_4905,N_4188);
nor U6334 (N_6334,N_4240,N_4683);
nand U6335 (N_6335,N_5932,N_5717);
and U6336 (N_6336,N_4825,N_5761);
nor U6337 (N_6337,N_5313,N_5207);
nand U6338 (N_6338,N_4540,N_4574);
nor U6339 (N_6339,N_5166,N_4296);
nand U6340 (N_6340,N_4099,N_4603);
nand U6341 (N_6341,N_4873,N_5975);
xnor U6342 (N_6342,N_4987,N_5109);
xnor U6343 (N_6343,N_5810,N_4000);
xnor U6344 (N_6344,N_5484,N_4154);
or U6345 (N_6345,N_4942,N_5017);
or U6346 (N_6346,N_5780,N_5503);
nand U6347 (N_6347,N_4477,N_5915);
or U6348 (N_6348,N_4836,N_4804);
xnor U6349 (N_6349,N_4920,N_5694);
nor U6350 (N_6350,N_4490,N_5964);
and U6351 (N_6351,N_5209,N_5393);
nor U6352 (N_6352,N_4114,N_5007);
xor U6353 (N_6353,N_5295,N_4127);
or U6354 (N_6354,N_4402,N_5084);
xnor U6355 (N_6355,N_5296,N_5626);
or U6356 (N_6356,N_5586,N_4883);
nor U6357 (N_6357,N_4464,N_5682);
nand U6358 (N_6358,N_4935,N_4446);
xor U6359 (N_6359,N_5372,N_4033);
nor U6360 (N_6360,N_5415,N_5576);
xnor U6361 (N_6361,N_4892,N_4860);
xor U6362 (N_6362,N_4235,N_4330);
or U6363 (N_6363,N_4983,N_4180);
xnor U6364 (N_6364,N_5325,N_4608);
nor U6365 (N_6365,N_4097,N_4522);
nor U6366 (N_6366,N_4943,N_4311);
nor U6367 (N_6367,N_5140,N_4611);
and U6368 (N_6368,N_4292,N_4041);
nor U6369 (N_6369,N_4710,N_4993);
xnor U6370 (N_6370,N_4068,N_4578);
nor U6371 (N_6371,N_4681,N_4417);
or U6372 (N_6372,N_5578,N_4201);
xnor U6373 (N_6373,N_4162,N_5094);
or U6374 (N_6374,N_4184,N_5063);
or U6375 (N_6375,N_5142,N_5143);
xor U6376 (N_6376,N_5145,N_5144);
nor U6377 (N_6377,N_4499,N_5650);
nor U6378 (N_6378,N_4383,N_5534);
nor U6379 (N_6379,N_5957,N_4777);
nor U6380 (N_6380,N_5730,N_5002);
and U6381 (N_6381,N_4764,N_4103);
nand U6382 (N_6382,N_4906,N_5951);
and U6383 (N_6383,N_5492,N_4164);
and U6384 (N_6384,N_5294,N_5933);
xnor U6385 (N_6385,N_5202,N_4721);
nor U6386 (N_6386,N_5992,N_5191);
or U6387 (N_6387,N_4216,N_4555);
and U6388 (N_6388,N_5137,N_5817);
nor U6389 (N_6389,N_5111,N_4457);
xor U6390 (N_6390,N_4845,N_4552);
nand U6391 (N_6391,N_5687,N_5819);
nand U6392 (N_6392,N_4706,N_4209);
nor U6393 (N_6393,N_5835,N_4742);
or U6394 (N_6394,N_5112,N_4743);
and U6395 (N_6395,N_5509,N_5100);
nor U6396 (N_6396,N_4850,N_5373);
nor U6397 (N_6397,N_4451,N_4854);
xor U6398 (N_6398,N_4381,N_5857);
nand U6399 (N_6399,N_4758,N_5736);
or U6400 (N_6400,N_5494,N_4276);
nor U6401 (N_6401,N_5351,N_4031);
or U6402 (N_6402,N_4771,N_5044);
nor U6403 (N_6403,N_5432,N_5211);
nor U6404 (N_6404,N_4588,N_4469);
and U6405 (N_6405,N_5726,N_5955);
nor U6406 (N_6406,N_4072,N_4089);
and U6407 (N_6407,N_5647,N_5259);
xor U6408 (N_6408,N_5012,N_5121);
nand U6409 (N_6409,N_4620,N_5554);
nand U6410 (N_6410,N_4027,N_4305);
nand U6411 (N_6411,N_5227,N_4273);
or U6412 (N_6412,N_4699,N_5524);
xnor U6413 (N_6413,N_5078,N_5255);
nand U6414 (N_6414,N_4621,N_4115);
nor U6415 (N_6415,N_5091,N_5839);
xor U6416 (N_6416,N_4370,N_5462);
nor U6417 (N_6417,N_5437,N_5088);
xnor U6418 (N_6418,N_5567,N_4364);
nand U6419 (N_6419,N_4849,N_5850);
nor U6420 (N_6420,N_5984,N_4268);
nor U6421 (N_6421,N_4138,N_4961);
or U6422 (N_6422,N_4907,N_4261);
or U6423 (N_6423,N_5231,N_4707);
or U6424 (N_6424,N_5673,N_5952);
xor U6425 (N_6425,N_5219,N_4030);
nor U6426 (N_6426,N_4838,N_4975);
xnor U6427 (N_6427,N_4672,N_4790);
xnor U6428 (N_6428,N_5659,N_4814);
and U6429 (N_6429,N_5522,N_4819);
nor U6430 (N_6430,N_5045,N_4569);
or U6431 (N_6431,N_5257,N_4856);
nand U6432 (N_6432,N_5341,N_5434);
nor U6433 (N_6433,N_5050,N_5036);
xnor U6434 (N_6434,N_4350,N_4977);
nand U6435 (N_6435,N_5677,N_5213);
and U6436 (N_6436,N_5067,N_5172);
and U6437 (N_6437,N_5389,N_4470);
nand U6438 (N_6438,N_5895,N_4355);
nor U6439 (N_6439,N_4840,N_5072);
or U6440 (N_6440,N_5608,N_4004);
xor U6441 (N_6441,N_4959,N_4738);
or U6442 (N_6442,N_4282,N_4442);
and U6443 (N_6443,N_4787,N_4322);
and U6444 (N_6444,N_4177,N_4941);
nand U6445 (N_6445,N_5929,N_4454);
nand U6446 (N_6446,N_5994,N_5329);
nand U6447 (N_6447,N_5059,N_5083);
and U6448 (N_6448,N_4182,N_5577);
nor U6449 (N_6449,N_5438,N_5916);
nor U6450 (N_6450,N_4249,N_5651);
nor U6451 (N_6451,N_5444,N_5164);
and U6452 (N_6452,N_4171,N_5974);
and U6453 (N_6453,N_5026,N_5733);
and U6454 (N_6454,N_4734,N_5266);
nor U6455 (N_6455,N_5532,N_4582);
and U6456 (N_6456,N_5448,N_5472);
nand U6457 (N_6457,N_4577,N_4367);
or U6458 (N_6458,N_4712,N_4636);
xnor U6459 (N_6459,N_4152,N_5703);
and U6460 (N_6460,N_4669,N_4161);
or U6461 (N_6461,N_4834,N_4735);
or U6462 (N_6462,N_4119,N_5195);
nor U6463 (N_6463,N_4071,N_4246);
xor U6464 (N_6464,N_5048,N_5711);
nor U6465 (N_6465,N_5447,N_5671);
nor U6466 (N_6466,N_5115,N_5339);
and U6467 (N_6467,N_4563,N_5724);
and U6468 (N_6468,N_5858,N_5010);
or U6469 (N_6469,N_5288,N_4530);
and U6470 (N_6470,N_5862,N_5281);
nand U6471 (N_6471,N_5727,N_5284);
nor U6472 (N_6472,N_5097,N_4017);
or U6473 (N_6473,N_4095,N_4396);
nor U6474 (N_6474,N_4190,N_5125);
nand U6475 (N_6475,N_4265,N_5362);
or U6476 (N_6476,N_4739,N_4867);
xor U6477 (N_6477,N_5193,N_4294);
and U6478 (N_6478,N_4730,N_5924);
nand U6479 (N_6479,N_4986,N_5105);
or U6480 (N_6480,N_4220,N_4090);
nand U6481 (N_6481,N_5901,N_4726);
xnor U6482 (N_6482,N_4085,N_4897);
xnor U6483 (N_6483,N_5381,N_4985);
nand U6484 (N_6484,N_4111,N_4397);
xor U6485 (N_6485,N_5499,N_4420);
and U6486 (N_6486,N_5369,N_4340);
nor U6487 (N_6487,N_5089,N_4310);
nand U6488 (N_6488,N_4142,N_5594);
or U6489 (N_6489,N_5315,N_4479);
xnor U6490 (N_6490,N_4317,N_4826);
nor U6491 (N_6491,N_5079,N_5749);
xor U6492 (N_6492,N_5865,N_5945);
nand U6493 (N_6493,N_5778,N_4212);
and U6494 (N_6494,N_4964,N_5833);
or U6495 (N_6495,N_5011,N_4062);
and U6496 (N_6496,N_4658,N_5836);
or U6497 (N_6497,N_5184,N_5512);
xnor U6498 (N_6498,N_4044,N_4337);
and U6499 (N_6499,N_5679,N_5103);
nor U6500 (N_6500,N_5278,N_4298);
nand U6501 (N_6501,N_4093,N_5134);
nand U6502 (N_6502,N_4705,N_4178);
or U6503 (N_6503,N_4118,N_5396);
nor U6504 (N_6504,N_5205,N_5672);
nor U6505 (N_6505,N_5871,N_5383);
or U6506 (N_6506,N_5500,N_4996);
xnor U6507 (N_6507,N_5956,N_4616);
xor U6508 (N_6508,N_5192,N_5937);
nand U6509 (N_6509,N_4512,N_5800);
or U6510 (N_6510,N_4732,N_5681);
xnor U6511 (N_6511,N_4837,N_4084);
or U6512 (N_6512,N_4801,N_5575);
nor U6513 (N_6513,N_4174,N_4237);
and U6514 (N_6514,N_4222,N_5275);
nor U6515 (N_6515,N_5163,N_5868);
nor U6516 (N_6516,N_4629,N_4911);
xnor U6517 (N_6517,N_5520,N_4067);
xor U6518 (N_6518,N_5634,N_4215);
xnor U6519 (N_6519,N_4514,N_4908);
nor U6520 (N_6520,N_4932,N_4403);
or U6521 (N_6521,N_5197,N_5496);
xor U6522 (N_6522,N_5533,N_4881);
and U6523 (N_6523,N_5293,N_5660);
nor U6524 (N_6524,N_4963,N_4244);
or U6525 (N_6525,N_5430,N_5361);
and U6526 (N_6526,N_5943,N_4919);
xor U6527 (N_6527,N_5147,N_4461);
nor U6528 (N_6528,N_5872,N_5664);
or U6529 (N_6529,N_5918,N_5573);
or U6530 (N_6530,N_4362,N_4585);
or U6531 (N_6531,N_4553,N_4680);
or U6532 (N_6532,N_5829,N_4422);
and U6533 (N_6533,N_4481,N_5323);
xnor U6534 (N_6534,N_5692,N_5119);
or U6535 (N_6535,N_5998,N_5400);
and U6536 (N_6536,N_4824,N_5136);
xnor U6537 (N_6537,N_5863,N_5080);
or U6538 (N_6538,N_4025,N_5306);
xnor U6539 (N_6539,N_5543,N_4272);
or U6540 (N_6540,N_4394,N_4851);
and U6541 (N_6541,N_5098,N_5613);
nand U6542 (N_6542,N_4525,N_5229);
nand U6543 (N_6543,N_5037,N_4200);
and U6544 (N_6544,N_5410,N_5967);
xor U6545 (N_6545,N_4756,N_4121);
and U6546 (N_6546,N_5830,N_4789);
and U6547 (N_6547,N_4704,N_4775);
nor U6548 (N_6548,N_4795,N_5340);
nor U6549 (N_6549,N_5821,N_5788);
or U6550 (N_6550,N_4995,N_4326);
xor U6551 (N_6551,N_5873,N_5605);
nor U6552 (N_6552,N_4832,N_5645);
or U6553 (N_6553,N_5034,N_4698);
nor U6554 (N_6554,N_4811,N_5310);
xnor U6555 (N_6555,N_5506,N_5489);
nor U6556 (N_6556,N_4087,N_5911);
and U6557 (N_6557,N_4915,N_5851);
or U6558 (N_6558,N_5907,N_4316);
nand U6559 (N_6559,N_5146,N_5790);
nand U6560 (N_6560,N_5917,N_4657);
xnor U6561 (N_6561,N_5170,N_4537);
or U6562 (N_6562,N_5734,N_5417);
and U6563 (N_6563,N_5633,N_4833);
or U6564 (N_6564,N_4747,N_4277);
nor U6565 (N_6565,N_5267,N_5805);
nor U6566 (N_6566,N_4153,N_5801);
nand U6567 (N_6567,N_5363,N_5013);
xor U6568 (N_6568,N_5225,N_5882);
nand U6569 (N_6569,N_4970,N_4809);
nand U6570 (N_6570,N_4969,N_5842);
xor U6571 (N_6571,N_4810,N_5849);
xor U6572 (N_6572,N_5887,N_4803);
and U6573 (N_6573,N_4562,N_5662);
or U6574 (N_6574,N_4315,N_5423);
nand U6575 (N_6575,N_5476,N_4348);
and U6576 (N_6576,N_5241,N_4823);
and U6577 (N_6577,N_4206,N_4500);
xor U6578 (N_6578,N_4207,N_5798);
and U6579 (N_6579,N_4379,N_4231);
xnor U6580 (N_6580,N_4491,N_4321);
nor U6581 (N_6581,N_5129,N_4247);
or U6582 (N_6582,N_5451,N_5452);
nand U6583 (N_6583,N_5117,N_5203);
xnor U6584 (N_6584,N_4519,N_5018);
and U6585 (N_6585,N_5212,N_4763);
or U6586 (N_6586,N_4158,N_4971);
and U6587 (N_6587,N_5789,N_5978);
and U6588 (N_6588,N_5547,N_4685);
xnor U6589 (N_6589,N_4080,N_5263);
and U6590 (N_6590,N_5840,N_4893);
or U6591 (N_6591,N_4375,N_5110);
nand U6592 (N_6592,N_5421,N_4301);
and U6593 (N_6593,N_5237,N_5467);
nor U6594 (N_6594,N_5667,N_5990);
and U6595 (N_6595,N_5905,N_4117);
or U6596 (N_6596,N_4746,N_4439);
or U6597 (N_6597,N_5611,N_5864);
nor U6598 (N_6598,N_4533,N_5966);
and U6599 (N_6599,N_5847,N_4728);
and U6600 (N_6600,N_4211,N_4999);
xor U6601 (N_6601,N_5460,N_5944);
nor U6602 (N_6602,N_4270,N_4320);
nor U6603 (N_6603,N_4160,N_5983);
xor U6604 (N_6604,N_4917,N_4304);
nor U6605 (N_6605,N_5030,N_4926);
or U6606 (N_6606,N_5409,N_5149);
or U6607 (N_6607,N_5630,N_5831);
xor U6608 (N_6608,N_4465,N_5020);
nand U6609 (N_6609,N_5553,N_5804);
and U6610 (N_6610,N_4703,N_5563);
nand U6611 (N_6611,N_4297,N_4981);
or U6612 (N_6612,N_5618,N_4494);
or U6613 (N_6613,N_5770,N_4901);
and U6614 (N_6614,N_4626,N_4082);
and U6615 (N_6615,N_4661,N_5334);
nor U6616 (N_6616,N_5968,N_5068);
or U6617 (N_6617,N_4473,N_5232);
or U6618 (N_6618,N_5216,N_5152);
or U6619 (N_6619,N_4572,N_5979);
nor U6620 (N_6620,N_5904,N_4976);
nor U6621 (N_6621,N_4202,N_5395);
and U6622 (N_6622,N_4543,N_5003);
nand U6623 (N_6623,N_4679,N_4876);
nor U6624 (N_6624,N_5938,N_5996);
and U6625 (N_6625,N_5023,N_4766);
nand U6626 (N_6626,N_4940,N_5517);
or U6627 (N_6627,N_4488,N_4772);
and U6628 (N_6628,N_4018,N_4520);
nor U6629 (N_6629,N_5876,N_4405);
nor U6630 (N_6630,N_4872,N_5379);
and U6631 (N_6631,N_5425,N_4938);
or U6632 (N_6632,N_5699,N_5368);
or U6633 (N_6633,N_4760,N_5962);
nor U6634 (N_6634,N_5970,N_5291);
nor U6635 (N_6635,N_4913,N_5856);
or U6636 (N_6636,N_4347,N_4568);
nor U6637 (N_6637,N_5382,N_4798);
nand U6638 (N_6638,N_4226,N_5562);
nor U6639 (N_6639,N_4144,N_4925);
and U6640 (N_6640,N_4484,N_5525);
or U6641 (N_6641,N_5028,N_5077);
xor U6642 (N_6642,N_4048,N_4544);
xor U6643 (N_6643,N_5866,N_5224);
nand U6644 (N_6644,N_4275,N_4633);
nand U6645 (N_6645,N_5560,N_4418);
or U6646 (N_6646,N_4020,N_5652);
nor U6647 (N_6647,N_5958,N_4692);
nand U6648 (N_6648,N_5449,N_4132);
and U6649 (N_6649,N_5530,N_5355);
xnor U6650 (N_6650,N_5190,N_4990);
and U6651 (N_6651,N_5511,N_5702);
nand U6652 (N_6652,N_5930,N_5741);
and U6653 (N_6653,N_4489,N_4290);
nand U6654 (N_6654,N_5320,N_5301);
nor U6655 (N_6655,N_5150,N_4125);
xor U6656 (N_6656,N_4556,N_5784);
xnor U6657 (N_6657,N_5704,N_4711);
and U6658 (N_6658,N_4797,N_4054);
nor U6659 (N_6659,N_4024,N_5228);
xor U6660 (N_6660,N_4596,N_5182);
and U6661 (N_6661,N_5926,N_4744);
and U6662 (N_6662,N_4581,N_4006);
xnor U6663 (N_6663,N_5407,N_4214);
nor U6664 (N_6664,N_4722,N_4430);
nand U6665 (N_6665,N_4822,N_4288);
or U6666 (N_6666,N_5478,N_4369);
and U6667 (N_6667,N_5106,N_5550);
xnor U6668 (N_6668,N_4427,N_5380);
nand U6669 (N_6669,N_5985,N_4641);
nand U6670 (N_6670,N_5813,N_5546);
and U6671 (N_6671,N_4627,N_5740);
nand U6672 (N_6672,N_5128,N_4952);
nor U6673 (N_6673,N_4884,N_4378);
xor U6674 (N_6674,N_4287,N_5588);
nand U6675 (N_6675,N_4624,N_4754);
nor U6676 (N_6676,N_4808,N_5809);
nor U6677 (N_6677,N_5279,N_5609);
or U6678 (N_6678,N_4487,N_5549);
and U6679 (N_6679,N_4516,N_4113);
xnor U6680 (N_6680,N_4238,N_4714);
or U6681 (N_6681,N_4813,N_5386);
and U6682 (N_6682,N_5256,N_4243);
nand U6683 (N_6683,N_5118,N_4194);
or U6684 (N_6684,N_4438,N_4561);
nor U6685 (N_6685,N_5963,N_4792);
or U6686 (N_6686,N_5877,N_5120);
xor U6687 (N_6687,N_5552,N_4129);
nand U6688 (N_6688,N_4416,N_4083);
nand U6689 (N_6689,N_4725,N_4639);
or U6690 (N_6690,N_5378,N_5126);
nor U6691 (N_6691,N_5510,N_4593);
xnor U6692 (N_6692,N_5706,N_5544);
nor U6693 (N_6693,N_5698,N_5041);
and U6694 (N_6694,N_4914,N_5601);
xnor U6695 (N_6695,N_4126,N_4844);
and U6696 (N_6696,N_4156,N_5501);
and U6697 (N_6697,N_4234,N_4625);
and U6698 (N_6698,N_4086,N_5176);
and U6699 (N_6699,N_4609,N_4931);
nor U6700 (N_6700,N_5796,N_5980);
nor U6701 (N_6701,N_5403,N_4966);
xnor U6702 (N_6702,N_4149,N_5700);
and U6703 (N_6703,N_4192,N_4102);
nand U6704 (N_6704,N_5965,N_4005);
or U6705 (N_6705,N_4767,N_5042);
nor U6706 (N_6706,N_5536,N_4377);
and U6707 (N_6707,N_5878,N_4955);
nor U6708 (N_6708,N_4769,N_4173);
or U6709 (N_6709,N_4697,N_4286);
or U6710 (N_6710,N_5572,N_4583);
nor U6711 (N_6711,N_5657,N_5617);
or U6712 (N_6712,N_4070,N_4962);
nand U6713 (N_6713,N_4245,N_5697);
nor U6714 (N_6714,N_4828,N_4753);
xnor U6715 (N_6715,N_4143,N_5541);
nand U6716 (N_6716,N_5753,N_4289);
and U6717 (N_6717,N_5316,N_4199);
and U6718 (N_6718,N_4008,N_4363);
nor U6719 (N_6719,N_5000,N_5468);
nand U6720 (N_6720,N_5359,N_4576);
or U6721 (N_6721,N_4806,N_5936);
and U6722 (N_6722,N_5646,N_5004);
xnor U6723 (N_6723,N_5159,N_4327);
or U6724 (N_6724,N_4436,N_5308);
nor U6725 (N_6725,N_5912,N_4302);
and U6726 (N_6726,N_5537,N_4197);
nand U6727 (N_6727,N_4496,N_5391);
nand U6728 (N_6728,N_5062,N_5025);
or U6729 (N_6729,N_5328,N_4887);
nand U6730 (N_6730,N_4037,N_5461);
or U6731 (N_6731,N_4042,N_5843);
nor U6732 (N_6732,N_5854,N_5344);
or U6733 (N_6733,N_4227,N_4724);
xor U6734 (N_6734,N_4980,N_4944);
xor U6735 (N_6735,N_5688,N_5559);
nand U6736 (N_6736,N_4431,N_5762);
xor U6737 (N_6737,N_5971,N_4064);
nand U6738 (N_6738,N_5360,N_4653);
or U6739 (N_6739,N_5838,N_4345);
xnor U6740 (N_6740,N_4684,N_4112);
nor U6741 (N_6741,N_4472,N_4432);
nand U6742 (N_6742,N_5528,N_5453);
xnor U6743 (N_6743,N_4433,N_5345);
xnor U6744 (N_6744,N_4830,N_5332);
nor U6745 (N_6745,N_4412,N_5927);
xor U6746 (N_6746,N_4664,N_5317);
or U6747 (N_6747,N_4333,N_5055);
nand U6748 (N_6748,N_5750,N_4063);
xnor U6749 (N_6749,N_4415,N_4128);
nand U6750 (N_6750,N_5114,N_5716);
and U6751 (N_6751,N_5348,N_5719);
or U6752 (N_6752,N_4580,N_4135);
xor U6753 (N_6753,N_4718,N_4668);
nand U6754 (N_6754,N_5488,N_4617);
nor U6755 (N_6755,N_5502,N_5783);
nand U6756 (N_6756,N_4571,N_4535);
nor U6757 (N_6757,N_4175,N_4463);
or U6758 (N_6758,N_4600,N_5199);
nor U6759 (N_6759,N_5469,N_5558);
and U6760 (N_6760,N_4676,N_5995);
and U6761 (N_6761,N_4040,N_5986);
xor U6762 (N_6762,N_4059,N_5766);
or U6763 (N_6763,N_5811,N_4429);
nor U6764 (N_6764,N_5571,N_4647);
and U6765 (N_6765,N_5521,N_5569);
nor U6766 (N_6766,N_4816,N_4979);
nor U6767 (N_6767,N_5156,N_5178);
or U6768 (N_6768,N_5442,N_4291);
nor U6769 (N_6769,N_4538,N_5818);
nand U6770 (N_6770,N_4262,N_5347);
nor U6771 (N_6771,N_5458,N_5999);
and U6772 (N_6772,N_5708,N_5756);
nor U6773 (N_6773,N_4939,N_5690);
nor U6774 (N_6774,N_5874,N_5884);
nor U6775 (N_6775,N_4109,N_4902);
or U6776 (N_6776,N_5635,N_5539);
xnor U6777 (N_6777,N_4501,N_4309);
xor U6778 (N_6778,N_4166,N_5596);
xor U6779 (N_6779,N_4776,N_5663);
nor U6780 (N_6780,N_5235,N_5685);
nand U6781 (N_6781,N_5568,N_4342);
nor U6782 (N_6782,N_4203,N_5896);
or U6783 (N_6783,N_5935,N_5299);
and U6784 (N_6784,N_5802,N_5426);
or U6785 (N_6785,N_5435,N_4868);
or U6786 (N_6786,N_5991,N_5433);
and U6787 (N_6787,N_5031,N_4502);
xor U6788 (N_6788,N_4716,N_4049);
and U6789 (N_6789,N_5791,N_5388);
or U6790 (N_6790,N_5107,N_5053);
or U6791 (N_6791,N_5130,N_5261);
and U6792 (N_6792,N_5401,N_5123);
nor U6793 (N_6793,N_5828,N_4607);
and U6794 (N_6794,N_5889,N_4453);
nand U6795 (N_6795,N_4414,N_4176);
nand U6796 (N_6796,N_4120,N_5262);
nor U6797 (N_6797,N_4773,N_4662);
and U6798 (N_6798,N_5358,N_5440);
nand U6799 (N_6799,N_5675,N_5777);
nor U6800 (N_6800,N_5913,N_4546);
nand U6801 (N_6801,N_4230,N_4424);
and U6802 (N_6802,N_4677,N_4542);
or U6803 (N_6803,N_4968,N_4228);
nor U6804 (N_6804,N_5397,N_5200);
nor U6805 (N_6805,N_4545,N_4667);
or U6806 (N_6806,N_5709,N_4660);
xnor U6807 (N_6807,N_5201,N_5165);
or U6808 (N_6808,N_4991,N_4462);
nor U6809 (N_6809,N_4258,N_4923);
nand U6810 (N_6810,N_5054,N_4467);
and U6811 (N_6811,N_5888,N_5290);
or U6812 (N_6812,N_5082,N_5069);
and U6813 (N_6813,N_4740,N_5772);
nor U6814 (N_6814,N_4515,N_4741);
or U6815 (N_6815,N_5581,N_5891);
xnor U6816 (N_6816,N_5739,N_4736);
and U6817 (N_6817,N_5245,N_4179);
or U6818 (N_6818,N_4853,N_4651);
xnor U6819 (N_6819,N_5218,N_5574);
nor U6820 (N_6820,N_5019,N_5167);
or U6821 (N_6821,N_5269,N_5376);
xor U6822 (N_6822,N_5827,N_4852);
or U6823 (N_6823,N_5515,N_4448);
nor U6824 (N_6824,N_4255,N_4997);
nand U6825 (N_6825,N_4761,N_5535);
nor U6826 (N_6826,N_4186,N_4619);
nor U6827 (N_6827,N_4903,N_5234);
or U6828 (N_6828,N_4857,N_4597);
or U6829 (N_6829,N_5092,N_4338);
nor U6830 (N_6830,N_5280,N_4455);
and U6831 (N_6831,N_5364,N_5542);
xnor U6832 (N_6832,N_4930,N_5845);
xor U6833 (N_6833,N_4257,N_4376);
nor U6834 (N_6834,N_4413,N_5942);
and U6835 (N_6835,N_5322,N_5464);
nand U6836 (N_6836,N_5330,N_4727);
nand U6837 (N_6837,N_5436,N_4098);
nor U6838 (N_6838,N_4036,N_4936);
nor U6839 (N_6839,N_4693,N_5622);
nand U6840 (N_6840,N_5183,N_5015);
or U6841 (N_6841,N_4012,N_5751);
xor U6842 (N_6842,N_5861,N_5210);
xor U6843 (N_6843,N_4483,N_5208);
xor U6844 (N_6844,N_4329,N_4638);
or U6845 (N_6845,N_4408,N_4614);
nor U6846 (N_6846,N_4217,N_4656);
nand U6847 (N_6847,N_5808,N_4933);
nor U6848 (N_6848,N_5096,N_5413);
and U6849 (N_6849,N_4768,N_4871);
nand U6850 (N_6850,N_5032,N_5540);
nor U6851 (N_6851,N_4663,N_4687);
and U6852 (N_6852,N_4028,N_5035);
or U6853 (N_6853,N_5298,N_4612);
nor U6854 (N_6854,N_5570,N_5061);
or U6855 (N_6855,N_5180,N_5931);
and U6856 (N_6856,N_5922,N_4644);
nand U6857 (N_6857,N_5321,N_4848);
or U6858 (N_6858,N_5564,N_4870);
xor U6859 (N_6859,N_5624,N_5006);
nor U6860 (N_6860,N_4353,N_5265);
nand U6861 (N_6861,N_5073,N_5722);
xnor U6862 (N_6862,N_4136,N_5799);
or U6863 (N_6863,N_4140,N_5133);
nand U6864 (N_6864,N_5056,N_5823);
xor U6865 (N_6865,N_5198,N_5404);
and U6866 (N_6866,N_4486,N_4283);
or U6867 (N_6867,N_5049,N_4251);
or U6868 (N_6868,N_5365,N_4332);
or U6869 (N_6869,N_5253,N_5815);
or U6870 (N_6870,N_4052,N_5374);
nand U6871 (N_6871,N_4096,N_4421);
or U6872 (N_6872,N_4232,N_5375);
or U6873 (N_6873,N_5354,N_5335);
xnor U6874 (N_6874,N_4263,N_4480);
or U6875 (N_6875,N_5001,N_4720);
or U6876 (N_6876,N_5721,N_4972);
and U6877 (N_6877,N_4815,N_4368);
xor U6878 (N_6878,N_4133,N_4751);
and U6879 (N_6879,N_4269,N_4130);
and U6880 (N_6880,N_4013,N_4978);
or U6881 (N_6881,N_4518,N_4361);
or U6882 (N_6882,N_5039,N_4755);
or U6883 (N_6883,N_4242,N_5644);
and U6884 (N_6884,N_4105,N_5903);
xnor U6885 (N_6885,N_4295,N_5270);
and U6886 (N_6886,N_5718,N_5312);
nor U6887 (N_6887,N_5639,N_4558);
nor U6888 (N_6888,N_4869,N_5016);
nor U6889 (N_6889,N_4528,N_5272);
nor U6890 (N_6890,N_4392,N_4882);
nor U6891 (N_6891,N_4428,N_5221);
xnor U6892 (N_6892,N_4839,N_5138);
nor U6893 (N_6893,N_4069,N_5406);
xor U6894 (N_6894,N_4523,N_4492);
or U6895 (N_6895,N_5899,N_4967);
nor U6896 (N_6896,N_4009,N_4352);
nor U6897 (N_6897,N_4862,N_5385);
nor U6898 (N_6898,N_4536,N_5988);
nor U6899 (N_6899,N_5981,N_4456);
xnor U6900 (N_6900,N_4678,N_4482);
or U6901 (N_6901,N_4783,N_4382);
and U6902 (N_6902,N_5024,N_4444);
or U6903 (N_6903,N_5820,N_5771);
and U6904 (N_6904,N_5021,N_4640);
and U6905 (N_6905,N_5529,N_5186);
and U6906 (N_6906,N_4812,N_4785);
nand U6907 (N_6907,N_4799,N_4831);
nand U6908 (N_6908,N_4630,N_5122);
xnor U6909 (N_6909,N_5695,N_4547);
nor U6910 (N_6910,N_5116,N_5162);
or U6911 (N_6911,N_4749,N_4458);
nand U6912 (N_6912,N_4280,N_5941);
nor U6913 (N_6913,N_4169,N_5841);
nor U6914 (N_6914,N_5982,N_5390);
nand U6915 (N_6915,N_5658,N_5244);
nand U6916 (N_6916,N_4074,N_4575);
nand U6917 (N_6917,N_5014,N_4688);
nand U6918 (N_6918,N_5600,N_4675);
nand U6919 (N_6919,N_4829,N_4306);
nand U6920 (N_6920,N_5302,N_5243);
nor U6921 (N_6921,N_4511,N_5029);
nand U6922 (N_6922,N_4400,N_4434);
or U6923 (N_6923,N_5273,N_5890);
nand U6924 (N_6924,N_4341,N_4198);
nand U6925 (N_6925,N_4946,N_5940);
nor U6926 (N_6926,N_5398,N_4155);
and U6927 (N_6927,N_4702,N_5648);
xnor U6928 (N_6928,N_5768,N_5370);
nand U6929 (N_6929,N_5997,N_4584);
nor U6930 (N_6930,N_4019,N_5909);
nand U6931 (N_6931,N_4043,N_5669);
nand U6932 (N_6932,N_4324,N_4051);
nand U6933 (N_6933,N_5040,N_5337);
and U6934 (N_6934,N_5271,N_5870);
or U6935 (N_6935,N_4654,N_4497);
nor U6936 (N_6936,N_4748,N_5470);
xnor U6937 (N_6937,N_5246,N_5158);
xor U6938 (N_6938,N_4527,N_4604);
nor U6939 (N_6939,N_5816,N_4723);
xnor U6940 (N_6940,N_5636,N_5656);
xor U6941 (N_6941,N_4912,N_4780);
and U6942 (N_6942,N_4303,N_5251);
nor U6943 (N_6943,N_5242,N_4504);
and U6944 (N_6944,N_4689,N_5477);
or U6945 (N_6945,N_4891,N_4700);
nand U6946 (N_6946,N_5456,N_5620);
and U6947 (N_6947,N_5474,N_4335);
nand U6948 (N_6948,N_5746,N_4788);
or U6949 (N_6949,N_5074,N_5885);
nand U6950 (N_6950,N_4351,N_4770);
nor U6951 (N_6951,N_5276,N_4343);
xor U6952 (N_6952,N_5160,N_4949);
xnor U6953 (N_6953,N_4974,N_5124);
and U6954 (N_6954,N_4425,N_5196);
nor U6955 (N_6955,N_5844,N_5168);
nand U6956 (N_6956,N_4992,N_4252);
nand U6957 (N_6957,N_5475,N_5728);
nand U6958 (N_6958,N_4011,N_5769);
and U6959 (N_6959,N_5086,N_5580);
nor U6960 (N_6960,N_5621,N_4419);
and U6961 (N_6961,N_5939,N_4410);
or U6962 (N_6962,N_4894,N_5519);
xnor U6963 (N_6963,N_4278,N_5674);
or U6964 (N_6964,N_4594,N_4890);
nor U6965 (N_6965,N_4116,N_5713);
nand U6966 (N_6966,N_4945,N_4323);
nand U6967 (N_6967,N_5428,N_5022);
xnor U6968 (N_6968,N_5763,N_5631);
and U6969 (N_6969,N_4729,N_5538);
xor U6970 (N_6970,N_5258,N_5948);
or U6971 (N_6971,N_4032,N_4994);
xnor U6972 (N_6972,N_4279,N_4691);
and U6973 (N_6973,N_5471,N_4842);
and U6974 (N_6974,N_4163,N_4498);
xnor U6975 (N_6975,N_5071,N_5405);
nand U6976 (N_6976,N_4508,N_5135);
xnor U6977 (N_6977,N_4141,N_5754);
and U6978 (N_6978,N_4185,N_4733);
or U6979 (N_6979,N_5371,N_5483);
nand U6980 (N_6980,N_5283,N_5893);
nand U6981 (N_6981,N_5482,N_4731);
nor U6982 (N_6982,N_5683,N_5686);
nand U6983 (N_6983,N_4618,N_5033);
or U6984 (N_6984,N_4440,N_4110);
nand U6985 (N_6985,N_4696,N_5566);
xor U6986 (N_6986,N_5420,N_4224);
nor U6987 (N_6987,N_4266,N_4313);
and U6988 (N_6988,N_5782,N_5825);
xor U6989 (N_6989,N_5342,N_5628);
nor U6990 (N_6990,N_5691,N_4794);
or U6991 (N_6991,N_5696,N_4750);
nand U6992 (N_6992,N_5587,N_5774);
nor U6993 (N_6993,N_4924,N_4984);
nor U6994 (N_6994,N_4210,N_5707);
xor U6995 (N_6995,N_5806,N_4998);
and U6996 (N_6996,N_4682,N_4393);
xnor U6997 (N_6997,N_5441,N_5416);
and U6998 (N_6998,N_4595,N_5236);
and U6999 (N_6999,N_4476,N_4437);
nor U7000 (N_7000,N_4995,N_5446);
and U7001 (N_7001,N_5608,N_4580);
xor U7002 (N_7002,N_5055,N_4773);
or U7003 (N_7003,N_4010,N_5732);
xnor U7004 (N_7004,N_4568,N_4631);
nand U7005 (N_7005,N_4580,N_4076);
or U7006 (N_7006,N_4256,N_5793);
nand U7007 (N_7007,N_5290,N_5941);
and U7008 (N_7008,N_5731,N_5849);
and U7009 (N_7009,N_5917,N_5201);
nand U7010 (N_7010,N_5848,N_5292);
xor U7011 (N_7011,N_5819,N_4574);
nand U7012 (N_7012,N_4458,N_4440);
and U7013 (N_7013,N_4329,N_5154);
or U7014 (N_7014,N_4077,N_5544);
or U7015 (N_7015,N_5243,N_4638);
or U7016 (N_7016,N_5920,N_4547);
or U7017 (N_7017,N_5765,N_4918);
nand U7018 (N_7018,N_4273,N_4114);
nor U7019 (N_7019,N_5391,N_4429);
or U7020 (N_7020,N_5650,N_5164);
nor U7021 (N_7021,N_5511,N_4329);
nor U7022 (N_7022,N_4819,N_4384);
or U7023 (N_7023,N_5661,N_5432);
or U7024 (N_7024,N_5823,N_4275);
or U7025 (N_7025,N_4167,N_5176);
or U7026 (N_7026,N_4594,N_4537);
or U7027 (N_7027,N_4876,N_5167);
nand U7028 (N_7028,N_4080,N_5356);
nor U7029 (N_7029,N_5429,N_4521);
and U7030 (N_7030,N_4811,N_5232);
or U7031 (N_7031,N_5705,N_5086);
and U7032 (N_7032,N_5355,N_4126);
or U7033 (N_7033,N_4798,N_5158);
nand U7034 (N_7034,N_5212,N_5507);
xor U7035 (N_7035,N_4004,N_5170);
nor U7036 (N_7036,N_5809,N_5273);
nand U7037 (N_7037,N_5166,N_4279);
and U7038 (N_7038,N_4394,N_5946);
or U7039 (N_7039,N_4349,N_5693);
and U7040 (N_7040,N_5975,N_4777);
nand U7041 (N_7041,N_4821,N_5282);
nor U7042 (N_7042,N_5401,N_5264);
nor U7043 (N_7043,N_4576,N_4175);
xnor U7044 (N_7044,N_4909,N_4104);
xor U7045 (N_7045,N_4215,N_4311);
and U7046 (N_7046,N_4749,N_5370);
or U7047 (N_7047,N_5769,N_5938);
xor U7048 (N_7048,N_5234,N_5090);
xnor U7049 (N_7049,N_4535,N_5639);
and U7050 (N_7050,N_5181,N_5233);
or U7051 (N_7051,N_4593,N_4671);
or U7052 (N_7052,N_4860,N_4945);
nand U7053 (N_7053,N_5037,N_5758);
nor U7054 (N_7054,N_5433,N_5163);
xnor U7055 (N_7055,N_4871,N_4778);
nand U7056 (N_7056,N_4958,N_5091);
nand U7057 (N_7057,N_5370,N_5719);
nor U7058 (N_7058,N_5205,N_4139);
xor U7059 (N_7059,N_5644,N_4980);
or U7060 (N_7060,N_5871,N_5878);
nor U7061 (N_7061,N_4888,N_5273);
nor U7062 (N_7062,N_4188,N_5509);
and U7063 (N_7063,N_4444,N_4753);
nand U7064 (N_7064,N_4788,N_5828);
nand U7065 (N_7065,N_4961,N_4188);
and U7066 (N_7066,N_4295,N_4163);
xor U7067 (N_7067,N_4097,N_4908);
and U7068 (N_7068,N_4261,N_5431);
and U7069 (N_7069,N_5914,N_4474);
or U7070 (N_7070,N_4780,N_5035);
and U7071 (N_7071,N_5843,N_5479);
xnor U7072 (N_7072,N_4995,N_4688);
and U7073 (N_7073,N_4847,N_5772);
nor U7074 (N_7074,N_4450,N_4912);
and U7075 (N_7075,N_4263,N_5932);
nor U7076 (N_7076,N_5541,N_4754);
nand U7077 (N_7077,N_4987,N_5764);
nor U7078 (N_7078,N_4736,N_4342);
nor U7079 (N_7079,N_4357,N_5201);
nand U7080 (N_7080,N_5702,N_4683);
or U7081 (N_7081,N_4538,N_4126);
xnor U7082 (N_7082,N_4213,N_4401);
nor U7083 (N_7083,N_5325,N_5439);
nand U7084 (N_7084,N_5275,N_4132);
nor U7085 (N_7085,N_4226,N_4323);
nor U7086 (N_7086,N_4806,N_4284);
or U7087 (N_7087,N_4242,N_5593);
nand U7088 (N_7088,N_4868,N_5136);
nor U7089 (N_7089,N_4068,N_5167);
nor U7090 (N_7090,N_5435,N_4264);
and U7091 (N_7091,N_4805,N_4734);
nor U7092 (N_7092,N_5197,N_5497);
nand U7093 (N_7093,N_4684,N_4213);
and U7094 (N_7094,N_5885,N_5668);
and U7095 (N_7095,N_5204,N_4244);
and U7096 (N_7096,N_4789,N_4583);
nor U7097 (N_7097,N_5161,N_5134);
nand U7098 (N_7098,N_4842,N_5206);
or U7099 (N_7099,N_4543,N_5835);
or U7100 (N_7100,N_4370,N_4746);
nor U7101 (N_7101,N_5404,N_5759);
nand U7102 (N_7102,N_5906,N_5090);
xor U7103 (N_7103,N_4352,N_4526);
or U7104 (N_7104,N_4692,N_4209);
xnor U7105 (N_7105,N_5296,N_5604);
nor U7106 (N_7106,N_4679,N_4251);
nor U7107 (N_7107,N_4019,N_5512);
nor U7108 (N_7108,N_5913,N_5426);
and U7109 (N_7109,N_4810,N_4831);
or U7110 (N_7110,N_5901,N_4596);
and U7111 (N_7111,N_5292,N_4990);
or U7112 (N_7112,N_5804,N_4650);
nand U7113 (N_7113,N_4208,N_5576);
or U7114 (N_7114,N_5165,N_5595);
or U7115 (N_7115,N_5108,N_4094);
nor U7116 (N_7116,N_5151,N_5299);
nand U7117 (N_7117,N_4901,N_4873);
nand U7118 (N_7118,N_5073,N_4250);
and U7119 (N_7119,N_4794,N_4898);
or U7120 (N_7120,N_5444,N_5491);
nand U7121 (N_7121,N_4943,N_5541);
xnor U7122 (N_7122,N_4638,N_5689);
nor U7123 (N_7123,N_4720,N_5820);
or U7124 (N_7124,N_4713,N_5150);
nand U7125 (N_7125,N_5823,N_4122);
nand U7126 (N_7126,N_5665,N_5718);
xor U7127 (N_7127,N_4982,N_5685);
and U7128 (N_7128,N_4736,N_5401);
nand U7129 (N_7129,N_4154,N_5051);
xnor U7130 (N_7130,N_5235,N_4352);
or U7131 (N_7131,N_4009,N_4533);
and U7132 (N_7132,N_5934,N_5781);
and U7133 (N_7133,N_5356,N_5448);
and U7134 (N_7134,N_4846,N_5866);
nor U7135 (N_7135,N_5838,N_5386);
and U7136 (N_7136,N_5526,N_5241);
or U7137 (N_7137,N_5085,N_4202);
or U7138 (N_7138,N_4287,N_5916);
or U7139 (N_7139,N_4983,N_5740);
xor U7140 (N_7140,N_5785,N_4555);
nand U7141 (N_7141,N_4144,N_4598);
nand U7142 (N_7142,N_5035,N_5939);
or U7143 (N_7143,N_4620,N_4181);
and U7144 (N_7144,N_4025,N_5250);
nand U7145 (N_7145,N_4172,N_4638);
or U7146 (N_7146,N_5425,N_5994);
and U7147 (N_7147,N_5623,N_4099);
nand U7148 (N_7148,N_5184,N_5014);
or U7149 (N_7149,N_5249,N_5204);
or U7150 (N_7150,N_4742,N_4048);
nor U7151 (N_7151,N_4591,N_5829);
nand U7152 (N_7152,N_4582,N_5290);
xor U7153 (N_7153,N_4754,N_4475);
nand U7154 (N_7154,N_4574,N_4389);
or U7155 (N_7155,N_4563,N_4305);
nor U7156 (N_7156,N_5746,N_4028);
xnor U7157 (N_7157,N_4147,N_5359);
xor U7158 (N_7158,N_5363,N_5405);
nor U7159 (N_7159,N_5239,N_4061);
nand U7160 (N_7160,N_4702,N_5435);
or U7161 (N_7161,N_4699,N_4616);
xnor U7162 (N_7162,N_5955,N_5837);
nand U7163 (N_7163,N_4866,N_5613);
nor U7164 (N_7164,N_5783,N_5950);
nand U7165 (N_7165,N_5173,N_5482);
nand U7166 (N_7166,N_4422,N_5533);
xnor U7167 (N_7167,N_4295,N_5247);
nand U7168 (N_7168,N_4073,N_4172);
or U7169 (N_7169,N_5730,N_5796);
nor U7170 (N_7170,N_4004,N_5924);
nor U7171 (N_7171,N_4898,N_4583);
and U7172 (N_7172,N_4188,N_4998);
nand U7173 (N_7173,N_4881,N_5697);
nor U7174 (N_7174,N_5586,N_5507);
nand U7175 (N_7175,N_4315,N_4700);
nor U7176 (N_7176,N_5005,N_5686);
and U7177 (N_7177,N_5610,N_4307);
or U7178 (N_7178,N_5524,N_5074);
xnor U7179 (N_7179,N_4784,N_4054);
nand U7180 (N_7180,N_4831,N_5990);
nand U7181 (N_7181,N_4177,N_5956);
nor U7182 (N_7182,N_5850,N_4368);
nand U7183 (N_7183,N_5551,N_4883);
xnor U7184 (N_7184,N_4282,N_5558);
and U7185 (N_7185,N_4404,N_4568);
or U7186 (N_7186,N_4921,N_4141);
or U7187 (N_7187,N_4287,N_5847);
or U7188 (N_7188,N_5181,N_4821);
and U7189 (N_7189,N_4950,N_4198);
nor U7190 (N_7190,N_4122,N_5606);
xor U7191 (N_7191,N_5143,N_4751);
or U7192 (N_7192,N_4182,N_4052);
or U7193 (N_7193,N_4632,N_5700);
nor U7194 (N_7194,N_5071,N_4637);
nand U7195 (N_7195,N_5752,N_4020);
and U7196 (N_7196,N_4172,N_5346);
or U7197 (N_7197,N_4470,N_5202);
and U7198 (N_7198,N_5818,N_4060);
and U7199 (N_7199,N_5464,N_4661);
or U7200 (N_7200,N_4693,N_5462);
and U7201 (N_7201,N_5555,N_4862);
xor U7202 (N_7202,N_4055,N_5136);
nand U7203 (N_7203,N_5824,N_4778);
and U7204 (N_7204,N_4179,N_4862);
nand U7205 (N_7205,N_5167,N_5072);
and U7206 (N_7206,N_4535,N_4240);
and U7207 (N_7207,N_5658,N_5806);
and U7208 (N_7208,N_4217,N_5513);
xor U7209 (N_7209,N_4443,N_5513);
and U7210 (N_7210,N_5586,N_4655);
and U7211 (N_7211,N_4112,N_4110);
xor U7212 (N_7212,N_5461,N_4147);
or U7213 (N_7213,N_5518,N_4494);
nor U7214 (N_7214,N_5894,N_5880);
nand U7215 (N_7215,N_5286,N_4734);
nor U7216 (N_7216,N_5858,N_5581);
nand U7217 (N_7217,N_4628,N_4827);
or U7218 (N_7218,N_4218,N_5260);
and U7219 (N_7219,N_4904,N_5044);
and U7220 (N_7220,N_4845,N_4203);
nand U7221 (N_7221,N_4991,N_4941);
or U7222 (N_7222,N_4128,N_4095);
or U7223 (N_7223,N_4791,N_5023);
xor U7224 (N_7224,N_5836,N_5817);
xnor U7225 (N_7225,N_4780,N_5706);
and U7226 (N_7226,N_4637,N_4478);
xnor U7227 (N_7227,N_5112,N_5717);
and U7228 (N_7228,N_5788,N_5780);
or U7229 (N_7229,N_4593,N_4182);
nand U7230 (N_7230,N_5592,N_5977);
nor U7231 (N_7231,N_4892,N_4592);
nand U7232 (N_7232,N_5625,N_4030);
xnor U7233 (N_7233,N_4398,N_4308);
xnor U7234 (N_7234,N_5921,N_5338);
and U7235 (N_7235,N_5815,N_4921);
and U7236 (N_7236,N_4246,N_4510);
xnor U7237 (N_7237,N_4951,N_4396);
nand U7238 (N_7238,N_5300,N_5703);
or U7239 (N_7239,N_4513,N_5541);
xor U7240 (N_7240,N_5500,N_5012);
xnor U7241 (N_7241,N_5529,N_4319);
and U7242 (N_7242,N_4644,N_4438);
and U7243 (N_7243,N_4858,N_4232);
xnor U7244 (N_7244,N_5651,N_5134);
nand U7245 (N_7245,N_4915,N_5774);
nor U7246 (N_7246,N_5052,N_5695);
and U7247 (N_7247,N_4879,N_5489);
nor U7248 (N_7248,N_5109,N_4809);
nor U7249 (N_7249,N_4337,N_5663);
and U7250 (N_7250,N_4512,N_5936);
or U7251 (N_7251,N_4455,N_5656);
xnor U7252 (N_7252,N_5226,N_4189);
or U7253 (N_7253,N_5057,N_5914);
nor U7254 (N_7254,N_5826,N_5959);
xnor U7255 (N_7255,N_4170,N_4661);
or U7256 (N_7256,N_5441,N_4469);
or U7257 (N_7257,N_4654,N_4713);
or U7258 (N_7258,N_5849,N_5743);
xnor U7259 (N_7259,N_4765,N_4826);
nand U7260 (N_7260,N_5543,N_5885);
nand U7261 (N_7261,N_4440,N_5653);
nand U7262 (N_7262,N_4334,N_4200);
and U7263 (N_7263,N_5925,N_5428);
nor U7264 (N_7264,N_4767,N_4882);
xnor U7265 (N_7265,N_4730,N_5637);
xor U7266 (N_7266,N_5304,N_4019);
or U7267 (N_7267,N_5176,N_5646);
nor U7268 (N_7268,N_5412,N_5941);
xnor U7269 (N_7269,N_4004,N_4587);
or U7270 (N_7270,N_5181,N_4548);
xnor U7271 (N_7271,N_4719,N_4611);
xor U7272 (N_7272,N_4771,N_4512);
nor U7273 (N_7273,N_5522,N_5074);
or U7274 (N_7274,N_5202,N_4560);
and U7275 (N_7275,N_5921,N_5411);
nand U7276 (N_7276,N_4956,N_5953);
or U7277 (N_7277,N_5826,N_4528);
xor U7278 (N_7278,N_4665,N_4975);
xor U7279 (N_7279,N_4889,N_5175);
xnor U7280 (N_7280,N_5385,N_5618);
xor U7281 (N_7281,N_4950,N_5500);
nor U7282 (N_7282,N_5238,N_5788);
nor U7283 (N_7283,N_4611,N_5784);
xnor U7284 (N_7284,N_4774,N_5234);
and U7285 (N_7285,N_5643,N_4060);
and U7286 (N_7286,N_4164,N_5544);
or U7287 (N_7287,N_4469,N_4410);
xnor U7288 (N_7288,N_5650,N_5563);
nand U7289 (N_7289,N_4984,N_4898);
nand U7290 (N_7290,N_4816,N_4093);
nand U7291 (N_7291,N_5695,N_4279);
or U7292 (N_7292,N_4089,N_5641);
xor U7293 (N_7293,N_4714,N_4346);
and U7294 (N_7294,N_5771,N_5089);
xnor U7295 (N_7295,N_4058,N_5063);
nand U7296 (N_7296,N_4121,N_5415);
or U7297 (N_7297,N_4517,N_5671);
nand U7298 (N_7298,N_5324,N_5172);
and U7299 (N_7299,N_5908,N_5190);
nor U7300 (N_7300,N_5322,N_5227);
nand U7301 (N_7301,N_5495,N_4590);
or U7302 (N_7302,N_4210,N_4181);
and U7303 (N_7303,N_5420,N_5604);
nand U7304 (N_7304,N_4198,N_4344);
xor U7305 (N_7305,N_5650,N_4068);
xnor U7306 (N_7306,N_5796,N_4337);
nor U7307 (N_7307,N_5723,N_4833);
or U7308 (N_7308,N_4551,N_4073);
nand U7309 (N_7309,N_4521,N_5172);
nand U7310 (N_7310,N_4097,N_5365);
nand U7311 (N_7311,N_5405,N_4988);
and U7312 (N_7312,N_5411,N_5242);
and U7313 (N_7313,N_5814,N_5490);
nand U7314 (N_7314,N_5095,N_4610);
or U7315 (N_7315,N_4750,N_5857);
and U7316 (N_7316,N_4817,N_4033);
xnor U7317 (N_7317,N_5507,N_5268);
nand U7318 (N_7318,N_4300,N_4215);
nor U7319 (N_7319,N_5318,N_5585);
nor U7320 (N_7320,N_5428,N_5167);
and U7321 (N_7321,N_5297,N_5367);
nand U7322 (N_7322,N_5845,N_4482);
xnor U7323 (N_7323,N_5622,N_5616);
or U7324 (N_7324,N_4803,N_5540);
or U7325 (N_7325,N_4982,N_5477);
and U7326 (N_7326,N_5097,N_5864);
nand U7327 (N_7327,N_4076,N_5153);
and U7328 (N_7328,N_4664,N_5199);
and U7329 (N_7329,N_5042,N_4467);
or U7330 (N_7330,N_5771,N_4430);
or U7331 (N_7331,N_5354,N_5676);
nand U7332 (N_7332,N_5431,N_4245);
nor U7333 (N_7333,N_4658,N_5228);
nand U7334 (N_7334,N_5710,N_4380);
xor U7335 (N_7335,N_4725,N_4942);
and U7336 (N_7336,N_5931,N_5162);
nor U7337 (N_7337,N_5629,N_5164);
xor U7338 (N_7338,N_5033,N_5452);
xnor U7339 (N_7339,N_4941,N_5820);
nand U7340 (N_7340,N_5243,N_4389);
and U7341 (N_7341,N_5505,N_4971);
and U7342 (N_7342,N_4992,N_5877);
and U7343 (N_7343,N_5646,N_5787);
nand U7344 (N_7344,N_5216,N_5266);
nand U7345 (N_7345,N_5387,N_5621);
and U7346 (N_7346,N_5870,N_4262);
xor U7347 (N_7347,N_5582,N_5295);
nor U7348 (N_7348,N_5661,N_5015);
or U7349 (N_7349,N_5333,N_5330);
or U7350 (N_7350,N_4355,N_4899);
nand U7351 (N_7351,N_5597,N_5494);
nor U7352 (N_7352,N_5466,N_5836);
nor U7353 (N_7353,N_5539,N_4558);
or U7354 (N_7354,N_5067,N_5968);
or U7355 (N_7355,N_4245,N_4739);
nand U7356 (N_7356,N_4421,N_5094);
or U7357 (N_7357,N_4600,N_5941);
or U7358 (N_7358,N_5883,N_5777);
or U7359 (N_7359,N_5966,N_5135);
nor U7360 (N_7360,N_5748,N_4377);
and U7361 (N_7361,N_4897,N_4263);
and U7362 (N_7362,N_4715,N_5252);
or U7363 (N_7363,N_4803,N_5827);
xor U7364 (N_7364,N_4091,N_5614);
or U7365 (N_7365,N_5197,N_4421);
nand U7366 (N_7366,N_4502,N_5173);
xor U7367 (N_7367,N_5971,N_5894);
or U7368 (N_7368,N_4572,N_4942);
xor U7369 (N_7369,N_5144,N_4170);
or U7370 (N_7370,N_4783,N_5644);
nor U7371 (N_7371,N_5977,N_5784);
or U7372 (N_7372,N_4164,N_4331);
xor U7373 (N_7373,N_4279,N_5925);
and U7374 (N_7374,N_4607,N_4248);
or U7375 (N_7375,N_4907,N_4464);
nand U7376 (N_7376,N_4197,N_4111);
or U7377 (N_7377,N_4216,N_5238);
or U7378 (N_7378,N_4105,N_4701);
xor U7379 (N_7379,N_5636,N_4717);
and U7380 (N_7380,N_5769,N_5883);
nand U7381 (N_7381,N_4892,N_5681);
nor U7382 (N_7382,N_4693,N_5543);
nor U7383 (N_7383,N_4180,N_4738);
nand U7384 (N_7384,N_5571,N_5869);
nor U7385 (N_7385,N_4082,N_5119);
and U7386 (N_7386,N_4105,N_4704);
or U7387 (N_7387,N_4696,N_4605);
xnor U7388 (N_7388,N_4423,N_4583);
xor U7389 (N_7389,N_5747,N_5760);
and U7390 (N_7390,N_4189,N_4407);
or U7391 (N_7391,N_5422,N_5672);
xor U7392 (N_7392,N_4509,N_5278);
nor U7393 (N_7393,N_5298,N_5740);
and U7394 (N_7394,N_5440,N_4879);
or U7395 (N_7395,N_5109,N_5747);
xnor U7396 (N_7396,N_4319,N_4937);
nor U7397 (N_7397,N_5758,N_5481);
xor U7398 (N_7398,N_5084,N_4703);
and U7399 (N_7399,N_4642,N_5916);
and U7400 (N_7400,N_4402,N_5753);
nor U7401 (N_7401,N_5827,N_5673);
nand U7402 (N_7402,N_4256,N_4735);
nand U7403 (N_7403,N_4714,N_4299);
and U7404 (N_7404,N_5786,N_5911);
and U7405 (N_7405,N_5762,N_4513);
or U7406 (N_7406,N_4758,N_5323);
xnor U7407 (N_7407,N_5102,N_5008);
nor U7408 (N_7408,N_5022,N_5636);
nand U7409 (N_7409,N_4282,N_4860);
xnor U7410 (N_7410,N_4175,N_5665);
nor U7411 (N_7411,N_4097,N_4562);
nand U7412 (N_7412,N_5038,N_5943);
nand U7413 (N_7413,N_5162,N_5104);
nor U7414 (N_7414,N_4223,N_5538);
nand U7415 (N_7415,N_5131,N_5668);
nand U7416 (N_7416,N_5203,N_4291);
nor U7417 (N_7417,N_5009,N_4710);
or U7418 (N_7418,N_4050,N_4236);
xnor U7419 (N_7419,N_4520,N_4501);
nor U7420 (N_7420,N_4427,N_4248);
xnor U7421 (N_7421,N_5147,N_5457);
and U7422 (N_7422,N_4045,N_4531);
xor U7423 (N_7423,N_5500,N_4485);
nor U7424 (N_7424,N_5761,N_4521);
xnor U7425 (N_7425,N_5172,N_4622);
or U7426 (N_7426,N_5211,N_5895);
xnor U7427 (N_7427,N_4729,N_5523);
and U7428 (N_7428,N_5318,N_5415);
and U7429 (N_7429,N_5791,N_5060);
nor U7430 (N_7430,N_5241,N_5332);
and U7431 (N_7431,N_5964,N_4797);
nor U7432 (N_7432,N_5088,N_5166);
xor U7433 (N_7433,N_5700,N_4686);
or U7434 (N_7434,N_5327,N_4809);
nor U7435 (N_7435,N_5707,N_4091);
and U7436 (N_7436,N_4111,N_5998);
and U7437 (N_7437,N_4118,N_5362);
nor U7438 (N_7438,N_5767,N_5599);
xnor U7439 (N_7439,N_5714,N_5268);
nor U7440 (N_7440,N_4797,N_5251);
nor U7441 (N_7441,N_5967,N_5790);
or U7442 (N_7442,N_4855,N_4771);
or U7443 (N_7443,N_4182,N_4424);
xnor U7444 (N_7444,N_4309,N_5097);
nor U7445 (N_7445,N_4014,N_4681);
nand U7446 (N_7446,N_5002,N_4208);
or U7447 (N_7447,N_5057,N_4908);
nor U7448 (N_7448,N_4853,N_5485);
xor U7449 (N_7449,N_4416,N_4887);
nor U7450 (N_7450,N_4455,N_4197);
nor U7451 (N_7451,N_4359,N_5710);
nor U7452 (N_7452,N_5335,N_4711);
nand U7453 (N_7453,N_4249,N_5747);
xor U7454 (N_7454,N_5002,N_5397);
and U7455 (N_7455,N_4715,N_4297);
nand U7456 (N_7456,N_5590,N_4811);
and U7457 (N_7457,N_4783,N_5902);
nor U7458 (N_7458,N_5161,N_5657);
and U7459 (N_7459,N_4338,N_5562);
nor U7460 (N_7460,N_5951,N_4518);
nand U7461 (N_7461,N_4971,N_5990);
xor U7462 (N_7462,N_5341,N_4832);
or U7463 (N_7463,N_4132,N_4817);
nor U7464 (N_7464,N_5982,N_5850);
nand U7465 (N_7465,N_4498,N_5443);
nor U7466 (N_7466,N_4701,N_4983);
nor U7467 (N_7467,N_4159,N_4219);
xor U7468 (N_7468,N_4073,N_5302);
xnor U7469 (N_7469,N_4852,N_5447);
xnor U7470 (N_7470,N_5775,N_4461);
and U7471 (N_7471,N_4230,N_4725);
and U7472 (N_7472,N_5442,N_4800);
or U7473 (N_7473,N_5318,N_4195);
xor U7474 (N_7474,N_4619,N_5072);
nor U7475 (N_7475,N_5310,N_4747);
nand U7476 (N_7476,N_5912,N_5183);
or U7477 (N_7477,N_5724,N_4380);
nand U7478 (N_7478,N_5063,N_5726);
nor U7479 (N_7479,N_4235,N_4524);
nand U7480 (N_7480,N_5602,N_5843);
and U7481 (N_7481,N_5353,N_4871);
or U7482 (N_7482,N_5277,N_4078);
nand U7483 (N_7483,N_4852,N_5746);
nor U7484 (N_7484,N_4286,N_5869);
nor U7485 (N_7485,N_4945,N_5913);
nor U7486 (N_7486,N_4858,N_5526);
and U7487 (N_7487,N_4745,N_4697);
xnor U7488 (N_7488,N_4652,N_4743);
or U7489 (N_7489,N_4761,N_4160);
nor U7490 (N_7490,N_4081,N_4975);
nand U7491 (N_7491,N_5208,N_5340);
xor U7492 (N_7492,N_4905,N_5465);
nand U7493 (N_7493,N_5221,N_5145);
xor U7494 (N_7494,N_5153,N_4801);
or U7495 (N_7495,N_5690,N_5304);
nor U7496 (N_7496,N_4555,N_4885);
and U7497 (N_7497,N_4026,N_4439);
or U7498 (N_7498,N_4716,N_5905);
and U7499 (N_7499,N_5419,N_4938);
or U7500 (N_7500,N_4305,N_4030);
nor U7501 (N_7501,N_4795,N_5683);
and U7502 (N_7502,N_5954,N_4474);
xor U7503 (N_7503,N_4408,N_5525);
xnor U7504 (N_7504,N_5612,N_4739);
or U7505 (N_7505,N_5374,N_4067);
nand U7506 (N_7506,N_4359,N_4852);
nor U7507 (N_7507,N_4599,N_4180);
and U7508 (N_7508,N_4857,N_5611);
and U7509 (N_7509,N_4486,N_5332);
nor U7510 (N_7510,N_5632,N_4987);
nor U7511 (N_7511,N_5545,N_5553);
and U7512 (N_7512,N_4492,N_5912);
and U7513 (N_7513,N_4406,N_5024);
nor U7514 (N_7514,N_5031,N_5846);
nor U7515 (N_7515,N_5293,N_5701);
nand U7516 (N_7516,N_5625,N_4693);
nor U7517 (N_7517,N_4077,N_5414);
or U7518 (N_7518,N_5206,N_5948);
or U7519 (N_7519,N_5632,N_5504);
nand U7520 (N_7520,N_4947,N_5735);
or U7521 (N_7521,N_4528,N_4969);
and U7522 (N_7522,N_4064,N_5128);
nor U7523 (N_7523,N_4083,N_4371);
and U7524 (N_7524,N_4858,N_5229);
or U7525 (N_7525,N_4543,N_5909);
nand U7526 (N_7526,N_4736,N_4151);
nor U7527 (N_7527,N_4997,N_4387);
and U7528 (N_7528,N_5314,N_5012);
or U7529 (N_7529,N_5102,N_4197);
and U7530 (N_7530,N_5858,N_5619);
and U7531 (N_7531,N_4808,N_5174);
or U7532 (N_7532,N_5272,N_4978);
or U7533 (N_7533,N_5553,N_5708);
and U7534 (N_7534,N_5859,N_4508);
and U7535 (N_7535,N_4539,N_5944);
and U7536 (N_7536,N_5590,N_5768);
nand U7537 (N_7537,N_5250,N_5953);
nand U7538 (N_7538,N_4106,N_5743);
nor U7539 (N_7539,N_5062,N_5716);
and U7540 (N_7540,N_5540,N_5502);
nor U7541 (N_7541,N_4723,N_4455);
xor U7542 (N_7542,N_5789,N_5157);
xnor U7543 (N_7543,N_5690,N_4361);
or U7544 (N_7544,N_5998,N_4038);
or U7545 (N_7545,N_4345,N_4429);
xnor U7546 (N_7546,N_5458,N_4485);
xor U7547 (N_7547,N_5311,N_5054);
and U7548 (N_7548,N_5842,N_4197);
and U7549 (N_7549,N_4689,N_4179);
and U7550 (N_7550,N_5998,N_4091);
nand U7551 (N_7551,N_4170,N_5362);
nand U7552 (N_7552,N_4075,N_4531);
xnor U7553 (N_7553,N_5195,N_5876);
and U7554 (N_7554,N_4870,N_4309);
or U7555 (N_7555,N_5082,N_5565);
nor U7556 (N_7556,N_4302,N_5700);
and U7557 (N_7557,N_5930,N_4325);
and U7558 (N_7558,N_5431,N_4013);
xor U7559 (N_7559,N_4597,N_5631);
and U7560 (N_7560,N_4697,N_5803);
xnor U7561 (N_7561,N_5282,N_5881);
and U7562 (N_7562,N_5645,N_5774);
and U7563 (N_7563,N_4995,N_4098);
and U7564 (N_7564,N_4734,N_4373);
nor U7565 (N_7565,N_5503,N_5981);
xor U7566 (N_7566,N_5881,N_4007);
and U7567 (N_7567,N_5638,N_5345);
nand U7568 (N_7568,N_4457,N_5668);
or U7569 (N_7569,N_4162,N_5754);
xor U7570 (N_7570,N_4271,N_4310);
xnor U7571 (N_7571,N_4743,N_5272);
or U7572 (N_7572,N_4723,N_4315);
nand U7573 (N_7573,N_5191,N_4517);
nand U7574 (N_7574,N_5558,N_5804);
xnor U7575 (N_7575,N_4956,N_5345);
and U7576 (N_7576,N_5673,N_5102);
and U7577 (N_7577,N_5772,N_5930);
or U7578 (N_7578,N_5690,N_4132);
nor U7579 (N_7579,N_4811,N_5930);
nor U7580 (N_7580,N_5549,N_4290);
nand U7581 (N_7581,N_5775,N_4742);
and U7582 (N_7582,N_4886,N_5324);
xnor U7583 (N_7583,N_5932,N_4099);
or U7584 (N_7584,N_4965,N_5449);
or U7585 (N_7585,N_4595,N_5184);
xnor U7586 (N_7586,N_5886,N_4477);
xnor U7587 (N_7587,N_4855,N_4554);
nor U7588 (N_7588,N_5172,N_4901);
xnor U7589 (N_7589,N_5598,N_5400);
or U7590 (N_7590,N_5337,N_4179);
xnor U7591 (N_7591,N_5867,N_5240);
and U7592 (N_7592,N_4218,N_5728);
and U7593 (N_7593,N_4780,N_5531);
nand U7594 (N_7594,N_4597,N_5850);
nor U7595 (N_7595,N_5643,N_5308);
nor U7596 (N_7596,N_5687,N_4693);
and U7597 (N_7597,N_5924,N_4182);
nor U7598 (N_7598,N_4833,N_5328);
or U7599 (N_7599,N_4751,N_4921);
nor U7600 (N_7600,N_4297,N_4161);
nor U7601 (N_7601,N_4546,N_4843);
and U7602 (N_7602,N_4272,N_4881);
xnor U7603 (N_7603,N_4755,N_5255);
nand U7604 (N_7604,N_4761,N_5631);
nand U7605 (N_7605,N_5720,N_5190);
or U7606 (N_7606,N_4838,N_5840);
nor U7607 (N_7607,N_5174,N_5281);
xor U7608 (N_7608,N_4122,N_5218);
or U7609 (N_7609,N_5005,N_5569);
or U7610 (N_7610,N_5905,N_5301);
nand U7611 (N_7611,N_5416,N_4022);
xnor U7612 (N_7612,N_4994,N_5116);
xor U7613 (N_7613,N_5573,N_5697);
nand U7614 (N_7614,N_4091,N_4495);
nand U7615 (N_7615,N_4483,N_5424);
or U7616 (N_7616,N_4957,N_4802);
xnor U7617 (N_7617,N_4742,N_4982);
and U7618 (N_7618,N_4057,N_4016);
or U7619 (N_7619,N_5259,N_4342);
xnor U7620 (N_7620,N_5685,N_4013);
nor U7621 (N_7621,N_4337,N_4391);
or U7622 (N_7622,N_5866,N_4639);
xor U7623 (N_7623,N_4180,N_5589);
nand U7624 (N_7624,N_4706,N_5742);
nor U7625 (N_7625,N_4836,N_5720);
or U7626 (N_7626,N_5756,N_4478);
and U7627 (N_7627,N_4657,N_5641);
xnor U7628 (N_7628,N_4227,N_5172);
xor U7629 (N_7629,N_4081,N_5586);
nand U7630 (N_7630,N_5344,N_5154);
xnor U7631 (N_7631,N_4507,N_5289);
and U7632 (N_7632,N_4218,N_4806);
or U7633 (N_7633,N_4332,N_4776);
xnor U7634 (N_7634,N_5693,N_4253);
or U7635 (N_7635,N_4154,N_5113);
xnor U7636 (N_7636,N_5702,N_5298);
or U7637 (N_7637,N_5902,N_5690);
nor U7638 (N_7638,N_5251,N_4173);
and U7639 (N_7639,N_4974,N_4958);
nor U7640 (N_7640,N_5402,N_5220);
xnor U7641 (N_7641,N_4789,N_5133);
nand U7642 (N_7642,N_5710,N_4279);
nand U7643 (N_7643,N_5130,N_5539);
nor U7644 (N_7644,N_4262,N_4298);
nor U7645 (N_7645,N_5283,N_5384);
and U7646 (N_7646,N_5857,N_5140);
or U7647 (N_7647,N_5402,N_5017);
nand U7648 (N_7648,N_5572,N_4679);
nand U7649 (N_7649,N_4732,N_5513);
xor U7650 (N_7650,N_5590,N_4838);
or U7651 (N_7651,N_4412,N_5397);
nand U7652 (N_7652,N_4169,N_5867);
xnor U7653 (N_7653,N_5015,N_5600);
and U7654 (N_7654,N_4123,N_5544);
and U7655 (N_7655,N_5542,N_5141);
or U7656 (N_7656,N_4648,N_4264);
xor U7657 (N_7657,N_4245,N_5797);
nor U7658 (N_7658,N_5600,N_4459);
xnor U7659 (N_7659,N_4952,N_4867);
and U7660 (N_7660,N_4809,N_5626);
nand U7661 (N_7661,N_5311,N_5758);
xnor U7662 (N_7662,N_5226,N_4529);
and U7663 (N_7663,N_5223,N_4235);
or U7664 (N_7664,N_5449,N_5003);
and U7665 (N_7665,N_4024,N_4348);
and U7666 (N_7666,N_4485,N_5425);
or U7667 (N_7667,N_4604,N_4860);
or U7668 (N_7668,N_5845,N_5074);
or U7669 (N_7669,N_5748,N_5581);
nand U7670 (N_7670,N_4087,N_5093);
and U7671 (N_7671,N_5602,N_5445);
nor U7672 (N_7672,N_4792,N_5909);
xor U7673 (N_7673,N_5379,N_4284);
or U7674 (N_7674,N_5411,N_5874);
or U7675 (N_7675,N_5387,N_5296);
nor U7676 (N_7676,N_4896,N_4794);
nand U7677 (N_7677,N_5267,N_4541);
nor U7678 (N_7678,N_4845,N_4110);
nand U7679 (N_7679,N_4046,N_4665);
xor U7680 (N_7680,N_5516,N_5688);
nor U7681 (N_7681,N_4492,N_4477);
or U7682 (N_7682,N_5112,N_4911);
nor U7683 (N_7683,N_5781,N_5637);
xor U7684 (N_7684,N_5059,N_4114);
nor U7685 (N_7685,N_4515,N_4658);
and U7686 (N_7686,N_4510,N_5947);
xnor U7687 (N_7687,N_4161,N_5245);
or U7688 (N_7688,N_5700,N_4598);
and U7689 (N_7689,N_5670,N_5657);
and U7690 (N_7690,N_4194,N_4453);
nand U7691 (N_7691,N_5932,N_5702);
nor U7692 (N_7692,N_4760,N_5442);
or U7693 (N_7693,N_5459,N_4750);
or U7694 (N_7694,N_4487,N_5570);
nor U7695 (N_7695,N_5938,N_5689);
xor U7696 (N_7696,N_5768,N_5749);
nand U7697 (N_7697,N_5428,N_4837);
or U7698 (N_7698,N_4755,N_4960);
or U7699 (N_7699,N_4022,N_4202);
and U7700 (N_7700,N_4547,N_5015);
xnor U7701 (N_7701,N_4722,N_4227);
nand U7702 (N_7702,N_4754,N_5615);
nor U7703 (N_7703,N_4581,N_5401);
and U7704 (N_7704,N_5127,N_5716);
or U7705 (N_7705,N_4021,N_4578);
nor U7706 (N_7706,N_4470,N_5977);
nor U7707 (N_7707,N_5044,N_4238);
and U7708 (N_7708,N_4371,N_4191);
or U7709 (N_7709,N_4872,N_4176);
or U7710 (N_7710,N_5254,N_5619);
xnor U7711 (N_7711,N_4981,N_4160);
nand U7712 (N_7712,N_5786,N_5364);
xor U7713 (N_7713,N_5871,N_4119);
nand U7714 (N_7714,N_5477,N_5880);
and U7715 (N_7715,N_4625,N_5631);
xnor U7716 (N_7716,N_4758,N_4321);
nor U7717 (N_7717,N_4232,N_5017);
xor U7718 (N_7718,N_5168,N_4118);
nor U7719 (N_7719,N_4794,N_4233);
nor U7720 (N_7720,N_5721,N_4742);
nor U7721 (N_7721,N_5337,N_4239);
nor U7722 (N_7722,N_5951,N_4381);
or U7723 (N_7723,N_4856,N_5295);
nand U7724 (N_7724,N_5139,N_5548);
nand U7725 (N_7725,N_4876,N_5222);
nand U7726 (N_7726,N_5021,N_5201);
nor U7727 (N_7727,N_5821,N_5676);
or U7728 (N_7728,N_5066,N_5710);
nor U7729 (N_7729,N_4271,N_4053);
and U7730 (N_7730,N_4893,N_5279);
or U7731 (N_7731,N_5760,N_4263);
and U7732 (N_7732,N_4297,N_5094);
and U7733 (N_7733,N_5619,N_4733);
nor U7734 (N_7734,N_5860,N_5901);
xor U7735 (N_7735,N_5675,N_5372);
xnor U7736 (N_7736,N_4756,N_4128);
nand U7737 (N_7737,N_4760,N_4886);
and U7738 (N_7738,N_5786,N_4406);
xnor U7739 (N_7739,N_4606,N_4331);
nand U7740 (N_7740,N_5914,N_5510);
or U7741 (N_7741,N_5631,N_4969);
xor U7742 (N_7742,N_5155,N_4054);
or U7743 (N_7743,N_4492,N_5934);
nor U7744 (N_7744,N_4293,N_5385);
nand U7745 (N_7745,N_4628,N_5489);
nor U7746 (N_7746,N_4661,N_4573);
nor U7747 (N_7747,N_5032,N_4013);
and U7748 (N_7748,N_5969,N_4168);
nor U7749 (N_7749,N_5676,N_4953);
nand U7750 (N_7750,N_5233,N_5512);
xor U7751 (N_7751,N_5924,N_5827);
xor U7752 (N_7752,N_5380,N_4799);
and U7753 (N_7753,N_5121,N_5966);
nor U7754 (N_7754,N_5706,N_4290);
and U7755 (N_7755,N_5393,N_5932);
nand U7756 (N_7756,N_4422,N_4641);
and U7757 (N_7757,N_5029,N_5099);
nand U7758 (N_7758,N_4289,N_4272);
and U7759 (N_7759,N_4874,N_5926);
xor U7760 (N_7760,N_5352,N_5452);
nand U7761 (N_7761,N_4996,N_5721);
or U7762 (N_7762,N_4711,N_4815);
and U7763 (N_7763,N_5100,N_5660);
and U7764 (N_7764,N_4281,N_5913);
and U7765 (N_7765,N_5011,N_5662);
nand U7766 (N_7766,N_5940,N_4929);
or U7767 (N_7767,N_4483,N_4999);
nor U7768 (N_7768,N_4884,N_4375);
and U7769 (N_7769,N_5925,N_5287);
nor U7770 (N_7770,N_5279,N_5804);
xnor U7771 (N_7771,N_4440,N_5693);
and U7772 (N_7772,N_4121,N_5466);
or U7773 (N_7773,N_4182,N_5546);
or U7774 (N_7774,N_5034,N_4652);
xor U7775 (N_7775,N_5145,N_4471);
or U7776 (N_7776,N_5882,N_5394);
nand U7777 (N_7777,N_4199,N_5284);
and U7778 (N_7778,N_4084,N_5604);
nand U7779 (N_7779,N_5662,N_5076);
and U7780 (N_7780,N_4604,N_5301);
and U7781 (N_7781,N_4319,N_5863);
nand U7782 (N_7782,N_5595,N_5951);
and U7783 (N_7783,N_4862,N_5303);
and U7784 (N_7784,N_4113,N_5201);
nand U7785 (N_7785,N_5106,N_4670);
xor U7786 (N_7786,N_4621,N_4078);
nand U7787 (N_7787,N_4200,N_5875);
and U7788 (N_7788,N_5411,N_4556);
nand U7789 (N_7789,N_4855,N_4389);
and U7790 (N_7790,N_4505,N_5692);
xnor U7791 (N_7791,N_5645,N_4775);
nor U7792 (N_7792,N_4634,N_5370);
or U7793 (N_7793,N_5500,N_5528);
and U7794 (N_7794,N_4196,N_4463);
nand U7795 (N_7795,N_5137,N_4439);
and U7796 (N_7796,N_4192,N_5004);
nand U7797 (N_7797,N_5456,N_4359);
nor U7798 (N_7798,N_4099,N_5471);
nor U7799 (N_7799,N_4918,N_5218);
nand U7800 (N_7800,N_5602,N_4854);
xnor U7801 (N_7801,N_5797,N_4851);
xor U7802 (N_7802,N_4829,N_4889);
nor U7803 (N_7803,N_4302,N_4719);
nand U7804 (N_7804,N_4609,N_5372);
xnor U7805 (N_7805,N_4822,N_4642);
nand U7806 (N_7806,N_4446,N_5625);
nor U7807 (N_7807,N_5316,N_5449);
and U7808 (N_7808,N_5146,N_5921);
xor U7809 (N_7809,N_4475,N_4962);
or U7810 (N_7810,N_4018,N_4924);
nor U7811 (N_7811,N_4068,N_4625);
and U7812 (N_7812,N_5608,N_4326);
nor U7813 (N_7813,N_5325,N_5317);
xor U7814 (N_7814,N_4215,N_5339);
and U7815 (N_7815,N_5018,N_4805);
and U7816 (N_7816,N_5058,N_4927);
xor U7817 (N_7817,N_4907,N_4094);
and U7818 (N_7818,N_4112,N_4304);
xor U7819 (N_7819,N_5346,N_4281);
nand U7820 (N_7820,N_5949,N_5825);
nand U7821 (N_7821,N_5790,N_4692);
nor U7822 (N_7822,N_5714,N_5530);
or U7823 (N_7823,N_5962,N_5166);
and U7824 (N_7824,N_4330,N_5257);
nor U7825 (N_7825,N_4545,N_4089);
nor U7826 (N_7826,N_5638,N_4628);
nor U7827 (N_7827,N_4047,N_5314);
and U7828 (N_7828,N_5904,N_5614);
xnor U7829 (N_7829,N_5024,N_4336);
or U7830 (N_7830,N_4700,N_4035);
nor U7831 (N_7831,N_5859,N_4768);
or U7832 (N_7832,N_4025,N_5054);
and U7833 (N_7833,N_4891,N_5947);
nor U7834 (N_7834,N_4440,N_4850);
nand U7835 (N_7835,N_4945,N_4797);
xor U7836 (N_7836,N_4483,N_5864);
nand U7837 (N_7837,N_5340,N_4876);
or U7838 (N_7838,N_5172,N_4787);
nand U7839 (N_7839,N_5895,N_5366);
nor U7840 (N_7840,N_4554,N_5465);
nand U7841 (N_7841,N_5408,N_4151);
and U7842 (N_7842,N_5849,N_5041);
or U7843 (N_7843,N_4732,N_4746);
nand U7844 (N_7844,N_5620,N_4538);
or U7845 (N_7845,N_5489,N_4415);
and U7846 (N_7846,N_4452,N_4372);
or U7847 (N_7847,N_5754,N_5239);
nand U7848 (N_7848,N_5066,N_5922);
xnor U7849 (N_7849,N_5157,N_5970);
nand U7850 (N_7850,N_5717,N_4493);
or U7851 (N_7851,N_4869,N_5528);
xor U7852 (N_7852,N_4146,N_5764);
and U7853 (N_7853,N_4255,N_4733);
xnor U7854 (N_7854,N_5870,N_5527);
and U7855 (N_7855,N_4407,N_4234);
or U7856 (N_7856,N_4648,N_4616);
and U7857 (N_7857,N_5007,N_5355);
or U7858 (N_7858,N_4199,N_4316);
nor U7859 (N_7859,N_4489,N_4932);
nor U7860 (N_7860,N_4567,N_4809);
xor U7861 (N_7861,N_4338,N_5617);
xnor U7862 (N_7862,N_5596,N_5069);
nor U7863 (N_7863,N_5153,N_4219);
and U7864 (N_7864,N_4097,N_4867);
or U7865 (N_7865,N_4219,N_4371);
nor U7866 (N_7866,N_5990,N_4511);
nor U7867 (N_7867,N_5328,N_4190);
and U7868 (N_7868,N_4500,N_4536);
and U7869 (N_7869,N_5210,N_4804);
nand U7870 (N_7870,N_4465,N_5632);
nand U7871 (N_7871,N_5371,N_5701);
nand U7872 (N_7872,N_5156,N_4815);
nor U7873 (N_7873,N_4339,N_5562);
and U7874 (N_7874,N_4402,N_5823);
xnor U7875 (N_7875,N_5936,N_5440);
xor U7876 (N_7876,N_4507,N_4340);
nor U7877 (N_7877,N_5138,N_4215);
nor U7878 (N_7878,N_4097,N_5947);
nand U7879 (N_7879,N_5767,N_5274);
or U7880 (N_7880,N_4257,N_5082);
nor U7881 (N_7881,N_5506,N_4571);
nor U7882 (N_7882,N_5121,N_5679);
or U7883 (N_7883,N_5299,N_4288);
or U7884 (N_7884,N_5145,N_5226);
and U7885 (N_7885,N_4218,N_5800);
and U7886 (N_7886,N_5287,N_4070);
nor U7887 (N_7887,N_5720,N_5257);
xor U7888 (N_7888,N_4838,N_4919);
or U7889 (N_7889,N_5872,N_4111);
xnor U7890 (N_7890,N_5572,N_4234);
nand U7891 (N_7891,N_4672,N_5022);
nand U7892 (N_7892,N_4033,N_5610);
or U7893 (N_7893,N_4995,N_4362);
nand U7894 (N_7894,N_5579,N_4173);
or U7895 (N_7895,N_5476,N_4857);
and U7896 (N_7896,N_5574,N_5853);
or U7897 (N_7897,N_5343,N_4240);
or U7898 (N_7898,N_4773,N_5402);
and U7899 (N_7899,N_4789,N_5220);
or U7900 (N_7900,N_4571,N_5364);
or U7901 (N_7901,N_5235,N_5148);
nor U7902 (N_7902,N_4543,N_5079);
nor U7903 (N_7903,N_5573,N_5752);
xnor U7904 (N_7904,N_4257,N_4878);
or U7905 (N_7905,N_4389,N_4706);
and U7906 (N_7906,N_5060,N_4490);
or U7907 (N_7907,N_5001,N_5635);
and U7908 (N_7908,N_5938,N_5199);
xnor U7909 (N_7909,N_4612,N_5823);
nand U7910 (N_7910,N_5407,N_4444);
and U7911 (N_7911,N_5494,N_4870);
and U7912 (N_7912,N_4341,N_5948);
nand U7913 (N_7913,N_5026,N_4946);
and U7914 (N_7914,N_4165,N_5425);
xor U7915 (N_7915,N_4847,N_4990);
or U7916 (N_7916,N_5315,N_5140);
xor U7917 (N_7917,N_5234,N_5183);
and U7918 (N_7918,N_4025,N_5967);
nor U7919 (N_7919,N_5690,N_4423);
xnor U7920 (N_7920,N_4416,N_4464);
or U7921 (N_7921,N_5597,N_4546);
nand U7922 (N_7922,N_5540,N_4253);
and U7923 (N_7923,N_4957,N_4209);
nand U7924 (N_7924,N_4903,N_5569);
nor U7925 (N_7925,N_5859,N_5799);
or U7926 (N_7926,N_4708,N_5154);
and U7927 (N_7927,N_4812,N_4568);
or U7928 (N_7928,N_4640,N_5288);
nand U7929 (N_7929,N_5689,N_5484);
xor U7930 (N_7930,N_5064,N_5021);
nand U7931 (N_7931,N_4696,N_4716);
or U7932 (N_7932,N_4722,N_5963);
xnor U7933 (N_7933,N_5214,N_5567);
nor U7934 (N_7934,N_4407,N_4396);
xor U7935 (N_7935,N_4713,N_4704);
and U7936 (N_7936,N_4212,N_5671);
and U7937 (N_7937,N_5989,N_4385);
nand U7938 (N_7938,N_5186,N_4510);
and U7939 (N_7939,N_4679,N_5618);
or U7940 (N_7940,N_5763,N_4835);
nor U7941 (N_7941,N_4029,N_4987);
nor U7942 (N_7942,N_5519,N_4666);
or U7943 (N_7943,N_5284,N_4125);
nor U7944 (N_7944,N_4885,N_5613);
xnor U7945 (N_7945,N_5774,N_4158);
xor U7946 (N_7946,N_4244,N_4692);
xor U7947 (N_7947,N_5821,N_5369);
and U7948 (N_7948,N_5877,N_4427);
nor U7949 (N_7949,N_5972,N_5019);
or U7950 (N_7950,N_5290,N_4083);
nand U7951 (N_7951,N_4988,N_5848);
nor U7952 (N_7952,N_4361,N_5536);
or U7953 (N_7953,N_4734,N_5127);
or U7954 (N_7954,N_4668,N_4524);
nor U7955 (N_7955,N_4331,N_5254);
nand U7956 (N_7956,N_4238,N_4329);
nor U7957 (N_7957,N_4390,N_5308);
or U7958 (N_7958,N_4760,N_5277);
or U7959 (N_7959,N_5693,N_5003);
nand U7960 (N_7960,N_5632,N_4801);
nor U7961 (N_7961,N_4183,N_5443);
nor U7962 (N_7962,N_4038,N_4395);
or U7963 (N_7963,N_5785,N_5587);
and U7964 (N_7964,N_5460,N_5764);
nor U7965 (N_7965,N_4072,N_5899);
nand U7966 (N_7966,N_5208,N_4976);
nor U7967 (N_7967,N_5556,N_4098);
nor U7968 (N_7968,N_5216,N_4638);
and U7969 (N_7969,N_4203,N_4289);
nand U7970 (N_7970,N_5131,N_4846);
xor U7971 (N_7971,N_5869,N_4708);
or U7972 (N_7972,N_4085,N_4710);
nor U7973 (N_7973,N_5007,N_5794);
nor U7974 (N_7974,N_5462,N_4132);
and U7975 (N_7975,N_5692,N_5043);
nor U7976 (N_7976,N_4523,N_5699);
nand U7977 (N_7977,N_5508,N_4191);
or U7978 (N_7978,N_5604,N_5642);
nor U7979 (N_7979,N_5053,N_4771);
or U7980 (N_7980,N_5158,N_5194);
and U7981 (N_7981,N_5607,N_5653);
xnor U7982 (N_7982,N_5550,N_5618);
xnor U7983 (N_7983,N_4270,N_4570);
and U7984 (N_7984,N_5365,N_5451);
and U7985 (N_7985,N_4170,N_5761);
xor U7986 (N_7986,N_4896,N_4105);
nor U7987 (N_7987,N_5090,N_5943);
or U7988 (N_7988,N_4780,N_5205);
xnor U7989 (N_7989,N_4226,N_5096);
xnor U7990 (N_7990,N_4255,N_5477);
and U7991 (N_7991,N_4347,N_4528);
or U7992 (N_7992,N_5296,N_4448);
nand U7993 (N_7993,N_5034,N_5210);
or U7994 (N_7994,N_4036,N_5878);
or U7995 (N_7995,N_4036,N_4044);
and U7996 (N_7996,N_4661,N_4483);
or U7997 (N_7997,N_5007,N_4554);
xnor U7998 (N_7998,N_5950,N_5260);
and U7999 (N_7999,N_5405,N_5107);
nor U8000 (N_8000,N_7055,N_6168);
and U8001 (N_8001,N_7626,N_6859);
and U8002 (N_8002,N_7360,N_7272);
nand U8003 (N_8003,N_6441,N_7015);
xnor U8004 (N_8004,N_6698,N_7357);
nor U8005 (N_8005,N_6406,N_6788);
nand U8006 (N_8006,N_6391,N_6479);
nor U8007 (N_8007,N_7530,N_7314);
nor U8008 (N_8008,N_7579,N_6880);
nand U8009 (N_8009,N_6066,N_6561);
and U8010 (N_8010,N_7044,N_6936);
nand U8011 (N_8011,N_6443,N_7446);
or U8012 (N_8012,N_7866,N_7521);
nor U8013 (N_8013,N_7518,N_6491);
nor U8014 (N_8014,N_7769,N_7766);
and U8015 (N_8015,N_6907,N_7648);
nor U8016 (N_8016,N_6404,N_6694);
or U8017 (N_8017,N_7546,N_6985);
xnor U8018 (N_8018,N_7730,N_6917);
or U8019 (N_8019,N_6972,N_6112);
or U8020 (N_8020,N_6298,N_7768);
and U8021 (N_8021,N_7217,N_7149);
and U8022 (N_8022,N_6249,N_7379);
and U8023 (N_8023,N_7981,N_7673);
xnor U8024 (N_8024,N_7230,N_6199);
xor U8025 (N_8025,N_7133,N_7231);
nand U8026 (N_8026,N_6158,N_7414);
or U8027 (N_8027,N_6733,N_7285);
and U8028 (N_8028,N_7096,N_7065);
xor U8029 (N_8029,N_6242,N_7721);
or U8030 (N_8030,N_7980,N_7933);
nand U8031 (N_8031,N_7099,N_7745);
xor U8032 (N_8032,N_6332,N_6606);
nand U8033 (N_8033,N_7457,N_7195);
or U8034 (N_8034,N_6954,N_6812);
nand U8035 (N_8035,N_7443,N_6712);
or U8036 (N_8036,N_6446,N_6463);
and U8037 (N_8037,N_7860,N_7525);
nor U8038 (N_8038,N_7193,N_6350);
xor U8039 (N_8039,N_7047,N_6292);
xor U8040 (N_8040,N_6182,N_7815);
xnor U8041 (N_8041,N_7958,N_6452);
nand U8042 (N_8042,N_7354,N_7909);
or U8043 (N_8043,N_7078,N_6870);
and U8044 (N_8044,N_6757,N_7853);
and U8045 (N_8045,N_6689,N_6590);
xnor U8046 (N_8046,N_7654,N_7585);
nor U8047 (N_8047,N_6418,N_6204);
and U8048 (N_8048,N_7510,N_6197);
or U8049 (N_8049,N_7083,N_6001);
nand U8050 (N_8050,N_6504,N_6819);
xnor U8051 (N_8051,N_7009,N_6500);
nand U8052 (N_8052,N_7394,N_7624);
xor U8053 (N_8053,N_7448,N_6223);
nand U8054 (N_8054,N_6251,N_7582);
and U8055 (N_8055,N_6594,N_7651);
or U8056 (N_8056,N_7978,N_6064);
nor U8057 (N_8057,N_7556,N_6351);
xor U8058 (N_8058,N_6358,N_7608);
nand U8059 (N_8059,N_6167,N_6850);
nand U8060 (N_8060,N_7577,N_6854);
xnor U8061 (N_8061,N_6513,N_6841);
nand U8062 (N_8062,N_7506,N_7552);
nor U8063 (N_8063,N_6287,N_7772);
nor U8064 (N_8064,N_6727,N_6004);
or U8065 (N_8065,N_6497,N_6495);
and U8066 (N_8066,N_7807,N_6597);
xor U8067 (N_8067,N_7680,N_6960);
xnor U8068 (N_8068,N_7486,N_6533);
and U8069 (N_8069,N_6417,N_7180);
or U8070 (N_8070,N_6373,N_7256);
nand U8071 (N_8071,N_6834,N_7074);
or U8072 (N_8072,N_6011,N_7794);
nand U8073 (N_8073,N_6370,N_6244);
and U8074 (N_8074,N_7062,N_6737);
or U8075 (N_8075,N_7841,N_6282);
and U8076 (N_8076,N_6920,N_7676);
xor U8077 (N_8077,N_7959,N_6840);
and U8078 (N_8078,N_7182,N_7692);
and U8079 (N_8079,N_6403,N_6780);
nor U8080 (N_8080,N_7233,N_7066);
nor U8081 (N_8081,N_7928,N_7305);
xnor U8082 (N_8082,N_7121,N_7063);
xor U8083 (N_8083,N_7811,N_6857);
nor U8084 (N_8084,N_6706,N_6569);
and U8085 (N_8085,N_7198,N_7384);
and U8086 (N_8086,N_6067,N_6746);
and U8087 (N_8087,N_7007,N_7787);
nor U8088 (N_8088,N_7235,N_7310);
nor U8089 (N_8089,N_6277,N_6033);
xnor U8090 (N_8090,N_6240,N_7125);
nor U8091 (N_8091,N_6359,N_7422);
nor U8092 (N_8092,N_6440,N_7567);
nand U8093 (N_8093,N_6486,N_7242);
nor U8094 (N_8094,N_6335,N_6666);
or U8095 (N_8095,N_6255,N_7499);
xnor U8096 (N_8096,N_6133,N_7176);
or U8097 (N_8097,N_7684,N_6631);
xnor U8098 (N_8098,N_7442,N_6794);
and U8099 (N_8099,N_6553,N_7051);
nor U8100 (N_8100,N_6316,N_7327);
nand U8101 (N_8101,N_6580,N_6238);
and U8102 (N_8102,N_6690,N_6506);
or U8103 (N_8103,N_7709,N_6604);
xnor U8104 (N_8104,N_6509,N_7924);
nand U8105 (N_8105,N_6871,N_6341);
nand U8106 (N_8106,N_7631,N_6865);
xnor U8107 (N_8107,N_6113,N_6967);
or U8108 (N_8108,N_6892,N_6600);
or U8109 (N_8109,N_7126,N_6475);
xor U8110 (N_8110,N_6900,N_7090);
or U8111 (N_8111,N_7696,N_6123);
and U8112 (N_8112,N_6888,N_6534);
xnor U8113 (N_8113,N_6328,N_7480);
nand U8114 (N_8114,N_6275,N_6056);
and U8115 (N_8115,N_6237,N_6775);
and U8116 (N_8116,N_7087,N_6020);
nor U8117 (N_8117,N_6924,N_6320);
nand U8118 (N_8118,N_6827,N_7398);
and U8119 (N_8119,N_6709,N_7297);
nor U8120 (N_8120,N_6037,N_6667);
nor U8121 (N_8121,N_7473,N_6602);
and U8122 (N_8122,N_6648,N_7010);
nand U8123 (N_8123,N_6679,N_7560);
nand U8124 (N_8124,N_7376,N_7395);
nor U8125 (N_8125,N_7254,N_6609);
or U8126 (N_8126,N_7966,N_6863);
and U8127 (N_8127,N_6550,N_6318);
or U8128 (N_8128,N_6405,N_7344);
and U8129 (N_8129,N_6633,N_6085);
nand U8130 (N_8130,N_7955,N_6266);
nor U8131 (N_8131,N_6490,N_7349);
or U8132 (N_8132,N_6458,N_6416);
nand U8133 (N_8133,N_6129,N_6838);
nor U8134 (N_8134,N_7904,N_7366);
xnor U8135 (N_8135,N_6473,N_7819);
and U8136 (N_8136,N_6055,N_7323);
xnor U8137 (N_8137,N_6540,N_7914);
xor U8138 (N_8138,N_6544,N_7814);
nand U8139 (N_8139,N_7246,N_7210);
nand U8140 (N_8140,N_7779,N_7412);
nor U8141 (N_8141,N_6369,N_7653);
xnor U8142 (N_8142,N_6673,N_6505);
nor U8143 (N_8143,N_6869,N_7979);
and U8144 (N_8144,N_7754,N_7547);
nor U8145 (N_8145,N_7257,N_7565);
nand U8146 (N_8146,N_6754,N_6315);
or U8147 (N_8147,N_6984,N_7559);
nor U8148 (N_8148,N_6937,N_6658);
xor U8149 (N_8149,N_6312,N_7963);
nor U8150 (N_8150,N_7408,N_7820);
nand U8151 (N_8151,N_7570,N_6045);
xnor U8152 (N_8152,N_7250,N_6245);
or U8153 (N_8153,N_6239,N_6778);
xor U8154 (N_8154,N_7621,N_6567);
or U8155 (N_8155,N_6512,N_7620);
xor U8156 (N_8156,N_7377,N_6231);
nand U8157 (N_8157,N_6285,N_6736);
and U8158 (N_8158,N_6910,N_6090);
nor U8159 (N_8159,N_7759,N_6467);
nor U8160 (N_8160,N_6217,N_7645);
nand U8161 (N_8161,N_7659,N_6683);
nor U8162 (N_8162,N_7699,N_7861);
and U8163 (N_8163,N_6030,N_7564);
and U8164 (N_8164,N_6041,N_6200);
nor U8165 (N_8165,N_7497,N_6205);
xor U8166 (N_8166,N_7163,N_7846);
nand U8167 (N_8167,N_7590,N_6799);
xor U8168 (N_8168,N_6570,N_6568);
nand U8169 (N_8169,N_6691,N_7054);
nand U8170 (N_8170,N_7165,N_6970);
nor U8171 (N_8171,N_6957,N_7484);
nor U8172 (N_8172,N_6088,N_7939);
nor U8173 (N_8173,N_7469,N_7736);
or U8174 (N_8174,N_6319,N_6574);
nand U8175 (N_8175,N_7781,N_7409);
and U8176 (N_8176,N_6524,N_6198);
nand U8177 (N_8177,N_6248,N_6881);
and U8178 (N_8178,N_7622,N_6148);
and U8179 (N_8179,N_6010,N_6966);
and U8180 (N_8180,N_6246,N_6663);
xnor U8181 (N_8181,N_6224,N_6081);
or U8182 (N_8182,N_6147,N_6087);
nand U8183 (N_8183,N_6571,N_7361);
or U8184 (N_8184,N_7027,N_6848);
and U8185 (N_8185,N_6708,N_6686);
xor U8186 (N_8186,N_6145,N_6276);
and U8187 (N_8187,N_6034,N_7840);
nand U8188 (N_8188,N_6955,N_6435);
nor U8189 (N_8189,N_6053,N_7304);
nand U8190 (N_8190,N_6759,N_7464);
or U8191 (N_8191,N_7971,N_7568);
or U8192 (N_8192,N_6127,N_7399);
and U8193 (N_8193,N_7501,N_7184);
nand U8194 (N_8194,N_7378,N_6563);
and U8195 (N_8195,N_6024,N_7527);
and U8196 (N_8196,N_7786,N_7161);
or U8197 (N_8197,N_6998,N_6517);
nor U8198 (N_8198,N_6894,N_6449);
or U8199 (N_8199,N_7474,N_7397);
and U8200 (N_8200,N_7504,N_6201);
xnor U8201 (N_8201,N_6921,N_6846);
nand U8202 (N_8202,N_7940,N_6372);
nor U8203 (N_8203,N_6185,N_6539);
xor U8204 (N_8204,N_6395,N_6329);
and U8205 (N_8205,N_7531,N_7538);
nor U8206 (N_8206,N_7902,N_6161);
or U8207 (N_8207,N_7179,N_6125);
xnor U8208 (N_8208,N_6742,N_7459);
nor U8209 (N_8209,N_6430,N_6758);
and U8210 (N_8210,N_6236,N_7657);
xor U8211 (N_8211,N_6766,N_7910);
nand U8212 (N_8212,N_6194,N_7701);
nor U8213 (N_8213,N_6434,N_7028);
xor U8214 (N_8214,N_7875,N_6585);
and U8215 (N_8215,N_7211,N_7308);
xor U8216 (N_8216,N_7893,N_6054);
nand U8217 (N_8217,N_6280,N_6428);
nand U8218 (N_8218,N_7346,N_6906);
or U8219 (N_8219,N_6284,N_7957);
xor U8220 (N_8220,N_7338,N_6557);
xnor U8221 (N_8221,N_7762,N_7301);
or U8222 (N_8222,N_6962,N_6288);
and U8223 (N_8223,N_6904,N_6617);
xnor U8224 (N_8224,N_6000,N_6105);
and U8225 (N_8225,N_6106,N_7899);
or U8226 (N_8226,N_7618,N_7625);
or U8227 (N_8227,N_6741,N_6187);
nand U8228 (N_8228,N_6172,N_7000);
nand U8229 (N_8229,N_6485,N_7404);
or U8230 (N_8230,N_6950,N_7452);
nand U8231 (N_8231,N_7136,N_6809);
or U8232 (N_8232,N_6965,N_6656);
xor U8233 (N_8233,N_6987,N_6971);
and U8234 (N_8234,N_7646,N_7302);
nor U8235 (N_8235,N_6747,N_7502);
nor U8236 (N_8236,N_7453,N_7528);
or U8237 (N_8237,N_7091,N_7732);
nor U8238 (N_8238,N_6547,N_6649);
xnor U8239 (N_8239,N_7386,N_7401);
and U8240 (N_8240,N_6993,N_6979);
or U8241 (N_8241,N_7061,N_7444);
and U8242 (N_8242,N_6379,N_7849);
nand U8243 (N_8243,N_6877,N_6636);
nand U8244 (N_8244,N_7471,N_7884);
nand U8245 (N_8245,N_6577,N_7333);
xnor U8246 (N_8246,N_6874,N_7148);
or U8247 (N_8247,N_7557,N_6908);
or U8248 (N_8248,N_6218,N_6589);
nand U8249 (N_8249,N_7870,N_7783);
and U8250 (N_8250,N_7192,N_7705);
nor U8251 (N_8251,N_6228,N_7277);
or U8252 (N_8252,N_6879,N_6815);
or U8253 (N_8253,N_6327,N_7877);
or U8254 (N_8254,N_6437,N_6143);
nand U8255 (N_8255,N_7587,N_6952);
xor U8256 (N_8256,N_6535,N_7809);
nor U8257 (N_8257,N_7319,N_7005);
xnor U8258 (N_8258,N_6104,N_6501);
nor U8259 (N_8259,N_6009,N_6029);
nand U8260 (N_8260,N_7837,N_7454);
xor U8261 (N_8261,N_6492,N_7985);
nor U8262 (N_8262,N_7173,N_6233);
nand U8263 (N_8263,N_6890,N_6202);
nor U8264 (N_8264,N_6752,N_7220);
and U8265 (N_8265,N_7868,N_7381);
or U8266 (N_8266,N_6885,N_6750);
nand U8267 (N_8267,N_7773,N_7503);
or U8268 (N_8268,N_6420,N_7390);
xnor U8269 (N_8269,N_7019,N_7239);
nand U8270 (N_8270,N_7498,N_7900);
or U8271 (N_8271,N_7132,N_7389);
nor U8272 (N_8272,N_6257,N_7418);
and U8273 (N_8273,N_6447,N_6873);
nand U8274 (N_8274,N_7923,N_7135);
and U8275 (N_8275,N_6831,N_7992);
or U8276 (N_8276,N_7864,N_7831);
and U8277 (N_8277,N_7541,N_7104);
nand U8278 (N_8278,N_6933,N_7533);
and U8279 (N_8279,N_6072,N_7611);
xor U8280 (N_8280,N_7094,N_7101);
nor U8281 (N_8281,N_6387,N_6942);
nand U8282 (N_8282,N_7874,N_7403);
nor U8283 (N_8283,N_6682,N_6354);
nor U8284 (N_8284,N_7245,N_7388);
and U8285 (N_8285,N_6426,N_6414);
and U8286 (N_8286,N_6536,N_7964);
nor U8287 (N_8287,N_7679,N_7013);
nand U8288 (N_8288,N_6652,N_7002);
and U8289 (N_8289,N_7725,N_7563);
and U8290 (N_8290,N_7986,N_7895);
nor U8291 (N_8291,N_6355,N_7150);
xor U8292 (N_8292,N_7001,N_6456);
nor U8293 (N_8293,N_6300,N_6849);
xor U8294 (N_8294,N_6400,N_7634);
and U8295 (N_8295,N_6681,N_6520);
or U8296 (N_8296,N_6804,N_6175);
nand U8297 (N_8297,N_6660,N_7727);
and U8298 (N_8298,N_7458,N_6362);
nand U8299 (N_8299,N_7993,N_6675);
or U8300 (N_8300,N_7279,N_7025);
nor U8301 (N_8301,N_6272,N_7850);
xor U8302 (N_8302,N_6502,N_7463);
or U8303 (N_8303,N_7115,N_7778);
nor U8304 (N_8304,N_7050,N_6796);
nand U8305 (N_8305,N_6707,N_6614);
nor U8306 (N_8306,N_7347,N_6012);
nand U8307 (N_8307,N_7919,N_7224);
nand U8308 (N_8308,N_7812,N_7669);
and U8309 (N_8309,N_6605,N_7298);
nor U8310 (N_8310,N_7561,N_6186);
and U8311 (N_8311,N_7908,N_6554);
and U8312 (N_8312,N_6220,N_7507);
or U8313 (N_8313,N_6940,N_6058);
xor U8314 (N_8314,N_6408,N_6964);
and U8315 (N_8315,N_6532,N_6668);
xnor U8316 (N_8316,N_6619,N_6260);
xor U8317 (N_8317,N_6091,N_6719);
xor U8318 (N_8318,N_6717,N_6922);
and U8319 (N_8319,N_6883,N_6703);
xor U8320 (N_8320,N_6803,N_6586);
nor U8321 (N_8321,N_7177,N_6325);
and U8322 (N_8322,N_7894,N_7380);
nor U8323 (N_8323,N_7470,N_6165);
xnor U8324 (N_8324,N_6474,N_7689);
nand U8325 (N_8325,N_6762,N_7977);
or U8326 (N_8326,N_6089,N_7070);
xor U8327 (N_8327,N_6286,N_6084);
nand U8328 (N_8328,N_7273,N_7006);
and U8329 (N_8329,N_6781,N_6195);
and U8330 (N_8330,N_7776,N_6499);
xnor U8331 (N_8331,N_7041,N_7640);
nor U8332 (N_8332,N_6525,N_6862);
nor U8333 (N_8333,N_6575,N_7374);
and U8334 (N_8334,N_6530,N_7243);
xor U8335 (N_8335,N_6232,N_7675);
xor U8336 (N_8336,N_7566,N_7915);
and U8337 (N_8337,N_6748,N_7606);
xnor U8338 (N_8338,N_6203,N_7822);
nand U8339 (N_8339,N_7667,N_6121);
or U8340 (N_8340,N_6969,N_6538);
and U8341 (N_8341,N_6496,N_6612);
xor U8342 (N_8342,N_7584,N_7854);
nand U8343 (N_8343,N_7712,N_6137);
nor U8344 (N_8344,N_6744,N_7797);
xnor U8345 (N_8345,N_7268,N_7748);
nor U8346 (N_8346,N_6444,N_7828);
nor U8347 (N_8347,N_7529,N_6025);
nor U8348 (N_8348,N_6386,N_6896);
or U8349 (N_8349,N_6753,N_6839);
or U8350 (N_8350,N_7810,N_6262);
nand U8351 (N_8351,N_6323,N_6982);
nand U8352 (N_8352,N_7800,N_6156);
and U8353 (N_8353,N_6886,N_6626);
and U8354 (N_8354,N_6738,N_7367);
xor U8355 (N_8355,N_6837,N_7229);
xor U8356 (N_8356,N_7102,N_7953);
or U8357 (N_8357,N_6996,N_6192);
nand U8358 (N_8358,N_7545,N_7283);
nor U8359 (N_8359,N_6043,N_6776);
nand U8360 (N_8360,N_6322,N_6770);
and U8361 (N_8361,N_7335,N_7973);
xor U8362 (N_8362,N_7665,N_7801);
or U8363 (N_8363,N_7802,N_6346);
or U8364 (N_8364,N_7260,N_7432);
or U8365 (N_8365,N_7972,N_6075);
or U8366 (N_8366,N_6047,N_7716);
nand U8367 (N_8367,N_6740,N_7630);
and U8368 (N_8368,N_7505,N_6716);
or U8369 (N_8369,N_6378,N_7071);
nand U8370 (N_8370,N_7097,N_7643);
or U8371 (N_8371,N_6992,N_6432);
nor U8372 (N_8372,N_6274,N_7700);
xnor U8373 (N_8373,N_6642,N_7312);
nand U8374 (N_8374,N_7780,N_6234);
or U8375 (N_8375,N_7281,N_6270);
nor U8376 (N_8376,N_7826,N_6273);
nand U8377 (N_8377,N_6258,N_6542);
nor U8378 (N_8378,N_7106,N_6196);
or U8379 (N_8379,N_7652,N_6613);
xnor U8380 (N_8380,N_6431,N_6986);
nand U8381 (N_8381,N_7903,N_7076);
or U8382 (N_8382,N_6817,N_6450);
nor U8383 (N_8383,N_6082,N_7629);
nor U8384 (N_8384,N_6134,N_6665);
or U8385 (N_8385,N_7449,N_6289);
nor U8386 (N_8386,N_7107,N_6988);
nor U8387 (N_8387,N_6564,N_6396);
nand U8388 (N_8388,N_7479,N_7987);
and U8389 (N_8389,N_7114,N_7290);
xor U8390 (N_8390,N_6810,N_7823);
nand U8391 (N_8391,N_6478,N_6730);
or U8392 (N_8392,N_7931,N_6153);
and U8393 (N_8393,N_7164,N_6835);
nand U8394 (N_8394,N_6958,N_7770);
nand U8395 (N_8395,N_6909,N_6997);
and U8396 (N_8396,N_6808,N_6773);
nand U8397 (N_8397,N_7535,N_6206);
and U8398 (N_8398,N_6647,N_7553);
nor U8399 (N_8399,N_6935,N_6421);
or U8400 (N_8400,N_6844,N_7049);
nor U8401 (N_8401,N_7219,N_6704);
nand U8402 (N_8402,N_6402,N_6603);
and U8403 (N_8403,N_7048,N_6928);
or U8404 (N_8404,N_6664,N_7543);
and U8405 (N_8405,N_6826,N_6424);
nand U8406 (N_8406,N_7738,N_7269);
nand U8407 (N_8407,N_7183,N_7339);
nand U8408 (N_8408,N_7155,N_7300);
nand U8409 (N_8409,N_7542,N_7171);
or U8410 (N_8410,N_6410,N_7156);
or U8411 (N_8411,N_7789,N_6913);
and U8412 (N_8412,N_7270,N_6162);
and U8413 (N_8413,N_7859,N_6036);
nand U8414 (N_8414,N_7969,N_6281);
nor U8415 (N_8415,N_7166,N_7878);
or U8416 (N_8416,N_7441,N_7882);
nand U8417 (N_8417,N_6864,N_7571);
xnor U8418 (N_8418,N_6157,N_6477);
nor U8419 (N_8419,N_7843,N_7392);
nand U8420 (N_8420,N_6584,N_6677);
xor U8421 (N_8421,N_7796,N_7004);
and U8422 (N_8422,N_7747,N_7169);
and U8423 (N_8423,N_6930,N_6077);
and U8424 (N_8424,N_7127,N_7580);
and U8425 (N_8425,N_6523,N_7352);
nand U8426 (N_8426,N_7075,N_6301);
and U8427 (N_8427,N_6639,N_7942);
nor U8428 (N_8428,N_6189,N_7282);
nor U8429 (N_8429,N_7003,N_6466);
and U8430 (N_8430,N_6774,N_6763);
and U8431 (N_8431,N_7737,N_7375);
nor U8432 (N_8432,N_7046,N_7739);
xor U8433 (N_8433,N_7920,N_7334);
and U8434 (N_8434,N_7678,N_7633);
or U8435 (N_8435,N_6813,N_7143);
xor U8436 (N_8436,N_7313,N_7317);
nor U8437 (N_8437,N_6498,N_6710);
nor U8438 (N_8438,N_7662,N_7291);
xor U8439 (N_8439,N_7137,N_7687);
and U8440 (N_8440,N_7337,N_7467);
or U8441 (N_8441,N_6313,N_6822);
or U8442 (N_8442,N_6385,N_7370);
xor U8443 (N_8443,N_7039,N_6784);
or U8444 (N_8444,N_7550,N_6901);
xor U8445 (N_8445,N_7461,N_7990);
or U8446 (N_8446,N_7632,N_7068);
or U8447 (N_8447,N_6311,N_6227);
nor U8448 (N_8448,N_7834,N_7941);
xnor U8449 (N_8449,N_7194,N_7974);
nand U8450 (N_8450,N_6638,N_6407);
xnor U8451 (N_8451,N_7214,N_7487);
or U8452 (N_8452,N_6229,N_6915);
xor U8453 (N_8453,N_7753,N_7213);
or U8454 (N_8454,N_7142,N_7212);
nor U8455 (N_8455,N_6916,N_7575);
nand U8456 (N_8456,N_6261,N_6259);
xnor U8457 (N_8457,N_7331,N_7294);
or U8458 (N_8458,N_7330,N_6180);
and U8459 (N_8459,N_7240,N_6887);
nor U8460 (N_8460,N_6096,N_6039);
nor U8461 (N_8461,N_6696,N_6163);
or U8462 (N_8462,N_7022,N_6304);
nand U8463 (N_8463,N_7430,N_6720);
and U8464 (N_8464,N_7615,N_7207);
and U8465 (N_8465,N_6149,N_6295);
and U8466 (N_8466,N_7160,N_6654);
and U8467 (N_8467,N_7650,N_7690);
and U8468 (N_8468,N_7481,N_7715);
xor U8469 (N_8469,N_6061,N_6062);
or U8470 (N_8470,N_6789,N_6761);
nand U8471 (N_8471,N_6023,N_7788);
and U8472 (N_8472,N_7704,N_7594);
xor U8473 (N_8473,N_7572,N_6650);
nor U8474 (N_8474,N_7021,N_7206);
nor U8475 (N_8475,N_7734,N_6963);
nor U8476 (N_8476,N_7706,N_6637);
and U8477 (N_8477,N_7286,N_7623);
and U8478 (N_8478,N_6939,N_6990);
nor U8479 (N_8479,N_7057,N_7029);
and U8480 (N_8480,N_7159,N_7888);
xor U8481 (N_8481,N_7296,N_6383);
or U8482 (N_8482,N_7598,N_7350);
nand U8483 (N_8483,N_7806,N_6307);
and U8484 (N_8484,N_7813,N_6419);
nand U8485 (N_8485,N_7512,N_6546);
or U8486 (N_8486,N_7947,N_7760);
nor U8487 (N_8487,N_7351,N_6050);
nand U8488 (N_8488,N_7905,N_6481);
nor U8489 (N_8489,N_6482,N_7867);
nor U8490 (N_8490,N_7082,N_6427);
or U8491 (N_8491,N_6063,N_7236);
and U8492 (N_8492,N_6715,N_6772);
xnor U8493 (N_8493,N_6688,N_7872);
xor U8494 (N_8494,N_6057,N_6177);
nor U8495 (N_8495,N_6680,N_6035);
xnor U8496 (N_8496,N_7656,N_6537);
and U8497 (N_8497,N_6166,N_7551);
and U8498 (N_8498,N_7140,N_6120);
nand U8499 (N_8499,N_6695,N_6830);
xor U8500 (N_8500,N_6454,N_7170);
xnor U8501 (N_8501,N_7253,N_7897);
or U8502 (N_8502,N_6135,N_6644);
or U8503 (N_8503,N_6949,N_7569);
nor U8504 (N_8504,N_7876,N_6676);
nand U8505 (N_8505,N_6925,N_6413);
or U8506 (N_8506,N_6174,N_6074);
nand U8507 (N_8507,N_6583,N_7103);
and U8508 (N_8508,N_7856,N_6760);
nand U8509 (N_8509,N_6728,N_7707);
or U8510 (N_8510,N_6599,N_7221);
nor U8511 (N_8511,N_7916,N_6208);
and U8512 (N_8512,N_7583,N_7405);
nand U8513 (N_8513,N_6578,N_7758);
or U8514 (N_8514,N_7280,N_7336);
and U8515 (N_8515,N_7508,N_6832);
or U8516 (N_8516,N_7108,N_7713);
xnor U8517 (N_8517,N_7244,N_6548);
nor U8518 (N_8518,N_6828,N_7287);
or U8519 (N_8519,N_7299,N_7666);
nand U8520 (N_8520,N_7764,N_7355);
and U8521 (N_8521,N_7356,N_7948);
xor U8522 (N_8522,N_7597,N_7791);
nor U8523 (N_8523,N_7478,N_6488);
and U8524 (N_8524,N_7638,N_6718);
nor U8525 (N_8525,N_7614,N_7586);
or U8526 (N_8526,N_7775,N_7427);
and U8527 (N_8527,N_6725,N_7952);
and U8528 (N_8528,N_6618,N_6902);
and U8529 (N_8529,N_7549,N_6438);
nor U8530 (N_8530,N_7731,N_6122);
nor U8531 (N_8531,N_6582,N_6805);
and U8532 (N_8532,N_7671,N_7862);
nand U8533 (N_8533,N_7119,N_7724);
or U8534 (N_8534,N_7428,N_7756);
xor U8535 (N_8535,N_7267,N_6337);
nand U8536 (N_8536,N_6471,N_6032);
and U8537 (N_8537,N_7729,N_7733);
nor U8538 (N_8538,N_7134,N_6005);
and U8539 (N_8539,N_7491,N_6390);
xor U8540 (N_8540,N_6433,N_6493);
nor U8541 (N_8541,N_7517,N_6661);
and U8542 (N_8542,N_6627,N_6324);
or U8543 (N_8543,N_6139,N_6006);
xnor U8544 (N_8544,N_7519,N_7237);
or U8545 (N_8545,N_7886,N_7416);
nor U8546 (N_8546,N_7326,N_6836);
or U8547 (N_8547,N_7682,N_6976);
and U8548 (N_8548,N_7146,N_6116);
nand U8549 (N_8549,N_6545,N_7989);
and U8550 (N_8550,N_6843,N_6212);
nor U8551 (N_8551,N_7588,N_6598);
nor U8552 (N_8552,N_7603,N_7555);
and U8553 (N_8553,N_6210,N_6207);
nor U8554 (N_8554,N_7111,N_6184);
and U8555 (N_8555,N_7303,N_6591);
nor U8556 (N_8556,N_6305,N_7954);
nor U8557 (N_8557,N_7639,N_7098);
or U8558 (N_8558,N_6398,N_6008);
or U8559 (N_8559,N_6083,N_6086);
nor U8560 (N_8560,N_7827,N_7918);
and U8561 (N_8561,N_6787,N_6179);
or U8562 (N_8562,N_7472,N_7128);
nand U8563 (N_8563,N_6076,N_6461);
nand U8564 (N_8564,N_6521,N_7020);
xor U8565 (N_8565,N_7836,N_6562);
nand U8566 (N_8566,N_7373,N_7685);
or U8567 (N_8567,N_7289,N_6022);
or U8568 (N_8568,N_6283,N_6136);
xor U8569 (N_8569,N_6171,N_7641);
and U8570 (N_8570,N_6209,N_6144);
xnor U8571 (N_8571,N_6038,N_7493);
or U8572 (N_8572,N_6070,N_7495);
and U8573 (N_8573,N_7263,N_7130);
xnor U8574 (N_8574,N_6847,N_7536);
or U8575 (N_8575,N_7741,N_6154);
xnor U8576 (N_8576,N_6108,N_6103);
or U8577 (N_8577,N_6559,N_6107);
and U8578 (N_8578,N_7628,N_7197);
and U8579 (N_8579,N_7901,N_7642);
or U8580 (N_8580,N_7693,N_7329);
or U8581 (N_8581,N_7785,N_6016);
and U8582 (N_8582,N_6007,N_6051);
nor U8583 (N_8583,N_7938,N_7292);
xor U8584 (N_8584,N_7649,N_6308);
or U8585 (N_8585,N_6994,N_7970);
or U8586 (N_8586,N_7189,N_6518);
nor U8587 (N_8587,N_7249,N_6401);
or U8588 (N_8588,N_7369,N_7147);
nor U8589 (N_8589,N_6342,N_7869);
and U8590 (N_8590,N_6999,N_7309);
nand U8591 (N_8591,N_7994,N_7426);
xor U8592 (N_8592,N_6356,N_7295);
nor U8593 (N_8593,N_7073,N_6150);
xor U8594 (N_8594,N_6230,N_7591);
nor U8595 (N_8595,N_7668,N_6959);
xor U8596 (N_8596,N_7885,N_6141);
nor U8597 (N_8597,N_7548,N_7723);
or U8598 (N_8598,N_7718,N_6455);
nand U8599 (N_8599,N_6643,N_6527);
nor U8600 (N_8600,N_6867,N_7433);
nand U8601 (N_8601,N_7225,N_7613);
nand U8602 (N_8602,N_6181,N_6659);
nor U8603 (N_8603,N_7095,N_6601);
or U8604 (N_8604,N_6825,N_7186);
nor U8605 (N_8605,N_6046,N_6140);
nand U8606 (N_8606,N_7514,N_6309);
or U8607 (N_8607,N_7961,N_7117);
nand U8608 (N_8608,N_7227,N_6884);
nor U8609 (N_8609,N_7848,N_6845);
xnor U8610 (N_8610,N_7275,N_7944);
or U8611 (N_8611,N_6394,N_6480);
xor U8612 (N_8612,N_6243,N_7100);
nand U8613 (N_8613,N_6911,N_7014);
nand U8614 (N_8614,N_6357,N_6267);
nor U8615 (N_8615,N_6934,N_7316);
nor U8616 (N_8616,N_7307,N_7060);
xnor U8617 (N_8617,N_6019,N_6268);
nand U8618 (N_8618,N_7262,N_6336);
nor U8619 (N_8619,N_6556,N_7683);
xor U8620 (N_8620,N_6097,N_6801);
nor U8621 (N_8621,N_6098,N_6795);
nor U8622 (N_8622,N_7576,N_7799);
xor U8623 (N_8623,N_6607,N_6611);
nand U8624 (N_8624,N_6003,N_7907);
xor U8625 (N_8625,N_7997,N_7852);
nor U8626 (N_8626,N_6078,N_7601);
or U8627 (N_8627,N_6290,N_7202);
or U8628 (N_8628,N_7602,N_6729);
and U8629 (N_8629,N_6214,N_6735);
nand U8630 (N_8630,N_7540,N_7832);
xor U8631 (N_8631,N_6655,N_7016);
nand U8632 (N_8632,N_6811,N_6634);
nor U8633 (N_8633,N_6065,N_7691);
or U8634 (N_8634,N_7708,N_7965);
xnor U8635 (N_8635,N_6330,N_6353);
xor U8636 (N_8636,N_6363,N_7085);
or U8637 (N_8637,N_7496,N_6645);
nor U8638 (N_8638,N_6823,N_7241);
or U8639 (N_8639,N_7744,N_6059);
or U8640 (N_8640,N_6615,N_6899);
nor U8641 (N_8641,N_7081,N_7199);
nor U8642 (N_8642,N_6549,N_6824);
nand U8643 (N_8643,N_6344,N_6093);
nand U8644 (N_8644,N_7092,N_6340);
nor U8645 (N_8645,N_7110,N_6953);
nand U8646 (N_8646,N_7228,N_7857);
nor U8647 (N_8647,N_7129,N_7751);
xor U8648 (N_8648,N_7086,N_7113);
and U8649 (N_8649,N_7795,N_7175);
and U8650 (N_8650,N_6114,N_6422);
xor U8651 (N_8651,N_6349,N_6079);
and U8652 (N_8652,N_7943,N_7596);
xnor U8653 (N_8653,N_6415,N_6632);
nand U8654 (N_8654,N_7911,N_7865);
nor U8655 (N_8655,N_7526,N_7742);
xnor U8656 (N_8656,N_7936,N_7674);
xnor U8657 (N_8657,N_6903,N_6635);
or U8658 (N_8658,N_6579,N_6291);
and U8659 (N_8659,N_6095,N_6138);
nor U8660 (N_8660,N_6995,N_7663);
or U8661 (N_8661,N_7537,N_6543);
xor U8662 (N_8662,N_7842,N_7396);
nand U8663 (N_8663,N_6713,N_7205);
nor U8664 (N_8664,N_6678,N_7883);
and U8665 (N_8665,N_7466,N_7429);
or U8666 (N_8666,N_7968,N_6069);
xor U8667 (N_8667,N_7532,N_7363);
nand U8668 (N_8668,N_6503,N_6384);
and U8669 (N_8669,N_7476,N_6221);
nor U8670 (N_8670,N_6861,N_7203);
nor U8671 (N_8671,N_7949,N_7784);
nand U8672 (N_8672,N_6222,N_7364);
xnor U8673 (N_8673,N_7956,N_7157);
or U8674 (N_8674,N_7332,N_6566);
nor U8675 (N_8675,N_7818,N_6769);
and U8676 (N_8676,N_7698,N_6573);
and U8677 (N_8677,N_7012,N_7950);
or U8678 (N_8678,N_6851,N_7581);
or U8679 (N_8679,N_6326,N_6792);
nand U8680 (N_8680,N_7534,N_6929);
nand U8681 (N_8681,N_7222,N_7482);
xnor U8682 (N_8682,N_6219,N_6216);
or U8683 (N_8683,N_6640,N_7516);
or U8684 (N_8684,N_6651,N_6723);
nor U8685 (N_8685,N_7036,N_7382);
nor U8686 (N_8686,N_6352,N_7695);
and U8687 (N_8687,N_6610,N_7991);
nor U8688 (N_8688,N_7607,N_7144);
and U8689 (N_8689,N_6519,N_6947);
nand U8690 (N_8690,N_6592,N_6013);
xor U8691 (N_8691,N_6250,N_6367);
and U8692 (N_8692,N_6178,N_7410);
nor U8693 (N_8693,N_7413,N_7757);
nand U8694 (N_8694,N_6465,N_7328);
nor U8695 (N_8695,N_6853,N_6365);
xnor U8696 (N_8696,N_7320,N_7752);
or U8697 (N_8697,N_7670,N_6302);
xnor U8698 (N_8698,N_6978,N_7131);
nor U8699 (N_8699,N_7520,N_7702);
nand U8700 (N_8700,N_6945,N_7726);
and U8701 (N_8701,N_7763,N_7703);
nand U8702 (N_8702,N_7605,N_7248);
and U8703 (N_8703,N_6510,N_6397);
or U8704 (N_8704,N_7185,N_6923);
xnor U8705 (N_8705,N_7200,N_7926);
and U8706 (N_8706,N_6256,N_7342);
and U8707 (N_8707,N_6779,N_6816);
xnor U8708 (N_8708,N_7168,N_6891);
and U8709 (N_8709,N_6252,N_7644);
nor U8710 (N_8710,N_6856,N_6820);
nand U8711 (N_8711,N_6968,N_6170);
xor U8712 (N_8712,N_7743,N_6684);
nand U8713 (N_8713,N_6464,N_6018);
and U8714 (N_8714,N_6119,N_7322);
nand U8715 (N_8715,N_7825,N_7122);
xor U8716 (N_8716,N_6670,N_6687);
and U8717 (N_8717,N_7031,N_7341);
or U8718 (N_8718,N_6641,N_7321);
and U8719 (N_8719,N_6293,N_7247);
nor U8720 (N_8720,N_7187,N_7999);
xor U8721 (N_8721,N_7523,N_6693);
or U8722 (N_8722,N_7821,N_6278);
xnor U8723 (N_8723,N_7998,N_6371);
and U8724 (N_8724,N_7018,N_6348);
nor U8725 (N_8725,N_7460,N_6983);
nor U8726 (N_8726,N_7930,N_6241);
or U8727 (N_8727,N_7554,N_7072);
nand U8728 (N_8728,N_7483,N_6265);
and U8729 (N_8729,N_7892,N_7714);
or U8730 (N_8730,N_6596,N_7434);
or U8731 (N_8731,N_6476,N_7879);
nor U8732 (N_8732,N_6732,N_6948);
nand U8733 (N_8733,N_7024,N_6818);
or U8734 (N_8734,N_6508,N_6299);
or U8735 (N_8735,N_6470,N_6361);
nor U8736 (N_8736,N_6782,N_6991);
and U8737 (N_8737,N_7647,N_7059);
and U8738 (N_8738,N_7962,N_6646);
nor U8739 (N_8739,N_7138,N_7609);
and U8740 (N_8740,N_7423,N_6927);
nor U8741 (N_8741,N_7816,N_6814);
nand U8742 (N_8742,N_6271,N_7951);
nand U8743 (N_8743,N_7191,N_7251);
nor U8744 (N_8744,N_7040,N_7515);
or U8745 (N_8745,N_6511,N_7844);
and U8746 (N_8746,N_6739,N_7490);
nor U8747 (N_8747,N_7172,N_6526);
nor U8748 (N_8748,N_6731,N_7255);
nor U8749 (N_8749,N_7798,N_6484);
and U8750 (N_8750,N_6176,N_7717);
and U8751 (N_8751,N_6630,N_6132);
xor U8752 (N_8752,N_7358,N_6697);
nor U8753 (N_8753,N_7672,N_6489);
xnor U8754 (N_8754,N_7881,N_6866);
nand U8755 (N_8755,N_6294,N_7077);
nand U8756 (N_8756,N_6528,N_6102);
xnor U8757 (N_8757,N_7562,N_6459);
and U8758 (N_8758,N_6565,N_6588);
xor U8759 (N_8759,N_7340,N_6015);
nand U8760 (N_8760,N_6791,N_7226);
nand U8761 (N_8761,N_7891,N_7439);
nor U8762 (N_8762,N_7921,N_6026);
and U8763 (N_8763,N_7790,N_7873);
and U8764 (N_8764,N_6375,N_6918);
and U8765 (N_8765,N_6875,N_7069);
or U8766 (N_8766,N_6783,N_7468);
xnor U8767 (N_8767,N_7627,N_6980);
nor U8768 (N_8768,N_7477,N_6699);
or U8769 (N_8769,N_6938,N_6572);
nor U8770 (N_8770,N_7445,N_7153);
nand U8771 (N_8771,N_7343,N_7419);
and U8772 (N_8772,N_7406,N_6700);
and U8773 (N_8773,N_7158,N_7151);
or U8774 (N_8774,N_7440,N_7511);
or U8775 (N_8775,N_7318,N_6620);
and U8776 (N_8776,N_7805,N_7407);
and U8777 (N_8777,N_7139,N_7056);
and U8778 (N_8778,N_6462,N_7817);
and U8779 (N_8779,N_7697,N_7089);
xor U8780 (N_8780,N_7324,N_7084);
nor U8781 (N_8781,N_6412,N_6722);
or U8782 (N_8782,N_7424,N_7190);
nor U8783 (N_8783,N_7042,N_7088);
nor U8784 (N_8784,N_6616,N_6897);
nand U8785 (N_8785,N_7365,N_7658);
or U8786 (N_8786,N_7118,N_6932);
and U8787 (N_8787,N_6049,N_7686);
and U8788 (N_8788,N_6975,N_6868);
or U8789 (N_8789,N_6117,N_6188);
nand U8790 (N_8790,N_6515,N_6800);
or U8791 (N_8791,N_7371,N_6701);
nor U8792 (N_8792,N_7402,N_7359);
xor U8793 (N_8793,N_6961,N_7932);
nand U8794 (N_8794,N_7793,N_6073);
xnor U8795 (N_8795,N_6068,N_7887);
xnor U8796 (N_8796,N_7271,N_7635);
and U8797 (N_8797,N_7400,N_7774);
xnor U8798 (N_8798,N_7513,N_6002);
nand U8799 (N_8799,N_7201,N_7234);
and U8800 (N_8800,N_7655,N_6893);
or U8801 (N_8801,N_7539,N_6989);
nor U8802 (N_8802,N_7353,N_7934);
nor U8803 (N_8803,N_6751,N_7694);
and U8804 (N_8804,N_6027,N_7573);
nand U8805 (N_8805,N_6100,N_6388);
nor U8806 (N_8806,N_7593,N_6247);
nand U8807 (N_8807,N_7735,N_7509);
nor U8808 (N_8808,N_7777,N_6882);
and U8809 (N_8809,N_6721,N_6399);
nand U8810 (N_8810,N_6622,N_7578);
and U8811 (N_8811,N_6124,N_6951);
and U8812 (N_8812,N_7711,N_7661);
nor U8813 (N_8813,N_7259,N_7677);
nand U8814 (N_8814,N_6333,N_7284);
or U8815 (N_8815,N_6516,N_6469);
nor U8816 (N_8816,N_6743,N_7619);
xnor U8817 (N_8817,N_6164,N_6514);
nand U8818 (N_8818,N_6558,N_7946);
nor U8819 (N_8819,N_7913,N_6653);
nor U8820 (N_8820,N_6472,N_6052);
nand U8821 (N_8821,N_6889,N_6487);
and U8822 (N_8822,N_6858,N_6755);
nand U8823 (N_8823,N_6842,N_7720);
xor U8824 (N_8824,N_7393,N_6726);
nand U8825 (N_8825,N_7995,N_6852);
nor U8826 (N_8826,N_6802,N_6507);
nand U8827 (N_8827,N_7345,N_6211);
or U8828 (N_8828,N_7437,N_7311);
nand U8829 (N_8829,N_6798,N_6411);
xor U8830 (N_8830,N_7833,N_6253);
nand U8831 (N_8831,N_6031,N_7178);
nand U8832 (N_8832,N_6368,N_6629);
or U8833 (N_8833,N_6806,N_6235);
or U8834 (N_8834,N_7500,N_6360);
nand U8835 (N_8835,N_7362,N_6905);
xor U8836 (N_8836,N_7045,N_6080);
nand U8837 (N_8837,N_7218,N_7456);
or U8838 (N_8838,N_7033,N_6028);
or U8839 (N_8839,N_6442,N_6685);
nor U8840 (N_8840,N_7223,N_7306);
nand U8841 (N_8841,N_7417,N_6745);
nor U8842 (N_8842,N_7937,N_6130);
nor U8843 (N_8843,N_6071,N_6017);
or U8844 (N_8844,N_6541,N_7485);
or U8845 (N_8845,N_7982,N_7851);
nor U8846 (N_8846,N_7975,N_6494);
or U8847 (N_8847,N_7746,N_7890);
nor U8848 (N_8848,N_6674,N_6531);
nor U8849 (N_8849,N_6173,N_7996);
or U8850 (N_8850,N_7372,N_6381);
and U8851 (N_8851,N_6926,N_7368);
xor U8852 (N_8852,N_6956,N_6334);
and U8853 (N_8853,N_7488,N_7765);
nor U8854 (N_8854,N_7767,N_6974);
xnor U8855 (N_8855,N_7425,N_7927);
xnor U8856 (N_8856,N_6560,N_7589);
or U8857 (N_8857,N_6860,N_7824);
nand U8858 (N_8858,N_7436,N_7035);
or U8859 (N_8859,N_6409,N_7258);
nand U8860 (N_8860,N_7415,N_7208);
xor U8861 (N_8861,N_6946,N_6705);
and U8862 (N_8862,N_6833,N_7420);
nor U8863 (N_8863,N_6764,N_7265);
or U8864 (N_8864,N_7196,N_7238);
nand U8865 (N_8865,N_7181,N_7906);
nor U8866 (N_8866,N_6576,N_6451);
nor U8867 (N_8867,N_7855,N_6624);
nor U8868 (N_8868,N_6155,N_6376);
or U8869 (N_8869,N_7935,N_7431);
xnor U8870 (N_8870,N_6587,N_7945);
xnor U8871 (N_8871,N_7984,N_7174);
nor U8872 (N_8872,N_6366,N_7917);
or U8873 (N_8873,N_6931,N_6919);
and U8874 (N_8874,N_6392,N_6448);
and U8875 (N_8875,N_6749,N_7612);
nor U8876 (N_8876,N_7080,N_6159);
xor U8877 (N_8877,N_7558,N_7053);
nand U8878 (N_8878,N_6608,N_6263);
or U8879 (N_8879,N_6042,N_7889);
nand U8880 (N_8880,N_6628,N_6339);
nand U8881 (N_8881,N_7167,N_6393);
and U8882 (N_8882,N_7592,N_6522);
or U8883 (N_8883,N_6110,N_6213);
and U8884 (N_8884,N_7880,N_6439);
xnor U8885 (N_8885,N_7079,N_7276);
xnor U8886 (N_8886,N_6436,N_6215);
xor U8887 (N_8887,N_7188,N_6126);
and U8888 (N_8888,N_6714,N_6183);
xnor U8889 (N_8889,N_7293,N_7216);
or U8890 (N_8890,N_6790,N_6191);
and U8891 (N_8891,N_6807,N_7450);
nand U8892 (N_8892,N_7960,N_7462);
nand U8893 (N_8893,N_6529,N_6555);
xor U8894 (N_8894,N_6895,N_6672);
nand U8895 (N_8895,N_7922,N_6702);
and U8896 (N_8896,N_7023,N_6483);
xnor U8897 (N_8897,N_7266,N_7385);
xnor U8898 (N_8898,N_7710,N_6226);
nor U8899 (N_8899,N_6321,N_7792);
nor U8900 (N_8900,N_6941,N_7116);
xnor U8901 (N_8901,N_6279,N_6765);
nor U8902 (N_8902,N_7052,N_7782);
and U8903 (N_8903,N_6118,N_7983);
xor U8904 (N_8904,N_6382,N_7383);
and U8905 (N_8905,N_7838,N_7835);
and U8906 (N_8906,N_7524,N_7610);
or U8907 (N_8907,N_6146,N_6460);
and U8908 (N_8908,N_7600,N_7288);
and U8909 (N_8909,N_7750,N_7348);
or U8910 (N_8910,N_7617,N_7847);
nor U8911 (N_8911,N_6389,N_7037);
nor U8912 (N_8912,N_6048,N_6254);
nor U8913 (N_8913,N_7447,N_7030);
xnor U8914 (N_8914,N_7038,N_7064);
nor U8915 (N_8915,N_7034,N_7043);
and U8916 (N_8916,N_6429,N_6793);
or U8917 (N_8917,N_6131,N_6160);
nand U8918 (N_8918,N_6876,N_6374);
and U8919 (N_8919,N_7898,N_6128);
nand U8920 (N_8920,N_7599,N_6044);
nand U8921 (N_8921,N_7925,N_6092);
nand U8922 (N_8922,N_7264,N_6453);
or U8923 (N_8923,N_7475,N_7719);
nor U8924 (N_8924,N_7109,N_7152);
and U8925 (N_8925,N_6115,N_6457);
or U8926 (N_8926,N_7112,N_6771);
nor U8927 (N_8927,N_6380,N_6021);
or U8928 (N_8928,N_6898,N_7232);
xor U8929 (N_8929,N_6269,N_7595);
or U8930 (N_8930,N_7141,N_7387);
xnor U8931 (N_8931,N_6581,N_6797);
or U8932 (N_8932,N_7489,N_7145);
or U8933 (N_8933,N_7761,N_7912);
and U8934 (N_8934,N_6657,N_7252);
nand U8935 (N_8935,N_6878,N_7863);
nor U8936 (N_8936,N_7755,N_6551);
xnor U8937 (N_8937,N_7124,N_6625);
and U8938 (N_8938,N_6310,N_6468);
or U8939 (N_8939,N_6821,N_7215);
and U8940 (N_8940,N_7858,N_6872);
xor U8941 (N_8941,N_6193,N_6331);
nand U8942 (N_8942,N_6669,N_7032);
and U8943 (N_8943,N_6981,N_7808);
nor U8944 (N_8944,N_7728,N_6711);
xnor U8945 (N_8945,N_6734,N_6296);
nand U8946 (N_8946,N_7544,N_6111);
nand U8947 (N_8947,N_6094,N_7451);
xnor U8948 (N_8948,N_7522,N_6423);
or U8949 (N_8949,N_7492,N_6040);
xnor U8950 (N_8950,N_7105,N_7017);
or U8951 (N_8951,N_6724,N_6829);
nand U8952 (N_8952,N_6364,N_7616);
xnor U8953 (N_8953,N_7154,N_7465);
and U8954 (N_8954,N_7839,N_7803);
xor U8955 (N_8955,N_6151,N_7636);
xor U8956 (N_8956,N_6977,N_7067);
or U8957 (N_8957,N_7722,N_7829);
nor U8958 (N_8958,N_7740,N_6190);
nor U8959 (N_8959,N_7435,N_6943);
xnor U8960 (N_8960,N_7988,N_6595);
and U8961 (N_8961,N_6445,N_7261);
nand U8962 (N_8962,N_7274,N_6314);
xor U8963 (N_8963,N_7845,N_6306);
nor U8964 (N_8964,N_7771,N_7411);
nor U8965 (N_8965,N_6671,N_6060);
nor U8966 (N_8966,N_7204,N_7120);
nand U8967 (N_8967,N_7438,N_6264);
or U8968 (N_8968,N_7058,N_7896);
xnor U8969 (N_8969,N_7494,N_6345);
nand U8970 (N_8970,N_7637,N_7967);
or U8971 (N_8971,N_6142,N_7093);
nor U8972 (N_8972,N_7574,N_7688);
or U8973 (N_8973,N_6343,N_7278);
nand U8974 (N_8974,N_6377,N_6338);
and U8975 (N_8975,N_6944,N_6692);
and U8976 (N_8976,N_7123,N_6317);
xor U8977 (N_8977,N_6101,N_6777);
and U8978 (N_8978,N_6152,N_7008);
nand U8979 (N_8979,N_6914,N_6767);
nor U8980 (N_8980,N_7660,N_6855);
or U8981 (N_8981,N_6621,N_6623);
nor U8982 (N_8982,N_7455,N_6225);
and U8983 (N_8983,N_7749,N_7681);
and U8984 (N_8984,N_6169,N_7976);
or U8985 (N_8985,N_6347,N_7664);
nand U8986 (N_8986,N_7929,N_7604);
or U8987 (N_8987,N_6973,N_7804);
and U8988 (N_8988,N_7162,N_7011);
nor U8989 (N_8989,N_7315,N_6785);
nor U8990 (N_8990,N_6014,N_6099);
and U8991 (N_8991,N_7026,N_6593);
xnor U8992 (N_8992,N_7325,N_7871);
nand U8993 (N_8993,N_6662,N_6552);
or U8994 (N_8994,N_6297,N_7391);
and U8995 (N_8995,N_6786,N_7421);
and U8996 (N_8996,N_7830,N_6768);
nand U8997 (N_8997,N_6303,N_6425);
nor U8998 (N_8998,N_7209,N_6109);
nor U8999 (N_8999,N_6756,N_6912);
and U9000 (N_9000,N_7496,N_6386);
xnor U9001 (N_9001,N_7928,N_6534);
nor U9002 (N_9002,N_7788,N_7976);
xor U9003 (N_9003,N_7663,N_6723);
xnor U9004 (N_9004,N_6256,N_7368);
xor U9005 (N_9005,N_7021,N_7347);
nor U9006 (N_9006,N_6486,N_7934);
xnor U9007 (N_9007,N_7491,N_7537);
and U9008 (N_9008,N_6244,N_6953);
nand U9009 (N_9009,N_7004,N_7648);
nor U9010 (N_9010,N_7650,N_6559);
nand U9011 (N_9011,N_6322,N_6297);
or U9012 (N_9012,N_6991,N_6911);
nand U9013 (N_9013,N_7814,N_7935);
nor U9014 (N_9014,N_6555,N_7104);
xnor U9015 (N_9015,N_6971,N_7632);
nor U9016 (N_9016,N_6608,N_6146);
or U9017 (N_9017,N_6825,N_7647);
and U9018 (N_9018,N_6463,N_7284);
or U9019 (N_9019,N_7812,N_7368);
nand U9020 (N_9020,N_7921,N_6381);
xnor U9021 (N_9021,N_7784,N_7455);
xnor U9022 (N_9022,N_7162,N_6910);
xor U9023 (N_9023,N_7804,N_7222);
and U9024 (N_9024,N_7181,N_6696);
nor U9025 (N_9025,N_6885,N_7863);
nor U9026 (N_9026,N_6638,N_7552);
and U9027 (N_9027,N_7092,N_6665);
nand U9028 (N_9028,N_7162,N_6501);
nor U9029 (N_9029,N_6919,N_6298);
or U9030 (N_9030,N_7937,N_6229);
nor U9031 (N_9031,N_6046,N_7517);
xor U9032 (N_9032,N_6729,N_6201);
nor U9033 (N_9033,N_6992,N_7324);
or U9034 (N_9034,N_7994,N_7040);
or U9035 (N_9035,N_6789,N_7734);
xnor U9036 (N_9036,N_7339,N_7970);
nand U9037 (N_9037,N_6347,N_6925);
nand U9038 (N_9038,N_6972,N_7206);
nor U9039 (N_9039,N_7044,N_7147);
nand U9040 (N_9040,N_6910,N_6221);
xor U9041 (N_9041,N_7630,N_7040);
or U9042 (N_9042,N_7900,N_6439);
xnor U9043 (N_9043,N_6736,N_7980);
and U9044 (N_9044,N_6119,N_7689);
nor U9045 (N_9045,N_6898,N_6816);
and U9046 (N_9046,N_6623,N_7883);
or U9047 (N_9047,N_6468,N_7883);
and U9048 (N_9048,N_6028,N_7338);
xor U9049 (N_9049,N_6679,N_7164);
nor U9050 (N_9050,N_6187,N_6817);
xnor U9051 (N_9051,N_6709,N_7937);
and U9052 (N_9052,N_6533,N_6735);
nand U9053 (N_9053,N_7875,N_7029);
xnor U9054 (N_9054,N_7035,N_6479);
nand U9055 (N_9055,N_7061,N_7517);
xnor U9056 (N_9056,N_6808,N_7516);
nand U9057 (N_9057,N_6399,N_7556);
or U9058 (N_9058,N_7670,N_6246);
and U9059 (N_9059,N_6272,N_6822);
nand U9060 (N_9060,N_7050,N_7755);
and U9061 (N_9061,N_7923,N_6519);
and U9062 (N_9062,N_7257,N_6283);
and U9063 (N_9063,N_6313,N_7260);
and U9064 (N_9064,N_7752,N_6223);
nor U9065 (N_9065,N_6081,N_6466);
or U9066 (N_9066,N_6553,N_7403);
xor U9067 (N_9067,N_7836,N_6660);
nor U9068 (N_9068,N_6212,N_6654);
or U9069 (N_9069,N_6982,N_7333);
and U9070 (N_9070,N_7538,N_6469);
nor U9071 (N_9071,N_6061,N_7411);
nand U9072 (N_9072,N_6072,N_7192);
nand U9073 (N_9073,N_6880,N_6978);
xor U9074 (N_9074,N_7901,N_6768);
nand U9075 (N_9075,N_6603,N_7417);
or U9076 (N_9076,N_6624,N_6773);
xnor U9077 (N_9077,N_6015,N_6046);
xnor U9078 (N_9078,N_7698,N_7100);
nor U9079 (N_9079,N_6912,N_6353);
and U9080 (N_9080,N_6039,N_6687);
nor U9081 (N_9081,N_7009,N_6287);
and U9082 (N_9082,N_6087,N_6697);
nor U9083 (N_9083,N_6805,N_6438);
xnor U9084 (N_9084,N_7525,N_7346);
nor U9085 (N_9085,N_7572,N_7306);
and U9086 (N_9086,N_7317,N_7421);
nand U9087 (N_9087,N_6110,N_6720);
nand U9088 (N_9088,N_7481,N_6529);
nand U9089 (N_9089,N_7970,N_7953);
and U9090 (N_9090,N_6337,N_7158);
xnor U9091 (N_9091,N_6976,N_6486);
or U9092 (N_9092,N_6946,N_7856);
and U9093 (N_9093,N_6647,N_7850);
nor U9094 (N_9094,N_6259,N_6606);
and U9095 (N_9095,N_7500,N_7662);
nor U9096 (N_9096,N_6581,N_7320);
and U9097 (N_9097,N_7774,N_7976);
nand U9098 (N_9098,N_6323,N_7547);
and U9099 (N_9099,N_7002,N_6793);
or U9100 (N_9100,N_6884,N_6246);
xnor U9101 (N_9101,N_7891,N_7572);
nand U9102 (N_9102,N_7392,N_6981);
xor U9103 (N_9103,N_6734,N_6938);
nor U9104 (N_9104,N_7962,N_6101);
and U9105 (N_9105,N_6132,N_7069);
and U9106 (N_9106,N_6547,N_7385);
and U9107 (N_9107,N_7167,N_7077);
nand U9108 (N_9108,N_7680,N_7138);
and U9109 (N_9109,N_7366,N_6596);
nand U9110 (N_9110,N_7129,N_6805);
nand U9111 (N_9111,N_7643,N_6731);
and U9112 (N_9112,N_7509,N_6906);
nand U9113 (N_9113,N_6625,N_7444);
xor U9114 (N_9114,N_6962,N_7939);
xnor U9115 (N_9115,N_6623,N_6156);
xnor U9116 (N_9116,N_6950,N_7082);
and U9117 (N_9117,N_6938,N_6194);
nand U9118 (N_9118,N_6586,N_6502);
and U9119 (N_9119,N_7108,N_6565);
nand U9120 (N_9120,N_6411,N_6192);
nand U9121 (N_9121,N_6709,N_6338);
nor U9122 (N_9122,N_7359,N_6361);
xor U9123 (N_9123,N_6797,N_6266);
nand U9124 (N_9124,N_7765,N_6497);
and U9125 (N_9125,N_7354,N_7223);
xor U9126 (N_9126,N_7256,N_7555);
or U9127 (N_9127,N_7764,N_7368);
nand U9128 (N_9128,N_6794,N_6057);
xnor U9129 (N_9129,N_7577,N_7418);
nand U9130 (N_9130,N_7173,N_6237);
nor U9131 (N_9131,N_7336,N_7373);
xor U9132 (N_9132,N_7537,N_6215);
nor U9133 (N_9133,N_6205,N_6152);
and U9134 (N_9134,N_6500,N_6226);
nand U9135 (N_9135,N_7782,N_7949);
and U9136 (N_9136,N_7038,N_6576);
xnor U9137 (N_9137,N_6701,N_7826);
xor U9138 (N_9138,N_6658,N_6064);
or U9139 (N_9139,N_6700,N_7534);
nand U9140 (N_9140,N_6397,N_7125);
or U9141 (N_9141,N_7907,N_6599);
nor U9142 (N_9142,N_6777,N_6668);
and U9143 (N_9143,N_6523,N_6432);
or U9144 (N_9144,N_6308,N_7191);
nand U9145 (N_9145,N_6584,N_7370);
or U9146 (N_9146,N_6731,N_6140);
and U9147 (N_9147,N_6822,N_7586);
nor U9148 (N_9148,N_7199,N_6119);
and U9149 (N_9149,N_6720,N_6103);
nor U9150 (N_9150,N_7908,N_7191);
nand U9151 (N_9151,N_7253,N_6493);
xor U9152 (N_9152,N_6263,N_6991);
and U9153 (N_9153,N_7620,N_7196);
nand U9154 (N_9154,N_6534,N_7901);
or U9155 (N_9155,N_7445,N_7134);
xor U9156 (N_9156,N_6347,N_7596);
xor U9157 (N_9157,N_7056,N_6422);
nor U9158 (N_9158,N_7700,N_7567);
xor U9159 (N_9159,N_7510,N_6748);
or U9160 (N_9160,N_6645,N_6435);
and U9161 (N_9161,N_6098,N_6875);
nor U9162 (N_9162,N_6377,N_7025);
or U9163 (N_9163,N_7297,N_7335);
nor U9164 (N_9164,N_7163,N_7736);
nor U9165 (N_9165,N_7700,N_7698);
and U9166 (N_9166,N_6781,N_6075);
and U9167 (N_9167,N_7817,N_7161);
nor U9168 (N_9168,N_6886,N_7141);
and U9169 (N_9169,N_7485,N_6385);
or U9170 (N_9170,N_7451,N_7167);
nand U9171 (N_9171,N_6831,N_7302);
nor U9172 (N_9172,N_7566,N_6283);
and U9173 (N_9173,N_6011,N_6851);
nand U9174 (N_9174,N_7520,N_7332);
and U9175 (N_9175,N_7235,N_6766);
nor U9176 (N_9176,N_7498,N_7196);
nand U9177 (N_9177,N_6362,N_6683);
or U9178 (N_9178,N_7821,N_6416);
xor U9179 (N_9179,N_6572,N_6968);
nor U9180 (N_9180,N_6527,N_6703);
nand U9181 (N_9181,N_6796,N_6223);
nand U9182 (N_9182,N_7296,N_7484);
xnor U9183 (N_9183,N_6568,N_6470);
or U9184 (N_9184,N_6618,N_6194);
or U9185 (N_9185,N_6952,N_7073);
xnor U9186 (N_9186,N_6597,N_7118);
xor U9187 (N_9187,N_7701,N_7710);
nor U9188 (N_9188,N_6182,N_6456);
nand U9189 (N_9189,N_7245,N_7186);
or U9190 (N_9190,N_7832,N_6815);
nor U9191 (N_9191,N_7106,N_7656);
nand U9192 (N_9192,N_6921,N_6838);
xnor U9193 (N_9193,N_6529,N_7610);
nor U9194 (N_9194,N_6743,N_6285);
xor U9195 (N_9195,N_7429,N_6432);
or U9196 (N_9196,N_7084,N_7880);
and U9197 (N_9197,N_7676,N_7922);
nor U9198 (N_9198,N_7435,N_6986);
nand U9199 (N_9199,N_7303,N_6881);
xor U9200 (N_9200,N_7709,N_7792);
nand U9201 (N_9201,N_6004,N_7691);
nand U9202 (N_9202,N_7740,N_6311);
xnor U9203 (N_9203,N_6533,N_6319);
or U9204 (N_9204,N_6824,N_7698);
nor U9205 (N_9205,N_6729,N_6664);
nand U9206 (N_9206,N_6565,N_6905);
or U9207 (N_9207,N_7791,N_6144);
or U9208 (N_9208,N_6467,N_7416);
and U9209 (N_9209,N_6479,N_6414);
nand U9210 (N_9210,N_7361,N_7811);
nand U9211 (N_9211,N_6241,N_7981);
and U9212 (N_9212,N_7245,N_6644);
or U9213 (N_9213,N_7776,N_7916);
nor U9214 (N_9214,N_6932,N_6518);
xor U9215 (N_9215,N_6903,N_7168);
xnor U9216 (N_9216,N_7455,N_7605);
and U9217 (N_9217,N_7063,N_7819);
nor U9218 (N_9218,N_7505,N_7672);
nand U9219 (N_9219,N_7836,N_6302);
nand U9220 (N_9220,N_7884,N_6759);
nand U9221 (N_9221,N_6045,N_6165);
and U9222 (N_9222,N_6725,N_7121);
nand U9223 (N_9223,N_6297,N_6722);
nand U9224 (N_9224,N_6849,N_7278);
xor U9225 (N_9225,N_6631,N_7388);
nor U9226 (N_9226,N_6414,N_6268);
or U9227 (N_9227,N_6786,N_6394);
or U9228 (N_9228,N_6700,N_6351);
xor U9229 (N_9229,N_7205,N_7891);
and U9230 (N_9230,N_7945,N_6986);
and U9231 (N_9231,N_6445,N_6101);
xnor U9232 (N_9232,N_6107,N_7620);
and U9233 (N_9233,N_6911,N_6214);
xor U9234 (N_9234,N_6110,N_7984);
or U9235 (N_9235,N_6870,N_7537);
and U9236 (N_9236,N_6001,N_7307);
nand U9237 (N_9237,N_6730,N_7415);
and U9238 (N_9238,N_7964,N_6614);
nand U9239 (N_9239,N_6947,N_7333);
nor U9240 (N_9240,N_7577,N_6907);
or U9241 (N_9241,N_7511,N_6849);
or U9242 (N_9242,N_6326,N_6459);
xnor U9243 (N_9243,N_7034,N_6358);
or U9244 (N_9244,N_6076,N_7079);
and U9245 (N_9245,N_6903,N_7050);
or U9246 (N_9246,N_6261,N_6678);
nand U9247 (N_9247,N_7447,N_7444);
nand U9248 (N_9248,N_6595,N_7715);
or U9249 (N_9249,N_7757,N_6807);
or U9250 (N_9250,N_6466,N_6427);
nor U9251 (N_9251,N_6251,N_6986);
and U9252 (N_9252,N_7336,N_7388);
and U9253 (N_9253,N_6386,N_7116);
or U9254 (N_9254,N_7502,N_7675);
or U9255 (N_9255,N_7245,N_7683);
or U9256 (N_9256,N_6831,N_7814);
nand U9257 (N_9257,N_7318,N_7322);
nor U9258 (N_9258,N_6345,N_7463);
nor U9259 (N_9259,N_6934,N_6955);
xnor U9260 (N_9260,N_7239,N_6778);
nand U9261 (N_9261,N_7070,N_7547);
xor U9262 (N_9262,N_6379,N_6502);
and U9263 (N_9263,N_7488,N_6753);
and U9264 (N_9264,N_6756,N_7769);
or U9265 (N_9265,N_7989,N_6451);
nand U9266 (N_9266,N_7532,N_7394);
nand U9267 (N_9267,N_7967,N_7047);
or U9268 (N_9268,N_6629,N_7671);
nand U9269 (N_9269,N_7970,N_7563);
nand U9270 (N_9270,N_6668,N_7031);
and U9271 (N_9271,N_6934,N_6018);
nand U9272 (N_9272,N_6043,N_6961);
or U9273 (N_9273,N_6014,N_6495);
xor U9274 (N_9274,N_6345,N_6993);
xor U9275 (N_9275,N_6903,N_7186);
xor U9276 (N_9276,N_6384,N_7944);
nor U9277 (N_9277,N_6920,N_7165);
and U9278 (N_9278,N_7559,N_6083);
and U9279 (N_9279,N_6646,N_7915);
or U9280 (N_9280,N_6172,N_7935);
or U9281 (N_9281,N_6588,N_6377);
nand U9282 (N_9282,N_7381,N_7871);
nor U9283 (N_9283,N_6869,N_7457);
nand U9284 (N_9284,N_6065,N_6033);
nand U9285 (N_9285,N_7468,N_6561);
nor U9286 (N_9286,N_7866,N_6584);
nand U9287 (N_9287,N_7824,N_6874);
nand U9288 (N_9288,N_7589,N_6696);
nor U9289 (N_9289,N_6951,N_6752);
nor U9290 (N_9290,N_6750,N_7464);
nand U9291 (N_9291,N_6787,N_6957);
nor U9292 (N_9292,N_7180,N_7542);
xor U9293 (N_9293,N_7856,N_6007);
and U9294 (N_9294,N_7630,N_7974);
and U9295 (N_9295,N_7061,N_7206);
nand U9296 (N_9296,N_7445,N_7573);
nor U9297 (N_9297,N_6975,N_6176);
nor U9298 (N_9298,N_6032,N_7840);
or U9299 (N_9299,N_6543,N_7799);
nor U9300 (N_9300,N_7046,N_7697);
xor U9301 (N_9301,N_6930,N_7562);
and U9302 (N_9302,N_6379,N_6215);
or U9303 (N_9303,N_7219,N_6515);
nand U9304 (N_9304,N_6689,N_6662);
xor U9305 (N_9305,N_6907,N_6989);
nand U9306 (N_9306,N_7000,N_7457);
nor U9307 (N_9307,N_7228,N_7778);
nand U9308 (N_9308,N_7530,N_7744);
xnor U9309 (N_9309,N_6228,N_6234);
xnor U9310 (N_9310,N_6572,N_7019);
nand U9311 (N_9311,N_7458,N_7173);
nand U9312 (N_9312,N_6890,N_7824);
nand U9313 (N_9313,N_7054,N_7810);
xnor U9314 (N_9314,N_6727,N_7655);
xnor U9315 (N_9315,N_6263,N_7957);
xor U9316 (N_9316,N_7465,N_6563);
nand U9317 (N_9317,N_7019,N_7434);
xor U9318 (N_9318,N_7533,N_7410);
xor U9319 (N_9319,N_7741,N_7161);
and U9320 (N_9320,N_7732,N_6925);
nand U9321 (N_9321,N_7652,N_7694);
nand U9322 (N_9322,N_7136,N_6739);
xor U9323 (N_9323,N_6641,N_6258);
or U9324 (N_9324,N_7969,N_6062);
nand U9325 (N_9325,N_7033,N_7482);
or U9326 (N_9326,N_6528,N_7176);
xnor U9327 (N_9327,N_7938,N_6127);
or U9328 (N_9328,N_6454,N_7122);
or U9329 (N_9329,N_6300,N_7475);
or U9330 (N_9330,N_6186,N_7262);
nor U9331 (N_9331,N_7730,N_6780);
and U9332 (N_9332,N_7791,N_7201);
nor U9333 (N_9333,N_7720,N_7142);
nor U9334 (N_9334,N_6556,N_6337);
xnor U9335 (N_9335,N_7352,N_7966);
nand U9336 (N_9336,N_6714,N_7630);
and U9337 (N_9337,N_7664,N_7039);
and U9338 (N_9338,N_6624,N_6780);
nor U9339 (N_9339,N_7281,N_6185);
nand U9340 (N_9340,N_6300,N_7744);
or U9341 (N_9341,N_6687,N_7430);
nand U9342 (N_9342,N_6638,N_6168);
xor U9343 (N_9343,N_6300,N_7278);
and U9344 (N_9344,N_7756,N_6076);
nand U9345 (N_9345,N_6338,N_7046);
and U9346 (N_9346,N_6597,N_6553);
nand U9347 (N_9347,N_7431,N_6738);
and U9348 (N_9348,N_6087,N_7973);
nor U9349 (N_9349,N_6021,N_7870);
nor U9350 (N_9350,N_7206,N_7253);
or U9351 (N_9351,N_6054,N_6037);
or U9352 (N_9352,N_6318,N_7401);
and U9353 (N_9353,N_6950,N_7234);
and U9354 (N_9354,N_7429,N_6705);
nor U9355 (N_9355,N_7014,N_7331);
and U9356 (N_9356,N_6106,N_7231);
or U9357 (N_9357,N_7410,N_7972);
and U9358 (N_9358,N_7318,N_7197);
xnor U9359 (N_9359,N_6525,N_6488);
or U9360 (N_9360,N_6383,N_6489);
nand U9361 (N_9361,N_6585,N_7939);
or U9362 (N_9362,N_6582,N_6329);
nor U9363 (N_9363,N_7275,N_6525);
or U9364 (N_9364,N_6605,N_6220);
nand U9365 (N_9365,N_7011,N_6164);
and U9366 (N_9366,N_7061,N_7253);
or U9367 (N_9367,N_6829,N_6963);
or U9368 (N_9368,N_7604,N_7092);
and U9369 (N_9369,N_6808,N_6087);
nand U9370 (N_9370,N_6761,N_7716);
nor U9371 (N_9371,N_6317,N_7781);
nand U9372 (N_9372,N_6855,N_7910);
nand U9373 (N_9373,N_6214,N_6489);
nand U9374 (N_9374,N_6053,N_7790);
nor U9375 (N_9375,N_7925,N_6916);
and U9376 (N_9376,N_7442,N_7612);
nand U9377 (N_9377,N_7268,N_7028);
xor U9378 (N_9378,N_7829,N_7685);
and U9379 (N_9379,N_7557,N_7388);
or U9380 (N_9380,N_7120,N_7824);
nand U9381 (N_9381,N_6029,N_6531);
nor U9382 (N_9382,N_6809,N_6202);
or U9383 (N_9383,N_6360,N_7157);
xnor U9384 (N_9384,N_6642,N_6021);
nand U9385 (N_9385,N_7693,N_7257);
and U9386 (N_9386,N_6817,N_7183);
nand U9387 (N_9387,N_6313,N_7881);
nor U9388 (N_9388,N_7953,N_7565);
nand U9389 (N_9389,N_7372,N_6796);
nand U9390 (N_9390,N_7701,N_7303);
or U9391 (N_9391,N_6979,N_7277);
and U9392 (N_9392,N_6072,N_6098);
and U9393 (N_9393,N_7163,N_6130);
xnor U9394 (N_9394,N_6529,N_6327);
and U9395 (N_9395,N_7748,N_6614);
or U9396 (N_9396,N_7415,N_6418);
and U9397 (N_9397,N_7622,N_7032);
and U9398 (N_9398,N_6186,N_6136);
and U9399 (N_9399,N_6413,N_7662);
or U9400 (N_9400,N_6238,N_7542);
or U9401 (N_9401,N_7844,N_6275);
and U9402 (N_9402,N_6475,N_7554);
and U9403 (N_9403,N_7763,N_7203);
and U9404 (N_9404,N_6458,N_7463);
xnor U9405 (N_9405,N_7999,N_7527);
xnor U9406 (N_9406,N_6850,N_6199);
or U9407 (N_9407,N_6065,N_6036);
and U9408 (N_9408,N_6381,N_7514);
or U9409 (N_9409,N_7353,N_6789);
xnor U9410 (N_9410,N_7630,N_7936);
or U9411 (N_9411,N_6419,N_6294);
xnor U9412 (N_9412,N_7631,N_6529);
nand U9413 (N_9413,N_7580,N_6545);
nand U9414 (N_9414,N_6135,N_7139);
and U9415 (N_9415,N_6400,N_6753);
and U9416 (N_9416,N_6711,N_6100);
and U9417 (N_9417,N_6428,N_6533);
nand U9418 (N_9418,N_6832,N_7458);
nor U9419 (N_9419,N_7605,N_6697);
nor U9420 (N_9420,N_7219,N_7514);
or U9421 (N_9421,N_6989,N_7401);
or U9422 (N_9422,N_6278,N_7560);
or U9423 (N_9423,N_6152,N_7755);
xnor U9424 (N_9424,N_6457,N_7065);
nand U9425 (N_9425,N_6977,N_7517);
or U9426 (N_9426,N_7799,N_7240);
and U9427 (N_9427,N_6654,N_7577);
or U9428 (N_9428,N_6002,N_6976);
xnor U9429 (N_9429,N_6791,N_6632);
nand U9430 (N_9430,N_7951,N_7381);
nor U9431 (N_9431,N_6204,N_6937);
nor U9432 (N_9432,N_7688,N_7554);
and U9433 (N_9433,N_6787,N_7736);
and U9434 (N_9434,N_7595,N_7550);
xnor U9435 (N_9435,N_7409,N_6704);
nand U9436 (N_9436,N_7720,N_6534);
xnor U9437 (N_9437,N_6263,N_6244);
nor U9438 (N_9438,N_7919,N_6645);
xor U9439 (N_9439,N_6691,N_7926);
and U9440 (N_9440,N_7366,N_7825);
or U9441 (N_9441,N_7913,N_6011);
nand U9442 (N_9442,N_7228,N_7499);
and U9443 (N_9443,N_7814,N_6057);
xnor U9444 (N_9444,N_7837,N_7858);
xor U9445 (N_9445,N_7251,N_7418);
nand U9446 (N_9446,N_7784,N_6357);
nand U9447 (N_9447,N_7149,N_7942);
or U9448 (N_9448,N_7493,N_6079);
or U9449 (N_9449,N_6142,N_7927);
nor U9450 (N_9450,N_7332,N_7595);
xnor U9451 (N_9451,N_6588,N_7489);
or U9452 (N_9452,N_7636,N_7124);
nor U9453 (N_9453,N_6388,N_6613);
and U9454 (N_9454,N_7082,N_7912);
and U9455 (N_9455,N_6144,N_6811);
or U9456 (N_9456,N_7687,N_6840);
and U9457 (N_9457,N_7924,N_6174);
and U9458 (N_9458,N_6726,N_7248);
xor U9459 (N_9459,N_7513,N_7305);
and U9460 (N_9460,N_6939,N_6869);
xor U9461 (N_9461,N_7427,N_6849);
nand U9462 (N_9462,N_6612,N_6704);
nand U9463 (N_9463,N_6766,N_7747);
nand U9464 (N_9464,N_7945,N_7497);
nand U9465 (N_9465,N_6468,N_7022);
nor U9466 (N_9466,N_7067,N_6802);
and U9467 (N_9467,N_6661,N_7372);
and U9468 (N_9468,N_7135,N_6902);
or U9469 (N_9469,N_6791,N_7926);
nand U9470 (N_9470,N_6040,N_6100);
xor U9471 (N_9471,N_6565,N_7749);
and U9472 (N_9472,N_7171,N_7049);
nor U9473 (N_9473,N_6542,N_6171);
and U9474 (N_9474,N_6718,N_6273);
nor U9475 (N_9475,N_7845,N_6401);
and U9476 (N_9476,N_6364,N_7867);
nor U9477 (N_9477,N_6831,N_7321);
nor U9478 (N_9478,N_7972,N_6068);
or U9479 (N_9479,N_6497,N_7553);
nand U9480 (N_9480,N_7346,N_6250);
nand U9481 (N_9481,N_7044,N_6169);
and U9482 (N_9482,N_7380,N_7767);
and U9483 (N_9483,N_6128,N_6217);
or U9484 (N_9484,N_7605,N_7688);
nand U9485 (N_9485,N_6487,N_6337);
nand U9486 (N_9486,N_6438,N_6953);
nand U9487 (N_9487,N_6542,N_7227);
nor U9488 (N_9488,N_7516,N_6453);
xor U9489 (N_9489,N_6067,N_7005);
and U9490 (N_9490,N_7322,N_7712);
or U9491 (N_9491,N_6558,N_7696);
nor U9492 (N_9492,N_6454,N_6389);
or U9493 (N_9493,N_6431,N_7596);
nor U9494 (N_9494,N_6198,N_6032);
and U9495 (N_9495,N_6911,N_6901);
xor U9496 (N_9496,N_6939,N_7563);
nor U9497 (N_9497,N_7546,N_6321);
or U9498 (N_9498,N_6578,N_6042);
nand U9499 (N_9499,N_6472,N_7887);
xor U9500 (N_9500,N_7699,N_6475);
xnor U9501 (N_9501,N_7025,N_6863);
nor U9502 (N_9502,N_7376,N_6189);
nand U9503 (N_9503,N_7071,N_7266);
and U9504 (N_9504,N_6593,N_7511);
and U9505 (N_9505,N_6473,N_7006);
nand U9506 (N_9506,N_7429,N_6180);
nor U9507 (N_9507,N_7560,N_6434);
nand U9508 (N_9508,N_7457,N_7528);
nor U9509 (N_9509,N_7807,N_7494);
and U9510 (N_9510,N_7053,N_7013);
nand U9511 (N_9511,N_6290,N_6164);
xnor U9512 (N_9512,N_6193,N_6440);
or U9513 (N_9513,N_6266,N_7038);
and U9514 (N_9514,N_7049,N_6190);
nand U9515 (N_9515,N_6902,N_6495);
and U9516 (N_9516,N_6673,N_6297);
xor U9517 (N_9517,N_6065,N_6713);
or U9518 (N_9518,N_6055,N_7714);
xor U9519 (N_9519,N_6500,N_6025);
nor U9520 (N_9520,N_6387,N_7300);
nand U9521 (N_9521,N_6076,N_7193);
or U9522 (N_9522,N_6792,N_7236);
and U9523 (N_9523,N_7255,N_6269);
xnor U9524 (N_9524,N_7419,N_6686);
or U9525 (N_9525,N_6575,N_6055);
nand U9526 (N_9526,N_7219,N_6154);
or U9527 (N_9527,N_7925,N_6594);
nand U9528 (N_9528,N_7802,N_7898);
or U9529 (N_9529,N_6794,N_7693);
xor U9530 (N_9530,N_6276,N_7849);
or U9531 (N_9531,N_6907,N_6761);
or U9532 (N_9532,N_6104,N_6466);
xor U9533 (N_9533,N_6784,N_6966);
nand U9534 (N_9534,N_6087,N_7805);
or U9535 (N_9535,N_7924,N_6523);
and U9536 (N_9536,N_7920,N_6859);
or U9537 (N_9537,N_6538,N_6950);
nand U9538 (N_9538,N_7179,N_7301);
nand U9539 (N_9539,N_6979,N_7837);
or U9540 (N_9540,N_6528,N_6913);
xnor U9541 (N_9541,N_7898,N_6124);
nor U9542 (N_9542,N_6159,N_6072);
xnor U9543 (N_9543,N_6679,N_6677);
nand U9544 (N_9544,N_7795,N_7058);
or U9545 (N_9545,N_7310,N_7894);
or U9546 (N_9546,N_6014,N_6714);
and U9547 (N_9547,N_6381,N_7064);
and U9548 (N_9548,N_6540,N_6977);
or U9549 (N_9549,N_6789,N_6179);
or U9550 (N_9550,N_6209,N_7510);
and U9551 (N_9551,N_6686,N_6632);
and U9552 (N_9552,N_7762,N_7006);
or U9553 (N_9553,N_7136,N_7912);
and U9554 (N_9554,N_6116,N_7055);
xor U9555 (N_9555,N_6507,N_7492);
xor U9556 (N_9556,N_6919,N_7262);
xnor U9557 (N_9557,N_6573,N_6460);
or U9558 (N_9558,N_6200,N_6881);
and U9559 (N_9559,N_7572,N_7971);
xnor U9560 (N_9560,N_6161,N_7693);
nand U9561 (N_9561,N_6284,N_6168);
and U9562 (N_9562,N_7430,N_7978);
and U9563 (N_9563,N_7764,N_7531);
nor U9564 (N_9564,N_7857,N_7647);
and U9565 (N_9565,N_7189,N_7445);
and U9566 (N_9566,N_7989,N_6292);
nor U9567 (N_9567,N_6746,N_6139);
nor U9568 (N_9568,N_6941,N_7294);
nand U9569 (N_9569,N_7333,N_7138);
or U9570 (N_9570,N_6548,N_7325);
nor U9571 (N_9571,N_7942,N_6996);
nand U9572 (N_9572,N_7372,N_6716);
or U9573 (N_9573,N_6278,N_7350);
nor U9574 (N_9574,N_6114,N_7875);
or U9575 (N_9575,N_6045,N_6460);
xor U9576 (N_9576,N_7591,N_6502);
nand U9577 (N_9577,N_6932,N_6394);
or U9578 (N_9578,N_6495,N_7873);
or U9579 (N_9579,N_6968,N_7754);
and U9580 (N_9580,N_6119,N_6459);
nor U9581 (N_9581,N_7482,N_7239);
nand U9582 (N_9582,N_7529,N_7290);
or U9583 (N_9583,N_6330,N_7951);
nand U9584 (N_9584,N_6512,N_6753);
nor U9585 (N_9585,N_7602,N_6484);
xor U9586 (N_9586,N_6983,N_6482);
xor U9587 (N_9587,N_7982,N_7058);
and U9588 (N_9588,N_7948,N_7805);
nand U9589 (N_9589,N_7717,N_6746);
nor U9590 (N_9590,N_6738,N_6683);
and U9591 (N_9591,N_6366,N_6734);
nor U9592 (N_9592,N_6340,N_6730);
xor U9593 (N_9593,N_6467,N_6044);
nand U9594 (N_9594,N_6797,N_6828);
and U9595 (N_9595,N_7500,N_6572);
nand U9596 (N_9596,N_6620,N_6053);
nor U9597 (N_9597,N_6799,N_7363);
and U9598 (N_9598,N_7233,N_6613);
nor U9599 (N_9599,N_6709,N_7103);
and U9600 (N_9600,N_7456,N_7397);
or U9601 (N_9601,N_6914,N_6385);
nand U9602 (N_9602,N_7651,N_7136);
or U9603 (N_9603,N_6666,N_6968);
xnor U9604 (N_9604,N_6427,N_7804);
or U9605 (N_9605,N_6290,N_6444);
xnor U9606 (N_9606,N_6867,N_7234);
or U9607 (N_9607,N_7286,N_6073);
nand U9608 (N_9608,N_7790,N_6120);
xnor U9609 (N_9609,N_6525,N_7964);
nand U9610 (N_9610,N_6214,N_6017);
and U9611 (N_9611,N_7196,N_7069);
xor U9612 (N_9612,N_7517,N_7659);
or U9613 (N_9613,N_6684,N_7767);
nand U9614 (N_9614,N_6347,N_7883);
xnor U9615 (N_9615,N_7171,N_6718);
nand U9616 (N_9616,N_6098,N_7273);
and U9617 (N_9617,N_6379,N_6748);
nor U9618 (N_9618,N_6069,N_7776);
or U9619 (N_9619,N_6044,N_7685);
nand U9620 (N_9620,N_6349,N_6930);
or U9621 (N_9621,N_7582,N_7707);
nor U9622 (N_9622,N_7876,N_6561);
nand U9623 (N_9623,N_7925,N_7722);
or U9624 (N_9624,N_6020,N_6938);
and U9625 (N_9625,N_7612,N_7105);
nand U9626 (N_9626,N_6534,N_6018);
nand U9627 (N_9627,N_6346,N_7161);
nor U9628 (N_9628,N_7003,N_6820);
nand U9629 (N_9629,N_7157,N_6458);
or U9630 (N_9630,N_6286,N_6976);
xor U9631 (N_9631,N_7056,N_6195);
xnor U9632 (N_9632,N_7551,N_7393);
or U9633 (N_9633,N_6027,N_7892);
nand U9634 (N_9634,N_6859,N_7857);
and U9635 (N_9635,N_6791,N_7601);
and U9636 (N_9636,N_6683,N_7907);
xor U9637 (N_9637,N_7312,N_6431);
or U9638 (N_9638,N_6727,N_6102);
and U9639 (N_9639,N_7381,N_6457);
and U9640 (N_9640,N_6285,N_6711);
nand U9641 (N_9641,N_6658,N_6222);
xnor U9642 (N_9642,N_6618,N_7577);
nor U9643 (N_9643,N_7955,N_6475);
nand U9644 (N_9644,N_6614,N_7617);
nand U9645 (N_9645,N_7363,N_7680);
nor U9646 (N_9646,N_7681,N_7888);
or U9647 (N_9647,N_7434,N_7218);
nor U9648 (N_9648,N_6486,N_6169);
and U9649 (N_9649,N_7024,N_7130);
nand U9650 (N_9650,N_7948,N_7568);
nor U9651 (N_9651,N_6507,N_7727);
xnor U9652 (N_9652,N_6055,N_6221);
nand U9653 (N_9653,N_7175,N_6732);
and U9654 (N_9654,N_7669,N_7558);
nand U9655 (N_9655,N_7137,N_6501);
and U9656 (N_9656,N_7184,N_7533);
or U9657 (N_9657,N_7437,N_7931);
or U9658 (N_9658,N_7621,N_7667);
or U9659 (N_9659,N_7942,N_7006);
nand U9660 (N_9660,N_6033,N_6566);
or U9661 (N_9661,N_7861,N_6953);
or U9662 (N_9662,N_7847,N_6315);
xor U9663 (N_9663,N_7213,N_6915);
or U9664 (N_9664,N_6688,N_7780);
nor U9665 (N_9665,N_6596,N_6300);
and U9666 (N_9666,N_6728,N_6971);
or U9667 (N_9667,N_7347,N_7041);
or U9668 (N_9668,N_7436,N_6732);
xor U9669 (N_9669,N_7813,N_6825);
nor U9670 (N_9670,N_6409,N_7361);
and U9671 (N_9671,N_6563,N_7868);
or U9672 (N_9672,N_6986,N_7538);
nor U9673 (N_9673,N_7203,N_7849);
or U9674 (N_9674,N_6694,N_7481);
xor U9675 (N_9675,N_6252,N_7829);
xor U9676 (N_9676,N_7918,N_6346);
and U9677 (N_9677,N_6802,N_7469);
xnor U9678 (N_9678,N_6134,N_7122);
nand U9679 (N_9679,N_7689,N_6476);
nand U9680 (N_9680,N_6081,N_6492);
and U9681 (N_9681,N_6897,N_7540);
and U9682 (N_9682,N_6338,N_7705);
nor U9683 (N_9683,N_6256,N_7006);
nor U9684 (N_9684,N_7292,N_6288);
nand U9685 (N_9685,N_7596,N_7235);
and U9686 (N_9686,N_7187,N_7676);
or U9687 (N_9687,N_6171,N_7551);
or U9688 (N_9688,N_7237,N_7266);
nor U9689 (N_9689,N_6403,N_6927);
and U9690 (N_9690,N_6461,N_6128);
nand U9691 (N_9691,N_6408,N_6588);
nor U9692 (N_9692,N_7769,N_6257);
and U9693 (N_9693,N_7185,N_7235);
or U9694 (N_9694,N_7332,N_6807);
nand U9695 (N_9695,N_7193,N_7908);
and U9696 (N_9696,N_6143,N_7754);
xor U9697 (N_9697,N_6517,N_6891);
or U9698 (N_9698,N_7335,N_7041);
nor U9699 (N_9699,N_6473,N_6973);
or U9700 (N_9700,N_6915,N_6578);
nand U9701 (N_9701,N_7318,N_6949);
nor U9702 (N_9702,N_7972,N_7865);
nand U9703 (N_9703,N_6836,N_6792);
xnor U9704 (N_9704,N_7651,N_7520);
and U9705 (N_9705,N_7983,N_7318);
or U9706 (N_9706,N_6358,N_6272);
nand U9707 (N_9707,N_7966,N_7384);
or U9708 (N_9708,N_7418,N_6040);
nand U9709 (N_9709,N_7497,N_6375);
and U9710 (N_9710,N_6977,N_6994);
or U9711 (N_9711,N_6596,N_6162);
nand U9712 (N_9712,N_6627,N_6105);
or U9713 (N_9713,N_6593,N_6180);
nand U9714 (N_9714,N_7028,N_6737);
nor U9715 (N_9715,N_7967,N_7652);
nand U9716 (N_9716,N_7536,N_7786);
nor U9717 (N_9717,N_7011,N_6417);
and U9718 (N_9718,N_6693,N_6391);
nor U9719 (N_9719,N_7233,N_7582);
nand U9720 (N_9720,N_7373,N_7537);
nor U9721 (N_9721,N_7330,N_6541);
or U9722 (N_9722,N_7464,N_7978);
or U9723 (N_9723,N_7049,N_7227);
nand U9724 (N_9724,N_6274,N_7632);
or U9725 (N_9725,N_7298,N_6561);
and U9726 (N_9726,N_7691,N_6429);
nor U9727 (N_9727,N_7861,N_6907);
nor U9728 (N_9728,N_6630,N_7961);
xnor U9729 (N_9729,N_7014,N_7038);
nand U9730 (N_9730,N_6101,N_6593);
nand U9731 (N_9731,N_6172,N_7593);
nor U9732 (N_9732,N_6657,N_7682);
or U9733 (N_9733,N_6944,N_7945);
xnor U9734 (N_9734,N_7264,N_7028);
or U9735 (N_9735,N_7414,N_7282);
or U9736 (N_9736,N_7288,N_6649);
or U9737 (N_9737,N_6363,N_7064);
or U9738 (N_9738,N_7394,N_7185);
or U9739 (N_9739,N_6917,N_7038);
xor U9740 (N_9740,N_6992,N_7080);
nor U9741 (N_9741,N_6498,N_6145);
nor U9742 (N_9742,N_7400,N_6440);
xnor U9743 (N_9743,N_7590,N_7994);
xor U9744 (N_9744,N_6513,N_7550);
or U9745 (N_9745,N_7883,N_6481);
or U9746 (N_9746,N_7947,N_6621);
xor U9747 (N_9747,N_6015,N_6494);
xnor U9748 (N_9748,N_6170,N_6174);
xnor U9749 (N_9749,N_6072,N_6707);
or U9750 (N_9750,N_6107,N_7938);
nor U9751 (N_9751,N_7559,N_7462);
nor U9752 (N_9752,N_7748,N_6043);
or U9753 (N_9753,N_7293,N_6216);
and U9754 (N_9754,N_7784,N_7934);
or U9755 (N_9755,N_6604,N_6110);
nor U9756 (N_9756,N_6549,N_6893);
nand U9757 (N_9757,N_6349,N_6520);
xnor U9758 (N_9758,N_7817,N_6589);
or U9759 (N_9759,N_6117,N_7993);
nand U9760 (N_9760,N_7548,N_7001);
xnor U9761 (N_9761,N_7602,N_6658);
nand U9762 (N_9762,N_6270,N_7599);
or U9763 (N_9763,N_6340,N_7822);
nor U9764 (N_9764,N_6880,N_7727);
nor U9765 (N_9765,N_6664,N_6848);
and U9766 (N_9766,N_7271,N_6505);
nor U9767 (N_9767,N_6996,N_6780);
xnor U9768 (N_9768,N_6702,N_7606);
xnor U9769 (N_9769,N_6262,N_7298);
xor U9770 (N_9770,N_6561,N_7279);
or U9771 (N_9771,N_6342,N_6987);
nor U9772 (N_9772,N_6437,N_6086);
and U9773 (N_9773,N_6348,N_7992);
or U9774 (N_9774,N_6917,N_7150);
or U9775 (N_9775,N_7652,N_7565);
nand U9776 (N_9776,N_7895,N_7161);
or U9777 (N_9777,N_6746,N_7233);
nor U9778 (N_9778,N_6877,N_7857);
nand U9779 (N_9779,N_7516,N_6756);
or U9780 (N_9780,N_7234,N_6953);
xnor U9781 (N_9781,N_6470,N_6410);
or U9782 (N_9782,N_7456,N_6021);
nand U9783 (N_9783,N_6760,N_6055);
or U9784 (N_9784,N_6320,N_6294);
and U9785 (N_9785,N_7741,N_7142);
xnor U9786 (N_9786,N_6584,N_6258);
nor U9787 (N_9787,N_7274,N_6395);
nand U9788 (N_9788,N_7966,N_7493);
and U9789 (N_9789,N_7754,N_7743);
nand U9790 (N_9790,N_6803,N_7036);
or U9791 (N_9791,N_6928,N_6173);
xnor U9792 (N_9792,N_7990,N_7580);
or U9793 (N_9793,N_6309,N_6267);
and U9794 (N_9794,N_6526,N_7185);
nand U9795 (N_9795,N_6944,N_6021);
or U9796 (N_9796,N_6911,N_6330);
and U9797 (N_9797,N_7155,N_6997);
or U9798 (N_9798,N_6864,N_6446);
or U9799 (N_9799,N_6455,N_7642);
nor U9800 (N_9800,N_7308,N_6968);
or U9801 (N_9801,N_6352,N_6914);
nand U9802 (N_9802,N_7347,N_6288);
nor U9803 (N_9803,N_7999,N_6342);
nand U9804 (N_9804,N_6475,N_6752);
nor U9805 (N_9805,N_7934,N_6976);
nand U9806 (N_9806,N_6972,N_6010);
nand U9807 (N_9807,N_7941,N_7215);
nand U9808 (N_9808,N_7629,N_7760);
nand U9809 (N_9809,N_7396,N_6383);
nor U9810 (N_9810,N_6023,N_7090);
xnor U9811 (N_9811,N_7345,N_7813);
nor U9812 (N_9812,N_7181,N_6291);
and U9813 (N_9813,N_6114,N_6135);
or U9814 (N_9814,N_7515,N_7255);
and U9815 (N_9815,N_7308,N_6534);
xor U9816 (N_9816,N_6548,N_6784);
nor U9817 (N_9817,N_7448,N_7136);
xnor U9818 (N_9818,N_7011,N_6124);
nand U9819 (N_9819,N_7356,N_6171);
or U9820 (N_9820,N_7771,N_6170);
or U9821 (N_9821,N_6255,N_7151);
or U9822 (N_9822,N_7359,N_6812);
and U9823 (N_9823,N_6468,N_7331);
and U9824 (N_9824,N_6035,N_7517);
xnor U9825 (N_9825,N_6252,N_6113);
nor U9826 (N_9826,N_7521,N_7279);
and U9827 (N_9827,N_7406,N_6259);
or U9828 (N_9828,N_7461,N_6675);
xor U9829 (N_9829,N_7726,N_6833);
or U9830 (N_9830,N_6025,N_6071);
xnor U9831 (N_9831,N_7456,N_7105);
nor U9832 (N_9832,N_7397,N_7787);
nand U9833 (N_9833,N_7082,N_7077);
nor U9834 (N_9834,N_6047,N_7433);
and U9835 (N_9835,N_6426,N_6854);
xnor U9836 (N_9836,N_6242,N_6911);
xnor U9837 (N_9837,N_6455,N_6393);
nor U9838 (N_9838,N_7073,N_6770);
xnor U9839 (N_9839,N_7838,N_6840);
and U9840 (N_9840,N_7780,N_6655);
xor U9841 (N_9841,N_6333,N_6472);
nor U9842 (N_9842,N_7644,N_7135);
xor U9843 (N_9843,N_6381,N_7196);
nor U9844 (N_9844,N_6606,N_7009);
nand U9845 (N_9845,N_6222,N_7776);
or U9846 (N_9846,N_6528,N_6236);
nand U9847 (N_9847,N_7631,N_6232);
xor U9848 (N_9848,N_7953,N_6881);
or U9849 (N_9849,N_7689,N_7794);
or U9850 (N_9850,N_6497,N_7038);
xnor U9851 (N_9851,N_6284,N_7974);
nor U9852 (N_9852,N_7194,N_7143);
nand U9853 (N_9853,N_7361,N_7637);
nor U9854 (N_9854,N_6693,N_6652);
or U9855 (N_9855,N_6129,N_7291);
and U9856 (N_9856,N_6970,N_7225);
or U9857 (N_9857,N_7538,N_6630);
or U9858 (N_9858,N_6996,N_6111);
nor U9859 (N_9859,N_6589,N_7242);
xor U9860 (N_9860,N_6037,N_6686);
or U9861 (N_9861,N_6827,N_6327);
or U9862 (N_9862,N_6104,N_7959);
or U9863 (N_9863,N_6522,N_6563);
nor U9864 (N_9864,N_6885,N_6126);
or U9865 (N_9865,N_6437,N_6999);
nor U9866 (N_9866,N_7796,N_7356);
nand U9867 (N_9867,N_6805,N_7618);
nand U9868 (N_9868,N_6944,N_7135);
nor U9869 (N_9869,N_7076,N_7552);
xnor U9870 (N_9870,N_6643,N_6087);
nand U9871 (N_9871,N_7543,N_6740);
xor U9872 (N_9872,N_7320,N_6894);
xnor U9873 (N_9873,N_6310,N_7655);
xor U9874 (N_9874,N_7190,N_7614);
nand U9875 (N_9875,N_6580,N_7819);
or U9876 (N_9876,N_6846,N_6775);
nor U9877 (N_9877,N_6572,N_7885);
and U9878 (N_9878,N_6364,N_6969);
xnor U9879 (N_9879,N_6421,N_7274);
nor U9880 (N_9880,N_6689,N_7145);
xnor U9881 (N_9881,N_7189,N_6623);
or U9882 (N_9882,N_6292,N_6082);
or U9883 (N_9883,N_6031,N_7078);
nand U9884 (N_9884,N_7704,N_7182);
or U9885 (N_9885,N_7509,N_6582);
nor U9886 (N_9886,N_7201,N_7764);
xor U9887 (N_9887,N_7230,N_7722);
or U9888 (N_9888,N_7548,N_7287);
and U9889 (N_9889,N_7482,N_6580);
nor U9890 (N_9890,N_6355,N_7376);
nor U9891 (N_9891,N_6438,N_6407);
xor U9892 (N_9892,N_6479,N_7086);
nand U9893 (N_9893,N_6477,N_7966);
nand U9894 (N_9894,N_7079,N_7511);
xor U9895 (N_9895,N_6379,N_7814);
nand U9896 (N_9896,N_6319,N_7992);
nand U9897 (N_9897,N_6820,N_7631);
xnor U9898 (N_9898,N_7521,N_7511);
nand U9899 (N_9899,N_7989,N_6345);
or U9900 (N_9900,N_6369,N_7015);
and U9901 (N_9901,N_6431,N_6301);
or U9902 (N_9902,N_7040,N_6152);
nand U9903 (N_9903,N_6173,N_6183);
xnor U9904 (N_9904,N_6485,N_7762);
nand U9905 (N_9905,N_6752,N_7259);
xor U9906 (N_9906,N_6639,N_6491);
nor U9907 (N_9907,N_6402,N_7458);
nand U9908 (N_9908,N_6127,N_7841);
nor U9909 (N_9909,N_7062,N_7132);
and U9910 (N_9910,N_6831,N_6350);
nand U9911 (N_9911,N_6969,N_7300);
xnor U9912 (N_9912,N_7408,N_7977);
and U9913 (N_9913,N_6371,N_7984);
or U9914 (N_9914,N_7301,N_6789);
or U9915 (N_9915,N_6958,N_6984);
or U9916 (N_9916,N_6661,N_7985);
or U9917 (N_9917,N_7147,N_7872);
xor U9918 (N_9918,N_6466,N_6051);
nor U9919 (N_9919,N_7862,N_7614);
nor U9920 (N_9920,N_6890,N_6266);
or U9921 (N_9921,N_6728,N_7061);
nor U9922 (N_9922,N_6820,N_6434);
or U9923 (N_9923,N_7652,N_6773);
xor U9924 (N_9924,N_6977,N_6698);
or U9925 (N_9925,N_7968,N_6518);
nand U9926 (N_9926,N_7700,N_7169);
or U9927 (N_9927,N_6243,N_7742);
nor U9928 (N_9928,N_7277,N_7534);
nand U9929 (N_9929,N_7169,N_7879);
nand U9930 (N_9930,N_6813,N_7433);
nand U9931 (N_9931,N_6833,N_6099);
xor U9932 (N_9932,N_7872,N_6378);
and U9933 (N_9933,N_6479,N_6492);
xor U9934 (N_9934,N_7357,N_7995);
nand U9935 (N_9935,N_6314,N_6734);
nor U9936 (N_9936,N_6587,N_6284);
and U9937 (N_9937,N_6939,N_7401);
nand U9938 (N_9938,N_7361,N_6502);
nand U9939 (N_9939,N_6919,N_6121);
and U9940 (N_9940,N_7087,N_7123);
or U9941 (N_9941,N_6111,N_7919);
nand U9942 (N_9942,N_7146,N_7628);
nand U9943 (N_9943,N_7683,N_6177);
nand U9944 (N_9944,N_6933,N_6756);
nand U9945 (N_9945,N_7252,N_6524);
xnor U9946 (N_9946,N_6647,N_7865);
and U9947 (N_9947,N_6045,N_7190);
xnor U9948 (N_9948,N_7312,N_7119);
and U9949 (N_9949,N_7224,N_7745);
nor U9950 (N_9950,N_7068,N_6829);
xnor U9951 (N_9951,N_7294,N_7296);
nand U9952 (N_9952,N_7303,N_7529);
nor U9953 (N_9953,N_7256,N_7487);
nand U9954 (N_9954,N_7624,N_6183);
or U9955 (N_9955,N_6993,N_6360);
and U9956 (N_9956,N_7158,N_6363);
nor U9957 (N_9957,N_7830,N_7959);
or U9958 (N_9958,N_7464,N_6993);
nor U9959 (N_9959,N_7005,N_7515);
or U9960 (N_9960,N_7191,N_6338);
nand U9961 (N_9961,N_6774,N_6068);
xor U9962 (N_9962,N_6197,N_7172);
and U9963 (N_9963,N_7031,N_7699);
xor U9964 (N_9964,N_7008,N_6544);
and U9965 (N_9965,N_7794,N_6187);
or U9966 (N_9966,N_7778,N_6720);
nand U9967 (N_9967,N_6493,N_6898);
or U9968 (N_9968,N_6428,N_7869);
xnor U9969 (N_9969,N_7206,N_7382);
xor U9970 (N_9970,N_7338,N_7984);
and U9971 (N_9971,N_7809,N_7819);
nand U9972 (N_9972,N_7925,N_7668);
and U9973 (N_9973,N_6728,N_7668);
xnor U9974 (N_9974,N_7643,N_6744);
xnor U9975 (N_9975,N_7458,N_6926);
or U9976 (N_9976,N_6607,N_6299);
and U9977 (N_9977,N_6254,N_6187);
nor U9978 (N_9978,N_6037,N_7442);
and U9979 (N_9979,N_7420,N_6488);
or U9980 (N_9980,N_7904,N_7363);
or U9981 (N_9981,N_7654,N_7595);
xor U9982 (N_9982,N_7041,N_7428);
or U9983 (N_9983,N_6512,N_6676);
and U9984 (N_9984,N_6938,N_7338);
or U9985 (N_9985,N_7793,N_6048);
nor U9986 (N_9986,N_6677,N_6778);
xnor U9987 (N_9987,N_7046,N_7992);
nand U9988 (N_9988,N_6121,N_6637);
or U9989 (N_9989,N_6777,N_7363);
and U9990 (N_9990,N_7067,N_7357);
and U9991 (N_9991,N_6551,N_7057);
nor U9992 (N_9992,N_7404,N_7079);
xor U9993 (N_9993,N_7466,N_6109);
xor U9994 (N_9994,N_6711,N_6477);
nand U9995 (N_9995,N_6644,N_6528);
and U9996 (N_9996,N_6024,N_6979);
and U9997 (N_9997,N_6371,N_6561);
xnor U9998 (N_9998,N_6683,N_7882);
nand U9999 (N_9999,N_7083,N_6167);
xnor UO_0 (O_0,N_9044,N_9813);
or UO_1 (O_1,N_9099,N_8169);
nand UO_2 (O_2,N_9041,N_8899);
nand UO_3 (O_3,N_8655,N_8506);
nor UO_4 (O_4,N_8880,N_8119);
nor UO_5 (O_5,N_8473,N_9994);
nor UO_6 (O_6,N_8626,N_8988);
nand UO_7 (O_7,N_8415,N_8080);
xnor UO_8 (O_8,N_8448,N_9562);
or UO_9 (O_9,N_9823,N_8563);
or UO_10 (O_10,N_9262,N_8553);
nand UO_11 (O_11,N_9997,N_9481);
or UO_12 (O_12,N_9820,N_9977);
nand UO_13 (O_13,N_9479,N_8271);
xor UO_14 (O_14,N_9443,N_9129);
and UO_15 (O_15,N_9606,N_8973);
nor UO_16 (O_16,N_8363,N_8590);
nor UO_17 (O_17,N_9593,N_8310);
and UO_18 (O_18,N_9970,N_9101);
and UO_19 (O_19,N_9386,N_9419);
or UO_20 (O_20,N_9538,N_8199);
xnor UO_21 (O_21,N_9374,N_8830);
nand UO_22 (O_22,N_9080,N_9581);
or UO_23 (O_23,N_9328,N_8218);
nand UO_24 (O_24,N_8738,N_8766);
and UO_25 (O_25,N_8995,N_9445);
xor UO_26 (O_26,N_9746,N_8859);
or UO_27 (O_27,N_9310,N_8051);
or UO_28 (O_28,N_8798,N_8581);
or UO_29 (O_29,N_9449,N_9156);
nand UO_30 (O_30,N_9227,N_8166);
nor UO_31 (O_31,N_9621,N_8542);
and UO_32 (O_32,N_9467,N_9781);
nor UO_33 (O_33,N_9671,N_9319);
nor UO_34 (O_34,N_9709,N_8290);
nor UO_35 (O_35,N_9003,N_9791);
or UO_36 (O_36,N_9808,N_9806);
xor UO_37 (O_37,N_9002,N_8243);
nand UO_38 (O_38,N_8047,N_9726);
nand UO_39 (O_39,N_8374,N_9821);
or UO_40 (O_40,N_9687,N_9889);
nand UO_41 (O_41,N_8433,N_8191);
nand UO_42 (O_42,N_8979,N_8055);
xor UO_43 (O_43,N_9368,N_9351);
nand UO_44 (O_44,N_9852,N_8726);
nor UO_45 (O_45,N_9789,N_9498);
nor UO_46 (O_46,N_9412,N_8855);
nand UO_47 (O_47,N_9814,N_9798);
or UO_48 (O_48,N_9656,N_9858);
nor UO_49 (O_49,N_8355,N_8361);
xor UO_50 (O_50,N_9552,N_9846);
or UO_51 (O_51,N_8193,N_9308);
nor UO_52 (O_52,N_8320,N_9250);
and UO_53 (O_53,N_8638,N_8325);
nor UO_54 (O_54,N_8931,N_9468);
and UO_55 (O_55,N_9465,N_8593);
xnor UO_56 (O_56,N_8485,N_9578);
nand UO_57 (O_57,N_9038,N_8665);
or UO_58 (O_58,N_8965,N_8058);
nor UO_59 (O_59,N_8424,N_8216);
nand UO_60 (O_60,N_8226,N_9140);
and UO_61 (O_61,N_9408,N_9117);
and UO_62 (O_62,N_9064,N_8804);
and UO_63 (O_63,N_8969,N_8627);
xor UO_64 (O_64,N_8913,N_8941);
nor UO_65 (O_65,N_8690,N_8545);
and UO_66 (O_66,N_9513,N_9034);
or UO_67 (O_67,N_9484,N_8881);
and UO_68 (O_68,N_9131,N_8440);
nor UO_69 (O_69,N_8050,N_9097);
nand UO_70 (O_70,N_9017,N_9841);
or UO_71 (O_71,N_9198,N_8641);
nand UO_72 (O_72,N_9608,N_8777);
and UO_73 (O_73,N_9924,N_8173);
nor UO_74 (O_74,N_9204,N_9116);
nor UO_75 (O_75,N_9990,N_8745);
nand UO_76 (O_76,N_8444,N_9396);
or UO_77 (O_77,N_9486,N_8113);
xor UO_78 (O_78,N_8518,N_8032);
xor UO_79 (O_79,N_9167,N_8044);
xnor UO_80 (O_80,N_9657,N_8073);
xnor UO_81 (O_81,N_8114,N_9127);
or UO_82 (O_82,N_8452,N_9021);
and UO_83 (O_83,N_9298,N_8062);
or UO_84 (O_84,N_9502,N_9752);
nand UO_85 (O_85,N_8522,N_8749);
nor UO_86 (O_86,N_8295,N_9570);
and UO_87 (O_87,N_8213,N_9891);
nand UO_88 (O_88,N_9734,N_8399);
nor UO_89 (O_89,N_8413,N_8364);
or UO_90 (O_90,N_8237,N_8223);
xor UO_91 (O_91,N_9141,N_8352);
or UO_92 (O_92,N_8708,N_8577);
or UO_93 (O_93,N_9278,N_9337);
or UO_94 (O_94,N_9978,N_9497);
xor UO_95 (O_95,N_8875,N_8315);
or UO_96 (O_96,N_9886,N_9345);
nand UO_97 (O_97,N_9910,N_9272);
nand UO_98 (O_98,N_9215,N_8842);
or UO_99 (O_99,N_9059,N_8664);
nand UO_100 (O_100,N_8688,N_9106);
or UO_101 (O_101,N_9398,N_9880);
nand UO_102 (O_102,N_8680,N_9218);
and UO_103 (O_103,N_9194,N_9875);
or UO_104 (O_104,N_9955,N_8771);
and UO_105 (O_105,N_9762,N_9695);
and UO_106 (O_106,N_9890,N_8395);
nor UO_107 (O_107,N_9348,N_8342);
and UO_108 (O_108,N_9874,N_8697);
or UO_109 (O_109,N_8538,N_8873);
nor UO_110 (O_110,N_8872,N_9030);
xnor UO_111 (O_111,N_9123,N_9669);
nor UO_112 (O_112,N_9799,N_9268);
and UO_113 (O_113,N_8387,N_9810);
and UO_114 (O_114,N_9933,N_8784);
and UO_115 (O_115,N_9023,N_8095);
and UO_116 (O_116,N_9591,N_8858);
nor UO_117 (O_117,N_9359,N_8728);
or UO_118 (O_118,N_9190,N_8084);
or UO_119 (O_119,N_8061,N_9115);
or UO_120 (O_120,N_8662,N_8565);
or UO_121 (O_121,N_8279,N_9893);
nand UO_122 (O_122,N_8029,N_8006);
or UO_123 (O_123,N_9622,N_8645);
nand UO_124 (O_124,N_9232,N_8052);
nor UO_125 (O_125,N_9401,N_8706);
nand UO_126 (O_126,N_8103,N_9338);
and UO_127 (O_127,N_8510,N_8887);
and UO_128 (O_128,N_8249,N_9639);
or UO_129 (O_129,N_9664,N_9714);
nand UO_130 (O_130,N_9316,N_8098);
nor UO_131 (O_131,N_8512,N_9940);
nand UO_132 (O_132,N_8228,N_8631);
and UO_133 (O_133,N_9912,N_9847);
xnor UO_134 (O_134,N_9378,N_9981);
or UO_135 (O_135,N_9046,N_8280);
or UO_136 (O_136,N_8498,N_9773);
or UO_137 (O_137,N_9558,N_9674);
or UO_138 (O_138,N_9514,N_8704);
and UO_139 (O_139,N_8617,N_8238);
nand UO_140 (O_140,N_8319,N_8871);
nand UO_141 (O_141,N_9224,N_8588);
nand UO_142 (O_142,N_9913,N_9866);
nand UO_143 (O_143,N_8940,N_9837);
nand UO_144 (O_144,N_8524,N_8480);
and UO_145 (O_145,N_8849,N_9540);
nor UO_146 (O_146,N_9922,N_9584);
nor UO_147 (O_147,N_9731,N_8847);
and UO_148 (O_148,N_8862,N_9435);
or UO_149 (O_149,N_9843,N_9026);
xnor UO_150 (O_150,N_8264,N_9377);
nor UO_151 (O_151,N_8710,N_9960);
or UO_152 (O_152,N_8539,N_9546);
or UO_153 (O_153,N_9666,N_9066);
and UO_154 (O_154,N_9031,N_9133);
nand UO_155 (O_155,N_9221,N_8456);
and UO_156 (O_156,N_8391,N_8041);
nand UO_157 (O_157,N_9462,N_9701);
nand UO_158 (O_158,N_9554,N_8230);
and UO_159 (O_159,N_9984,N_8414);
or UO_160 (O_160,N_8164,N_9915);
and UO_161 (O_161,N_8020,N_8381);
or UO_162 (O_162,N_9958,N_9261);
xnor UO_163 (O_163,N_9119,N_8576);
nor UO_164 (O_164,N_8247,N_8868);
nand UO_165 (O_165,N_9177,N_9085);
or UO_166 (O_166,N_8852,N_9640);
and UO_167 (O_167,N_9289,N_9599);
nor UO_168 (O_168,N_8551,N_9055);
or UO_169 (O_169,N_9077,N_8469);
xnor UO_170 (O_170,N_9052,N_9779);
nand UO_171 (O_171,N_9950,N_8145);
or UO_172 (O_172,N_8770,N_9304);
xnor UO_173 (O_173,N_9132,N_9534);
xor UO_174 (O_174,N_9020,N_8287);
or UO_175 (O_175,N_9597,N_9094);
nor UO_176 (O_176,N_8813,N_8289);
and UO_177 (O_177,N_8916,N_9483);
nand UO_178 (O_178,N_8422,N_9499);
and UO_179 (O_179,N_8718,N_8479);
or UO_180 (O_180,N_8435,N_9393);
or UO_181 (O_181,N_8179,N_8333);
nor UO_182 (O_182,N_8729,N_9312);
xor UO_183 (O_183,N_9456,N_8416);
or UO_184 (O_184,N_9057,N_8412);
and UO_185 (O_185,N_8393,N_8097);
nand UO_186 (O_186,N_8453,N_9469);
xnor UO_187 (O_187,N_9180,N_9580);
xnor UO_188 (O_188,N_8186,N_9192);
or UO_189 (O_189,N_8863,N_8520);
xnor UO_190 (O_190,N_9281,N_9983);
nor UO_191 (O_191,N_8116,N_8261);
nand UO_192 (O_192,N_8225,N_9440);
xor UO_193 (O_193,N_8040,N_8937);
xnor UO_194 (O_194,N_8754,N_8076);
and UO_195 (O_195,N_9182,N_9536);
nand UO_196 (O_196,N_9004,N_8764);
and UO_197 (O_197,N_9800,N_9371);
nand UO_198 (O_198,N_8094,N_8304);
xor UO_199 (O_199,N_9457,N_8953);
or UO_200 (O_200,N_8924,N_9925);
and UO_201 (O_201,N_9557,N_8550);
and UO_202 (O_202,N_9394,N_8282);
or UO_203 (O_203,N_8370,N_9501);
or UO_204 (O_204,N_9200,N_8669);
nand UO_205 (O_205,N_8011,N_9504);
or UO_206 (O_206,N_8671,N_8668);
xor UO_207 (O_207,N_8724,N_9700);
nand UO_208 (O_208,N_8244,N_9561);
nor UO_209 (O_209,N_8936,N_8908);
and UO_210 (O_210,N_8928,N_8944);
nor UO_211 (O_211,N_8752,N_8093);
nor UO_212 (O_212,N_8486,N_9815);
or UO_213 (O_213,N_9551,N_9128);
xnor UO_214 (O_214,N_9697,N_8144);
nor UO_215 (O_215,N_9191,N_8330);
nor UO_216 (O_216,N_8468,N_9474);
xor UO_217 (O_217,N_9860,N_9850);
nand UO_218 (O_218,N_9476,N_8968);
nand UO_219 (O_219,N_9176,N_9114);
nor UO_220 (O_220,N_9539,N_9964);
and UO_221 (O_221,N_9336,N_9838);
or UO_222 (O_222,N_8929,N_9676);
or UO_223 (O_223,N_8254,N_9299);
and UO_224 (O_224,N_9206,N_9317);
and UO_225 (O_225,N_8778,N_8188);
nand UO_226 (O_226,N_8568,N_9305);
xnor UO_227 (O_227,N_9906,N_9069);
and UO_228 (O_228,N_8975,N_9022);
or UO_229 (O_229,N_9965,N_9189);
xnor UO_230 (O_230,N_9638,N_8323);
xor UO_231 (O_231,N_9225,N_9226);
and UO_232 (O_232,N_9556,N_8702);
and UO_233 (O_233,N_8999,N_9845);
nand UO_234 (O_234,N_9724,N_8611);
or UO_235 (O_235,N_8720,N_8721);
and UO_236 (O_236,N_9411,N_9859);
xor UO_237 (O_237,N_9919,N_9945);
and UO_238 (O_238,N_9526,N_9384);
nand UO_239 (O_239,N_8850,N_8366);
xor UO_240 (O_240,N_9856,N_9938);
xor UO_241 (O_241,N_9611,N_8077);
nand UO_242 (O_242,N_9730,N_8744);
or UO_243 (O_243,N_9753,N_9690);
nand UO_244 (O_244,N_9529,N_8065);
or UO_245 (O_245,N_9001,N_8864);
nand UO_246 (O_246,N_9488,N_8552);
and UO_247 (O_247,N_9704,N_8151);
and UO_248 (O_248,N_9908,N_8499);
nor UO_249 (O_249,N_8652,N_8821);
and UO_250 (O_250,N_8501,N_9573);
and UO_251 (O_251,N_8088,N_8909);
or UO_252 (O_252,N_9610,N_9087);
nor UO_253 (O_253,N_8423,N_9618);
or UO_254 (O_254,N_8496,N_9683);
and UO_255 (O_255,N_9899,N_9260);
nand UO_256 (O_256,N_8786,N_8684);
nand UO_257 (O_257,N_9027,N_8483);
nand UO_258 (O_258,N_9314,N_8848);
and UO_259 (O_259,N_8439,N_9146);
xnor UO_260 (O_260,N_9433,N_8630);
nor UO_261 (O_261,N_8207,N_9187);
nand UO_262 (O_262,N_8102,N_8066);
or UO_263 (O_263,N_9313,N_9450);
nor UO_264 (O_264,N_9110,N_8951);
nor UO_265 (O_265,N_9461,N_9842);
and UO_266 (O_266,N_8385,N_9006);
xnor UO_267 (O_267,N_9492,N_9356);
xnor UO_268 (O_268,N_8014,N_8796);
and UO_269 (O_269,N_9632,N_9205);
nor UO_270 (O_270,N_8070,N_9968);
xnor UO_271 (O_271,N_9986,N_9409);
nor UO_272 (O_272,N_9559,N_8340);
or UO_273 (O_273,N_9160,N_8826);
nand UO_274 (O_274,N_9712,N_8344);
or UO_275 (O_275,N_8131,N_9809);
nand UO_276 (O_276,N_8240,N_9234);
and UO_277 (O_277,N_9475,N_9315);
xnor UO_278 (O_278,N_8886,N_8396);
nor UO_279 (O_279,N_8075,N_9757);
nand UO_280 (O_280,N_9869,N_8554);
xnor UO_281 (O_281,N_8201,N_9949);
and UO_282 (O_282,N_9222,N_8765);
nand UO_283 (O_283,N_8016,N_9231);
xnor UO_284 (O_284,N_9705,N_8128);
or UO_285 (O_285,N_9971,N_8607);
nor UO_286 (O_286,N_8168,N_9742);
nor UO_287 (O_287,N_9517,N_8907);
or UO_288 (O_288,N_9975,N_9532);
or UO_289 (O_289,N_8118,N_8298);
and UO_290 (O_290,N_9793,N_9873);
nor UO_291 (O_291,N_9954,N_8825);
nand UO_292 (O_292,N_9266,N_8782);
or UO_293 (O_293,N_8807,N_9060);
and UO_294 (O_294,N_8541,N_8241);
and UO_295 (O_295,N_8354,N_8252);
or UO_296 (O_296,N_8418,N_9086);
xor UO_297 (O_297,N_9024,N_8489);
and UO_298 (O_298,N_8682,N_8829);
nor UO_299 (O_299,N_8383,N_9832);
nor UO_300 (O_300,N_8935,N_9145);
and UO_301 (O_301,N_9427,N_8582);
nor UO_302 (O_302,N_9966,N_9203);
and UO_303 (O_303,N_9755,N_8629);
or UO_304 (O_304,N_9733,N_8599);
nor UO_305 (O_305,N_8827,N_8274);
and UO_306 (O_306,N_8775,N_8170);
nor UO_307 (O_307,N_8753,N_9211);
or UO_308 (O_308,N_8699,N_9416);
or UO_309 (O_309,N_9564,N_8734);
xnor UO_310 (O_310,N_9170,N_9091);
and UO_311 (O_311,N_8768,N_9230);
and UO_312 (O_312,N_8947,N_9329);
nor UO_313 (O_313,N_9238,N_8705);
nand UO_314 (O_314,N_8291,N_9589);
nand UO_315 (O_315,N_9171,N_9962);
nand UO_316 (O_316,N_9719,N_8962);
nor UO_317 (O_317,N_9068,N_9452);
nor UO_318 (O_318,N_8234,N_8063);
nor UO_319 (O_319,N_8272,N_8150);
nand UO_320 (O_320,N_8527,N_8269);
or UO_321 (O_321,N_9078,N_8059);
nand UO_322 (O_322,N_8376,N_8471);
nand UO_323 (O_323,N_9152,N_8187);
xor UO_324 (O_324,N_8981,N_8123);
nand UO_325 (O_325,N_9749,N_8991);
nand UO_326 (O_326,N_9207,N_8160);
nand UO_327 (O_327,N_9344,N_9372);
nand UO_328 (O_328,N_9598,N_8637);
xnor UO_329 (O_329,N_8785,N_8152);
nand UO_330 (O_330,N_8870,N_8488);
nand UO_331 (O_331,N_8893,N_9918);
and UO_332 (O_332,N_9349,N_8491);
and UO_333 (O_333,N_8009,N_8475);
xor UO_334 (O_334,N_8008,N_8819);
xnor UO_335 (O_335,N_9183,N_8747);
xor UO_336 (O_336,N_8996,N_8198);
nand UO_337 (O_337,N_8389,N_9121);
nor UO_338 (O_338,N_9202,N_8019);
nand UO_339 (O_339,N_8514,N_8096);
nand UO_340 (O_340,N_8197,N_8037);
xor UO_341 (O_341,N_9615,N_9721);
and UO_342 (O_342,N_8183,N_8108);
or UO_343 (O_343,N_8823,N_8679);
nor UO_344 (O_344,N_9596,N_9609);
nand UO_345 (O_345,N_8557,N_8712);
or UO_346 (O_346,N_8616,N_9375);
nand UO_347 (O_347,N_9273,N_9357);
or UO_348 (O_348,N_9645,N_9729);
nor UO_349 (O_349,N_8661,N_8492);
xor UO_350 (O_350,N_8606,N_8987);
or UO_351 (O_351,N_8772,N_8153);
nand UO_352 (O_352,N_9533,N_9587);
xor UO_353 (O_353,N_8540,N_8956);
and UO_354 (O_354,N_8203,N_9446);
nand UO_355 (O_355,N_9029,N_8619);
and UO_356 (O_356,N_9716,N_8544);
nand UO_357 (O_357,N_8656,N_8949);
nand UO_358 (O_358,N_9051,N_9453);
or UO_359 (O_359,N_8876,N_8334);
nor UO_360 (O_360,N_9223,N_8429);
and UO_361 (O_361,N_9049,N_8356);
nand UO_362 (O_362,N_8474,N_9784);
and UO_363 (O_363,N_9431,N_9074);
nand UO_364 (O_364,N_8214,N_8809);
xnor UO_365 (O_365,N_8653,N_8537);
and UO_366 (O_366,N_8614,N_9699);
or UO_367 (O_367,N_8647,N_8436);
or UO_368 (O_368,N_9139,N_9153);
nand UO_369 (O_369,N_8003,N_9169);
nor UO_370 (O_370,N_8185,N_9048);
nor UO_371 (O_371,N_8209,N_8329);
or UO_372 (O_372,N_8731,N_9459);
nand UO_373 (O_373,N_9485,N_8124);
or UO_374 (O_374,N_9667,N_9567);
or UO_375 (O_375,N_9290,N_9340);
nand UO_376 (O_376,N_8998,N_9917);
nor UO_377 (O_377,N_8017,N_9947);
xnor UO_378 (O_378,N_8392,N_8115);
nand UO_379 (O_379,N_9025,N_9415);
xor UO_380 (O_380,N_9787,N_8380);
nand UO_381 (O_381,N_8659,N_9967);
xor UO_382 (O_382,N_9770,N_9295);
nand UO_383 (O_383,N_9619,N_8285);
xor UO_384 (O_384,N_9296,N_8036);
xnor UO_385 (O_385,N_9015,N_8945);
and UO_386 (O_386,N_9948,N_9565);
nor UO_387 (O_387,N_9604,N_8622);
nand UO_388 (O_388,N_8977,N_8405);
nor UO_389 (O_389,N_9493,N_9330);
nand UO_390 (O_390,N_9905,N_8901);
or UO_391 (O_391,N_9658,N_9424);
xor UO_392 (O_392,N_9100,N_8331);
and UO_393 (O_393,N_8709,N_9527);
xor UO_394 (O_394,N_9627,N_8676);
and UO_395 (O_395,N_8950,N_8265);
or UO_396 (O_396,N_9804,N_8722);
nand UO_397 (O_397,N_9648,N_8211);
nor UO_398 (O_398,N_9681,N_8643);
or UO_399 (O_399,N_9659,N_9936);
and UO_400 (O_400,N_8918,N_9723);
or UO_401 (O_401,N_8171,N_8466);
or UO_402 (O_402,N_8589,N_8814);
nor UO_403 (O_403,N_9436,N_8028);
and UO_404 (O_404,N_9710,N_9840);
and UO_405 (O_405,N_9258,N_8297);
or UO_406 (O_406,N_8681,N_9271);
nand UO_407 (O_407,N_8314,N_8903);
nand UO_408 (O_408,N_9142,N_8038);
nand UO_409 (O_409,N_9072,N_9923);
nor UO_410 (O_410,N_8189,N_9545);
nor UO_411 (O_411,N_9014,N_9898);
xnor UO_412 (O_412,N_9745,N_9780);
xor UO_413 (O_413,N_9568,N_8365);
xor UO_414 (O_414,N_9686,N_8042);
or UO_415 (O_415,N_8739,N_9969);
and UO_416 (O_416,N_8674,N_8046);
nand UO_417 (O_417,N_9879,N_9229);
nand UO_418 (O_418,N_8800,N_8672);
nand UO_419 (O_419,N_8445,N_8367);
nand UO_420 (O_420,N_8902,N_8311);
xor UO_421 (O_421,N_9595,N_8454);
or UO_422 (O_422,N_9876,N_8140);
xnor UO_423 (O_423,N_9122,N_8202);
nand UO_424 (O_424,N_8253,N_8043);
nand UO_425 (O_425,N_8182,N_8157);
or UO_426 (O_426,N_9463,N_9601);
nor UO_427 (O_427,N_8683,N_8603);
nor UO_428 (O_428,N_9976,N_8426);
and UO_429 (O_429,N_9764,N_8368);
or UO_430 (O_430,N_9892,N_8215);
xnor UO_431 (O_431,N_8045,N_9061);
nor UO_432 (O_432,N_8451,N_9903);
nor UO_433 (O_433,N_8972,N_8428);
xor UO_434 (O_434,N_8815,N_8336);
nand UO_435 (O_435,N_9390,N_8034);
xnor UO_436 (O_436,N_8357,N_8284);
nor UO_437 (O_437,N_8258,N_9777);
or UO_438 (O_438,N_8733,N_8411);
nor UO_439 (O_439,N_9395,N_8547);
and UO_440 (O_440,N_9795,N_9172);
xnor UO_441 (O_441,N_8750,N_9016);
xor UO_442 (O_442,N_9071,N_8591);
xnor UO_443 (O_443,N_8419,N_9239);
or UO_444 (O_444,N_9149,N_9796);
nand UO_445 (O_445,N_9988,N_9735);
and UO_446 (O_446,N_8963,N_8696);
xor UO_447 (O_447,N_8343,N_8450);
xnor UO_448 (O_448,N_8634,N_8461);
xnor UO_449 (O_449,N_8455,N_9854);
nand UO_450 (O_450,N_8470,N_8580);
or UO_451 (O_451,N_9675,N_9366);
or UO_452 (O_452,N_9352,N_9201);
and UO_453 (O_453,N_8633,N_8923);
or UO_454 (O_454,N_8236,N_9163);
or UO_455 (O_455,N_8421,N_9033);
or UO_456 (O_456,N_9343,N_8528);
xor UO_457 (O_457,N_9603,N_9276);
or UO_458 (O_458,N_8494,N_9353);
or UO_459 (O_459,N_9042,N_9240);
xnor UO_460 (O_460,N_8231,N_9901);
xor UO_461 (O_461,N_9297,N_8472);
nor UO_462 (O_462,N_9228,N_8162);
and UO_463 (O_463,N_9439,N_8027);
and UO_464 (O_464,N_8586,N_8335);
or UO_465 (O_465,N_9358,N_8635);
or UO_466 (O_466,N_8976,N_8530);
or UO_467 (O_467,N_9897,N_8312);
nor UO_468 (O_468,N_8675,N_8110);
or UO_469 (O_469,N_8623,N_8099);
or UO_470 (O_470,N_9895,N_9523);
nor UO_471 (O_471,N_8313,N_8811);
and UO_472 (O_472,N_8256,N_9185);
nor UO_473 (O_473,N_8317,N_9644);
or UO_474 (O_474,N_9829,N_8639);
xnor UO_475 (O_475,N_9835,N_9429);
nand UO_476 (O_476,N_8158,N_9280);
nand UO_477 (O_477,N_8081,N_9065);
nor UO_478 (O_478,N_8837,N_9692);
and UO_479 (O_479,N_8229,N_8497);
or UO_480 (O_480,N_9095,N_9089);
and UO_481 (O_481,N_9614,N_8255);
or UO_482 (O_482,N_9819,N_9863);
or UO_483 (O_483,N_8914,N_8984);
nand UO_484 (O_484,N_9500,N_8477);
and UO_485 (O_485,N_8758,N_9706);
nand UO_486 (O_486,N_8134,N_8007);
and UO_487 (O_487,N_8262,N_8584);
nor UO_488 (O_488,N_9422,N_8163);
or UO_489 (O_489,N_9321,N_8505);
and UO_490 (O_490,N_8068,N_8318);
nand UO_491 (O_491,N_9935,N_9506);
nand UO_492 (O_492,N_9404,N_8447);
or UO_493 (O_493,N_9980,N_8693);
and UO_494 (O_494,N_9150,N_9574);
or UO_495 (O_495,N_8742,N_9548);
nand UO_496 (O_496,N_8670,N_9217);
nor UO_497 (O_497,N_8303,N_9489);
xnor UO_498 (O_498,N_9590,N_8574);
and UO_499 (O_499,N_8767,N_8172);
and UO_500 (O_500,N_8286,N_9264);
nand UO_501 (O_501,N_9711,N_8030);
nand UO_502 (O_502,N_9494,N_9547);
and UO_503 (O_503,N_9350,N_8649);
or UO_504 (O_504,N_9511,N_9790);
nand UO_505 (O_505,N_8787,N_9582);
xor UO_506 (O_506,N_9625,N_8579);
xor UO_507 (O_507,N_8082,N_8861);
or UO_508 (O_508,N_9047,N_9836);
nor UO_509 (O_509,N_9682,N_8024);
or UO_510 (O_510,N_8831,N_9037);
nand UO_511 (O_511,N_9322,N_8328);
nand UO_512 (O_512,N_9727,N_9294);
xnor UO_513 (O_513,N_8090,N_9113);
xor UO_514 (O_514,N_8462,N_8083);
nand UO_515 (O_515,N_8021,N_8657);
xor UO_516 (O_516,N_8056,N_9524);
nand UO_517 (O_517,N_8519,N_8865);
or UO_518 (O_518,N_9679,N_9549);
xor UO_519 (O_519,N_8667,N_8615);
xor UO_520 (O_520,N_9996,N_9515);
or UO_521 (O_521,N_9009,N_8857);
nand UO_522 (O_522,N_9293,N_8822);
xnor UO_523 (O_523,N_8717,N_9914);
and UO_524 (O_524,N_9728,N_9098);
and UO_525 (O_525,N_8911,N_8560);
or UO_526 (O_526,N_8122,N_8500);
xnor UO_527 (O_527,N_8281,N_9346);
xor UO_528 (O_528,N_9380,N_9165);
nor UO_529 (O_529,N_9179,N_8139);
nand UO_530 (O_530,N_9857,N_9339);
xnor UO_531 (O_531,N_9541,N_8339);
nor UO_532 (O_532,N_9233,N_9155);
or UO_533 (O_533,N_9216,N_9707);
nand UO_534 (O_534,N_8994,N_9235);
xor UO_535 (O_535,N_9011,N_8713);
nand UO_536 (O_536,N_8711,N_9364);
or UO_537 (O_537,N_8601,N_8898);
nor UO_538 (O_538,N_9812,N_9503);
and UO_539 (O_539,N_9956,N_8146);
or UO_540 (O_540,N_8434,N_9050);
xnor UO_541 (O_541,N_8790,N_8906);
xor UO_542 (O_542,N_9441,N_8362);
xor UO_543 (O_543,N_8874,N_8130);
nand UO_544 (O_544,N_8817,N_9542);
nor UO_545 (O_545,N_9320,N_9677);
or UO_546 (O_546,N_8879,N_9008);
nor UO_547 (O_547,N_8493,N_9107);
and UO_548 (O_548,N_8602,N_9387);
or UO_549 (O_549,N_9403,N_9028);
or UO_550 (O_550,N_9553,N_8853);
nand UO_551 (O_551,N_9932,N_9126);
and UO_552 (O_552,N_9473,N_8910);
xor UO_553 (O_553,N_8410,N_9407);
xnor UO_554 (O_554,N_9219,N_8358);
xnor UO_555 (O_555,N_8917,N_9855);
or UO_556 (O_556,N_9347,N_8259);
xnor UO_557 (O_557,N_9754,N_8386);
or UO_558 (O_558,N_9585,N_9566);
nand UO_559 (O_559,N_8983,N_9583);
nor UO_560 (O_560,N_8267,N_8206);
xnor UO_561 (O_561,N_8417,N_8845);
or UO_562 (O_562,N_8300,N_8978);
and UO_563 (O_563,N_8012,N_9148);
or UO_564 (O_564,N_8751,N_9884);
nand UO_565 (O_565,N_9630,N_9888);
nor UO_566 (O_566,N_8222,N_8232);
nand UO_567 (O_567,N_9118,N_9168);
and UO_568 (O_568,N_8239,N_8783);
nand UO_569 (O_569,N_9019,N_9342);
nor UO_570 (O_570,N_8467,N_9402);
nand UO_571 (O_571,N_8891,N_9451);
nand UO_572 (O_572,N_9594,N_9109);
nor UO_573 (O_573,N_8980,N_9760);
nor UO_574 (O_574,N_9642,N_8919);
xor UO_575 (O_575,N_9178,N_8628);
or UO_576 (O_576,N_8687,N_9778);
nor UO_577 (O_577,N_8402,N_8673);
nor UO_578 (O_578,N_8018,N_8525);
or UO_579 (O_579,N_9406,N_8308);
and UO_580 (O_580,N_8789,N_8005);
or UO_581 (O_581,N_8463,N_8840);
nor UO_582 (O_582,N_9607,N_8104);
nor UO_583 (O_583,N_9244,N_8517);
xnor UO_584 (O_584,N_8523,N_8561);
xor UO_585 (O_585,N_9267,N_9877);
xnor UO_586 (O_586,N_9663,N_9765);
xnor UO_587 (O_587,N_9743,N_9834);
nand UO_588 (O_588,N_9075,N_9269);
or UO_589 (O_589,N_8934,N_8882);
nand UO_590 (O_590,N_8154,N_9035);
nand UO_591 (O_591,N_9999,N_8459);
or UO_592 (O_592,N_8324,N_8860);
xnor UO_593 (O_593,N_8609,N_9470);
xnor UO_594 (O_594,N_8235,N_9058);
nor UO_595 (O_595,N_9039,N_8373);
nor UO_596 (O_596,N_8957,N_9332);
nand UO_597 (O_597,N_8177,N_9084);
nand UO_598 (O_598,N_9442,N_8723);
or UO_599 (O_599,N_8621,N_8100);
or UO_600 (O_600,N_8890,N_8912);
nand UO_601 (O_601,N_9751,N_9629);
and UO_602 (O_602,N_9054,N_8803);
nand UO_603 (O_603,N_8210,N_9495);
or UO_604 (O_604,N_8359,N_9909);
and UO_605 (O_605,N_8851,N_9828);
nor UO_606 (O_606,N_9848,N_8762);
and UO_607 (O_607,N_8835,N_9927);
nor UO_608 (O_608,N_9882,N_8268);
and UO_609 (O_609,N_8338,N_8757);
and UO_610 (O_610,N_9144,N_9505);
xnor UO_611 (O_611,N_9653,N_9894);
or UO_612 (O_612,N_9738,N_9641);
xnor UO_613 (O_613,N_9367,N_8884);
xor UO_614 (O_614,N_8925,N_9480);
nor UO_615 (O_615,N_9112,N_8091);
nor UO_616 (O_616,N_9881,N_8288);
nand UO_617 (O_617,N_8101,N_8535);
and UO_618 (O_618,N_9672,N_8138);
nand UO_619 (O_619,N_9257,N_8035);
nand UO_620 (O_620,N_8002,N_9602);
xnor UO_621 (O_621,N_9241,N_9053);
nor UO_622 (O_622,N_8646,N_9186);
nor UO_623 (O_623,N_8926,N_9702);
and UO_624 (O_624,N_8938,N_9673);
and UO_625 (O_625,N_9717,N_8054);
and UO_626 (O_626,N_8703,N_9421);
and UO_627 (O_627,N_9849,N_9005);
or UO_628 (O_628,N_8360,N_8127);
and UO_629 (O_629,N_8401,N_8689);
nand UO_630 (O_630,N_8587,N_9108);
or UO_631 (O_631,N_8307,N_9831);
and UO_632 (O_632,N_9105,N_8932);
and UO_633 (O_633,N_8349,N_8805);
nor UO_634 (O_634,N_9388,N_9196);
or UO_635 (O_635,N_8074,N_9939);
nor UO_636 (O_636,N_8534,N_9759);
xnor UO_637 (O_637,N_9720,N_9992);
xor UO_638 (O_638,N_8854,N_9373);
or UO_639 (O_639,N_8529,N_9665);
and UO_640 (O_640,N_8069,N_9082);
or UO_641 (O_641,N_9776,N_9993);
and UO_642 (O_642,N_8677,N_9438);
nor UO_643 (O_643,N_8596,N_9157);
nor UO_644 (O_644,N_8001,N_9588);
xor UO_645 (O_645,N_9867,N_8484);
and UO_646 (O_646,N_8952,N_9586);
nor UO_647 (O_647,N_8948,N_9125);
nand UO_648 (O_648,N_9208,N_8049);
nor UO_649 (O_649,N_9537,N_8900);
and UO_650 (O_650,N_8446,N_8922);
xor UO_651 (O_651,N_8135,N_8521);
nand UO_652 (O_652,N_9865,N_8799);
or UO_653 (O_653,N_8251,N_9959);
xnor UO_654 (O_654,N_9120,N_8309);
and UO_655 (O_655,N_8741,N_8149);
nor UO_656 (O_656,N_9376,N_8732);
nand UO_657 (O_657,N_8556,N_8839);
nand UO_658 (O_658,N_8326,N_8727);
xor UO_659 (O_659,N_8060,N_8369);
or UO_660 (O_660,N_8877,N_9655);
nor UO_661 (O_661,N_9696,N_8516);
and UO_662 (O_662,N_9725,N_8292);
xor UO_663 (O_663,N_8449,N_8573);
and UO_664 (O_664,N_8511,N_9056);
and UO_665 (O_665,N_9929,N_9036);
nand UO_666 (O_666,N_8549,N_9563);
and UO_667 (O_667,N_8294,N_8260);
and UO_668 (O_668,N_8161,N_9013);
nand UO_669 (O_669,N_9285,N_8701);
and UO_670 (O_670,N_8117,N_8666);
nand UO_671 (O_671,N_8175,N_9464);
nor UO_672 (O_672,N_9636,N_9466);
xor UO_673 (O_673,N_9460,N_9928);
or UO_674 (O_674,N_8509,N_8053);
xor UO_675 (O_675,N_9147,N_8618);
nand UO_676 (O_676,N_9942,N_8997);
and UO_677 (O_677,N_9635,N_8327);
nand UO_678 (O_678,N_9212,N_9637);
xor UO_679 (O_679,N_9678,N_9767);
or UO_680 (O_680,N_9124,N_8004);
xnor UO_681 (O_681,N_8504,N_9245);
nor UO_682 (O_682,N_8275,N_8299);
and UO_683 (O_683,N_8878,N_8347);
nor UO_684 (O_684,N_8812,N_8967);
or UO_685 (O_685,N_8594,N_8181);
or UO_686 (O_686,N_8691,N_8087);
nand UO_687 (O_687,N_9381,N_9739);
and UO_688 (O_688,N_8085,N_9951);
and UO_689 (O_689,N_9868,N_8337);
nand UO_690 (O_690,N_9323,N_9242);
and UO_691 (O_691,N_8136,N_9694);
nor UO_692 (O_692,N_8955,N_9750);
nor UO_693 (O_693,N_9768,N_9428);
or UO_694 (O_694,N_8397,N_8578);
and UO_695 (O_695,N_8802,N_9758);
xor UO_696 (O_696,N_9572,N_8400);
nand UO_697 (O_697,N_8283,N_8064);
and UO_698 (O_698,N_9430,N_9509);
nor UO_699 (O_699,N_8316,N_9210);
nand UO_700 (O_700,N_8067,N_8147);
nand UO_701 (O_701,N_9301,N_9284);
or UO_702 (O_702,N_9772,N_9136);
or UO_703 (O_703,N_8301,N_8608);
or UO_704 (O_704,N_9247,N_8625);
nand UO_705 (O_705,N_8109,N_9397);
nor UO_706 (O_706,N_9104,N_8985);
and UO_707 (O_707,N_8442,N_8250);
xor UO_708 (O_708,N_9444,N_8137);
nand UO_709 (O_709,N_8388,N_9154);
nand UO_710 (O_710,N_8915,N_9279);
xnor UO_711 (O_711,N_9646,N_8224);
nand UO_712 (O_712,N_9654,N_9418);
xor UO_713 (O_713,N_9691,N_8694);
or UO_714 (O_714,N_9531,N_9253);
nor UO_715 (O_715,N_8121,N_9649);
or UO_716 (O_716,N_9318,N_8933);
nand UO_717 (O_717,N_9405,N_8927);
nor UO_718 (O_718,N_9763,N_8219);
nand UO_719 (O_719,N_8546,N_9911);
xor UO_720 (O_720,N_9385,N_9916);
xor UO_721 (O_721,N_8660,N_9786);
and UO_722 (O_722,N_8921,N_9803);
or UO_723 (O_723,N_8548,N_8894);
nor UO_724 (O_724,N_8867,N_8844);
nor UO_725 (O_725,N_9326,N_9896);
xnor UO_726 (O_726,N_8427,N_9816);
nand UO_727 (O_727,N_9715,N_9543);
xor UO_728 (O_728,N_9698,N_9010);
and UO_729 (O_729,N_9944,N_9432);
nor UO_730 (O_730,N_8180,N_9661);
and UO_731 (O_731,N_8970,N_8178);
nand UO_732 (O_732,N_8966,N_9425);
xnor UO_733 (O_733,N_9188,N_9792);
xor UO_734 (O_734,N_9399,N_9785);
nand UO_735 (O_735,N_8515,N_8533);
and UO_736 (O_736,N_9410,N_9741);
and UO_737 (O_737,N_9825,N_8409);
nand UO_738 (O_738,N_9525,N_8377);
or UO_739 (O_739,N_8351,N_9575);
xnor UO_740 (O_740,N_8730,N_8801);
or UO_741 (O_741,N_9151,N_9341);
and UO_742 (O_742,N_8141,N_9252);
xnor UO_743 (O_743,N_9096,N_9973);
nor UO_744 (O_744,N_8959,N_8663);
nor UO_745 (O_745,N_8221,N_8896);
xor UO_746 (O_746,N_8905,N_8404);
xnor UO_747 (O_747,N_8398,N_8039);
nand UO_748 (O_748,N_9612,N_9363);
nor UO_749 (O_749,N_9920,N_8930);
and UO_750 (O_750,N_9718,N_9824);
and UO_751 (O_751,N_8375,N_8242);
xnor UO_752 (O_752,N_8227,N_8192);
or UO_753 (O_753,N_8725,N_9477);
and UO_754 (O_754,N_9083,N_8707);
nand UO_755 (O_755,N_9073,N_9807);
nor UO_756 (O_756,N_9472,N_9921);
or UO_757 (O_757,N_9274,N_8686);
nor UO_758 (O_758,N_9937,N_9067);
nor UO_759 (O_759,N_9199,N_9887);
or UO_760 (O_760,N_8564,N_9747);
and UO_761 (O_761,N_8856,N_8974);
or UO_762 (O_762,N_9291,N_9417);
xor UO_763 (O_763,N_8763,N_9111);
xnor UO_764 (O_764,N_9335,N_9788);
and UO_765 (O_765,N_8476,N_9783);
nand UO_766 (O_766,N_8592,N_8478);
and UO_767 (O_767,N_8624,N_8773);
and UO_768 (O_768,N_9685,N_9282);
xor UO_769 (O_769,N_8700,N_8612);
or UO_770 (O_770,N_8457,N_8828);
or UO_771 (O_771,N_9103,N_9817);
nor UO_772 (O_772,N_8895,N_9251);
or UO_773 (O_773,N_9774,N_9311);
and UO_774 (O_774,N_8685,N_9991);
nor UO_775 (O_775,N_9643,N_8107);
nor UO_776 (O_776,N_9040,N_9437);
nor UO_777 (O_777,N_9811,N_8836);
and UO_778 (O_778,N_9900,N_9592);
or UO_779 (O_779,N_8248,N_9516);
nor UO_780 (O_780,N_9826,N_8570);
or UO_781 (O_781,N_8438,N_8112);
or UO_782 (O_782,N_8532,N_9471);
or UO_783 (O_783,N_8196,N_9963);
or UO_784 (O_784,N_9458,N_9447);
or UO_785 (O_785,N_8559,N_9288);
nor UO_786 (O_786,N_9512,N_9275);
or UO_787 (O_787,N_9197,N_8960);
nor UO_788 (O_788,N_8425,N_8719);
and UO_789 (O_789,N_8885,N_8126);
and UO_790 (O_790,N_8348,N_9647);
nand UO_791 (O_791,N_8735,N_9987);
nand UO_792 (O_792,N_8806,N_8740);
or UO_793 (O_793,N_8971,N_9158);
or UO_794 (O_794,N_8033,N_9303);
nor UO_795 (O_795,N_8379,N_9652);
nand UO_796 (O_796,N_8942,N_9370);
nor UO_797 (O_797,N_8920,N_9827);
or UO_798 (O_798,N_9423,N_9740);
xor UO_799 (O_799,N_9620,N_9713);
and UO_800 (O_800,N_8408,N_9490);
xor UO_801 (O_801,N_8371,N_8946);
xor UO_802 (O_802,N_9617,N_8176);
or UO_803 (O_803,N_8394,N_9246);
or UO_804 (O_804,N_8986,N_8651);
nand UO_805 (O_805,N_8133,N_8888);
nor UO_806 (O_806,N_8715,N_9623);
nor UO_807 (O_807,N_9434,N_9162);
nand UO_808 (O_808,N_9530,N_9708);
xor UO_809 (O_809,N_8487,N_8620);
or UO_810 (O_810,N_8350,N_8321);
xnor UO_811 (O_811,N_9680,N_9383);
xnor UO_812 (O_812,N_8432,N_8443);
xnor UO_813 (O_813,N_9926,N_9334);
nor UO_814 (O_814,N_9769,N_9571);
xnor UO_815 (O_815,N_8212,N_8610);
xor UO_816 (O_816,N_8543,N_9508);
nor UO_817 (O_817,N_9998,N_8023);
nor UO_818 (O_818,N_9138,N_8266);
or UO_819 (O_819,N_9392,N_9365);
nand UO_820 (O_820,N_9519,N_9420);
or UO_821 (O_821,N_9018,N_9576);
nor UO_822 (O_822,N_9736,N_8597);
nor UO_823 (O_823,N_9045,N_9400);
xor UO_824 (O_824,N_8774,N_9902);
and UO_825 (O_825,N_9070,N_8263);
and UO_826 (O_826,N_9292,N_9507);
nor UO_827 (O_827,N_8111,N_9878);
and UO_828 (O_828,N_8585,N_9851);
xor UO_829 (O_829,N_9577,N_8174);
nand UO_830 (O_830,N_8759,N_8781);
xnor UO_831 (O_831,N_9236,N_8605);
or UO_832 (O_832,N_9520,N_8293);
and UO_833 (O_833,N_9616,N_8125);
nand UO_834 (O_834,N_9626,N_8302);
or UO_835 (O_835,N_8760,N_9775);
or UO_836 (O_836,N_8143,N_9818);
nor UO_837 (O_837,N_9455,N_8531);
nor UO_838 (O_838,N_8993,N_9628);
xnor UO_839 (O_839,N_8695,N_8650);
or UO_840 (O_840,N_9871,N_9953);
nor UO_841 (O_841,N_8820,N_8755);
nor UO_842 (O_842,N_9079,N_9088);
or UO_843 (O_843,N_8992,N_8644);
and UO_844 (O_844,N_9830,N_8273);
nand UO_845 (O_845,N_8756,N_8841);
and UO_846 (O_846,N_9137,N_8430);
nand UO_847 (O_847,N_9302,N_8598);
and UO_848 (O_848,N_8205,N_8503);
or UO_849 (O_849,N_9032,N_9801);
and UO_850 (O_850,N_9957,N_9872);
xor UO_851 (O_851,N_9985,N_9426);
xnor UO_852 (O_852,N_9904,N_8441);
and UO_853 (O_853,N_8220,N_8562);
or UO_854 (O_854,N_9722,N_8632);
nor UO_855 (O_855,N_8384,N_9306);
nor UO_856 (O_856,N_9283,N_9090);
nand UO_857 (O_857,N_9143,N_8658);
or UO_858 (O_858,N_9413,N_8378);
nor UO_859 (O_859,N_9193,N_8743);
xor UO_860 (O_860,N_8217,N_8078);
xor UO_861 (O_861,N_8072,N_8013);
nor UO_862 (O_862,N_8464,N_8195);
or UO_863 (O_863,N_9907,N_8420);
xor UO_864 (O_864,N_8277,N_8353);
xnor UO_865 (O_865,N_8092,N_9613);
nand UO_866 (O_866,N_8843,N_9522);
and UO_867 (O_867,N_9839,N_9062);
or UO_868 (O_868,N_9166,N_9518);
nor UO_869 (O_869,N_9448,N_9263);
nor UO_870 (O_870,N_9946,N_9737);
and UO_871 (O_871,N_8746,N_9012);
or UO_872 (O_872,N_9995,N_8595);
nand UO_873 (O_873,N_9688,N_9802);
and UO_874 (O_874,N_9600,N_9989);
nor UO_875 (O_875,N_9362,N_9521);
and UO_876 (O_876,N_9862,N_9355);
nand UO_877 (O_877,N_8026,N_9943);
nor UO_878 (O_878,N_8810,N_9631);
or UO_879 (O_879,N_9961,N_9883);
xnor UO_880 (O_880,N_9528,N_8982);
or UO_881 (O_881,N_9300,N_8636);
nand UO_882 (O_882,N_8372,N_8142);
or UO_883 (O_883,N_8184,N_8640);
nor UO_884 (O_884,N_8642,N_9569);
and UO_885 (O_885,N_8869,N_8567);
and UO_886 (O_886,N_9982,N_8031);
xnor UO_887 (O_887,N_8698,N_9161);
nand UO_888 (O_888,N_9650,N_9213);
xnor UO_889 (O_889,N_8167,N_8889);
nand UO_890 (O_890,N_8502,N_8572);
xor UO_891 (O_891,N_9478,N_8155);
xnor UO_892 (O_892,N_9243,N_9181);
xor UO_893 (O_893,N_8536,N_9092);
and UO_894 (O_894,N_9684,N_8156);
nand UO_895 (O_895,N_9130,N_8159);
nor UO_896 (O_896,N_9972,N_9853);
or UO_897 (O_897,N_8816,N_9979);
or UO_898 (O_898,N_9324,N_8437);
nor UO_899 (O_899,N_9327,N_8010);
nor UO_900 (O_900,N_9081,N_8769);
xnor UO_901 (O_901,N_9941,N_9000);
nor UO_902 (O_902,N_8204,N_9255);
and UO_903 (O_903,N_9248,N_9748);
or UO_904 (O_904,N_8086,N_9633);
and UO_905 (O_905,N_8600,N_9782);
and UO_906 (O_906,N_9535,N_9184);
xor UO_907 (O_907,N_8714,N_8748);
or UO_908 (O_908,N_8403,N_8482);
and UO_909 (O_909,N_8296,N_8332);
nand UO_910 (O_910,N_9668,N_9732);
or UO_911 (O_911,N_8737,N_9382);
xnor UO_912 (O_912,N_9805,N_9379);
nor UO_913 (O_913,N_8276,N_8346);
nand UO_914 (O_914,N_9414,N_8345);
xor UO_915 (O_915,N_8583,N_9159);
xor UO_916 (O_916,N_9214,N_9931);
xor UO_917 (O_917,N_8507,N_9579);
or UO_918 (O_918,N_8465,N_8892);
nand UO_919 (O_919,N_8961,N_9331);
or UO_920 (O_920,N_9256,N_8571);
or UO_921 (O_921,N_8322,N_8508);
nor UO_922 (O_922,N_9844,N_9209);
and UO_923 (O_923,N_8458,N_9703);
nor UO_924 (O_924,N_9391,N_9794);
xnor UO_925 (O_925,N_9309,N_8048);
nand UO_926 (O_926,N_9220,N_9660);
and UO_927 (O_927,N_9689,N_8190);
nor UO_928 (O_928,N_8245,N_8958);
or UO_929 (O_929,N_8808,N_8148);
nand UO_930 (O_930,N_8129,N_8015);
xnor UO_931 (O_931,N_9361,N_8257);
nor UO_932 (O_932,N_9605,N_8832);
nand UO_933 (O_933,N_9771,N_9325);
or UO_934 (O_934,N_9175,N_8939);
xor UO_935 (O_935,N_9369,N_8431);
xnor UO_936 (O_936,N_8490,N_8795);
nand UO_937 (O_937,N_9822,N_9560);
and UO_938 (O_938,N_9307,N_9833);
xor UO_939 (O_939,N_9974,N_8025);
and UO_940 (O_940,N_8555,N_8233);
nor UO_941 (O_941,N_8407,N_8079);
xor UO_942 (O_942,N_8791,N_9670);
xnor UO_943 (O_943,N_8513,N_8575);
and UO_944 (O_944,N_9510,N_8692);
nor UO_945 (O_945,N_9885,N_9744);
and UO_946 (O_946,N_8793,N_9766);
xor UO_947 (O_947,N_9164,N_8788);
xor UO_948 (O_948,N_8165,N_8943);
or UO_949 (O_949,N_9360,N_8460);
and UO_950 (O_950,N_8526,N_9693);
xnor UO_951 (O_951,N_8604,N_8481);
nand UO_952 (O_952,N_8990,N_8057);
or UO_953 (O_953,N_8341,N_8776);
or UO_954 (O_954,N_9270,N_9487);
and UO_955 (O_955,N_8838,N_8406);
or UO_956 (O_956,N_8904,N_9389);
nand UO_957 (O_957,N_8648,N_8833);
or UO_958 (O_958,N_9634,N_9624);
xor UO_959 (O_959,N_8954,N_9102);
and UO_960 (O_960,N_9333,N_9134);
nand UO_961 (O_961,N_8208,N_8390);
and UO_962 (O_962,N_9797,N_9555);
or UO_963 (O_963,N_8736,N_9135);
xnor UO_964 (O_964,N_9093,N_9482);
and UO_965 (O_965,N_8000,N_8071);
xor UO_966 (O_966,N_9761,N_8897);
nor UO_967 (O_967,N_8200,N_8989);
nor UO_968 (O_968,N_8797,N_8106);
nor UO_969 (O_969,N_9007,N_8846);
nand UO_970 (O_970,N_8964,N_8270);
or UO_971 (O_971,N_8382,N_8654);
nor UO_972 (O_972,N_9756,N_9076);
nor UO_973 (O_973,N_8613,N_9491);
nor UO_974 (O_974,N_8824,N_8278);
nand UO_975 (O_975,N_9930,N_9354);
xor UO_976 (O_976,N_8558,N_9550);
and UO_977 (O_977,N_8678,N_9265);
or UO_978 (O_978,N_9544,N_8132);
and UO_979 (O_979,N_9259,N_9870);
nor UO_980 (O_980,N_9277,N_9249);
nand UO_981 (O_981,N_8569,N_9864);
or UO_982 (O_982,N_8779,N_9195);
or UO_983 (O_983,N_9496,N_9651);
or UO_984 (O_984,N_9254,N_9662);
nor UO_985 (O_985,N_8305,N_9934);
nor UO_986 (O_986,N_8834,N_8022);
and UO_987 (O_987,N_8780,N_8792);
and UO_988 (O_988,N_9173,N_8866);
or UO_989 (O_989,N_9043,N_9237);
xor UO_990 (O_990,N_9861,N_9287);
nand UO_991 (O_991,N_9952,N_8566);
nor UO_992 (O_992,N_8105,N_8306);
xor UO_993 (O_993,N_8818,N_8089);
or UO_994 (O_994,N_9286,N_8716);
nand UO_995 (O_995,N_8194,N_8794);
xor UO_996 (O_996,N_8761,N_9454);
or UO_997 (O_997,N_9174,N_8246);
xnor UO_998 (O_998,N_9063,N_8495);
nor UO_999 (O_999,N_8883,N_8120);
and UO_1000 (O_1000,N_9485,N_9680);
nand UO_1001 (O_1001,N_9326,N_9993);
or UO_1002 (O_1002,N_8166,N_9898);
xnor UO_1003 (O_1003,N_8892,N_8755);
and UO_1004 (O_1004,N_9684,N_8572);
xnor UO_1005 (O_1005,N_8263,N_9503);
nor UO_1006 (O_1006,N_8684,N_8441);
and UO_1007 (O_1007,N_9055,N_9164);
nor UO_1008 (O_1008,N_8889,N_8201);
nand UO_1009 (O_1009,N_8868,N_9666);
nor UO_1010 (O_1010,N_9981,N_9225);
or UO_1011 (O_1011,N_9074,N_9077);
or UO_1012 (O_1012,N_8050,N_9200);
and UO_1013 (O_1013,N_9282,N_9252);
or UO_1014 (O_1014,N_9602,N_9331);
nand UO_1015 (O_1015,N_8202,N_8545);
xor UO_1016 (O_1016,N_9967,N_9918);
nor UO_1017 (O_1017,N_9204,N_8964);
or UO_1018 (O_1018,N_8418,N_9172);
or UO_1019 (O_1019,N_8183,N_8899);
xnor UO_1020 (O_1020,N_9654,N_8020);
or UO_1021 (O_1021,N_8913,N_9512);
or UO_1022 (O_1022,N_8417,N_9995);
xnor UO_1023 (O_1023,N_8609,N_8878);
nor UO_1024 (O_1024,N_9872,N_8891);
and UO_1025 (O_1025,N_8178,N_8824);
or UO_1026 (O_1026,N_8729,N_9519);
nor UO_1027 (O_1027,N_9489,N_8290);
nor UO_1028 (O_1028,N_8370,N_9868);
or UO_1029 (O_1029,N_9546,N_9565);
and UO_1030 (O_1030,N_9149,N_8360);
or UO_1031 (O_1031,N_9002,N_9534);
and UO_1032 (O_1032,N_8066,N_9650);
xor UO_1033 (O_1033,N_9442,N_8306);
nand UO_1034 (O_1034,N_8826,N_8675);
and UO_1035 (O_1035,N_9744,N_9645);
or UO_1036 (O_1036,N_8180,N_9248);
nor UO_1037 (O_1037,N_9063,N_9152);
nand UO_1038 (O_1038,N_8702,N_9839);
xnor UO_1039 (O_1039,N_8486,N_9646);
xor UO_1040 (O_1040,N_8443,N_9931);
or UO_1041 (O_1041,N_9153,N_9749);
nand UO_1042 (O_1042,N_8591,N_8206);
or UO_1043 (O_1043,N_9803,N_9780);
nor UO_1044 (O_1044,N_8000,N_9797);
or UO_1045 (O_1045,N_9393,N_9958);
or UO_1046 (O_1046,N_8760,N_8204);
nand UO_1047 (O_1047,N_9477,N_8599);
and UO_1048 (O_1048,N_8154,N_9236);
and UO_1049 (O_1049,N_9743,N_8316);
nand UO_1050 (O_1050,N_8185,N_8462);
xor UO_1051 (O_1051,N_8992,N_9089);
and UO_1052 (O_1052,N_8473,N_8681);
and UO_1053 (O_1053,N_8507,N_8310);
or UO_1054 (O_1054,N_8350,N_9760);
nand UO_1055 (O_1055,N_9679,N_8081);
xnor UO_1056 (O_1056,N_9848,N_8555);
and UO_1057 (O_1057,N_9643,N_9480);
nor UO_1058 (O_1058,N_9520,N_8424);
and UO_1059 (O_1059,N_9068,N_8441);
xnor UO_1060 (O_1060,N_8568,N_9032);
nand UO_1061 (O_1061,N_8650,N_9312);
or UO_1062 (O_1062,N_9969,N_9619);
nand UO_1063 (O_1063,N_9882,N_9886);
xnor UO_1064 (O_1064,N_8473,N_9775);
nand UO_1065 (O_1065,N_9144,N_9313);
and UO_1066 (O_1066,N_8529,N_8084);
nand UO_1067 (O_1067,N_8520,N_9188);
or UO_1068 (O_1068,N_8058,N_9277);
nor UO_1069 (O_1069,N_9864,N_8893);
xnor UO_1070 (O_1070,N_9214,N_9076);
xnor UO_1071 (O_1071,N_8391,N_8561);
and UO_1072 (O_1072,N_9637,N_8501);
or UO_1073 (O_1073,N_8383,N_9589);
xnor UO_1074 (O_1074,N_8306,N_9090);
or UO_1075 (O_1075,N_8158,N_8291);
and UO_1076 (O_1076,N_8624,N_8459);
xnor UO_1077 (O_1077,N_8749,N_8875);
nand UO_1078 (O_1078,N_8867,N_8192);
or UO_1079 (O_1079,N_9346,N_9505);
nand UO_1080 (O_1080,N_9763,N_8746);
and UO_1081 (O_1081,N_9166,N_8459);
xnor UO_1082 (O_1082,N_8028,N_9805);
nand UO_1083 (O_1083,N_8842,N_9957);
xnor UO_1084 (O_1084,N_8092,N_8768);
nor UO_1085 (O_1085,N_8441,N_9825);
xnor UO_1086 (O_1086,N_9228,N_9423);
nor UO_1087 (O_1087,N_9620,N_9270);
nor UO_1088 (O_1088,N_8030,N_8046);
nand UO_1089 (O_1089,N_8593,N_9649);
and UO_1090 (O_1090,N_8816,N_8868);
or UO_1091 (O_1091,N_9898,N_9026);
xnor UO_1092 (O_1092,N_8188,N_8262);
and UO_1093 (O_1093,N_9078,N_8574);
or UO_1094 (O_1094,N_8345,N_9000);
xor UO_1095 (O_1095,N_8065,N_9017);
or UO_1096 (O_1096,N_8634,N_8449);
and UO_1097 (O_1097,N_8667,N_9643);
nand UO_1098 (O_1098,N_8239,N_8174);
nand UO_1099 (O_1099,N_8767,N_9589);
nor UO_1100 (O_1100,N_9507,N_9625);
nand UO_1101 (O_1101,N_8933,N_8332);
and UO_1102 (O_1102,N_8684,N_8860);
and UO_1103 (O_1103,N_9335,N_9801);
xor UO_1104 (O_1104,N_8511,N_8784);
nor UO_1105 (O_1105,N_8225,N_9259);
nor UO_1106 (O_1106,N_8862,N_8895);
xor UO_1107 (O_1107,N_8359,N_9374);
and UO_1108 (O_1108,N_8486,N_9859);
xnor UO_1109 (O_1109,N_9032,N_9199);
or UO_1110 (O_1110,N_9802,N_8578);
nor UO_1111 (O_1111,N_8082,N_9558);
xnor UO_1112 (O_1112,N_8944,N_8417);
or UO_1113 (O_1113,N_8052,N_9716);
nor UO_1114 (O_1114,N_9110,N_8688);
or UO_1115 (O_1115,N_9173,N_8555);
nand UO_1116 (O_1116,N_9907,N_8450);
or UO_1117 (O_1117,N_8459,N_9487);
nand UO_1118 (O_1118,N_8671,N_8882);
nand UO_1119 (O_1119,N_9903,N_8568);
nand UO_1120 (O_1120,N_8420,N_8746);
xor UO_1121 (O_1121,N_8642,N_8657);
nor UO_1122 (O_1122,N_9042,N_9791);
xnor UO_1123 (O_1123,N_8269,N_8149);
xnor UO_1124 (O_1124,N_8350,N_8787);
or UO_1125 (O_1125,N_8434,N_9234);
nand UO_1126 (O_1126,N_9129,N_8427);
or UO_1127 (O_1127,N_8717,N_9221);
and UO_1128 (O_1128,N_9252,N_9939);
and UO_1129 (O_1129,N_9973,N_8573);
and UO_1130 (O_1130,N_8984,N_9209);
nor UO_1131 (O_1131,N_9201,N_9760);
or UO_1132 (O_1132,N_9335,N_9530);
nor UO_1133 (O_1133,N_8838,N_8294);
xnor UO_1134 (O_1134,N_9381,N_8188);
and UO_1135 (O_1135,N_9230,N_9978);
xor UO_1136 (O_1136,N_9726,N_9378);
nor UO_1137 (O_1137,N_9422,N_8582);
and UO_1138 (O_1138,N_8987,N_8574);
nor UO_1139 (O_1139,N_9254,N_9216);
and UO_1140 (O_1140,N_9138,N_9083);
and UO_1141 (O_1141,N_8273,N_9855);
or UO_1142 (O_1142,N_8730,N_8813);
or UO_1143 (O_1143,N_8694,N_9960);
nor UO_1144 (O_1144,N_8539,N_8499);
nor UO_1145 (O_1145,N_9267,N_9561);
nor UO_1146 (O_1146,N_8598,N_8597);
nand UO_1147 (O_1147,N_9262,N_9025);
nand UO_1148 (O_1148,N_9798,N_8454);
or UO_1149 (O_1149,N_8327,N_8594);
xnor UO_1150 (O_1150,N_9883,N_9240);
xnor UO_1151 (O_1151,N_9518,N_8330);
xnor UO_1152 (O_1152,N_9690,N_8012);
and UO_1153 (O_1153,N_8180,N_9495);
nand UO_1154 (O_1154,N_8546,N_8110);
nor UO_1155 (O_1155,N_9842,N_8794);
or UO_1156 (O_1156,N_9304,N_8786);
xor UO_1157 (O_1157,N_8835,N_9479);
nor UO_1158 (O_1158,N_9027,N_8114);
nor UO_1159 (O_1159,N_9775,N_9064);
xor UO_1160 (O_1160,N_8068,N_8997);
and UO_1161 (O_1161,N_8283,N_8769);
or UO_1162 (O_1162,N_8022,N_9383);
nor UO_1163 (O_1163,N_8369,N_9976);
xnor UO_1164 (O_1164,N_9370,N_9295);
nand UO_1165 (O_1165,N_9404,N_8580);
and UO_1166 (O_1166,N_9164,N_9872);
or UO_1167 (O_1167,N_9667,N_9779);
and UO_1168 (O_1168,N_8155,N_8347);
xnor UO_1169 (O_1169,N_8124,N_8121);
and UO_1170 (O_1170,N_9230,N_9317);
nor UO_1171 (O_1171,N_9246,N_9404);
xnor UO_1172 (O_1172,N_9939,N_8589);
nand UO_1173 (O_1173,N_8548,N_8623);
and UO_1174 (O_1174,N_8510,N_8010);
nand UO_1175 (O_1175,N_9511,N_8100);
and UO_1176 (O_1176,N_9822,N_8357);
nor UO_1177 (O_1177,N_9301,N_9249);
nor UO_1178 (O_1178,N_9159,N_8743);
nor UO_1179 (O_1179,N_8610,N_8316);
and UO_1180 (O_1180,N_9084,N_9835);
nand UO_1181 (O_1181,N_8657,N_9549);
or UO_1182 (O_1182,N_9962,N_8567);
and UO_1183 (O_1183,N_8753,N_8296);
or UO_1184 (O_1184,N_8645,N_9978);
and UO_1185 (O_1185,N_8011,N_8411);
nand UO_1186 (O_1186,N_9586,N_8864);
nand UO_1187 (O_1187,N_8745,N_9103);
nand UO_1188 (O_1188,N_8119,N_8159);
xnor UO_1189 (O_1189,N_9662,N_9581);
xor UO_1190 (O_1190,N_9527,N_9962);
or UO_1191 (O_1191,N_8550,N_9929);
xor UO_1192 (O_1192,N_8744,N_8763);
and UO_1193 (O_1193,N_9696,N_9197);
xnor UO_1194 (O_1194,N_9796,N_9123);
or UO_1195 (O_1195,N_9172,N_8326);
nand UO_1196 (O_1196,N_9904,N_9886);
and UO_1197 (O_1197,N_9558,N_8927);
xor UO_1198 (O_1198,N_8129,N_9017);
nand UO_1199 (O_1199,N_9613,N_8681);
nor UO_1200 (O_1200,N_9948,N_8330);
nor UO_1201 (O_1201,N_8394,N_9746);
or UO_1202 (O_1202,N_8134,N_9944);
or UO_1203 (O_1203,N_8721,N_8131);
or UO_1204 (O_1204,N_8941,N_8017);
nor UO_1205 (O_1205,N_8399,N_8207);
xnor UO_1206 (O_1206,N_9895,N_9397);
or UO_1207 (O_1207,N_9927,N_8720);
nand UO_1208 (O_1208,N_8682,N_9662);
xor UO_1209 (O_1209,N_8242,N_9003);
nor UO_1210 (O_1210,N_9503,N_8949);
nand UO_1211 (O_1211,N_9454,N_8746);
nor UO_1212 (O_1212,N_8229,N_8066);
and UO_1213 (O_1213,N_8805,N_8381);
nand UO_1214 (O_1214,N_8935,N_9603);
and UO_1215 (O_1215,N_9700,N_8282);
or UO_1216 (O_1216,N_8026,N_8535);
or UO_1217 (O_1217,N_9298,N_9415);
nor UO_1218 (O_1218,N_9652,N_8563);
and UO_1219 (O_1219,N_9174,N_9152);
and UO_1220 (O_1220,N_9116,N_8619);
xnor UO_1221 (O_1221,N_8653,N_8629);
nor UO_1222 (O_1222,N_9293,N_8979);
xor UO_1223 (O_1223,N_9300,N_8416);
nor UO_1224 (O_1224,N_9886,N_9101);
nor UO_1225 (O_1225,N_8658,N_8322);
nor UO_1226 (O_1226,N_9540,N_8316);
xnor UO_1227 (O_1227,N_8307,N_8369);
nand UO_1228 (O_1228,N_9029,N_9227);
or UO_1229 (O_1229,N_9707,N_9950);
and UO_1230 (O_1230,N_9731,N_9162);
xnor UO_1231 (O_1231,N_8802,N_9102);
and UO_1232 (O_1232,N_9007,N_9937);
xor UO_1233 (O_1233,N_8643,N_8473);
nor UO_1234 (O_1234,N_9211,N_9577);
or UO_1235 (O_1235,N_8426,N_8317);
nor UO_1236 (O_1236,N_8205,N_8889);
nand UO_1237 (O_1237,N_9212,N_8054);
or UO_1238 (O_1238,N_9210,N_9118);
nor UO_1239 (O_1239,N_8438,N_8108);
nor UO_1240 (O_1240,N_9774,N_9042);
and UO_1241 (O_1241,N_8839,N_9136);
or UO_1242 (O_1242,N_8727,N_9168);
or UO_1243 (O_1243,N_9685,N_8135);
xor UO_1244 (O_1244,N_9509,N_9505);
and UO_1245 (O_1245,N_8653,N_8057);
nor UO_1246 (O_1246,N_9908,N_9875);
nand UO_1247 (O_1247,N_9125,N_9079);
nand UO_1248 (O_1248,N_8885,N_9234);
nor UO_1249 (O_1249,N_8499,N_8254);
nor UO_1250 (O_1250,N_8855,N_9128);
nand UO_1251 (O_1251,N_9883,N_8784);
or UO_1252 (O_1252,N_8708,N_8836);
xnor UO_1253 (O_1253,N_8492,N_8207);
and UO_1254 (O_1254,N_8476,N_9813);
or UO_1255 (O_1255,N_8073,N_8280);
and UO_1256 (O_1256,N_9881,N_9809);
and UO_1257 (O_1257,N_9595,N_8688);
or UO_1258 (O_1258,N_9455,N_8606);
xor UO_1259 (O_1259,N_9682,N_8840);
xnor UO_1260 (O_1260,N_9719,N_8715);
nor UO_1261 (O_1261,N_9067,N_8989);
and UO_1262 (O_1262,N_8888,N_8969);
or UO_1263 (O_1263,N_9661,N_8459);
or UO_1264 (O_1264,N_8694,N_8658);
xnor UO_1265 (O_1265,N_9824,N_8082);
nor UO_1266 (O_1266,N_9451,N_8369);
nand UO_1267 (O_1267,N_8209,N_9482);
nor UO_1268 (O_1268,N_8037,N_8189);
or UO_1269 (O_1269,N_8034,N_8903);
and UO_1270 (O_1270,N_9125,N_8184);
and UO_1271 (O_1271,N_9697,N_9651);
nand UO_1272 (O_1272,N_9899,N_8146);
xnor UO_1273 (O_1273,N_8160,N_8364);
nand UO_1274 (O_1274,N_9665,N_9580);
nand UO_1275 (O_1275,N_9890,N_9366);
nor UO_1276 (O_1276,N_9276,N_9973);
xor UO_1277 (O_1277,N_8489,N_9222);
nor UO_1278 (O_1278,N_9680,N_8669);
or UO_1279 (O_1279,N_9521,N_9390);
nand UO_1280 (O_1280,N_8172,N_9453);
and UO_1281 (O_1281,N_9662,N_8986);
and UO_1282 (O_1282,N_9853,N_8006);
nor UO_1283 (O_1283,N_8564,N_9883);
and UO_1284 (O_1284,N_9206,N_8341);
or UO_1285 (O_1285,N_8136,N_9646);
nor UO_1286 (O_1286,N_8750,N_8326);
nand UO_1287 (O_1287,N_8837,N_9379);
nand UO_1288 (O_1288,N_9844,N_9095);
nand UO_1289 (O_1289,N_8880,N_9717);
or UO_1290 (O_1290,N_9508,N_9727);
or UO_1291 (O_1291,N_9410,N_9789);
nor UO_1292 (O_1292,N_9700,N_9870);
nor UO_1293 (O_1293,N_8645,N_8210);
or UO_1294 (O_1294,N_8707,N_9883);
xor UO_1295 (O_1295,N_9485,N_8932);
and UO_1296 (O_1296,N_9276,N_8912);
nand UO_1297 (O_1297,N_8945,N_9288);
nor UO_1298 (O_1298,N_9971,N_9514);
nand UO_1299 (O_1299,N_9749,N_8994);
and UO_1300 (O_1300,N_9322,N_8209);
nand UO_1301 (O_1301,N_9584,N_9131);
nor UO_1302 (O_1302,N_9682,N_9207);
nor UO_1303 (O_1303,N_8276,N_8094);
nand UO_1304 (O_1304,N_9464,N_8050);
or UO_1305 (O_1305,N_8686,N_9098);
nor UO_1306 (O_1306,N_9653,N_8147);
xor UO_1307 (O_1307,N_8254,N_8037);
and UO_1308 (O_1308,N_8552,N_8238);
or UO_1309 (O_1309,N_9978,N_9947);
nor UO_1310 (O_1310,N_8591,N_9309);
or UO_1311 (O_1311,N_8579,N_8591);
or UO_1312 (O_1312,N_8872,N_8644);
xor UO_1313 (O_1313,N_8445,N_9748);
xnor UO_1314 (O_1314,N_8820,N_9401);
nand UO_1315 (O_1315,N_8632,N_9526);
or UO_1316 (O_1316,N_9008,N_9097);
and UO_1317 (O_1317,N_9082,N_8983);
or UO_1318 (O_1318,N_8841,N_8107);
nand UO_1319 (O_1319,N_8785,N_8225);
or UO_1320 (O_1320,N_9270,N_8401);
nor UO_1321 (O_1321,N_8055,N_9128);
nor UO_1322 (O_1322,N_8144,N_8954);
xor UO_1323 (O_1323,N_9685,N_8819);
or UO_1324 (O_1324,N_9087,N_9911);
xor UO_1325 (O_1325,N_8039,N_9171);
nand UO_1326 (O_1326,N_9071,N_9353);
or UO_1327 (O_1327,N_9036,N_9987);
nor UO_1328 (O_1328,N_9629,N_9283);
and UO_1329 (O_1329,N_9320,N_9783);
xnor UO_1330 (O_1330,N_9203,N_9016);
xor UO_1331 (O_1331,N_8876,N_9760);
or UO_1332 (O_1332,N_9777,N_9981);
nor UO_1333 (O_1333,N_9640,N_8238);
nand UO_1334 (O_1334,N_8246,N_8178);
xor UO_1335 (O_1335,N_9644,N_8539);
or UO_1336 (O_1336,N_9720,N_8403);
nor UO_1337 (O_1337,N_8814,N_8642);
xnor UO_1338 (O_1338,N_8003,N_8316);
xor UO_1339 (O_1339,N_9832,N_9921);
nor UO_1340 (O_1340,N_9554,N_9003);
nand UO_1341 (O_1341,N_8065,N_8323);
nand UO_1342 (O_1342,N_9911,N_8676);
or UO_1343 (O_1343,N_9585,N_9944);
nand UO_1344 (O_1344,N_9380,N_9055);
xor UO_1345 (O_1345,N_9136,N_9879);
nor UO_1346 (O_1346,N_8316,N_8499);
nor UO_1347 (O_1347,N_9763,N_9668);
nor UO_1348 (O_1348,N_9454,N_9000);
nand UO_1349 (O_1349,N_9244,N_8285);
or UO_1350 (O_1350,N_8142,N_8566);
xor UO_1351 (O_1351,N_8950,N_8614);
xor UO_1352 (O_1352,N_9421,N_8338);
xnor UO_1353 (O_1353,N_9609,N_9344);
xnor UO_1354 (O_1354,N_9692,N_8167);
nor UO_1355 (O_1355,N_8820,N_8317);
or UO_1356 (O_1356,N_8347,N_9513);
nor UO_1357 (O_1357,N_9457,N_9257);
nor UO_1358 (O_1358,N_9803,N_8833);
nand UO_1359 (O_1359,N_9360,N_8374);
nor UO_1360 (O_1360,N_8656,N_9704);
and UO_1361 (O_1361,N_8976,N_9117);
and UO_1362 (O_1362,N_9135,N_9347);
and UO_1363 (O_1363,N_8380,N_8861);
nor UO_1364 (O_1364,N_8390,N_8158);
and UO_1365 (O_1365,N_8088,N_8996);
nor UO_1366 (O_1366,N_8552,N_9893);
nand UO_1367 (O_1367,N_9921,N_9038);
or UO_1368 (O_1368,N_8395,N_9124);
and UO_1369 (O_1369,N_8371,N_9601);
nor UO_1370 (O_1370,N_9916,N_8020);
or UO_1371 (O_1371,N_8484,N_9574);
or UO_1372 (O_1372,N_8943,N_9835);
nor UO_1373 (O_1373,N_8565,N_9261);
nand UO_1374 (O_1374,N_9123,N_9567);
nor UO_1375 (O_1375,N_8453,N_8808);
or UO_1376 (O_1376,N_9083,N_8048);
or UO_1377 (O_1377,N_9027,N_8282);
or UO_1378 (O_1378,N_8892,N_9446);
and UO_1379 (O_1379,N_8661,N_9910);
or UO_1380 (O_1380,N_8681,N_9071);
or UO_1381 (O_1381,N_8287,N_8472);
nand UO_1382 (O_1382,N_8058,N_9984);
or UO_1383 (O_1383,N_9013,N_8264);
and UO_1384 (O_1384,N_8947,N_8359);
or UO_1385 (O_1385,N_9411,N_9720);
or UO_1386 (O_1386,N_8447,N_8760);
nand UO_1387 (O_1387,N_8313,N_9474);
nor UO_1388 (O_1388,N_9708,N_8430);
xor UO_1389 (O_1389,N_9130,N_9472);
xor UO_1390 (O_1390,N_8663,N_9126);
and UO_1391 (O_1391,N_8711,N_8656);
nor UO_1392 (O_1392,N_9103,N_9498);
nor UO_1393 (O_1393,N_9485,N_8412);
or UO_1394 (O_1394,N_9424,N_8510);
and UO_1395 (O_1395,N_9823,N_9081);
and UO_1396 (O_1396,N_8465,N_9434);
nor UO_1397 (O_1397,N_9425,N_8995);
nand UO_1398 (O_1398,N_9662,N_9873);
nand UO_1399 (O_1399,N_9146,N_8595);
and UO_1400 (O_1400,N_8482,N_9192);
and UO_1401 (O_1401,N_9097,N_8842);
xnor UO_1402 (O_1402,N_8439,N_9828);
and UO_1403 (O_1403,N_8508,N_9538);
nand UO_1404 (O_1404,N_9160,N_9672);
nand UO_1405 (O_1405,N_8057,N_8092);
or UO_1406 (O_1406,N_8957,N_9692);
and UO_1407 (O_1407,N_9870,N_9472);
nor UO_1408 (O_1408,N_8244,N_9025);
and UO_1409 (O_1409,N_8505,N_9561);
nor UO_1410 (O_1410,N_9013,N_8431);
nor UO_1411 (O_1411,N_9127,N_9914);
nor UO_1412 (O_1412,N_8205,N_8306);
nor UO_1413 (O_1413,N_9657,N_9821);
nand UO_1414 (O_1414,N_8958,N_9103);
nor UO_1415 (O_1415,N_8418,N_8395);
or UO_1416 (O_1416,N_9640,N_9946);
or UO_1417 (O_1417,N_9175,N_9861);
nand UO_1418 (O_1418,N_8759,N_9767);
and UO_1419 (O_1419,N_8613,N_8884);
and UO_1420 (O_1420,N_9416,N_8993);
nor UO_1421 (O_1421,N_8105,N_9114);
and UO_1422 (O_1422,N_8907,N_9535);
nand UO_1423 (O_1423,N_8987,N_9553);
xnor UO_1424 (O_1424,N_8292,N_8844);
nor UO_1425 (O_1425,N_9927,N_9671);
or UO_1426 (O_1426,N_8048,N_9251);
xnor UO_1427 (O_1427,N_9226,N_8293);
xnor UO_1428 (O_1428,N_8985,N_8600);
or UO_1429 (O_1429,N_8356,N_9169);
or UO_1430 (O_1430,N_9113,N_8868);
xor UO_1431 (O_1431,N_8426,N_8034);
nand UO_1432 (O_1432,N_8159,N_9359);
xnor UO_1433 (O_1433,N_8329,N_9730);
nor UO_1434 (O_1434,N_8126,N_8246);
or UO_1435 (O_1435,N_8694,N_8852);
xnor UO_1436 (O_1436,N_8310,N_9470);
and UO_1437 (O_1437,N_8532,N_8680);
or UO_1438 (O_1438,N_9433,N_9616);
nor UO_1439 (O_1439,N_9702,N_9742);
nor UO_1440 (O_1440,N_9366,N_9206);
xor UO_1441 (O_1441,N_8307,N_8130);
and UO_1442 (O_1442,N_8842,N_8354);
xnor UO_1443 (O_1443,N_9059,N_8739);
and UO_1444 (O_1444,N_8780,N_8032);
nor UO_1445 (O_1445,N_8967,N_8989);
nand UO_1446 (O_1446,N_8097,N_8584);
xnor UO_1447 (O_1447,N_8337,N_8999);
xnor UO_1448 (O_1448,N_8995,N_9418);
xor UO_1449 (O_1449,N_9461,N_8962);
and UO_1450 (O_1450,N_9423,N_9151);
or UO_1451 (O_1451,N_8982,N_9421);
nand UO_1452 (O_1452,N_8660,N_9094);
nor UO_1453 (O_1453,N_8785,N_9052);
and UO_1454 (O_1454,N_9523,N_9670);
and UO_1455 (O_1455,N_9462,N_9847);
nand UO_1456 (O_1456,N_9513,N_9848);
nand UO_1457 (O_1457,N_8539,N_8389);
and UO_1458 (O_1458,N_9301,N_8068);
nand UO_1459 (O_1459,N_8128,N_9168);
xnor UO_1460 (O_1460,N_9420,N_9374);
nand UO_1461 (O_1461,N_8010,N_8514);
nand UO_1462 (O_1462,N_9597,N_8123);
nand UO_1463 (O_1463,N_8854,N_8838);
and UO_1464 (O_1464,N_9586,N_9181);
nor UO_1465 (O_1465,N_9745,N_8705);
nor UO_1466 (O_1466,N_8250,N_9167);
and UO_1467 (O_1467,N_9251,N_9319);
xnor UO_1468 (O_1468,N_9159,N_9723);
nand UO_1469 (O_1469,N_8303,N_9487);
nand UO_1470 (O_1470,N_8258,N_8686);
nor UO_1471 (O_1471,N_9927,N_8175);
and UO_1472 (O_1472,N_9828,N_9871);
xnor UO_1473 (O_1473,N_9496,N_8954);
nand UO_1474 (O_1474,N_9702,N_9874);
xnor UO_1475 (O_1475,N_8556,N_9083);
nand UO_1476 (O_1476,N_9666,N_8506);
or UO_1477 (O_1477,N_9663,N_8197);
nand UO_1478 (O_1478,N_9952,N_9121);
or UO_1479 (O_1479,N_8924,N_9382);
nor UO_1480 (O_1480,N_8344,N_8580);
nor UO_1481 (O_1481,N_9006,N_9654);
and UO_1482 (O_1482,N_9342,N_9903);
xor UO_1483 (O_1483,N_9333,N_9029);
nand UO_1484 (O_1484,N_9014,N_8845);
nor UO_1485 (O_1485,N_8183,N_9271);
nand UO_1486 (O_1486,N_8302,N_8578);
nand UO_1487 (O_1487,N_9110,N_9568);
xnor UO_1488 (O_1488,N_9793,N_9570);
and UO_1489 (O_1489,N_8108,N_8917);
nand UO_1490 (O_1490,N_9101,N_8415);
nor UO_1491 (O_1491,N_8511,N_8965);
and UO_1492 (O_1492,N_9655,N_9060);
xnor UO_1493 (O_1493,N_9736,N_9202);
nor UO_1494 (O_1494,N_8460,N_9216);
xnor UO_1495 (O_1495,N_8803,N_9212);
or UO_1496 (O_1496,N_9258,N_9483);
nand UO_1497 (O_1497,N_9047,N_8163);
or UO_1498 (O_1498,N_9077,N_8928);
and UO_1499 (O_1499,N_8267,N_9744);
endmodule