module basic_2000_20000_2500_25_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_1402,In_1522);
or U1 (N_1,In_268,In_1118);
and U2 (N_2,In_1550,In_709);
nand U3 (N_3,In_372,In_1670);
or U4 (N_4,In_1125,In_1327);
and U5 (N_5,In_985,In_137);
xor U6 (N_6,In_741,In_1986);
nor U7 (N_7,In_877,In_1300);
and U8 (N_8,In_1237,In_1396);
nor U9 (N_9,In_97,In_157);
xnor U10 (N_10,In_391,In_405);
xor U11 (N_11,In_250,In_382);
and U12 (N_12,In_959,In_418);
or U13 (N_13,In_213,In_1935);
or U14 (N_14,In_1874,In_1183);
xnor U15 (N_15,In_1005,In_758);
xor U16 (N_16,In_1859,In_200);
xor U17 (N_17,In_433,In_1565);
and U18 (N_18,In_617,In_1480);
xnor U19 (N_19,In_1971,In_1240);
nand U20 (N_20,In_605,In_156);
or U21 (N_21,In_839,In_152);
nor U22 (N_22,In_136,In_1852);
xnor U23 (N_23,In_1469,In_1764);
nand U24 (N_24,In_882,In_1766);
and U25 (N_25,In_1401,In_217);
xnor U26 (N_26,In_687,In_796);
and U27 (N_27,In_525,In_214);
and U28 (N_28,In_426,In_1673);
and U29 (N_29,In_1718,In_943);
nor U30 (N_30,In_122,In_380);
nor U31 (N_31,In_1280,In_1827);
or U32 (N_32,In_550,In_1387);
nor U33 (N_33,In_13,In_1890);
nor U34 (N_34,In_1832,In_1488);
and U35 (N_35,In_1729,In_1506);
or U36 (N_36,In_1624,In_1615);
or U37 (N_37,In_1957,In_823);
xor U38 (N_38,In_1574,In_423);
and U39 (N_39,In_1811,In_1163);
and U40 (N_40,In_932,In_743);
or U41 (N_41,In_303,In_1343);
nand U42 (N_42,In_917,In_1868);
nor U43 (N_43,In_72,In_20);
nand U44 (N_44,In_651,In_141);
nor U45 (N_45,In_7,In_507);
and U46 (N_46,In_689,In_1412);
nand U47 (N_47,In_1249,In_1558);
xor U48 (N_48,In_592,In_1323);
xnor U49 (N_49,In_1800,In_1638);
nor U50 (N_50,In_698,In_560);
xnor U51 (N_51,In_196,In_1593);
nor U52 (N_52,In_1353,In_1101);
or U53 (N_53,In_1499,In_276);
and U54 (N_54,In_1022,In_179);
nand U55 (N_55,In_1555,In_215);
or U56 (N_56,In_505,In_1862);
nand U57 (N_57,In_65,In_1326);
nor U58 (N_58,In_1011,In_1524);
and U59 (N_59,In_1568,In_103);
and U60 (N_60,In_623,In_814);
and U61 (N_61,In_767,In_1444);
and U62 (N_62,In_45,In_1683);
and U63 (N_63,In_1947,In_1846);
xnor U64 (N_64,In_580,In_1755);
nor U65 (N_65,In_1422,In_190);
xnor U66 (N_66,In_1225,In_1534);
xnor U67 (N_67,In_348,In_1503);
and U68 (N_68,In_1744,In_1067);
nand U69 (N_69,In_753,In_688);
nand U70 (N_70,In_569,In_1419);
nand U71 (N_71,In_311,In_519);
xnor U72 (N_72,In_1538,In_771);
nor U73 (N_73,In_696,In_585);
or U74 (N_74,In_1818,In_1404);
nor U75 (N_75,In_982,In_616);
xnor U76 (N_76,In_1308,In_610);
xor U77 (N_77,In_1675,In_778);
xnor U78 (N_78,In_1677,In_596);
nand U79 (N_79,In_869,In_1057);
or U80 (N_80,In_115,In_1625);
nand U81 (N_81,In_1620,In_1203);
nor U82 (N_82,In_1400,In_1315);
nor U83 (N_83,In_1247,In_455);
nand U84 (N_84,In_88,In_654);
nand U85 (N_85,In_1036,In_102);
and U86 (N_86,In_1934,In_544);
nor U87 (N_87,In_663,In_600);
xnor U88 (N_88,In_1951,In_1903);
xnor U89 (N_89,In_1206,In_1416);
nand U90 (N_90,In_735,In_304);
nand U91 (N_91,In_1687,In_1665);
nand U92 (N_92,In_1781,In_1445);
nor U93 (N_93,In_460,In_1093);
xor U94 (N_94,In_1543,In_1063);
and U95 (N_95,In_1960,In_960);
xor U96 (N_96,In_1805,In_759);
or U97 (N_97,In_449,In_318);
or U98 (N_98,In_642,In_360);
nor U99 (N_99,In_629,In_1429);
nor U100 (N_100,In_171,In_1569);
nand U101 (N_101,In_465,In_1398);
xor U102 (N_102,In_969,In_1342);
or U103 (N_103,In_637,In_697);
or U104 (N_104,In_1086,In_1804);
and U105 (N_105,In_1871,In_1000);
nand U106 (N_106,In_1532,In_1123);
xor U107 (N_107,In_189,In_992);
nand U108 (N_108,In_1196,In_524);
or U109 (N_109,In_515,In_664);
nand U110 (N_110,In_1201,In_227);
nor U111 (N_111,In_24,In_1495);
xnor U112 (N_112,In_1088,In_326);
nand U113 (N_113,In_85,In_1676);
or U114 (N_114,In_1334,In_1180);
and U115 (N_115,In_16,In_1984);
xnor U116 (N_116,In_1883,In_924);
xor U117 (N_117,In_257,In_602);
and U118 (N_118,In_1742,In_472);
or U119 (N_119,In_1454,In_1896);
nand U120 (N_120,In_96,In_1414);
or U121 (N_121,In_1390,In_1831);
or U122 (N_122,In_1710,In_568);
nor U123 (N_123,In_1816,In_1702);
nor U124 (N_124,In_716,In_952);
xor U125 (N_125,In_454,In_1750);
xor U126 (N_126,In_324,In_1113);
nand U127 (N_127,In_1441,In_1162);
xor U128 (N_128,In_191,In_22);
or U129 (N_129,In_691,In_1823);
nor U130 (N_130,In_1709,In_1245);
xnor U131 (N_131,In_618,In_973);
xor U132 (N_132,In_1104,In_135);
or U133 (N_133,In_1256,In_657);
nor U134 (N_134,In_1566,In_910);
nor U135 (N_135,In_206,In_599);
or U136 (N_136,In_1448,In_1160);
nor U137 (N_137,In_491,In_47);
xnor U138 (N_138,In_1255,In_784);
xnor U139 (N_139,In_720,In_949);
and U140 (N_140,In_1678,In_462);
xor U141 (N_141,In_708,In_723);
nor U142 (N_142,In_450,In_703);
nand U143 (N_143,In_1297,In_1187);
nor U144 (N_144,In_883,In_1777);
nand U145 (N_145,In_1937,In_6);
nand U146 (N_146,In_532,In_1640);
and U147 (N_147,In_1411,In_343);
xor U148 (N_148,In_1330,In_1092);
or U149 (N_149,In_417,In_939);
and U150 (N_150,In_1567,In_1803);
nand U151 (N_151,In_719,In_1784);
nand U152 (N_152,In_9,In_1873);
or U153 (N_153,In_1253,In_1318);
xor U154 (N_154,In_1779,In_1142);
and U155 (N_155,In_205,In_175);
or U156 (N_156,In_224,In_368);
xnor U157 (N_157,In_1878,In_369);
or U158 (N_158,In_1331,In_1027);
and U159 (N_159,In_1920,In_81);
xnor U160 (N_160,In_986,In_807);
or U161 (N_161,In_267,In_1476);
nand U162 (N_162,In_1577,In_1451);
nand U163 (N_163,In_17,In_764);
and U164 (N_164,In_1279,In_1660);
and U165 (N_165,In_1848,In_106);
and U166 (N_166,In_67,In_1587);
nor U167 (N_167,In_971,In_358);
nor U168 (N_168,In_1513,In_1529);
nand U169 (N_169,In_752,In_672);
and U170 (N_170,In_319,In_480);
nor U171 (N_171,In_306,In_1291);
or U172 (N_172,In_1371,In_641);
nor U173 (N_173,In_923,In_1303);
or U174 (N_174,In_1202,In_667);
nor U175 (N_175,In_1415,In_798);
and U176 (N_176,In_133,In_1970);
and U177 (N_177,In_1131,In_104);
xnor U178 (N_178,In_1186,In_1571);
or U179 (N_179,In_1712,In_105);
xnor U180 (N_180,In_1598,In_1156);
nor U181 (N_181,In_356,In_851);
xor U182 (N_182,In_363,In_1185);
xor U183 (N_183,In_808,In_576);
nor U184 (N_184,In_1599,In_389);
nor U185 (N_185,In_1737,In_1319);
xor U186 (N_186,In_1659,In_751);
nand U187 (N_187,In_1809,In_69);
nand U188 (N_188,In_1626,In_339);
nand U189 (N_189,In_328,In_1837);
xor U190 (N_190,In_1556,In_173);
and U191 (N_191,In_563,In_286);
or U192 (N_192,In_1273,In_1901);
nand U193 (N_193,In_1916,In_912);
nor U194 (N_194,In_979,In_1926);
or U195 (N_195,In_540,In_1305);
and U196 (N_196,In_8,In_1807);
and U197 (N_197,In_740,In_929);
and U198 (N_198,In_1796,In_577);
nand U199 (N_199,In_761,In_1149);
nor U200 (N_200,In_652,In_714);
nand U201 (N_201,In_1711,In_766);
and U202 (N_202,In_1606,In_1485);
nor U203 (N_203,In_11,In_1627);
nor U204 (N_204,In_1704,In_1374);
and U205 (N_205,In_1706,In_308);
xor U206 (N_206,In_290,In_464);
nand U207 (N_207,In_461,In_411);
xnor U208 (N_208,In_1719,In_590);
or U209 (N_209,In_1995,In_82);
nand U210 (N_210,In_1560,In_899);
xnor U211 (N_211,In_1126,In_564);
nor U212 (N_212,In_1211,In_158);
and U213 (N_213,In_296,In_1684);
nand U214 (N_214,In_1048,In_976);
and U215 (N_215,In_984,In_678);
nand U216 (N_216,In_1333,In_692);
nand U217 (N_217,In_1815,In_1337);
nand U218 (N_218,In_436,In_204);
and U219 (N_219,In_1136,In_1798);
and U220 (N_220,In_1952,In_167);
and U221 (N_221,In_791,In_1824);
and U222 (N_222,In_1214,In_1347);
and U223 (N_223,In_732,In_1685);
or U224 (N_224,In_333,In_1363);
nor U225 (N_225,In_188,In_941);
or U226 (N_226,In_867,In_1306);
xor U227 (N_227,In_1958,In_844);
and U228 (N_228,In_1325,In_1542);
nor U229 (N_229,In_1802,In_597);
and U230 (N_230,In_1295,In_134);
nand U231 (N_231,In_309,In_1872);
nor U232 (N_232,In_234,In_579);
nor U233 (N_233,In_1492,In_231);
and U234 (N_234,In_571,In_864);
or U235 (N_235,In_441,In_1288);
nor U236 (N_236,In_1435,In_1554);
nor U237 (N_237,In_1033,In_1754);
nor U238 (N_238,In_292,In_1046);
xnor U239 (N_239,In_340,In_1949);
xnor U240 (N_240,In_792,In_101);
and U241 (N_241,In_38,In_1270);
xor U242 (N_242,In_1413,In_1500);
nor U243 (N_243,In_876,In_422);
nand U244 (N_244,In_1405,In_542);
nand U245 (N_245,In_619,In_1658);
nand U246 (N_246,In_251,In_216);
or U247 (N_247,In_694,In_968);
nand U248 (N_248,In_146,In_1731);
xnor U249 (N_249,In_879,In_1924);
and U250 (N_250,In_481,In_1148);
nand U251 (N_251,In_230,In_1231);
or U252 (N_252,In_1917,In_1771);
and U253 (N_253,In_1228,In_1188);
xor U254 (N_254,In_742,In_1988);
or U255 (N_255,In_208,In_1084);
or U256 (N_256,In_1239,In_660);
nand U257 (N_257,In_1407,In_1431);
or U258 (N_258,In_377,In_859);
and U259 (N_259,In_1197,In_1586);
or U260 (N_260,In_355,In_1610);
or U261 (N_261,In_218,In_1474);
or U262 (N_262,In_140,In_457);
and U263 (N_263,In_1179,In_620);
nand U264 (N_264,In_896,In_384);
xnor U265 (N_265,In_1345,In_523);
and U266 (N_266,In_614,In_154);
xnor U267 (N_267,In_399,In_430);
nor U268 (N_268,In_1622,In_1498);
xor U269 (N_269,In_1623,In_484);
or U270 (N_270,In_647,In_1477);
or U271 (N_271,In_1030,In_1932);
or U272 (N_272,In_974,In_1207);
nand U273 (N_273,In_0,In_897);
and U274 (N_274,In_1521,In_1547);
nor U275 (N_275,In_565,In_955);
nand U276 (N_276,In_1009,In_359);
and U277 (N_277,In_888,In_1968);
or U278 (N_278,In_573,In_1320);
and U279 (N_279,In_1674,In_1286);
nor U280 (N_280,In_554,In_1355);
nor U281 (N_281,In_253,In_1468);
or U282 (N_282,In_852,In_1533);
xor U283 (N_283,In_1893,In_1362);
nor U284 (N_284,In_1695,In_32);
xnor U285 (N_285,In_375,In_337);
nand U286 (N_286,In_170,In_1793);
nand U287 (N_287,In_1551,In_827);
or U288 (N_288,In_1109,In_502);
or U289 (N_289,In_1631,In_349);
xor U290 (N_290,In_1941,In_1041);
or U291 (N_291,In_1613,In_1064);
nor U292 (N_292,In_279,In_1643);
or U293 (N_293,In_1921,In_172);
or U294 (N_294,In_62,In_780);
nor U295 (N_295,In_479,In_1655);
xnor U296 (N_296,In_1144,In_996);
and U297 (N_297,In_87,In_1434);
nor U298 (N_298,In_850,In_665);
xnor U299 (N_299,In_1649,In_983);
xor U300 (N_300,In_1739,In_420);
xor U301 (N_301,In_492,In_1950);
nand U302 (N_302,In_1298,In_1840);
nand U303 (N_303,In_834,In_1072);
xnor U304 (N_304,In_1130,In_1889);
xnor U305 (N_305,In_1176,In_1065);
nand U306 (N_306,In_1780,In_1894);
or U307 (N_307,In_829,In_1976);
nor U308 (N_308,In_736,In_1669);
and U309 (N_309,In_1034,In_1112);
xnor U310 (N_310,In_1020,In_1514);
nand U311 (N_311,In_643,In_159);
and U312 (N_312,In_1339,In_452);
or U313 (N_313,In_160,In_830);
nor U314 (N_314,In_1283,In_1437);
or U315 (N_315,In_1738,In_1508);
nor U316 (N_316,In_777,In_746);
or U317 (N_317,In_1996,In_832);
and U318 (N_318,In_1455,In_1356);
and U319 (N_319,In_89,In_1446);
nand U320 (N_320,In_1884,In_1511);
and U321 (N_321,In_1198,In_301);
xor U322 (N_322,In_111,In_887);
xnor U323 (N_323,In_421,In_1908);
xnor U324 (N_324,In_1962,In_769);
or U325 (N_325,In_265,In_578);
and U326 (N_326,In_693,In_329);
xnor U327 (N_327,In_506,In_1259);
xnor U328 (N_328,In_1735,In_1394);
nor U329 (N_329,In_1760,In_595);
nor U330 (N_330,In_621,In_843);
or U331 (N_331,In_682,In_645);
or U332 (N_332,In_497,In_946);
or U333 (N_333,In_169,In_1923);
or U334 (N_334,In_1668,In_717);
or U335 (N_335,In_608,In_275);
or U336 (N_336,In_627,In_1473);
xor U337 (N_337,In_486,In_1931);
nand U338 (N_338,In_1672,In_1489);
nor U339 (N_339,In_1461,In_1094);
and U340 (N_340,In_1467,In_226);
nor U341 (N_341,In_1043,In_1003);
xnor U342 (N_342,In_789,In_298);
xnor U343 (N_343,In_900,In_1799);
and U344 (N_344,In_1170,In_1375);
nor U345 (N_345,In_931,In_1154);
nand U346 (N_346,In_1458,In_671);
nor U347 (N_347,In_347,In_810);
nand U348 (N_348,In_1842,In_1716);
xor U349 (N_349,In_1369,In_1447);
nor U350 (N_350,In_750,In_95);
xor U351 (N_351,In_1209,In_315);
or U352 (N_352,In_30,In_601);
nand U353 (N_353,In_1867,In_1497);
and U354 (N_354,In_551,In_783);
nand U355 (N_355,In_1217,In_956);
or U356 (N_356,In_670,In_1096);
nand U357 (N_357,In_1794,In_29);
and U358 (N_358,In_1851,In_1652);
nand U359 (N_359,In_1481,In_593);
and U360 (N_360,In_50,In_1752);
or U361 (N_361,In_856,In_1050);
or U362 (N_362,In_533,In_799);
or U363 (N_363,In_634,In_1686);
nand U364 (N_364,In_28,In_395);
xor U365 (N_365,In_1153,In_1789);
nand U366 (N_366,In_366,In_1713);
xnor U367 (N_367,In_1292,In_414);
and U368 (N_368,In_1351,In_1733);
or U369 (N_369,In_287,In_1933);
xnor U370 (N_370,In_953,In_1397);
and U371 (N_371,In_1392,In_1026);
nor U372 (N_372,In_1496,In_1146);
nand U373 (N_373,In_53,In_1222);
xnor U374 (N_374,In_1863,In_40);
xnor U375 (N_375,In_555,In_1479);
xor U376 (N_376,In_730,In_1314);
or U377 (N_377,In_177,In_92);
nor U378 (N_378,In_1855,In_1159);
nor U379 (N_379,In_413,In_1083);
or U380 (N_380,In_197,In_155);
and U381 (N_381,In_1812,In_567);
or U382 (N_382,In_1376,In_517);
xor U383 (N_383,In_1531,In_1635);
nor U384 (N_384,In_1523,In_1352);
nand U385 (N_385,In_1858,In_302);
xor U386 (N_386,In_1462,In_1991);
xor U387 (N_387,In_1257,In_936);
and U388 (N_388,In_1930,In_680);
xor U389 (N_389,In_893,In_398);
nand U390 (N_390,In_557,In_142);
or U391 (N_391,In_396,In_1787);
nor U392 (N_392,In_1767,In_1205);
and U393 (N_393,In_966,In_198);
or U394 (N_394,In_675,In_763);
nor U395 (N_395,In_1282,In_1632);
nand U396 (N_396,In_1845,In_1681);
nor U397 (N_397,In_1002,In_1758);
nor U398 (N_398,In_453,In_1667);
xor U399 (N_399,In_1029,In_59);
nand U400 (N_400,In_415,In_1054);
and U401 (N_401,In_1783,In_1421);
xor U402 (N_402,In_1728,In_775);
xor U403 (N_403,In_451,In_335);
and U404 (N_404,In_1236,In_1472);
xnor U405 (N_405,In_727,In_646);
nand U406 (N_406,In_261,In_1466);
and U407 (N_407,In_818,In_1470);
nor U408 (N_408,In_71,In_779);
nor U409 (N_409,In_440,In_1108);
xnor U410 (N_410,In_1570,In_18);
nand U411 (N_411,In_1505,In_1490);
and U412 (N_412,In_1603,In_1417);
or U413 (N_413,In_1340,In_633);
nor U414 (N_414,In_531,In_1349);
and U415 (N_415,In_541,In_1723);
nand U416 (N_416,In_424,In_1129);
xnor U417 (N_417,In_1967,In_1990);
nand U418 (N_418,In_1328,In_636);
and U419 (N_419,In_1494,In_1060);
nand U420 (N_420,In_785,In_1382);
or U421 (N_421,In_937,In_1493);
xor U422 (N_422,In_121,In_184);
nand U423 (N_423,In_1220,In_1013);
and U424 (N_424,In_126,In_1510);
and U425 (N_425,In_1909,In_1992);
xor U426 (N_426,In_1006,In_988);
and U427 (N_427,In_1302,In_1945);
nand U428 (N_428,In_1252,In_794);
and U429 (N_429,In_1768,In_1575);
or U430 (N_430,In_285,In_1938);
xnor U431 (N_431,In_370,In_695);
nor U432 (N_432,In_1939,In_1810);
or U433 (N_433,In_781,In_1839);
xnor U434 (N_434,In_1634,In_556);
or U435 (N_435,In_473,In_1892);
and U436 (N_436,In_1482,In_288);
and U437 (N_437,In_733,In_958);
and U438 (N_438,In_351,In_1730);
nand U439 (N_439,In_371,In_903);
xnor U440 (N_440,In_760,In_222);
and U441 (N_441,In_1518,In_1090);
nor U442 (N_442,In_98,In_1790);
nand U443 (N_443,In_1311,In_12);
xnor U444 (N_444,In_786,In_1055);
nor U445 (N_445,In_1963,In_817);
and U446 (N_446,In_1776,In_1004);
xor U447 (N_447,In_1747,In_271);
or U448 (N_448,In_330,In_1483);
xnor U449 (N_449,In_1053,In_247);
or U450 (N_450,In_1132,In_1426);
xnor U451 (N_451,In_625,In_622);
or U452 (N_452,In_1221,In_1119);
nor U453 (N_453,In_707,In_131);
xor U454 (N_454,In_868,In_1385);
and U455 (N_455,In_442,In_1501);
nand U456 (N_456,In_857,In_768);
nand U457 (N_457,In_1701,In_416);
or U458 (N_458,In_1386,In_1830);
or U459 (N_459,In_1875,In_1853);
nor U460 (N_460,In_865,In_863);
nand U461 (N_461,In_1955,In_1487);
nand U462 (N_462,In_1049,In_1251);
nor U463 (N_463,In_933,In_1689);
or U464 (N_464,In_1350,In_683);
nor U465 (N_465,In_99,In_161);
or U466 (N_466,In_1456,In_930);
xor U467 (N_467,In_725,In_401);
and U468 (N_468,In_1087,In_1998);
or U469 (N_469,In_1114,In_1143);
and U470 (N_470,In_1595,In_997);
and U471 (N_471,In_125,In_1307);
xor U472 (N_472,In_991,In_242);
nand U473 (N_473,In_361,In_1745);
and U474 (N_474,In_4,In_90);
and U475 (N_475,In_467,In_787);
nor U476 (N_476,In_1707,In_164);
and U477 (N_477,In_635,In_378);
xnor U478 (N_478,In_561,In_1443);
nand U479 (N_479,In_1007,In_1765);
nand U480 (N_480,In_545,In_1366);
nand U481 (N_481,In_1233,In_1001);
or U482 (N_482,In_1227,In_1527);
xor U483 (N_483,In_1381,In_244);
or U484 (N_484,In_1696,In_1014);
and U485 (N_485,In_1212,In_987);
or U486 (N_486,In_112,In_1268);
or U487 (N_487,In_352,In_640);
nand U488 (N_488,In_738,In_980);
nor U489 (N_489,In_54,In_1912);
nor U490 (N_490,In_1942,In_1721);
nand U491 (N_491,In_58,In_1261);
and U492 (N_492,In_435,In_236);
or U493 (N_493,In_448,In_1038);
xnor U494 (N_494,In_1389,In_243);
and U495 (N_495,In_1365,In_901);
or U496 (N_496,In_954,In_566);
or U497 (N_497,In_1618,In_1509);
and U498 (N_498,In_1975,In_537);
or U499 (N_499,In_1699,In_195);
xnor U500 (N_500,In_344,In_1817);
nand U501 (N_501,In_1124,In_1418);
or U502 (N_502,In_386,In_1042);
and U503 (N_503,In_1700,In_1103);
xnor U504 (N_504,In_284,In_661);
nand U505 (N_505,In_521,In_649);
xnor U506 (N_506,In_336,In_1486);
nand U507 (N_507,In_612,In_393);
or U508 (N_508,In_278,In_892);
xor U509 (N_509,In_1128,In_365);
nor U510 (N_510,In_1321,In_1023);
nand U511 (N_511,In_475,In_1377);
xor U512 (N_512,In_1010,In_341);
nand U513 (N_513,In_848,In_1244);
and U514 (N_514,In_1152,In_1232);
nand U515 (N_515,In_130,In_407);
nand U516 (N_516,In_1174,In_731);
xor U517 (N_517,In_1044,In_489);
nor U518 (N_518,In_659,In_1994);
nand U519 (N_519,In_1993,In_842);
and U520 (N_520,In_1338,In_229);
or U521 (N_521,In_588,In_379);
xnor U522 (N_522,In_1727,In_999);
or U523 (N_523,In_1138,In_520);
or U524 (N_524,In_1062,In_1692);
xor U525 (N_525,In_1985,In_989);
or U526 (N_526,In_1539,In_724);
and U527 (N_527,In_885,In_711);
and U528 (N_528,In_412,In_166);
or U529 (N_529,In_262,In_34);
nor U530 (N_530,In_1047,In_207);
xor U531 (N_531,In_438,In_1165);
nand U532 (N_532,In_314,In_120);
and U533 (N_533,In_36,In_1019);
nor U534 (N_534,In_354,In_718);
nor U535 (N_535,In_662,In_252);
xor U536 (N_536,In_765,In_840);
or U537 (N_537,In_1682,In_403);
nand U538 (N_538,In_1639,In_1774);
nor U539 (N_539,In_891,In_1059);
nor U540 (N_540,In_993,In_273);
nand U541 (N_541,In_35,In_1806);
nand U542 (N_542,In_404,In_1161);
nor U543 (N_543,In_1761,In_770);
xnor U544 (N_544,In_1698,In_232);
and U545 (N_545,In_446,In_589);
nand U546 (N_546,In_1066,In_1145);
or U547 (N_547,In_1726,In_239);
nor U548 (N_548,In_1905,In_835);
and U549 (N_549,In_562,In_632);
nand U550 (N_550,In_168,In_1465);
nor U551 (N_551,In_1753,In_1579);
nand U552 (N_552,In_1559,In_926);
or U553 (N_553,In_237,In_797);
xnor U554 (N_554,In_1697,In_655);
xor U555 (N_555,In_1825,In_1645);
xnor U556 (N_556,In_726,In_1576);
nand U557 (N_557,In_1287,In_638);
or U558 (N_558,In_1238,In_1275);
or U559 (N_559,In_1778,In_1797);
or U560 (N_560,In_107,In_1572);
or U561 (N_561,In_26,In_1866);
and U562 (N_562,In_332,In_1316);
xor U563 (N_563,In_944,In_291);
nand U564 (N_564,In_1982,In_1722);
or U565 (N_565,In_263,In_447);
xnor U566 (N_566,In_1974,In_1502);
xor U567 (N_567,In_1324,In_1861);
nand U568 (N_568,In_1208,In_928);
nand U569 (N_569,In_1134,In_345);
and U570 (N_570,In_950,In_866);
or U571 (N_571,In_1978,In_1040);
or U572 (N_572,In_437,In_1581);
nor U573 (N_573,In_439,In_474);
nor U574 (N_574,In_1121,In_254);
xnor U575 (N_575,In_1313,In_128);
and U576 (N_576,In_1749,In_1267);
nor U577 (N_577,In_774,In_1304);
nand U578 (N_578,In_700,In_1822);
xor U579 (N_579,In_282,In_10);
nor U580 (N_580,In_1433,In_63);
xor U581 (N_581,In_591,In_1078);
or U582 (N_582,In_630,In_826);
and U583 (N_583,In_849,In_1956);
nand U584 (N_584,In_1368,In_1317);
xnor U585 (N_585,In_1388,In_1155);
and U586 (N_586,In_940,In_108);
and U587 (N_587,In_19,In_1182);
xor U588 (N_588,In_1881,In_1786);
nand U589 (N_589,In_755,In_1943);
and U590 (N_590,In_431,In_1666);
or U591 (N_591,In_913,In_1791);
and U592 (N_592,In_1589,In_219);
nor U593 (N_593,In_704,In_653);
or U594 (N_594,In_1061,In_203);
nor U595 (N_595,In_737,In_1705);
nand U596 (N_596,In_1929,In_425);
xnor U597 (N_597,In_1169,In_747);
nand U598 (N_598,In_93,In_1585);
xnor U599 (N_599,In_1600,In_1516);
nand U600 (N_600,In_174,In_1423);
nand U601 (N_601,In_1106,In_1269);
and U602 (N_602,In_1834,In_1463);
nand U603 (N_603,In_853,In_220);
nand U604 (N_604,In_788,In_1637);
xnor U605 (N_605,In_1367,In_176);
and U606 (N_606,In_2,In_880);
or U607 (N_607,In_1348,In_598);
or U608 (N_608,In_1897,In_1139);
nor U609 (N_609,In_990,In_685);
nand U610 (N_610,In_961,In_806);
or U611 (N_611,In_482,In_1910);
and U612 (N_612,In_1464,In_644);
or U613 (N_613,In_1869,In_772);
nand U614 (N_614,In_1904,In_1720);
xor U615 (N_615,In_48,In_186);
nand U616 (N_616,In_165,In_1032);
or U617 (N_617,In_739,In_478);
nor U618 (N_618,In_249,In_1122);
nand U619 (N_619,In_970,In_1335);
or U620 (N_620,In_1946,In_124);
and U621 (N_621,In_916,In_527);
xnor U622 (N_622,In_898,In_539);
nor U623 (N_623,In_1336,In_1953);
xnor U624 (N_624,In_1460,In_1299);
and U625 (N_625,In_1741,In_1919);
xor U626 (N_626,In_44,In_1184);
nand U627 (N_627,In_513,In_570);
and U628 (N_628,In_1117,In_534);
nand U629 (N_629,In_1070,In_925);
or U630 (N_630,In_824,In_295);
nand U631 (N_631,In_803,In_1242);
or U632 (N_632,In_225,In_1216);
and U633 (N_633,In_1332,In_221);
nor U634 (N_634,In_3,In_677);
nand U635 (N_635,In_1424,In_83);
xor U636 (N_636,In_193,In_1150);
nand U637 (N_637,In_488,In_1230);
or U638 (N_638,In_350,In_813);
nor U639 (N_639,In_918,In_1792);
nor U640 (N_640,In_1262,In_151);
or U641 (N_641,In_606,In_185);
or U642 (N_642,In_428,In_1195);
or U643 (N_643,In_1105,In_658);
or U644 (N_644,In_374,In_313);
nor U645 (N_645,In_1549,In_86);
or U646 (N_646,In_201,In_55);
xnor U647 (N_647,In_1715,In_495);
or U648 (N_648,In_631,In_582);
or U649 (N_649,In_1512,In_1641);
or U650 (N_650,In_1849,In_1954);
nand U651 (N_651,In_364,In_1588);
or U652 (N_652,In_907,In_1223);
nor U653 (N_653,In_1164,In_801);
and U654 (N_654,In_1724,In_429);
xnor U655 (N_655,In_114,In_1911);
and U656 (N_656,In_468,In_5);
xor U657 (N_657,In_1192,In_1346);
nor U658 (N_658,In_1821,In_1012);
or U659 (N_659,In_100,In_1944);
xnor U660 (N_660,In_1194,In_1880);
and U661 (N_661,In_1080,In_182);
and U662 (N_662,In_307,In_80);
nor U663 (N_663,In_322,In_1116);
nor U664 (N_664,In_594,In_15);
or U665 (N_665,In_855,In_1769);
or U666 (N_666,In_270,In_745);
or U667 (N_667,In_1838,In_317);
or U668 (N_668,In_927,In_1535);
or U669 (N_669,In_705,In_884);
nor U670 (N_670,In_1879,In_470);
nor U671 (N_671,In_1151,In_861);
nand U672 (N_672,In_1248,In_320);
nand U673 (N_673,In_1289,In_1999);
nand U674 (N_674,In_1359,In_1408);
xor U675 (N_675,In_409,In_1210);
and U676 (N_676,In_744,In_406);
or U677 (N_677,In_748,In_297);
nand U678 (N_678,In_500,In_1409);
or U679 (N_679,In_42,In_699);
xnor U680 (N_680,In_904,In_1969);
nor U681 (N_681,In_833,In_109);
and U682 (N_682,In_1907,In_1679);
nand U683 (N_683,In_639,In_181);
or U684 (N_684,In_1406,In_1358);
nand U685 (N_685,In_1621,In_362);
xor U686 (N_686,In_972,In_240);
and U687 (N_687,In_650,In_1378);
nand U688 (N_688,In_183,In_514);
or U689 (N_689,In_825,In_228);
nand U690 (N_690,In_1076,In_1137);
nor U691 (N_691,In_624,In_1085);
and U692 (N_692,In_310,In_858);
nand U693 (N_693,In_1656,In_1616);
and U694 (N_694,In_199,In_1438);
nand U695 (N_695,In_400,In_1876);
nor U696 (N_696,In_76,In_776);
or U697 (N_697,In_1762,In_819);
nand U698 (N_698,In_1854,In_1383);
xor U699 (N_699,In_269,In_1329);
nand U700 (N_700,In_1959,In_1052);
nand U701 (N_701,In_79,In_690);
nor U702 (N_702,In_1813,In_1828);
nor U703 (N_703,In_1788,In_1561);
or U704 (N_704,In_212,In_1016);
or U705 (N_705,In_1141,In_1265);
nor U706 (N_706,In_1918,In_994);
nand U707 (N_707,In_1384,In_1536);
nand U708 (N_708,In_1922,In_469);
xnor U709 (N_709,In_511,In_153);
nand U710 (N_710,In_1399,In_1364);
xor U711 (N_711,In_376,In_70);
nand U712 (N_712,In_526,In_1120);
xnor U713 (N_713,In_1987,In_1650);
and U714 (N_714,In_1814,In_162);
and U715 (N_715,In_129,In_485);
nand U716 (N_716,In_518,In_1847);
xor U717 (N_717,In_493,In_558);
nand U718 (N_718,In_1293,In_1900);
xor U719 (N_719,In_61,In_1177);
xor U720 (N_720,In_1189,In_1484);
nand U721 (N_721,In_615,In_1642);
xnor U722 (N_722,In_503,In_316);
or U723 (N_723,In_712,In_1074);
nand U724 (N_724,In_274,In_1051);
nor U725 (N_725,In_552,In_1081);
xor U726 (N_726,In_729,In_1100);
nand U727 (N_727,In_1617,In_110);
nand U728 (N_728,In_1258,In_1099);
or U729 (N_729,In_1979,In_1850);
nor U730 (N_730,In_1562,In_1564);
xor U731 (N_731,In_1902,In_1602);
nor U732 (N_732,In_535,In_1018);
and U733 (N_733,In_804,In_1361);
nand U734 (N_734,In_862,In_701);
nand U735 (N_735,In_1770,In_1671);
nor U736 (N_736,In_1629,In_145);
or U737 (N_737,In_408,In_1591);
xnor U738 (N_738,In_873,In_1661);
or U739 (N_739,In_1190,In_1925);
nor U740 (N_740,In_805,In_1775);
xnor U741 (N_741,In_1578,In_46);
nand U742 (N_742,In_1173,In_1243);
nand U743 (N_743,In_1819,In_458);
or U744 (N_744,In_846,In_1436);
nor U745 (N_745,In_1427,In_902);
and U746 (N_746,In_1546,In_938);
xor U747 (N_747,In_1964,In_1235);
xor U748 (N_748,In_1580,In_66);
nor U749 (N_749,In_1147,In_1037);
xnor U750 (N_750,In_1452,In_1940);
nor U751 (N_751,In_113,In_1633);
or U752 (N_752,In_860,In_800);
or U753 (N_753,In_1795,In_210);
xnor U754 (N_754,In_367,In_945);
or U755 (N_755,In_1605,In_211);
nand U756 (N_756,In_1420,In_1517);
and U757 (N_757,In_1111,In_1457);
nor U758 (N_758,In_385,In_39);
nor U759 (N_759,In_1545,In_668);
nor U760 (N_760,In_575,In_836);
and U761 (N_761,In_1557,In_1301);
nand U762 (N_762,In_676,In_1746);
xor U763 (N_763,In_1928,In_1608);
nor U764 (N_764,In_878,In_1276);
nor U765 (N_765,In_529,In_272);
nand U766 (N_766,In_975,In_456);
xor U767 (N_767,In_1835,In_1844);
nor U768 (N_768,In_78,In_871);
nand U769 (N_769,In_444,In_1354);
nor U770 (N_770,In_790,In_419);
nand U771 (N_771,In_1224,In_14);
or U772 (N_772,In_1888,In_1653);
or U773 (N_773,In_1860,In_1663);
or U774 (N_774,In_911,In_962);
nand U775 (N_775,In_1972,In_1541);
and U776 (N_776,In_1133,In_530);
or U777 (N_777,In_381,In_1260);
xor U778 (N_778,In_1757,In_1773);
or U779 (N_779,In_981,In_281);
nand U780 (N_780,In_60,In_1703);
nand U781 (N_781,In_266,In_1218);
nor U782 (N_782,In_1073,In_1264);
nor U783 (N_783,In_1344,In_387);
and U784 (N_784,In_1596,In_1604);
or U785 (N_785,In_559,In_1690);
and U786 (N_786,In_150,In_1552);
nor U787 (N_787,In_721,In_1648);
or U788 (N_788,In_728,In_1841);
xor U789 (N_789,In_1763,In_1548);
and U790 (N_790,In_119,In_209);
and U791 (N_791,In_1583,In_872);
xnor U792 (N_792,In_1507,In_289);
and U793 (N_793,In_1736,In_132);
or U794 (N_794,In_870,In_163);
nor U795 (N_795,In_1285,In_1887);
xor U796 (N_796,In_756,In_1274);
and U797 (N_797,In_68,In_1039);
and U798 (N_798,In_607,In_27);
and U799 (N_799,In_1607,In_1597);
xor U800 (N_800,In_1157,N_595);
nand U801 (N_801,N_744,N_355);
xor U802 (N_802,In_264,N_256);
nand U803 (N_803,In_192,N_771);
xnor U804 (N_804,N_180,In_77);
and U805 (N_805,N_456,N_659);
xnor U806 (N_806,N_725,N_275);
nor U807 (N_807,N_208,In_73);
nor U808 (N_808,N_214,N_67);
or U809 (N_809,In_41,In_1743);
nor U810 (N_810,N_370,N_110);
or U811 (N_811,N_40,N_547);
xor U812 (N_812,N_391,In_1717);
nand U813 (N_813,In_1836,N_198);
nor U814 (N_814,N_70,N_592);
xnor U815 (N_815,In_1058,N_133);
or U816 (N_816,In_43,In_1290);
xnor U817 (N_817,N_346,N_269);
xnor U818 (N_818,N_21,N_295);
xnor U819 (N_819,In_1540,N_611);
and U820 (N_820,In_459,In_1654);
or U821 (N_821,In_327,In_1725);
or U822 (N_822,N_336,In_21);
or U823 (N_823,N_340,N_93);
nor U824 (N_824,In_1662,N_733);
nor U825 (N_825,In_321,In_1520);
and U826 (N_826,In_434,In_1594);
nor U827 (N_827,N_378,N_749);
or U828 (N_828,N_85,In_845);
nor U829 (N_829,N_278,In_1425);
xnor U830 (N_830,N_743,In_1172);
or U831 (N_831,N_219,N_712);
nand U832 (N_832,N_577,In_1450);
nand U833 (N_833,N_294,In_300);
or U834 (N_834,N_151,N_35);
xnor U835 (N_835,N_588,N_648);
nor U836 (N_836,N_361,N_663);
or U837 (N_837,N_349,N_624);
nand U838 (N_838,In_1158,N_292);
nor U839 (N_839,N_508,N_538);
and U840 (N_840,N_128,N_548);
and U841 (N_841,N_0,N_350);
nand U842 (N_842,N_96,In_1936);
xor U843 (N_843,In_957,N_480);
or U844 (N_844,N_37,N_652);
nor U845 (N_845,In_1573,N_451);
xor U846 (N_846,In_669,In_536);
and U847 (N_847,N_258,In_1281);
or U848 (N_848,N_728,N_715);
or U849 (N_849,N_625,N_750);
or U850 (N_850,In_241,In_383);
nor U851 (N_851,N_50,In_886);
xnor U852 (N_852,In_443,N_684);
xor U853 (N_853,In_233,N_754);
nand U854 (N_854,In_1544,N_656);
and U855 (N_855,N_136,N_57);
and U856 (N_856,N_621,N_720);
xnor U857 (N_857,In_1504,N_542);
and U858 (N_858,N_513,In_1045);
and U859 (N_859,N_170,N_518);
nor U860 (N_860,In_1895,N_384);
nor U861 (N_861,In_1973,N_245);
xor U862 (N_862,N_468,In_656);
or U863 (N_863,N_443,N_783);
nand U864 (N_864,N_407,N_182);
nand U865 (N_865,In_1647,N_432);
and U866 (N_866,In_466,N_168);
or U867 (N_867,N_490,N_41);
or U868 (N_868,N_619,In_1782);
and U869 (N_869,N_660,N_319);
and U870 (N_870,N_446,N_273);
or U871 (N_871,N_34,N_778);
and U872 (N_872,In_762,N_109);
nand U873 (N_873,N_234,N_306);
xor U874 (N_874,In_666,N_729);
and U875 (N_875,N_314,N_97);
and U876 (N_876,N_790,N_132);
nand U877 (N_877,In_915,N_47);
or U878 (N_878,In_238,N_647);
or U879 (N_879,N_487,N_147);
nor U880 (N_880,N_390,In_1609);
nand U881 (N_881,N_442,In_802);
nand U882 (N_882,N_463,N_495);
nor U883 (N_883,N_516,N_484);
nand U884 (N_884,N_669,In_1178);
or U885 (N_885,N_531,N_260);
or U886 (N_886,In_246,N_575);
xnor U887 (N_887,N_427,In_1219);
xor U888 (N_888,N_231,In_749);
or U889 (N_889,In_710,In_1168);
or U890 (N_890,N_604,N_543);
and U891 (N_891,In_1175,In_626);
or U892 (N_892,N_488,N_503);
nor U893 (N_893,In_1614,N_158);
and U894 (N_894,N_679,In_722);
nor U895 (N_895,In_1948,N_765);
xnor U896 (N_896,In_1199,In_299);
or U897 (N_897,N_287,In_1772);
nor U898 (N_898,N_82,In_782);
nand U899 (N_899,In_1478,In_1089);
or U900 (N_900,N_546,N_402);
xnor U901 (N_901,N_244,N_581);
or U902 (N_902,In_854,N_724);
or U903 (N_903,N_593,In_342);
and U904 (N_904,N_166,N_413);
nand U905 (N_905,In_1864,N_140);
nand U906 (N_906,N_458,In_609);
nand U907 (N_907,N_429,In_334);
nor U908 (N_908,N_742,In_504);
nor U909 (N_909,N_60,N_524);
or U910 (N_910,N_134,N_63);
and U911 (N_911,In_483,N_731);
or U912 (N_912,In_934,In_144);
xor U913 (N_913,N_573,N_686);
xor U914 (N_914,In_679,In_1537);
nand U915 (N_915,N_795,In_543);
nor U916 (N_916,N_130,N_551);
and U917 (N_917,N_223,In_1530);
nor U918 (N_918,In_510,N_562);
xnor U919 (N_919,In_978,N_641);
nand U920 (N_920,N_83,N_525);
or U921 (N_921,N_172,N_31);
xnor U922 (N_922,N_552,N_455);
nor U923 (N_923,In_1296,N_98);
nand U924 (N_924,N_101,In_1865);
nor U925 (N_925,In_838,In_223);
and U926 (N_926,N_603,N_33);
nand U927 (N_927,N_86,N_705);
and U928 (N_928,N_123,N_474);
nor U929 (N_929,In_1171,N_261);
nor U930 (N_930,N_8,N_325);
nor U931 (N_931,In_967,N_745);
xnor U932 (N_932,N_175,In_1430);
nand U933 (N_933,In_947,In_889);
xor U934 (N_934,N_78,N_544);
xor U935 (N_935,N_354,N_666);
nor U936 (N_936,N_334,N_420);
and U937 (N_937,N_233,In_1740);
nand U938 (N_938,N_788,In_1628);
xnor U939 (N_939,N_775,In_353);
and U940 (N_940,N_87,N_760);
or U941 (N_941,In_1528,In_116);
or U942 (N_942,N_300,N_107);
and U943 (N_943,N_30,N_117);
or U944 (N_944,N_554,N_126);
nor U945 (N_945,N_371,N_363);
nand U946 (N_946,N_122,N_191);
or U947 (N_947,N_194,N_321);
xnor U948 (N_948,N_138,N_173);
nor U949 (N_949,In_1263,N_397);
xnor U950 (N_950,N_557,N_382);
xnor U951 (N_951,N_36,In_628);
nor U952 (N_952,N_475,N_17);
or U953 (N_953,N_598,N_764);
xnor U954 (N_954,N_145,N_752);
xor U955 (N_955,N_307,In_1732);
nor U956 (N_956,N_630,In_245);
nand U957 (N_957,N_64,N_367);
or U958 (N_958,N_673,N_496);
and U959 (N_959,N_634,N_165);
xor U960 (N_960,In_1630,N_448);
nor U961 (N_961,N_61,In_1357);
xnor U962 (N_962,N_520,In_1127);
or U963 (N_963,In_572,N_661);
nand U964 (N_964,N_746,N_4);
and U965 (N_965,N_44,In_1590);
or U966 (N_966,In_965,In_1310);
nor U967 (N_967,In_586,N_206);
xor U968 (N_968,In_325,N_365);
and U969 (N_969,N_710,In_522);
or U970 (N_970,N_787,In_1250);
nor U971 (N_971,In_1611,In_323);
and U972 (N_972,N_709,N_436);
nor U973 (N_973,In_1075,N_246);
or U974 (N_974,In_684,N_687);
xor U975 (N_975,In_1898,In_1024);
or U976 (N_976,N_84,N_254);
nand U977 (N_977,N_376,In_890);
xor U978 (N_978,In_906,N_626);
and U979 (N_979,In_445,N_736);
nand U980 (N_980,In_1395,N_609);
and U981 (N_981,In_394,N_302);
and U982 (N_982,N_711,N_237);
xor U983 (N_983,N_777,In_1379);
xnor U984 (N_984,N_276,N_576);
nand U985 (N_985,N_309,N_671);
nand U986 (N_986,N_755,N_617);
or U987 (N_987,N_615,N_250);
nand U988 (N_988,In_248,N_797);
nor U989 (N_989,N_42,In_392);
nor U990 (N_990,N_209,N_331);
or U991 (N_991,In_1181,In_948);
nor U992 (N_992,N_235,In_1636);
xnor U993 (N_993,In_235,In_1082);
and U994 (N_994,In_812,N_58);
nor U995 (N_995,In_1965,N_270);
nand U996 (N_996,N_568,In_1241);
or U997 (N_997,In_508,N_396);
xnor U998 (N_998,In_37,In_331);
and U999 (N_999,N_649,N_449);
and U1000 (N_1000,N_618,N_399);
or U1001 (N_1001,In_1071,N_221);
nand U1002 (N_1002,In_581,In_1294);
xnor U1003 (N_1003,N_32,N_774);
or U1004 (N_1004,N_483,In_516);
nor U1005 (N_1005,N_784,In_1584);
xnor U1006 (N_1006,N_640,N_763);
nand U1007 (N_1007,N_181,N_789);
and U1008 (N_1008,N_620,N_698);
nand U1009 (N_1009,N_457,N_105);
xnor U1010 (N_1010,In_1563,In_1226);
and U1011 (N_1011,N_515,N_124);
nor U1012 (N_1012,In_603,N_434);
or U1013 (N_1013,N_338,N_594);
nor U1014 (N_1014,N_741,In_33);
nand U1015 (N_1015,N_726,N_322);
or U1016 (N_1016,N_7,N_418);
or U1017 (N_1017,N_111,In_1229);
and U1018 (N_1018,N_737,N_424);
xor U1019 (N_1019,N_121,In_793);
nor U1020 (N_1020,In_681,N_556);
or U1021 (N_1021,In_490,N_230);
xor U1022 (N_1022,N_584,In_1035);
and U1023 (N_1023,N_676,N_257);
and U1024 (N_1024,N_668,N_591);
xnor U1025 (N_1025,In_1440,N_131);
xor U1026 (N_1026,In_1166,In_706);
nor U1027 (N_1027,N_500,N_757);
xor U1028 (N_1028,In_256,In_1857);
nand U1029 (N_1029,N_348,N_433);
nand U1030 (N_1030,In_1651,N_464);
nor U1031 (N_1031,In_56,In_674);
nor U1032 (N_1032,N_185,In_1442);
nand U1033 (N_1033,In_1785,N_430);
xor U1034 (N_1034,In_1471,N_716);
or U1035 (N_1035,N_772,N_431);
and U1036 (N_1036,N_727,N_517);
and U1037 (N_1037,N_414,In_1886);
and U1038 (N_1038,N_342,N_441);
xor U1039 (N_1039,In_1961,N_71);
and U1040 (N_1040,N_723,N_739);
xor U1041 (N_1041,N_466,N_578);
nand U1042 (N_1042,N_706,N_312);
or U1043 (N_1043,In_1360,In_1031);
nor U1044 (N_1044,In_734,N_425);
nand U1045 (N_1045,In_809,N_232);
and U1046 (N_1046,N_150,N_310);
nor U1047 (N_1047,N_639,N_318);
nor U1048 (N_1048,N_606,N_685);
xnor U1049 (N_1049,In_648,N_196);
xor U1050 (N_1050,N_69,N_357);
nand U1051 (N_1051,In_757,N_422);
nor U1052 (N_1052,In_1284,N_445);
nor U1053 (N_1053,N_732,N_279);
xor U1054 (N_1054,N_26,N_601);
or U1055 (N_1055,In_1515,In_1997);
and U1056 (N_1056,N_154,N_608);
xor U1057 (N_1057,N_19,N_259);
xor U1058 (N_1058,N_296,N_220);
and U1059 (N_1059,In_1914,N_329);
nor U1060 (N_1060,N_437,In_427);
nor U1061 (N_1061,In_1102,In_1519);
nand U1062 (N_1062,N_199,N_146);
or U1063 (N_1063,In_1734,N_493);
xnor U1064 (N_1064,N_226,N_670);
xnor U1065 (N_1065,N_127,In_1693);
and U1066 (N_1066,N_758,N_143);
nand U1067 (N_1067,N_574,In_1135);
xnor U1068 (N_1068,N_388,N_74);
nand U1069 (N_1069,N_459,N_409);
and U1070 (N_1070,In_604,N_633);
nor U1071 (N_1071,In_1826,N_205);
xor U1072 (N_1072,In_1309,In_149);
nand U1073 (N_1073,In_75,N_323);
and U1074 (N_1074,In_1592,In_538);
nand U1075 (N_1075,N_247,N_561);
and U1076 (N_1076,In_964,N_192);
or U1077 (N_1077,N_103,N_360);
nor U1078 (N_1078,In_1980,N_665);
or U1079 (N_1079,N_730,N_532);
and U1080 (N_1080,N_635,N_65);
and U1081 (N_1081,N_162,N_629);
xnor U1082 (N_1082,N_189,N_2);
xnor U1083 (N_1083,In_471,N_560);
or U1084 (N_1084,N_406,N_766);
and U1085 (N_1085,In_1432,N_20);
nand U1086 (N_1086,N_650,N_682);
nand U1087 (N_1087,N_528,In_118);
or U1088 (N_1088,N_693,N_571);
and U1089 (N_1089,N_423,N_389);
nand U1090 (N_1090,In_1808,N_597);
xnor U1091 (N_1091,N_80,N_529);
nor U1092 (N_1092,N_225,N_505);
and U1093 (N_1093,In_1167,In_138);
xnor U1094 (N_1094,N_337,N_438);
and U1095 (N_1095,N_510,N_535);
nand U1096 (N_1096,N_489,N_211);
or U1097 (N_1097,N_697,In_1272);
xor U1098 (N_1098,N_672,N_216);
nand U1099 (N_1099,In_1553,N_317);
nor U1100 (N_1100,N_401,N_638);
xor U1101 (N_1101,N_49,N_79);
xor U1102 (N_1102,N_527,N_22);
or U1103 (N_1103,N_335,N_10);
nand U1104 (N_1104,In_1246,In_998);
nand U1105 (N_1105,N_627,In_23);
and U1106 (N_1106,N_285,N_13);
or U1107 (N_1107,N_286,N_703);
or U1108 (N_1108,In_1234,N_303);
nand U1109 (N_1109,N_66,N_102);
nand U1110 (N_1110,N_164,N_631);
nor U1111 (N_1111,N_73,N_379);
and U1112 (N_1112,In_498,In_1644);
and U1113 (N_1113,In_549,In_1525);
or U1114 (N_1114,N_264,N_118);
xor U1115 (N_1115,N_613,In_1915);
nand U1116 (N_1116,In_895,N_253);
or U1117 (N_1117,In_1278,N_512);
nor U1118 (N_1118,In_894,In_258);
or U1119 (N_1119,N_228,N_761);
nand U1120 (N_1120,N_696,In_942);
xnor U1121 (N_1121,N_347,N_252);
and U1122 (N_1122,N_550,In_881);
xor U1123 (N_1123,In_1410,N_91);
nand U1124 (N_1124,N_115,In_1380);
xor U1125 (N_1125,In_1906,In_180);
or U1126 (N_1126,N_100,In_1820);
nor U1127 (N_1127,N_700,N_161);
xnor U1128 (N_1128,N_453,N_229);
nor U1129 (N_1129,N_6,N_653);
xnor U1130 (N_1130,In_1191,In_283);
xor U1131 (N_1131,N_572,N_171);
xnor U1132 (N_1132,N_89,In_187);
xor U1133 (N_1133,N_714,N_215);
nor U1134 (N_1134,N_51,N_526);
nand U1135 (N_1135,N_461,In_1322);
nor U1136 (N_1136,N_770,N_677);
and U1137 (N_1137,N_267,In_31);
nand U1138 (N_1138,In_875,In_52);
xnor U1139 (N_1139,N_28,N_202);
nor U1140 (N_1140,In_837,N_112);
nand U1141 (N_1141,N_600,N_636);
xor U1142 (N_1142,N_263,N_472);
nor U1143 (N_1143,N_55,N_227);
or U1144 (N_1144,N_266,In_1107);
nor U1145 (N_1145,N_190,N_667);
and U1146 (N_1146,In_1582,N_564);
nor U1147 (N_1147,In_1691,N_582);
nand U1148 (N_1148,In_1056,In_1843);
nor U1149 (N_1149,N_343,N_265);
and U1150 (N_1150,N_454,In_202);
xnor U1151 (N_1151,N_794,N_203);
xor U1152 (N_1152,In_259,In_1439);
nor U1153 (N_1153,N_486,In_1204);
nor U1154 (N_1154,N_522,N_341);
nand U1155 (N_1155,N_569,N_169);
nor U1156 (N_1156,N_756,In_1271);
and U1157 (N_1157,N_288,In_1312);
and U1158 (N_1158,N_694,N_632);
nor U1159 (N_1159,N_460,N_119);
nand U1160 (N_1160,In_476,N_184);
and U1161 (N_1161,N_690,N_559);
nor U1162 (N_1162,N_392,N_646);
and U1163 (N_1163,N_751,N_224);
nand U1164 (N_1164,N_735,In_1856);
xor U1165 (N_1165,N_54,N_477);
or U1166 (N_1166,N_514,In_397);
and U1167 (N_1167,N_482,N_563);
nor U1168 (N_1168,N_471,In_1115);
or U1169 (N_1169,N_502,N_351);
and U1170 (N_1170,N_27,N_654);
nand U1171 (N_1171,N_394,N_419);
or U1172 (N_1172,In_1254,N_602);
nor U1173 (N_1173,In_1097,N_293);
nor U1174 (N_1174,N_153,N_137);
nand U1175 (N_1175,In_1913,N_702);
and U1176 (N_1176,N_545,N_781);
and U1177 (N_1177,N_773,In_496);
nor U1178 (N_1178,In_831,N_148);
nor U1179 (N_1179,In_1277,N_5);
xnor U1180 (N_1180,N_149,N_320);
nor U1181 (N_1181,N_405,N_776);
xnor U1182 (N_1182,In_49,In_512);
nor U1183 (N_1183,N_692,N_447);
xor U1184 (N_1184,In_847,In_1028);
or U1185 (N_1185,N_298,N_521);
xor U1186 (N_1186,N_281,N_479);
and U1187 (N_1187,In_1266,N_274);
or U1188 (N_1188,N_497,N_385);
and U1189 (N_1189,N_645,In_1077);
nor U1190 (N_1190,N_683,N_374);
or U1191 (N_1191,N_450,N_791);
and U1192 (N_1192,N_481,N_210);
or U1193 (N_1193,In_509,N_125);
or U1194 (N_1194,N_327,In_402);
or U1195 (N_1195,In_1714,N_330);
nand U1196 (N_1196,N_583,In_1966);
nand U1197 (N_1197,In_811,In_1882);
nor U1198 (N_1198,In_494,N_415);
and U1199 (N_1199,N_616,In_1393);
and U1200 (N_1200,In_255,N_747);
or U1201 (N_1201,N_236,In_501);
or U1202 (N_1202,In_1688,N_586);
or U1203 (N_1203,N_62,N_155);
xnor U1204 (N_1204,N_381,N_691);
and U1205 (N_1205,N_539,N_179);
nand U1206 (N_1206,In_935,N_23);
xor U1207 (N_1207,N_291,In_1428);
and U1208 (N_1208,N_410,N_3);
nand U1209 (N_1209,N_193,In_546);
or U1210 (N_1210,In_357,In_1449);
xor U1211 (N_1211,In_390,In_821);
and U1212 (N_1212,N_664,In_74);
xnor U1213 (N_1213,N_43,In_1391);
or U1214 (N_1214,N_536,In_584);
or U1215 (N_1215,N_476,N_38);
or U1216 (N_1216,N_651,In_139);
nand U1217 (N_1217,N_222,N_280);
nand U1218 (N_1218,N_167,In_795);
or U1219 (N_1219,In_816,N_416);
xor U1220 (N_1220,N_704,N_129);
nor U1221 (N_1221,N_589,In_1098);
nand U1222 (N_1222,N_242,In_1526);
nor U1223 (N_1223,N_768,N_509);
or U1224 (N_1224,N_271,N_299);
xnor U1225 (N_1225,In_1095,N_45);
or U1226 (N_1226,N_106,In_1475);
nor U1227 (N_1227,In_1657,N_144);
and U1228 (N_1228,In_477,N_753);
nor U1229 (N_1229,N_570,N_39);
xnor U1230 (N_1230,N_217,N_722);
nand U1231 (N_1231,In_548,In_84);
and U1232 (N_1232,N_779,In_1748);
or U1233 (N_1233,N_386,In_280);
and U1234 (N_1234,In_147,In_919);
and U1235 (N_1235,N_177,In_57);
nand U1236 (N_1236,In_613,N_344);
nor U1237 (N_1237,In_587,N_607);
and U1238 (N_1238,N_304,N_799);
nor U1239 (N_1239,In_1981,In_1977);
and U1240 (N_1240,N_689,N_92);
xor U1241 (N_1241,N_695,N_94);
and U1242 (N_1242,In_1140,N_792);
or U1243 (N_1243,N_218,N_9);
xor U1244 (N_1244,N_77,N_99);
nor U1245 (N_1245,N_284,In_1079);
and U1246 (N_1246,In_815,N_174);
and U1247 (N_1247,N_637,N_241);
or U1248 (N_1248,In_1215,N_339);
or U1249 (N_1249,In_905,In_1885);
nand U1250 (N_1250,N_786,N_734);
xor U1251 (N_1251,N_12,In_294);
and U1252 (N_1252,In_1459,N_567);
or U1253 (N_1253,N_311,In_686);
and U1254 (N_1254,N_485,N_359);
or U1255 (N_1255,N_657,N_213);
or U1256 (N_1256,In_1341,N_796);
nand U1257 (N_1257,N_400,In_293);
and U1258 (N_1258,N_462,N_717);
nor U1259 (N_1259,N_421,N_88);
nor U1260 (N_1260,In_178,N_762);
or U1261 (N_1261,In_951,N_555);
and U1262 (N_1262,N_249,N_114);
and U1263 (N_1263,N_297,N_643);
xor U1264 (N_1264,In_1989,N_655);
nand U1265 (N_1265,N_362,N_501);
or U1266 (N_1266,In_94,N_358);
and U1267 (N_1267,N_333,In_1829);
and U1268 (N_1268,N_610,N_553);
and U1269 (N_1269,In_820,N_622);
nor U1270 (N_1270,In_194,In_64);
or U1271 (N_1271,N_506,N_798);
or U1272 (N_1272,In_574,N_395);
nand U1273 (N_1273,N_707,In_1193);
nor U1274 (N_1274,In_260,N_439);
nor U1275 (N_1275,In_91,N_56);
or U1276 (N_1276,In_1870,In_1801);
nor U1277 (N_1277,In_611,In_1);
nand U1278 (N_1278,N_541,In_1646);
nand U1279 (N_1279,In_922,N_780);
nand U1280 (N_1280,N_658,N_519);
or U1281 (N_1281,In_432,N_491);
nand U1282 (N_1282,N_372,In_1612);
nor U1283 (N_1283,N_580,N_53);
nor U1284 (N_1284,N_113,In_1069);
nor U1285 (N_1285,N_240,In_117);
nor U1286 (N_1286,N_377,N_590);
and U1287 (N_1287,N_579,N_678);
nand U1288 (N_1288,N_156,In_921);
xor U1289 (N_1289,N_315,N_675);
or U1290 (N_1290,In_673,N_195);
and U1291 (N_1291,In_148,N_767);
nor U1292 (N_1292,N_782,N_674);
nand U1293 (N_1293,N_537,N_176);
xor U1294 (N_1294,N_207,N_494);
or U1295 (N_1295,In_909,In_1751);
nor U1296 (N_1296,In_1680,N_473);
nand U1297 (N_1297,N_76,N_478);
and U1298 (N_1298,In_1927,N_534);
or U1299 (N_1299,N_785,N_404);
nor U1300 (N_1300,In_1373,In_305);
nor U1301 (N_1301,N_24,N_499);
or U1302 (N_1302,N_248,N_721);
and U1303 (N_1303,N_313,N_614);
and U1304 (N_1304,N_644,N_282);
and U1305 (N_1305,N_398,In_410);
and U1306 (N_1306,N_272,N_688);
xnor U1307 (N_1307,In_1370,In_51);
nor U1308 (N_1308,In_1372,N_452);
nor U1309 (N_1309,N_605,N_290);
and U1310 (N_1310,N_25,N_139);
or U1311 (N_1311,N_15,In_499);
nor U1312 (N_1312,In_1983,N_75);
and U1313 (N_1313,In_1877,N_238);
and U1314 (N_1314,N_18,N_243);
nand U1315 (N_1315,N_316,N_587);
xor U1316 (N_1316,N_412,N_373);
or U1317 (N_1317,In_1021,N_29);
or U1318 (N_1318,N_204,N_163);
or U1319 (N_1319,In_702,N_68);
or U1320 (N_1320,In_143,N_393);
nor U1321 (N_1321,N_708,N_46);
xor U1322 (N_1322,N_152,N_440);
nand U1323 (N_1323,In_373,N_200);
or U1324 (N_1324,N_187,N_375);
nor U1325 (N_1325,In_25,N_178);
or U1326 (N_1326,N_411,N_623);
and U1327 (N_1327,N_492,N_188);
xor U1328 (N_1328,N_549,In_1213);
and U1329 (N_1329,N_680,In_1491);
nor U1330 (N_1330,In_908,N_467);
or U1331 (N_1331,In_1664,N_701);
nor U1332 (N_1332,In_822,In_528);
nand U1333 (N_1333,N_681,In_754);
xnor U1334 (N_1334,N_251,N_59);
nor U1335 (N_1335,In_914,In_1619);
or U1336 (N_1336,N_380,In_1899);
nand U1337 (N_1337,N_507,N_52);
or U1338 (N_1338,N_120,N_183);
or U1339 (N_1339,N_511,In_1708);
xnor U1340 (N_1340,In_338,N_262);
nor U1341 (N_1341,In_1403,N_14);
or U1342 (N_1342,In_920,N_368);
and U1343 (N_1343,In_995,N_504);
xnor U1344 (N_1344,N_612,N_498);
nor U1345 (N_1345,In_388,N_523);
or U1346 (N_1346,In_1891,In_123);
and U1347 (N_1347,N_308,N_699);
and U1348 (N_1348,N_444,In_127);
nand U1349 (N_1349,N_255,N_324);
nor U1350 (N_1350,N_212,N_596);
nor U1351 (N_1351,N_277,N_345);
and U1352 (N_1352,N_793,In_463);
or U1353 (N_1353,N_142,In_977);
xor U1354 (N_1354,N_72,N_387);
nand U1355 (N_1355,N_268,In_841);
nor U1356 (N_1356,In_312,N_159);
and U1357 (N_1357,In_1110,In_1015);
and U1358 (N_1358,N_95,N_465);
nand U1359 (N_1359,N_566,N_201);
nand U1360 (N_1360,N_403,N_718);
and U1361 (N_1361,N_470,N_748);
nor U1362 (N_1362,In_1017,In_715);
nor U1363 (N_1363,N_662,In_1068);
or U1364 (N_1364,N_104,N_332);
or U1365 (N_1365,In_1756,N_11);
xor U1366 (N_1366,N_90,N_197);
xor U1367 (N_1367,N_533,In_874);
xor U1368 (N_1368,In_1200,In_713);
or U1369 (N_1369,N_356,N_599);
or U1370 (N_1370,N_366,N_160);
or U1371 (N_1371,N_530,N_353);
xnor U1372 (N_1372,In_1759,In_1453);
and U1373 (N_1373,N_628,N_435);
nand U1374 (N_1374,N_642,N_108);
or U1375 (N_1375,N_305,N_328);
or U1376 (N_1376,N_408,In_487);
xnor U1377 (N_1377,In_828,N_352);
nand U1378 (N_1378,N_565,N_759);
or U1379 (N_1379,N_769,N_369);
xnor U1380 (N_1380,N_239,N_116);
or U1381 (N_1381,N_383,N_428);
or U1382 (N_1382,N_738,N_301);
xor U1383 (N_1383,In_1091,In_346);
and U1384 (N_1384,In_963,In_277);
xnor U1385 (N_1385,In_1833,N_540);
nand U1386 (N_1386,N_289,In_1008);
or U1387 (N_1387,N_283,N_364);
and U1388 (N_1388,N_16,N_585);
nor U1389 (N_1389,N_141,In_547);
and U1390 (N_1390,N_417,In_553);
or U1391 (N_1391,N_81,In_1694);
nand U1392 (N_1392,In_1601,In_773);
or U1393 (N_1393,N_1,N_426);
or U1394 (N_1394,N_719,N_740);
nor U1395 (N_1395,N_326,N_713);
xnor U1396 (N_1396,N_186,N_558);
nand U1397 (N_1397,In_1025,N_157);
xnor U1398 (N_1398,In_583,N_469);
nand U1399 (N_1399,N_48,N_135);
and U1400 (N_1400,N_587,N_195);
and U1401 (N_1401,In_178,In_1833);
or U1402 (N_1402,N_487,N_729);
nand U1403 (N_1403,N_16,N_31);
or U1404 (N_1404,N_580,N_592);
nor U1405 (N_1405,N_97,N_561);
or U1406 (N_1406,N_310,In_538);
or U1407 (N_1407,N_175,N_49);
and U1408 (N_1408,N_464,N_236);
nand U1409 (N_1409,N_196,N_424);
nand U1410 (N_1410,N_175,In_1069);
and U1411 (N_1411,N_264,N_126);
nor U1412 (N_1412,N_426,N_686);
and U1413 (N_1413,N_493,N_500);
nor U1414 (N_1414,N_78,N_693);
and U1415 (N_1415,In_1725,N_566);
xor U1416 (N_1416,In_1836,N_169);
nand U1417 (N_1417,In_21,In_820);
nor U1418 (N_1418,In_1449,N_188);
nand U1419 (N_1419,N_482,In_117);
or U1420 (N_1420,N_199,N_54);
nor U1421 (N_1421,In_1271,In_1284);
nor U1422 (N_1422,N_19,In_394);
and U1423 (N_1423,N_525,N_452);
and U1424 (N_1424,N_372,In_300);
xor U1425 (N_1425,N_400,N_504);
nand U1426 (N_1426,N_463,In_581);
xor U1427 (N_1427,N_191,In_957);
and U1428 (N_1428,In_669,N_748);
nor U1429 (N_1429,In_1826,In_574);
nand U1430 (N_1430,In_138,N_314);
nor U1431 (N_1431,N_361,In_1644);
xor U1432 (N_1432,N_576,In_1664);
nand U1433 (N_1433,N_31,N_316);
and U1434 (N_1434,In_293,N_25);
and U1435 (N_1435,N_567,N_425);
xor U1436 (N_1436,In_1204,In_74);
and U1437 (N_1437,In_1980,In_919);
nand U1438 (N_1438,In_1899,In_138);
nand U1439 (N_1439,N_762,N_95);
nor U1440 (N_1440,In_1028,N_311);
and U1441 (N_1441,N_628,N_363);
nand U1442 (N_1442,N_495,In_1213);
or U1443 (N_1443,In_1647,N_471);
xor U1444 (N_1444,N_86,N_286);
or U1445 (N_1445,N_546,In_1158);
nand U1446 (N_1446,N_516,N_215);
nand U1447 (N_1447,N_173,In_905);
xor U1448 (N_1448,N_229,N_554);
nand U1449 (N_1449,N_97,N_285);
nor U1450 (N_1450,In_504,In_1391);
nand U1451 (N_1451,N_473,N_480);
nor U1452 (N_1452,N_770,In_1428);
xnor U1453 (N_1453,In_1826,In_963);
nor U1454 (N_1454,In_648,In_793);
or U1455 (N_1455,In_1403,N_463);
xnor U1456 (N_1456,In_1097,In_1646);
nor U1457 (N_1457,N_430,N_509);
nand U1458 (N_1458,N_699,N_559);
nor U1459 (N_1459,N_683,N_426);
xnor U1460 (N_1460,In_245,In_91);
and U1461 (N_1461,In_471,N_615);
nor U1462 (N_1462,N_326,In_75);
xnor U1463 (N_1463,In_1857,N_199);
or U1464 (N_1464,In_1168,N_732);
and U1465 (N_1465,N_313,N_140);
xor U1466 (N_1466,N_339,N_569);
xor U1467 (N_1467,N_207,In_845);
nand U1468 (N_1468,N_159,N_51);
or U1469 (N_1469,In_1836,N_664);
xor U1470 (N_1470,N_6,In_443);
or U1471 (N_1471,In_1403,N_752);
nand U1472 (N_1472,N_350,N_596);
and U1473 (N_1473,N_736,In_1915);
and U1474 (N_1474,In_1075,In_1614);
nand U1475 (N_1475,N_436,N_508);
or U1476 (N_1476,N_733,N_32);
nor U1477 (N_1477,N_73,N_497);
nand U1478 (N_1478,N_427,N_604);
or U1479 (N_1479,N_360,In_1630);
nand U1480 (N_1480,N_15,N_559);
and U1481 (N_1481,In_1833,N_265);
and U1482 (N_1482,In_1636,N_195);
nor U1483 (N_1483,N_250,In_845);
or U1484 (N_1484,N_717,N_490);
nor U1485 (N_1485,In_1592,N_290);
nand U1486 (N_1486,N_691,N_34);
nand U1487 (N_1487,N_420,N_101);
or U1488 (N_1488,N_10,N_688);
xnor U1489 (N_1489,N_532,In_259);
and U1490 (N_1490,In_572,N_630);
and U1491 (N_1491,N_150,N_107);
nand U1492 (N_1492,In_802,In_572);
and U1493 (N_1493,In_139,In_1471);
xor U1494 (N_1494,N_567,N_431);
or U1495 (N_1495,N_674,N_279);
nand U1496 (N_1496,In_1158,N_528);
xor U1497 (N_1497,In_1428,In_258);
nor U1498 (N_1498,N_412,N_248);
and U1499 (N_1499,In_1069,N_795);
xor U1500 (N_1500,In_1785,N_100);
xor U1501 (N_1501,In_820,In_734);
xnor U1502 (N_1502,N_483,N_737);
nor U1503 (N_1503,In_21,In_1379);
xor U1504 (N_1504,N_370,N_66);
nor U1505 (N_1505,N_401,N_291);
or U1506 (N_1506,N_645,N_636);
or U1507 (N_1507,In_553,In_613);
and U1508 (N_1508,N_125,In_845);
or U1509 (N_1509,In_1045,In_1250);
xor U1510 (N_1510,In_353,In_117);
xnor U1511 (N_1511,N_504,N_34);
nand U1512 (N_1512,N_332,N_680);
nor U1513 (N_1513,In_713,N_396);
nand U1514 (N_1514,N_279,N_181);
and U1515 (N_1515,N_314,N_769);
nor U1516 (N_1516,N_678,In_1997);
and U1517 (N_1517,N_592,N_700);
or U1518 (N_1518,In_1977,In_762);
nand U1519 (N_1519,N_73,In_1662);
or U1520 (N_1520,N_241,N_717);
nor U1521 (N_1521,N_42,N_126);
nor U1522 (N_1522,N_703,N_278);
and U1523 (N_1523,N_392,N_572);
xor U1524 (N_1524,N_306,In_734);
or U1525 (N_1525,N_551,N_447);
nor U1526 (N_1526,In_1820,N_240);
or U1527 (N_1527,N_723,N_30);
and U1528 (N_1528,In_383,N_274);
and U1529 (N_1529,N_147,N_233);
xnor U1530 (N_1530,N_232,N_742);
nand U1531 (N_1531,N_348,N_769);
xor U1532 (N_1532,N_61,N_464);
or U1533 (N_1533,In_490,N_118);
and U1534 (N_1534,In_1277,N_247);
nor U1535 (N_1535,In_1229,In_1309);
nand U1536 (N_1536,N_321,N_57);
and U1537 (N_1537,N_359,In_1927);
or U1538 (N_1538,In_256,N_659);
or U1539 (N_1539,In_1526,N_517);
nand U1540 (N_1540,N_610,In_260);
xnor U1541 (N_1541,N_405,In_477);
and U1542 (N_1542,N_363,In_603);
xnor U1543 (N_1543,N_735,N_161);
xnor U1544 (N_1544,N_784,N_335);
nor U1545 (N_1545,N_446,N_556);
nand U1546 (N_1546,N_640,N_261);
or U1547 (N_1547,N_570,N_737);
nor U1548 (N_1548,N_454,N_229);
xnor U1549 (N_1549,In_1614,In_874);
nand U1550 (N_1550,In_795,N_778);
nand U1551 (N_1551,N_141,N_71);
or U1552 (N_1552,In_548,In_581);
nand U1553 (N_1553,N_280,N_784);
and U1554 (N_1554,In_1296,In_1647);
nor U1555 (N_1555,N_703,N_528);
and U1556 (N_1556,In_1601,In_656);
and U1557 (N_1557,N_155,In_1175);
nor U1558 (N_1558,N_177,In_1820);
or U1559 (N_1559,N_555,N_136);
nand U1560 (N_1560,N_326,N_50);
nand U1561 (N_1561,In_255,N_110);
nor U1562 (N_1562,N_153,In_118);
and U1563 (N_1563,N_449,In_816);
or U1564 (N_1564,N_172,N_776);
xor U1565 (N_1565,N_762,N_489);
and U1566 (N_1566,In_934,N_747);
or U1567 (N_1567,N_793,In_906);
nand U1568 (N_1568,N_69,N_477);
nor U1569 (N_1569,N_133,In_1284);
xnor U1570 (N_1570,N_336,In_604);
or U1571 (N_1571,In_1882,N_476);
nand U1572 (N_1572,N_319,N_584);
nand U1573 (N_1573,N_427,N_628);
and U1574 (N_1574,N_696,N_110);
nor U1575 (N_1575,N_370,In_1891);
and U1576 (N_1576,In_734,N_418);
or U1577 (N_1577,N_308,N_279);
nand U1578 (N_1578,N_703,N_61);
and U1579 (N_1579,In_427,N_782);
or U1580 (N_1580,N_129,N_622);
or U1581 (N_1581,N_44,N_99);
nand U1582 (N_1582,In_299,N_482);
and U1583 (N_1583,N_423,N_169);
xor U1584 (N_1584,In_1229,N_637);
and U1585 (N_1585,In_1528,N_785);
and U1586 (N_1586,N_301,N_607);
and U1587 (N_1587,N_578,In_890);
and U1588 (N_1588,N_557,In_1611);
or U1589 (N_1589,N_0,N_531);
or U1590 (N_1590,N_109,In_845);
xnor U1591 (N_1591,N_126,N_483);
nand U1592 (N_1592,N_347,N_781);
and U1593 (N_1593,N_404,N_726);
xor U1594 (N_1594,N_498,N_465);
and U1595 (N_1595,N_633,In_1826);
nand U1596 (N_1596,In_1808,N_220);
xnor U1597 (N_1597,N_663,N_161);
nand U1598 (N_1598,N_794,N_291);
xnor U1599 (N_1599,N_384,In_914);
and U1600 (N_1600,N_1225,N_846);
nor U1601 (N_1601,N_1174,N_1037);
nor U1602 (N_1602,N_1502,N_1253);
nor U1603 (N_1603,N_1335,N_1558);
and U1604 (N_1604,N_1330,N_1126);
xor U1605 (N_1605,N_1471,N_1547);
xor U1606 (N_1606,N_1531,N_1185);
and U1607 (N_1607,N_843,N_873);
and U1608 (N_1608,N_1306,N_815);
and U1609 (N_1609,N_1570,N_1535);
xor U1610 (N_1610,N_1116,N_1396);
or U1611 (N_1611,N_1114,N_1493);
xnor U1612 (N_1612,N_1569,N_829);
nand U1613 (N_1613,N_915,N_1244);
nor U1614 (N_1614,N_1394,N_1473);
and U1615 (N_1615,N_1033,N_1053);
xor U1616 (N_1616,N_1424,N_1525);
and U1617 (N_1617,N_842,N_880);
and U1618 (N_1618,N_803,N_1044);
xor U1619 (N_1619,N_1428,N_1011);
nand U1620 (N_1620,N_1417,N_1405);
xnor U1621 (N_1621,N_805,N_824);
nor U1622 (N_1622,N_1338,N_1071);
nor U1623 (N_1623,N_1314,N_1495);
and U1624 (N_1624,N_865,N_1410);
nand U1625 (N_1625,N_1542,N_897);
xnor U1626 (N_1626,N_812,N_1197);
or U1627 (N_1627,N_1040,N_917);
nor U1628 (N_1628,N_1256,N_976);
xnor U1629 (N_1629,N_1128,N_1597);
xnor U1630 (N_1630,N_1595,N_832);
xnor U1631 (N_1631,N_935,N_1492);
and U1632 (N_1632,N_1389,N_1453);
or U1633 (N_1633,N_1480,N_1586);
nand U1634 (N_1634,N_1085,N_1333);
nand U1635 (N_1635,N_1252,N_1274);
nor U1636 (N_1636,N_1002,N_979);
nor U1637 (N_1637,N_1401,N_1121);
nand U1638 (N_1638,N_1235,N_826);
nor U1639 (N_1639,N_1350,N_949);
xnor U1640 (N_1640,N_1519,N_1248);
and U1641 (N_1641,N_1233,N_1251);
xor U1642 (N_1642,N_964,N_1474);
or U1643 (N_1643,N_877,N_1568);
xor U1644 (N_1644,N_958,N_867);
xnor U1645 (N_1645,N_1511,N_982);
or U1646 (N_1646,N_1107,N_1022);
or U1647 (N_1647,N_1392,N_1470);
or U1648 (N_1648,N_888,N_1352);
and U1649 (N_1649,N_990,N_1269);
and U1650 (N_1650,N_1412,N_1151);
and U1651 (N_1651,N_1211,N_1052);
or U1652 (N_1652,N_1353,N_1305);
or U1653 (N_1653,N_1099,N_1489);
nor U1654 (N_1654,N_1245,N_1193);
and U1655 (N_1655,N_1092,N_942);
nor U1656 (N_1656,N_1190,N_1295);
xor U1657 (N_1657,N_1021,N_1390);
nand U1658 (N_1658,N_1215,N_1501);
nor U1659 (N_1659,N_1342,N_1194);
and U1660 (N_1660,N_1339,N_1458);
nor U1661 (N_1661,N_1210,N_1195);
xor U1662 (N_1662,N_1323,N_893);
and U1663 (N_1663,N_1157,N_866);
nor U1664 (N_1664,N_831,N_1036);
xnor U1665 (N_1665,N_1191,N_927);
or U1666 (N_1666,N_1562,N_1388);
nor U1667 (N_1667,N_1178,N_890);
and U1668 (N_1668,N_965,N_1315);
nor U1669 (N_1669,N_951,N_1540);
xor U1670 (N_1670,N_1188,N_1443);
and U1671 (N_1671,N_1187,N_827);
or U1672 (N_1672,N_1283,N_1205);
and U1673 (N_1673,N_1346,N_1119);
nor U1674 (N_1674,N_1160,N_1059);
and U1675 (N_1675,N_910,N_1219);
nand U1676 (N_1676,N_941,N_1249);
nor U1677 (N_1677,N_845,N_1406);
and U1678 (N_1678,N_889,N_1578);
or U1679 (N_1679,N_1364,N_1423);
and U1680 (N_1680,N_1148,N_852);
or U1681 (N_1681,N_948,N_1505);
or U1682 (N_1682,N_1538,N_1327);
xnor U1683 (N_1683,N_804,N_1290);
xnor U1684 (N_1684,N_1476,N_820);
and U1685 (N_1685,N_901,N_1276);
and U1686 (N_1686,N_1477,N_981);
nor U1687 (N_1687,N_1077,N_836);
or U1688 (N_1688,N_977,N_1436);
nand U1689 (N_1689,N_1220,N_1294);
or U1690 (N_1690,N_1045,N_1017);
xor U1691 (N_1691,N_1367,N_1361);
or U1692 (N_1692,N_1204,N_1246);
or U1693 (N_1693,N_851,N_1432);
nand U1694 (N_1694,N_1326,N_1387);
nand U1695 (N_1695,N_1563,N_1241);
and U1696 (N_1696,N_1167,N_1213);
xnor U1697 (N_1697,N_878,N_1403);
xnor U1698 (N_1698,N_1302,N_1025);
nand U1699 (N_1699,N_973,N_1574);
and U1700 (N_1700,N_1583,N_819);
xor U1701 (N_1701,N_1529,N_1404);
or U1702 (N_1702,N_1226,N_997);
nand U1703 (N_1703,N_1012,N_1334);
xor U1704 (N_1704,N_1242,N_859);
nor U1705 (N_1705,N_929,N_811);
nor U1706 (N_1706,N_985,N_1081);
or U1707 (N_1707,N_1561,N_1039);
or U1708 (N_1708,N_1023,N_924);
or U1709 (N_1709,N_808,N_969);
and U1710 (N_1710,N_1196,N_1240);
xor U1711 (N_1711,N_1008,N_908);
or U1712 (N_1712,N_1451,N_1509);
and U1713 (N_1713,N_1236,N_986);
or U1714 (N_1714,N_926,N_800);
xor U1715 (N_1715,N_925,N_1309);
or U1716 (N_1716,N_974,N_984);
xnor U1717 (N_1717,N_892,N_1180);
nor U1718 (N_1718,N_1091,N_1299);
nand U1719 (N_1719,N_1170,N_1397);
nor U1720 (N_1720,N_874,N_922);
or U1721 (N_1721,N_1541,N_904);
nor U1722 (N_1722,N_1006,N_998);
or U1723 (N_1723,N_839,N_1445);
and U1724 (N_1724,N_1175,N_1238);
and U1725 (N_1725,N_1065,N_857);
nor U1726 (N_1726,N_1115,N_1186);
and U1727 (N_1727,N_1227,N_817);
or U1728 (N_1728,N_1551,N_1153);
xnor U1729 (N_1729,N_1325,N_1136);
xnor U1730 (N_1730,N_863,N_1328);
xor U1731 (N_1731,N_813,N_1166);
or U1732 (N_1732,N_1499,N_1588);
xnor U1733 (N_1733,N_1598,N_900);
or U1734 (N_1734,N_1014,N_1061);
and U1735 (N_1735,N_907,N_1035);
and U1736 (N_1736,N_1019,N_1341);
nor U1737 (N_1737,N_967,N_809);
and U1738 (N_1738,N_911,N_1377);
xor U1739 (N_1739,N_1265,N_828);
or U1740 (N_1740,N_1144,N_1078);
xor U1741 (N_1741,N_838,N_1552);
xnor U1742 (N_1742,N_1056,N_1123);
nor U1743 (N_1743,N_980,N_1366);
nor U1744 (N_1744,N_1537,N_1281);
or U1745 (N_1745,N_1169,N_1267);
xor U1746 (N_1746,N_1082,N_1332);
nor U1747 (N_1747,N_930,N_1047);
nor U1748 (N_1748,N_1407,N_1359);
nand U1749 (N_1749,N_834,N_850);
nor U1750 (N_1750,N_899,N_960);
xor U1751 (N_1751,N_1516,N_989);
nand U1752 (N_1752,N_1369,N_1110);
or U1753 (N_1753,N_1310,N_818);
nor U1754 (N_1754,N_1032,N_1468);
nand U1755 (N_1755,N_1182,N_1321);
and U1756 (N_1756,N_1122,N_1523);
and U1757 (N_1757,N_1076,N_1273);
xor U1758 (N_1758,N_1582,N_1447);
and U1759 (N_1759,N_1254,N_1429);
or U1760 (N_1760,N_928,N_1131);
and U1761 (N_1761,N_1408,N_1336);
and U1762 (N_1762,N_1046,N_1137);
and U1763 (N_1763,N_821,N_1420);
and U1764 (N_1764,N_1132,N_1030);
xnor U1765 (N_1765,N_1209,N_1288);
or U1766 (N_1766,N_1100,N_1101);
or U1767 (N_1767,N_1097,N_946);
nor U1768 (N_1768,N_1400,N_1293);
and U1769 (N_1769,N_1120,N_1413);
and U1770 (N_1770,N_1374,N_1015);
or U1771 (N_1771,N_1340,N_991);
and U1772 (N_1772,N_1384,N_1064);
xor U1773 (N_1773,N_1434,N_1171);
and U1774 (N_1774,N_1522,N_1347);
xor U1775 (N_1775,N_870,N_921);
and U1776 (N_1776,N_1286,N_1319);
xnor U1777 (N_1777,N_995,N_896);
or U1778 (N_1778,N_1393,N_1284);
and U1779 (N_1779,N_1356,N_1221);
or U1780 (N_1780,N_970,N_1010);
xor U1781 (N_1781,N_1557,N_1280);
nor U1782 (N_1782,N_1231,N_1318);
and U1783 (N_1783,N_894,N_1192);
nand U1784 (N_1784,N_1165,N_1460);
or U1785 (N_1785,N_835,N_1358);
nor U1786 (N_1786,N_1093,N_1088);
and U1787 (N_1787,N_1202,N_1313);
nor U1788 (N_1788,N_1365,N_1544);
nand U1789 (N_1789,N_1060,N_1150);
or U1790 (N_1790,N_1255,N_1571);
and U1791 (N_1791,N_1034,N_1592);
and U1792 (N_1792,N_1074,N_884);
and U1793 (N_1793,N_1376,N_1134);
and U1794 (N_1794,N_1243,N_876);
or U1795 (N_1795,N_840,N_833);
nor U1796 (N_1796,N_1285,N_1158);
or U1797 (N_1797,N_1068,N_1520);
nor U1798 (N_1798,N_919,N_822);
xnor U1799 (N_1799,N_1380,N_1534);
xnor U1800 (N_1800,N_1168,N_1536);
xor U1801 (N_1801,N_903,N_905);
xor U1802 (N_1802,N_923,N_1086);
and U1803 (N_1803,N_871,N_841);
or U1804 (N_1804,N_1257,N_1062);
and U1805 (N_1805,N_1512,N_933);
xnor U1806 (N_1806,N_1431,N_1289);
nand U1807 (N_1807,N_1018,N_1212);
nor U1808 (N_1808,N_1222,N_1138);
or U1809 (N_1809,N_1206,N_1362);
xnor U1810 (N_1810,N_1312,N_1133);
nor U1811 (N_1811,N_1503,N_1539);
nor U1812 (N_1812,N_1456,N_961);
xnor U1813 (N_1813,N_1268,N_1108);
or U1814 (N_1814,N_1141,N_1135);
or U1815 (N_1815,N_1223,N_1435);
and U1816 (N_1816,N_1024,N_1229);
and U1817 (N_1817,N_1363,N_1079);
and U1818 (N_1818,N_1069,N_955);
and U1819 (N_1819,N_1430,N_993);
or U1820 (N_1820,N_1467,N_1560);
or U1821 (N_1821,N_1016,N_1200);
or U1822 (N_1822,N_1442,N_1124);
nor U1823 (N_1823,N_1103,N_1344);
nand U1824 (N_1824,N_1043,N_1510);
or U1825 (N_1825,N_1308,N_1084);
xor U1826 (N_1826,N_1438,N_1130);
nand U1827 (N_1827,N_1360,N_895);
nand U1828 (N_1828,N_875,N_1567);
or U1829 (N_1829,N_1409,N_1482);
and U1830 (N_1830,N_1232,N_883);
or U1831 (N_1831,N_914,N_1080);
nor U1832 (N_1832,N_1096,N_1524);
and U1833 (N_1833,N_988,N_1263);
or U1834 (N_1834,N_1398,N_1465);
xnor U1835 (N_1835,N_1070,N_1307);
nor U1836 (N_1836,N_1304,N_1581);
nor U1837 (N_1837,N_1508,N_1322);
and U1838 (N_1838,N_1565,N_1147);
or U1839 (N_1839,N_1426,N_856);
and U1840 (N_1840,N_1207,N_952);
or U1841 (N_1841,N_1298,N_978);
xor U1842 (N_1842,N_1452,N_802);
xnor U1843 (N_1843,N_1320,N_1555);
and U1844 (N_1844,N_1554,N_1441);
or U1845 (N_1845,N_1262,N_1464);
or U1846 (N_1846,N_1593,N_1486);
xor U1847 (N_1847,N_855,N_1585);
nor U1848 (N_1848,N_1007,N_1031);
nor U1849 (N_1849,N_1083,N_1282);
or U1850 (N_1850,N_934,N_1026);
xor U1851 (N_1851,N_1425,N_1051);
nor U1852 (N_1852,N_887,N_1479);
nand U1853 (N_1853,N_1278,N_1041);
and U1854 (N_1854,N_1530,N_1533);
nand U1855 (N_1855,N_810,N_1230);
nand U1856 (N_1856,N_1239,N_848);
and U1857 (N_1857,N_1004,N_971);
or U1858 (N_1858,N_1543,N_1378);
and U1859 (N_1859,N_814,N_1020);
or U1860 (N_1860,N_1548,N_1275);
or U1861 (N_1861,N_860,N_1271);
xnor U1862 (N_1862,N_1348,N_1472);
and U1863 (N_1863,N_1549,N_1528);
and U1864 (N_1864,N_1237,N_1422);
nand U1865 (N_1865,N_906,N_847);
or U1866 (N_1866,N_972,N_1500);
or U1867 (N_1867,N_1596,N_1573);
nor U1868 (N_1868,N_937,N_1514);
and U1869 (N_1869,N_1439,N_1487);
or U1870 (N_1870,N_956,N_1095);
nand U1871 (N_1871,N_1279,N_1556);
nand U1872 (N_1872,N_1264,N_1457);
or U1873 (N_1873,N_1090,N_1550);
or U1874 (N_1874,N_1161,N_1001);
xor U1875 (N_1875,N_1112,N_1266);
xnor U1876 (N_1876,N_1559,N_1507);
or U1877 (N_1877,N_1277,N_891);
xor U1878 (N_1878,N_1444,N_1216);
nor U1879 (N_1879,N_1349,N_1203);
nor U1880 (N_1880,N_1357,N_1272);
or U1881 (N_1881,N_944,N_909);
and U1882 (N_1882,N_1475,N_1270);
nor U1883 (N_1883,N_885,N_872);
or U1884 (N_1884,N_1139,N_1433);
xor U1885 (N_1885,N_1201,N_1485);
or U1886 (N_1886,N_1454,N_1427);
xnor U1887 (N_1887,N_807,N_1504);
or U1888 (N_1888,N_1234,N_1189);
xor U1889 (N_1889,N_1466,N_1580);
or U1890 (N_1890,N_1129,N_1117);
and U1891 (N_1891,N_912,N_940);
nand U1892 (N_1892,N_837,N_1073);
and U1893 (N_1893,N_1446,N_1553);
and U1894 (N_1894,N_879,N_1156);
and U1895 (N_1895,N_1164,N_1013);
nor U1896 (N_1896,N_1143,N_1455);
xnor U1897 (N_1897,N_1584,N_1214);
nor U1898 (N_1898,N_1411,N_1145);
and U1899 (N_1899,N_950,N_806);
and U1900 (N_1900,N_1048,N_1337);
xor U1901 (N_1901,N_918,N_1343);
nor U1902 (N_1902,N_1055,N_1478);
nor U1903 (N_1903,N_869,N_1247);
or U1904 (N_1904,N_1149,N_987);
or U1905 (N_1905,N_1217,N_1414);
and U1906 (N_1906,N_954,N_1513);
or U1907 (N_1907,N_1009,N_1463);
and U1908 (N_1908,N_881,N_1259);
or U1909 (N_1909,N_1483,N_994);
xnor U1910 (N_1910,N_1449,N_1075);
nor U1911 (N_1911,N_862,N_939);
nor U1912 (N_1912,N_1515,N_1375);
or U1913 (N_1913,N_999,N_1029);
nand U1914 (N_1914,N_849,N_1287);
nor U1915 (N_1915,N_1459,N_1526);
nand U1916 (N_1916,N_1163,N_1419);
nand U1917 (N_1917,N_1300,N_1106);
and U1918 (N_1918,N_936,N_1368);
xor U1919 (N_1919,N_957,N_1498);
nand U1920 (N_1920,N_1575,N_913);
nand U1921 (N_1921,N_1506,N_853);
nand U1922 (N_1922,N_1317,N_1469);
xor U1923 (N_1923,N_1000,N_1146);
xnor U1924 (N_1924,N_1228,N_1354);
nand U1925 (N_1925,N_1104,N_1003);
nand U1926 (N_1926,N_1379,N_1329);
or U1927 (N_1927,N_1291,N_1049);
nand U1928 (N_1928,N_1564,N_1102);
nand U1929 (N_1929,N_1373,N_1311);
nor U1930 (N_1930,N_1415,N_1181);
xor U1931 (N_1931,N_1301,N_1063);
nand U1932 (N_1932,N_1050,N_1518);
or U1933 (N_1933,N_1027,N_1572);
nand U1934 (N_1934,N_1038,N_1589);
nand U1935 (N_1935,N_1587,N_1261);
or U1936 (N_1936,N_1395,N_1067);
xnor U1937 (N_1937,N_1383,N_1494);
nor U1938 (N_1938,N_931,N_1058);
nand U1939 (N_1939,N_916,N_1042);
and U1940 (N_1940,N_1224,N_983);
nand U1941 (N_1941,N_1385,N_1517);
xnor U1942 (N_1942,N_1154,N_1303);
nor U1943 (N_1943,N_844,N_1546);
and U1944 (N_1944,N_1527,N_1028);
nor U1945 (N_1945,N_1316,N_886);
xor U1946 (N_1946,N_1250,N_1450);
and U1947 (N_1947,N_1297,N_1142);
and U1948 (N_1948,N_1576,N_882);
nor U1949 (N_1949,N_1066,N_1173);
and U1950 (N_1950,N_1094,N_920);
nand U1951 (N_1951,N_1462,N_1098);
and U1952 (N_1952,N_1416,N_1109);
nor U1953 (N_1953,N_1448,N_1199);
and U1954 (N_1954,N_1198,N_1345);
xnor U1955 (N_1955,N_962,N_1176);
nand U1956 (N_1956,N_963,N_1496);
and U1957 (N_1957,N_823,N_1497);
and U1958 (N_1958,N_1545,N_1391);
xnor U1959 (N_1959,N_1057,N_801);
and U1960 (N_1960,N_1159,N_1566);
or U1961 (N_1961,N_1111,N_992);
or U1962 (N_1962,N_1437,N_1488);
and U1963 (N_1963,N_1208,N_1292);
xor U1964 (N_1964,N_1118,N_1127);
nand U1965 (N_1965,N_902,N_1183);
nand U1966 (N_1966,N_830,N_968);
nor U1967 (N_1967,N_861,N_1440);
and U1968 (N_1968,N_1590,N_898);
or U1969 (N_1969,N_1105,N_932);
nand U1970 (N_1970,N_953,N_1152);
xor U1971 (N_1971,N_1577,N_959);
xnor U1972 (N_1972,N_1532,N_1072);
xnor U1973 (N_1973,N_1418,N_1054);
and U1974 (N_1974,N_975,N_1386);
nor U1975 (N_1975,N_868,N_1113);
or U1976 (N_1976,N_966,N_1579);
or U1977 (N_1977,N_1421,N_1491);
xnor U1978 (N_1978,N_1490,N_858);
nand U1979 (N_1979,N_1481,N_1399);
nor U1980 (N_1980,N_854,N_1461);
or U1981 (N_1981,N_1179,N_1599);
nand U1982 (N_1982,N_864,N_1324);
or U1983 (N_1983,N_1140,N_1162);
and U1984 (N_1984,N_1370,N_1087);
nand U1985 (N_1985,N_1382,N_1260);
xnor U1986 (N_1986,N_945,N_1521);
nand U1987 (N_1987,N_1591,N_1184);
nor U1988 (N_1988,N_1402,N_825);
or U1989 (N_1989,N_1594,N_1177);
or U1990 (N_1990,N_816,N_1155);
nand U1991 (N_1991,N_938,N_1351);
nor U1992 (N_1992,N_1125,N_1371);
xnor U1993 (N_1993,N_1381,N_996);
nor U1994 (N_1994,N_1258,N_1331);
nor U1995 (N_1995,N_1296,N_1355);
nor U1996 (N_1996,N_943,N_1005);
and U1997 (N_1997,N_1372,N_1484);
xnor U1998 (N_1998,N_1218,N_947);
and U1999 (N_1999,N_1089,N_1172);
and U2000 (N_2000,N_1303,N_1196);
xor U2001 (N_2001,N_1445,N_874);
nand U2002 (N_2002,N_1375,N_1251);
xnor U2003 (N_2003,N_1192,N_1257);
nor U2004 (N_2004,N_888,N_1023);
nor U2005 (N_2005,N_1010,N_1197);
nand U2006 (N_2006,N_1562,N_890);
and U2007 (N_2007,N_1352,N_896);
nand U2008 (N_2008,N_1013,N_948);
or U2009 (N_2009,N_1494,N_1584);
and U2010 (N_2010,N_906,N_1348);
and U2011 (N_2011,N_1276,N_1272);
nand U2012 (N_2012,N_1490,N_1472);
xor U2013 (N_2013,N_979,N_1140);
xnor U2014 (N_2014,N_1406,N_1519);
nor U2015 (N_2015,N_1511,N_866);
nor U2016 (N_2016,N_1084,N_1273);
xnor U2017 (N_2017,N_1277,N_992);
and U2018 (N_2018,N_1355,N_935);
or U2019 (N_2019,N_1586,N_1237);
and U2020 (N_2020,N_1305,N_1392);
xnor U2021 (N_2021,N_879,N_1250);
nor U2022 (N_2022,N_1547,N_1513);
xor U2023 (N_2023,N_1504,N_1394);
or U2024 (N_2024,N_1049,N_1474);
nand U2025 (N_2025,N_1206,N_1302);
and U2026 (N_2026,N_1399,N_1296);
nand U2027 (N_2027,N_1512,N_1544);
and U2028 (N_2028,N_1514,N_817);
nand U2029 (N_2029,N_1499,N_1364);
nor U2030 (N_2030,N_1443,N_1410);
nor U2031 (N_2031,N_928,N_946);
or U2032 (N_2032,N_1077,N_880);
nand U2033 (N_2033,N_1551,N_1488);
nand U2034 (N_2034,N_806,N_1450);
xor U2035 (N_2035,N_1147,N_1069);
xnor U2036 (N_2036,N_1064,N_1054);
nor U2037 (N_2037,N_1435,N_1072);
xor U2038 (N_2038,N_1173,N_828);
nand U2039 (N_2039,N_1159,N_1595);
and U2040 (N_2040,N_1030,N_1278);
and U2041 (N_2041,N_1460,N_1157);
and U2042 (N_2042,N_1391,N_983);
xnor U2043 (N_2043,N_943,N_1470);
nand U2044 (N_2044,N_1358,N_1386);
nor U2045 (N_2045,N_1117,N_808);
nand U2046 (N_2046,N_1382,N_1252);
and U2047 (N_2047,N_1122,N_1534);
xnor U2048 (N_2048,N_1262,N_1041);
nand U2049 (N_2049,N_1072,N_1007);
nor U2050 (N_2050,N_959,N_971);
and U2051 (N_2051,N_856,N_1065);
xnor U2052 (N_2052,N_1561,N_1598);
xor U2053 (N_2053,N_1116,N_1301);
nor U2054 (N_2054,N_1344,N_1503);
or U2055 (N_2055,N_994,N_1367);
xor U2056 (N_2056,N_1484,N_1104);
and U2057 (N_2057,N_1395,N_1518);
and U2058 (N_2058,N_1197,N_1287);
nor U2059 (N_2059,N_1437,N_1571);
xnor U2060 (N_2060,N_1064,N_1546);
nand U2061 (N_2061,N_1122,N_1525);
or U2062 (N_2062,N_1451,N_1090);
nor U2063 (N_2063,N_1089,N_910);
nor U2064 (N_2064,N_1084,N_803);
or U2065 (N_2065,N_814,N_847);
nand U2066 (N_2066,N_1008,N_1424);
xnor U2067 (N_2067,N_1008,N_1160);
nor U2068 (N_2068,N_1303,N_1272);
nor U2069 (N_2069,N_883,N_1527);
xor U2070 (N_2070,N_993,N_812);
or U2071 (N_2071,N_825,N_842);
and U2072 (N_2072,N_1438,N_1175);
or U2073 (N_2073,N_1059,N_955);
and U2074 (N_2074,N_1070,N_906);
nor U2075 (N_2075,N_898,N_936);
or U2076 (N_2076,N_923,N_1323);
xnor U2077 (N_2077,N_974,N_1585);
nand U2078 (N_2078,N_1343,N_1203);
or U2079 (N_2079,N_1203,N_1559);
and U2080 (N_2080,N_1031,N_1368);
nand U2081 (N_2081,N_1001,N_805);
nor U2082 (N_2082,N_1060,N_1552);
xnor U2083 (N_2083,N_1147,N_842);
or U2084 (N_2084,N_841,N_1328);
or U2085 (N_2085,N_1479,N_1476);
or U2086 (N_2086,N_1001,N_1356);
nor U2087 (N_2087,N_1241,N_1274);
nand U2088 (N_2088,N_1335,N_1261);
nand U2089 (N_2089,N_1244,N_1304);
nor U2090 (N_2090,N_1294,N_1119);
nor U2091 (N_2091,N_833,N_986);
and U2092 (N_2092,N_938,N_1547);
nand U2093 (N_2093,N_1546,N_1178);
or U2094 (N_2094,N_1372,N_1516);
or U2095 (N_2095,N_1515,N_838);
xnor U2096 (N_2096,N_1307,N_1504);
nand U2097 (N_2097,N_1236,N_926);
and U2098 (N_2098,N_856,N_1433);
and U2099 (N_2099,N_1154,N_1311);
and U2100 (N_2100,N_975,N_1180);
nand U2101 (N_2101,N_1262,N_956);
nand U2102 (N_2102,N_970,N_1206);
nor U2103 (N_2103,N_1021,N_1195);
nor U2104 (N_2104,N_923,N_1565);
xnor U2105 (N_2105,N_1534,N_1541);
or U2106 (N_2106,N_909,N_839);
or U2107 (N_2107,N_867,N_1324);
nand U2108 (N_2108,N_1549,N_1272);
nand U2109 (N_2109,N_1567,N_1297);
or U2110 (N_2110,N_830,N_1371);
xnor U2111 (N_2111,N_1120,N_1343);
nand U2112 (N_2112,N_1467,N_1165);
nand U2113 (N_2113,N_993,N_936);
nor U2114 (N_2114,N_1484,N_1231);
or U2115 (N_2115,N_1327,N_1563);
xor U2116 (N_2116,N_1236,N_1291);
nand U2117 (N_2117,N_1308,N_806);
and U2118 (N_2118,N_1476,N_1253);
xnor U2119 (N_2119,N_1352,N_1521);
xor U2120 (N_2120,N_1478,N_1341);
or U2121 (N_2121,N_1004,N_1349);
nor U2122 (N_2122,N_1214,N_839);
nand U2123 (N_2123,N_806,N_1054);
xnor U2124 (N_2124,N_1423,N_1000);
nand U2125 (N_2125,N_1041,N_1157);
nor U2126 (N_2126,N_1258,N_1502);
nand U2127 (N_2127,N_1320,N_953);
xnor U2128 (N_2128,N_1004,N_1042);
xor U2129 (N_2129,N_1291,N_1527);
and U2130 (N_2130,N_1400,N_1359);
xnor U2131 (N_2131,N_1203,N_1303);
nor U2132 (N_2132,N_1043,N_861);
xor U2133 (N_2133,N_1218,N_1246);
and U2134 (N_2134,N_1116,N_865);
or U2135 (N_2135,N_1381,N_1150);
xor U2136 (N_2136,N_1009,N_1126);
nor U2137 (N_2137,N_1301,N_1041);
xor U2138 (N_2138,N_992,N_949);
nand U2139 (N_2139,N_1065,N_1532);
nor U2140 (N_2140,N_1533,N_964);
xor U2141 (N_2141,N_1309,N_1142);
xnor U2142 (N_2142,N_1434,N_984);
or U2143 (N_2143,N_1540,N_989);
nand U2144 (N_2144,N_903,N_1190);
and U2145 (N_2145,N_1539,N_964);
and U2146 (N_2146,N_1391,N_1195);
nor U2147 (N_2147,N_1548,N_847);
and U2148 (N_2148,N_871,N_1232);
nor U2149 (N_2149,N_1273,N_978);
xor U2150 (N_2150,N_916,N_1505);
xor U2151 (N_2151,N_1510,N_1128);
nor U2152 (N_2152,N_873,N_828);
nand U2153 (N_2153,N_1507,N_1435);
or U2154 (N_2154,N_1251,N_1395);
xor U2155 (N_2155,N_1157,N_1092);
xnor U2156 (N_2156,N_1093,N_880);
nand U2157 (N_2157,N_1059,N_1484);
and U2158 (N_2158,N_1005,N_844);
or U2159 (N_2159,N_1050,N_1085);
and U2160 (N_2160,N_1469,N_1543);
or U2161 (N_2161,N_1455,N_1224);
nor U2162 (N_2162,N_903,N_867);
nand U2163 (N_2163,N_1228,N_1550);
and U2164 (N_2164,N_1462,N_1582);
nor U2165 (N_2165,N_1353,N_1078);
and U2166 (N_2166,N_1047,N_951);
xnor U2167 (N_2167,N_927,N_1181);
and U2168 (N_2168,N_1177,N_1113);
nor U2169 (N_2169,N_1004,N_1065);
nor U2170 (N_2170,N_1120,N_1529);
nand U2171 (N_2171,N_1471,N_1135);
nand U2172 (N_2172,N_1422,N_1302);
nand U2173 (N_2173,N_1404,N_1332);
or U2174 (N_2174,N_1382,N_869);
and U2175 (N_2175,N_1049,N_1524);
and U2176 (N_2176,N_1047,N_1235);
or U2177 (N_2177,N_1393,N_1306);
nor U2178 (N_2178,N_1030,N_1545);
xor U2179 (N_2179,N_888,N_1584);
nand U2180 (N_2180,N_1381,N_972);
nand U2181 (N_2181,N_1115,N_974);
xnor U2182 (N_2182,N_980,N_971);
nor U2183 (N_2183,N_1459,N_1101);
nor U2184 (N_2184,N_1528,N_1305);
or U2185 (N_2185,N_1213,N_1513);
and U2186 (N_2186,N_1572,N_1460);
nor U2187 (N_2187,N_1149,N_889);
nand U2188 (N_2188,N_1028,N_1065);
or U2189 (N_2189,N_896,N_1129);
xor U2190 (N_2190,N_1400,N_1014);
nor U2191 (N_2191,N_1301,N_888);
nor U2192 (N_2192,N_1038,N_1065);
and U2193 (N_2193,N_1287,N_1078);
nand U2194 (N_2194,N_1187,N_1490);
or U2195 (N_2195,N_817,N_1270);
xor U2196 (N_2196,N_1353,N_965);
and U2197 (N_2197,N_1252,N_1123);
xor U2198 (N_2198,N_1346,N_1007);
nand U2199 (N_2199,N_1219,N_1212);
and U2200 (N_2200,N_1396,N_1554);
nand U2201 (N_2201,N_1251,N_924);
nand U2202 (N_2202,N_1554,N_985);
nor U2203 (N_2203,N_1429,N_1027);
nor U2204 (N_2204,N_944,N_1563);
nand U2205 (N_2205,N_1100,N_814);
nand U2206 (N_2206,N_1266,N_883);
or U2207 (N_2207,N_1457,N_1410);
nor U2208 (N_2208,N_887,N_936);
nor U2209 (N_2209,N_961,N_1122);
and U2210 (N_2210,N_1099,N_1575);
xnor U2211 (N_2211,N_1230,N_1486);
nand U2212 (N_2212,N_906,N_809);
or U2213 (N_2213,N_1449,N_1566);
xnor U2214 (N_2214,N_942,N_1065);
and U2215 (N_2215,N_1260,N_989);
xnor U2216 (N_2216,N_1146,N_1520);
and U2217 (N_2217,N_1515,N_836);
nand U2218 (N_2218,N_1339,N_972);
nand U2219 (N_2219,N_1188,N_1298);
and U2220 (N_2220,N_1238,N_1347);
nor U2221 (N_2221,N_1400,N_1267);
nor U2222 (N_2222,N_907,N_1213);
or U2223 (N_2223,N_1240,N_903);
or U2224 (N_2224,N_874,N_1564);
nor U2225 (N_2225,N_1021,N_1225);
nor U2226 (N_2226,N_903,N_1468);
or U2227 (N_2227,N_1129,N_1306);
xor U2228 (N_2228,N_1013,N_996);
or U2229 (N_2229,N_859,N_1394);
nand U2230 (N_2230,N_931,N_1192);
and U2231 (N_2231,N_908,N_1348);
nor U2232 (N_2232,N_910,N_1218);
and U2233 (N_2233,N_1070,N_1034);
or U2234 (N_2234,N_848,N_1490);
xor U2235 (N_2235,N_1394,N_1578);
xnor U2236 (N_2236,N_1256,N_890);
xnor U2237 (N_2237,N_847,N_919);
nand U2238 (N_2238,N_1346,N_1311);
xor U2239 (N_2239,N_986,N_861);
xnor U2240 (N_2240,N_1223,N_1330);
nor U2241 (N_2241,N_1592,N_1426);
and U2242 (N_2242,N_1504,N_1239);
and U2243 (N_2243,N_910,N_973);
and U2244 (N_2244,N_1436,N_1253);
and U2245 (N_2245,N_1090,N_1057);
xor U2246 (N_2246,N_1388,N_1286);
xor U2247 (N_2247,N_1347,N_1305);
or U2248 (N_2248,N_1228,N_941);
and U2249 (N_2249,N_1483,N_1364);
and U2250 (N_2250,N_1386,N_964);
nand U2251 (N_2251,N_1508,N_1483);
nor U2252 (N_2252,N_1080,N_1142);
or U2253 (N_2253,N_968,N_1213);
nand U2254 (N_2254,N_1321,N_1476);
and U2255 (N_2255,N_1390,N_948);
nor U2256 (N_2256,N_1040,N_1568);
or U2257 (N_2257,N_1453,N_1324);
xor U2258 (N_2258,N_941,N_1518);
xor U2259 (N_2259,N_1462,N_1424);
and U2260 (N_2260,N_1548,N_802);
and U2261 (N_2261,N_1460,N_1077);
xnor U2262 (N_2262,N_817,N_1292);
nor U2263 (N_2263,N_1163,N_887);
nand U2264 (N_2264,N_1013,N_880);
or U2265 (N_2265,N_1238,N_1458);
or U2266 (N_2266,N_830,N_1142);
nand U2267 (N_2267,N_993,N_1237);
or U2268 (N_2268,N_1505,N_1033);
or U2269 (N_2269,N_1032,N_905);
or U2270 (N_2270,N_1070,N_884);
or U2271 (N_2271,N_1434,N_895);
and U2272 (N_2272,N_1086,N_836);
xor U2273 (N_2273,N_1248,N_1020);
nor U2274 (N_2274,N_1072,N_1057);
nor U2275 (N_2275,N_1037,N_1066);
xnor U2276 (N_2276,N_1323,N_1293);
nand U2277 (N_2277,N_1539,N_887);
nand U2278 (N_2278,N_1511,N_958);
or U2279 (N_2279,N_1581,N_831);
and U2280 (N_2280,N_922,N_1039);
or U2281 (N_2281,N_1242,N_1571);
and U2282 (N_2282,N_1091,N_1386);
xor U2283 (N_2283,N_964,N_1403);
or U2284 (N_2284,N_928,N_1278);
nand U2285 (N_2285,N_1425,N_1210);
or U2286 (N_2286,N_1438,N_1578);
and U2287 (N_2287,N_1234,N_1164);
nand U2288 (N_2288,N_967,N_1521);
nand U2289 (N_2289,N_980,N_863);
nor U2290 (N_2290,N_1146,N_1334);
or U2291 (N_2291,N_950,N_1054);
xor U2292 (N_2292,N_1391,N_1315);
and U2293 (N_2293,N_1578,N_885);
or U2294 (N_2294,N_1186,N_1094);
xor U2295 (N_2295,N_1580,N_1093);
or U2296 (N_2296,N_969,N_1308);
nand U2297 (N_2297,N_1268,N_856);
and U2298 (N_2298,N_1250,N_1040);
nor U2299 (N_2299,N_1577,N_1359);
nor U2300 (N_2300,N_1272,N_1050);
and U2301 (N_2301,N_1498,N_1066);
xnor U2302 (N_2302,N_1214,N_1056);
or U2303 (N_2303,N_1521,N_1121);
nand U2304 (N_2304,N_1418,N_1282);
nand U2305 (N_2305,N_897,N_1192);
nand U2306 (N_2306,N_1440,N_887);
nand U2307 (N_2307,N_1243,N_1395);
and U2308 (N_2308,N_1040,N_1062);
xor U2309 (N_2309,N_901,N_920);
nand U2310 (N_2310,N_1163,N_1298);
xnor U2311 (N_2311,N_1451,N_1070);
xnor U2312 (N_2312,N_1402,N_1554);
nor U2313 (N_2313,N_1287,N_894);
or U2314 (N_2314,N_1512,N_1319);
and U2315 (N_2315,N_873,N_1071);
nor U2316 (N_2316,N_1120,N_1373);
nand U2317 (N_2317,N_1486,N_1146);
and U2318 (N_2318,N_1175,N_998);
nand U2319 (N_2319,N_1113,N_1267);
nand U2320 (N_2320,N_927,N_1424);
xnor U2321 (N_2321,N_1294,N_849);
and U2322 (N_2322,N_1287,N_1262);
nor U2323 (N_2323,N_1325,N_951);
nand U2324 (N_2324,N_1408,N_1214);
or U2325 (N_2325,N_1049,N_918);
and U2326 (N_2326,N_1422,N_1115);
or U2327 (N_2327,N_1365,N_1240);
and U2328 (N_2328,N_951,N_1090);
or U2329 (N_2329,N_1223,N_1109);
and U2330 (N_2330,N_1441,N_1352);
and U2331 (N_2331,N_1033,N_1238);
nand U2332 (N_2332,N_1412,N_1334);
or U2333 (N_2333,N_1044,N_1302);
nor U2334 (N_2334,N_869,N_1287);
or U2335 (N_2335,N_1372,N_940);
xnor U2336 (N_2336,N_1051,N_1122);
xnor U2337 (N_2337,N_1092,N_1579);
and U2338 (N_2338,N_1591,N_1100);
and U2339 (N_2339,N_1584,N_901);
and U2340 (N_2340,N_1342,N_1473);
nor U2341 (N_2341,N_1350,N_1367);
nor U2342 (N_2342,N_1120,N_978);
or U2343 (N_2343,N_1323,N_845);
or U2344 (N_2344,N_1585,N_1517);
or U2345 (N_2345,N_1071,N_1343);
nand U2346 (N_2346,N_1497,N_1546);
and U2347 (N_2347,N_955,N_1364);
or U2348 (N_2348,N_1410,N_1518);
xnor U2349 (N_2349,N_1578,N_1351);
or U2350 (N_2350,N_1144,N_1041);
nor U2351 (N_2351,N_1053,N_896);
nand U2352 (N_2352,N_1150,N_1102);
nor U2353 (N_2353,N_1331,N_1423);
xnor U2354 (N_2354,N_1130,N_1419);
nor U2355 (N_2355,N_1534,N_1495);
nand U2356 (N_2356,N_1565,N_1142);
xnor U2357 (N_2357,N_1194,N_1377);
nor U2358 (N_2358,N_1458,N_872);
xnor U2359 (N_2359,N_907,N_1300);
or U2360 (N_2360,N_853,N_1289);
and U2361 (N_2361,N_1280,N_1357);
and U2362 (N_2362,N_1193,N_1417);
or U2363 (N_2363,N_1224,N_915);
nor U2364 (N_2364,N_1418,N_939);
nor U2365 (N_2365,N_1584,N_1536);
nor U2366 (N_2366,N_1492,N_1079);
and U2367 (N_2367,N_1020,N_1312);
xnor U2368 (N_2368,N_1547,N_953);
nand U2369 (N_2369,N_1348,N_1565);
xnor U2370 (N_2370,N_1045,N_1439);
nand U2371 (N_2371,N_1214,N_882);
nor U2372 (N_2372,N_1051,N_1228);
and U2373 (N_2373,N_1116,N_1171);
xor U2374 (N_2374,N_870,N_1018);
nand U2375 (N_2375,N_1150,N_1174);
and U2376 (N_2376,N_1068,N_862);
nand U2377 (N_2377,N_1160,N_873);
nor U2378 (N_2378,N_1453,N_1488);
and U2379 (N_2379,N_1596,N_1119);
or U2380 (N_2380,N_1276,N_964);
xor U2381 (N_2381,N_1596,N_995);
nand U2382 (N_2382,N_1379,N_1584);
or U2383 (N_2383,N_813,N_1393);
xnor U2384 (N_2384,N_1225,N_1396);
xor U2385 (N_2385,N_1136,N_809);
nand U2386 (N_2386,N_1046,N_838);
nand U2387 (N_2387,N_885,N_1314);
nor U2388 (N_2388,N_1419,N_1157);
and U2389 (N_2389,N_803,N_1573);
and U2390 (N_2390,N_1131,N_1360);
nand U2391 (N_2391,N_1184,N_1049);
and U2392 (N_2392,N_888,N_1434);
or U2393 (N_2393,N_1253,N_1046);
nor U2394 (N_2394,N_1313,N_891);
and U2395 (N_2395,N_1259,N_1597);
nand U2396 (N_2396,N_805,N_1107);
nand U2397 (N_2397,N_1339,N_1051);
and U2398 (N_2398,N_994,N_1258);
or U2399 (N_2399,N_901,N_827);
nor U2400 (N_2400,N_1961,N_2218);
nand U2401 (N_2401,N_1867,N_1635);
or U2402 (N_2402,N_1841,N_2310);
nand U2403 (N_2403,N_1860,N_1825);
nand U2404 (N_2404,N_1744,N_2240);
nor U2405 (N_2405,N_1763,N_1950);
nand U2406 (N_2406,N_1812,N_1994);
nor U2407 (N_2407,N_2050,N_1944);
or U2408 (N_2408,N_1746,N_2217);
nor U2409 (N_2409,N_1875,N_1956);
and U2410 (N_2410,N_1965,N_2270);
or U2411 (N_2411,N_2332,N_1690);
xnor U2412 (N_2412,N_1783,N_1991);
nand U2413 (N_2413,N_1854,N_1692);
xnor U2414 (N_2414,N_1630,N_2047);
nand U2415 (N_2415,N_2336,N_2243);
nor U2416 (N_2416,N_1925,N_1805);
nand U2417 (N_2417,N_1636,N_1664);
and U2418 (N_2418,N_2251,N_1884);
nor U2419 (N_2419,N_2343,N_2358);
nor U2420 (N_2420,N_2054,N_2271);
xor U2421 (N_2421,N_2290,N_1703);
nor U2422 (N_2422,N_1622,N_2393);
or U2423 (N_2423,N_1959,N_1842);
or U2424 (N_2424,N_1643,N_2394);
xor U2425 (N_2425,N_1649,N_1935);
xnor U2426 (N_2426,N_1928,N_2044);
nand U2427 (N_2427,N_1730,N_1981);
xnor U2428 (N_2428,N_1696,N_1788);
xnor U2429 (N_2429,N_1702,N_1764);
nor U2430 (N_2430,N_1918,N_1762);
nor U2431 (N_2431,N_1971,N_2201);
or U2432 (N_2432,N_2179,N_1931);
and U2433 (N_2433,N_1992,N_2286);
xor U2434 (N_2434,N_1821,N_1851);
and U2435 (N_2435,N_2184,N_1939);
xor U2436 (N_2436,N_2162,N_2022);
and U2437 (N_2437,N_2362,N_2302);
nor U2438 (N_2438,N_2386,N_1794);
xnor U2439 (N_2439,N_2320,N_2357);
or U2440 (N_2440,N_2204,N_1914);
xnor U2441 (N_2441,N_1778,N_2387);
nor U2442 (N_2442,N_2331,N_1653);
nor U2443 (N_2443,N_2323,N_1648);
nor U2444 (N_2444,N_1849,N_2152);
and U2445 (N_2445,N_1732,N_2131);
xnor U2446 (N_2446,N_2113,N_1674);
xnor U2447 (N_2447,N_1632,N_1752);
xnor U2448 (N_2448,N_2074,N_1930);
nand U2449 (N_2449,N_2057,N_2288);
nor U2450 (N_2450,N_1745,N_2071);
xor U2451 (N_2451,N_2158,N_2212);
or U2452 (N_2452,N_1739,N_2134);
nor U2453 (N_2453,N_1819,N_2335);
and U2454 (N_2454,N_1657,N_1640);
xor U2455 (N_2455,N_1892,N_2304);
nor U2456 (N_2456,N_2368,N_1682);
nor U2457 (N_2457,N_2048,N_2367);
and U2458 (N_2458,N_1871,N_1617);
nor U2459 (N_2459,N_2051,N_2155);
and U2460 (N_2460,N_1665,N_2352);
and U2461 (N_2461,N_2116,N_1968);
and U2462 (N_2462,N_1853,N_2333);
and U2463 (N_2463,N_2282,N_1877);
nand U2464 (N_2464,N_1896,N_2062);
or U2465 (N_2465,N_2183,N_2385);
and U2466 (N_2466,N_1986,N_1796);
nor U2467 (N_2467,N_1618,N_1667);
nand U2468 (N_2468,N_2366,N_2244);
nand U2469 (N_2469,N_2127,N_2058);
nand U2470 (N_2470,N_2287,N_1684);
and U2471 (N_2471,N_1862,N_2000);
nor U2472 (N_2472,N_2164,N_1721);
xor U2473 (N_2473,N_1737,N_2225);
or U2474 (N_2474,N_2242,N_1609);
and U2475 (N_2475,N_2035,N_1698);
nor U2476 (N_2476,N_2137,N_2149);
nand U2477 (N_2477,N_1814,N_2086);
nand U2478 (N_2478,N_2095,N_2019);
and U2479 (N_2479,N_1754,N_2125);
xnor U2480 (N_2480,N_2147,N_2023);
nor U2481 (N_2481,N_1685,N_1772);
or U2482 (N_2482,N_1834,N_1779);
xnor U2483 (N_2483,N_2001,N_2031);
and U2484 (N_2484,N_2092,N_2206);
nor U2485 (N_2485,N_2009,N_1999);
or U2486 (N_2486,N_2325,N_1985);
or U2487 (N_2487,N_2205,N_2021);
nor U2488 (N_2488,N_1908,N_2289);
and U2489 (N_2489,N_2375,N_1786);
and U2490 (N_2490,N_2055,N_2075);
and U2491 (N_2491,N_2042,N_2157);
and U2492 (N_2492,N_2292,N_2046);
or U2493 (N_2493,N_2254,N_1839);
and U2494 (N_2494,N_1680,N_1784);
or U2495 (N_2495,N_2117,N_2033);
and U2496 (N_2496,N_1962,N_1937);
xnor U2497 (N_2497,N_2061,N_1615);
xnor U2498 (N_2498,N_2284,N_1611);
nor U2499 (N_2499,N_2052,N_1824);
or U2500 (N_2500,N_1888,N_2199);
and U2501 (N_2501,N_1700,N_2169);
or U2502 (N_2502,N_2280,N_2353);
nor U2503 (N_2503,N_2166,N_1910);
nand U2504 (N_2504,N_2148,N_2102);
xor U2505 (N_2505,N_1946,N_2014);
nor U2506 (N_2506,N_2040,N_1738);
and U2507 (N_2507,N_2180,N_2010);
or U2508 (N_2508,N_1624,N_2161);
nand U2509 (N_2509,N_1610,N_2049);
nor U2510 (N_2510,N_1952,N_2070);
xnor U2511 (N_2511,N_1977,N_1942);
and U2512 (N_2512,N_1616,N_1826);
and U2513 (N_2513,N_2322,N_1974);
xnor U2514 (N_2514,N_2235,N_1715);
nand U2515 (N_2515,N_2239,N_2344);
nand U2516 (N_2516,N_2281,N_2297);
nand U2517 (N_2517,N_1614,N_2296);
nor U2518 (N_2518,N_1724,N_2099);
nand U2519 (N_2519,N_2027,N_2112);
and U2520 (N_2520,N_2312,N_2246);
and U2521 (N_2521,N_1912,N_1829);
xor U2522 (N_2522,N_1642,N_1727);
nor U2523 (N_2523,N_1602,N_2255);
nor U2524 (N_2524,N_2136,N_1921);
nand U2525 (N_2525,N_2265,N_2156);
or U2526 (N_2526,N_1874,N_2278);
or U2527 (N_2527,N_2274,N_2256);
or U2528 (N_2528,N_1883,N_1911);
xnor U2529 (N_2529,N_1701,N_2091);
nor U2530 (N_2530,N_1924,N_2233);
nand U2531 (N_2531,N_2364,N_2305);
nor U2532 (N_2532,N_1756,N_2203);
xor U2533 (N_2533,N_1673,N_2309);
or U2534 (N_2534,N_2030,N_2337);
xor U2535 (N_2535,N_2151,N_2372);
xnor U2536 (N_2536,N_2143,N_1634);
xor U2537 (N_2537,N_2346,N_1964);
nand U2538 (N_2538,N_1646,N_2196);
xnor U2539 (N_2539,N_2163,N_1975);
and U2540 (N_2540,N_2324,N_2081);
xor U2541 (N_2541,N_2124,N_2090);
xnor U2542 (N_2542,N_1933,N_2038);
and U2543 (N_2543,N_2359,N_1857);
nand U2544 (N_2544,N_2083,N_1720);
nor U2545 (N_2545,N_1781,N_2089);
or U2546 (N_2546,N_1706,N_1856);
xnor U2547 (N_2547,N_2024,N_2041);
or U2548 (N_2548,N_2094,N_1855);
xor U2549 (N_2549,N_1887,N_1936);
and U2550 (N_2550,N_1714,N_1947);
and U2551 (N_2551,N_2017,N_1980);
xor U2552 (N_2552,N_1929,N_1852);
xor U2553 (N_2553,N_1775,N_2029);
and U2554 (N_2554,N_2300,N_1903);
and U2555 (N_2555,N_2214,N_2069);
nand U2556 (N_2556,N_1963,N_1750);
nand U2557 (N_2557,N_1713,N_2252);
nand U2558 (N_2558,N_1861,N_1807);
nand U2559 (N_2559,N_1656,N_1777);
nor U2560 (N_2560,N_1880,N_1827);
or U2561 (N_2561,N_2347,N_2178);
xor U2562 (N_2562,N_2084,N_1718);
or U2563 (N_2563,N_1920,N_2108);
and U2564 (N_2564,N_1916,N_2032);
nand U2565 (N_2565,N_2327,N_2228);
nand U2566 (N_2566,N_1889,N_2103);
nand U2567 (N_2567,N_2221,N_2341);
xnor U2568 (N_2568,N_1662,N_1678);
nand U2569 (N_2569,N_1726,N_2007);
nand U2570 (N_2570,N_1976,N_2260);
nand U2571 (N_2571,N_1832,N_2096);
xnor U2572 (N_2572,N_1753,N_2130);
or U2573 (N_2573,N_1709,N_2340);
or U2574 (N_2574,N_2053,N_2195);
nand U2575 (N_2575,N_2187,N_2261);
and U2576 (N_2576,N_1785,N_1913);
nand U2577 (N_2577,N_2238,N_2115);
nand U2578 (N_2578,N_2060,N_1719);
and U2579 (N_2579,N_2371,N_1633);
xnor U2580 (N_2580,N_2277,N_1603);
and U2581 (N_2581,N_2085,N_1716);
or U2582 (N_2582,N_1945,N_1865);
and U2583 (N_2583,N_1661,N_1847);
or U2584 (N_2584,N_1978,N_1943);
xor U2585 (N_2585,N_2082,N_1987);
nand U2586 (N_2586,N_2273,N_2349);
or U2587 (N_2587,N_1787,N_1810);
xnor U2588 (N_2588,N_1631,N_1881);
nand U2589 (N_2589,N_2330,N_1795);
nor U2590 (N_2590,N_2128,N_2208);
nor U2591 (N_2591,N_1802,N_1932);
xor U2592 (N_2592,N_2381,N_2043);
xnor U2593 (N_2593,N_2307,N_2230);
or U2594 (N_2594,N_2384,N_2391);
xnor U2595 (N_2595,N_2272,N_2259);
xnor U2596 (N_2596,N_2220,N_2306);
nor U2597 (N_2597,N_1792,N_1679);
nand U2598 (N_2598,N_2068,N_1808);
nor U2599 (N_2599,N_2174,N_2018);
or U2600 (N_2600,N_2293,N_1647);
nor U2601 (N_2601,N_1793,N_2185);
or U2602 (N_2602,N_1809,N_2093);
nor U2603 (N_2603,N_2073,N_2379);
and U2604 (N_2604,N_1815,N_1972);
nor U2605 (N_2605,N_1823,N_1740);
or U2606 (N_2606,N_2173,N_1686);
or U2607 (N_2607,N_2175,N_1695);
nor U2608 (N_2608,N_1704,N_2295);
xnor U2609 (N_2609,N_1863,N_1604);
or U2610 (N_2610,N_1958,N_1837);
nor U2611 (N_2611,N_2192,N_2126);
nand U2612 (N_2612,N_1765,N_2241);
xnor U2613 (N_2613,N_2129,N_2299);
xnor U2614 (N_2614,N_2186,N_2361);
nand U2615 (N_2615,N_1607,N_2382);
or U2616 (N_2616,N_2076,N_2026);
and U2617 (N_2617,N_1866,N_1890);
or U2618 (N_2618,N_2170,N_1669);
or U2619 (N_2619,N_2020,N_1940);
nor U2620 (N_2620,N_1905,N_1687);
or U2621 (N_2621,N_2015,N_1651);
and U2622 (N_2622,N_2249,N_2168);
and U2623 (N_2623,N_2013,N_2308);
xor U2624 (N_2624,N_1899,N_2006);
xor U2625 (N_2625,N_2266,N_2059);
or U2626 (N_2626,N_1743,N_1758);
xor U2627 (N_2627,N_2121,N_2189);
nor U2628 (N_2628,N_1897,N_2248);
nor U2629 (N_2629,N_1782,N_1670);
nor U2630 (N_2630,N_2236,N_1838);
xor U2631 (N_2631,N_1878,N_2350);
or U2632 (N_2632,N_1938,N_1844);
and U2633 (N_2633,N_2104,N_2224);
nor U2634 (N_2634,N_2373,N_1710);
xor U2635 (N_2635,N_2219,N_2165);
xnor U2636 (N_2636,N_2097,N_2245);
nor U2637 (N_2637,N_2153,N_1953);
nor U2638 (N_2638,N_2338,N_1858);
nor U2639 (N_2639,N_1922,N_1605);
nor U2640 (N_2640,N_1663,N_1659);
or U2641 (N_2641,N_2025,N_2313);
nor U2642 (N_2642,N_1791,N_2159);
xnor U2643 (N_2643,N_1728,N_1731);
and U2644 (N_2644,N_2231,N_1689);
nand U2645 (N_2645,N_2138,N_2144);
and U2646 (N_2646,N_1749,N_2374);
nor U2647 (N_2647,N_2388,N_2037);
and U2648 (N_2648,N_1742,N_1818);
xnor U2649 (N_2649,N_2182,N_1898);
and U2650 (N_2650,N_2321,N_2264);
nand U2651 (N_2651,N_1906,N_1934);
nand U2652 (N_2652,N_1672,N_1900);
nand U2653 (N_2653,N_1723,N_2045);
nor U2654 (N_2654,N_1612,N_1629);
xnor U2655 (N_2655,N_2122,N_1660);
and U2656 (N_2656,N_2016,N_2363);
nand U2657 (N_2657,N_2279,N_1820);
or U2658 (N_2658,N_1893,N_1813);
or U2659 (N_2659,N_1748,N_2263);
or U2660 (N_2660,N_1627,N_1641);
or U2661 (N_2661,N_2298,N_2355);
nor U2662 (N_2662,N_1904,N_1666);
nor U2663 (N_2663,N_1652,N_1619);
xnor U2664 (N_2664,N_1736,N_1828);
or U2665 (N_2665,N_2190,N_2109);
nor U2666 (N_2666,N_1966,N_1869);
nand U2667 (N_2667,N_2188,N_2399);
nand U2668 (N_2668,N_2039,N_1768);
xnor U2669 (N_2669,N_1850,N_1955);
xnor U2670 (N_2670,N_2120,N_2319);
nand U2671 (N_2671,N_2334,N_2193);
or U2672 (N_2672,N_1683,N_2234);
or U2673 (N_2673,N_2088,N_2067);
and U2674 (N_2674,N_1891,N_1606);
and U2675 (N_2675,N_2326,N_2145);
or U2676 (N_2676,N_1804,N_1915);
nand U2677 (N_2677,N_2257,N_1835);
or U2678 (N_2678,N_1747,N_1846);
nand U2679 (N_2679,N_2114,N_2118);
xor U2680 (N_2680,N_2198,N_2395);
nor U2681 (N_2681,N_2253,N_2133);
or U2682 (N_2682,N_1873,N_2197);
nor U2683 (N_2683,N_2191,N_2100);
and U2684 (N_2684,N_1620,N_2028);
xor U2685 (N_2685,N_2285,N_1801);
xor U2686 (N_2686,N_1725,N_1822);
and U2687 (N_2687,N_2369,N_1717);
xor U2688 (N_2688,N_1995,N_2316);
nand U2689 (N_2689,N_2329,N_2398);
nor U2690 (N_2690,N_1840,N_2140);
nor U2691 (N_2691,N_2002,N_1879);
and U2692 (N_2692,N_2247,N_1637);
nor U2693 (N_2693,N_1859,N_2167);
or U2694 (N_2694,N_1876,N_1623);
nand U2695 (N_2695,N_2150,N_2004);
xor U2696 (N_2696,N_1771,N_1761);
xnor U2697 (N_2697,N_1848,N_1712);
or U2698 (N_2698,N_2063,N_1766);
or U2699 (N_2699,N_2011,N_2079);
nand U2700 (N_2700,N_2301,N_2200);
xor U2701 (N_2701,N_1733,N_1677);
and U2702 (N_2702,N_2080,N_1885);
or U2703 (N_2703,N_2276,N_1895);
nor U2704 (N_2704,N_1694,N_2132);
nor U2705 (N_2705,N_1969,N_2003);
nor U2706 (N_2706,N_1811,N_1836);
xor U2707 (N_2707,N_2262,N_1601);
nand U2708 (N_2708,N_1691,N_2356);
or U2709 (N_2709,N_1886,N_1676);
nor U2710 (N_2710,N_1982,N_2077);
and U2711 (N_2711,N_2211,N_2345);
nor U2712 (N_2712,N_1996,N_2232);
xnor U2713 (N_2713,N_2227,N_1997);
nand U2714 (N_2714,N_2226,N_1927);
nor U2715 (N_2715,N_2268,N_1806);
nand U2716 (N_2716,N_1845,N_2267);
xor U2717 (N_2717,N_2348,N_2056);
nor U2718 (N_2718,N_2107,N_1882);
or U2719 (N_2719,N_2223,N_1957);
or U2720 (N_2720,N_1989,N_2171);
and U2721 (N_2721,N_1917,N_2065);
xor U2722 (N_2722,N_1780,N_1960);
nand U2723 (N_2723,N_1799,N_1751);
nand U2724 (N_2724,N_1800,N_2111);
or U2725 (N_2725,N_1625,N_1868);
and U2726 (N_2726,N_2177,N_1954);
or U2727 (N_2727,N_2202,N_2314);
nand U2728 (N_2728,N_1708,N_2119);
or U2729 (N_2729,N_1755,N_2318);
xnor U2730 (N_2730,N_2008,N_1655);
or U2731 (N_2731,N_2106,N_1901);
nand U2732 (N_2732,N_2383,N_1833);
nor U2733 (N_2733,N_2380,N_1843);
and U2734 (N_2734,N_1872,N_1613);
nand U2735 (N_2735,N_2250,N_1681);
xor U2736 (N_2736,N_1711,N_1639);
nand U2737 (N_2737,N_2339,N_2378);
or U2738 (N_2738,N_1949,N_2370);
and U2739 (N_2739,N_1817,N_1688);
and U2740 (N_2740,N_1628,N_1990);
nor U2741 (N_2741,N_1816,N_2354);
xor U2742 (N_2742,N_1645,N_1870);
nor U2743 (N_2743,N_1759,N_1948);
nor U2744 (N_2744,N_2283,N_2105);
or U2745 (N_2745,N_2160,N_1830);
nand U2746 (N_2746,N_2389,N_1769);
nor U2747 (N_2747,N_2181,N_2229);
xor U2748 (N_2748,N_2139,N_2172);
xnor U2749 (N_2749,N_1675,N_2216);
and U2750 (N_2750,N_1773,N_1638);
nand U2751 (N_2751,N_1626,N_2064);
and U2752 (N_2752,N_1650,N_1729);
nor U2753 (N_2753,N_2154,N_2209);
and U2754 (N_2754,N_1983,N_1988);
nand U2755 (N_2755,N_1797,N_1697);
nor U2756 (N_2756,N_2377,N_2101);
nor U2757 (N_2757,N_1998,N_2258);
nor U2758 (N_2758,N_2237,N_2360);
nor U2759 (N_2759,N_2005,N_1671);
nand U2760 (N_2760,N_1790,N_1926);
xnor U2761 (N_2761,N_2135,N_1774);
or U2762 (N_2762,N_1621,N_1707);
xor U2763 (N_2763,N_1668,N_2034);
nor U2764 (N_2764,N_1979,N_1984);
nand U2765 (N_2765,N_1658,N_1970);
nor U2766 (N_2766,N_1741,N_1907);
or U2767 (N_2767,N_2142,N_1776);
nand U2768 (N_2768,N_1967,N_2123);
nand U2769 (N_2769,N_2275,N_2351);
xor U2770 (N_2770,N_2365,N_1864);
nor U2771 (N_2771,N_1654,N_2210);
nor U2772 (N_2772,N_1789,N_1803);
or U2773 (N_2773,N_2303,N_1798);
and U2774 (N_2774,N_1923,N_2397);
and U2775 (N_2775,N_2207,N_1902);
nand U2776 (N_2776,N_2146,N_2194);
xor U2777 (N_2777,N_2294,N_1760);
or U2778 (N_2778,N_2012,N_2317);
or U2779 (N_2779,N_1894,N_1734);
and U2780 (N_2780,N_2098,N_1767);
nor U2781 (N_2781,N_1600,N_1993);
or U2782 (N_2782,N_1705,N_2396);
xor U2783 (N_2783,N_2110,N_2222);
or U2784 (N_2784,N_2215,N_2311);
xnor U2785 (N_2785,N_1770,N_2315);
and U2786 (N_2786,N_1644,N_2072);
or U2787 (N_2787,N_1757,N_1941);
nor U2788 (N_2788,N_1951,N_1919);
or U2789 (N_2789,N_1831,N_2066);
nor U2790 (N_2790,N_2269,N_2291);
and U2791 (N_2791,N_1699,N_2176);
xnor U2792 (N_2792,N_2390,N_2213);
and U2793 (N_2793,N_1909,N_2078);
xnor U2794 (N_2794,N_1722,N_1735);
and U2795 (N_2795,N_2376,N_1693);
and U2796 (N_2796,N_2036,N_2141);
or U2797 (N_2797,N_1608,N_2087);
nand U2798 (N_2798,N_2392,N_2328);
and U2799 (N_2799,N_2342,N_1973);
nor U2800 (N_2800,N_2281,N_2089);
nand U2801 (N_2801,N_2090,N_1625);
nor U2802 (N_2802,N_2330,N_2219);
or U2803 (N_2803,N_1672,N_1881);
xnor U2804 (N_2804,N_2325,N_2276);
xnor U2805 (N_2805,N_2033,N_2045);
or U2806 (N_2806,N_2387,N_2256);
or U2807 (N_2807,N_2062,N_2256);
nor U2808 (N_2808,N_1717,N_2009);
and U2809 (N_2809,N_2390,N_2250);
or U2810 (N_2810,N_2309,N_2386);
and U2811 (N_2811,N_1712,N_1900);
nor U2812 (N_2812,N_2366,N_1979);
xor U2813 (N_2813,N_2395,N_2144);
nor U2814 (N_2814,N_1873,N_2139);
nand U2815 (N_2815,N_2190,N_1619);
nor U2816 (N_2816,N_1886,N_2150);
xnor U2817 (N_2817,N_2153,N_2385);
nor U2818 (N_2818,N_2317,N_2088);
xor U2819 (N_2819,N_2188,N_1774);
xnor U2820 (N_2820,N_1711,N_1920);
nand U2821 (N_2821,N_2236,N_2314);
or U2822 (N_2822,N_2211,N_1826);
or U2823 (N_2823,N_1690,N_2083);
or U2824 (N_2824,N_2249,N_2050);
nand U2825 (N_2825,N_1893,N_2359);
nand U2826 (N_2826,N_1940,N_1646);
nor U2827 (N_2827,N_1753,N_1802);
and U2828 (N_2828,N_1628,N_2348);
nand U2829 (N_2829,N_1745,N_2265);
or U2830 (N_2830,N_2121,N_2149);
and U2831 (N_2831,N_1694,N_1805);
xor U2832 (N_2832,N_2079,N_2107);
or U2833 (N_2833,N_1879,N_2198);
nor U2834 (N_2834,N_2356,N_2391);
nand U2835 (N_2835,N_1960,N_2342);
nand U2836 (N_2836,N_2051,N_1657);
nand U2837 (N_2837,N_2066,N_1640);
or U2838 (N_2838,N_2123,N_2246);
xnor U2839 (N_2839,N_1932,N_1724);
nor U2840 (N_2840,N_2183,N_1852);
or U2841 (N_2841,N_2311,N_1770);
or U2842 (N_2842,N_1784,N_2126);
xor U2843 (N_2843,N_2354,N_1764);
and U2844 (N_2844,N_2092,N_1955);
or U2845 (N_2845,N_2226,N_2363);
nand U2846 (N_2846,N_2111,N_2142);
xnor U2847 (N_2847,N_1666,N_2116);
or U2848 (N_2848,N_1630,N_1785);
or U2849 (N_2849,N_1874,N_2006);
nor U2850 (N_2850,N_1796,N_2352);
nor U2851 (N_2851,N_2031,N_1774);
or U2852 (N_2852,N_1924,N_1830);
or U2853 (N_2853,N_1899,N_2328);
xor U2854 (N_2854,N_1715,N_2074);
nor U2855 (N_2855,N_1826,N_1637);
or U2856 (N_2856,N_2130,N_2346);
and U2857 (N_2857,N_2252,N_1813);
and U2858 (N_2858,N_2184,N_1892);
nor U2859 (N_2859,N_2064,N_2023);
xor U2860 (N_2860,N_2154,N_1969);
and U2861 (N_2861,N_2241,N_2091);
and U2862 (N_2862,N_1716,N_1757);
nor U2863 (N_2863,N_2287,N_2349);
or U2864 (N_2864,N_2060,N_2059);
and U2865 (N_2865,N_2342,N_1670);
and U2866 (N_2866,N_1888,N_1795);
nor U2867 (N_2867,N_2069,N_1703);
xor U2868 (N_2868,N_1695,N_1971);
xor U2869 (N_2869,N_2396,N_1836);
xor U2870 (N_2870,N_1799,N_2146);
nor U2871 (N_2871,N_2017,N_1680);
or U2872 (N_2872,N_1743,N_1906);
nor U2873 (N_2873,N_1887,N_2135);
and U2874 (N_2874,N_2146,N_2204);
xnor U2875 (N_2875,N_2361,N_2032);
and U2876 (N_2876,N_2154,N_1739);
and U2877 (N_2877,N_1966,N_2098);
nand U2878 (N_2878,N_2303,N_2284);
or U2879 (N_2879,N_2384,N_1856);
nor U2880 (N_2880,N_1925,N_1797);
nor U2881 (N_2881,N_2241,N_1884);
nor U2882 (N_2882,N_1744,N_2069);
or U2883 (N_2883,N_2181,N_1945);
or U2884 (N_2884,N_1618,N_2156);
nand U2885 (N_2885,N_1652,N_2309);
nor U2886 (N_2886,N_2055,N_1932);
nor U2887 (N_2887,N_1731,N_1805);
nand U2888 (N_2888,N_1619,N_2156);
nor U2889 (N_2889,N_1650,N_2111);
nand U2890 (N_2890,N_1973,N_2272);
nand U2891 (N_2891,N_1610,N_2091);
and U2892 (N_2892,N_2380,N_1627);
nand U2893 (N_2893,N_2201,N_1793);
and U2894 (N_2894,N_1754,N_2262);
and U2895 (N_2895,N_1951,N_2306);
xnor U2896 (N_2896,N_1737,N_2191);
nor U2897 (N_2897,N_1893,N_2354);
xnor U2898 (N_2898,N_2041,N_1742);
nand U2899 (N_2899,N_2377,N_2017);
xor U2900 (N_2900,N_2334,N_1619);
nand U2901 (N_2901,N_2390,N_2330);
nor U2902 (N_2902,N_1686,N_2003);
and U2903 (N_2903,N_2334,N_1739);
nand U2904 (N_2904,N_1651,N_1605);
or U2905 (N_2905,N_2136,N_2113);
nor U2906 (N_2906,N_2368,N_2292);
and U2907 (N_2907,N_2345,N_2062);
or U2908 (N_2908,N_2198,N_1663);
xnor U2909 (N_2909,N_2385,N_2027);
nor U2910 (N_2910,N_1642,N_1828);
nor U2911 (N_2911,N_1646,N_2348);
nand U2912 (N_2912,N_1909,N_2193);
nand U2913 (N_2913,N_2073,N_2318);
nand U2914 (N_2914,N_1967,N_1844);
nand U2915 (N_2915,N_1805,N_2237);
or U2916 (N_2916,N_1979,N_1970);
or U2917 (N_2917,N_1807,N_1778);
or U2918 (N_2918,N_1615,N_1974);
nor U2919 (N_2919,N_1796,N_2181);
or U2920 (N_2920,N_1871,N_2278);
and U2921 (N_2921,N_2125,N_2278);
nand U2922 (N_2922,N_2318,N_1797);
and U2923 (N_2923,N_2220,N_2391);
nor U2924 (N_2924,N_2381,N_2302);
and U2925 (N_2925,N_1938,N_1955);
nand U2926 (N_2926,N_2364,N_2180);
nand U2927 (N_2927,N_2217,N_1638);
or U2928 (N_2928,N_1911,N_2237);
nor U2929 (N_2929,N_1672,N_2121);
xor U2930 (N_2930,N_2209,N_1787);
and U2931 (N_2931,N_1841,N_1999);
nor U2932 (N_2932,N_2115,N_2219);
and U2933 (N_2933,N_1681,N_1801);
or U2934 (N_2934,N_2080,N_1882);
nand U2935 (N_2935,N_1727,N_1955);
and U2936 (N_2936,N_2258,N_1680);
nor U2937 (N_2937,N_1955,N_1962);
and U2938 (N_2938,N_1673,N_2110);
nor U2939 (N_2939,N_1957,N_1671);
or U2940 (N_2940,N_2179,N_1781);
or U2941 (N_2941,N_2022,N_1891);
and U2942 (N_2942,N_2042,N_1926);
xor U2943 (N_2943,N_1602,N_1948);
or U2944 (N_2944,N_2042,N_2271);
xor U2945 (N_2945,N_1744,N_2093);
or U2946 (N_2946,N_1915,N_2384);
nand U2947 (N_2947,N_1758,N_2311);
nor U2948 (N_2948,N_2086,N_1615);
and U2949 (N_2949,N_1826,N_2040);
xnor U2950 (N_2950,N_2342,N_2250);
nand U2951 (N_2951,N_1950,N_1669);
xnor U2952 (N_2952,N_2306,N_1737);
xnor U2953 (N_2953,N_1853,N_1946);
or U2954 (N_2954,N_1992,N_1743);
nand U2955 (N_2955,N_1865,N_1682);
and U2956 (N_2956,N_1958,N_2186);
nor U2957 (N_2957,N_1952,N_1681);
or U2958 (N_2958,N_2018,N_2353);
nand U2959 (N_2959,N_2104,N_2356);
nor U2960 (N_2960,N_1602,N_1829);
nor U2961 (N_2961,N_2066,N_1762);
and U2962 (N_2962,N_1949,N_2125);
or U2963 (N_2963,N_2379,N_2283);
nand U2964 (N_2964,N_1686,N_1764);
or U2965 (N_2965,N_2223,N_1670);
nor U2966 (N_2966,N_2169,N_2134);
nor U2967 (N_2967,N_2042,N_1720);
xnor U2968 (N_2968,N_1737,N_2210);
nor U2969 (N_2969,N_2028,N_2307);
xnor U2970 (N_2970,N_2353,N_1716);
and U2971 (N_2971,N_2185,N_2369);
nand U2972 (N_2972,N_2358,N_1905);
xnor U2973 (N_2973,N_2187,N_1994);
xnor U2974 (N_2974,N_2282,N_2266);
nor U2975 (N_2975,N_2226,N_2320);
nor U2976 (N_2976,N_2093,N_1709);
and U2977 (N_2977,N_1780,N_1720);
nand U2978 (N_2978,N_1825,N_2083);
and U2979 (N_2979,N_1610,N_2117);
nor U2980 (N_2980,N_2150,N_1755);
xnor U2981 (N_2981,N_2027,N_2231);
nand U2982 (N_2982,N_1770,N_2352);
and U2983 (N_2983,N_1675,N_1664);
or U2984 (N_2984,N_2042,N_2268);
nand U2985 (N_2985,N_2102,N_1669);
nor U2986 (N_2986,N_1659,N_2268);
and U2987 (N_2987,N_2110,N_1796);
nor U2988 (N_2988,N_2068,N_1927);
xnor U2989 (N_2989,N_1800,N_1964);
nand U2990 (N_2990,N_1759,N_2046);
or U2991 (N_2991,N_2259,N_1791);
xor U2992 (N_2992,N_2023,N_1916);
xor U2993 (N_2993,N_1691,N_2079);
and U2994 (N_2994,N_2396,N_2073);
xor U2995 (N_2995,N_1618,N_2053);
and U2996 (N_2996,N_2242,N_2183);
nor U2997 (N_2997,N_2001,N_1753);
nand U2998 (N_2998,N_2236,N_1968);
nand U2999 (N_2999,N_1848,N_1837);
nand U3000 (N_3000,N_2391,N_1920);
xor U3001 (N_3001,N_1730,N_2034);
or U3002 (N_3002,N_1967,N_1769);
nand U3003 (N_3003,N_2087,N_1739);
or U3004 (N_3004,N_1976,N_2325);
or U3005 (N_3005,N_2112,N_2050);
and U3006 (N_3006,N_1675,N_1697);
nand U3007 (N_3007,N_1972,N_2214);
nor U3008 (N_3008,N_1800,N_2307);
nand U3009 (N_3009,N_2258,N_1819);
nand U3010 (N_3010,N_2024,N_2086);
nand U3011 (N_3011,N_2084,N_2020);
or U3012 (N_3012,N_2306,N_2180);
or U3013 (N_3013,N_1657,N_2192);
xor U3014 (N_3014,N_1845,N_2363);
nor U3015 (N_3015,N_2038,N_1927);
or U3016 (N_3016,N_1864,N_2107);
nand U3017 (N_3017,N_2378,N_1938);
nor U3018 (N_3018,N_1764,N_1724);
xor U3019 (N_3019,N_2380,N_2187);
xor U3020 (N_3020,N_1880,N_1900);
nor U3021 (N_3021,N_2089,N_1789);
or U3022 (N_3022,N_1999,N_2162);
xor U3023 (N_3023,N_1773,N_1842);
xnor U3024 (N_3024,N_2314,N_2055);
or U3025 (N_3025,N_2156,N_2221);
nor U3026 (N_3026,N_2358,N_1983);
nor U3027 (N_3027,N_1779,N_2338);
or U3028 (N_3028,N_2120,N_1832);
nor U3029 (N_3029,N_2048,N_2384);
and U3030 (N_3030,N_1622,N_2077);
and U3031 (N_3031,N_2266,N_1874);
and U3032 (N_3032,N_2176,N_1902);
or U3033 (N_3033,N_1956,N_2115);
xor U3034 (N_3034,N_1685,N_1799);
nand U3035 (N_3035,N_2178,N_2016);
and U3036 (N_3036,N_1797,N_2284);
xnor U3037 (N_3037,N_1763,N_2333);
nor U3038 (N_3038,N_1843,N_2097);
or U3039 (N_3039,N_2299,N_2174);
nand U3040 (N_3040,N_1859,N_2133);
nor U3041 (N_3041,N_2024,N_2251);
or U3042 (N_3042,N_1690,N_1829);
nor U3043 (N_3043,N_2093,N_2281);
xnor U3044 (N_3044,N_2305,N_1605);
or U3045 (N_3045,N_1742,N_1822);
nor U3046 (N_3046,N_2349,N_2108);
and U3047 (N_3047,N_1612,N_2327);
and U3048 (N_3048,N_2074,N_2352);
nand U3049 (N_3049,N_1726,N_2085);
nor U3050 (N_3050,N_2015,N_2137);
and U3051 (N_3051,N_2143,N_1823);
or U3052 (N_3052,N_2231,N_2391);
and U3053 (N_3053,N_1680,N_1781);
nor U3054 (N_3054,N_1790,N_1605);
nand U3055 (N_3055,N_2294,N_1873);
or U3056 (N_3056,N_2226,N_1677);
and U3057 (N_3057,N_1647,N_2196);
nand U3058 (N_3058,N_2308,N_1634);
xnor U3059 (N_3059,N_1989,N_2370);
nand U3060 (N_3060,N_2184,N_2387);
xor U3061 (N_3061,N_1670,N_2252);
nor U3062 (N_3062,N_1923,N_2275);
nand U3063 (N_3063,N_1691,N_1701);
and U3064 (N_3064,N_1889,N_1709);
or U3065 (N_3065,N_2038,N_1831);
or U3066 (N_3066,N_2279,N_2079);
and U3067 (N_3067,N_1749,N_2344);
and U3068 (N_3068,N_2268,N_1604);
xor U3069 (N_3069,N_1840,N_1878);
nand U3070 (N_3070,N_2275,N_2070);
or U3071 (N_3071,N_2312,N_1811);
or U3072 (N_3072,N_1710,N_1690);
xnor U3073 (N_3073,N_1620,N_1792);
nand U3074 (N_3074,N_1979,N_2019);
nand U3075 (N_3075,N_1704,N_1810);
nand U3076 (N_3076,N_1710,N_2154);
or U3077 (N_3077,N_2047,N_1696);
xnor U3078 (N_3078,N_1685,N_1838);
and U3079 (N_3079,N_1727,N_2195);
nor U3080 (N_3080,N_2350,N_2143);
xnor U3081 (N_3081,N_2279,N_1741);
and U3082 (N_3082,N_1834,N_2316);
nand U3083 (N_3083,N_2158,N_2384);
nand U3084 (N_3084,N_2062,N_2324);
xnor U3085 (N_3085,N_1808,N_1758);
or U3086 (N_3086,N_1975,N_1782);
nor U3087 (N_3087,N_2253,N_1633);
and U3088 (N_3088,N_1685,N_1751);
and U3089 (N_3089,N_2042,N_2053);
or U3090 (N_3090,N_2284,N_2344);
nand U3091 (N_3091,N_1827,N_1688);
and U3092 (N_3092,N_2227,N_1711);
or U3093 (N_3093,N_1863,N_2206);
or U3094 (N_3094,N_1824,N_1781);
nor U3095 (N_3095,N_2342,N_2141);
xor U3096 (N_3096,N_1694,N_2336);
and U3097 (N_3097,N_1972,N_2301);
nand U3098 (N_3098,N_1816,N_1766);
nor U3099 (N_3099,N_1916,N_1920);
nand U3100 (N_3100,N_1701,N_1783);
and U3101 (N_3101,N_1806,N_2029);
nor U3102 (N_3102,N_1627,N_1696);
nand U3103 (N_3103,N_1968,N_2352);
or U3104 (N_3104,N_1900,N_1752);
nor U3105 (N_3105,N_2021,N_1740);
or U3106 (N_3106,N_2297,N_2310);
xnor U3107 (N_3107,N_1717,N_2060);
or U3108 (N_3108,N_1626,N_2042);
and U3109 (N_3109,N_1609,N_1858);
or U3110 (N_3110,N_1890,N_1768);
nand U3111 (N_3111,N_1655,N_1995);
or U3112 (N_3112,N_1632,N_1898);
or U3113 (N_3113,N_1879,N_2162);
nor U3114 (N_3114,N_1890,N_2278);
and U3115 (N_3115,N_1627,N_1667);
nand U3116 (N_3116,N_1903,N_1954);
nor U3117 (N_3117,N_2048,N_1954);
nand U3118 (N_3118,N_2381,N_2241);
xor U3119 (N_3119,N_2369,N_2138);
and U3120 (N_3120,N_2204,N_1652);
xor U3121 (N_3121,N_1915,N_1743);
nor U3122 (N_3122,N_1617,N_1768);
nor U3123 (N_3123,N_2169,N_2078);
and U3124 (N_3124,N_2032,N_2078);
and U3125 (N_3125,N_1676,N_2286);
nor U3126 (N_3126,N_1726,N_2201);
or U3127 (N_3127,N_1885,N_1604);
xor U3128 (N_3128,N_2036,N_2285);
or U3129 (N_3129,N_1866,N_2292);
nand U3130 (N_3130,N_2067,N_2258);
nand U3131 (N_3131,N_1751,N_1695);
nor U3132 (N_3132,N_1726,N_2204);
xor U3133 (N_3133,N_1889,N_2011);
xnor U3134 (N_3134,N_1711,N_2204);
or U3135 (N_3135,N_1954,N_2167);
nor U3136 (N_3136,N_2343,N_1931);
nand U3137 (N_3137,N_1677,N_2097);
nor U3138 (N_3138,N_2305,N_1944);
and U3139 (N_3139,N_1825,N_1842);
xor U3140 (N_3140,N_1803,N_1951);
xnor U3141 (N_3141,N_2209,N_1997);
and U3142 (N_3142,N_2150,N_1932);
xor U3143 (N_3143,N_1977,N_2381);
or U3144 (N_3144,N_2228,N_2351);
nand U3145 (N_3145,N_1844,N_1724);
or U3146 (N_3146,N_2178,N_2166);
xnor U3147 (N_3147,N_1757,N_2163);
nand U3148 (N_3148,N_2191,N_1637);
xor U3149 (N_3149,N_2303,N_1738);
nand U3150 (N_3150,N_2052,N_1981);
xnor U3151 (N_3151,N_2178,N_1937);
or U3152 (N_3152,N_1816,N_1794);
nand U3153 (N_3153,N_2384,N_1755);
xor U3154 (N_3154,N_2302,N_1800);
and U3155 (N_3155,N_2291,N_1669);
nand U3156 (N_3156,N_1645,N_1634);
or U3157 (N_3157,N_2038,N_1752);
or U3158 (N_3158,N_2360,N_2076);
nor U3159 (N_3159,N_1831,N_1738);
and U3160 (N_3160,N_2279,N_2150);
nor U3161 (N_3161,N_2390,N_1652);
nor U3162 (N_3162,N_2092,N_2093);
xor U3163 (N_3163,N_1866,N_1887);
xor U3164 (N_3164,N_2301,N_2056);
and U3165 (N_3165,N_2358,N_1961);
xnor U3166 (N_3166,N_1763,N_1662);
nand U3167 (N_3167,N_1622,N_1855);
xor U3168 (N_3168,N_2373,N_1832);
nor U3169 (N_3169,N_1651,N_1754);
nand U3170 (N_3170,N_2312,N_1641);
or U3171 (N_3171,N_1939,N_1996);
nor U3172 (N_3172,N_2392,N_2124);
nor U3173 (N_3173,N_1717,N_2027);
and U3174 (N_3174,N_2074,N_2326);
nand U3175 (N_3175,N_1644,N_1949);
and U3176 (N_3176,N_2383,N_1660);
and U3177 (N_3177,N_1983,N_1865);
and U3178 (N_3178,N_2174,N_1911);
nor U3179 (N_3179,N_2107,N_1729);
and U3180 (N_3180,N_2318,N_2384);
xnor U3181 (N_3181,N_1662,N_2396);
or U3182 (N_3182,N_1944,N_1638);
and U3183 (N_3183,N_2260,N_2065);
nor U3184 (N_3184,N_1977,N_2380);
nor U3185 (N_3185,N_2369,N_1734);
nor U3186 (N_3186,N_2091,N_1650);
nand U3187 (N_3187,N_2294,N_1688);
xor U3188 (N_3188,N_1746,N_2140);
and U3189 (N_3189,N_2170,N_2075);
nand U3190 (N_3190,N_2013,N_1754);
nor U3191 (N_3191,N_2326,N_2139);
or U3192 (N_3192,N_1705,N_2055);
xor U3193 (N_3193,N_2231,N_2375);
xor U3194 (N_3194,N_1622,N_2241);
nand U3195 (N_3195,N_2278,N_2030);
xor U3196 (N_3196,N_1733,N_2048);
nor U3197 (N_3197,N_2010,N_1667);
or U3198 (N_3198,N_2184,N_1963);
or U3199 (N_3199,N_1720,N_2051);
xnor U3200 (N_3200,N_2519,N_3047);
nand U3201 (N_3201,N_2682,N_3190);
and U3202 (N_3202,N_2902,N_3168);
nor U3203 (N_3203,N_2948,N_2827);
nor U3204 (N_3204,N_2495,N_2570);
and U3205 (N_3205,N_2459,N_3073);
xor U3206 (N_3206,N_2724,N_3016);
xor U3207 (N_3207,N_2956,N_3003);
xor U3208 (N_3208,N_3082,N_2668);
xor U3209 (N_3209,N_2634,N_3198);
xor U3210 (N_3210,N_2759,N_2700);
nand U3211 (N_3211,N_2811,N_3043);
nand U3212 (N_3212,N_2661,N_2665);
and U3213 (N_3213,N_2981,N_3086);
nand U3214 (N_3214,N_2691,N_2573);
and U3215 (N_3215,N_2653,N_2507);
nor U3216 (N_3216,N_2584,N_2806);
nand U3217 (N_3217,N_2767,N_2518);
or U3218 (N_3218,N_2589,N_2600);
nand U3219 (N_3219,N_3171,N_2404);
and U3220 (N_3220,N_2962,N_2963);
or U3221 (N_3221,N_2987,N_2477);
nor U3222 (N_3222,N_3014,N_2802);
nand U3223 (N_3223,N_2999,N_2539);
xor U3224 (N_3224,N_2763,N_2428);
and U3225 (N_3225,N_2636,N_2852);
nor U3226 (N_3226,N_2672,N_3040);
and U3227 (N_3227,N_2936,N_2747);
xnor U3228 (N_3228,N_2451,N_2940);
nor U3229 (N_3229,N_2647,N_2909);
or U3230 (N_3230,N_2410,N_2533);
and U3231 (N_3231,N_2833,N_2580);
and U3232 (N_3232,N_2403,N_3091);
and U3233 (N_3233,N_2897,N_3013);
nand U3234 (N_3234,N_3195,N_2844);
nand U3235 (N_3235,N_2860,N_2591);
nor U3236 (N_3236,N_2719,N_2671);
or U3237 (N_3237,N_2438,N_2406);
and U3238 (N_3238,N_3020,N_2854);
and U3239 (N_3239,N_3167,N_3093);
or U3240 (N_3240,N_2498,N_2540);
xnor U3241 (N_3241,N_2468,N_2456);
nor U3242 (N_3242,N_2474,N_2701);
or U3243 (N_3243,N_2819,N_2486);
nand U3244 (N_3244,N_2548,N_2933);
and U3245 (N_3245,N_2556,N_2654);
xnor U3246 (N_3246,N_3126,N_2890);
nor U3247 (N_3247,N_2554,N_3054);
and U3248 (N_3248,N_3011,N_2828);
xor U3249 (N_3249,N_3042,N_2640);
nor U3250 (N_3250,N_2775,N_2632);
and U3251 (N_3251,N_2513,N_2972);
nor U3252 (N_3252,N_2530,N_2746);
nand U3253 (N_3253,N_2889,N_3085);
and U3254 (N_3254,N_2749,N_2786);
or U3255 (N_3255,N_2740,N_2947);
xor U3256 (N_3256,N_3092,N_2764);
nor U3257 (N_3257,N_2483,N_2470);
or U3258 (N_3258,N_2583,N_2969);
nand U3259 (N_3259,N_3046,N_3111);
nand U3260 (N_3260,N_2585,N_2955);
xnor U3261 (N_3261,N_3109,N_3138);
nor U3262 (N_3262,N_2912,N_2801);
xor U3263 (N_3263,N_3050,N_2644);
nor U3264 (N_3264,N_3017,N_2941);
nor U3265 (N_3265,N_2447,N_2566);
and U3266 (N_3266,N_3112,N_2505);
nand U3267 (N_3267,N_2893,N_2508);
or U3268 (N_3268,N_2810,N_2820);
xnor U3269 (N_3269,N_3100,N_2750);
and U3270 (N_3270,N_2953,N_2516);
nor U3271 (N_3271,N_2843,N_2465);
xnor U3272 (N_3272,N_2718,N_3142);
nor U3273 (N_3273,N_2710,N_2723);
or U3274 (N_3274,N_2450,N_2496);
and U3275 (N_3275,N_2778,N_3137);
nor U3276 (N_3276,N_2887,N_2920);
nand U3277 (N_3277,N_2702,N_2419);
nand U3278 (N_3278,N_2721,N_3166);
xnor U3279 (N_3279,N_2576,N_2777);
xnor U3280 (N_3280,N_2954,N_3065);
nand U3281 (N_3281,N_2907,N_3118);
nor U3282 (N_3282,N_2814,N_2931);
or U3283 (N_3283,N_3180,N_2871);
nor U3284 (N_3284,N_3072,N_2880);
nand U3285 (N_3285,N_3056,N_2448);
or U3286 (N_3286,N_2679,N_3110);
or U3287 (N_3287,N_2524,N_2625);
nand U3288 (N_3288,N_2944,N_2864);
and U3289 (N_3289,N_3023,N_3045);
xor U3290 (N_3290,N_2908,N_2503);
nand U3291 (N_3291,N_2689,N_2607);
xor U3292 (N_3292,N_2731,N_2841);
nand U3293 (N_3293,N_2872,N_2703);
nand U3294 (N_3294,N_3121,N_2532);
nor U3295 (N_3295,N_2641,N_2582);
and U3296 (N_3296,N_3117,N_2413);
nand U3297 (N_3297,N_2652,N_2840);
xor U3298 (N_3298,N_3032,N_3162);
and U3299 (N_3299,N_2990,N_2735);
nor U3300 (N_3300,N_3015,N_2825);
nor U3301 (N_3301,N_2690,N_2432);
or U3302 (N_3302,N_2514,N_2903);
xnor U3303 (N_3303,N_3084,N_2568);
nand U3304 (N_3304,N_2858,N_3033);
and U3305 (N_3305,N_2961,N_2587);
and U3306 (N_3306,N_2541,N_2742);
nor U3307 (N_3307,N_2934,N_3172);
nor U3308 (N_3308,N_2949,N_2537);
nand U3309 (N_3309,N_2555,N_2717);
and U3310 (N_3310,N_2832,N_2957);
xnor U3311 (N_3311,N_2939,N_2744);
nand U3312 (N_3312,N_3150,N_2741);
nand U3313 (N_3313,N_2673,N_3035);
nor U3314 (N_3314,N_2462,N_2722);
or U3315 (N_3315,N_2433,N_2497);
nand U3316 (N_3316,N_2697,N_3107);
xnor U3317 (N_3317,N_2562,N_2688);
xnor U3318 (N_3318,N_2464,N_2423);
and U3319 (N_3319,N_2831,N_2895);
nor U3320 (N_3320,N_2984,N_2736);
nor U3321 (N_3321,N_2500,N_2793);
and U3322 (N_3322,N_2604,N_2886);
xor U3323 (N_3323,N_3146,N_2838);
nand U3324 (N_3324,N_3196,N_2856);
xnor U3325 (N_3325,N_2899,N_2463);
or U3326 (N_3326,N_3153,N_2935);
and U3327 (N_3327,N_2563,N_2715);
nand U3328 (N_3328,N_2928,N_3140);
nand U3329 (N_3329,N_3152,N_2845);
or U3330 (N_3330,N_3141,N_2528);
nor U3331 (N_3331,N_2996,N_2637);
and U3332 (N_3332,N_2734,N_2753);
and U3333 (N_3333,N_2476,N_3163);
and U3334 (N_3334,N_3120,N_2628);
nand U3335 (N_3335,N_2693,N_2914);
xnor U3336 (N_3336,N_3165,N_2650);
nor U3337 (N_3337,N_2453,N_3024);
xnor U3338 (N_3338,N_2593,N_2492);
and U3339 (N_3339,N_2575,N_2745);
and U3340 (N_3340,N_2992,N_2977);
nor U3341 (N_3341,N_2611,N_2817);
nand U3342 (N_3342,N_2904,N_2598);
xor U3343 (N_3343,N_2623,N_2439);
xor U3344 (N_3344,N_3041,N_2517);
nor U3345 (N_3345,N_2577,N_2445);
nand U3346 (N_3346,N_2437,N_3189);
and U3347 (N_3347,N_2752,N_3128);
or U3348 (N_3348,N_2449,N_2816);
nor U3349 (N_3349,N_3044,N_2815);
or U3350 (N_3350,N_2616,N_3078);
and U3351 (N_3351,N_3096,N_2918);
and U3352 (N_3352,N_3192,N_3057);
xor U3353 (N_3353,N_2882,N_2952);
and U3354 (N_3354,N_3133,N_3076);
nor U3355 (N_3355,N_2785,N_2620);
nand U3356 (N_3356,N_3053,N_2705);
or U3357 (N_3357,N_2642,N_2966);
or U3358 (N_3358,N_2751,N_2475);
nand U3359 (N_3359,N_2510,N_2834);
or U3360 (N_3360,N_2666,N_3185);
nand U3361 (N_3361,N_3063,N_2771);
nand U3362 (N_3362,N_2599,N_2967);
nor U3363 (N_3363,N_2624,N_3030);
or U3364 (N_3364,N_2979,N_2824);
nand U3365 (N_3365,N_3181,N_2971);
and U3366 (N_3366,N_2866,N_2557);
nor U3367 (N_3367,N_2643,N_2635);
nand U3368 (N_3368,N_2714,N_2919);
xnor U3369 (N_3369,N_2923,N_3176);
xor U3370 (N_3370,N_3036,N_2472);
or U3371 (N_3371,N_2830,N_3131);
xnor U3372 (N_3372,N_2489,N_2894);
xor U3373 (N_3373,N_2756,N_2425);
xnor U3374 (N_3374,N_3143,N_2772);
nand U3375 (N_3375,N_2869,N_3187);
nor U3376 (N_3376,N_2565,N_2482);
or U3377 (N_3377,N_2631,N_2501);
or U3378 (N_3378,N_2601,N_2687);
and U3379 (N_3379,N_2426,N_2848);
xor U3380 (N_3380,N_2846,N_2900);
nand U3381 (N_3381,N_2727,N_2658);
xor U3382 (N_3382,N_2695,N_2704);
and U3383 (N_3383,N_2603,N_3049);
nand U3384 (N_3384,N_3182,N_2946);
nor U3385 (N_3385,N_3018,N_3094);
nor U3386 (N_3386,N_2619,N_2504);
xor U3387 (N_3387,N_2991,N_2708);
nor U3388 (N_3388,N_2906,N_2862);
and U3389 (N_3389,N_3028,N_3113);
nor U3390 (N_3390,N_3037,N_2709);
xnor U3391 (N_3391,N_3157,N_2733);
xor U3392 (N_3392,N_3067,N_2592);
or U3393 (N_3393,N_2974,N_2527);
xnor U3394 (N_3394,N_2538,N_2626);
and U3395 (N_3395,N_2552,N_2629);
nor U3396 (N_3396,N_2660,N_3122);
or U3397 (N_3397,N_3199,N_2926);
nor U3398 (N_3398,N_3183,N_3048);
and U3399 (N_3399,N_2612,N_2441);
nand U3400 (N_3400,N_2546,N_2400);
nand U3401 (N_3401,N_2891,N_3031);
and U3402 (N_3402,N_2916,N_2766);
nand U3403 (N_3403,N_3005,N_2484);
nor U3404 (N_3404,N_3038,N_2706);
xnor U3405 (N_3405,N_3174,N_3064);
nor U3406 (N_3406,N_2412,N_2561);
and U3407 (N_3407,N_2473,N_2525);
and U3408 (N_3408,N_2536,N_2588);
and U3409 (N_3409,N_2932,N_2522);
and U3410 (N_3410,N_2550,N_2610);
xnor U3411 (N_3411,N_3103,N_2596);
or U3412 (N_3412,N_3097,N_2809);
xor U3413 (N_3413,N_2898,N_3124);
and U3414 (N_3414,N_2606,N_2417);
nor U3415 (N_3415,N_2595,N_2685);
xnor U3416 (N_3416,N_2659,N_2780);
nand U3417 (N_3417,N_2789,N_2427);
xnor U3418 (N_3418,N_2422,N_2922);
xor U3419 (N_3419,N_3130,N_3022);
xnor U3420 (N_3420,N_2980,N_2863);
nand U3421 (N_3421,N_3156,N_2559);
nand U3422 (N_3422,N_3188,N_2434);
or U3423 (N_3423,N_2648,N_2874);
or U3424 (N_3424,N_2558,N_2812);
nand U3425 (N_3425,N_2466,N_3001);
nor U3426 (N_3426,N_2769,N_2509);
nand U3427 (N_3427,N_2680,N_2460);
nor U3428 (N_3428,N_2711,N_2480);
and U3429 (N_3429,N_3007,N_3134);
xor U3430 (N_3430,N_2564,N_2925);
nand U3431 (N_3431,N_2681,N_2485);
and U3432 (N_3432,N_2892,N_2402);
or U3433 (N_3433,N_2535,N_2760);
xnor U3434 (N_3434,N_2859,N_2645);
nand U3435 (N_3435,N_3101,N_2618);
or U3436 (N_3436,N_2430,N_3029);
nor U3437 (N_3437,N_3164,N_2964);
nor U3438 (N_3438,N_3069,N_3108);
nand U3439 (N_3439,N_3139,N_2674);
and U3440 (N_3440,N_2797,N_3088);
xnor U3441 (N_3441,N_2849,N_2927);
and U3442 (N_3442,N_2549,N_3173);
nor U3443 (N_3443,N_2788,N_3055);
nand U3444 (N_3444,N_2888,N_2488);
xnor U3445 (N_3445,N_2782,N_2826);
and U3446 (N_3446,N_2471,N_3000);
xor U3447 (N_3447,N_2458,N_2521);
nand U3448 (N_3448,N_3068,N_3061);
xnor U3449 (N_3449,N_2790,N_3177);
and U3450 (N_3450,N_2960,N_2657);
nand U3451 (N_3451,N_2543,N_2917);
or U3452 (N_3452,N_2452,N_2855);
xor U3453 (N_3453,N_2446,N_2861);
or U3454 (N_3454,N_2885,N_2942);
or U3455 (N_3455,N_2523,N_3062);
or U3456 (N_3456,N_2959,N_2867);
or U3457 (N_3457,N_2569,N_2545);
nor U3458 (N_3458,N_2761,N_2613);
nor U3459 (N_3459,N_3051,N_2930);
xor U3460 (N_3460,N_2853,N_3116);
or U3461 (N_3461,N_3004,N_2408);
or U3462 (N_3462,N_2622,N_2779);
or U3463 (N_3463,N_2455,N_2664);
and U3464 (N_3464,N_2683,N_2416);
and U3465 (N_3465,N_2993,N_2594);
xnor U3466 (N_3466,N_2829,N_2667);
or U3467 (N_3467,N_2881,N_3147);
or U3468 (N_3468,N_2684,N_2421);
and U3469 (N_3469,N_2803,N_2454);
xnor U3470 (N_3470,N_2958,N_2968);
nor U3471 (N_3471,N_2970,N_2534);
nand U3472 (N_3472,N_3021,N_2581);
and U3473 (N_3473,N_3184,N_2478);
and U3474 (N_3474,N_2481,N_2997);
and U3475 (N_3475,N_3158,N_2847);
nor U3476 (N_3476,N_2656,N_2544);
and U3477 (N_3477,N_2879,N_2418);
xor U3478 (N_3478,N_3161,N_2865);
and U3479 (N_3479,N_2823,N_2995);
nand U3480 (N_3480,N_2526,N_3081);
and U3481 (N_3481,N_2586,N_2929);
nand U3482 (N_3482,N_2835,N_3194);
and U3483 (N_3483,N_3179,N_2499);
and U3484 (N_3484,N_2663,N_3149);
nand U3485 (N_3485,N_2884,N_3089);
and U3486 (N_3486,N_2726,N_3154);
nand U3487 (N_3487,N_2739,N_2553);
or U3488 (N_3488,N_2873,N_2945);
nor U3489 (N_3489,N_2877,N_2692);
or U3490 (N_3490,N_3095,N_3009);
or U3491 (N_3491,N_2986,N_2795);
nand U3492 (N_3492,N_3160,N_2783);
and U3493 (N_3493,N_2913,N_2560);
xnor U3494 (N_3494,N_2713,N_2567);
and U3495 (N_3495,N_2698,N_2662);
nor U3496 (N_3496,N_2608,N_2531);
xnor U3497 (N_3497,N_2633,N_2639);
or U3498 (N_3498,N_2494,N_2515);
nor U3499 (N_3499,N_3074,N_3039);
and U3500 (N_3500,N_2579,N_2405);
or U3501 (N_3501,N_2975,N_2988);
and U3502 (N_3502,N_2511,N_2768);
nor U3503 (N_3503,N_2551,N_2983);
nand U3504 (N_3504,N_2937,N_2738);
nand U3505 (N_3505,N_2730,N_2765);
and U3506 (N_3506,N_3144,N_2699);
nor U3507 (N_3507,N_2444,N_3136);
nor U3508 (N_3508,N_3075,N_2651);
or U3509 (N_3509,N_3080,N_2737);
or U3510 (N_3510,N_2813,N_2807);
xor U3511 (N_3511,N_3155,N_2951);
nand U3512 (N_3512,N_2414,N_2924);
or U3513 (N_3513,N_2716,N_3002);
and U3514 (N_3514,N_2787,N_3151);
nand U3515 (N_3515,N_2982,N_2978);
and U3516 (N_3516,N_2490,N_2915);
nor U3517 (N_3517,N_3148,N_2520);
xor U3518 (N_3518,N_3106,N_3125);
or U3519 (N_3519,N_3027,N_2965);
nor U3520 (N_3520,N_3175,N_2415);
nor U3521 (N_3521,N_2804,N_3191);
xnor U3522 (N_3522,N_2896,N_2818);
xnor U3523 (N_3523,N_3105,N_2431);
nand U3524 (N_3524,N_2440,N_3129);
nand U3525 (N_3525,N_2821,N_2762);
or U3526 (N_3526,N_2638,N_2720);
nand U3527 (N_3527,N_2694,N_2547);
or U3528 (N_3528,N_3058,N_2943);
xor U3529 (N_3529,N_2770,N_3178);
nand U3530 (N_3530,N_2487,N_2910);
nand U3531 (N_3531,N_2732,N_2675);
nor U3532 (N_3532,N_3079,N_2800);
nand U3533 (N_3533,N_2836,N_2757);
and U3534 (N_3534,N_2670,N_3193);
xnor U3535 (N_3535,N_2677,N_2850);
xnor U3536 (N_3536,N_2868,N_2424);
nor U3537 (N_3537,N_2590,N_2506);
nand U3538 (N_3538,N_2435,N_2707);
nor U3539 (N_3539,N_2605,N_2678);
nand U3540 (N_3540,N_2911,N_2905);
nor U3541 (N_3541,N_2725,N_2743);
or U3542 (N_3542,N_3066,N_2429);
and U3543 (N_3543,N_2878,N_2748);
nand U3544 (N_3544,N_2676,N_2839);
nand U3545 (N_3545,N_2512,N_2883);
xor U3546 (N_3546,N_2574,N_2976);
nand U3547 (N_3547,N_3119,N_3135);
or U3548 (N_3548,N_3132,N_2851);
xor U3549 (N_3549,N_2467,N_3169);
and U3550 (N_3550,N_3104,N_2578);
nand U3551 (N_3551,N_2758,N_3186);
and U3552 (N_3552,N_2621,N_2411);
or U3553 (N_3553,N_2938,N_2502);
and U3554 (N_3554,N_2822,N_3197);
and U3555 (N_3555,N_2798,N_3010);
xnor U3556 (N_3556,N_2443,N_2998);
or U3557 (N_3557,N_2627,N_3087);
or U3558 (N_3558,N_3025,N_3012);
xor U3559 (N_3559,N_2712,N_2875);
nand U3560 (N_3560,N_3060,N_2773);
xor U3561 (N_3561,N_2776,N_2542);
xor U3562 (N_3562,N_3114,N_3083);
nand U3563 (N_3563,N_2989,N_2597);
or U3564 (N_3564,N_2401,N_2729);
and U3565 (N_3565,N_3077,N_2842);
nand U3566 (N_3566,N_2409,N_3070);
or U3567 (N_3567,N_3102,N_2799);
and U3568 (N_3568,N_2529,N_2457);
and U3569 (N_3569,N_2870,N_2420);
and U3570 (N_3570,N_2784,N_2973);
and U3571 (N_3571,N_2493,N_2754);
nor U3572 (N_3572,N_2617,N_3071);
or U3573 (N_3573,N_2614,N_2876);
and U3574 (N_3574,N_2728,N_2436);
nor U3575 (N_3575,N_2857,N_2461);
nand U3576 (N_3576,N_2655,N_3123);
and U3577 (N_3577,N_2615,N_2602);
and U3578 (N_3578,N_2994,N_2808);
or U3579 (N_3579,N_2686,N_2921);
or U3580 (N_3580,N_3008,N_2805);
xnor U3581 (N_3581,N_2901,N_2669);
or U3582 (N_3582,N_2407,N_2794);
or U3583 (N_3583,N_2950,N_2609);
or U3584 (N_3584,N_2630,N_2837);
or U3585 (N_3585,N_3019,N_3127);
and U3586 (N_3586,N_3026,N_2442);
or U3587 (N_3587,N_2649,N_2792);
nor U3588 (N_3588,N_3145,N_3034);
nand U3589 (N_3589,N_2572,N_2791);
and U3590 (N_3590,N_3090,N_2985);
nor U3591 (N_3591,N_3006,N_2774);
and U3592 (N_3592,N_2696,N_3115);
nand U3593 (N_3593,N_2479,N_2796);
nor U3594 (N_3594,N_3059,N_3098);
xnor U3595 (N_3595,N_2571,N_3170);
and U3596 (N_3596,N_3052,N_2755);
or U3597 (N_3597,N_3099,N_3159);
and U3598 (N_3598,N_2646,N_2781);
and U3599 (N_3599,N_2491,N_2469);
or U3600 (N_3600,N_2810,N_2920);
nor U3601 (N_3601,N_2647,N_3020);
nor U3602 (N_3602,N_2693,N_2846);
xnor U3603 (N_3603,N_2523,N_2424);
nand U3604 (N_3604,N_2906,N_2861);
nor U3605 (N_3605,N_3006,N_2978);
xor U3606 (N_3606,N_2778,N_2966);
nor U3607 (N_3607,N_2901,N_2953);
nor U3608 (N_3608,N_3049,N_3151);
nand U3609 (N_3609,N_2408,N_3089);
nor U3610 (N_3610,N_3123,N_3122);
and U3611 (N_3611,N_2639,N_3158);
xor U3612 (N_3612,N_3077,N_3094);
or U3613 (N_3613,N_3031,N_2669);
and U3614 (N_3614,N_3196,N_3187);
nor U3615 (N_3615,N_2931,N_2961);
nor U3616 (N_3616,N_2998,N_3128);
or U3617 (N_3617,N_2765,N_2606);
or U3618 (N_3618,N_2447,N_2730);
xnor U3619 (N_3619,N_2727,N_2444);
nand U3620 (N_3620,N_3073,N_2553);
and U3621 (N_3621,N_3116,N_2886);
or U3622 (N_3622,N_2426,N_2833);
and U3623 (N_3623,N_2596,N_3168);
or U3624 (N_3624,N_2902,N_3179);
xnor U3625 (N_3625,N_2608,N_2677);
nand U3626 (N_3626,N_2465,N_3092);
xnor U3627 (N_3627,N_2476,N_3145);
or U3628 (N_3628,N_2744,N_2415);
and U3629 (N_3629,N_2909,N_2906);
or U3630 (N_3630,N_2887,N_2979);
nor U3631 (N_3631,N_3037,N_2664);
nand U3632 (N_3632,N_2409,N_2555);
xor U3633 (N_3633,N_3173,N_3194);
nand U3634 (N_3634,N_2442,N_2703);
xnor U3635 (N_3635,N_2734,N_3160);
xor U3636 (N_3636,N_2895,N_2787);
nand U3637 (N_3637,N_3036,N_2469);
nor U3638 (N_3638,N_2528,N_2455);
or U3639 (N_3639,N_2904,N_2778);
nor U3640 (N_3640,N_2956,N_2642);
or U3641 (N_3641,N_2813,N_2956);
nand U3642 (N_3642,N_2748,N_2458);
nand U3643 (N_3643,N_2765,N_2976);
xor U3644 (N_3644,N_2710,N_2562);
or U3645 (N_3645,N_2821,N_2940);
nand U3646 (N_3646,N_2547,N_2544);
xnor U3647 (N_3647,N_3131,N_2608);
nor U3648 (N_3648,N_2622,N_2903);
nand U3649 (N_3649,N_2620,N_2443);
nor U3650 (N_3650,N_2767,N_2867);
and U3651 (N_3651,N_2614,N_2415);
nand U3652 (N_3652,N_3172,N_2944);
or U3653 (N_3653,N_2510,N_3111);
or U3654 (N_3654,N_2992,N_2659);
nor U3655 (N_3655,N_2759,N_2492);
nand U3656 (N_3656,N_3134,N_2724);
xnor U3657 (N_3657,N_2830,N_3136);
xnor U3658 (N_3658,N_2476,N_2776);
nand U3659 (N_3659,N_2452,N_2420);
xnor U3660 (N_3660,N_2531,N_3010);
nand U3661 (N_3661,N_3130,N_2466);
xor U3662 (N_3662,N_2442,N_3030);
nand U3663 (N_3663,N_2453,N_3038);
and U3664 (N_3664,N_3197,N_2435);
nor U3665 (N_3665,N_2948,N_3092);
xor U3666 (N_3666,N_2729,N_2810);
nor U3667 (N_3667,N_3198,N_2519);
xor U3668 (N_3668,N_2692,N_2859);
xnor U3669 (N_3669,N_3086,N_2541);
nand U3670 (N_3670,N_2662,N_2643);
nor U3671 (N_3671,N_2826,N_3157);
or U3672 (N_3672,N_3072,N_2716);
and U3673 (N_3673,N_2980,N_2658);
xor U3674 (N_3674,N_2563,N_2748);
nor U3675 (N_3675,N_2626,N_3024);
or U3676 (N_3676,N_3122,N_2413);
nand U3677 (N_3677,N_3185,N_2813);
or U3678 (N_3678,N_2917,N_3044);
xor U3679 (N_3679,N_3159,N_2638);
and U3680 (N_3680,N_3031,N_2702);
and U3681 (N_3681,N_2836,N_2584);
and U3682 (N_3682,N_3085,N_2507);
and U3683 (N_3683,N_2759,N_2712);
xor U3684 (N_3684,N_2877,N_2576);
nor U3685 (N_3685,N_2618,N_2885);
nand U3686 (N_3686,N_2767,N_2967);
nand U3687 (N_3687,N_2409,N_3093);
nor U3688 (N_3688,N_2412,N_2949);
or U3689 (N_3689,N_3096,N_2937);
and U3690 (N_3690,N_3158,N_2852);
nor U3691 (N_3691,N_3033,N_2777);
nand U3692 (N_3692,N_2899,N_3004);
and U3693 (N_3693,N_3047,N_3143);
nor U3694 (N_3694,N_3114,N_2870);
nor U3695 (N_3695,N_2626,N_2753);
or U3696 (N_3696,N_2448,N_2915);
xnor U3697 (N_3697,N_2435,N_3025);
nor U3698 (N_3698,N_3179,N_2584);
nor U3699 (N_3699,N_2554,N_2540);
nand U3700 (N_3700,N_2717,N_2537);
nor U3701 (N_3701,N_3123,N_2879);
nor U3702 (N_3702,N_2889,N_2679);
xnor U3703 (N_3703,N_3070,N_2632);
or U3704 (N_3704,N_2492,N_3093);
nor U3705 (N_3705,N_3116,N_2951);
nand U3706 (N_3706,N_2451,N_2419);
xor U3707 (N_3707,N_2741,N_2811);
and U3708 (N_3708,N_2979,N_2563);
or U3709 (N_3709,N_2681,N_2625);
xnor U3710 (N_3710,N_2886,N_3085);
nand U3711 (N_3711,N_2509,N_2598);
nor U3712 (N_3712,N_3192,N_2984);
nor U3713 (N_3713,N_2457,N_2410);
nor U3714 (N_3714,N_2809,N_2543);
or U3715 (N_3715,N_3077,N_3152);
nor U3716 (N_3716,N_2820,N_2747);
nand U3717 (N_3717,N_2473,N_2915);
or U3718 (N_3718,N_3180,N_2699);
xor U3719 (N_3719,N_3104,N_2614);
nand U3720 (N_3720,N_2563,N_2549);
nand U3721 (N_3721,N_2776,N_2638);
or U3722 (N_3722,N_2435,N_2956);
nand U3723 (N_3723,N_3037,N_2693);
xnor U3724 (N_3724,N_2876,N_2773);
nor U3725 (N_3725,N_2941,N_2622);
and U3726 (N_3726,N_3122,N_2777);
and U3727 (N_3727,N_3090,N_2885);
or U3728 (N_3728,N_3152,N_2842);
or U3729 (N_3729,N_2847,N_2699);
xor U3730 (N_3730,N_2500,N_3061);
xor U3731 (N_3731,N_2437,N_2742);
xnor U3732 (N_3732,N_2484,N_2893);
nand U3733 (N_3733,N_2466,N_2852);
nand U3734 (N_3734,N_2929,N_2474);
nand U3735 (N_3735,N_2725,N_3033);
and U3736 (N_3736,N_2471,N_3191);
nand U3737 (N_3737,N_2426,N_3071);
or U3738 (N_3738,N_2952,N_2859);
and U3739 (N_3739,N_2550,N_2844);
xor U3740 (N_3740,N_2454,N_2901);
nor U3741 (N_3741,N_2745,N_3047);
nand U3742 (N_3742,N_2705,N_2664);
nor U3743 (N_3743,N_2400,N_2873);
nand U3744 (N_3744,N_2673,N_2796);
nand U3745 (N_3745,N_2539,N_2569);
nor U3746 (N_3746,N_2685,N_2429);
nor U3747 (N_3747,N_2494,N_2896);
nand U3748 (N_3748,N_2511,N_2610);
and U3749 (N_3749,N_2457,N_2433);
xnor U3750 (N_3750,N_2793,N_2978);
nand U3751 (N_3751,N_2992,N_2796);
nor U3752 (N_3752,N_3198,N_2590);
or U3753 (N_3753,N_2980,N_3099);
nor U3754 (N_3754,N_2599,N_2868);
or U3755 (N_3755,N_2976,N_3144);
nand U3756 (N_3756,N_2918,N_3150);
nor U3757 (N_3757,N_3181,N_3164);
or U3758 (N_3758,N_2607,N_2544);
xnor U3759 (N_3759,N_3078,N_2401);
xor U3760 (N_3760,N_2717,N_2781);
and U3761 (N_3761,N_2413,N_2552);
nand U3762 (N_3762,N_2435,N_2745);
or U3763 (N_3763,N_2745,N_3005);
nand U3764 (N_3764,N_2580,N_2430);
nor U3765 (N_3765,N_3029,N_2981);
or U3766 (N_3766,N_2999,N_2662);
nor U3767 (N_3767,N_3068,N_3188);
xor U3768 (N_3768,N_2770,N_2510);
or U3769 (N_3769,N_3167,N_2985);
nor U3770 (N_3770,N_2714,N_2893);
nor U3771 (N_3771,N_2438,N_3162);
or U3772 (N_3772,N_2895,N_2800);
nor U3773 (N_3773,N_2923,N_2562);
and U3774 (N_3774,N_2875,N_2775);
nand U3775 (N_3775,N_2763,N_2501);
nand U3776 (N_3776,N_2554,N_2736);
xor U3777 (N_3777,N_2449,N_2586);
nor U3778 (N_3778,N_2665,N_2954);
and U3779 (N_3779,N_2719,N_2464);
xnor U3780 (N_3780,N_2981,N_3159);
nand U3781 (N_3781,N_3095,N_3007);
nor U3782 (N_3782,N_2629,N_3188);
and U3783 (N_3783,N_2529,N_2833);
nor U3784 (N_3784,N_2553,N_3052);
or U3785 (N_3785,N_3111,N_2621);
and U3786 (N_3786,N_2537,N_2567);
or U3787 (N_3787,N_3047,N_2548);
nand U3788 (N_3788,N_2996,N_2826);
and U3789 (N_3789,N_3178,N_2849);
nor U3790 (N_3790,N_2705,N_2532);
nor U3791 (N_3791,N_3142,N_2641);
nor U3792 (N_3792,N_2421,N_2895);
and U3793 (N_3793,N_2614,N_2482);
xnor U3794 (N_3794,N_2452,N_2902);
nand U3795 (N_3795,N_2688,N_2623);
nor U3796 (N_3796,N_2479,N_2655);
and U3797 (N_3797,N_2424,N_2491);
nand U3798 (N_3798,N_3034,N_2799);
and U3799 (N_3799,N_2658,N_2993);
xnor U3800 (N_3800,N_3029,N_2916);
nor U3801 (N_3801,N_2470,N_2463);
and U3802 (N_3802,N_2899,N_2487);
nor U3803 (N_3803,N_3160,N_2526);
xor U3804 (N_3804,N_2420,N_3087);
and U3805 (N_3805,N_2885,N_2483);
and U3806 (N_3806,N_2408,N_2510);
nor U3807 (N_3807,N_3183,N_3058);
xor U3808 (N_3808,N_3155,N_2465);
nand U3809 (N_3809,N_3131,N_2980);
xnor U3810 (N_3810,N_2775,N_3154);
or U3811 (N_3811,N_2637,N_2837);
and U3812 (N_3812,N_2409,N_2513);
nor U3813 (N_3813,N_2669,N_2516);
nand U3814 (N_3814,N_2768,N_2890);
xnor U3815 (N_3815,N_3129,N_2912);
nand U3816 (N_3816,N_2570,N_2403);
nand U3817 (N_3817,N_2825,N_2470);
xnor U3818 (N_3818,N_2682,N_2998);
xnor U3819 (N_3819,N_3091,N_2793);
and U3820 (N_3820,N_2896,N_2663);
xnor U3821 (N_3821,N_2516,N_2584);
or U3822 (N_3822,N_2962,N_2561);
and U3823 (N_3823,N_3077,N_2589);
xor U3824 (N_3824,N_2851,N_2848);
and U3825 (N_3825,N_2419,N_3065);
nor U3826 (N_3826,N_2684,N_3110);
nand U3827 (N_3827,N_2926,N_2900);
nand U3828 (N_3828,N_3190,N_3174);
nor U3829 (N_3829,N_2414,N_2858);
nand U3830 (N_3830,N_2689,N_2662);
nor U3831 (N_3831,N_2569,N_2737);
nand U3832 (N_3832,N_3084,N_3178);
nand U3833 (N_3833,N_2733,N_2687);
nor U3834 (N_3834,N_3057,N_2561);
nand U3835 (N_3835,N_2978,N_2720);
xnor U3836 (N_3836,N_2687,N_3114);
nor U3837 (N_3837,N_2429,N_3114);
nor U3838 (N_3838,N_2652,N_2955);
and U3839 (N_3839,N_3162,N_2483);
xor U3840 (N_3840,N_3116,N_2450);
nand U3841 (N_3841,N_3196,N_2999);
nand U3842 (N_3842,N_2421,N_2869);
xnor U3843 (N_3843,N_2880,N_3152);
and U3844 (N_3844,N_2522,N_2623);
nand U3845 (N_3845,N_2681,N_2632);
nor U3846 (N_3846,N_2526,N_3020);
nand U3847 (N_3847,N_3102,N_2951);
xor U3848 (N_3848,N_2470,N_2623);
nand U3849 (N_3849,N_2665,N_2783);
xnor U3850 (N_3850,N_2503,N_2888);
xnor U3851 (N_3851,N_2561,N_2696);
and U3852 (N_3852,N_2917,N_3107);
or U3853 (N_3853,N_2745,N_2523);
nor U3854 (N_3854,N_2952,N_2731);
or U3855 (N_3855,N_2405,N_2848);
and U3856 (N_3856,N_2666,N_3182);
and U3857 (N_3857,N_2526,N_2552);
nor U3858 (N_3858,N_3006,N_2431);
nand U3859 (N_3859,N_2609,N_2660);
nor U3860 (N_3860,N_2872,N_3099);
nand U3861 (N_3861,N_2502,N_3090);
and U3862 (N_3862,N_3136,N_2892);
nand U3863 (N_3863,N_2745,N_2805);
nor U3864 (N_3864,N_3005,N_2900);
or U3865 (N_3865,N_2715,N_2555);
or U3866 (N_3866,N_2586,N_2985);
or U3867 (N_3867,N_2471,N_2644);
or U3868 (N_3868,N_2661,N_2987);
xnor U3869 (N_3869,N_3000,N_2753);
xnor U3870 (N_3870,N_3092,N_2861);
nor U3871 (N_3871,N_2783,N_2423);
or U3872 (N_3872,N_3027,N_3150);
and U3873 (N_3873,N_2813,N_3008);
nand U3874 (N_3874,N_2424,N_2631);
and U3875 (N_3875,N_2795,N_3164);
and U3876 (N_3876,N_2837,N_2910);
nor U3877 (N_3877,N_2527,N_2720);
and U3878 (N_3878,N_2646,N_2926);
or U3879 (N_3879,N_2866,N_2560);
nor U3880 (N_3880,N_3024,N_2513);
nor U3881 (N_3881,N_2886,N_2603);
nand U3882 (N_3882,N_3127,N_2885);
xnor U3883 (N_3883,N_2847,N_2617);
or U3884 (N_3884,N_2755,N_2806);
nor U3885 (N_3885,N_3196,N_3169);
xnor U3886 (N_3886,N_3131,N_3183);
nand U3887 (N_3887,N_3147,N_2416);
or U3888 (N_3888,N_2888,N_2801);
nor U3889 (N_3889,N_2645,N_2976);
xor U3890 (N_3890,N_3188,N_2524);
nand U3891 (N_3891,N_3041,N_3125);
or U3892 (N_3892,N_2476,N_2679);
and U3893 (N_3893,N_2815,N_2862);
or U3894 (N_3894,N_2928,N_3049);
and U3895 (N_3895,N_2806,N_3070);
or U3896 (N_3896,N_2464,N_3087);
nor U3897 (N_3897,N_2456,N_2494);
nor U3898 (N_3898,N_2589,N_2836);
and U3899 (N_3899,N_3100,N_2787);
xnor U3900 (N_3900,N_2906,N_2986);
nor U3901 (N_3901,N_2488,N_2441);
xor U3902 (N_3902,N_2643,N_3020);
and U3903 (N_3903,N_2796,N_3109);
and U3904 (N_3904,N_2549,N_2600);
or U3905 (N_3905,N_2420,N_2960);
nor U3906 (N_3906,N_3007,N_2866);
nor U3907 (N_3907,N_3083,N_2920);
nor U3908 (N_3908,N_2883,N_2550);
and U3909 (N_3909,N_2568,N_2561);
xor U3910 (N_3910,N_2622,N_2416);
and U3911 (N_3911,N_2934,N_2937);
and U3912 (N_3912,N_2932,N_2610);
nand U3913 (N_3913,N_3099,N_2735);
or U3914 (N_3914,N_2711,N_2967);
nand U3915 (N_3915,N_3146,N_2602);
and U3916 (N_3916,N_2962,N_3164);
nand U3917 (N_3917,N_2500,N_2428);
and U3918 (N_3918,N_2774,N_2939);
xor U3919 (N_3919,N_3142,N_2939);
xnor U3920 (N_3920,N_2693,N_2526);
and U3921 (N_3921,N_2406,N_2815);
and U3922 (N_3922,N_2867,N_3012);
and U3923 (N_3923,N_3169,N_2469);
xor U3924 (N_3924,N_2560,N_2610);
nand U3925 (N_3925,N_2851,N_2488);
nor U3926 (N_3926,N_2865,N_2873);
xnor U3927 (N_3927,N_2759,N_2709);
or U3928 (N_3928,N_2706,N_2782);
nand U3929 (N_3929,N_2690,N_2960);
xnor U3930 (N_3930,N_2423,N_2996);
nor U3931 (N_3931,N_3073,N_2887);
nand U3932 (N_3932,N_2972,N_2964);
nand U3933 (N_3933,N_3089,N_3014);
or U3934 (N_3934,N_2533,N_2632);
or U3935 (N_3935,N_2725,N_2767);
xor U3936 (N_3936,N_2792,N_2558);
xor U3937 (N_3937,N_2478,N_3127);
or U3938 (N_3938,N_2541,N_2770);
or U3939 (N_3939,N_2933,N_2461);
and U3940 (N_3940,N_3027,N_2420);
xor U3941 (N_3941,N_2886,N_2580);
xnor U3942 (N_3942,N_3134,N_2493);
nand U3943 (N_3943,N_3007,N_3180);
or U3944 (N_3944,N_3144,N_2825);
nor U3945 (N_3945,N_3109,N_3085);
and U3946 (N_3946,N_3155,N_3082);
nand U3947 (N_3947,N_2821,N_3000);
and U3948 (N_3948,N_2785,N_2426);
or U3949 (N_3949,N_2579,N_2546);
and U3950 (N_3950,N_2712,N_2858);
nand U3951 (N_3951,N_2735,N_3030);
and U3952 (N_3952,N_3105,N_2428);
and U3953 (N_3953,N_2956,N_3069);
nand U3954 (N_3954,N_2882,N_3003);
xnor U3955 (N_3955,N_2830,N_2899);
xor U3956 (N_3956,N_3147,N_2625);
and U3957 (N_3957,N_2876,N_3024);
and U3958 (N_3958,N_2561,N_2863);
nor U3959 (N_3959,N_3057,N_2746);
xnor U3960 (N_3960,N_2800,N_3144);
or U3961 (N_3961,N_2757,N_2860);
or U3962 (N_3962,N_2510,N_3155);
or U3963 (N_3963,N_2837,N_2931);
nand U3964 (N_3964,N_2654,N_3126);
xor U3965 (N_3965,N_2722,N_2858);
nand U3966 (N_3966,N_3087,N_2620);
nor U3967 (N_3967,N_2559,N_2640);
xnor U3968 (N_3968,N_2416,N_2950);
nor U3969 (N_3969,N_2989,N_3091);
and U3970 (N_3970,N_2485,N_2934);
nor U3971 (N_3971,N_2411,N_2925);
and U3972 (N_3972,N_2766,N_2502);
nand U3973 (N_3973,N_2876,N_3090);
xnor U3974 (N_3974,N_2788,N_2783);
nor U3975 (N_3975,N_2920,N_2574);
and U3976 (N_3976,N_2556,N_2510);
nor U3977 (N_3977,N_3050,N_2654);
and U3978 (N_3978,N_2964,N_2657);
nand U3979 (N_3979,N_2941,N_2795);
or U3980 (N_3980,N_2997,N_3035);
or U3981 (N_3981,N_2484,N_3169);
nand U3982 (N_3982,N_2466,N_3160);
xor U3983 (N_3983,N_2662,N_3158);
nand U3984 (N_3984,N_2560,N_2897);
or U3985 (N_3985,N_2419,N_2405);
nand U3986 (N_3986,N_2694,N_2909);
nor U3987 (N_3987,N_2606,N_2815);
xor U3988 (N_3988,N_2464,N_3080);
and U3989 (N_3989,N_3051,N_2843);
xor U3990 (N_3990,N_2424,N_2499);
xor U3991 (N_3991,N_3088,N_3194);
xnor U3992 (N_3992,N_3172,N_2512);
nor U3993 (N_3993,N_2598,N_3061);
and U3994 (N_3994,N_2717,N_2948);
and U3995 (N_3995,N_2820,N_2693);
nor U3996 (N_3996,N_2742,N_3114);
and U3997 (N_3997,N_3081,N_2841);
and U3998 (N_3998,N_2476,N_3006);
nand U3999 (N_3999,N_2528,N_2563);
xnor U4000 (N_4000,N_3495,N_3617);
or U4001 (N_4001,N_3968,N_3484);
xnor U4002 (N_4002,N_3881,N_3685);
nand U4003 (N_4003,N_3777,N_3566);
nand U4004 (N_4004,N_3594,N_3438);
or U4005 (N_4005,N_3596,N_3900);
xor U4006 (N_4006,N_3887,N_3750);
and U4007 (N_4007,N_3783,N_3318);
or U4008 (N_4008,N_3207,N_3742);
nand U4009 (N_4009,N_3591,N_3980);
nand U4010 (N_4010,N_3612,N_3333);
nor U4011 (N_4011,N_3278,N_3850);
nand U4012 (N_4012,N_3841,N_3236);
nor U4013 (N_4013,N_3509,N_3354);
and U4014 (N_4014,N_3677,N_3827);
and U4015 (N_4015,N_3398,N_3544);
xnor U4016 (N_4016,N_3905,N_3849);
and U4017 (N_4017,N_3523,N_3731);
xnor U4018 (N_4018,N_3532,N_3434);
or U4019 (N_4019,N_3796,N_3671);
or U4020 (N_4020,N_3504,N_3978);
nor U4021 (N_4021,N_3325,N_3952);
xnor U4022 (N_4022,N_3763,N_3656);
and U4023 (N_4023,N_3366,N_3793);
xnor U4024 (N_4024,N_3308,N_3744);
nor U4025 (N_4025,N_3652,N_3700);
nor U4026 (N_4026,N_3792,N_3466);
nand U4027 (N_4027,N_3762,N_3292);
nand U4028 (N_4028,N_3365,N_3340);
xor U4029 (N_4029,N_3926,N_3680);
nor U4030 (N_4030,N_3898,N_3737);
xnor U4031 (N_4031,N_3277,N_3956);
nor U4032 (N_4032,N_3991,N_3595);
or U4033 (N_4033,N_3561,N_3773);
or U4034 (N_4034,N_3997,N_3706);
and U4035 (N_4035,N_3672,N_3515);
nand U4036 (N_4036,N_3942,N_3752);
nand U4037 (N_4037,N_3444,N_3441);
nor U4038 (N_4038,N_3688,N_3824);
or U4039 (N_4039,N_3353,N_3713);
xnor U4040 (N_4040,N_3306,N_3804);
nand U4041 (N_4041,N_3897,N_3368);
or U4042 (N_4042,N_3349,N_3859);
nor U4043 (N_4043,N_3470,N_3663);
nor U4044 (N_4044,N_3243,N_3225);
and U4045 (N_4045,N_3920,N_3604);
and U4046 (N_4046,N_3985,N_3704);
xor U4047 (N_4047,N_3878,N_3265);
and U4048 (N_4048,N_3862,N_3969);
nor U4049 (N_4049,N_3312,N_3579);
nand U4050 (N_4050,N_3975,N_3399);
or U4051 (N_4051,N_3838,N_3716);
and U4052 (N_4052,N_3487,N_3778);
or U4053 (N_4053,N_3965,N_3915);
nand U4054 (N_4054,N_3720,N_3735);
or U4055 (N_4055,N_3201,N_3809);
or U4056 (N_4056,N_3469,N_3902);
nand U4057 (N_4057,N_3806,N_3380);
nor U4058 (N_4058,N_3304,N_3315);
nor U4059 (N_4059,N_3632,N_3247);
and U4060 (N_4060,N_3821,N_3275);
nor U4061 (N_4061,N_3414,N_3914);
xnor U4062 (N_4062,N_3831,N_3458);
and U4063 (N_4063,N_3732,N_3291);
nor U4064 (N_4064,N_3733,N_3896);
nor U4065 (N_4065,N_3981,N_3427);
nand U4066 (N_4066,N_3326,N_3760);
and U4067 (N_4067,N_3852,N_3223);
nand U4068 (N_4068,N_3369,N_3381);
and U4069 (N_4069,N_3683,N_3955);
nand U4070 (N_4070,N_3626,N_3238);
or U4071 (N_4071,N_3943,N_3425);
xnor U4072 (N_4072,N_3846,N_3334);
xor U4073 (N_4073,N_3734,N_3547);
xor U4074 (N_4074,N_3511,N_3941);
xnor U4075 (N_4075,N_3830,N_3736);
and U4076 (N_4076,N_3376,N_3933);
nor U4077 (N_4077,N_3320,N_3745);
nor U4078 (N_4078,N_3578,N_3242);
or U4079 (N_4079,N_3437,N_3814);
xnor U4080 (N_4080,N_3577,N_3455);
xnor U4081 (N_4081,N_3257,N_3541);
nor U4082 (N_4082,N_3330,N_3345);
xnor U4083 (N_4083,N_3987,N_3606);
or U4084 (N_4084,N_3298,N_3227);
and U4085 (N_4085,N_3605,N_3880);
or U4086 (N_4086,N_3485,N_3934);
or U4087 (N_4087,N_3241,N_3508);
nor U4088 (N_4088,N_3216,N_3857);
xor U4089 (N_4089,N_3367,N_3299);
nand U4090 (N_4090,N_3749,N_3855);
or U4091 (N_4091,N_3217,N_3373);
or U4092 (N_4092,N_3754,N_3383);
xnor U4093 (N_4093,N_3614,N_3634);
or U4094 (N_4094,N_3507,N_3296);
xor U4095 (N_4095,N_3667,N_3935);
or U4096 (N_4096,N_3769,N_3894);
nand U4097 (N_4097,N_3525,N_3442);
xnor U4098 (N_4098,N_3418,N_3843);
and U4099 (N_4099,N_3601,N_3562);
or U4100 (N_4100,N_3530,N_3213);
and U4101 (N_4101,N_3516,N_3989);
and U4102 (N_4102,N_3833,N_3925);
xnor U4103 (N_4103,N_3903,N_3267);
or U4104 (N_4104,N_3270,N_3839);
or U4105 (N_4105,N_3430,N_3829);
xor U4106 (N_4106,N_3992,N_3725);
nand U4107 (N_4107,N_3641,N_3271);
nor U4108 (N_4108,N_3708,N_3599);
nor U4109 (N_4109,N_3853,N_3653);
nor U4110 (N_4110,N_3401,N_3932);
nand U4111 (N_4111,N_3826,N_3245);
nand U4112 (N_4112,N_3772,N_3260);
xor U4113 (N_4113,N_3959,N_3410);
xor U4114 (N_4114,N_3906,N_3681);
xnor U4115 (N_4115,N_3983,N_3633);
or U4116 (N_4116,N_3502,N_3480);
and U4117 (N_4117,N_3222,N_3813);
nor U4118 (N_4118,N_3538,N_3627);
nor U4119 (N_4119,N_3288,N_3563);
and U4120 (N_4120,N_3553,N_3620);
or U4121 (N_4121,N_3501,N_3726);
nand U4122 (N_4122,N_3479,N_3232);
nor U4123 (N_4123,N_3715,N_3951);
nand U4124 (N_4124,N_3891,N_3347);
or U4125 (N_4125,N_3256,N_3660);
xor U4126 (N_4126,N_3283,N_3348);
nor U4127 (N_4127,N_3422,N_3739);
and U4128 (N_4128,N_3690,N_3486);
and U4129 (N_4129,N_3823,N_3861);
nand U4130 (N_4130,N_3568,N_3436);
or U4131 (N_4131,N_3886,N_3939);
or U4132 (N_4132,N_3864,N_3820);
nand U4133 (N_4133,N_3409,N_3549);
or U4134 (N_4134,N_3753,N_3305);
nand U4135 (N_4135,N_3776,N_3872);
xnor U4136 (N_4136,N_3912,N_3884);
xnor U4137 (N_4137,N_3570,N_3329);
or U4138 (N_4138,N_3473,N_3211);
nor U4139 (N_4139,N_3432,N_3361);
xnor U4140 (N_4140,N_3676,N_3250);
and U4141 (N_4141,N_3755,N_3930);
and U4142 (N_4142,N_3286,N_3865);
nand U4143 (N_4143,N_3384,N_3701);
nor U4144 (N_4144,N_3647,N_3842);
nor U4145 (N_4145,N_3684,N_3335);
xnor U4146 (N_4146,N_3874,N_3481);
xor U4147 (N_4147,N_3678,N_3764);
nand U4148 (N_4148,N_3866,N_3264);
xnor U4149 (N_4149,N_3397,N_3837);
or U4150 (N_4150,N_3822,N_3527);
xor U4151 (N_4151,N_3494,N_3575);
or U4152 (N_4152,N_3729,N_3988);
xnor U4153 (N_4153,N_3451,N_3395);
and U4154 (N_4154,N_3202,N_3537);
nand U4155 (N_4155,N_3832,N_3738);
or U4156 (N_4156,N_3248,N_3583);
or U4157 (N_4157,N_3556,N_3730);
xnor U4158 (N_4158,N_3582,N_3558);
and U4159 (N_4159,N_3311,N_3274);
or U4160 (N_4160,N_3816,N_3597);
and U4161 (N_4161,N_3616,N_3707);
and U4162 (N_4162,N_3477,N_3885);
and U4163 (N_4163,N_3328,N_3757);
xnor U4164 (N_4164,N_3807,N_3293);
nor U4165 (N_4165,N_3927,N_3374);
nand U4166 (N_4166,N_3510,N_3341);
xor U4167 (N_4167,N_3958,N_3351);
and U4168 (N_4168,N_3404,N_3372);
nor U4169 (N_4169,N_3476,N_3869);
or U4170 (N_4170,N_3603,N_3423);
and U4171 (N_4171,N_3518,N_3230);
or U4172 (N_4172,N_3393,N_3608);
nor U4173 (N_4173,N_3966,N_3724);
or U4174 (N_4174,N_3209,N_3559);
xor U4175 (N_4175,N_3836,N_3613);
or U4176 (N_4176,N_3917,N_3767);
nand U4177 (N_4177,N_3908,N_3206);
or U4178 (N_4178,N_3268,N_3825);
xor U4179 (N_4179,N_3565,N_3686);
nor U4180 (N_4180,N_3402,N_3396);
or U4181 (N_4181,N_3482,N_3560);
nand U4182 (N_4182,N_3557,N_3637);
xnor U4183 (N_4183,N_3723,N_3300);
and U4184 (N_4184,N_3623,N_3643);
nor U4185 (N_4185,N_3431,N_3665);
xor U4186 (N_4186,N_3743,N_3937);
and U4187 (N_4187,N_3710,N_3649);
nor U4188 (N_4188,N_3923,N_3948);
or U4189 (N_4189,N_3654,N_3871);
xor U4190 (N_4190,N_3600,N_3835);
nor U4191 (N_4191,N_3779,N_3440);
nor U4192 (N_4192,N_3998,N_3364);
or U4193 (N_4193,N_3635,N_3585);
or U4194 (N_4194,N_3203,N_3931);
xnor U4195 (N_4195,N_3618,N_3666);
xnor U4196 (N_4196,N_3491,N_3717);
nor U4197 (N_4197,N_3587,N_3322);
nand U4198 (N_4198,N_3357,N_3664);
or U4199 (N_4199,N_3574,N_3818);
or U4200 (N_4200,N_3448,N_3791);
xnor U4201 (N_4201,N_3815,N_3858);
nor U4202 (N_4202,N_3674,N_3963);
and U4203 (N_4203,N_3994,N_3790);
or U4204 (N_4204,N_3741,N_3419);
and U4205 (N_4205,N_3798,N_3645);
and U4206 (N_4206,N_3651,N_3503);
and U4207 (N_4207,N_3412,N_3758);
nand U4208 (N_4208,N_3655,N_3911);
xor U4209 (N_4209,N_3233,N_3276);
nor U4210 (N_4210,N_3450,N_3281);
nand U4211 (N_4211,N_3215,N_3982);
nor U4212 (N_4212,N_3533,N_3788);
xor U4213 (N_4213,N_3382,N_3789);
xnor U4214 (N_4214,N_3999,N_3615);
and U4215 (N_4215,N_3851,N_3928);
nand U4216 (N_4216,N_3949,N_3478);
nor U4217 (N_4217,N_3695,N_3593);
xnor U4218 (N_4218,N_3590,N_3475);
nand U4219 (N_4219,N_3840,N_3512);
and U4220 (N_4220,N_3317,N_3868);
nor U4221 (N_4221,N_3536,N_3648);
nand U4222 (N_4222,N_3636,N_3258);
nor U4223 (N_4223,N_3520,N_3234);
nand U4224 (N_4224,N_3882,N_3890);
nor U4225 (N_4225,N_3879,N_3255);
or U4226 (N_4226,N_3658,N_3922);
and U4227 (N_4227,N_3580,N_3554);
or U4228 (N_4228,N_3218,N_3940);
nor U4229 (N_4229,N_3456,N_3889);
nand U4230 (N_4230,N_3214,N_3429);
or U4231 (N_4231,N_3531,N_3331);
xnor U4232 (N_4232,N_3521,N_3787);
or U4233 (N_4233,N_3379,N_3629);
xor U4234 (N_4234,N_3819,N_3411);
and U4235 (N_4235,N_3355,N_3447);
xor U4236 (N_4236,N_3426,N_3498);
and U4237 (N_4237,N_3493,N_3524);
and U4238 (N_4238,N_3343,N_3768);
nand U4239 (N_4239,N_3628,N_3252);
nand U4240 (N_4240,N_3490,N_3204);
xnor U4241 (N_4241,N_3625,N_3698);
nand U4242 (N_4242,N_3619,N_3542);
nor U4243 (N_4243,N_3659,N_3705);
xnor U4244 (N_4244,N_3918,N_3443);
nor U4245 (N_4245,N_3200,N_3433);
and U4246 (N_4246,N_3550,N_3586);
nand U4247 (N_4247,N_3319,N_3513);
and U4248 (N_4248,N_3224,N_3314);
nand U4249 (N_4249,N_3282,N_3237);
xnor U4250 (N_4250,N_3888,N_3460);
xnor U4251 (N_4251,N_3766,N_3468);
xor U4252 (N_4252,N_3362,N_3370);
nand U4253 (N_4253,N_3387,N_3576);
xnor U4254 (N_4254,N_3488,N_3718);
xor U4255 (N_4255,N_3506,N_3385);
nand U4256 (N_4256,N_3971,N_3756);
nand U4257 (N_4257,N_3699,N_3295);
xor U4258 (N_4258,N_3785,N_3679);
and U4259 (N_4259,N_3309,N_3719);
or U4260 (N_4260,N_3728,N_3799);
and U4261 (N_4261,N_3212,N_3848);
or U4262 (N_4262,N_3539,N_3350);
nor U4263 (N_4263,N_3421,N_3463);
xor U4264 (N_4264,N_3548,N_3953);
xor U4265 (N_4265,N_3435,N_3239);
xnor U4266 (N_4266,N_3976,N_3472);
or U4267 (N_4267,N_3621,N_3938);
or U4268 (N_4268,N_3970,N_3904);
nand U4269 (N_4269,N_3428,N_3921);
nand U4270 (N_4270,N_3564,N_3784);
nand U4271 (N_4271,N_3415,N_3555);
xor U4272 (N_4272,N_3413,N_3316);
xor U4273 (N_4273,N_3346,N_3638);
and U4274 (N_4274,N_3406,N_3289);
or U4275 (N_4275,N_3294,N_3205);
or U4276 (N_4276,N_3377,N_3834);
and U4277 (N_4277,N_3417,N_3860);
xor U4278 (N_4278,N_3817,N_3721);
and U4279 (N_4279,N_3913,N_3803);
and U4280 (N_4280,N_3584,N_3572);
or U4281 (N_4281,N_3944,N_3901);
and U4282 (N_4282,N_3474,N_3244);
or U4283 (N_4283,N_3420,N_3356);
or U4284 (N_4284,N_3961,N_3254);
nor U4285 (N_4285,N_3781,N_3573);
nand U4286 (N_4286,N_3811,N_3446);
xor U4287 (N_4287,N_3973,N_3588);
or U4288 (N_4288,N_3893,N_3877);
or U4289 (N_4289,N_3492,N_3386);
and U4290 (N_4290,N_3499,N_3714);
and U4291 (N_4291,N_3774,N_3797);
xnor U4292 (N_4292,N_3876,N_3363);
nor U4293 (N_4293,N_3337,N_3226);
nor U4294 (N_4294,N_3895,N_3747);
and U4295 (N_4295,N_3800,N_3697);
or U4296 (N_4296,N_3529,N_3828);
or U4297 (N_4297,N_3471,N_3313);
nand U4298 (N_4298,N_3307,N_3449);
and U4299 (N_4299,N_3770,N_3727);
nand U4300 (N_4300,N_3854,N_3310);
nand U4301 (N_4301,N_3646,N_3977);
nor U4302 (N_4302,N_3936,N_3229);
xnor U4303 (N_4303,N_3266,N_3235);
and U4304 (N_4304,N_3269,N_3461);
nand U4305 (N_4305,N_3251,N_3360);
nor U4306 (N_4306,N_3602,N_3240);
nand U4307 (N_4307,N_3445,N_3657);
or U4308 (N_4308,N_3517,N_3545);
or U4309 (N_4309,N_3929,N_3543);
and U4310 (N_4310,N_3500,N_3467);
or U4311 (N_4311,N_3694,N_3624);
nor U4312 (N_4312,N_3535,N_3262);
nand U4313 (N_4313,N_3287,N_3540);
or U4314 (N_4314,N_3775,N_3795);
nor U4315 (N_4315,N_3622,N_3974);
and U4316 (N_4316,N_3650,N_3883);
or U4317 (N_4317,N_3640,N_3552);
nor U4318 (N_4318,N_3993,N_3371);
xor U4319 (N_4319,N_3870,N_3592);
xnor U4320 (N_4320,N_3505,N_3263);
xor U4321 (N_4321,N_3297,N_3465);
xnor U4322 (N_4322,N_3711,N_3452);
or U4323 (N_4323,N_3390,N_3391);
or U4324 (N_4324,N_3496,N_3551);
and U4325 (N_4325,N_3761,N_3534);
and U4326 (N_4326,N_3810,N_3327);
or U4327 (N_4327,N_3909,N_3693);
or U4328 (N_4328,N_3301,N_3332);
nand U4329 (N_4329,N_3589,N_3682);
and U4330 (N_4330,N_3454,N_3748);
and U4331 (N_4331,N_3220,N_3668);
nor U4332 (N_4332,N_3709,N_3497);
nand U4333 (N_4333,N_3352,N_3528);
nand U4334 (N_4334,N_3919,N_3990);
xnor U4335 (N_4335,N_3388,N_3273);
xnor U4336 (N_4336,N_3261,N_3867);
xnor U4337 (N_4337,N_3995,N_3669);
xor U4338 (N_4338,N_3812,N_3687);
or U4339 (N_4339,N_3514,N_3324);
nand U4340 (N_4340,N_3794,N_3910);
xor U4341 (N_4341,N_3394,N_3336);
xor U4342 (N_4342,N_3740,N_3712);
nor U4343 (N_4343,N_3546,N_3375);
and U4344 (N_4344,N_3957,N_3210);
xnor U4345 (N_4345,N_3946,N_3285);
nor U4346 (N_4346,N_3321,N_3691);
nand U4347 (N_4347,N_3359,N_3221);
nor U4348 (N_4348,N_3323,N_3892);
nor U4349 (N_4349,N_3907,N_3610);
xor U4350 (N_4350,N_3986,N_3284);
nand U4351 (N_4351,N_3899,N_3392);
and U4352 (N_4352,N_3400,N_3462);
nor U4353 (N_4353,N_3950,N_3453);
nand U4354 (N_4354,N_3786,N_3661);
xnor U4355 (N_4355,N_3962,N_3598);
xnor U4356 (N_4356,N_3702,N_3303);
and U4357 (N_4357,N_3782,N_3249);
and U4358 (N_4358,N_3457,N_3996);
or U4359 (N_4359,N_3416,N_3759);
xnor U4360 (N_4360,N_3662,N_3389);
and U4361 (N_4361,N_3526,N_3208);
and U4362 (N_4362,N_3571,N_3670);
xnor U4363 (N_4363,N_3424,N_3689);
or U4364 (N_4364,N_3405,N_3924);
nor U4365 (N_4365,N_3259,N_3358);
nand U4366 (N_4366,N_3960,N_3280);
nor U4367 (N_4367,N_3863,N_3407);
nor U4368 (N_4368,N_3967,N_3378);
nor U4369 (N_4369,N_3228,N_3464);
xor U4370 (N_4370,N_3642,N_3845);
or U4371 (N_4371,N_3272,N_3408);
nand U4372 (N_4372,N_3231,N_3581);
xnor U4373 (N_4373,N_3611,N_3847);
and U4374 (N_4374,N_3703,N_3339);
nor U4375 (N_4375,N_3219,N_3746);
and U4376 (N_4376,N_3692,N_3338);
or U4377 (N_4377,N_3805,N_3801);
and U4378 (N_4378,N_3569,N_3253);
nand U4379 (N_4379,N_3439,N_3631);
nand U4380 (N_4380,N_3945,N_3630);
and U4381 (N_4381,N_3489,N_3639);
nand U4382 (N_4382,N_3279,N_3954);
nand U4383 (N_4383,N_3771,N_3609);
or U4384 (N_4384,N_3873,N_3947);
xnor U4385 (N_4385,N_3765,N_3984);
xnor U4386 (N_4386,N_3644,N_3751);
nor U4387 (N_4387,N_3844,N_3290);
nor U4388 (N_4388,N_3808,N_3522);
nand U4389 (N_4389,N_3856,N_3342);
and U4390 (N_4390,N_3780,N_3964);
nor U4391 (N_4391,N_3344,N_3302);
nor U4392 (N_4392,N_3802,N_3972);
xor U4393 (N_4393,N_3403,N_3696);
nor U4394 (N_4394,N_3567,N_3916);
or U4395 (N_4395,N_3246,N_3722);
nand U4396 (N_4396,N_3483,N_3459);
and U4397 (N_4397,N_3673,N_3979);
or U4398 (N_4398,N_3519,N_3607);
nor U4399 (N_4399,N_3675,N_3875);
and U4400 (N_4400,N_3546,N_3596);
and U4401 (N_4401,N_3801,N_3429);
nor U4402 (N_4402,N_3856,N_3851);
and U4403 (N_4403,N_3705,N_3224);
and U4404 (N_4404,N_3928,N_3521);
or U4405 (N_4405,N_3362,N_3206);
nor U4406 (N_4406,N_3484,N_3351);
nor U4407 (N_4407,N_3843,N_3817);
or U4408 (N_4408,N_3680,N_3446);
nor U4409 (N_4409,N_3646,N_3501);
and U4410 (N_4410,N_3644,N_3511);
and U4411 (N_4411,N_3490,N_3568);
nand U4412 (N_4412,N_3633,N_3397);
nor U4413 (N_4413,N_3255,N_3552);
xor U4414 (N_4414,N_3568,N_3962);
and U4415 (N_4415,N_3460,N_3865);
nor U4416 (N_4416,N_3568,N_3317);
xor U4417 (N_4417,N_3445,N_3696);
nand U4418 (N_4418,N_3450,N_3651);
and U4419 (N_4419,N_3777,N_3861);
xnor U4420 (N_4420,N_3818,N_3480);
nor U4421 (N_4421,N_3287,N_3955);
xor U4422 (N_4422,N_3938,N_3488);
nor U4423 (N_4423,N_3913,N_3711);
and U4424 (N_4424,N_3249,N_3707);
and U4425 (N_4425,N_3387,N_3379);
nand U4426 (N_4426,N_3717,N_3450);
nor U4427 (N_4427,N_3503,N_3435);
xor U4428 (N_4428,N_3229,N_3849);
and U4429 (N_4429,N_3302,N_3565);
xor U4430 (N_4430,N_3212,N_3962);
xnor U4431 (N_4431,N_3982,N_3730);
xnor U4432 (N_4432,N_3461,N_3441);
or U4433 (N_4433,N_3232,N_3248);
or U4434 (N_4434,N_3322,N_3348);
nor U4435 (N_4435,N_3481,N_3838);
nor U4436 (N_4436,N_3663,N_3571);
or U4437 (N_4437,N_3964,N_3498);
nand U4438 (N_4438,N_3276,N_3632);
and U4439 (N_4439,N_3536,N_3749);
xor U4440 (N_4440,N_3415,N_3761);
or U4441 (N_4441,N_3738,N_3916);
xor U4442 (N_4442,N_3337,N_3796);
nor U4443 (N_4443,N_3854,N_3998);
nor U4444 (N_4444,N_3782,N_3705);
nor U4445 (N_4445,N_3210,N_3397);
xnor U4446 (N_4446,N_3622,N_3303);
or U4447 (N_4447,N_3711,N_3827);
or U4448 (N_4448,N_3804,N_3834);
nand U4449 (N_4449,N_3281,N_3641);
xnor U4450 (N_4450,N_3578,N_3587);
nand U4451 (N_4451,N_3269,N_3299);
nor U4452 (N_4452,N_3617,N_3216);
and U4453 (N_4453,N_3295,N_3561);
nor U4454 (N_4454,N_3352,N_3772);
nand U4455 (N_4455,N_3507,N_3434);
nor U4456 (N_4456,N_3848,N_3293);
xor U4457 (N_4457,N_3908,N_3492);
nand U4458 (N_4458,N_3847,N_3624);
or U4459 (N_4459,N_3745,N_3393);
nor U4460 (N_4460,N_3485,N_3288);
or U4461 (N_4461,N_3640,N_3682);
nor U4462 (N_4462,N_3370,N_3541);
nand U4463 (N_4463,N_3947,N_3269);
and U4464 (N_4464,N_3497,N_3554);
nand U4465 (N_4465,N_3301,N_3482);
xor U4466 (N_4466,N_3338,N_3724);
nor U4467 (N_4467,N_3979,N_3685);
xnor U4468 (N_4468,N_3993,N_3747);
xor U4469 (N_4469,N_3420,N_3807);
or U4470 (N_4470,N_3298,N_3262);
or U4471 (N_4471,N_3308,N_3479);
and U4472 (N_4472,N_3672,N_3869);
xor U4473 (N_4473,N_3587,N_3594);
or U4474 (N_4474,N_3584,N_3301);
xor U4475 (N_4475,N_3826,N_3689);
and U4476 (N_4476,N_3666,N_3261);
nand U4477 (N_4477,N_3798,N_3469);
nor U4478 (N_4478,N_3737,N_3371);
nor U4479 (N_4479,N_3536,N_3675);
nand U4480 (N_4480,N_3271,N_3494);
or U4481 (N_4481,N_3639,N_3930);
nor U4482 (N_4482,N_3641,N_3773);
and U4483 (N_4483,N_3862,N_3565);
nor U4484 (N_4484,N_3935,N_3455);
and U4485 (N_4485,N_3978,N_3378);
and U4486 (N_4486,N_3453,N_3591);
and U4487 (N_4487,N_3643,N_3339);
nand U4488 (N_4488,N_3776,N_3947);
and U4489 (N_4489,N_3641,N_3379);
xor U4490 (N_4490,N_3325,N_3438);
xnor U4491 (N_4491,N_3237,N_3973);
nor U4492 (N_4492,N_3832,N_3210);
or U4493 (N_4493,N_3554,N_3626);
nor U4494 (N_4494,N_3319,N_3657);
nor U4495 (N_4495,N_3540,N_3655);
nand U4496 (N_4496,N_3917,N_3735);
or U4497 (N_4497,N_3949,N_3578);
nor U4498 (N_4498,N_3436,N_3856);
nand U4499 (N_4499,N_3954,N_3913);
xnor U4500 (N_4500,N_3363,N_3751);
xor U4501 (N_4501,N_3801,N_3854);
nand U4502 (N_4502,N_3705,N_3931);
nand U4503 (N_4503,N_3308,N_3228);
nand U4504 (N_4504,N_3421,N_3749);
and U4505 (N_4505,N_3790,N_3341);
xnor U4506 (N_4506,N_3264,N_3257);
and U4507 (N_4507,N_3955,N_3917);
or U4508 (N_4508,N_3768,N_3458);
or U4509 (N_4509,N_3415,N_3570);
nand U4510 (N_4510,N_3818,N_3259);
and U4511 (N_4511,N_3473,N_3611);
nor U4512 (N_4512,N_3903,N_3551);
nor U4513 (N_4513,N_3271,N_3307);
nor U4514 (N_4514,N_3877,N_3948);
xnor U4515 (N_4515,N_3959,N_3628);
nand U4516 (N_4516,N_3526,N_3545);
and U4517 (N_4517,N_3681,N_3546);
and U4518 (N_4518,N_3779,N_3965);
or U4519 (N_4519,N_3977,N_3972);
or U4520 (N_4520,N_3375,N_3532);
nand U4521 (N_4521,N_3723,N_3985);
and U4522 (N_4522,N_3519,N_3358);
or U4523 (N_4523,N_3717,N_3482);
nand U4524 (N_4524,N_3431,N_3572);
or U4525 (N_4525,N_3665,N_3727);
and U4526 (N_4526,N_3400,N_3842);
or U4527 (N_4527,N_3204,N_3465);
nor U4528 (N_4528,N_3369,N_3898);
xor U4529 (N_4529,N_3771,N_3320);
nor U4530 (N_4530,N_3850,N_3906);
nand U4531 (N_4531,N_3910,N_3250);
or U4532 (N_4532,N_3674,N_3552);
or U4533 (N_4533,N_3999,N_3525);
and U4534 (N_4534,N_3366,N_3468);
nor U4535 (N_4535,N_3277,N_3696);
xnor U4536 (N_4536,N_3352,N_3884);
xnor U4537 (N_4537,N_3751,N_3764);
and U4538 (N_4538,N_3320,N_3927);
or U4539 (N_4539,N_3734,N_3640);
xor U4540 (N_4540,N_3655,N_3658);
nor U4541 (N_4541,N_3940,N_3751);
or U4542 (N_4542,N_3677,N_3713);
or U4543 (N_4543,N_3814,N_3963);
xor U4544 (N_4544,N_3910,N_3727);
xor U4545 (N_4545,N_3239,N_3708);
xnor U4546 (N_4546,N_3410,N_3342);
or U4547 (N_4547,N_3957,N_3242);
xnor U4548 (N_4548,N_3522,N_3248);
or U4549 (N_4549,N_3515,N_3342);
xnor U4550 (N_4550,N_3933,N_3331);
xor U4551 (N_4551,N_3413,N_3337);
or U4552 (N_4552,N_3976,N_3720);
and U4553 (N_4553,N_3295,N_3471);
nor U4554 (N_4554,N_3567,N_3314);
nand U4555 (N_4555,N_3522,N_3834);
and U4556 (N_4556,N_3235,N_3865);
or U4557 (N_4557,N_3333,N_3833);
xor U4558 (N_4558,N_3723,N_3724);
nand U4559 (N_4559,N_3430,N_3906);
nand U4560 (N_4560,N_3802,N_3429);
or U4561 (N_4561,N_3272,N_3688);
or U4562 (N_4562,N_3244,N_3798);
and U4563 (N_4563,N_3511,N_3583);
nor U4564 (N_4564,N_3973,N_3415);
nand U4565 (N_4565,N_3766,N_3579);
and U4566 (N_4566,N_3368,N_3410);
and U4567 (N_4567,N_3321,N_3365);
nand U4568 (N_4568,N_3602,N_3593);
nand U4569 (N_4569,N_3667,N_3652);
and U4570 (N_4570,N_3997,N_3369);
and U4571 (N_4571,N_3545,N_3424);
or U4572 (N_4572,N_3296,N_3573);
and U4573 (N_4573,N_3555,N_3456);
and U4574 (N_4574,N_3247,N_3693);
and U4575 (N_4575,N_3447,N_3947);
or U4576 (N_4576,N_3449,N_3462);
and U4577 (N_4577,N_3845,N_3741);
xnor U4578 (N_4578,N_3204,N_3995);
nor U4579 (N_4579,N_3697,N_3527);
and U4580 (N_4580,N_3231,N_3994);
nand U4581 (N_4581,N_3510,N_3979);
or U4582 (N_4582,N_3481,N_3593);
xnor U4583 (N_4583,N_3714,N_3685);
nor U4584 (N_4584,N_3936,N_3768);
or U4585 (N_4585,N_3418,N_3852);
nand U4586 (N_4586,N_3512,N_3905);
xnor U4587 (N_4587,N_3499,N_3219);
nand U4588 (N_4588,N_3205,N_3302);
and U4589 (N_4589,N_3874,N_3310);
nand U4590 (N_4590,N_3889,N_3772);
xnor U4591 (N_4591,N_3354,N_3380);
nor U4592 (N_4592,N_3869,N_3588);
xor U4593 (N_4593,N_3811,N_3404);
and U4594 (N_4594,N_3855,N_3801);
or U4595 (N_4595,N_3227,N_3497);
xnor U4596 (N_4596,N_3750,N_3451);
and U4597 (N_4597,N_3504,N_3498);
nor U4598 (N_4598,N_3341,N_3834);
nor U4599 (N_4599,N_3891,N_3282);
or U4600 (N_4600,N_3350,N_3817);
nor U4601 (N_4601,N_3726,N_3316);
nor U4602 (N_4602,N_3256,N_3339);
xnor U4603 (N_4603,N_3360,N_3866);
or U4604 (N_4604,N_3589,N_3360);
or U4605 (N_4605,N_3516,N_3888);
and U4606 (N_4606,N_3521,N_3474);
nand U4607 (N_4607,N_3951,N_3414);
nor U4608 (N_4608,N_3310,N_3660);
nand U4609 (N_4609,N_3402,N_3524);
and U4610 (N_4610,N_3980,N_3448);
and U4611 (N_4611,N_3359,N_3626);
xnor U4612 (N_4612,N_3726,N_3673);
xor U4613 (N_4613,N_3834,N_3592);
or U4614 (N_4614,N_3538,N_3887);
or U4615 (N_4615,N_3979,N_3636);
nand U4616 (N_4616,N_3268,N_3788);
nand U4617 (N_4617,N_3860,N_3258);
and U4618 (N_4618,N_3271,N_3888);
nor U4619 (N_4619,N_3767,N_3728);
and U4620 (N_4620,N_3277,N_3999);
nand U4621 (N_4621,N_3305,N_3556);
xor U4622 (N_4622,N_3687,N_3576);
or U4623 (N_4623,N_3996,N_3750);
xor U4624 (N_4624,N_3800,N_3449);
nand U4625 (N_4625,N_3341,N_3902);
nand U4626 (N_4626,N_3864,N_3433);
nor U4627 (N_4627,N_3583,N_3741);
and U4628 (N_4628,N_3926,N_3454);
nand U4629 (N_4629,N_3445,N_3461);
or U4630 (N_4630,N_3916,N_3860);
and U4631 (N_4631,N_3791,N_3671);
nor U4632 (N_4632,N_3882,N_3214);
or U4633 (N_4633,N_3502,N_3777);
and U4634 (N_4634,N_3635,N_3424);
or U4635 (N_4635,N_3360,N_3602);
or U4636 (N_4636,N_3573,N_3908);
xnor U4637 (N_4637,N_3601,N_3250);
nor U4638 (N_4638,N_3730,N_3718);
nor U4639 (N_4639,N_3258,N_3857);
xnor U4640 (N_4640,N_3419,N_3796);
nand U4641 (N_4641,N_3689,N_3335);
nor U4642 (N_4642,N_3379,N_3532);
nand U4643 (N_4643,N_3389,N_3285);
or U4644 (N_4644,N_3377,N_3802);
or U4645 (N_4645,N_3729,N_3463);
nand U4646 (N_4646,N_3374,N_3623);
or U4647 (N_4647,N_3572,N_3351);
nand U4648 (N_4648,N_3671,N_3407);
nand U4649 (N_4649,N_3876,N_3371);
nor U4650 (N_4650,N_3452,N_3684);
and U4651 (N_4651,N_3390,N_3310);
nor U4652 (N_4652,N_3394,N_3635);
or U4653 (N_4653,N_3265,N_3613);
nand U4654 (N_4654,N_3205,N_3423);
nor U4655 (N_4655,N_3401,N_3843);
xor U4656 (N_4656,N_3924,N_3279);
nand U4657 (N_4657,N_3403,N_3481);
nand U4658 (N_4658,N_3211,N_3435);
nor U4659 (N_4659,N_3633,N_3319);
nor U4660 (N_4660,N_3225,N_3726);
xnor U4661 (N_4661,N_3225,N_3434);
xor U4662 (N_4662,N_3386,N_3583);
and U4663 (N_4663,N_3752,N_3458);
xor U4664 (N_4664,N_3916,N_3294);
xor U4665 (N_4665,N_3860,N_3865);
xnor U4666 (N_4666,N_3421,N_3791);
or U4667 (N_4667,N_3862,N_3246);
nor U4668 (N_4668,N_3457,N_3292);
or U4669 (N_4669,N_3489,N_3633);
xor U4670 (N_4670,N_3521,N_3625);
and U4671 (N_4671,N_3929,N_3677);
xor U4672 (N_4672,N_3437,N_3468);
xnor U4673 (N_4673,N_3815,N_3374);
xor U4674 (N_4674,N_3797,N_3280);
and U4675 (N_4675,N_3990,N_3967);
xor U4676 (N_4676,N_3505,N_3413);
nor U4677 (N_4677,N_3208,N_3868);
nor U4678 (N_4678,N_3849,N_3449);
or U4679 (N_4679,N_3384,N_3799);
xor U4680 (N_4680,N_3485,N_3947);
and U4681 (N_4681,N_3210,N_3956);
or U4682 (N_4682,N_3596,N_3389);
or U4683 (N_4683,N_3612,N_3526);
nand U4684 (N_4684,N_3524,N_3483);
or U4685 (N_4685,N_3617,N_3828);
and U4686 (N_4686,N_3789,N_3507);
or U4687 (N_4687,N_3290,N_3262);
or U4688 (N_4688,N_3505,N_3742);
nor U4689 (N_4689,N_3432,N_3385);
and U4690 (N_4690,N_3500,N_3622);
nor U4691 (N_4691,N_3421,N_3644);
and U4692 (N_4692,N_3619,N_3486);
and U4693 (N_4693,N_3872,N_3346);
nand U4694 (N_4694,N_3475,N_3716);
xor U4695 (N_4695,N_3681,N_3900);
xnor U4696 (N_4696,N_3442,N_3926);
nor U4697 (N_4697,N_3631,N_3258);
and U4698 (N_4698,N_3231,N_3264);
or U4699 (N_4699,N_3610,N_3638);
or U4700 (N_4700,N_3987,N_3711);
nand U4701 (N_4701,N_3357,N_3496);
xnor U4702 (N_4702,N_3615,N_3439);
xnor U4703 (N_4703,N_3375,N_3630);
or U4704 (N_4704,N_3974,N_3220);
nor U4705 (N_4705,N_3753,N_3399);
and U4706 (N_4706,N_3710,N_3229);
nor U4707 (N_4707,N_3556,N_3387);
nor U4708 (N_4708,N_3697,N_3568);
and U4709 (N_4709,N_3291,N_3774);
or U4710 (N_4710,N_3424,N_3268);
nand U4711 (N_4711,N_3773,N_3924);
or U4712 (N_4712,N_3680,N_3818);
and U4713 (N_4713,N_3892,N_3475);
and U4714 (N_4714,N_3495,N_3234);
xor U4715 (N_4715,N_3260,N_3939);
nand U4716 (N_4716,N_3636,N_3847);
or U4717 (N_4717,N_3807,N_3663);
nor U4718 (N_4718,N_3854,N_3688);
xor U4719 (N_4719,N_3528,N_3958);
xnor U4720 (N_4720,N_3727,N_3389);
xor U4721 (N_4721,N_3286,N_3647);
nand U4722 (N_4722,N_3675,N_3454);
xor U4723 (N_4723,N_3806,N_3667);
nand U4724 (N_4724,N_3546,N_3732);
nor U4725 (N_4725,N_3259,N_3307);
xnor U4726 (N_4726,N_3467,N_3936);
xnor U4727 (N_4727,N_3658,N_3294);
and U4728 (N_4728,N_3897,N_3469);
or U4729 (N_4729,N_3966,N_3744);
nor U4730 (N_4730,N_3620,N_3660);
nand U4731 (N_4731,N_3829,N_3271);
and U4732 (N_4732,N_3946,N_3661);
and U4733 (N_4733,N_3209,N_3233);
nand U4734 (N_4734,N_3290,N_3959);
or U4735 (N_4735,N_3648,N_3224);
or U4736 (N_4736,N_3815,N_3224);
nor U4737 (N_4737,N_3622,N_3260);
xor U4738 (N_4738,N_3738,N_3202);
xor U4739 (N_4739,N_3997,N_3268);
nor U4740 (N_4740,N_3602,N_3580);
and U4741 (N_4741,N_3745,N_3443);
nand U4742 (N_4742,N_3361,N_3276);
xor U4743 (N_4743,N_3719,N_3803);
and U4744 (N_4744,N_3269,N_3796);
xnor U4745 (N_4745,N_3727,N_3225);
xnor U4746 (N_4746,N_3747,N_3704);
or U4747 (N_4747,N_3851,N_3502);
nand U4748 (N_4748,N_3435,N_3420);
xnor U4749 (N_4749,N_3500,N_3715);
and U4750 (N_4750,N_3470,N_3503);
and U4751 (N_4751,N_3876,N_3375);
nand U4752 (N_4752,N_3804,N_3875);
and U4753 (N_4753,N_3683,N_3988);
or U4754 (N_4754,N_3229,N_3933);
nor U4755 (N_4755,N_3735,N_3314);
xor U4756 (N_4756,N_3519,N_3934);
and U4757 (N_4757,N_3980,N_3665);
or U4758 (N_4758,N_3539,N_3351);
and U4759 (N_4759,N_3739,N_3908);
xnor U4760 (N_4760,N_3504,N_3731);
and U4761 (N_4761,N_3696,N_3900);
xnor U4762 (N_4762,N_3701,N_3523);
nand U4763 (N_4763,N_3992,N_3344);
xnor U4764 (N_4764,N_3850,N_3904);
nand U4765 (N_4765,N_3788,N_3589);
nand U4766 (N_4766,N_3722,N_3480);
nor U4767 (N_4767,N_3275,N_3681);
or U4768 (N_4768,N_3525,N_3602);
and U4769 (N_4769,N_3267,N_3227);
nor U4770 (N_4770,N_3237,N_3917);
xor U4771 (N_4771,N_3447,N_3883);
xnor U4772 (N_4772,N_3279,N_3732);
and U4773 (N_4773,N_3727,N_3871);
and U4774 (N_4774,N_3397,N_3385);
nor U4775 (N_4775,N_3814,N_3528);
nand U4776 (N_4776,N_3970,N_3354);
nand U4777 (N_4777,N_3342,N_3242);
nand U4778 (N_4778,N_3803,N_3830);
or U4779 (N_4779,N_3265,N_3252);
xor U4780 (N_4780,N_3840,N_3564);
nor U4781 (N_4781,N_3561,N_3237);
nor U4782 (N_4782,N_3501,N_3810);
nor U4783 (N_4783,N_3402,N_3772);
or U4784 (N_4784,N_3746,N_3647);
xnor U4785 (N_4785,N_3845,N_3721);
nor U4786 (N_4786,N_3974,N_3244);
nor U4787 (N_4787,N_3720,N_3248);
or U4788 (N_4788,N_3758,N_3701);
nand U4789 (N_4789,N_3813,N_3680);
and U4790 (N_4790,N_3932,N_3373);
or U4791 (N_4791,N_3829,N_3551);
and U4792 (N_4792,N_3799,N_3453);
or U4793 (N_4793,N_3934,N_3437);
and U4794 (N_4794,N_3961,N_3410);
or U4795 (N_4795,N_3310,N_3422);
nand U4796 (N_4796,N_3786,N_3604);
nand U4797 (N_4797,N_3438,N_3850);
or U4798 (N_4798,N_3920,N_3570);
xor U4799 (N_4799,N_3854,N_3799);
nand U4800 (N_4800,N_4042,N_4354);
xor U4801 (N_4801,N_4716,N_4294);
and U4802 (N_4802,N_4481,N_4761);
xnor U4803 (N_4803,N_4231,N_4096);
nor U4804 (N_4804,N_4623,N_4588);
xor U4805 (N_4805,N_4631,N_4023);
nor U4806 (N_4806,N_4007,N_4678);
and U4807 (N_4807,N_4650,N_4253);
xnor U4808 (N_4808,N_4159,N_4664);
nand U4809 (N_4809,N_4649,N_4302);
xnor U4810 (N_4810,N_4483,N_4503);
and U4811 (N_4811,N_4757,N_4372);
nand U4812 (N_4812,N_4728,N_4148);
xor U4813 (N_4813,N_4699,N_4085);
nor U4814 (N_4814,N_4020,N_4144);
nor U4815 (N_4815,N_4622,N_4250);
nor U4816 (N_4816,N_4799,N_4292);
nor U4817 (N_4817,N_4127,N_4640);
xor U4818 (N_4818,N_4666,N_4457);
xor U4819 (N_4819,N_4154,N_4196);
and U4820 (N_4820,N_4143,N_4531);
xnor U4821 (N_4821,N_4347,N_4610);
and U4822 (N_4822,N_4073,N_4165);
or U4823 (N_4823,N_4095,N_4147);
nand U4824 (N_4824,N_4319,N_4743);
nor U4825 (N_4825,N_4104,N_4018);
xor U4826 (N_4826,N_4607,N_4193);
nand U4827 (N_4827,N_4512,N_4580);
and U4828 (N_4828,N_4459,N_4507);
xor U4829 (N_4829,N_4390,N_4693);
or U4830 (N_4830,N_4792,N_4222);
nand U4831 (N_4831,N_4199,N_4052);
xor U4832 (N_4832,N_4557,N_4476);
or U4833 (N_4833,N_4489,N_4167);
or U4834 (N_4834,N_4559,N_4269);
nor U4835 (N_4835,N_4209,N_4644);
nor U4836 (N_4836,N_4415,N_4658);
and U4837 (N_4837,N_4471,N_4609);
nand U4838 (N_4838,N_4194,N_4352);
or U4839 (N_4839,N_4564,N_4568);
or U4840 (N_4840,N_4139,N_4674);
nor U4841 (N_4841,N_4562,N_4395);
or U4842 (N_4842,N_4525,N_4560);
or U4843 (N_4843,N_4259,N_4326);
nor U4844 (N_4844,N_4594,N_4409);
xnor U4845 (N_4845,N_4331,N_4472);
xnor U4846 (N_4846,N_4175,N_4389);
or U4847 (N_4847,N_4388,N_4367);
nor U4848 (N_4848,N_4432,N_4092);
and U4849 (N_4849,N_4789,N_4592);
or U4850 (N_4850,N_4318,N_4323);
and U4851 (N_4851,N_4527,N_4405);
nor U4852 (N_4852,N_4549,N_4229);
or U4853 (N_4853,N_4279,N_4463);
or U4854 (N_4854,N_4673,N_4049);
and U4855 (N_4855,N_4679,N_4083);
or U4856 (N_4856,N_4293,N_4370);
and U4857 (N_4857,N_4638,N_4698);
nand U4858 (N_4858,N_4363,N_4730);
nor U4859 (N_4859,N_4455,N_4060);
and U4860 (N_4860,N_4100,N_4101);
and U4861 (N_4861,N_4702,N_4632);
xor U4862 (N_4862,N_4106,N_4039);
and U4863 (N_4863,N_4089,N_4791);
and U4864 (N_4864,N_4569,N_4627);
and U4865 (N_4865,N_4449,N_4747);
nand U4866 (N_4866,N_4491,N_4350);
or U4867 (N_4867,N_4080,N_4377);
and U4868 (N_4868,N_4307,N_4320);
or U4869 (N_4869,N_4171,N_4027);
nand U4870 (N_4870,N_4133,N_4735);
nor U4871 (N_4871,N_4308,N_4356);
nand U4872 (N_4872,N_4493,N_4335);
xnor U4873 (N_4873,N_4671,N_4461);
nand U4874 (N_4874,N_4176,N_4777);
nor U4875 (N_4875,N_4291,N_4164);
or U4876 (N_4876,N_4305,N_4474);
and U4877 (N_4877,N_4152,N_4538);
xor U4878 (N_4878,N_4097,N_4517);
nand U4879 (N_4879,N_4417,N_4346);
nand U4880 (N_4880,N_4072,N_4620);
and U4881 (N_4881,N_4540,N_4412);
nand U4882 (N_4882,N_4486,N_4442);
xor U4883 (N_4883,N_4779,N_4379);
nand U4884 (N_4884,N_4059,N_4450);
nor U4885 (N_4885,N_4603,N_4077);
nor U4886 (N_4886,N_4636,N_4391);
and U4887 (N_4887,N_4286,N_4596);
nand U4888 (N_4888,N_4197,N_4754);
or U4889 (N_4889,N_4396,N_4581);
nand U4890 (N_4890,N_4790,N_4753);
nor U4891 (N_4891,N_4465,N_4469);
xnor U4892 (N_4892,N_4103,N_4187);
or U4893 (N_4893,N_4445,N_4502);
nor U4894 (N_4894,N_4722,N_4136);
and U4895 (N_4895,N_4715,N_4506);
and U4896 (N_4896,N_4665,N_4254);
xnor U4897 (N_4897,N_4621,N_4441);
nand U4898 (N_4898,N_4499,N_4251);
nor U4899 (N_4899,N_4773,N_4265);
and U4900 (N_4900,N_4266,N_4076);
xor U4901 (N_4901,N_4212,N_4706);
and U4902 (N_4902,N_4374,N_4583);
nor U4903 (N_4903,N_4301,N_4659);
or U4904 (N_4904,N_4406,N_4119);
or U4905 (N_4905,N_4386,N_4227);
and U4906 (N_4906,N_4672,N_4282);
nand U4907 (N_4907,N_4695,N_4509);
nand U4908 (N_4908,N_4545,N_4566);
nand U4909 (N_4909,N_4703,N_4794);
nand U4910 (N_4910,N_4369,N_4273);
nor U4911 (N_4911,N_4694,N_4578);
xnor U4912 (N_4912,N_4008,N_4041);
nand U4913 (N_4913,N_4189,N_4132);
nor U4914 (N_4914,N_4543,N_4551);
nand U4915 (N_4915,N_4523,N_4263);
or U4916 (N_4916,N_4121,N_4242);
nor U4917 (N_4917,N_4032,N_4344);
xor U4918 (N_4918,N_4456,N_4516);
nor U4919 (N_4919,N_4070,N_4325);
nand U4920 (N_4920,N_4797,N_4230);
nand U4921 (N_4921,N_4107,N_4040);
xor U4922 (N_4922,N_4138,N_4487);
and U4923 (N_4923,N_4524,N_4561);
or U4924 (N_4924,N_4030,N_4676);
and U4925 (N_4925,N_4198,N_4241);
nand U4926 (N_4926,N_4641,N_4563);
nor U4927 (N_4927,N_4435,N_4394);
and U4928 (N_4928,N_4741,N_4422);
nor U4929 (N_4929,N_4739,N_4793);
and U4930 (N_4930,N_4084,N_4617);
xnor U4931 (N_4931,N_4764,N_4766);
nor U4932 (N_4932,N_4093,N_4012);
nor U4933 (N_4933,N_4324,N_4683);
nand U4934 (N_4934,N_4329,N_4166);
nor U4935 (N_4935,N_4190,N_4338);
nor U4936 (N_4936,N_4750,N_4726);
and U4937 (N_4937,N_4724,N_4454);
xor U4938 (N_4938,N_4718,N_4280);
and U4939 (N_4939,N_4003,N_4289);
xnor U4940 (N_4940,N_4629,N_4590);
nor U4941 (N_4941,N_4426,N_4208);
and U4942 (N_4942,N_4633,N_4428);
xnor U4943 (N_4943,N_4383,N_4238);
nand U4944 (N_4944,N_4772,N_4371);
nor U4945 (N_4945,N_4400,N_4321);
nor U4946 (N_4946,N_4734,N_4157);
or U4947 (N_4947,N_4274,N_4351);
or U4948 (N_4948,N_4360,N_4681);
or U4949 (N_4949,N_4662,N_4717);
or U4950 (N_4950,N_4556,N_4425);
and U4951 (N_4951,N_4542,N_4221);
xnor U4952 (N_4952,N_4539,N_4243);
and U4953 (N_4953,N_4498,N_4290);
nand U4954 (N_4954,N_4206,N_4065);
nor U4955 (N_4955,N_4480,N_4785);
nor U4956 (N_4956,N_4168,N_4494);
nand U4957 (N_4957,N_4174,N_4748);
and U4958 (N_4958,N_4366,N_4156);
nand U4959 (N_4959,N_4223,N_4408);
nand U4960 (N_4960,N_4200,N_4054);
and U4961 (N_4961,N_4576,N_4064);
and U4962 (N_4962,N_4648,N_4098);
nand U4963 (N_4963,N_4670,N_4186);
nor U4964 (N_4964,N_4645,N_4439);
and U4965 (N_4965,N_4034,N_4384);
or U4966 (N_4966,N_4146,N_4142);
nand U4967 (N_4967,N_4765,N_4532);
or U4968 (N_4968,N_4605,N_4654);
nor U4969 (N_4969,N_4047,N_4236);
nor U4970 (N_4970,N_4416,N_4541);
nor U4971 (N_4971,N_4604,N_4528);
and U4972 (N_4972,N_4205,N_4704);
xor U4973 (N_4973,N_4624,N_4399);
or U4974 (N_4974,N_4262,N_4711);
nor U4975 (N_4975,N_4029,N_4057);
nor U4976 (N_4976,N_4075,N_4546);
nor U4977 (N_4977,N_4213,N_4477);
xor U4978 (N_4978,N_4697,N_4710);
nor U4979 (N_4979,N_4690,N_4519);
and U4980 (N_4980,N_4462,N_4210);
and U4981 (N_4981,N_4062,N_4179);
nor U4982 (N_4982,N_4478,N_4550);
or U4983 (N_4983,N_4071,N_4207);
nand U4984 (N_4984,N_4767,N_4732);
nor U4985 (N_4985,N_4203,N_4705);
and U4986 (N_4986,N_4284,N_4028);
nand U4987 (N_4987,N_4783,N_4501);
nor U4988 (N_4988,N_4328,N_4191);
and U4989 (N_4989,N_4736,N_4429);
and U4990 (N_4990,N_4411,N_4050);
and U4991 (N_4991,N_4482,N_4567);
and U4992 (N_4992,N_4788,N_4019);
nor U4993 (N_4993,N_4586,N_4385);
nor U4994 (N_4994,N_4714,N_4744);
nand U4995 (N_4995,N_4689,N_4602);
or U4996 (N_4996,N_4033,N_4639);
nor U4997 (N_4997,N_4402,N_4087);
nand U4998 (N_4998,N_4696,N_4233);
xnor U4999 (N_4999,N_4088,N_4466);
nand U5000 (N_5000,N_4646,N_4036);
or U5001 (N_5001,N_4283,N_4656);
nor U5002 (N_5002,N_4615,N_4781);
nor U5003 (N_5003,N_4061,N_4460);
nand U5004 (N_5004,N_4359,N_4264);
nand U5005 (N_5005,N_4109,N_4163);
nand U5006 (N_5006,N_4270,N_4513);
xnor U5007 (N_5007,N_4520,N_4045);
xor U5008 (N_5008,N_4745,N_4332);
or U5009 (N_5009,N_4358,N_4544);
nand U5010 (N_5010,N_4521,N_4642);
xor U5011 (N_5011,N_4635,N_4118);
and U5012 (N_5012,N_4473,N_4117);
xnor U5013 (N_5013,N_4496,N_4063);
nor U5014 (N_5014,N_4306,N_4081);
or U5015 (N_5015,N_4733,N_4130);
xnor U5016 (N_5016,N_4484,N_4184);
nor U5017 (N_5017,N_4558,N_4468);
nand U5018 (N_5018,N_4091,N_4720);
nor U5019 (N_5019,N_4625,N_4614);
nor U5020 (N_5020,N_4701,N_4452);
nor U5021 (N_5021,N_4414,N_4267);
or U5022 (N_5022,N_4464,N_4719);
xor U5023 (N_5023,N_4613,N_4707);
nor U5024 (N_5024,N_4214,N_4756);
and U5025 (N_5025,N_4006,N_4522);
nand U5026 (N_5026,N_4573,N_4303);
and U5027 (N_5027,N_4407,N_4158);
nor U5028 (N_5028,N_4505,N_4099);
or U5029 (N_5029,N_4239,N_4479);
or U5030 (N_5030,N_4141,N_4271);
and U5031 (N_5031,N_4255,N_4224);
and U5032 (N_5032,N_4288,N_4295);
nor U5033 (N_5033,N_4444,N_4608);
and U5034 (N_5034,N_4630,N_4298);
nor U5035 (N_5035,N_4069,N_4795);
nand U5036 (N_5036,N_4713,N_4433);
or U5037 (N_5037,N_4430,N_4067);
or U5038 (N_5038,N_4552,N_4131);
or U5039 (N_5039,N_4438,N_4181);
nand U5040 (N_5040,N_4322,N_4774);
nor U5041 (N_5041,N_4110,N_4361);
or U5042 (N_5042,N_4137,N_4688);
or U5043 (N_5043,N_4046,N_4637);
and U5044 (N_5044,N_4074,N_4111);
and U5045 (N_5045,N_4443,N_4490);
nand U5046 (N_5046,N_4281,N_4277);
nor U5047 (N_5047,N_4188,N_4185);
xnor U5048 (N_5048,N_4312,N_4330);
nor U5049 (N_5049,N_4125,N_4353);
nor U5050 (N_5050,N_4285,N_4170);
nand U5051 (N_5051,N_4304,N_4579);
nand U5052 (N_5052,N_4025,N_4173);
xnor U5053 (N_5053,N_4066,N_4013);
and U5054 (N_5054,N_4378,N_4218);
and U5055 (N_5055,N_4548,N_4037);
and U5056 (N_5056,N_4112,N_4183);
and U5057 (N_5057,N_4009,N_4628);
nor U5058 (N_5058,N_4453,N_4192);
nand U5059 (N_5059,N_4348,N_4577);
nand U5060 (N_5060,N_4599,N_4404);
and U5061 (N_5061,N_4235,N_4553);
nor U5062 (N_5062,N_4446,N_4740);
or U5063 (N_5063,N_4217,N_4387);
xnor U5064 (N_5064,N_4780,N_4510);
nand U5065 (N_5065,N_4297,N_4169);
xnor U5066 (N_5066,N_4226,N_4763);
and U5067 (N_5067,N_4752,N_4220);
and U5068 (N_5068,N_4458,N_4150);
nor U5069 (N_5069,N_4078,N_4016);
xor U5070 (N_5070,N_4675,N_4669);
nor U5071 (N_5071,N_4434,N_4436);
and U5072 (N_5072,N_4355,N_4215);
nor U5073 (N_5073,N_4260,N_4368);
or U5074 (N_5074,N_4145,N_4655);
or U5075 (N_5075,N_4587,N_4643);
nand U5076 (N_5076,N_4742,N_4612);
xor U5077 (N_5077,N_4668,N_4014);
or U5078 (N_5078,N_4575,N_4011);
xnor U5079 (N_5079,N_4300,N_4467);
xor U5080 (N_5080,N_4334,N_4336);
or U5081 (N_5081,N_4775,N_4657);
and U5082 (N_5082,N_4258,N_4272);
nand U5083 (N_5083,N_4341,N_4245);
and U5084 (N_5084,N_4015,N_4626);
nand U5085 (N_5085,N_4031,N_4349);
nand U5086 (N_5086,N_4392,N_4122);
or U5087 (N_5087,N_4035,N_4339);
or U5088 (N_5088,N_4682,N_4533);
nor U5089 (N_5089,N_4364,N_4410);
nand U5090 (N_5090,N_4309,N_4237);
nand U5091 (N_5091,N_4616,N_4002);
xor U5092 (N_5092,N_4381,N_4677);
and U5093 (N_5093,N_4114,N_4086);
nor U5094 (N_5094,N_4619,N_4079);
and U5095 (N_5095,N_4327,N_4153);
nor U5096 (N_5096,N_4749,N_4504);
nor U5097 (N_5097,N_4005,N_4149);
nand U5098 (N_5098,N_4337,N_4535);
xor U5099 (N_5099,N_4204,N_4058);
xor U5100 (N_5100,N_4500,N_4043);
nand U5101 (N_5101,N_4311,N_4762);
and U5102 (N_5102,N_4424,N_4257);
nor U5103 (N_5103,N_4299,N_4345);
and U5104 (N_5104,N_4249,N_4684);
nor U5105 (N_5105,N_4128,N_4554);
or U5106 (N_5106,N_4514,N_4437);
nand U5107 (N_5107,N_4782,N_4240);
or U5108 (N_5108,N_4247,N_4447);
and U5109 (N_5109,N_4140,N_4000);
xnor U5110 (N_5110,N_4090,N_4151);
nand U5111 (N_5111,N_4228,N_4536);
nand U5112 (N_5112,N_4182,N_4343);
or U5113 (N_5113,N_4180,N_4278);
nand U5114 (N_5114,N_4252,N_4663);
xnor U5115 (N_5115,N_4310,N_4102);
xnor U5116 (N_5116,N_4244,N_4518);
nor U5117 (N_5117,N_4248,N_4511);
and U5118 (N_5118,N_4155,N_4373);
nand U5119 (N_5119,N_4547,N_4618);
and U5120 (N_5120,N_4022,N_4124);
nor U5121 (N_5121,N_4776,N_4202);
nand U5122 (N_5122,N_4001,N_4232);
xnor U5123 (N_5123,N_4729,N_4094);
nand U5124 (N_5124,N_4448,N_4647);
or U5125 (N_5125,N_4055,N_4275);
nand U5126 (N_5126,N_4420,N_4485);
xnor U5127 (N_5127,N_4760,N_4771);
and U5128 (N_5128,N_4314,N_4634);
nand U5129 (N_5129,N_4796,N_4113);
xnor U5130 (N_5130,N_4686,N_4082);
or U5131 (N_5131,N_4600,N_4401);
or U5132 (N_5132,N_4529,N_4606);
and U5133 (N_5133,N_4423,N_4598);
or U5134 (N_5134,N_4440,N_4362);
nand U5135 (N_5135,N_4727,N_4526);
and U5136 (N_5136,N_4162,N_4570);
nor U5137 (N_5137,N_4708,N_4584);
xor U5138 (N_5138,N_4397,N_4555);
and U5139 (N_5139,N_4010,N_4571);
nand U5140 (N_5140,N_4123,N_4115);
nor U5141 (N_5141,N_4768,N_4530);
xor U5142 (N_5142,N_4611,N_4135);
or U5143 (N_5143,N_4365,N_4725);
xnor U5144 (N_5144,N_4585,N_4161);
and U5145 (N_5145,N_4316,N_4056);
nor U5146 (N_5146,N_4313,N_4759);
nor U5147 (N_5147,N_4017,N_4475);
nor U5148 (N_5148,N_4709,N_4201);
and U5149 (N_5149,N_4692,N_4652);
nand U5150 (N_5150,N_4582,N_4296);
and U5151 (N_5151,N_4376,N_4680);
xor U5152 (N_5152,N_4256,N_4340);
or U5153 (N_5153,N_4382,N_4225);
xor U5154 (N_5154,N_4660,N_4534);
or U5155 (N_5155,N_4246,N_4403);
or U5156 (N_5156,N_4287,N_4195);
and U5157 (N_5157,N_4357,N_4451);
nor U5158 (N_5158,N_4755,N_4268);
or U5159 (N_5159,N_4597,N_4778);
and U5160 (N_5160,N_4026,N_4770);
nand U5161 (N_5161,N_4427,N_4787);
nor U5162 (N_5162,N_4492,N_4134);
or U5163 (N_5163,N_4784,N_4172);
nand U5164 (N_5164,N_4421,N_4413);
xor U5165 (N_5165,N_4601,N_4431);
nand U5166 (N_5166,N_4572,N_4068);
nor U5167 (N_5167,N_4048,N_4653);
nor U5168 (N_5168,N_4315,N_4418);
or U5169 (N_5169,N_4591,N_4751);
xnor U5170 (N_5170,N_4691,N_4574);
or U5171 (N_5171,N_4234,N_4798);
or U5172 (N_5172,N_4595,N_4160);
and U5173 (N_5173,N_4105,N_4024);
xor U5174 (N_5174,N_4342,N_4508);
and U5175 (N_5175,N_4053,N_4700);
and U5176 (N_5176,N_4178,N_4687);
and U5177 (N_5177,N_4565,N_4723);
and U5178 (N_5178,N_4116,N_4380);
or U5179 (N_5179,N_4667,N_4515);
nand U5180 (N_5180,N_4758,N_4333);
and U5181 (N_5181,N_4177,N_4712);
or U5182 (N_5182,N_4593,N_4261);
nor U5183 (N_5183,N_4470,N_4276);
nor U5184 (N_5184,N_4393,N_4661);
nand U5185 (N_5185,N_4317,N_4051);
nand U5186 (N_5186,N_4129,N_4126);
or U5187 (N_5187,N_4419,N_4021);
and U5188 (N_5188,N_4721,N_4488);
nand U5189 (N_5189,N_4038,N_4004);
or U5190 (N_5190,N_4219,N_4537);
or U5191 (N_5191,N_4495,N_4738);
or U5192 (N_5192,N_4731,N_4651);
or U5193 (N_5193,N_4375,N_4211);
nand U5194 (N_5194,N_4497,N_4746);
nor U5195 (N_5195,N_4120,N_4589);
nand U5196 (N_5196,N_4044,N_4216);
and U5197 (N_5197,N_4685,N_4108);
and U5198 (N_5198,N_4398,N_4786);
nand U5199 (N_5199,N_4737,N_4769);
and U5200 (N_5200,N_4368,N_4060);
or U5201 (N_5201,N_4069,N_4454);
or U5202 (N_5202,N_4303,N_4506);
or U5203 (N_5203,N_4695,N_4445);
nor U5204 (N_5204,N_4218,N_4665);
or U5205 (N_5205,N_4600,N_4273);
xor U5206 (N_5206,N_4197,N_4209);
nand U5207 (N_5207,N_4458,N_4305);
or U5208 (N_5208,N_4130,N_4109);
nor U5209 (N_5209,N_4720,N_4578);
or U5210 (N_5210,N_4513,N_4680);
and U5211 (N_5211,N_4574,N_4316);
nor U5212 (N_5212,N_4206,N_4692);
nand U5213 (N_5213,N_4758,N_4345);
nor U5214 (N_5214,N_4544,N_4089);
and U5215 (N_5215,N_4345,N_4681);
nor U5216 (N_5216,N_4279,N_4097);
xnor U5217 (N_5217,N_4771,N_4671);
xnor U5218 (N_5218,N_4001,N_4291);
and U5219 (N_5219,N_4439,N_4785);
and U5220 (N_5220,N_4441,N_4528);
or U5221 (N_5221,N_4033,N_4531);
xnor U5222 (N_5222,N_4771,N_4419);
nor U5223 (N_5223,N_4650,N_4301);
xnor U5224 (N_5224,N_4794,N_4049);
and U5225 (N_5225,N_4735,N_4480);
and U5226 (N_5226,N_4511,N_4169);
or U5227 (N_5227,N_4762,N_4014);
xor U5228 (N_5228,N_4310,N_4599);
and U5229 (N_5229,N_4452,N_4538);
nand U5230 (N_5230,N_4595,N_4090);
nand U5231 (N_5231,N_4216,N_4039);
or U5232 (N_5232,N_4102,N_4194);
nand U5233 (N_5233,N_4060,N_4001);
and U5234 (N_5234,N_4576,N_4532);
and U5235 (N_5235,N_4772,N_4103);
xor U5236 (N_5236,N_4545,N_4642);
or U5237 (N_5237,N_4589,N_4692);
or U5238 (N_5238,N_4455,N_4508);
or U5239 (N_5239,N_4162,N_4251);
or U5240 (N_5240,N_4523,N_4319);
nand U5241 (N_5241,N_4129,N_4299);
nand U5242 (N_5242,N_4761,N_4416);
nand U5243 (N_5243,N_4685,N_4311);
or U5244 (N_5244,N_4118,N_4198);
xnor U5245 (N_5245,N_4497,N_4020);
or U5246 (N_5246,N_4798,N_4220);
nand U5247 (N_5247,N_4152,N_4208);
nor U5248 (N_5248,N_4149,N_4128);
nand U5249 (N_5249,N_4382,N_4008);
and U5250 (N_5250,N_4222,N_4240);
nor U5251 (N_5251,N_4505,N_4423);
and U5252 (N_5252,N_4764,N_4251);
or U5253 (N_5253,N_4053,N_4263);
xnor U5254 (N_5254,N_4342,N_4253);
nor U5255 (N_5255,N_4363,N_4018);
nand U5256 (N_5256,N_4290,N_4782);
nand U5257 (N_5257,N_4524,N_4233);
or U5258 (N_5258,N_4175,N_4268);
xnor U5259 (N_5259,N_4768,N_4634);
and U5260 (N_5260,N_4188,N_4462);
nand U5261 (N_5261,N_4086,N_4731);
nor U5262 (N_5262,N_4635,N_4218);
and U5263 (N_5263,N_4551,N_4297);
xor U5264 (N_5264,N_4759,N_4294);
nor U5265 (N_5265,N_4470,N_4393);
and U5266 (N_5266,N_4323,N_4643);
and U5267 (N_5267,N_4443,N_4088);
or U5268 (N_5268,N_4102,N_4653);
nor U5269 (N_5269,N_4615,N_4329);
nand U5270 (N_5270,N_4554,N_4046);
and U5271 (N_5271,N_4038,N_4433);
xnor U5272 (N_5272,N_4566,N_4399);
and U5273 (N_5273,N_4097,N_4154);
and U5274 (N_5274,N_4019,N_4116);
or U5275 (N_5275,N_4504,N_4073);
nand U5276 (N_5276,N_4425,N_4493);
or U5277 (N_5277,N_4239,N_4477);
and U5278 (N_5278,N_4717,N_4787);
xnor U5279 (N_5279,N_4765,N_4635);
nor U5280 (N_5280,N_4590,N_4621);
xnor U5281 (N_5281,N_4171,N_4089);
or U5282 (N_5282,N_4230,N_4356);
nand U5283 (N_5283,N_4541,N_4356);
or U5284 (N_5284,N_4249,N_4651);
nor U5285 (N_5285,N_4303,N_4170);
nor U5286 (N_5286,N_4351,N_4639);
nor U5287 (N_5287,N_4061,N_4242);
or U5288 (N_5288,N_4617,N_4645);
and U5289 (N_5289,N_4594,N_4489);
nand U5290 (N_5290,N_4058,N_4323);
nor U5291 (N_5291,N_4027,N_4279);
nand U5292 (N_5292,N_4266,N_4667);
nand U5293 (N_5293,N_4226,N_4724);
nand U5294 (N_5294,N_4646,N_4648);
or U5295 (N_5295,N_4412,N_4464);
and U5296 (N_5296,N_4659,N_4011);
xnor U5297 (N_5297,N_4393,N_4476);
or U5298 (N_5298,N_4431,N_4662);
nor U5299 (N_5299,N_4595,N_4002);
and U5300 (N_5300,N_4191,N_4627);
and U5301 (N_5301,N_4556,N_4521);
or U5302 (N_5302,N_4401,N_4455);
nand U5303 (N_5303,N_4100,N_4002);
or U5304 (N_5304,N_4602,N_4478);
nand U5305 (N_5305,N_4152,N_4444);
or U5306 (N_5306,N_4086,N_4256);
or U5307 (N_5307,N_4469,N_4544);
xor U5308 (N_5308,N_4745,N_4393);
or U5309 (N_5309,N_4191,N_4571);
xor U5310 (N_5310,N_4343,N_4125);
nand U5311 (N_5311,N_4734,N_4031);
and U5312 (N_5312,N_4429,N_4319);
xnor U5313 (N_5313,N_4187,N_4054);
nor U5314 (N_5314,N_4414,N_4216);
nor U5315 (N_5315,N_4152,N_4635);
nor U5316 (N_5316,N_4170,N_4621);
xnor U5317 (N_5317,N_4362,N_4395);
or U5318 (N_5318,N_4618,N_4724);
nand U5319 (N_5319,N_4048,N_4391);
nor U5320 (N_5320,N_4672,N_4610);
or U5321 (N_5321,N_4396,N_4674);
or U5322 (N_5322,N_4774,N_4671);
or U5323 (N_5323,N_4786,N_4383);
xnor U5324 (N_5324,N_4631,N_4691);
xnor U5325 (N_5325,N_4481,N_4778);
nand U5326 (N_5326,N_4252,N_4061);
nand U5327 (N_5327,N_4744,N_4544);
or U5328 (N_5328,N_4316,N_4177);
or U5329 (N_5329,N_4648,N_4790);
nor U5330 (N_5330,N_4302,N_4048);
and U5331 (N_5331,N_4605,N_4115);
nor U5332 (N_5332,N_4515,N_4103);
xnor U5333 (N_5333,N_4785,N_4457);
and U5334 (N_5334,N_4674,N_4407);
xor U5335 (N_5335,N_4395,N_4297);
nor U5336 (N_5336,N_4690,N_4018);
nand U5337 (N_5337,N_4399,N_4616);
nand U5338 (N_5338,N_4354,N_4693);
xnor U5339 (N_5339,N_4342,N_4416);
xnor U5340 (N_5340,N_4265,N_4657);
nor U5341 (N_5341,N_4039,N_4507);
nand U5342 (N_5342,N_4008,N_4491);
or U5343 (N_5343,N_4553,N_4664);
nand U5344 (N_5344,N_4428,N_4341);
nor U5345 (N_5345,N_4032,N_4451);
and U5346 (N_5346,N_4058,N_4356);
or U5347 (N_5347,N_4734,N_4788);
nor U5348 (N_5348,N_4110,N_4045);
nand U5349 (N_5349,N_4162,N_4730);
nor U5350 (N_5350,N_4203,N_4320);
nor U5351 (N_5351,N_4330,N_4268);
and U5352 (N_5352,N_4108,N_4212);
xnor U5353 (N_5353,N_4356,N_4078);
and U5354 (N_5354,N_4245,N_4277);
xnor U5355 (N_5355,N_4257,N_4267);
nand U5356 (N_5356,N_4263,N_4789);
nor U5357 (N_5357,N_4656,N_4799);
or U5358 (N_5358,N_4776,N_4437);
nand U5359 (N_5359,N_4087,N_4442);
nor U5360 (N_5360,N_4478,N_4127);
xnor U5361 (N_5361,N_4076,N_4141);
nand U5362 (N_5362,N_4444,N_4198);
nor U5363 (N_5363,N_4620,N_4590);
xor U5364 (N_5364,N_4161,N_4465);
nand U5365 (N_5365,N_4530,N_4715);
nand U5366 (N_5366,N_4652,N_4428);
xor U5367 (N_5367,N_4681,N_4527);
and U5368 (N_5368,N_4792,N_4718);
xor U5369 (N_5369,N_4595,N_4779);
nor U5370 (N_5370,N_4690,N_4669);
nor U5371 (N_5371,N_4580,N_4611);
xnor U5372 (N_5372,N_4277,N_4455);
and U5373 (N_5373,N_4575,N_4030);
or U5374 (N_5374,N_4760,N_4636);
and U5375 (N_5375,N_4038,N_4317);
and U5376 (N_5376,N_4541,N_4226);
or U5377 (N_5377,N_4419,N_4722);
nor U5378 (N_5378,N_4498,N_4076);
nor U5379 (N_5379,N_4645,N_4265);
or U5380 (N_5380,N_4068,N_4217);
nor U5381 (N_5381,N_4310,N_4481);
or U5382 (N_5382,N_4262,N_4249);
nor U5383 (N_5383,N_4022,N_4333);
or U5384 (N_5384,N_4017,N_4617);
xor U5385 (N_5385,N_4533,N_4219);
or U5386 (N_5386,N_4236,N_4575);
nand U5387 (N_5387,N_4539,N_4701);
and U5388 (N_5388,N_4246,N_4437);
nor U5389 (N_5389,N_4562,N_4181);
and U5390 (N_5390,N_4329,N_4103);
nand U5391 (N_5391,N_4752,N_4316);
nand U5392 (N_5392,N_4795,N_4564);
xnor U5393 (N_5393,N_4327,N_4739);
xor U5394 (N_5394,N_4720,N_4483);
nand U5395 (N_5395,N_4148,N_4598);
or U5396 (N_5396,N_4076,N_4694);
xnor U5397 (N_5397,N_4388,N_4461);
nand U5398 (N_5398,N_4500,N_4041);
xor U5399 (N_5399,N_4481,N_4397);
nand U5400 (N_5400,N_4447,N_4473);
or U5401 (N_5401,N_4579,N_4004);
or U5402 (N_5402,N_4788,N_4165);
and U5403 (N_5403,N_4299,N_4727);
and U5404 (N_5404,N_4791,N_4677);
nand U5405 (N_5405,N_4443,N_4327);
and U5406 (N_5406,N_4664,N_4377);
nor U5407 (N_5407,N_4085,N_4122);
xnor U5408 (N_5408,N_4082,N_4370);
nand U5409 (N_5409,N_4289,N_4738);
or U5410 (N_5410,N_4498,N_4270);
nor U5411 (N_5411,N_4287,N_4118);
xnor U5412 (N_5412,N_4445,N_4318);
nor U5413 (N_5413,N_4270,N_4395);
or U5414 (N_5414,N_4225,N_4243);
nor U5415 (N_5415,N_4607,N_4441);
xnor U5416 (N_5416,N_4437,N_4658);
nor U5417 (N_5417,N_4235,N_4472);
xnor U5418 (N_5418,N_4097,N_4021);
or U5419 (N_5419,N_4413,N_4262);
xnor U5420 (N_5420,N_4073,N_4524);
or U5421 (N_5421,N_4171,N_4326);
and U5422 (N_5422,N_4148,N_4039);
nand U5423 (N_5423,N_4074,N_4010);
xnor U5424 (N_5424,N_4101,N_4364);
or U5425 (N_5425,N_4144,N_4291);
nand U5426 (N_5426,N_4470,N_4408);
nand U5427 (N_5427,N_4447,N_4386);
nand U5428 (N_5428,N_4726,N_4010);
nor U5429 (N_5429,N_4211,N_4790);
xnor U5430 (N_5430,N_4776,N_4675);
and U5431 (N_5431,N_4443,N_4441);
nand U5432 (N_5432,N_4389,N_4624);
xor U5433 (N_5433,N_4180,N_4026);
nor U5434 (N_5434,N_4456,N_4679);
nand U5435 (N_5435,N_4729,N_4579);
xnor U5436 (N_5436,N_4332,N_4145);
nand U5437 (N_5437,N_4490,N_4668);
or U5438 (N_5438,N_4579,N_4710);
and U5439 (N_5439,N_4145,N_4582);
nand U5440 (N_5440,N_4684,N_4739);
and U5441 (N_5441,N_4788,N_4577);
nand U5442 (N_5442,N_4335,N_4263);
xnor U5443 (N_5443,N_4442,N_4004);
nand U5444 (N_5444,N_4673,N_4449);
nand U5445 (N_5445,N_4594,N_4675);
nor U5446 (N_5446,N_4440,N_4005);
or U5447 (N_5447,N_4370,N_4142);
nor U5448 (N_5448,N_4384,N_4379);
or U5449 (N_5449,N_4771,N_4081);
nor U5450 (N_5450,N_4444,N_4005);
and U5451 (N_5451,N_4046,N_4686);
or U5452 (N_5452,N_4654,N_4581);
nor U5453 (N_5453,N_4493,N_4455);
or U5454 (N_5454,N_4280,N_4267);
nand U5455 (N_5455,N_4164,N_4795);
or U5456 (N_5456,N_4753,N_4324);
nor U5457 (N_5457,N_4669,N_4322);
xor U5458 (N_5458,N_4348,N_4656);
or U5459 (N_5459,N_4590,N_4044);
nand U5460 (N_5460,N_4689,N_4548);
xnor U5461 (N_5461,N_4107,N_4364);
or U5462 (N_5462,N_4639,N_4254);
nand U5463 (N_5463,N_4481,N_4176);
nand U5464 (N_5464,N_4615,N_4767);
and U5465 (N_5465,N_4656,N_4772);
nand U5466 (N_5466,N_4336,N_4501);
nor U5467 (N_5467,N_4708,N_4206);
xor U5468 (N_5468,N_4387,N_4115);
or U5469 (N_5469,N_4675,N_4172);
and U5470 (N_5470,N_4556,N_4382);
xor U5471 (N_5471,N_4548,N_4791);
or U5472 (N_5472,N_4204,N_4503);
nor U5473 (N_5473,N_4628,N_4339);
nand U5474 (N_5474,N_4693,N_4279);
or U5475 (N_5475,N_4304,N_4135);
nand U5476 (N_5476,N_4431,N_4282);
or U5477 (N_5477,N_4583,N_4573);
nand U5478 (N_5478,N_4247,N_4391);
or U5479 (N_5479,N_4397,N_4337);
or U5480 (N_5480,N_4422,N_4176);
nor U5481 (N_5481,N_4334,N_4742);
nand U5482 (N_5482,N_4325,N_4249);
or U5483 (N_5483,N_4510,N_4137);
and U5484 (N_5484,N_4605,N_4119);
nor U5485 (N_5485,N_4166,N_4776);
xnor U5486 (N_5486,N_4050,N_4448);
xor U5487 (N_5487,N_4613,N_4435);
or U5488 (N_5488,N_4569,N_4254);
or U5489 (N_5489,N_4014,N_4786);
nor U5490 (N_5490,N_4761,N_4425);
or U5491 (N_5491,N_4144,N_4495);
or U5492 (N_5492,N_4123,N_4240);
xnor U5493 (N_5493,N_4212,N_4626);
or U5494 (N_5494,N_4562,N_4223);
or U5495 (N_5495,N_4468,N_4482);
or U5496 (N_5496,N_4532,N_4780);
xnor U5497 (N_5497,N_4584,N_4401);
nand U5498 (N_5498,N_4575,N_4451);
or U5499 (N_5499,N_4080,N_4714);
and U5500 (N_5500,N_4573,N_4687);
or U5501 (N_5501,N_4398,N_4683);
xnor U5502 (N_5502,N_4003,N_4469);
nand U5503 (N_5503,N_4057,N_4382);
xor U5504 (N_5504,N_4113,N_4492);
nand U5505 (N_5505,N_4150,N_4487);
nand U5506 (N_5506,N_4072,N_4295);
or U5507 (N_5507,N_4362,N_4699);
and U5508 (N_5508,N_4479,N_4601);
nand U5509 (N_5509,N_4230,N_4386);
and U5510 (N_5510,N_4140,N_4261);
nor U5511 (N_5511,N_4621,N_4757);
and U5512 (N_5512,N_4463,N_4668);
or U5513 (N_5513,N_4131,N_4282);
and U5514 (N_5514,N_4311,N_4623);
or U5515 (N_5515,N_4356,N_4223);
nor U5516 (N_5516,N_4258,N_4238);
nand U5517 (N_5517,N_4279,N_4445);
xor U5518 (N_5518,N_4706,N_4670);
nor U5519 (N_5519,N_4706,N_4198);
nand U5520 (N_5520,N_4374,N_4467);
nand U5521 (N_5521,N_4225,N_4183);
or U5522 (N_5522,N_4683,N_4562);
nand U5523 (N_5523,N_4734,N_4638);
xor U5524 (N_5524,N_4258,N_4347);
nand U5525 (N_5525,N_4187,N_4051);
nand U5526 (N_5526,N_4537,N_4284);
nor U5527 (N_5527,N_4308,N_4617);
nand U5528 (N_5528,N_4549,N_4171);
or U5529 (N_5529,N_4526,N_4543);
and U5530 (N_5530,N_4590,N_4669);
xnor U5531 (N_5531,N_4026,N_4502);
nand U5532 (N_5532,N_4601,N_4034);
nand U5533 (N_5533,N_4506,N_4070);
nor U5534 (N_5534,N_4109,N_4307);
xor U5535 (N_5535,N_4055,N_4406);
or U5536 (N_5536,N_4088,N_4699);
xor U5537 (N_5537,N_4434,N_4482);
and U5538 (N_5538,N_4547,N_4668);
and U5539 (N_5539,N_4143,N_4136);
nand U5540 (N_5540,N_4609,N_4787);
xnor U5541 (N_5541,N_4413,N_4088);
and U5542 (N_5542,N_4739,N_4397);
nand U5543 (N_5543,N_4177,N_4042);
xnor U5544 (N_5544,N_4007,N_4582);
or U5545 (N_5545,N_4225,N_4184);
or U5546 (N_5546,N_4132,N_4237);
nand U5547 (N_5547,N_4116,N_4247);
and U5548 (N_5548,N_4495,N_4137);
xor U5549 (N_5549,N_4404,N_4282);
xor U5550 (N_5550,N_4733,N_4105);
nor U5551 (N_5551,N_4701,N_4389);
xnor U5552 (N_5552,N_4515,N_4586);
nor U5553 (N_5553,N_4509,N_4544);
xor U5554 (N_5554,N_4253,N_4465);
nor U5555 (N_5555,N_4212,N_4642);
xnor U5556 (N_5556,N_4434,N_4005);
xor U5557 (N_5557,N_4470,N_4637);
nor U5558 (N_5558,N_4552,N_4532);
nor U5559 (N_5559,N_4527,N_4224);
and U5560 (N_5560,N_4259,N_4573);
xnor U5561 (N_5561,N_4629,N_4502);
or U5562 (N_5562,N_4618,N_4435);
and U5563 (N_5563,N_4773,N_4172);
nor U5564 (N_5564,N_4663,N_4053);
xor U5565 (N_5565,N_4295,N_4167);
or U5566 (N_5566,N_4568,N_4581);
and U5567 (N_5567,N_4405,N_4008);
nand U5568 (N_5568,N_4499,N_4582);
nor U5569 (N_5569,N_4107,N_4020);
and U5570 (N_5570,N_4535,N_4349);
and U5571 (N_5571,N_4385,N_4376);
or U5572 (N_5572,N_4172,N_4684);
nand U5573 (N_5573,N_4771,N_4198);
and U5574 (N_5574,N_4116,N_4647);
or U5575 (N_5575,N_4357,N_4052);
and U5576 (N_5576,N_4603,N_4438);
and U5577 (N_5577,N_4181,N_4045);
and U5578 (N_5578,N_4529,N_4017);
and U5579 (N_5579,N_4197,N_4753);
and U5580 (N_5580,N_4188,N_4687);
nand U5581 (N_5581,N_4683,N_4627);
xnor U5582 (N_5582,N_4735,N_4232);
nand U5583 (N_5583,N_4133,N_4120);
nand U5584 (N_5584,N_4453,N_4175);
or U5585 (N_5585,N_4447,N_4783);
and U5586 (N_5586,N_4054,N_4170);
nor U5587 (N_5587,N_4386,N_4166);
and U5588 (N_5588,N_4317,N_4000);
nor U5589 (N_5589,N_4242,N_4345);
xor U5590 (N_5590,N_4716,N_4661);
nand U5591 (N_5591,N_4179,N_4751);
or U5592 (N_5592,N_4133,N_4334);
nor U5593 (N_5593,N_4087,N_4354);
nor U5594 (N_5594,N_4176,N_4780);
nor U5595 (N_5595,N_4393,N_4150);
or U5596 (N_5596,N_4398,N_4755);
nor U5597 (N_5597,N_4533,N_4152);
nor U5598 (N_5598,N_4548,N_4460);
and U5599 (N_5599,N_4516,N_4144);
nand U5600 (N_5600,N_4849,N_5408);
nor U5601 (N_5601,N_5098,N_4936);
nor U5602 (N_5602,N_5120,N_4812);
xnor U5603 (N_5603,N_4894,N_4945);
and U5604 (N_5604,N_5497,N_4911);
and U5605 (N_5605,N_4922,N_5506);
and U5606 (N_5606,N_4895,N_5326);
xor U5607 (N_5607,N_5006,N_4928);
and U5608 (N_5608,N_5243,N_4829);
xor U5609 (N_5609,N_5110,N_5448);
nand U5610 (N_5610,N_5552,N_4968);
nand U5611 (N_5611,N_5030,N_4824);
nor U5612 (N_5612,N_4846,N_5165);
nand U5613 (N_5613,N_5079,N_5330);
or U5614 (N_5614,N_5474,N_4946);
xnor U5615 (N_5615,N_5286,N_5278);
and U5616 (N_5616,N_4979,N_5238);
nor U5617 (N_5617,N_5227,N_5137);
xor U5618 (N_5618,N_5477,N_5437);
and U5619 (N_5619,N_5240,N_5595);
and U5620 (N_5620,N_5528,N_4943);
xnor U5621 (N_5621,N_5212,N_5094);
xnor U5622 (N_5622,N_4863,N_4896);
xor U5623 (N_5623,N_4834,N_5460);
xnor U5624 (N_5624,N_4951,N_4926);
or U5625 (N_5625,N_5185,N_4980);
nor U5626 (N_5626,N_4913,N_5307);
nand U5627 (N_5627,N_5572,N_5491);
or U5628 (N_5628,N_4978,N_4967);
or U5629 (N_5629,N_5438,N_4817);
or U5630 (N_5630,N_4907,N_5095);
nor U5631 (N_5631,N_4814,N_5260);
or U5632 (N_5632,N_5369,N_5266);
nor U5633 (N_5633,N_5591,N_5256);
or U5634 (N_5634,N_4971,N_5249);
and U5635 (N_5635,N_5596,N_5075);
nand U5636 (N_5636,N_5464,N_5233);
nor U5637 (N_5637,N_5017,N_4827);
nand U5638 (N_5638,N_5034,N_4972);
nor U5639 (N_5639,N_5005,N_5194);
and U5640 (N_5640,N_4871,N_5329);
and U5641 (N_5641,N_5028,N_5139);
xnor U5642 (N_5642,N_4995,N_5411);
nor U5643 (N_5643,N_5415,N_4805);
and U5644 (N_5644,N_5259,N_4800);
and U5645 (N_5645,N_5308,N_5353);
nand U5646 (N_5646,N_4937,N_5085);
nand U5647 (N_5647,N_5090,N_5401);
nand U5648 (N_5648,N_4899,N_5253);
nor U5649 (N_5649,N_5068,N_5056);
and U5650 (N_5650,N_5398,N_4906);
or U5651 (N_5651,N_4981,N_5053);
and U5652 (N_5652,N_5523,N_5208);
nand U5653 (N_5653,N_5275,N_5323);
nor U5654 (N_5654,N_5502,N_5381);
xnor U5655 (N_5655,N_4813,N_5407);
nand U5656 (N_5656,N_4925,N_5132);
nor U5657 (N_5657,N_4873,N_5232);
nor U5658 (N_5658,N_5190,N_5347);
or U5659 (N_5659,N_5453,N_5380);
and U5660 (N_5660,N_4898,N_5403);
nor U5661 (N_5661,N_4857,N_5527);
xor U5662 (N_5662,N_5131,N_5024);
nand U5663 (N_5663,N_5004,N_4944);
nand U5664 (N_5664,N_5057,N_5443);
and U5665 (N_5665,N_4958,N_4869);
nand U5666 (N_5666,N_5333,N_5588);
and U5667 (N_5667,N_4858,N_5292);
nand U5668 (N_5668,N_4825,N_5385);
xor U5669 (N_5669,N_4885,N_5488);
or U5670 (N_5670,N_5417,N_5136);
nand U5671 (N_5671,N_5200,N_4961);
and U5672 (N_5672,N_5064,N_5317);
xnor U5673 (N_5673,N_4986,N_5039);
xor U5674 (N_5674,N_5164,N_5166);
or U5675 (N_5675,N_4838,N_4847);
or U5676 (N_5676,N_5390,N_5172);
or U5677 (N_5677,N_5069,N_5533);
nand U5678 (N_5678,N_5519,N_5283);
xnor U5679 (N_5679,N_5360,N_5269);
nor U5680 (N_5680,N_5117,N_5092);
nand U5681 (N_5681,N_5456,N_4920);
nor U5682 (N_5682,N_5322,N_5141);
nand U5683 (N_5683,N_5044,N_5300);
or U5684 (N_5684,N_4973,N_5454);
xor U5685 (N_5685,N_4924,N_5134);
nor U5686 (N_5686,N_5178,N_5433);
nand U5687 (N_5687,N_5224,N_5237);
xnor U5688 (N_5688,N_5346,N_4853);
nand U5689 (N_5689,N_5100,N_5078);
or U5690 (N_5690,N_5109,N_4884);
nand U5691 (N_5691,N_5305,N_5501);
or U5692 (N_5692,N_4888,N_5220);
nand U5693 (N_5693,N_5143,N_5507);
or U5694 (N_5694,N_5222,N_4855);
and U5695 (N_5695,N_4820,N_4864);
xnor U5696 (N_5696,N_5435,N_4993);
nor U5697 (N_5697,N_5434,N_4874);
nor U5698 (N_5698,N_5549,N_5146);
and U5699 (N_5699,N_5402,N_5421);
and U5700 (N_5700,N_4878,N_5129);
and U5701 (N_5701,N_5036,N_5587);
nor U5702 (N_5702,N_5127,N_5444);
xnor U5703 (N_5703,N_5344,N_5512);
and U5704 (N_5704,N_4938,N_5458);
or U5705 (N_5705,N_5379,N_5348);
and U5706 (N_5706,N_5043,N_5149);
and U5707 (N_5707,N_5001,N_5545);
nor U5708 (N_5708,N_5280,N_5350);
and U5709 (N_5709,N_5555,N_5213);
xnor U5710 (N_5710,N_4999,N_5067);
and U5711 (N_5711,N_5032,N_5331);
nand U5712 (N_5712,N_5535,N_5008);
and U5713 (N_5713,N_5514,N_5257);
nor U5714 (N_5714,N_4970,N_5550);
nand U5715 (N_5715,N_5375,N_5383);
and U5716 (N_5716,N_5084,N_5291);
or U5717 (N_5717,N_5371,N_4890);
or U5718 (N_5718,N_5176,N_5461);
nand U5719 (N_5719,N_5066,N_4832);
and U5720 (N_5720,N_5060,N_5562);
nor U5721 (N_5721,N_4856,N_5026);
nor U5722 (N_5722,N_5374,N_5569);
and U5723 (N_5723,N_5116,N_5387);
nand U5724 (N_5724,N_5288,N_5503);
or U5725 (N_5725,N_5018,N_4991);
and U5726 (N_5726,N_4974,N_4892);
nand U5727 (N_5727,N_5386,N_5103);
and U5728 (N_5728,N_5570,N_5351);
nor U5729 (N_5729,N_5123,N_4960);
or U5730 (N_5730,N_5363,N_4949);
nand U5731 (N_5731,N_5585,N_5155);
nor U5732 (N_5732,N_4964,N_5590);
and U5733 (N_5733,N_4982,N_4833);
nand U5734 (N_5734,N_4839,N_4891);
and U5735 (N_5735,N_5483,N_5184);
xor U5736 (N_5736,N_5599,N_5097);
nand U5737 (N_5737,N_5573,N_5239);
xor U5738 (N_5738,N_5541,N_5251);
and U5739 (N_5739,N_5513,N_4917);
nand U5740 (N_5740,N_5175,N_5193);
xor U5741 (N_5741,N_5153,N_4963);
nor U5742 (N_5742,N_5357,N_5538);
and U5743 (N_5743,N_4870,N_5158);
and U5744 (N_5744,N_5582,N_5508);
nand U5745 (N_5745,N_5478,N_5135);
xor U5746 (N_5746,N_4996,N_5581);
nand U5747 (N_5747,N_5526,N_5480);
and U5748 (N_5748,N_5180,N_5159);
and U5749 (N_5749,N_5367,N_5225);
nand U5750 (N_5750,N_5575,N_4952);
and U5751 (N_5751,N_5261,N_5309);
and U5752 (N_5752,N_5577,N_5274);
and U5753 (N_5753,N_5424,N_5107);
nand U5754 (N_5754,N_5148,N_5082);
and U5755 (N_5755,N_5061,N_5365);
nor U5756 (N_5756,N_5262,N_5485);
or U5757 (N_5757,N_4914,N_5228);
and U5758 (N_5758,N_4923,N_4865);
xor U5759 (N_5759,N_4909,N_5567);
nand U5760 (N_5760,N_5049,N_4860);
xor U5761 (N_5761,N_5258,N_5336);
or U5762 (N_5762,N_5469,N_5396);
and U5763 (N_5763,N_5169,N_5389);
nor U5764 (N_5764,N_5204,N_5510);
nand U5765 (N_5765,N_5203,N_4830);
xnor U5766 (N_5766,N_4897,N_5349);
xnor U5767 (N_5767,N_5284,N_5509);
xnor U5768 (N_5768,N_5548,N_5201);
or U5769 (N_5769,N_4984,N_5393);
nand U5770 (N_5770,N_5406,N_5167);
nor U5771 (N_5771,N_5559,N_4910);
or U5772 (N_5772,N_5031,N_5161);
and U5773 (N_5773,N_5242,N_5042);
xnor U5774 (N_5774,N_5229,N_4994);
or U5775 (N_5775,N_5188,N_5250);
xnor U5776 (N_5776,N_5293,N_5035);
and U5777 (N_5777,N_5128,N_5086);
or U5778 (N_5778,N_5440,N_5499);
or U5779 (N_5779,N_5231,N_5553);
nor U5780 (N_5780,N_5270,N_5295);
or U5781 (N_5781,N_4818,N_4831);
nand U5782 (N_5782,N_5029,N_4880);
xnor U5783 (N_5783,N_5170,N_5163);
and U5784 (N_5784,N_5314,N_5074);
xnor U5785 (N_5785,N_5486,N_5122);
and U5786 (N_5786,N_5471,N_5530);
or U5787 (N_5787,N_5126,N_5304);
or U5788 (N_5788,N_5400,N_4806);
or U5789 (N_5789,N_5459,N_5140);
xnor U5790 (N_5790,N_4802,N_5397);
and U5791 (N_5791,N_5101,N_5425);
xnor U5792 (N_5792,N_5558,N_5455);
or U5793 (N_5793,N_5327,N_5119);
or U5794 (N_5794,N_5306,N_5505);
and U5795 (N_5795,N_5422,N_5112);
nand U5796 (N_5796,N_5209,N_4861);
and U5797 (N_5797,N_5125,N_5152);
nor U5798 (N_5798,N_5298,N_5010);
nor U5799 (N_5799,N_5529,N_5426);
nand U5800 (N_5800,N_5554,N_5248);
xor U5801 (N_5801,N_5564,N_5160);
and U5802 (N_5802,N_4959,N_5038);
nand U5803 (N_5803,N_5279,N_4953);
and U5804 (N_5804,N_5334,N_5054);
xor U5805 (N_5805,N_5059,N_4866);
nand U5806 (N_5806,N_5187,N_5504);
nor U5807 (N_5807,N_5579,N_5568);
nand U5808 (N_5808,N_5083,N_5009);
xor U5809 (N_5809,N_5446,N_5332);
and U5810 (N_5810,N_5593,N_5565);
nor U5811 (N_5811,N_4810,N_5432);
and U5812 (N_5812,N_4886,N_4988);
or U5813 (N_5813,N_4900,N_5356);
xor U5814 (N_5814,N_4989,N_4941);
nand U5815 (N_5815,N_5003,N_5431);
and U5816 (N_5816,N_4876,N_5002);
nand U5817 (N_5817,N_5518,N_4842);
or U5818 (N_5818,N_4882,N_5156);
nor U5819 (N_5819,N_5179,N_5532);
nor U5820 (N_5820,N_5484,N_4841);
nor U5821 (N_5821,N_5047,N_5466);
nor U5822 (N_5822,N_5359,N_5487);
nand U5823 (N_5823,N_5445,N_5021);
or U5824 (N_5824,N_4826,N_4992);
and U5825 (N_5825,N_5252,N_4815);
xor U5826 (N_5826,N_5055,N_5181);
nor U5827 (N_5827,N_5162,N_5467);
nand U5828 (N_5828,N_5521,N_5320);
xnor U5829 (N_5829,N_5276,N_5087);
nand U5830 (N_5830,N_5493,N_5543);
nand U5831 (N_5831,N_4836,N_5197);
xnor U5832 (N_5832,N_4843,N_5576);
and U5833 (N_5833,N_5272,N_5404);
and U5834 (N_5834,N_5151,N_5303);
or U5835 (N_5835,N_4908,N_5150);
and U5836 (N_5836,N_5255,N_5451);
and U5837 (N_5837,N_5364,N_5277);
nand U5838 (N_5838,N_4930,N_5247);
xnor U5839 (N_5839,N_5168,N_5366);
nor U5840 (N_5840,N_5007,N_5073);
xor U5841 (N_5841,N_5391,N_5267);
or U5842 (N_5842,N_5537,N_5598);
and U5843 (N_5843,N_5378,N_5210);
nor U5844 (N_5844,N_5594,N_5016);
and U5845 (N_5845,N_5195,N_5586);
nor U5846 (N_5846,N_5318,N_5345);
nor U5847 (N_5847,N_5312,N_5539);
and U5848 (N_5848,N_5515,N_5102);
or U5849 (N_5849,N_5273,N_4819);
and U5850 (N_5850,N_5234,N_5093);
nand U5851 (N_5851,N_5045,N_5462);
and U5852 (N_5852,N_5089,N_5072);
xor U5853 (N_5853,N_5392,N_4854);
nand U5854 (N_5854,N_5281,N_5423);
nor U5855 (N_5855,N_4845,N_5511);
nor U5856 (N_5856,N_5362,N_5547);
nor U5857 (N_5857,N_5182,N_4921);
and U5858 (N_5858,N_5215,N_5321);
or U5859 (N_5859,N_5409,N_5335);
xnor U5860 (N_5860,N_5382,N_5070);
xnor U5861 (N_5861,N_4852,N_5520);
xor U5862 (N_5862,N_5081,N_4867);
nand U5863 (N_5863,N_4942,N_4823);
nor U5864 (N_5864,N_5235,N_4940);
and U5865 (N_5865,N_4948,N_4889);
nand U5866 (N_5866,N_5157,N_4933);
nor U5867 (N_5867,N_5196,N_5427);
and U5868 (N_5868,N_5524,N_5589);
nand U5869 (N_5869,N_5566,N_5463);
nand U5870 (N_5870,N_4932,N_4850);
and U5871 (N_5871,N_4879,N_5027);
nand U5872 (N_5872,N_4955,N_4837);
and U5873 (N_5873,N_5439,N_5492);
nand U5874 (N_5874,N_5370,N_5494);
nand U5875 (N_5875,N_5338,N_5557);
and U5876 (N_5876,N_4828,N_5241);
xnor U5877 (N_5877,N_5145,N_5022);
nor U5878 (N_5878,N_4962,N_5144);
xnor U5879 (N_5879,N_5516,N_5058);
nand U5880 (N_5880,N_4862,N_5405);
xnor U5881 (N_5881,N_4915,N_5000);
nand U5882 (N_5882,N_5372,N_4809);
or U5883 (N_5883,N_5263,N_5413);
xnor U5884 (N_5884,N_5419,N_5546);
and U5885 (N_5885,N_5174,N_5498);
nand U5886 (N_5886,N_5302,N_5012);
or U5887 (N_5887,N_5342,N_4903);
nor U5888 (N_5888,N_5219,N_5481);
xor U5889 (N_5889,N_4905,N_5449);
nor U5890 (N_5890,N_5050,N_5388);
nand U5891 (N_5891,N_4803,N_5358);
and U5892 (N_5892,N_5289,N_5341);
or U5893 (N_5893,N_5414,N_5536);
nor U5894 (N_5894,N_4821,N_5465);
or U5895 (N_5895,N_5418,N_5230);
nand U5896 (N_5896,N_5121,N_5325);
or U5897 (N_5897,N_4840,N_5416);
nand U5898 (N_5898,N_5412,N_5096);
nand U5899 (N_5899,N_5099,N_5221);
xnor U5900 (N_5900,N_5297,N_5063);
and U5901 (N_5901,N_5337,N_4877);
nor U5902 (N_5902,N_5118,N_4902);
or U5903 (N_5903,N_5368,N_5216);
and U5904 (N_5904,N_4976,N_4918);
or U5905 (N_5905,N_5091,N_5597);
xnor U5906 (N_5906,N_5246,N_5111);
nand U5907 (N_5907,N_4893,N_5352);
or U5908 (N_5908,N_5282,N_5019);
nand U5909 (N_5909,N_5113,N_5339);
nand U5910 (N_5910,N_5583,N_5355);
nand U5911 (N_5911,N_4851,N_5025);
nand U5912 (N_5912,N_5399,N_5108);
nor U5913 (N_5913,N_4848,N_5065);
and U5914 (N_5914,N_4887,N_5052);
and U5915 (N_5915,N_5154,N_5441);
nor U5916 (N_5916,N_5580,N_5534);
or U5917 (N_5917,N_5207,N_4916);
xnor U5918 (N_5918,N_4919,N_5592);
xor U5919 (N_5919,N_5561,N_5015);
nand U5920 (N_5920,N_5033,N_5476);
nor U5921 (N_5921,N_4977,N_5522);
and U5922 (N_5922,N_5430,N_4947);
xnor U5923 (N_5923,N_5011,N_4816);
or U5924 (N_5924,N_5315,N_5147);
xor U5925 (N_5925,N_4801,N_4975);
xor U5926 (N_5926,N_5214,N_5489);
nand U5927 (N_5927,N_4883,N_5177);
or U5928 (N_5928,N_4956,N_4912);
xor U5929 (N_5929,N_5531,N_5077);
and U5930 (N_5930,N_5447,N_5354);
or U5931 (N_5931,N_5473,N_5479);
and U5932 (N_5932,N_5490,N_4957);
and U5933 (N_5933,N_5205,N_5544);
or U5934 (N_5934,N_4875,N_5223);
nand U5935 (N_5935,N_4904,N_4935);
xor U5936 (N_5936,N_5496,N_4807);
or U5937 (N_5937,N_4901,N_5236);
or U5938 (N_5938,N_5254,N_5517);
xor U5939 (N_5939,N_5563,N_5429);
xnor U5940 (N_5940,N_5500,N_4804);
or U5941 (N_5941,N_4969,N_5574);
nand U5942 (N_5942,N_5340,N_5245);
nand U5943 (N_5943,N_5062,N_5189);
nand U5944 (N_5944,N_4872,N_5217);
and U5945 (N_5945,N_5023,N_5173);
xor U5946 (N_5946,N_5076,N_5301);
xnor U5947 (N_5947,N_5271,N_5183);
xnor U5948 (N_5948,N_5287,N_4939);
and U5949 (N_5949,N_4950,N_5395);
nor U5950 (N_5950,N_5124,N_5560);
xnor U5951 (N_5951,N_5048,N_5051);
or U5952 (N_5952,N_5442,N_5265);
and U5953 (N_5953,N_5268,N_5376);
nand U5954 (N_5954,N_4931,N_5202);
xor U5955 (N_5955,N_5285,N_5578);
and U5956 (N_5956,N_5296,N_5115);
xor U5957 (N_5957,N_4934,N_5218);
nor U5958 (N_5958,N_5046,N_5482);
xnor U5959 (N_5959,N_5294,N_5104);
and U5960 (N_5960,N_5014,N_5244);
nand U5961 (N_5961,N_5071,N_5114);
nor U5962 (N_5962,N_4965,N_5468);
xor U5963 (N_5963,N_5428,N_5206);
nand U5964 (N_5964,N_4987,N_5584);
xor U5965 (N_5965,N_5457,N_4990);
or U5966 (N_5966,N_4822,N_4927);
or U5967 (N_5967,N_4835,N_5525);
xor U5968 (N_5968,N_5343,N_5450);
and U5969 (N_5969,N_5470,N_5420);
nand U5970 (N_5970,N_5542,N_5186);
nor U5971 (N_5971,N_5199,N_5138);
or U5972 (N_5972,N_4929,N_5142);
or U5973 (N_5973,N_4998,N_4868);
nor U5974 (N_5974,N_5310,N_5130);
nor U5975 (N_5975,N_5299,N_5452);
or U5976 (N_5976,N_5041,N_5088);
and U5977 (N_5977,N_5556,N_5290);
nor U5978 (N_5978,N_5211,N_5226);
xnor U5979 (N_5979,N_5475,N_4985);
xnor U5980 (N_5980,N_5324,N_5316);
nor U5981 (N_5981,N_5410,N_5020);
and U5982 (N_5982,N_5080,N_4859);
nand U5983 (N_5983,N_5313,N_5133);
and U5984 (N_5984,N_4808,N_5373);
nand U5985 (N_5985,N_5105,N_5436);
nor U5986 (N_5986,N_5394,N_5551);
xor U5987 (N_5987,N_4983,N_5191);
xnor U5988 (N_5988,N_5106,N_5264);
nand U5989 (N_5989,N_5495,N_4997);
nor U5990 (N_5990,N_4966,N_5540);
xor U5991 (N_5991,N_5171,N_5328);
and U5992 (N_5992,N_5384,N_5319);
xor U5993 (N_5993,N_5472,N_5361);
and U5994 (N_5994,N_4844,N_5198);
and U5995 (N_5995,N_5040,N_5037);
xor U5996 (N_5996,N_5192,N_4954);
nand U5997 (N_5997,N_4811,N_5571);
and U5998 (N_5998,N_5311,N_4881);
xor U5999 (N_5999,N_5377,N_5013);
xor U6000 (N_6000,N_4938,N_4889);
and U6001 (N_6001,N_5335,N_4817);
and U6002 (N_6002,N_5431,N_5168);
and U6003 (N_6003,N_5392,N_5015);
nor U6004 (N_6004,N_5595,N_5202);
nor U6005 (N_6005,N_5232,N_4817);
xor U6006 (N_6006,N_5031,N_5003);
and U6007 (N_6007,N_5290,N_4826);
nor U6008 (N_6008,N_5499,N_5095);
nand U6009 (N_6009,N_5069,N_5106);
or U6010 (N_6010,N_4881,N_5477);
nor U6011 (N_6011,N_4842,N_5029);
or U6012 (N_6012,N_5084,N_4829);
xor U6013 (N_6013,N_4881,N_5068);
xor U6014 (N_6014,N_5392,N_4883);
and U6015 (N_6015,N_5007,N_4976);
nand U6016 (N_6016,N_5012,N_5388);
nor U6017 (N_6017,N_5187,N_5505);
nor U6018 (N_6018,N_5044,N_5442);
nor U6019 (N_6019,N_5178,N_4813);
nand U6020 (N_6020,N_5106,N_5380);
nor U6021 (N_6021,N_4897,N_5014);
or U6022 (N_6022,N_5238,N_5547);
nand U6023 (N_6023,N_5146,N_5376);
or U6024 (N_6024,N_4982,N_4959);
or U6025 (N_6025,N_5232,N_5044);
or U6026 (N_6026,N_5461,N_5464);
nor U6027 (N_6027,N_4870,N_5278);
xor U6028 (N_6028,N_5538,N_5396);
nor U6029 (N_6029,N_4956,N_5170);
nand U6030 (N_6030,N_5375,N_5288);
or U6031 (N_6031,N_5189,N_5103);
nor U6032 (N_6032,N_5463,N_5150);
or U6033 (N_6033,N_4998,N_5454);
or U6034 (N_6034,N_5580,N_5026);
nor U6035 (N_6035,N_5221,N_4954);
or U6036 (N_6036,N_5194,N_5097);
nor U6037 (N_6037,N_5377,N_4930);
xor U6038 (N_6038,N_5098,N_4893);
or U6039 (N_6039,N_4800,N_5147);
nor U6040 (N_6040,N_5161,N_5281);
nor U6041 (N_6041,N_4917,N_5522);
xnor U6042 (N_6042,N_5178,N_5188);
nor U6043 (N_6043,N_5465,N_4955);
nand U6044 (N_6044,N_5418,N_5400);
nor U6045 (N_6045,N_4958,N_5525);
xor U6046 (N_6046,N_5330,N_5580);
and U6047 (N_6047,N_5170,N_4958);
or U6048 (N_6048,N_4906,N_4976);
or U6049 (N_6049,N_5504,N_5528);
and U6050 (N_6050,N_5085,N_4950);
xor U6051 (N_6051,N_5568,N_5376);
xnor U6052 (N_6052,N_4942,N_5216);
xnor U6053 (N_6053,N_4809,N_5434);
or U6054 (N_6054,N_5225,N_5525);
or U6055 (N_6055,N_5550,N_5113);
xnor U6056 (N_6056,N_5001,N_5012);
or U6057 (N_6057,N_5136,N_5009);
or U6058 (N_6058,N_4984,N_5424);
xor U6059 (N_6059,N_4896,N_5389);
or U6060 (N_6060,N_5310,N_5074);
or U6061 (N_6061,N_4916,N_5474);
and U6062 (N_6062,N_5579,N_5205);
xnor U6063 (N_6063,N_5495,N_5255);
nand U6064 (N_6064,N_5038,N_5391);
nor U6065 (N_6065,N_5571,N_5088);
nor U6066 (N_6066,N_5490,N_5331);
xnor U6067 (N_6067,N_5334,N_5484);
nand U6068 (N_6068,N_5167,N_5061);
and U6069 (N_6069,N_5382,N_5366);
and U6070 (N_6070,N_4888,N_5269);
nor U6071 (N_6071,N_5128,N_5058);
nor U6072 (N_6072,N_5154,N_5096);
and U6073 (N_6073,N_5528,N_5205);
nor U6074 (N_6074,N_5174,N_4922);
or U6075 (N_6075,N_5587,N_5124);
nand U6076 (N_6076,N_5464,N_5323);
and U6077 (N_6077,N_5400,N_4903);
nand U6078 (N_6078,N_5478,N_5514);
or U6079 (N_6079,N_4851,N_5083);
or U6080 (N_6080,N_5575,N_5256);
nor U6081 (N_6081,N_5185,N_5198);
xnor U6082 (N_6082,N_5110,N_5513);
or U6083 (N_6083,N_5025,N_4912);
xnor U6084 (N_6084,N_4965,N_5004);
nand U6085 (N_6085,N_5000,N_5555);
nand U6086 (N_6086,N_5583,N_5076);
and U6087 (N_6087,N_5518,N_4865);
nor U6088 (N_6088,N_5352,N_5283);
nor U6089 (N_6089,N_5568,N_5267);
and U6090 (N_6090,N_4973,N_5200);
nor U6091 (N_6091,N_4812,N_5357);
nand U6092 (N_6092,N_4943,N_5153);
or U6093 (N_6093,N_5093,N_5210);
and U6094 (N_6094,N_5101,N_5292);
nor U6095 (N_6095,N_5188,N_5181);
nand U6096 (N_6096,N_5359,N_4824);
nand U6097 (N_6097,N_5085,N_5514);
or U6098 (N_6098,N_5346,N_5456);
xnor U6099 (N_6099,N_5402,N_5487);
or U6100 (N_6100,N_5534,N_5434);
and U6101 (N_6101,N_4837,N_5039);
and U6102 (N_6102,N_4933,N_5285);
nand U6103 (N_6103,N_5111,N_5544);
and U6104 (N_6104,N_5449,N_5188);
nand U6105 (N_6105,N_4846,N_5515);
nor U6106 (N_6106,N_5588,N_5164);
xnor U6107 (N_6107,N_4976,N_4915);
nand U6108 (N_6108,N_5399,N_5112);
or U6109 (N_6109,N_5302,N_5476);
or U6110 (N_6110,N_5246,N_5408);
xor U6111 (N_6111,N_5534,N_5293);
and U6112 (N_6112,N_5491,N_4938);
nand U6113 (N_6113,N_5191,N_5241);
xnor U6114 (N_6114,N_5222,N_5098);
xnor U6115 (N_6115,N_5575,N_4935);
nand U6116 (N_6116,N_5280,N_5299);
xnor U6117 (N_6117,N_5154,N_4977);
xnor U6118 (N_6118,N_4942,N_4934);
or U6119 (N_6119,N_5505,N_5590);
nand U6120 (N_6120,N_5009,N_5488);
nand U6121 (N_6121,N_5349,N_5406);
nor U6122 (N_6122,N_5240,N_5580);
nand U6123 (N_6123,N_5261,N_5274);
xnor U6124 (N_6124,N_5216,N_5045);
or U6125 (N_6125,N_4843,N_5282);
and U6126 (N_6126,N_5169,N_5326);
xnor U6127 (N_6127,N_4910,N_5487);
nor U6128 (N_6128,N_4986,N_5059);
and U6129 (N_6129,N_5131,N_5289);
xnor U6130 (N_6130,N_5346,N_5263);
nor U6131 (N_6131,N_5193,N_5413);
xnor U6132 (N_6132,N_5084,N_5158);
or U6133 (N_6133,N_5216,N_5416);
nor U6134 (N_6134,N_5179,N_5450);
and U6135 (N_6135,N_5453,N_5267);
nand U6136 (N_6136,N_5529,N_4970);
nor U6137 (N_6137,N_5055,N_5159);
nor U6138 (N_6138,N_5022,N_5201);
xnor U6139 (N_6139,N_5354,N_5198);
xnor U6140 (N_6140,N_5392,N_5084);
nand U6141 (N_6141,N_5211,N_5443);
and U6142 (N_6142,N_5509,N_5147);
xor U6143 (N_6143,N_5415,N_4982);
or U6144 (N_6144,N_5194,N_4876);
xor U6145 (N_6145,N_5444,N_4834);
nor U6146 (N_6146,N_5071,N_5268);
nor U6147 (N_6147,N_5587,N_5563);
or U6148 (N_6148,N_5006,N_5198);
or U6149 (N_6149,N_5257,N_4933);
and U6150 (N_6150,N_5461,N_5449);
and U6151 (N_6151,N_5246,N_5005);
nand U6152 (N_6152,N_5477,N_5562);
and U6153 (N_6153,N_4897,N_4957);
or U6154 (N_6154,N_4882,N_4933);
and U6155 (N_6155,N_5117,N_4940);
xnor U6156 (N_6156,N_4800,N_4939);
and U6157 (N_6157,N_5143,N_5062);
and U6158 (N_6158,N_5308,N_5115);
or U6159 (N_6159,N_5335,N_5338);
and U6160 (N_6160,N_5148,N_5010);
nand U6161 (N_6161,N_5157,N_5249);
or U6162 (N_6162,N_5145,N_4815);
or U6163 (N_6163,N_5345,N_5371);
xnor U6164 (N_6164,N_5072,N_5397);
nor U6165 (N_6165,N_5323,N_5116);
nor U6166 (N_6166,N_4983,N_5002);
or U6167 (N_6167,N_5155,N_5091);
nor U6168 (N_6168,N_5438,N_5365);
nor U6169 (N_6169,N_5067,N_5478);
xnor U6170 (N_6170,N_4801,N_4931);
xnor U6171 (N_6171,N_5445,N_4952);
nor U6172 (N_6172,N_5077,N_5512);
nor U6173 (N_6173,N_4841,N_5453);
nor U6174 (N_6174,N_5309,N_5300);
or U6175 (N_6175,N_5299,N_4856);
and U6176 (N_6176,N_5168,N_5344);
xor U6177 (N_6177,N_5378,N_5560);
nor U6178 (N_6178,N_5476,N_5465);
nor U6179 (N_6179,N_5117,N_5459);
nor U6180 (N_6180,N_5169,N_5480);
nor U6181 (N_6181,N_5567,N_5430);
nand U6182 (N_6182,N_5236,N_5303);
xor U6183 (N_6183,N_5520,N_5513);
xnor U6184 (N_6184,N_5175,N_4984);
nor U6185 (N_6185,N_5275,N_5142);
nand U6186 (N_6186,N_4821,N_5190);
nand U6187 (N_6187,N_5049,N_5257);
or U6188 (N_6188,N_5218,N_4829);
and U6189 (N_6189,N_5463,N_5160);
or U6190 (N_6190,N_5369,N_4800);
and U6191 (N_6191,N_4894,N_5377);
nor U6192 (N_6192,N_4904,N_5278);
and U6193 (N_6193,N_4839,N_5283);
or U6194 (N_6194,N_4896,N_4830);
nand U6195 (N_6195,N_5091,N_5027);
or U6196 (N_6196,N_5339,N_5252);
nor U6197 (N_6197,N_5483,N_5047);
and U6198 (N_6198,N_5317,N_5599);
or U6199 (N_6199,N_4846,N_5482);
xnor U6200 (N_6200,N_5497,N_5307);
nor U6201 (N_6201,N_4867,N_4848);
nand U6202 (N_6202,N_5193,N_4817);
xnor U6203 (N_6203,N_5536,N_5106);
or U6204 (N_6204,N_5272,N_5433);
nand U6205 (N_6205,N_4878,N_5181);
nand U6206 (N_6206,N_5099,N_5578);
xor U6207 (N_6207,N_4939,N_4859);
nor U6208 (N_6208,N_5429,N_5328);
and U6209 (N_6209,N_5589,N_5478);
nor U6210 (N_6210,N_5347,N_5460);
nor U6211 (N_6211,N_5029,N_5003);
and U6212 (N_6212,N_5035,N_5117);
or U6213 (N_6213,N_5415,N_4874);
xnor U6214 (N_6214,N_5530,N_5293);
and U6215 (N_6215,N_4944,N_5424);
and U6216 (N_6216,N_4831,N_5564);
or U6217 (N_6217,N_5489,N_5285);
nor U6218 (N_6218,N_5058,N_4830);
nand U6219 (N_6219,N_5193,N_4945);
or U6220 (N_6220,N_5147,N_5256);
or U6221 (N_6221,N_5527,N_5128);
and U6222 (N_6222,N_4906,N_5505);
nor U6223 (N_6223,N_5367,N_5288);
xnor U6224 (N_6224,N_5503,N_5046);
nand U6225 (N_6225,N_4842,N_4984);
nand U6226 (N_6226,N_5578,N_5592);
or U6227 (N_6227,N_4815,N_5516);
nor U6228 (N_6228,N_4872,N_5314);
or U6229 (N_6229,N_5451,N_4935);
nand U6230 (N_6230,N_5028,N_5505);
and U6231 (N_6231,N_5594,N_4933);
nor U6232 (N_6232,N_5115,N_4955);
nor U6233 (N_6233,N_5579,N_5068);
nand U6234 (N_6234,N_5035,N_5464);
or U6235 (N_6235,N_5347,N_4946);
nor U6236 (N_6236,N_5334,N_5394);
and U6237 (N_6237,N_4839,N_5389);
or U6238 (N_6238,N_4853,N_5130);
xor U6239 (N_6239,N_5157,N_4884);
and U6240 (N_6240,N_4942,N_5579);
xnor U6241 (N_6241,N_5331,N_5596);
xor U6242 (N_6242,N_4823,N_5519);
xnor U6243 (N_6243,N_4954,N_5224);
and U6244 (N_6244,N_5558,N_5008);
nand U6245 (N_6245,N_5067,N_5039);
xnor U6246 (N_6246,N_4980,N_5289);
or U6247 (N_6247,N_5260,N_5053);
xor U6248 (N_6248,N_5563,N_5072);
nand U6249 (N_6249,N_5568,N_5404);
or U6250 (N_6250,N_5557,N_5107);
or U6251 (N_6251,N_5028,N_5402);
xor U6252 (N_6252,N_5511,N_5361);
nor U6253 (N_6253,N_5101,N_4869);
or U6254 (N_6254,N_5357,N_5359);
or U6255 (N_6255,N_5491,N_5507);
or U6256 (N_6256,N_5584,N_5026);
or U6257 (N_6257,N_4920,N_5095);
nor U6258 (N_6258,N_5285,N_5016);
nor U6259 (N_6259,N_4967,N_5308);
xor U6260 (N_6260,N_5293,N_4857);
nand U6261 (N_6261,N_5303,N_5127);
nand U6262 (N_6262,N_4919,N_5417);
or U6263 (N_6263,N_4882,N_5256);
and U6264 (N_6264,N_5312,N_5225);
nand U6265 (N_6265,N_5126,N_5103);
and U6266 (N_6266,N_5371,N_5545);
xnor U6267 (N_6267,N_4823,N_4883);
or U6268 (N_6268,N_5037,N_5088);
nor U6269 (N_6269,N_4994,N_5433);
xor U6270 (N_6270,N_5597,N_5000);
xnor U6271 (N_6271,N_5567,N_5080);
and U6272 (N_6272,N_5563,N_4958);
nor U6273 (N_6273,N_5269,N_5304);
or U6274 (N_6274,N_5334,N_5521);
nor U6275 (N_6275,N_5001,N_5146);
xor U6276 (N_6276,N_4905,N_5289);
and U6277 (N_6277,N_5070,N_5554);
nor U6278 (N_6278,N_5548,N_5371);
or U6279 (N_6279,N_5184,N_5338);
xor U6280 (N_6280,N_5330,N_5150);
nor U6281 (N_6281,N_5158,N_5268);
nor U6282 (N_6282,N_4986,N_5386);
and U6283 (N_6283,N_5358,N_5049);
nand U6284 (N_6284,N_5549,N_4880);
nand U6285 (N_6285,N_5490,N_5188);
and U6286 (N_6286,N_5567,N_5435);
xnor U6287 (N_6287,N_5574,N_5503);
nor U6288 (N_6288,N_5271,N_5392);
nand U6289 (N_6289,N_5373,N_5211);
nor U6290 (N_6290,N_5100,N_4911);
nor U6291 (N_6291,N_5566,N_4802);
nand U6292 (N_6292,N_4912,N_5574);
and U6293 (N_6293,N_4850,N_5554);
or U6294 (N_6294,N_5533,N_5358);
or U6295 (N_6295,N_4939,N_5477);
nand U6296 (N_6296,N_5196,N_4918);
nor U6297 (N_6297,N_5024,N_4957);
nor U6298 (N_6298,N_5429,N_5289);
nor U6299 (N_6299,N_4934,N_5229);
nor U6300 (N_6300,N_5265,N_4852);
or U6301 (N_6301,N_5131,N_5305);
and U6302 (N_6302,N_5467,N_5215);
and U6303 (N_6303,N_5586,N_5410);
and U6304 (N_6304,N_4962,N_4935);
nand U6305 (N_6305,N_4814,N_5444);
and U6306 (N_6306,N_5162,N_4842);
nor U6307 (N_6307,N_5506,N_4828);
or U6308 (N_6308,N_4867,N_5409);
and U6309 (N_6309,N_5438,N_5085);
xnor U6310 (N_6310,N_5059,N_5272);
nand U6311 (N_6311,N_4856,N_5012);
xor U6312 (N_6312,N_5201,N_5312);
or U6313 (N_6313,N_5109,N_5166);
xnor U6314 (N_6314,N_5524,N_5432);
nor U6315 (N_6315,N_5460,N_5582);
or U6316 (N_6316,N_4856,N_5121);
nor U6317 (N_6317,N_5419,N_5333);
nor U6318 (N_6318,N_5582,N_5529);
nand U6319 (N_6319,N_5510,N_5021);
and U6320 (N_6320,N_5094,N_5255);
or U6321 (N_6321,N_5319,N_5265);
nor U6322 (N_6322,N_4880,N_5344);
nor U6323 (N_6323,N_5042,N_5539);
and U6324 (N_6324,N_5514,N_5317);
nand U6325 (N_6325,N_4997,N_5048);
nand U6326 (N_6326,N_5019,N_5508);
and U6327 (N_6327,N_5472,N_4957);
xnor U6328 (N_6328,N_5137,N_5469);
or U6329 (N_6329,N_5095,N_4981);
and U6330 (N_6330,N_5599,N_5099);
xnor U6331 (N_6331,N_5366,N_4940);
or U6332 (N_6332,N_4885,N_5434);
nand U6333 (N_6333,N_5126,N_5259);
nor U6334 (N_6334,N_4932,N_5453);
nand U6335 (N_6335,N_5377,N_4808);
nand U6336 (N_6336,N_4828,N_4823);
nor U6337 (N_6337,N_5336,N_5210);
or U6338 (N_6338,N_5338,N_4995);
or U6339 (N_6339,N_4952,N_5250);
nand U6340 (N_6340,N_5026,N_5070);
xor U6341 (N_6341,N_4973,N_5119);
or U6342 (N_6342,N_5379,N_5399);
xor U6343 (N_6343,N_5477,N_5532);
nand U6344 (N_6344,N_5378,N_5283);
nor U6345 (N_6345,N_5561,N_4829);
nand U6346 (N_6346,N_4977,N_4967);
and U6347 (N_6347,N_5045,N_5170);
xor U6348 (N_6348,N_5285,N_5205);
or U6349 (N_6349,N_5571,N_5496);
nor U6350 (N_6350,N_4866,N_5468);
and U6351 (N_6351,N_5236,N_4972);
and U6352 (N_6352,N_5444,N_5137);
xnor U6353 (N_6353,N_5544,N_5585);
nand U6354 (N_6354,N_5374,N_4822);
and U6355 (N_6355,N_5033,N_4905);
xnor U6356 (N_6356,N_4957,N_5383);
nand U6357 (N_6357,N_4906,N_5068);
and U6358 (N_6358,N_4960,N_4820);
nor U6359 (N_6359,N_5141,N_5475);
and U6360 (N_6360,N_4961,N_5392);
and U6361 (N_6361,N_4865,N_4981);
and U6362 (N_6362,N_4823,N_5018);
nor U6363 (N_6363,N_4956,N_4897);
nand U6364 (N_6364,N_5466,N_5586);
or U6365 (N_6365,N_4871,N_5228);
nand U6366 (N_6366,N_5284,N_5546);
nand U6367 (N_6367,N_5211,N_5550);
xnor U6368 (N_6368,N_5261,N_5568);
nor U6369 (N_6369,N_4977,N_5580);
or U6370 (N_6370,N_5323,N_5212);
or U6371 (N_6371,N_5430,N_5276);
nor U6372 (N_6372,N_5060,N_5192);
nand U6373 (N_6373,N_5266,N_5505);
xor U6374 (N_6374,N_5228,N_5051);
nor U6375 (N_6375,N_4882,N_5453);
nor U6376 (N_6376,N_5377,N_5536);
or U6377 (N_6377,N_4932,N_5599);
xor U6378 (N_6378,N_4834,N_4917);
nand U6379 (N_6379,N_5425,N_5200);
xor U6380 (N_6380,N_5060,N_4911);
nor U6381 (N_6381,N_5422,N_5571);
or U6382 (N_6382,N_5234,N_5473);
xor U6383 (N_6383,N_4849,N_5465);
nand U6384 (N_6384,N_4951,N_5164);
or U6385 (N_6385,N_4877,N_5366);
xnor U6386 (N_6386,N_5172,N_5181);
or U6387 (N_6387,N_5512,N_4975);
or U6388 (N_6388,N_5037,N_5536);
or U6389 (N_6389,N_5126,N_5255);
and U6390 (N_6390,N_5577,N_5049);
nand U6391 (N_6391,N_5215,N_5208);
or U6392 (N_6392,N_5411,N_5149);
xor U6393 (N_6393,N_5395,N_4817);
nand U6394 (N_6394,N_5317,N_5396);
xor U6395 (N_6395,N_5280,N_5545);
or U6396 (N_6396,N_5515,N_5570);
or U6397 (N_6397,N_4975,N_5002);
or U6398 (N_6398,N_5443,N_5116);
xor U6399 (N_6399,N_5248,N_5427);
nand U6400 (N_6400,N_5972,N_6202);
nor U6401 (N_6401,N_6266,N_6075);
or U6402 (N_6402,N_5956,N_5736);
xnor U6403 (N_6403,N_6107,N_6271);
nand U6404 (N_6404,N_5893,N_6272);
and U6405 (N_6405,N_6285,N_6101);
xnor U6406 (N_6406,N_5809,N_6389);
nor U6407 (N_6407,N_5955,N_6180);
and U6408 (N_6408,N_6134,N_6123);
xnor U6409 (N_6409,N_5984,N_6380);
or U6410 (N_6410,N_6236,N_6035);
or U6411 (N_6411,N_6304,N_6197);
nor U6412 (N_6412,N_6033,N_6296);
or U6413 (N_6413,N_5768,N_6354);
and U6414 (N_6414,N_5941,N_5989);
and U6415 (N_6415,N_5896,N_6032);
and U6416 (N_6416,N_5954,N_5745);
or U6417 (N_6417,N_5812,N_5654);
or U6418 (N_6418,N_6143,N_6251);
and U6419 (N_6419,N_5789,N_6394);
nor U6420 (N_6420,N_5651,N_5765);
or U6421 (N_6421,N_5904,N_5925);
nand U6422 (N_6422,N_6274,N_5773);
and U6423 (N_6423,N_5806,N_5817);
nand U6424 (N_6424,N_5769,N_6083);
or U6425 (N_6425,N_5946,N_6203);
or U6426 (N_6426,N_5790,N_5938);
and U6427 (N_6427,N_6163,N_6200);
and U6428 (N_6428,N_6284,N_5723);
nand U6429 (N_6429,N_6115,N_5646);
or U6430 (N_6430,N_5758,N_6239);
nor U6431 (N_6431,N_6315,N_6241);
nor U6432 (N_6432,N_5663,N_6109);
and U6433 (N_6433,N_6162,N_5625);
or U6434 (N_6434,N_6377,N_5604);
nor U6435 (N_6435,N_5726,N_6317);
xnor U6436 (N_6436,N_6055,N_6141);
nor U6437 (N_6437,N_6299,N_6145);
xnor U6438 (N_6438,N_6081,N_6137);
and U6439 (N_6439,N_5824,N_5650);
or U6440 (N_6440,N_6103,N_5722);
or U6441 (N_6441,N_6124,N_5831);
xnor U6442 (N_6442,N_6046,N_6228);
nand U6443 (N_6443,N_6015,N_5708);
xor U6444 (N_6444,N_5690,N_5832);
nor U6445 (N_6445,N_6003,N_5703);
nand U6446 (N_6446,N_5815,N_5655);
and U6447 (N_6447,N_5600,N_6392);
or U6448 (N_6448,N_6240,N_5905);
and U6449 (N_6449,N_5665,N_5866);
xnor U6450 (N_6450,N_5908,N_5803);
xor U6451 (N_6451,N_6211,N_6154);
nor U6452 (N_6452,N_5686,N_5825);
xor U6453 (N_6453,N_6378,N_5906);
or U6454 (N_6454,N_5672,N_6279);
nand U6455 (N_6455,N_5701,N_5776);
and U6456 (N_6456,N_5932,N_6136);
or U6457 (N_6457,N_5966,N_5627);
nand U6458 (N_6458,N_5673,N_5890);
nand U6459 (N_6459,N_5689,N_6070);
xor U6460 (N_6460,N_5977,N_6301);
or U6461 (N_6461,N_5878,N_5659);
and U6462 (N_6462,N_5747,N_5630);
and U6463 (N_6463,N_5664,N_6289);
or U6464 (N_6464,N_6018,N_5729);
nor U6465 (N_6465,N_5709,N_5897);
nand U6466 (N_6466,N_6077,N_6363);
or U6467 (N_6467,N_6269,N_6359);
or U6468 (N_6468,N_5999,N_5939);
nor U6469 (N_6469,N_6206,N_5711);
or U6470 (N_6470,N_6097,N_5800);
xnor U6471 (N_6471,N_5674,N_5828);
nand U6472 (N_6472,N_6059,N_5750);
and U6473 (N_6473,N_5784,N_5931);
nand U6474 (N_6474,N_5762,N_5850);
or U6475 (N_6475,N_6114,N_6256);
or U6476 (N_6476,N_5887,N_5614);
and U6477 (N_6477,N_5740,N_5732);
nor U6478 (N_6478,N_6370,N_6331);
or U6479 (N_6479,N_6342,N_6045);
nor U6480 (N_6480,N_6234,N_5872);
or U6481 (N_6481,N_6351,N_5863);
and U6482 (N_6482,N_5668,N_5691);
or U6483 (N_6483,N_5652,N_6156);
xnor U6484 (N_6484,N_5658,N_5678);
nor U6485 (N_6485,N_5751,N_5959);
nor U6486 (N_6486,N_6001,N_6335);
xnor U6487 (N_6487,N_6327,N_6017);
or U6488 (N_6488,N_6161,N_5763);
nor U6489 (N_6489,N_5934,N_5618);
or U6490 (N_6490,N_6312,N_6330);
and U6491 (N_6491,N_6339,N_6012);
nor U6492 (N_6492,N_5982,N_6082);
xor U6493 (N_6493,N_5936,N_6085);
nand U6494 (N_6494,N_6053,N_5877);
xor U6495 (N_6495,N_5929,N_6058);
xor U6496 (N_6496,N_6369,N_5834);
nor U6497 (N_6497,N_5759,N_6157);
nor U6498 (N_6498,N_5841,N_5707);
nand U6499 (N_6499,N_6158,N_6292);
nor U6500 (N_6500,N_6374,N_6334);
nor U6501 (N_6501,N_6128,N_5993);
xnor U6502 (N_6502,N_5653,N_5602);
and U6503 (N_6503,N_6006,N_5601);
and U6504 (N_6504,N_5608,N_5821);
xnor U6505 (N_6505,N_6386,N_6319);
xor U6506 (N_6506,N_6019,N_6298);
and U6507 (N_6507,N_6013,N_6261);
or U6508 (N_6508,N_5861,N_5813);
nand U6509 (N_6509,N_6125,N_5948);
nor U6510 (N_6510,N_6066,N_6036);
xnor U6511 (N_6511,N_6108,N_5749);
xnor U6512 (N_6512,N_6004,N_5901);
nor U6513 (N_6513,N_5923,N_5842);
xor U6514 (N_6514,N_5793,N_6345);
nor U6515 (N_6515,N_5677,N_6166);
xor U6516 (N_6516,N_6297,N_6350);
or U6517 (N_6517,N_5805,N_5802);
nor U6518 (N_6518,N_6325,N_5724);
nor U6519 (N_6519,N_6185,N_5868);
nand U6520 (N_6520,N_6028,N_6138);
and U6521 (N_6521,N_5730,N_5685);
nor U6522 (N_6522,N_6376,N_5657);
and U6523 (N_6523,N_5717,N_6218);
nor U6524 (N_6524,N_6153,N_6391);
nor U6525 (N_6525,N_5770,N_6179);
and U6526 (N_6526,N_5857,N_6048);
or U6527 (N_6527,N_5694,N_6144);
or U6528 (N_6528,N_6122,N_6183);
nand U6529 (N_6529,N_5808,N_5693);
or U6530 (N_6530,N_6398,N_6054);
xnor U6531 (N_6531,N_6191,N_5830);
nand U6532 (N_6532,N_6364,N_5943);
or U6533 (N_6533,N_5843,N_6399);
nor U6534 (N_6534,N_5788,N_6027);
nand U6535 (N_6535,N_6302,N_6135);
xor U6536 (N_6536,N_6201,N_5801);
and U6537 (N_6537,N_5715,N_6366);
or U6538 (N_6538,N_6352,N_6367);
and U6539 (N_6539,N_6341,N_5860);
xor U6540 (N_6540,N_6061,N_6190);
xor U6541 (N_6541,N_6009,N_6320);
nor U6542 (N_6542,N_5628,N_6076);
and U6543 (N_6543,N_5957,N_6310);
or U6544 (N_6544,N_5633,N_5835);
nand U6545 (N_6545,N_6385,N_5848);
xnor U6546 (N_6546,N_5675,N_5682);
nand U6547 (N_6547,N_5692,N_6287);
nor U6548 (N_6548,N_5649,N_6008);
and U6549 (N_6549,N_5629,N_6348);
and U6550 (N_6550,N_5699,N_5656);
xor U6551 (N_6551,N_6307,N_5944);
and U6552 (N_6552,N_6247,N_6333);
nand U6553 (N_6553,N_5615,N_6005);
nand U6554 (N_6554,N_6365,N_5710);
and U6555 (N_6555,N_5980,N_6071);
or U6556 (N_6556,N_5611,N_5937);
nor U6557 (N_6557,N_6324,N_6024);
nor U6558 (N_6558,N_5713,N_6002);
xnor U6559 (N_6559,N_6067,N_6209);
xnor U6560 (N_6560,N_5735,N_6252);
and U6561 (N_6561,N_6192,N_6074);
and U6562 (N_6562,N_6257,N_5919);
xnor U6563 (N_6563,N_6381,N_5823);
or U6564 (N_6564,N_5774,N_5852);
and U6565 (N_6565,N_5731,N_5643);
or U6566 (N_6566,N_6276,N_5928);
nand U6567 (N_6567,N_5609,N_6132);
or U6568 (N_6568,N_6152,N_5782);
xnor U6569 (N_6569,N_5899,N_6196);
xnor U6570 (N_6570,N_5676,N_6208);
and U6571 (N_6571,N_6215,N_5873);
nor U6572 (N_6572,N_6283,N_5855);
nor U6573 (N_6573,N_6395,N_6250);
and U6574 (N_6574,N_6073,N_5869);
nor U6575 (N_6575,N_6321,N_5926);
or U6576 (N_6576,N_6273,N_6223);
and U6577 (N_6577,N_5666,N_5880);
xnor U6578 (N_6578,N_5916,N_6375);
or U6579 (N_6579,N_6245,N_6121);
nand U6580 (N_6580,N_6233,N_6072);
or U6581 (N_6581,N_5883,N_6219);
nand U6582 (N_6582,N_5617,N_5858);
nand U6583 (N_6583,N_6086,N_5992);
nand U6584 (N_6584,N_5720,N_6323);
or U6585 (N_6585,N_6280,N_6383);
nor U6586 (N_6586,N_5733,N_6170);
or U6587 (N_6587,N_6199,N_6393);
or U6588 (N_6588,N_5727,N_5838);
or U6589 (N_6589,N_5846,N_6328);
xnor U6590 (N_6590,N_5684,N_6133);
and U6591 (N_6591,N_6100,N_6318);
and U6592 (N_6592,N_6326,N_6357);
and U6593 (N_6593,N_5647,N_6249);
xor U6594 (N_6594,N_5623,N_6089);
nor U6595 (N_6595,N_5990,N_6300);
nor U6596 (N_6596,N_5799,N_6104);
and U6597 (N_6597,N_6131,N_5621);
nand U6598 (N_6598,N_5741,N_5661);
xor U6599 (N_6599,N_5968,N_6142);
xor U6600 (N_6600,N_5914,N_6155);
or U6601 (N_6601,N_6244,N_6237);
nor U6602 (N_6602,N_5854,N_6217);
nor U6603 (N_6603,N_5780,N_6288);
xor U6604 (N_6604,N_6396,N_5620);
or U6605 (N_6605,N_5986,N_5764);
nor U6606 (N_6606,N_5697,N_5795);
and U6607 (N_6607,N_6255,N_5997);
xnor U6608 (N_6608,N_5920,N_5907);
xnor U6609 (N_6609,N_6322,N_5882);
nand U6610 (N_6610,N_6204,N_6338);
nand U6611 (N_6611,N_6306,N_5881);
or U6612 (N_6612,N_5744,N_5874);
xnor U6613 (N_6613,N_5639,N_6213);
nand U6614 (N_6614,N_6043,N_6216);
or U6615 (N_6615,N_5965,N_6181);
and U6616 (N_6616,N_6106,N_5777);
xor U6617 (N_6617,N_6177,N_6016);
nand U6618 (N_6618,N_5772,N_5903);
and U6619 (N_6619,N_5670,N_6308);
or U6620 (N_6620,N_6102,N_5819);
nand U6621 (N_6621,N_5760,N_6176);
nand U6622 (N_6622,N_5895,N_6096);
and U6623 (N_6623,N_5798,N_5753);
nand U6624 (N_6624,N_5644,N_5962);
or U6625 (N_6625,N_5859,N_6021);
xor U6626 (N_6626,N_6270,N_5702);
nor U6627 (N_6627,N_5851,N_6092);
nor U6628 (N_6628,N_5876,N_6091);
xnor U6629 (N_6629,N_6062,N_6022);
nor U6630 (N_6630,N_5910,N_5742);
nor U6631 (N_6631,N_5683,N_6212);
nand U6632 (N_6632,N_6011,N_5667);
or U6633 (N_6633,N_5743,N_6373);
or U6634 (N_6634,N_5947,N_5884);
and U6635 (N_6635,N_6172,N_5983);
nand U6636 (N_6636,N_5738,N_5756);
xnor U6637 (N_6637,N_5953,N_5626);
and U6638 (N_6638,N_6311,N_5721);
and U6639 (N_6639,N_6039,N_6242);
and U6640 (N_6640,N_5778,N_6064);
nor U6641 (N_6641,N_5839,N_5767);
xnor U6642 (N_6642,N_6260,N_5734);
nor U6643 (N_6643,N_5669,N_6079);
xor U6644 (N_6644,N_5960,N_6282);
nor U6645 (N_6645,N_5616,N_5818);
and U6646 (N_6646,N_6175,N_6355);
xor U6647 (N_6647,N_5791,N_6194);
nand U6648 (N_6648,N_6329,N_5642);
nor U6649 (N_6649,N_5648,N_5606);
nand U6650 (N_6650,N_6029,N_5900);
and U6651 (N_6651,N_6184,N_5787);
nand U6652 (N_6652,N_6160,N_5991);
xnor U6653 (N_6653,N_5775,N_6281);
nand U6654 (N_6654,N_6238,N_5797);
xor U6655 (N_6655,N_6034,N_5885);
and U6656 (N_6656,N_6253,N_5603);
xor U6657 (N_6657,N_6303,N_5949);
xnor U6658 (N_6658,N_5969,N_5892);
and U6659 (N_6659,N_5636,N_5624);
nor U6660 (N_6660,N_6278,N_6226);
or U6661 (N_6661,N_6093,N_6314);
xor U6662 (N_6662,N_6174,N_6056);
xor U6663 (N_6663,N_6313,N_6246);
and U6664 (N_6664,N_6353,N_5739);
nor U6665 (N_6665,N_6150,N_5902);
or U6666 (N_6666,N_6116,N_5631);
or U6667 (N_6667,N_5662,N_6340);
or U6668 (N_6668,N_5961,N_5725);
and U6669 (N_6669,N_6025,N_6263);
nand U6670 (N_6670,N_5958,N_6126);
xor U6671 (N_6671,N_5967,N_6294);
nand U6672 (N_6672,N_6205,N_5975);
or U6673 (N_6673,N_6254,N_6007);
or U6674 (N_6674,N_6235,N_6291);
nor U6675 (N_6675,N_6052,N_5964);
nand U6676 (N_6676,N_6265,N_5688);
or U6677 (N_6677,N_6182,N_5605);
nand U6678 (N_6678,N_5637,N_5783);
nand U6679 (N_6679,N_5706,N_6361);
and U6680 (N_6680,N_5640,N_5847);
xnor U6681 (N_6681,N_5864,N_6264);
and U6682 (N_6682,N_5870,N_5804);
nor U6683 (N_6683,N_6224,N_6095);
nor U6684 (N_6684,N_6368,N_6173);
nand U6685 (N_6685,N_5998,N_6069);
nor U6686 (N_6686,N_5974,N_5826);
nand U6687 (N_6687,N_6337,N_6065);
xnor U6688 (N_6688,N_6110,N_5865);
nor U6689 (N_6689,N_6305,N_5833);
nand U6690 (N_6690,N_5766,N_6127);
xnor U6691 (N_6691,N_6293,N_6198);
nand U6692 (N_6692,N_5971,N_6099);
nor U6693 (N_6693,N_6120,N_5814);
nand U6694 (N_6694,N_5716,N_6139);
nor U6695 (N_6695,N_5811,N_6068);
xor U6696 (N_6696,N_6010,N_6078);
and U6697 (N_6697,N_5718,N_6316);
or U6698 (N_6698,N_5779,N_5935);
and U6699 (N_6699,N_6372,N_6332);
or U6700 (N_6700,N_6047,N_5886);
nor U6701 (N_6701,N_5681,N_6087);
nor U6702 (N_6702,N_5719,N_5912);
nor U6703 (N_6703,N_5705,N_6189);
xor U6704 (N_6704,N_5862,N_6346);
xnor U6705 (N_6705,N_5822,N_6040);
nand U6706 (N_6706,N_6268,N_6113);
or U6707 (N_6707,N_6384,N_6397);
and U6708 (N_6708,N_5927,N_6038);
nor U6709 (N_6709,N_6230,N_6362);
nand U6710 (N_6710,N_6063,N_5695);
nor U6711 (N_6711,N_5728,N_6171);
nor U6712 (N_6712,N_5951,N_5911);
and U6713 (N_6713,N_6020,N_5660);
nor U6714 (N_6714,N_6210,N_5645);
or U6715 (N_6715,N_6258,N_5994);
and U6716 (N_6716,N_5849,N_5891);
xnor U6717 (N_6717,N_5700,N_6037);
and U6718 (N_6718,N_5755,N_6186);
and U6719 (N_6719,N_6358,N_6229);
or U6720 (N_6720,N_6275,N_5622);
nor U6721 (N_6721,N_6214,N_6050);
xnor U6722 (N_6722,N_6105,N_6388);
xnor U6723 (N_6723,N_5714,N_6243);
and U6724 (N_6724,N_6000,N_6387);
nand U6725 (N_6725,N_6031,N_6360);
and U6726 (N_6726,N_6207,N_5837);
or U6727 (N_6727,N_5856,N_5942);
nor U6728 (N_6728,N_5613,N_6231);
and U6729 (N_6729,N_5781,N_5829);
nand U6730 (N_6730,N_5634,N_6349);
xnor U6731 (N_6731,N_6051,N_6347);
or U6732 (N_6732,N_5638,N_6187);
xnor U6733 (N_6733,N_5752,N_6112);
nand U6734 (N_6734,N_5687,N_5921);
xnor U6735 (N_6735,N_5754,N_5922);
nor U6736 (N_6736,N_6232,N_6343);
or U6737 (N_6737,N_5924,N_6248);
and U6738 (N_6738,N_5940,N_6149);
nand U6739 (N_6739,N_5845,N_6111);
nor U6740 (N_6740,N_6193,N_6188);
or U6741 (N_6741,N_5836,N_5794);
or U6742 (N_6742,N_6041,N_5792);
xnor U6743 (N_6743,N_5950,N_5712);
nor U6744 (N_6744,N_6195,N_5827);
or U6745 (N_6745,N_5978,N_5748);
and U6746 (N_6746,N_6026,N_5820);
and U6747 (N_6747,N_5619,N_5796);
xnor U6748 (N_6748,N_5671,N_6165);
or U6749 (N_6749,N_6098,N_6042);
nor U6750 (N_6750,N_5879,N_5952);
or U6751 (N_6751,N_6030,N_6286);
and U6752 (N_6752,N_5889,N_6295);
nand U6753 (N_6753,N_5679,N_5632);
xnor U6754 (N_6754,N_6379,N_5963);
and U6755 (N_6755,N_6014,N_6023);
or U6756 (N_6756,N_5973,N_6119);
xnor U6757 (N_6757,N_6140,N_5981);
xnor U6758 (N_6758,N_6277,N_6080);
and U6759 (N_6759,N_5894,N_6262);
or U6760 (N_6760,N_6090,N_6390);
or U6761 (N_6761,N_5888,N_6344);
nor U6762 (N_6762,N_6221,N_5985);
nor U6763 (N_6763,N_6088,N_6147);
nor U6764 (N_6764,N_5786,N_6220);
nand U6765 (N_6765,N_6356,N_5945);
nor U6766 (N_6766,N_5875,N_6044);
xnor U6767 (N_6767,N_5680,N_6227);
or U6768 (N_6768,N_6267,N_5607);
or U6769 (N_6769,N_6129,N_5704);
and U6770 (N_6770,N_5641,N_5810);
xor U6771 (N_6771,N_6118,N_6057);
and U6772 (N_6772,N_5915,N_5635);
and U6773 (N_6773,N_5995,N_5816);
nor U6774 (N_6774,N_5771,N_6117);
and U6775 (N_6775,N_6222,N_6336);
xnor U6776 (N_6776,N_5871,N_6371);
and U6777 (N_6777,N_5840,N_6225);
nor U6778 (N_6778,N_5909,N_6151);
nand U6779 (N_6779,N_5746,N_6164);
nor U6780 (N_6780,N_5844,N_6060);
xor U6781 (N_6781,N_5898,N_6148);
xor U6782 (N_6782,N_5807,N_6168);
or U6783 (N_6783,N_5996,N_5696);
xor U6784 (N_6784,N_5698,N_5987);
and U6785 (N_6785,N_5917,N_5737);
nor U6786 (N_6786,N_5933,N_6382);
nor U6787 (N_6787,N_5867,N_6167);
xnor U6788 (N_6788,N_5976,N_6309);
and U6789 (N_6789,N_5913,N_5930);
or U6790 (N_6790,N_5988,N_6178);
nand U6791 (N_6791,N_5761,N_6146);
xor U6792 (N_6792,N_5979,N_6084);
and U6793 (N_6793,N_6290,N_6094);
nand U6794 (N_6794,N_5610,N_5918);
or U6795 (N_6795,N_5612,N_5970);
and U6796 (N_6796,N_6049,N_6159);
nand U6797 (N_6797,N_6169,N_6259);
and U6798 (N_6798,N_5785,N_6130);
nand U6799 (N_6799,N_5853,N_5757);
and U6800 (N_6800,N_6152,N_5887);
and U6801 (N_6801,N_6211,N_6383);
and U6802 (N_6802,N_5981,N_5926);
xnor U6803 (N_6803,N_6345,N_6101);
and U6804 (N_6804,N_6289,N_6105);
or U6805 (N_6805,N_5694,N_5957);
xnor U6806 (N_6806,N_5622,N_5742);
xor U6807 (N_6807,N_6297,N_5894);
and U6808 (N_6808,N_6368,N_5978);
nor U6809 (N_6809,N_6160,N_5760);
xnor U6810 (N_6810,N_5920,N_6356);
nand U6811 (N_6811,N_5795,N_6117);
or U6812 (N_6812,N_5797,N_6357);
nor U6813 (N_6813,N_5604,N_6087);
nor U6814 (N_6814,N_5904,N_5944);
nand U6815 (N_6815,N_6113,N_5676);
nor U6816 (N_6816,N_5898,N_5905);
and U6817 (N_6817,N_6313,N_6324);
nor U6818 (N_6818,N_5759,N_6293);
and U6819 (N_6819,N_5908,N_6162);
nor U6820 (N_6820,N_6067,N_5821);
or U6821 (N_6821,N_6239,N_5614);
and U6822 (N_6822,N_5627,N_5716);
or U6823 (N_6823,N_5666,N_5898);
and U6824 (N_6824,N_5675,N_5922);
or U6825 (N_6825,N_6228,N_5768);
or U6826 (N_6826,N_5698,N_5763);
nor U6827 (N_6827,N_5791,N_5624);
nand U6828 (N_6828,N_5994,N_6106);
and U6829 (N_6829,N_6214,N_6179);
xor U6830 (N_6830,N_6219,N_6243);
nand U6831 (N_6831,N_5695,N_6022);
nor U6832 (N_6832,N_6034,N_5746);
nand U6833 (N_6833,N_6211,N_6113);
nor U6834 (N_6834,N_5899,N_6273);
or U6835 (N_6835,N_5726,N_6037);
nor U6836 (N_6836,N_6158,N_5921);
nor U6837 (N_6837,N_6273,N_6149);
nand U6838 (N_6838,N_5986,N_5853);
or U6839 (N_6839,N_5895,N_6019);
nand U6840 (N_6840,N_6316,N_5968);
or U6841 (N_6841,N_5940,N_6017);
nor U6842 (N_6842,N_6196,N_6343);
or U6843 (N_6843,N_5739,N_6060);
or U6844 (N_6844,N_6301,N_6034);
or U6845 (N_6845,N_6125,N_5965);
xor U6846 (N_6846,N_5752,N_6060);
nor U6847 (N_6847,N_6240,N_5646);
nand U6848 (N_6848,N_6127,N_6092);
nor U6849 (N_6849,N_6188,N_5919);
nand U6850 (N_6850,N_5763,N_6198);
and U6851 (N_6851,N_5614,N_5645);
nor U6852 (N_6852,N_5832,N_5975);
or U6853 (N_6853,N_5902,N_5766);
nor U6854 (N_6854,N_5989,N_5791);
and U6855 (N_6855,N_5935,N_6265);
nand U6856 (N_6856,N_5652,N_5756);
and U6857 (N_6857,N_5849,N_5874);
or U6858 (N_6858,N_5769,N_6078);
nor U6859 (N_6859,N_6396,N_5713);
xnor U6860 (N_6860,N_6243,N_5822);
nor U6861 (N_6861,N_6192,N_6165);
and U6862 (N_6862,N_5892,N_5832);
and U6863 (N_6863,N_5852,N_6024);
nand U6864 (N_6864,N_5812,N_5741);
nor U6865 (N_6865,N_6252,N_5924);
xnor U6866 (N_6866,N_5931,N_5615);
and U6867 (N_6867,N_5614,N_5855);
or U6868 (N_6868,N_5718,N_5956);
nor U6869 (N_6869,N_5658,N_5786);
nor U6870 (N_6870,N_6339,N_5729);
or U6871 (N_6871,N_5967,N_5628);
nand U6872 (N_6872,N_6158,N_6285);
and U6873 (N_6873,N_6140,N_5819);
xnor U6874 (N_6874,N_6102,N_5828);
or U6875 (N_6875,N_5942,N_5960);
and U6876 (N_6876,N_5975,N_5615);
nor U6877 (N_6877,N_5792,N_5967);
or U6878 (N_6878,N_6156,N_5975);
xor U6879 (N_6879,N_6387,N_6067);
or U6880 (N_6880,N_6076,N_5648);
xnor U6881 (N_6881,N_5894,N_6087);
and U6882 (N_6882,N_6140,N_5997);
or U6883 (N_6883,N_6246,N_6176);
and U6884 (N_6884,N_5660,N_5655);
xnor U6885 (N_6885,N_6276,N_5637);
and U6886 (N_6886,N_5687,N_5795);
or U6887 (N_6887,N_5726,N_6166);
xor U6888 (N_6888,N_5744,N_6058);
xnor U6889 (N_6889,N_5970,N_6172);
xor U6890 (N_6890,N_6168,N_6150);
or U6891 (N_6891,N_5953,N_6077);
xnor U6892 (N_6892,N_5823,N_5695);
nand U6893 (N_6893,N_5890,N_5992);
nand U6894 (N_6894,N_5620,N_6025);
nor U6895 (N_6895,N_5670,N_5820);
and U6896 (N_6896,N_5655,N_5657);
or U6897 (N_6897,N_6152,N_5995);
and U6898 (N_6898,N_5625,N_6380);
or U6899 (N_6899,N_6384,N_6186);
xnor U6900 (N_6900,N_6038,N_6129);
nand U6901 (N_6901,N_5864,N_6237);
or U6902 (N_6902,N_5676,N_5874);
and U6903 (N_6903,N_6150,N_6084);
and U6904 (N_6904,N_6337,N_6315);
xor U6905 (N_6905,N_6014,N_5629);
and U6906 (N_6906,N_5978,N_5952);
or U6907 (N_6907,N_6062,N_6091);
xnor U6908 (N_6908,N_5952,N_5999);
and U6909 (N_6909,N_6064,N_5892);
and U6910 (N_6910,N_6144,N_5879);
xor U6911 (N_6911,N_5686,N_5817);
xnor U6912 (N_6912,N_6030,N_6252);
or U6913 (N_6913,N_5887,N_6096);
nand U6914 (N_6914,N_6300,N_6376);
or U6915 (N_6915,N_5761,N_6087);
xor U6916 (N_6916,N_5764,N_6186);
and U6917 (N_6917,N_6336,N_6356);
nand U6918 (N_6918,N_6090,N_6013);
xor U6919 (N_6919,N_5832,N_6143);
or U6920 (N_6920,N_6175,N_6031);
or U6921 (N_6921,N_5689,N_6088);
or U6922 (N_6922,N_6198,N_5757);
or U6923 (N_6923,N_6007,N_5912);
nand U6924 (N_6924,N_6366,N_6160);
xor U6925 (N_6925,N_5802,N_5900);
and U6926 (N_6926,N_5660,N_6121);
or U6927 (N_6927,N_6333,N_5995);
and U6928 (N_6928,N_5864,N_6044);
nand U6929 (N_6929,N_5893,N_6005);
nand U6930 (N_6930,N_6134,N_5731);
and U6931 (N_6931,N_6243,N_6253);
or U6932 (N_6932,N_6159,N_6082);
xor U6933 (N_6933,N_5990,N_5712);
or U6934 (N_6934,N_6129,N_6343);
nor U6935 (N_6935,N_6330,N_5884);
nand U6936 (N_6936,N_6289,N_6137);
and U6937 (N_6937,N_6030,N_6260);
or U6938 (N_6938,N_6123,N_6140);
nor U6939 (N_6939,N_6043,N_5624);
nor U6940 (N_6940,N_6065,N_6229);
or U6941 (N_6941,N_6142,N_6229);
nor U6942 (N_6942,N_6148,N_6038);
nor U6943 (N_6943,N_5884,N_6283);
nor U6944 (N_6944,N_6051,N_5871);
xor U6945 (N_6945,N_6365,N_6063);
nor U6946 (N_6946,N_5810,N_5794);
nor U6947 (N_6947,N_6130,N_6394);
nand U6948 (N_6948,N_6067,N_5865);
nand U6949 (N_6949,N_5651,N_5798);
nand U6950 (N_6950,N_5648,N_6119);
nor U6951 (N_6951,N_6009,N_6024);
nand U6952 (N_6952,N_6285,N_5977);
xnor U6953 (N_6953,N_6021,N_5892);
and U6954 (N_6954,N_5781,N_6278);
nor U6955 (N_6955,N_6337,N_6150);
or U6956 (N_6956,N_6356,N_5829);
and U6957 (N_6957,N_6303,N_5892);
xnor U6958 (N_6958,N_5865,N_6017);
nor U6959 (N_6959,N_6067,N_6392);
and U6960 (N_6960,N_5986,N_6090);
nand U6961 (N_6961,N_5957,N_5699);
or U6962 (N_6962,N_5843,N_6390);
nor U6963 (N_6963,N_5993,N_6058);
and U6964 (N_6964,N_5892,N_6234);
or U6965 (N_6965,N_5949,N_6030);
or U6966 (N_6966,N_5854,N_6244);
nand U6967 (N_6967,N_5828,N_5677);
nand U6968 (N_6968,N_6197,N_6094);
nand U6969 (N_6969,N_6270,N_5810);
nor U6970 (N_6970,N_5759,N_5886);
xor U6971 (N_6971,N_5608,N_6342);
and U6972 (N_6972,N_6160,N_6068);
or U6973 (N_6973,N_6213,N_6163);
nor U6974 (N_6974,N_6349,N_5774);
and U6975 (N_6975,N_5906,N_6051);
or U6976 (N_6976,N_5891,N_5692);
nor U6977 (N_6977,N_5980,N_5975);
and U6978 (N_6978,N_5915,N_6080);
and U6979 (N_6979,N_5999,N_5936);
or U6980 (N_6980,N_5644,N_5620);
or U6981 (N_6981,N_5704,N_5866);
or U6982 (N_6982,N_5996,N_6002);
or U6983 (N_6983,N_6202,N_5859);
nand U6984 (N_6984,N_5876,N_5630);
nor U6985 (N_6985,N_5722,N_5913);
nor U6986 (N_6986,N_5763,N_6230);
nor U6987 (N_6987,N_6391,N_5818);
xor U6988 (N_6988,N_6023,N_5951);
nand U6989 (N_6989,N_6213,N_6032);
xor U6990 (N_6990,N_6309,N_5836);
and U6991 (N_6991,N_5668,N_5640);
nand U6992 (N_6992,N_5832,N_5819);
nor U6993 (N_6993,N_5977,N_6173);
xnor U6994 (N_6994,N_6012,N_6176);
nand U6995 (N_6995,N_5894,N_5648);
nand U6996 (N_6996,N_6071,N_5618);
or U6997 (N_6997,N_6066,N_6330);
xor U6998 (N_6998,N_6338,N_5681);
or U6999 (N_6999,N_6045,N_5665);
or U7000 (N_7000,N_5645,N_5707);
and U7001 (N_7001,N_6242,N_5633);
xnor U7002 (N_7002,N_6296,N_6275);
or U7003 (N_7003,N_6038,N_6143);
and U7004 (N_7004,N_6027,N_6334);
nor U7005 (N_7005,N_6379,N_6145);
nand U7006 (N_7006,N_5675,N_6164);
and U7007 (N_7007,N_6241,N_6127);
nor U7008 (N_7008,N_5626,N_6090);
xnor U7009 (N_7009,N_6113,N_6315);
or U7010 (N_7010,N_6374,N_5938);
nor U7011 (N_7011,N_5813,N_5975);
or U7012 (N_7012,N_5612,N_5627);
xor U7013 (N_7013,N_6249,N_6226);
xnor U7014 (N_7014,N_5634,N_5904);
and U7015 (N_7015,N_6198,N_6245);
nor U7016 (N_7016,N_5894,N_5780);
or U7017 (N_7017,N_5769,N_5656);
nor U7018 (N_7018,N_6144,N_6152);
xnor U7019 (N_7019,N_6383,N_6065);
nor U7020 (N_7020,N_6341,N_6306);
nor U7021 (N_7021,N_6023,N_6082);
and U7022 (N_7022,N_6227,N_5844);
and U7023 (N_7023,N_5851,N_6124);
xor U7024 (N_7024,N_5986,N_5851);
nor U7025 (N_7025,N_6038,N_6181);
nand U7026 (N_7026,N_5902,N_5948);
xnor U7027 (N_7027,N_6040,N_5801);
nor U7028 (N_7028,N_5686,N_5857);
or U7029 (N_7029,N_5672,N_5899);
nor U7030 (N_7030,N_5881,N_5902);
xor U7031 (N_7031,N_6146,N_5776);
and U7032 (N_7032,N_5811,N_5682);
or U7033 (N_7033,N_6291,N_5694);
nor U7034 (N_7034,N_5656,N_6174);
or U7035 (N_7035,N_5608,N_5978);
nand U7036 (N_7036,N_6377,N_5689);
or U7037 (N_7037,N_6105,N_5871);
or U7038 (N_7038,N_6234,N_6210);
nand U7039 (N_7039,N_6303,N_5684);
nor U7040 (N_7040,N_6234,N_5662);
or U7041 (N_7041,N_5938,N_5840);
and U7042 (N_7042,N_6053,N_6365);
nor U7043 (N_7043,N_6067,N_5684);
nand U7044 (N_7044,N_6313,N_5859);
nor U7045 (N_7045,N_5812,N_6360);
nor U7046 (N_7046,N_5843,N_6196);
or U7047 (N_7047,N_5637,N_5605);
nor U7048 (N_7048,N_6102,N_5771);
nand U7049 (N_7049,N_5790,N_6352);
and U7050 (N_7050,N_6134,N_5751);
nor U7051 (N_7051,N_5898,N_5960);
and U7052 (N_7052,N_5766,N_5712);
nand U7053 (N_7053,N_5734,N_6339);
xnor U7054 (N_7054,N_5619,N_6135);
nor U7055 (N_7055,N_5917,N_5958);
nand U7056 (N_7056,N_6146,N_6122);
or U7057 (N_7057,N_6056,N_6020);
xnor U7058 (N_7058,N_6142,N_6061);
nand U7059 (N_7059,N_5710,N_5897);
or U7060 (N_7060,N_5615,N_5744);
or U7061 (N_7061,N_6165,N_6378);
nand U7062 (N_7062,N_6230,N_6311);
or U7063 (N_7063,N_6042,N_5991);
xor U7064 (N_7064,N_5998,N_5881);
or U7065 (N_7065,N_6193,N_5653);
or U7066 (N_7066,N_6115,N_5842);
and U7067 (N_7067,N_5810,N_5697);
and U7068 (N_7068,N_6249,N_6327);
and U7069 (N_7069,N_6161,N_6210);
or U7070 (N_7070,N_6197,N_6232);
nand U7071 (N_7071,N_5811,N_5878);
or U7072 (N_7072,N_5822,N_5608);
xnor U7073 (N_7073,N_5913,N_6249);
xor U7074 (N_7074,N_6363,N_5950);
or U7075 (N_7075,N_6222,N_5767);
or U7076 (N_7076,N_6197,N_6157);
and U7077 (N_7077,N_6143,N_6303);
nand U7078 (N_7078,N_5832,N_6149);
or U7079 (N_7079,N_6134,N_5846);
nor U7080 (N_7080,N_5693,N_6236);
nand U7081 (N_7081,N_5763,N_5729);
and U7082 (N_7082,N_5715,N_5893);
nor U7083 (N_7083,N_6291,N_5686);
nor U7084 (N_7084,N_5840,N_6121);
nor U7085 (N_7085,N_6281,N_5628);
xor U7086 (N_7086,N_5808,N_5959);
nor U7087 (N_7087,N_5733,N_6097);
nand U7088 (N_7088,N_6340,N_5971);
and U7089 (N_7089,N_6349,N_5860);
and U7090 (N_7090,N_6392,N_6329);
and U7091 (N_7091,N_5726,N_5913);
xor U7092 (N_7092,N_5808,N_6317);
and U7093 (N_7093,N_5803,N_5887);
xor U7094 (N_7094,N_5803,N_6148);
or U7095 (N_7095,N_5967,N_5658);
nor U7096 (N_7096,N_5683,N_5812);
nand U7097 (N_7097,N_5618,N_5623);
nand U7098 (N_7098,N_5614,N_5932);
nand U7099 (N_7099,N_5965,N_5875);
xor U7100 (N_7100,N_6342,N_6385);
xnor U7101 (N_7101,N_5761,N_6161);
and U7102 (N_7102,N_5802,N_5699);
and U7103 (N_7103,N_5668,N_5683);
xor U7104 (N_7104,N_5943,N_6094);
xnor U7105 (N_7105,N_6090,N_5834);
or U7106 (N_7106,N_6102,N_6157);
nor U7107 (N_7107,N_6382,N_5947);
xnor U7108 (N_7108,N_5628,N_5929);
xor U7109 (N_7109,N_6126,N_6047);
xor U7110 (N_7110,N_6180,N_5693);
nand U7111 (N_7111,N_5892,N_5707);
nand U7112 (N_7112,N_5981,N_5719);
and U7113 (N_7113,N_6102,N_6012);
nor U7114 (N_7114,N_5848,N_6135);
nor U7115 (N_7115,N_6042,N_6184);
nand U7116 (N_7116,N_5667,N_6355);
nand U7117 (N_7117,N_5961,N_6222);
nor U7118 (N_7118,N_6250,N_5768);
nor U7119 (N_7119,N_5991,N_6053);
xnor U7120 (N_7120,N_5992,N_5895);
and U7121 (N_7121,N_6312,N_5822);
nand U7122 (N_7122,N_5707,N_5960);
nor U7123 (N_7123,N_5724,N_5829);
xnor U7124 (N_7124,N_5917,N_6062);
and U7125 (N_7125,N_6322,N_6343);
and U7126 (N_7126,N_5677,N_5645);
or U7127 (N_7127,N_5773,N_6276);
and U7128 (N_7128,N_6339,N_5687);
and U7129 (N_7129,N_6359,N_6386);
nor U7130 (N_7130,N_6232,N_5945);
or U7131 (N_7131,N_5891,N_6323);
nor U7132 (N_7132,N_6049,N_6011);
and U7133 (N_7133,N_5969,N_6077);
and U7134 (N_7134,N_5756,N_5848);
xnor U7135 (N_7135,N_6103,N_6291);
nand U7136 (N_7136,N_6218,N_6267);
xor U7137 (N_7137,N_6121,N_6298);
xnor U7138 (N_7138,N_5844,N_5630);
nor U7139 (N_7139,N_6034,N_6245);
nor U7140 (N_7140,N_5695,N_5754);
nor U7141 (N_7141,N_5892,N_6012);
and U7142 (N_7142,N_6049,N_6315);
nor U7143 (N_7143,N_5664,N_6133);
nand U7144 (N_7144,N_6033,N_5634);
xor U7145 (N_7145,N_5751,N_6273);
nand U7146 (N_7146,N_6382,N_5718);
xnor U7147 (N_7147,N_5935,N_6026);
nand U7148 (N_7148,N_5721,N_5696);
nor U7149 (N_7149,N_5761,N_6175);
xor U7150 (N_7150,N_5755,N_6166);
or U7151 (N_7151,N_6376,N_6317);
and U7152 (N_7152,N_5789,N_6244);
nor U7153 (N_7153,N_5977,N_6384);
nor U7154 (N_7154,N_5731,N_5681);
xor U7155 (N_7155,N_5848,N_5793);
or U7156 (N_7156,N_5825,N_5894);
nor U7157 (N_7157,N_6242,N_6024);
nor U7158 (N_7158,N_6223,N_5886);
and U7159 (N_7159,N_5830,N_6357);
nand U7160 (N_7160,N_5800,N_5682);
or U7161 (N_7161,N_6197,N_6396);
and U7162 (N_7162,N_5825,N_5829);
xor U7163 (N_7163,N_5792,N_5889);
and U7164 (N_7164,N_6050,N_6309);
nor U7165 (N_7165,N_5665,N_6383);
and U7166 (N_7166,N_5806,N_6002);
nand U7167 (N_7167,N_6049,N_6072);
xnor U7168 (N_7168,N_5993,N_5858);
or U7169 (N_7169,N_6256,N_5738);
nor U7170 (N_7170,N_6338,N_6091);
nor U7171 (N_7171,N_5670,N_6316);
xnor U7172 (N_7172,N_5623,N_5942);
nor U7173 (N_7173,N_6316,N_6212);
or U7174 (N_7174,N_6350,N_5826);
nor U7175 (N_7175,N_6110,N_6023);
nor U7176 (N_7176,N_6225,N_6230);
nor U7177 (N_7177,N_5735,N_6010);
nand U7178 (N_7178,N_5879,N_5844);
nor U7179 (N_7179,N_5878,N_5962);
or U7180 (N_7180,N_6118,N_5783);
nor U7181 (N_7181,N_6010,N_6319);
or U7182 (N_7182,N_6077,N_5885);
nand U7183 (N_7183,N_5735,N_5749);
xnor U7184 (N_7184,N_5735,N_5722);
and U7185 (N_7185,N_6297,N_6343);
nand U7186 (N_7186,N_5808,N_6000);
nor U7187 (N_7187,N_5627,N_6064);
xnor U7188 (N_7188,N_6110,N_5632);
and U7189 (N_7189,N_5815,N_6028);
and U7190 (N_7190,N_5678,N_6301);
nand U7191 (N_7191,N_6080,N_6179);
and U7192 (N_7192,N_6318,N_6381);
and U7193 (N_7193,N_5702,N_5856);
and U7194 (N_7194,N_5673,N_6280);
nand U7195 (N_7195,N_5673,N_5934);
xor U7196 (N_7196,N_5871,N_5710);
nand U7197 (N_7197,N_5660,N_6096);
or U7198 (N_7198,N_6080,N_6030);
nor U7199 (N_7199,N_6222,N_6268);
xor U7200 (N_7200,N_7135,N_6602);
xor U7201 (N_7201,N_7120,N_6554);
nor U7202 (N_7202,N_6785,N_6679);
nor U7203 (N_7203,N_6509,N_6504);
nand U7204 (N_7204,N_6609,N_6889);
and U7205 (N_7205,N_6810,N_6695);
nand U7206 (N_7206,N_6674,N_6986);
xnor U7207 (N_7207,N_7102,N_6790);
or U7208 (N_7208,N_7137,N_6576);
xnor U7209 (N_7209,N_6783,N_6590);
nand U7210 (N_7210,N_7163,N_7042);
or U7211 (N_7211,N_6687,N_6725);
xor U7212 (N_7212,N_6424,N_6714);
or U7213 (N_7213,N_6622,N_6982);
and U7214 (N_7214,N_6448,N_6910);
nand U7215 (N_7215,N_7124,N_6870);
nand U7216 (N_7216,N_7062,N_7174);
nand U7217 (N_7217,N_6949,N_6856);
nand U7218 (N_7218,N_6902,N_7103);
nand U7219 (N_7219,N_6670,N_6942);
or U7220 (N_7220,N_6914,N_6897);
nor U7221 (N_7221,N_6626,N_7067);
nand U7222 (N_7222,N_7015,N_6850);
xor U7223 (N_7223,N_6467,N_6698);
nand U7224 (N_7224,N_6427,N_6820);
or U7225 (N_7225,N_6945,N_6912);
or U7226 (N_7226,N_6849,N_7101);
nand U7227 (N_7227,N_6441,N_6432);
or U7228 (N_7228,N_6979,N_6722);
xor U7229 (N_7229,N_7131,N_6781);
nor U7230 (N_7230,N_6573,N_6552);
and U7231 (N_7231,N_6638,N_7122);
or U7232 (N_7232,N_7006,N_6676);
nand U7233 (N_7233,N_6831,N_6694);
xor U7234 (N_7234,N_7087,N_6458);
or U7235 (N_7235,N_7050,N_6641);
and U7236 (N_7236,N_7011,N_6519);
nand U7237 (N_7237,N_6705,N_6579);
nor U7238 (N_7238,N_7021,N_6888);
nor U7239 (N_7239,N_6619,N_6816);
xnor U7240 (N_7240,N_6656,N_7108);
xnor U7241 (N_7241,N_6433,N_6672);
nor U7242 (N_7242,N_6689,N_7090);
nor U7243 (N_7243,N_6992,N_6791);
and U7244 (N_7244,N_6913,N_6421);
nor U7245 (N_7245,N_6699,N_6898);
xnor U7246 (N_7246,N_6815,N_6978);
or U7247 (N_7247,N_6911,N_7180);
and U7248 (N_7248,N_6776,N_6900);
xnor U7249 (N_7249,N_6806,N_6630);
nor U7250 (N_7250,N_6955,N_7002);
and U7251 (N_7251,N_6866,N_6901);
nor U7252 (N_7252,N_6419,N_6952);
xor U7253 (N_7253,N_7127,N_6594);
or U7254 (N_7254,N_6644,N_6526);
nor U7255 (N_7255,N_6530,N_6539);
nand U7256 (N_7256,N_6971,N_6643);
and U7257 (N_7257,N_6586,N_6498);
or U7258 (N_7258,N_6628,N_6686);
or U7259 (N_7259,N_7004,N_6891);
xnor U7260 (N_7260,N_6682,N_7094);
nor U7261 (N_7261,N_7194,N_6566);
xnor U7262 (N_7262,N_7162,N_6511);
or U7263 (N_7263,N_7008,N_6425);
xnor U7264 (N_7264,N_6871,N_6770);
nand U7265 (N_7265,N_6549,N_6943);
xor U7266 (N_7266,N_6933,N_6924);
nand U7267 (N_7267,N_7121,N_6751);
nand U7268 (N_7268,N_6516,N_7029);
or U7269 (N_7269,N_6431,N_6998);
nand U7270 (N_7270,N_6488,N_6972);
or U7271 (N_7271,N_6729,N_6771);
xnor U7272 (N_7272,N_6652,N_6838);
or U7273 (N_7273,N_7084,N_6975);
nor U7274 (N_7274,N_7145,N_7000);
nand U7275 (N_7275,N_6983,N_6525);
and U7276 (N_7276,N_7199,N_6589);
nand U7277 (N_7277,N_6520,N_6451);
xnor U7278 (N_7278,N_6565,N_6953);
and U7279 (N_7279,N_6449,N_7188);
nor U7280 (N_7280,N_7155,N_6627);
nand U7281 (N_7281,N_6747,N_6648);
or U7282 (N_7282,N_6446,N_6673);
and U7283 (N_7283,N_7097,N_7088);
nand U7284 (N_7284,N_7117,N_7140);
xnor U7285 (N_7285,N_6854,N_6802);
and U7286 (N_7286,N_6919,N_6957);
or U7287 (N_7287,N_6769,N_6584);
or U7288 (N_7288,N_6477,N_6890);
or U7289 (N_7289,N_7093,N_6631);
or U7290 (N_7290,N_7078,N_6796);
xor U7291 (N_7291,N_6855,N_6593);
nand U7292 (N_7292,N_6462,N_6899);
xor U7293 (N_7293,N_7092,N_6437);
and U7294 (N_7294,N_6809,N_7081);
and U7295 (N_7295,N_6755,N_6574);
or U7296 (N_7296,N_6610,N_6859);
or U7297 (N_7297,N_7023,N_6683);
nor U7298 (N_7298,N_7129,N_7100);
nor U7299 (N_7299,N_6882,N_6531);
nor U7300 (N_7300,N_7056,N_6829);
and U7301 (N_7301,N_6731,N_6591);
nor U7302 (N_7302,N_6614,N_6968);
or U7303 (N_7303,N_6557,N_7107);
and U7304 (N_7304,N_6487,N_6981);
xnor U7305 (N_7305,N_7150,N_6719);
or U7306 (N_7306,N_6764,N_6438);
nor U7307 (N_7307,N_6495,N_6455);
or U7308 (N_7308,N_6839,N_6443);
or U7309 (N_7309,N_7045,N_6570);
nand U7310 (N_7310,N_6478,N_7171);
and U7311 (N_7311,N_6693,N_7172);
nand U7312 (N_7312,N_6469,N_6601);
nand U7313 (N_7313,N_7071,N_6988);
nand U7314 (N_7314,N_6550,N_6775);
or U7315 (N_7315,N_6744,N_6896);
and U7316 (N_7316,N_6788,N_6606);
nand U7317 (N_7317,N_7133,N_6993);
nand U7318 (N_7318,N_7060,N_6440);
nor U7319 (N_7319,N_7178,N_6886);
xnor U7320 (N_7320,N_6822,N_6517);
nand U7321 (N_7321,N_6647,N_6843);
nand U7322 (N_7322,N_6653,N_6658);
nand U7323 (N_7323,N_6476,N_6585);
and U7324 (N_7324,N_6887,N_6436);
xor U7325 (N_7325,N_7123,N_6401);
or U7326 (N_7326,N_7086,N_6869);
or U7327 (N_7327,N_6501,N_6807);
nand U7328 (N_7328,N_6941,N_6571);
and U7329 (N_7329,N_6926,N_6999);
xnor U7330 (N_7330,N_6551,N_6684);
xnor U7331 (N_7331,N_6966,N_6713);
and U7332 (N_7332,N_6546,N_6750);
nand U7333 (N_7333,N_6406,N_7195);
xor U7334 (N_7334,N_6749,N_6878);
nand U7335 (N_7335,N_6930,N_7099);
or U7336 (N_7336,N_6580,N_6489);
or U7337 (N_7337,N_7080,N_6515);
nand U7338 (N_7338,N_7198,N_6618);
nand U7339 (N_7339,N_6490,N_6651);
and U7340 (N_7340,N_6721,N_6603);
nand U7341 (N_7341,N_6703,N_6430);
nor U7342 (N_7342,N_7096,N_7152);
and U7343 (N_7343,N_7168,N_6474);
nand U7344 (N_7344,N_7055,N_6928);
and U7345 (N_7345,N_7109,N_6667);
or U7346 (N_7346,N_7095,N_7089);
or U7347 (N_7347,N_7106,N_6600);
nand U7348 (N_7348,N_6834,N_6905);
and U7349 (N_7349,N_7061,N_6454);
nor U7350 (N_7350,N_6632,N_7065);
xor U7351 (N_7351,N_7113,N_6872);
xor U7352 (N_7352,N_6918,N_7032);
xnor U7353 (N_7353,N_6464,N_6865);
and U7354 (N_7354,N_6635,N_6857);
nor U7355 (N_7355,N_6528,N_6678);
and U7356 (N_7356,N_6756,N_6403);
nor U7357 (N_7357,N_6964,N_6768);
and U7358 (N_7358,N_6450,N_6581);
and U7359 (N_7359,N_7037,N_7085);
and U7360 (N_7360,N_6936,N_6852);
or U7361 (N_7361,N_6418,N_7098);
or U7362 (N_7362,N_6479,N_6492);
or U7363 (N_7363,N_6720,N_6496);
nor U7364 (N_7364,N_6588,N_7105);
and U7365 (N_7365,N_6502,N_7186);
nand U7366 (N_7366,N_6757,N_6938);
or U7367 (N_7367,N_6961,N_6533);
nor U7368 (N_7368,N_6792,N_6409);
nor U7369 (N_7369,N_6818,N_7010);
and U7370 (N_7370,N_7057,N_6700);
nor U7371 (N_7371,N_7143,N_6803);
nand U7372 (N_7372,N_6841,N_6794);
nand U7373 (N_7373,N_7136,N_7160);
nand U7374 (N_7374,N_6860,N_6471);
nand U7375 (N_7375,N_7158,N_6445);
or U7376 (N_7376,N_6962,N_6759);
nor U7377 (N_7377,N_6877,N_6762);
xnor U7378 (N_7378,N_7020,N_6814);
nor U7379 (N_7379,N_7130,N_7068);
nand U7380 (N_7380,N_7049,N_6639);
nor U7381 (N_7381,N_7069,N_7157);
or U7382 (N_7382,N_6547,N_6944);
nand U7383 (N_7383,N_6697,N_6895);
and U7384 (N_7384,N_6795,N_6510);
nor U7385 (N_7385,N_6428,N_6948);
nor U7386 (N_7386,N_6407,N_6553);
or U7387 (N_7387,N_6696,N_7059);
nor U7388 (N_7388,N_7118,N_6845);
xnor U7389 (N_7389,N_6706,N_6991);
or U7390 (N_7390,N_6710,N_6715);
nor U7391 (N_7391,N_6408,N_6485);
nor U7392 (N_7392,N_7116,N_7063);
or U7393 (N_7393,N_6457,N_7189);
nand U7394 (N_7394,N_6723,N_6774);
and U7395 (N_7395,N_7058,N_6666);
nor U7396 (N_7396,N_6808,N_7017);
nor U7397 (N_7397,N_6415,N_7119);
and U7398 (N_7398,N_6650,N_6688);
or U7399 (N_7399,N_6567,N_7161);
xnor U7400 (N_7400,N_6417,N_6738);
or U7401 (N_7401,N_7142,N_6939);
nand U7402 (N_7402,N_7079,N_7024);
nor U7403 (N_7403,N_6671,N_6481);
nor U7404 (N_7404,N_6654,N_6691);
nor U7405 (N_7405,N_7076,N_7134);
or U7406 (N_7406,N_6578,N_6904);
and U7407 (N_7407,N_6617,N_6486);
and U7408 (N_7408,N_7104,N_7064);
or U7409 (N_7409,N_6465,N_6737);
and U7410 (N_7410,N_6611,N_7165);
or U7411 (N_7411,N_7190,N_6534);
or U7412 (N_7412,N_6420,N_6642);
nor U7413 (N_7413,N_6535,N_6836);
or U7414 (N_7414,N_6956,N_6784);
and U7415 (N_7415,N_7030,N_6995);
and U7416 (N_7416,N_6548,N_6493);
nor U7417 (N_7417,N_6506,N_7052);
nor U7418 (N_7418,N_6412,N_6921);
nand U7419 (N_7419,N_6940,N_6799);
xnor U7420 (N_7420,N_6655,N_7192);
xor U7421 (N_7421,N_6825,N_7125);
xor U7422 (N_7422,N_6793,N_6704);
xnor U7423 (N_7423,N_6976,N_6616);
nor U7424 (N_7424,N_6463,N_6996);
or U7425 (N_7425,N_7014,N_6660);
or U7426 (N_7426,N_6801,N_6435);
xnor U7427 (N_7427,N_6447,N_7183);
xor U7428 (N_7428,N_7151,N_7025);
xor U7429 (N_7429,N_6532,N_6935);
or U7430 (N_7430,N_6634,N_6572);
nor U7431 (N_7431,N_7016,N_6819);
or U7432 (N_7432,N_6665,N_6442);
and U7433 (N_7433,N_6766,N_7147);
nand U7434 (N_7434,N_6649,N_6633);
xor U7435 (N_7435,N_6527,N_7187);
nor U7436 (N_7436,N_6742,N_6405);
nor U7437 (N_7437,N_7177,N_7040);
nor U7438 (N_7438,N_6541,N_7046);
or U7439 (N_7439,N_6536,N_6592);
xor U7440 (N_7440,N_6482,N_7139);
and U7441 (N_7441,N_6508,N_7003);
and U7442 (N_7442,N_6568,N_7031);
xnor U7443 (N_7443,N_6669,N_7193);
nand U7444 (N_7444,N_6922,N_7156);
xor U7445 (N_7445,N_6514,N_6543);
nor U7446 (N_7446,N_6597,N_6797);
nand U7447 (N_7447,N_6959,N_6640);
nand U7448 (N_7448,N_7012,N_6934);
nand U7449 (N_7449,N_7027,N_7184);
or U7450 (N_7450,N_7054,N_6545);
and U7451 (N_7451,N_6734,N_6804);
and U7452 (N_7452,N_6690,N_6861);
xor U7453 (N_7453,N_6800,N_7026);
nor U7454 (N_7454,N_6522,N_6411);
and U7455 (N_7455,N_6468,N_6805);
nor U7456 (N_7456,N_6620,N_6717);
and U7457 (N_7457,N_6858,N_6880);
or U7458 (N_7458,N_6472,N_7005);
or U7459 (N_7459,N_6821,N_7181);
xnor U7460 (N_7460,N_6484,N_6833);
or U7461 (N_7461,N_6772,N_6937);
or U7462 (N_7462,N_6613,N_6728);
or U7463 (N_7463,N_6743,N_6452);
nor U7464 (N_7464,N_6960,N_7036);
and U7465 (N_7465,N_7082,N_6973);
xor U7466 (N_7466,N_6980,N_6503);
or U7467 (N_7467,N_6400,N_7144);
or U7468 (N_7468,N_6416,N_6916);
xor U7469 (N_7469,N_7182,N_6414);
nor U7470 (N_7470,N_6513,N_6760);
nor U7471 (N_7471,N_6677,N_6863);
xnor U7472 (N_7472,N_6518,N_6475);
and U7473 (N_7473,N_6680,N_6827);
or U7474 (N_7474,N_6466,N_7044);
or U7475 (N_7475,N_6681,N_6538);
nand U7476 (N_7476,N_6851,N_6608);
and U7477 (N_7477,N_6524,N_7018);
nor U7478 (N_7478,N_7175,N_7009);
nor U7479 (N_7479,N_6661,N_6997);
xnor U7480 (N_7480,N_6732,N_6473);
nand U7481 (N_7481,N_6542,N_6842);
nor U7482 (N_7482,N_7028,N_6577);
and U7483 (N_7483,N_6925,N_7007);
nor U7484 (N_7484,N_6958,N_6663);
nor U7485 (N_7485,N_6657,N_6830);
nand U7486 (N_7486,N_7166,N_6929);
nor U7487 (N_7487,N_6736,N_6582);
nand U7488 (N_7488,N_6894,N_7170);
and U7489 (N_7489,N_6823,N_6664);
or U7490 (N_7490,N_6779,N_6828);
nor U7491 (N_7491,N_6716,N_6599);
nand U7492 (N_7492,N_6873,N_6817);
nand U7493 (N_7493,N_6583,N_6556);
or U7494 (N_7494,N_7074,N_6727);
and U7495 (N_7495,N_6753,N_7075);
xor U7496 (N_7496,N_7149,N_6844);
nand U7497 (N_7497,N_7043,N_6562);
nor U7498 (N_7498,N_6946,N_7091);
and U7499 (N_7499,N_6702,N_6868);
xnor U7500 (N_7500,N_6621,N_6423);
xnor U7501 (N_7501,N_6470,N_6625);
nor U7502 (N_7502,N_6444,N_6637);
or U7503 (N_7503,N_7039,N_7141);
nor U7504 (N_7504,N_6846,N_6712);
nand U7505 (N_7505,N_6607,N_6777);
nor U7506 (N_7506,N_7191,N_6947);
nor U7507 (N_7507,N_6811,N_6984);
nor U7508 (N_7508,N_6954,N_6500);
and U7509 (N_7509,N_6410,N_6909);
nand U7510 (N_7510,N_6950,N_6835);
and U7511 (N_7511,N_6969,N_6453);
or U7512 (N_7512,N_6864,N_6615);
and U7513 (N_7513,N_6512,N_6733);
nor U7514 (N_7514,N_6707,N_7173);
nand U7515 (N_7515,N_6605,N_6917);
and U7516 (N_7516,N_6951,N_6701);
nand U7517 (N_7517,N_6529,N_6558);
or U7518 (N_7518,N_6885,N_7167);
and U7519 (N_7519,N_6903,N_6708);
xor U7520 (N_7520,N_6711,N_7019);
nand U7521 (N_7521,N_7048,N_6659);
xor U7522 (N_7522,N_6848,N_6507);
xnor U7523 (N_7523,N_6499,N_6985);
nor U7524 (N_7524,N_6879,N_6763);
xnor U7525 (N_7525,N_6853,N_6675);
nand U7526 (N_7526,N_6624,N_6994);
nor U7527 (N_7527,N_7138,N_6746);
nand U7528 (N_7528,N_6847,N_7022);
and U7529 (N_7529,N_6813,N_7053);
or U7530 (N_7530,N_6739,N_6990);
nor U7531 (N_7531,N_7013,N_7153);
nor U7532 (N_7532,N_6460,N_7035);
xnor U7533 (N_7533,N_6989,N_6559);
xnor U7534 (N_7534,N_6977,N_6881);
and U7535 (N_7535,N_6561,N_7001);
nand U7536 (N_7536,N_6596,N_6569);
nor U7537 (N_7537,N_7041,N_6461);
xor U7538 (N_7538,N_6718,N_6780);
or U7539 (N_7539,N_7176,N_6812);
nor U7540 (N_7540,N_6646,N_6893);
and U7541 (N_7541,N_6402,N_6798);
xor U7542 (N_7542,N_6892,N_7128);
and U7543 (N_7543,N_7077,N_6505);
nand U7544 (N_7544,N_6726,N_6965);
nor U7545 (N_7545,N_6970,N_6884);
or U7546 (N_7546,N_6587,N_7073);
nand U7547 (N_7547,N_6752,N_6563);
and U7548 (N_7548,N_6459,N_6429);
and U7549 (N_7549,N_6920,N_6786);
nand U7550 (N_7550,N_6604,N_6741);
nand U7551 (N_7551,N_6623,N_6497);
xor U7552 (N_7552,N_6483,N_7169);
xor U7553 (N_7553,N_6906,N_6837);
nor U7554 (N_7554,N_6840,N_7146);
nand U7555 (N_7555,N_6876,N_6537);
and U7556 (N_7556,N_7197,N_6778);
nor U7557 (N_7557,N_6575,N_6662);
and U7558 (N_7558,N_7051,N_7034);
nand U7559 (N_7559,N_6434,N_7033);
and U7560 (N_7560,N_6636,N_6521);
and U7561 (N_7561,N_6832,N_6974);
or U7562 (N_7562,N_6745,N_7148);
nor U7563 (N_7563,N_6422,N_6404);
xor U7564 (N_7564,N_6724,N_6426);
nor U7565 (N_7565,N_6782,N_6685);
or U7566 (N_7566,N_6787,N_7047);
xnor U7567 (N_7567,N_6915,N_6564);
nand U7568 (N_7568,N_7112,N_6555);
nand U7569 (N_7569,N_7164,N_6773);
or U7570 (N_7570,N_6544,N_6540);
xor U7571 (N_7571,N_6908,N_6612);
and U7572 (N_7572,N_6560,N_7110);
and U7573 (N_7573,N_7072,N_6413);
xor U7574 (N_7574,N_6761,N_6862);
and U7575 (N_7575,N_6765,N_6730);
xnor U7576 (N_7576,N_6963,N_6754);
nand U7577 (N_7577,N_6874,N_6867);
and U7578 (N_7578,N_7185,N_6709);
and U7579 (N_7579,N_6883,N_7126);
and U7580 (N_7580,N_7038,N_6456);
and U7581 (N_7581,N_6826,N_6740);
or U7582 (N_7582,N_6629,N_7114);
and U7583 (N_7583,N_6932,N_7083);
or U7584 (N_7584,N_7111,N_7070);
nand U7585 (N_7585,N_6645,N_7179);
nand U7586 (N_7586,N_6987,N_6927);
xor U7587 (N_7587,N_6923,N_6907);
xnor U7588 (N_7588,N_6598,N_7159);
xnor U7589 (N_7589,N_7115,N_6735);
or U7590 (N_7590,N_6439,N_6789);
and U7591 (N_7591,N_6595,N_7196);
and U7592 (N_7592,N_6748,N_6668);
xor U7593 (N_7593,N_6875,N_6767);
xnor U7594 (N_7594,N_6491,N_6523);
nor U7595 (N_7595,N_7132,N_7154);
nor U7596 (N_7596,N_6758,N_6480);
nand U7597 (N_7597,N_6692,N_6931);
nand U7598 (N_7598,N_7066,N_6494);
or U7599 (N_7599,N_6824,N_6967);
nor U7600 (N_7600,N_6894,N_7004);
xnor U7601 (N_7601,N_6898,N_7074);
nor U7602 (N_7602,N_6514,N_7031);
xor U7603 (N_7603,N_6449,N_6898);
and U7604 (N_7604,N_6702,N_6941);
nor U7605 (N_7605,N_6820,N_6782);
and U7606 (N_7606,N_6916,N_6419);
nand U7607 (N_7607,N_7149,N_6882);
xnor U7608 (N_7608,N_6634,N_6509);
nand U7609 (N_7609,N_7168,N_6958);
nand U7610 (N_7610,N_6912,N_6618);
xnor U7611 (N_7611,N_6801,N_7047);
xor U7612 (N_7612,N_6478,N_7193);
xor U7613 (N_7613,N_6849,N_7088);
and U7614 (N_7614,N_6907,N_6960);
or U7615 (N_7615,N_6587,N_6598);
nand U7616 (N_7616,N_6528,N_7167);
xnor U7617 (N_7617,N_6485,N_7165);
or U7618 (N_7618,N_7097,N_6571);
nand U7619 (N_7619,N_6808,N_7182);
and U7620 (N_7620,N_6899,N_6686);
xor U7621 (N_7621,N_6945,N_6603);
nor U7622 (N_7622,N_6488,N_6825);
and U7623 (N_7623,N_6723,N_6480);
and U7624 (N_7624,N_7071,N_6532);
nor U7625 (N_7625,N_6711,N_6759);
nand U7626 (N_7626,N_6444,N_7151);
nor U7627 (N_7627,N_6685,N_7074);
nor U7628 (N_7628,N_7036,N_6542);
and U7629 (N_7629,N_6993,N_7190);
and U7630 (N_7630,N_7181,N_7034);
nand U7631 (N_7631,N_6715,N_6858);
xnor U7632 (N_7632,N_6715,N_6641);
and U7633 (N_7633,N_6690,N_6421);
nand U7634 (N_7634,N_6583,N_7196);
xnor U7635 (N_7635,N_6664,N_6786);
nor U7636 (N_7636,N_6476,N_7018);
xor U7637 (N_7637,N_6856,N_6902);
or U7638 (N_7638,N_6554,N_6857);
or U7639 (N_7639,N_6842,N_7016);
and U7640 (N_7640,N_6639,N_6675);
and U7641 (N_7641,N_6543,N_6525);
and U7642 (N_7642,N_6534,N_6980);
nor U7643 (N_7643,N_6595,N_6694);
and U7644 (N_7644,N_6979,N_6933);
nor U7645 (N_7645,N_6550,N_6517);
xnor U7646 (N_7646,N_7141,N_6643);
nand U7647 (N_7647,N_6879,N_6922);
nand U7648 (N_7648,N_6569,N_6787);
xnor U7649 (N_7649,N_6424,N_6882);
nor U7650 (N_7650,N_6596,N_7118);
nand U7651 (N_7651,N_6642,N_6428);
nand U7652 (N_7652,N_7096,N_6579);
or U7653 (N_7653,N_6739,N_6917);
or U7654 (N_7654,N_6536,N_6930);
and U7655 (N_7655,N_6714,N_6515);
nor U7656 (N_7656,N_6859,N_7006);
nor U7657 (N_7657,N_6665,N_6712);
nand U7658 (N_7658,N_6837,N_6502);
nor U7659 (N_7659,N_6470,N_7141);
and U7660 (N_7660,N_7013,N_7146);
nand U7661 (N_7661,N_7003,N_6817);
or U7662 (N_7662,N_6972,N_6915);
xor U7663 (N_7663,N_6406,N_7193);
xnor U7664 (N_7664,N_6794,N_7155);
nand U7665 (N_7665,N_7002,N_7052);
xnor U7666 (N_7666,N_7071,N_6769);
nand U7667 (N_7667,N_6452,N_6760);
and U7668 (N_7668,N_7102,N_6728);
nor U7669 (N_7669,N_6982,N_6666);
and U7670 (N_7670,N_7098,N_6513);
or U7671 (N_7671,N_7132,N_7110);
nand U7672 (N_7672,N_6639,N_6502);
and U7673 (N_7673,N_6691,N_6945);
or U7674 (N_7674,N_6508,N_6830);
nand U7675 (N_7675,N_6683,N_6751);
nand U7676 (N_7676,N_6724,N_6943);
and U7677 (N_7677,N_6864,N_7061);
or U7678 (N_7678,N_7007,N_6887);
nand U7679 (N_7679,N_6880,N_7050);
or U7680 (N_7680,N_6745,N_6832);
and U7681 (N_7681,N_6995,N_6466);
or U7682 (N_7682,N_6745,N_6655);
nand U7683 (N_7683,N_7114,N_6964);
nand U7684 (N_7684,N_6686,N_6599);
or U7685 (N_7685,N_6411,N_6628);
nor U7686 (N_7686,N_6537,N_6803);
nor U7687 (N_7687,N_6418,N_7070);
nor U7688 (N_7688,N_6977,N_6441);
nor U7689 (N_7689,N_7132,N_6813);
xor U7690 (N_7690,N_7046,N_6588);
nor U7691 (N_7691,N_6599,N_6493);
and U7692 (N_7692,N_6467,N_7056);
nand U7693 (N_7693,N_7199,N_6537);
and U7694 (N_7694,N_7025,N_6998);
or U7695 (N_7695,N_6484,N_6853);
or U7696 (N_7696,N_6714,N_6530);
or U7697 (N_7697,N_6504,N_6670);
nand U7698 (N_7698,N_6887,N_6971);
nor U7699 (N_7699,N_6831,N_6907);
nand U7700 (N_7700,N_6471,N_6925);
nor U7701 (N_7701,N_6505,N_6653);
xnor U7702 (N_7702,N_7034,N_6969);
nor U7703 (N_7703,N_6659,N_6831);
nand U7704 (N_7704,N_7181,N_6670);
and U7705 (N_7705,N_7105,N_7066);
and U7706 (N_7706,N_6565,N_7177);
nand U7707 (N_7707,N_7064,N_6720);
xnor U7708 (N_7708,N_6447,N_6455);
or U7709 (N_7709,N_6778,N_6468);
nand U7710 (N_7710,N_6452,N_7148);
xnor U7711 (N_7711,N_6611,N_7056);
xor U7712 (N_7712,N_6732,N_7057);
nand U7713 (N_7713,N_6783,N_7056);
xnor U7714 (N_7714,N_6779,N_7075);
nor U7715 (N_7715,N_6678,N_6650);
and U7716 (N_7716,N_6732,N_6805);
xnor U7717 (N_7717,N_6416,N_6439);
and U7718 (N_7718,N_6981,N_6709);
or U7719 (N_7719,N_6846,N_6457);
nand U7720 (N_7720,N_6480,N_6557);
xor U7721 (N_7721,N_7052,N_6735);
xnor U7722 (N_7722,N_6622,N_7001);
xnor U7723 (N_7723,N_6795,N_6937);
nor U7724 (N_7724,N_6452,N_6861);
or U7725 (N_7725,N_7091,N_6544);
nor U7726 (N_7726,N_6650,N_6658);
and U7727 (N_7727,N_6889,N_6792);
nor U7728 (N_7728,N_6908,N_6896);
or U7729 (N_7729,N_6504,N_6989);
xor U7730 (N_7730,N_6916,N_6989);
nor U7731 (N_7731,N_6742,N_6955);
and U7732 (N_7732,N_6925,N_6626);
or U7733 (N_7733,N_7161,N_6415);
nand U7734 (N_7734,N_6584,N_7108);
nor U7735 (N_7735,N_7006,N_6443);
nor U7736 (N_7736,N_6789,N_6412);
and U7737 (N_7737,N_6917,N_7076);
nand U7738 (N_7738,N_6872,N_7075);
xor U7739 (N_7739,N_7069,N_6977);
and U7740 (N_7740,N_7051,N_6763);
nand U7741 (N_7741,N_6992,N_6909);
nand U7742 (N_7742,N_6694,N_7075);
xnor U7743 (N_7743,N_6779,N_6683);
nand U7744 (N_7744,N_7115,N_7172);
and U7745 (N_7745,N_7136,N_6690);
or U7746 (N_7746,N_7088,N_6931);
xnor U7747 (N_7747,N_6835,N_6441);
xor U7748 (N_7748,N_6450,N_6652);
xnor U7749 (N_7749,N_7135,N_6476);
xor U7750 (N_7750,N_6556,N_6802);
or U7751 (N_7751,N_7078,N_7190);
nor U7752 (N_7752,N_6817,N_6891);
xnor U7753 (N_7753,N_6904,N_7040);
nor U7754 (N_7754,N_6948,N_6417);
xnor U7755 (N_7755,N_6860,N_6957);
nand U7756 (N_7756,N_7091,N_6670);
nand U7757 (N_7757,N_6853,N_7044);
nand U7758 (N_7758,N_6885,N_6710);
nor U7759 (N_7759,N_6660,N_6509);
xor U7760 (N_7760,N_6588,N_6986);
nor U7761 (N_7761,N_7060,N_6695);
xnor U7762 (N_7762,N_6892,N_6504);
and U7763 (N_7763,N_6590,N_7099);
and U7764 (N_7764,N_6737,N_6545);
xnor U7765 (N_7765,N_6677,N_6533);
nand U7766 (N_7766,N_6817,N_7067);
or U7767 (N_7767,N_6716,N_6961);
nand U7768 (N_7768,N_7146,N_6945);
xor U7769 (N_7769,N_6790,N_6812);
or U7770 (N_7770,N_6930,N_6416);
xor U7771 (N_7771,N_6845,N_6948);
or U7772 (N_7772,N_6442,N_7101);
nor U7773 (N_7773,N_7180,N_6918);
nor U7774 (N_7774,N_6812,N_6806);
nand U7775 (N_7775,N_7158,N_6435);
or U7776 (N_7776,N_6760,N_6403);
nand U7777 (N_7777,N_6707,N_7074);
or U7778 (N_7778,N_7097,N_6448);
nor U7779 (N_7779,N_7080,N_6595);
and U7780 (N_7780,N_6701,N_6408);
nor U7781 (N_7781,N_7012,N_6435);
and U7782 (N_7782,N_6586,N_6985);
nor U7783 (N_7783,N_6571,N_6666);
xor U7784 (N_7784,N_6761,N_7112);
or U7785 (N_7785,N_7158,N_6606);
and U7786 (N_7786,N_6857,N_6692);
or U7787 (N_7787,N_6571,N_6670);
xnor U7788 (N_7788,N_6571,N_6450);
nor U7789 (N_7789,N_6739,N_7106);
nand U7790 (N_7790,N_7161,N_6972);
or U7791 (N_7791,N_7081,N_6531);
nand U7792 (N_7792,N_6647,N_6488);
xor U7793 (N_7793,N_6457,N_6884);
nand U7794 (N_7794,N_6678,N_6681);
xor U7795 (N_7795,N_6745,N_6725);
xor U7796 (N_7796,N_6838,N_6989);
nand U7797 (N_7797,N_6408,N_6760);
and U7798 (N_7798,N_6859,N_6906);
nand U7799 (N_7799,N_6845,N_6651);
or U7800 (N_7800,N_6746,N_7079);
or U7801 (N_7801,N_6736,N_6720);
xor U7802 (N_7802,N_6795,N_6483);
nor U7803 (N_7803,N_6878,N_6562);
xnor U7804 (N_7804,N_6946,N_6556);
or U7805 (N_7805,N_6482,N_6638);
or U7806 (N_7806,N_7146,N_6439);
or U7807 (N_7807,N_6901,N_7102);
xnor U7808 (N_7808,N_7013,N_6802);
nand U7809 (N_7809,N_6935,N_7169);
and U7810 (N_7810,N_6880,N_6966);
and U7811 (N_7811,N_6635,N_6613);
nand U7812 (N_7812,N_6929,N_6806);
and U7813 (N_7813,N_6854,N_6634);
and U7814 (N_7814,N_6547,N_7061);
nand U7815 (N_7815,N_6727,N_7194);
nand U7816 (N_7816,N_6937,N_6800);
xor U7817 (N_7817,N_6699,N_6863);
nor U7818 (N_7818,N_6564,N_6813);
or U7819 (N_7819,N_6528,N_6903);
or U7820 (N_7820,N_6981,N_6747);
and U7821 (N_7821,N_6887,N_6751);
xor U7822 (N_7822,N_7061,N_6878);
nand U7823 (N_7823,N_6834,N_6406);
or U7824 (N_7824,N_6594,N_7178);
nand U7825 (N_7825,N_6559,N_6915);
or U7826 (N_7826,N_6700,N_6794);
xnor U7827 (N_7827,N_6692,N_7120);
nor U7828 (N_7828,N_6943,N_7116);
nand U7829 (N_7829,N_6609,N_7024);
xor U7830 (N_7830,N_6601,N_7190);
and U7831 (N_7831,N_6916,N_6482);
nor U7832 (N_7832,N_6875,N_7081);
xnor U7833 (N_7833,N_7104,N_7058);
nand U7834 (N_7834,N_7157,N_6945);
nand U7835 (N_7835,N_6995,N_6668);
or U7836 (N_7836,N_6728,N_7036);
or U7837 (N_7837,N_6505,N_6788);
nor U7838 (N_7838,N_6783,N_7150);
nor U7839 (N_7839,N_6443,N_6522);
xnor U7840 (N_7840,N_7110,N_6910);
nor U7841 (N_7841,N_6863,N_6903);
xnor U7842 (N_7842,N_6792,N_6993);
nor U7843 (N_7843,N_6428,N_7170);
xor U7844 (N_7844,N_6523,N_6656);
xnor U7845 (N_7845,N_6805,N_6867);
nand U7846 (N_7846,N_7195,N_6777);
or U7847 (N_7847,N_7169,N_6628);
nor U7848 (N_7848,N_6595,N_6525);
nor U7849 (N_7849,N_6549,N_6947);
xor U7850 (N_7850,N_6694,N_6411);
xor U7851 (N_7851,N_7076,N_6465);
nand U7852 (N_7852,N_6602,N_7164);
or U7853 (N_7853,N_6787,N_6560);
xnor U7854 (N_7854,N_7092,N_6990);
nor U7855 (N_7855,N_6775,N_6504);
or U7856 (N_7856,N_6958,N_6473);
or U7857 (N_7857,N_7068,N_7002);
or U7858 (N_7858,N_7116,N_6644);
or U7859 (N_7859,N_6682,N_6753);
nor U7860 (N_7860,N_6454,N_6892);
and U7861 (N_7861,N_6647,N_7177);
nor U7862 (N_7862,N_6921,N_6995);
nand U7863 (N_7863,N_6725,N_6586);
nor U7864 (N_7864,N_6714,N_6776);
nand U7865 (N_7865,N_6724,N_7089);
xor U7866 (N_7866,N_6793,N_7060);
nand U7867 (N_7867,N_7093,N_6685);
nand U7868 (N_7868,N_6711,N_6609);
or U7869 (N_7869,N_6742,N_7008);
or U7870 (N_7870,N_7167,N_6734);
and U7871 (N_7871,N_7187,N_6531);
nand U7872 (N_7872,N_6786,N_6582);
nor U7873 (N_7873,N_6851,N_6978);
nand U7874 (N_7874,N_7075,N_6564);
nor U7875 (N_7875,N_6921,N_6764);
or U7876 (N_7876,N_6524,N_6798);
nor U7877 (N_7877,N_7050,N_6939);
and U7878 (N_7878,N_6659,N_6889);
xnor U7879 (N_7879,N_6801,N_6761);
or U7880 (N_7880,N_7027,N_6812);
and U7881 (N_7881,N_6635,N_7112);
and U7882 (N_7882,N_7056,N_7035);
nor U7883 (N_7883,N_6799,N_6560);
nand U7884 (N_7884,N_6499,N_7143);
and U7885 (N_7885,N_6722,N_6645);
and U7886 (N_7886,N_6675,N_7177);
nor U7887 (N_7887,N_7035,N_6827);
or U7888 (N_7888,N_7190,N_6538);
nand U7889 (N_7889,N_6805,N_6579);
nor U7890 (N_7890,N_6426,N_6834);
or U7891 (N_7891,N_6853,N_6578);
nand U7892 (N_7892,N_6841,N_6783);
xor U7893 (N_7893,N_6806,N_6567);
and U7894 (N_7894,N_6958,N_6785);
nand U7895 (N_7895,N_6606,N_6730);
and U7896 (N_7896,N_6844,N_6917);
xnor U7897 (N_7897,N_7148,N_6932);
nor U7898 (N_7898,N_7155,N_7049);
nand U7899 (N_7899,N_6990,N_6988);
nor U7900 (N_7900,N_6899,N_6789);
or U7901 (N_7901,N_6591,N_6965);
and U7902 (N_7902,N_6652,N_6731);
nor U7903 (N_7903,N_7037,N_6459);
nor U7904 (N_7904,N_6555,N_6850);
or U7905 (N_7905,N_6480,N_6879);
or U7906 (N_7906,N_6601,N_6991);
or U7907 (N_7907,N_6762,N_6716);
or U7908 (N_7908,N_7130,N_6929);
xnor U7909 (N_7909,N_7156,N_6569);
nand U7910 (N_7910,N_6755,N_6461);
nand U7911 (N_7911,N_6540,N_6449);
nand U7912 (N_7912,N_6439,N_7042);
and U7913 (N_7913,N_6865,N_6527);
and U7914 (N_7914,N_6733,N_7031);
nand U7915 (N_7915,N_6814,N_6520);
and U7916 (N_7916,N_7045,N_7157);
xnor U7917 (N_7917,N_7128,N_6645);
xor U7918 (N_7918,N_6824,N_6494);
or U7919 (N_7919,N_6951,N_6774);
nand U7920 (N_7920,N_6510,N_6691);
nand U7921 (N_7921,N_6534,N_7183);
and U7922 (N_7922,N_7021,N_6622);
and U7923 (N_7923,N_6573,N_6553);
xor U7924 (N_7924,N_6721,N_6753);
and U7925 (N_7925,N_6547,N_6590);
nor U7926 (N_7926,N_6654,N_6498);
or U7927 (N_7927,N_6808,N_6667);
nor U7928 (N_7928,N_6417,N_7068);
xnor U7929 (N_7929,N_6589,N_6551);
xor U7930 (N_7930,N_6524,N_6747);
nor U7931 (N_7931,N_6688,N_6485);
and U7932 (N_7932,N_6624,N_6861);
nand U7933 (N_7933,N_6711,N_7054);
xnor U7934 (N_7934,N_6915,N_6529);
or U7935 (N_7935,N_7033,N_6647);
and U7936 (N_7936,N_6617,N_6685);
and U7937 (N_7937,N_6840,N_7093);
nand U7938 (N_7938,N_6576,N_7178);
and U7939 (N_7939,N_7151,N_6913);
and U7940 (N_7940,N_6739,N_6902);
xor U7941 (N_7941,N_6542,N_6707);
or U7942 (N_7942,N_6906,N_6531);
nand U7943 (N_7943,N_6699,N_6745);
or U7944 (N_7944,N_6453,N_6758);
nand U7945 (N_7945,N_6544,N_6416);
nand U7946 (N_7946,N_6716,N_6973);
nor U7947 (N_7947,N_6675,N_6894);
nor U7948 (N_7948,N_6602,N_7154);
nand U7949 (N_7949,N_7029,N_6584);
nand U7950 (N_7950,N_6553,N_7129);
nor U7951 (N_7951,N_6440,N_6736);
or U7952 (N_7952,N_6813,N_6423);
and U7953 (N_7953,N_6662,N_6516);
and U7954 (N_7954,N_6783,N_6719);
and U7955 (N_7955,N_6504,N_6427);
xor U7956 (N_7956,N_6632,N_6602);
and U7957 (N_7957,N_7180,N_6845);
nor U7958 (N_7958,N_6495,N_7080);
and U7959 (N_7959,N_6861,N_6923);
or U7960 (N_7960,N_6421,N_6745);
nor U7961 (N_7961,N_6913,N_7016);
or U7962 (N_7962,N_7103,N_6767);
nand U7963 (N_7963,N_6515,N_6535);
and U7964 (N_7964,N_6551,N_6650);
or U7965 (N_7965,N_6549,N_6908);
nor U7966 (N_7966,N_6491,N_6617);
or U7967 (N_7967,N_6763,N_6725);
and U7968 (N_7968,N_7130,N_6401);
nor U7969 (N_7969,N_6453,N_7192);
nand U7970 (N_7970,N_7074,N_7184);
nor U7971 (N_7971,N_6521,N_6806);
nand U7972 (N_7972,N_7019,N_6992);
and U7973 (N_7973,N_7067,N_7125);
xor U7974 (N_7974,N_6447,N_6878);
xnor U7975 (N_7975,N_6718,N_6442);
and U7976 (N_7976,N_6656,N_7016);
and U7977 (N_7977,N_6875,N_6689);
or U7978 (N_7978,N_6747,N_7156);
or U7979 (N_7979,N_6408,N_6659);
nand U7980 (N_7980,N_6446,N_6556);
or U7981 (N_7981,N_7138,N_6632);
or U7982 (N_7982,N_6755,N_6667);
nand U7983 (N_7983,N_7120,N_6508);
xor U7984 (N_7984,N_6419,N_6462);
nand U7985 (N_7985,N_6768,N_6528);
xnor U7986 (N_7986,N_6421,N_7087);
xor U7987 (N_7987,N_6474,N_6590);
or U7988 (N_7988,N_6953,N_6746);
or U7989 (N_7989,N_6704,N_6900);
nor U7990 (N_7990,N_6866,N_6559);
or U7991 (N_7991,N_7143,N_7107);
and U7992 (N_7992,N_7117,N_6718);
nand U7993 (N_7993,N_6995,N_6577);
nand U7994 (N_7994,N_6465,N_6827);
nor U7995 (N_7995,N_6597,N_6613);
and U7996 (N_7996,N_7159,N_6745);
nand U7997 (N_7997,N_6824,N_6738);
nand U7998 (N_7998,N_6739,N_6685);
and U7999 (N_7999,N_7181,N_6864);
nor U8000 (N_8000,N_7319,N_7241);
or U8001 (N_8001,N_7846,N_7712);
nor U8002 (N_8002,N_7847,N_7737);
xnor U8003 (N_8003,N_7213,N_7885);
nand U8004 (N_8004,N_7332,N_7747);
xor U8005 (N_8005,N_7790,N_7946);
nor U8006 (N_8006,N_7732,N_7326);
xnor U8007 (N_8007,N_7504,N_7797);
or U8008 (N_8008,N_7222,N_7596);
and U8009 (N_8009,N_7677,N_7920);
and U8010 (N_8010,N_7625,N_7698);
nand U8011 (N_8011,N_7774,N_7320);
nand U8012 (N_8012,N_7741,N_7910);
xor U8013 (N_8013,N_7394,N_7526);
xor U8014 (N_8014,N_7338,N_7366);
nand U8015 (N_8015,N_7621,N_7610);
nor U8016 (N_8016,N_7909,N_7735);
and U8017 (N_8017,N_7646,N_7565);
nor U8018 (N_8018,N_7398,N_7551);
and U8019 (N_8019,N_7978,N_7809);
or U8020 (N_8020,N_7449,N_7690);
nor U8021 (N_8021,N_7363,N_7283);
nand U8022 (N_8022,N_7607,N_7364);
or U8023 (N_8023,N_7682,N_7440);
nand U8024 (N_8024,N_7888,N_7863);
nor U8025 (N_8025,N_7611,N_7348);
or U8026 (N_8026,N_7340,N_7518);
xor U8027 (N_8027,N_7490,N_7425);
and U8028 (N_8028,N_7552,N_7753);
nand U8029 (N_8029,N_7403,N_7681);
and U8030 (N_8030,N_7419,N_7255);
nand U8031 (N_8031,N_7870,N_7586);
xnor U8032 (N_8032,N_7520,N_7287);
and U8033 (N_8033,N_7308,N_7852);
and U8034 (N_8034,N_7994,N_7877);
or U8035 (N_8035,N_7421,N_7894);
xor U8036 (N_8036,N_7497,N_7921);
and U8037 (N_8037,N_7208,N_7907);
nand U8038 (N_8038,N_7923,N_7536);
nor U8039 (N_8039,N_7524,N_7715);
nor U8040 (N_8040,N_7508,N_7884);
xor U8041 (N_8041,N_7517,N_7349);
and U8042 (N_8042,N_7236,N_7322);
xor U8043 (N_8043,N_7751,N_7811);
and U8044 (N_8044,N_7861,N_7950);
nor U8045 (N_8045,N_7616,N_7478);
and U8046 (N_8046,N_7396,N_7391);
or U8047 (N_8047,N_7259,N_7588);
and U8048 (N_8048,N_7777,N_7395);
nor U8049 (N_8049,N_7325,N_7722);
xor U8050 (N_8050,N_7299,N_7702);
xor U8051 (N_8051,N_7428,N_7498);
and U8052 (N_8052,N_7678,N_7641);
xor U8053 (N_8053,N_7600,N_7873);
and U8054 (N_8054,N_7881,N_7868);
or U8055 (N_8055,N_7880,N_7848);
or U8056 (N_8056,N_7555,N_7265);
xnor U8057 (N_8057,N_7750,N_7965);
or U8058 (N_8058,N_7521,N_7765);
or U8059 (N_8059,N_7224,N_7619);
nor U8060 (N_8060,N_7392,N_7691);
and U8061 (N_8061,N_7709,N_7656);
xnor U8062 (N_8062,N_7358,N_7344);
xnor U8063 (N_8063,N_7952,N_7734);
nor U8064 (N_8064,N_7471,N_7294);
xnor U8065 (N_8065,N_7815,N_7372);
and U8066 (N_8066,N_7563,N_7399);
nor U8067 (N_8067,N_7666,N_7539);
or U8068 (N_8068,N_7875,N_7307);
or U8069 (N_8069,N_7464,N_7650);
nand U8070 (N_8070,N_7234,N_7988);
nand U8071 (N_8071,N_7817,N_7413);
and U8072 (N_8072,N_7627,N_7744);
and U8073 (N_8073,N_7467,N_7495);
or U8074 (N_8074,N_7785,N_7382);
and U8075 (N_8075,N_7446,N_7576);
nand U8076 (N_8076,N_7824,N_7913);
nor U8077 (N_8077,N_7414,N_7981);
and U8078 (N_8078,N_7511,N_7746);
nand U8079 (N_8079,N_7583,N_7639);
xnor U8080 (N_8080,N_7887,N_7231);
nand U8081 (N_8081,N_7537,N_7856);
or U8082 (N_8082,N_7664,N_7669);
nand U8083 (N_8083,N_7361,N_7886);
nand U8084 (N_8084,N_7312,N_7791);
nor U8085 (N_8085,N_7992,N_7476);
xor U8086 (N_8086,N_7356,N_7523);
and U8087 (N_8087,N_7221,N_7697);
nand U8088 (N_8088,N_7999,N_7529);
nand U8089 (N_8089,N_7595,N_7686);
or U8090 (N_8090,N_7762,N_7412);
nor U8091 (N_8091,N_7936,N_7778);
nor U8092 (N_8092,N_7959,N_7401);
nor U8093 (N_8093,N_7604,N_7728);
nand U8094 (N_8094,N_7632,N_7316);
nand U8095 (N_8095,N_7794,N_7987);
xnor U8096 (N_8096,N_7603,N_7284);
and U8097 (N_8097,N_7648,N_7764);
xor U8098 (N_8098,N_7757,N_7489);
or U8099 (N_8099,N_7397,N_7874);
xnor U8100 (N_8100,N_7384,N_7819);
nand U8101 (N_8101,N_7437,N_7273);
and U8102 (N_8102,N_7388,N_7422);
nand U8103 (N_8103,N_7816,N_7261);
nand U8104 (N_8104,N_7483,N_7651);
and U8105 (N_8105,N_7956,N_7461);
nor U8106 (N_8106,N_7716,N_7324);
or U8107 (N_8107,N_7561,N_7766);
or U8108 (N_8108,N_7674,N_7918);
xnor U8109 (N_8109,N_7351,N_7532);
or U8110 (N_8110,N_7493,N_7429);
or U8111 (N_8111,N_7642,N_7542);
and U8112 (N_8112,N_7843,N_7821);
xnor U8113 (N_8113,N_7772,N_7371);
or U8114 (N_8114,N_7754,N_7628);
xnor U8115 (N_8115,N_7767,N_7834);
and U8116 (N_8116,N_7662,N_7288);
nand U8117 (N_8117,N_7836,N_7788);
or U8118 (N_8118,N_7434,N_7763);
nand U8119 (N_8119,N_7380,N_7237);
and U8120 (N_8120,N_7919,N_7911);
and U8121 (N_8121,N_7644,N_7582);
nand U8122 (N_8122,N_7331,N_7612);
nand U8123 (N_8123,N_7971,N_7465);
nor U8124 (N_8124,N_7640,N_7771);
nor U8125 (N_8125,N_7845,N_7801);
nor U8126 (N_8126,N_7853,N_7339);
nor U8127 (N_8127,N_7564,N_7942);
nand U8128 (N_8128,N_7783,N_7330);
and U8129 (N_8129,N_7688,N_7906);
xor U8130 (N_8130,N_7983,N_7657);
or U8131 (N_8131,N_7713,N_7494);
or U8132 (N_8132,N_7280,N_7786);
nand U8133 (N_8133,N_7225,N_7314);
xor U8134 (N_8134,N_7577,N_7473);
or U8135 (N_8135,N_7296,N_7710);
xnor U8136 (N_8136,N_7304,N_7758);
xor U8137 (N_8137,N_7424,N_7411);
nand U8138 (N_8138,N_7985,N_7624);
nor U8139 (N_8139,N_7272,N_7718);
or U8140 (N_8140,N_7775,N_7321);
nand U8141 (N_8141,N_7381,N_7486);
nand U8142 (N_8142,N_7247,N_7243);
nand U8143 (N_8143,N_7472,N_7295);
xnor U8144 (N_8144,N_7974,N_7903);
nor U8145 (N_8145,N_7892,N_7447);
nand U8146 (N_8146,N_7776,N_7336);
nand U8147 (N_8147,N_7941,N_7967);
and U8148 (N_8148,N_7254,N_7851);
nor U8149 (N_8149,N_7680,N_7431);
and U8150 (N_8150,N_7647,N_7573);
and U8151 (N_8151,N_7643,N_7850);
or U8152 (N_8152,N_7742,N_7665);
or U8153 (N_8153,N_7675,N_7546);
xor U8154 (N_8154,N_7951,N_7773);
xor U8155 (N_8155,N_7379,N_7479);
nand U8156 (N_8156,N_7796,N_7622);
nor U8157 (N_8157,N_7822,N_7589);
or U8158 (N_8158,N_7825,N_7590);
xor U8159 (N_8159,N_7482,N_7645);
nor U8160 (N_8160,N_7352,N_7220);
or U8161 (N_8161,N_7389,N_7503);
or U8162 (N_8162,N_7488,N_7623);
xnor U8163 (N_8163,N_7263,N_7275);
nand U8164 (N_8164,N_7867,N_7350);
and U8165 (N_8165,N_7510,N_7426);
and U8166 (N_8166,N_7730,N_7671);
nor U8167 (N_8167,N_7736,N_7696);
and U8168 (N_8168,N_7219,N_7516);
or U8169 (N_8169,N_7327,N_7244);
and U8170 (N_8170,N_7368,N_7932);
nor U8171 (N_8171,N_7719,N_7292);
xor U8172 (N_8172,N_7705,N_7893);
or U8173 (N_8173,N_7699,N_7406);
and U8174 (N_8174,N_7585,N_7281);
nor U8175 (N_8175,N_7964,N_7779);
nor U8176 (N_8176,N_7966,N_7636);
or U8177 (N_8177,N_7238,N_7832);
or U8178 (N_8178,N_7420,N_7293);
and U8179 (N_8179,N_7575,N_7228);
and U8180 (N_8180,N_7842,N_7393);
nand U8181 (N_8181,N_7386,N_7729);
xor U8182 (N_8182,N_7335,N_7871);
and U8183 (N_8183,N_7835,N_7720);
nor U8184 (N_8184,N_7207,N_7997);
or U8185 (N_8185,N_7457,N_7223);
xnor U8186 (N_8186,N_7844,N_7313);
nand U8187 (N_8187,N_7883,N_7855);
nand U8188 (N_8188,N_7269,N_7854);
xnor U8189 (N_8189,N_7509,N_7970);
nor U8190 (N_8190,N_7830,N_7706);
nand U8191 (N_8191,N_7550,N_7303);
or U8192 (N_8192,N_7553,N_7692);
or U8193 (N_8193,N_7427,N_7306);
nand U8194 (N_8194,N_7579,N_7438);
nor U8195 (N_8195,N_7248,N_7390);
and U8196 (N_8196,N_7962,N_7374);
or U8197 (N_8197,N_7580,N_7333);
nand U8198 (N_8198,N_7738,N_7954);
nor U8199 (N_8199,N_7963,N_7458);
xnor U8200 (N_8200,N_7229,N_7840);
nor U8201 (N_8201,N_7492,N_7435);
nor U8202 (N_8202,N_7679,N_7469);
nand U8203 (N_8203,N_7748,N_7813);
nor U8204 (N_8204,N_7876,N_7752);
xor U8205 (N_8205,N_7598,N_7897);
nor U8206 (N_8206,N_7899,N_7803);
and U8207 (N_8207,N_7721,N_7500);
nand U8208 (N_8208,N_7806,N_7416);
or U8209 (N_8209,N_7301,N_7298);
xor U8210 (N_8210,N_7814,N_7556);
nor U8211 (N_8211,N_7933,N_7441);
and U8212 (N_8212,N_7463,N_7276);
or U8213 (N_8213,N_7466,N_7531);
nand U8214 (N_8214,N_7976,N_7342);
xor U8215 (N_8215,N_7972,N_7833);
xnor U8216 (N_8216,N_7896,N_7560);
or U8217 (N_8217,N_7869,N_7934);
nand U8218 (N_8218,N_7210,N_7442);
xnor U8219 (N_8219,N_7711,N_7620);
and U8220 (N_8220,N_7898,N_7947);
nor U8221 (N_8221,N_7761,N_7245);
xnor U8222 (N_8222,N_7828,N_7841);
and U8223 (N_8223,N_7759,N_7795);
or U8224 (N_8224,N_7957,N_7267);
or U8225 (N_8225,N_7701,N_7444);
and U8226 (N_8226,N_7726,N_7633);
and U8227 (N_8227,N_7481,N_7613);
or U8228 (N_8228,N_7649,N_7849);
nand U8229 (N_8229,N_7407,N_7459);
xnor U8230 (N_8230,N_7405,N_7538);
and U8231 (N_8231,N_7986,N_7235);
or U8232 (N_8232,N_7993,N_7377);
nor U8233 (N_8233,N_7347,N_7343);
nor U8234 (N_8234,N_7968,N_7979);
xor U8235 (N_8235,N_7895,N_7931);
xnor U8236 (N_8236,N_7926,N_7663);
and U8237 (N_8237,N_7996,N_7362);
and U8238 (N_8238,N_7689,N_7271);
and U8239 (N_8239,N_7973,N_7345);
nor U8240 (N_8240,N_7230,N_7291);
nand U8241 (N_8241,N_7700,N_7337);
and U8242 (N_8242,N_7548,N_7250);
or U8243 (N_8243,N_7249,N_7638);
and U8244 (N_8244,N_7925,N_7214);
nand U8245 (N_8245,N_7512,N_7535);
and U8246 (N_8246,N_7980,N_7456);
nor U8247 (N_8247,N_7443,N_7989);
and U8248 (N_8248,N_7792,N_7928);
xnor U8249 (N_8249,N_7995,N_7436);
or U8250 (N_8250,N_7502,N_7798);
xnor U8251 (N_8251,N_7206,N_7953);
and U8252 (N_8252,N_7547,N_7982);
nand U8253 (N_8253,N_7927,N_7297);
or U8254 (N_8254,N_7559,N_7807);
or U8255 (N_8255,N_7530,N_7725);
nor U8256 (N_8256,N_7262,N_7609);
nor U8257 (N_8257,N_7670,N_7346);
nor U8258 (N_8258,N_7258,N_7860);
nor U8259 (N_8259,N_7800,N_7891);
or U8260 (N_8260,N_7818,N_7499);
xor U8261 (N_8261,N_7901,N_7514);
xor U8262 (N_8262,N_7749,N_7484);
or U8263 (N_8263,N_7549,N_7404);
nor U8264 (N_8264,N_7507,N_7360);
nor U8265 (N_8265,N_7373,N_7597);
nand U8266 (N_8266,N_7599,N_7592);
or U8267 (N_8267,N_7318,N_7812);
nor U8268 (N_8268,N_7367,N_7782);
xor U8269 (N_8269,N_7279,N_7408);
and U8270 (N_8270,N_7415,N_7226);
nor U8271 (N_8271,N_7252,N_7543);
and U8272 (N_8272,N_7227,N_7939);
nor U8273 (N_8273,N_7658,N_7823);
or U8274 (N_8274,N_7630,N_7653);
and U8275 (N_8275,N_7454,N_7938);
or U8276 (N_8276,N_7285,N_7311);
nor U8277 (N_8277,N_7423,N_7866);
nand U8278 (N_8278,N_7365,N_7496);
nand U8279 (N_8279,N_7491,N_7282);
and U8280 (N_8280,N_7487,N_7202);
nand U8281 (N_8281,N_7944,N_7506);
nand U8282 (N_8282,N_7541,N_7935);
nand U8283 (N_8283,N_7274,N_7445);
and U8284 (N_8284,N_7432,N_7357);
nor U8285 (N_8285,N_7940,N_7882);
xnor U8286 (N_8286,N_7672,N_7385);
and U8287 (N_8287,N_7755,N_7889);
xor U8288 (N_8288,N_7717,N_7684);
or U8289 (N_8289,N_7960,N_7837);
nor U8290 (N_8290,N_7300,N_7557);
nor U8291 (N_8291,N_7286,N_7707);
nand U8292 (N_8292,N_7802,N_7584);
or U8293 (N_8293,N_7991,N_7570);
nand U8294 (N_8294,N_7501,N_7606);
nand U8295 (N_8295,N_7242,N_7246);
and U8296 (N_8296,N_7945,N_7278);
or U8297 (N_8297,N_7740,N_7890);
or U8298 (N_8298,N_7216,N_7949);
and U8299 (N_8299,N_7930,N_7417);
nand U8300 (N_8300,N_7264,N_7687);
or U8301 (N_8301,N_7659,N_7376);
and U8302 (N_8302,N_7924,N_7359);
xor U8303 (N_8303,N_7602,N_7475);
xnor U8304 (N_8304,N_7878,N_7756);
and U8305 (N_8305,N_7733,N_7914);
nor U8306 (N_8306,N_7685,N_7239);
nor U8307 (N_8307,N_7277,N_7410);
nand U8308 (N_8308,N_7354,N_7315);
nand U8309 (N_8309,N_7634,N_7270);
nand U8310 (N_8310,N_7341,N_7654);
or U8311 (N_8311,N_7594,N_7723);
nand U8312 (N_8312,N_7703,N_7902);
nand U8313 (N_8313,N_7568,N_7240);
and U8314 (N_8314,N_7232,N_7865);
or U8315 (N_8315,N_7578,N_7694);
xnor U8316 (N_8316,N_7310,N_7943);
or U8317 (N_8317,N_7793,N_7477);
xor U8318 (N_8318,N_7683,N_7605);
and U8319 (N_8319,N_7540,N_7808);
or U8320 (N_8320,N_7369,N_7724);
and U8321 (N_8321,N_7859,N_7562);
or U8322 (N_8322,N_7534,N_7289);
nor U8323 (N_8323,N_7810,N_7787);
and U8324 (N_8324,N_7317,N_7676);
and U8325 (N_8325,N_7998,N_7545);
and U8326 (N_8326,N_7569,N_7652);
nor U8327 (N_8327,N_7574,N_7922);
and U8328 (N_8328,N_7328,N_7587);
nor U8329 (N_8329,N_7618,N_7858);
xor U8330 (N_8330,N_7375,N_7215);
and U8331 (N_8331,N_7485,N_7418);
or U8332 (N_8332,N_7453,N_7731);
nor U8333 (N_8333,N_7760,N_7355);
xor U8334 (N_8334,N_7451,N_7455);
nor U8335 (N_8335,N_7201,N_7212);
xor U8336 (N_8336,N_7505,N_7862);
nor U8337 (N_8337,N_7515,N_7400);
nor U8338 (N_8338,N_7211,N_7839);
nor U8339 (N_8339,N_7629,N_7955);
xor U8340 (N_8340,N_7268,N_7260);
or U8341 (N_8341,N_7635,N_7581);
xor U8342 (N_8342,N_7799,N_7203);
and U8343 (N_8343,N_7969,N_7984);
nor U8344 (N_8344,N_7525,N_7554);
and U8345 (N_8345,N_7601,N_7480);
nor U8346 (N_8346,N_7378,N_7462);
and U8347 (N_8347,N_7566,N_7266);
or U8348 (N_8348,N_7290,N_7527);
or U8349 (N_8349,N_7838,N_7704);
nand U8350 (N_8350,N_7217,N_7450);
nor U8351 (N_8351,N_7353,N_7452);
nand U8352 (N_8352,N_7915,N_7470);
and U8353 (N_8353,N_7789,N_7770);
xnor U8354 (N_8354,N_7781,N_7533);
or U8355 (N_8355,N_7667,N_7708);
or U8356 (N_8356,N_7977,N_7693);
and U8357 (N_8357,N_7743,N_7544);
or U8358 (N_8358,N_7528,N_7329);
and U8359 (N_8359,N_7668,N_7831);
xor U8360 (N_8360,N_7302,N_7961);
and U8361 (N_8361,N_7253,N_7593);
xnor U8362 (N_8362,N_7387,N_7370);
nor U8363 (N_8363,N_7905,N_7558);
xnor U8364 (N_8364,N_7615,N_7879);
nand U8365 (N_8365,N_7768,N_7948);
or U8366 (N_8366,N_7614,N_7631);
xnor U8367 (N_8367,N_7637,N_7769);
xnor U8368 (N_8368,N_7519,N_7257);
or U8369 (N_8369,N_7805,N_7937);
or U8370 (N_8370,N_7829,N_7305);
nor U8371 (N_8371,N_7474,N_7780);
xor U8372 (N_8372,N_7826,N_7872);
nand U8373 (N_8373,N_7673,N_7745);
nand U8374 (N_8374,N_7334,N_7827);
nor U8375 (N_8375,N_7804,N_7916);
nor U8376 (N_8376,N_7784,N_7200);
xnor U8377 (N_8377,N_7975,N_7591);
and U8378 (N_8378,N_7571,N_7468);
xnor U8379 (N_8379,N_7661,N_7857);
or U8380 (N_8380,N_7900,N_7433);
and U8381 (N_8381,N_7256,N_7608);
or U8382 (N_8382,N_7617,N_7990);
and U8383 (N_8383,N_7917,N_7448);
xnor U8384 (N_8384,N_7820,N_7204);
nor U8385 (N_8385,N_7572,N_7309);
xnor U8386 (N_8386,N_7912,N_7409);
or U8387 (N_8387,N_7209,N_7430);
xor U8388 (N_8388,N_7908,N_7251);
or U8389 (N_8389,N_7323,N_7655);
or U8390 (N_8390,N_7695,N_7460);
xnor U8391 (N_8391,N_7233,N_7714);
nor U8392 (N_8392,N_7739,N_7402);
xnor U8393 (N_8393,N_7205,N_7958);
or U8394 (N_8394,N_7626,N_7727);
and U8395 (N_8395,N_7218,N_7929);
and U8396 (N_8396,N_7864,N_7522);
nor U8397 (N_8397,N_7567,N_7439);
and U8398 (N_8398,N_7383,N_7660);
and U8399 (N_8399,N_7904,N_7513);
nor U8400 (N_8400,N_7941,N_7353);
nand U8401 (N_8401,N_7778,N_7545);
nand U8402 (N_8402,N_7710,N_7843);
xor U8403 (N_8403,N_7430,N_7475);
nand U8404 (N_8404,N_7812,N_7751);
or U8405 (N_8405,N_7473,N_7723);
nor U8406 (N_8406,N_7551,N_7532);
xor U8407 (N_8407,N_7269,N_7437);
or U8408 (N_8408,N_7440,N_7469);
or U8409 (N_8409,N_7978,N_7933);
xor U8410 (N_8410,N_7816,N_7460);
or U8411 (N_8411,N_7774,N_7786);
nor U8412 (N_8412,N_7656,N_7640);
nand U8413 (N_8413,N_7216,N_7513);
nand U8414 (N_8414,N_7395,N_7890);
nor U8415 (N_8415,N_7464,N_7597);
nor U8416 (N_8416,N_7424,N_7535);
nand U8417 (N_8417,N_7217,N_7532);
nor U8418 (N_8418,N_7509,N_7576);
and U8419 (N_8419,N_7725,N_7684);
nor U8420 (N_8420,N_7695,N_7213);
and U8421 (N_8421,N_7348,N_7250);
or U8422 (N_8422,N_7488,N_7956);
nor U8423 (N_8423,N_7973,N_7806);
nor U8424 (N_8424,N_7560,N_7806);
and U8425 (N_8425,N_7329,N_7726);
and U8426 (N_8426,N_7877,N_7694);
and U8427 (N_8427,N_7213,N_7849);
nand U8428 (N_8428,N_7503,N_7324);
nand U8429 (N_8429,N_7943,N_7358);
or U8430 (N_8430,N_7450,N_7603);
nor U8431 (N_8431,N_7461,N_7209);
nor U8432 (N_8432,N_7446,N_7301);
xnor U8433 (N_8433,N_7689,N_7625);
nand U8434 (N_8434,N_7783,N_7263);
or U8435 (N_8435,N_7273,N_7705);
or U8436 (N_8436,N_7949,N_7323);
or U8437 (N_8437,N_7993,N_7688);
or U8438 (N_8438,N_7495,N_7776);
xor U8439 (N_8439,N_7620,N_7437);
nor U8440 (N_8440,N_7792,N_7948);
nand U8441 (N_8441,N_7880,N_7975);
nand U8442 (N_8442,N_7301,N_7904);
xor U8443 (N_8443,N_7363,N_7212);
or U8444 (N_8444,N_7903,N_7671);
xnor U8445 (N_8445,N_7794,N_7301);
nand U8446 (N_8446,N_7719,N_7213);
and U8447 (N_8447,N_7323,N_7712);
and U8448 (N_8448,N_7784,N_7816);
and U8449 (N_8449,N_7985,N_7556);
nor U8450 (N_8450,N_7639,N_7736);
xnor U8451 (N_8451,N_7516,N_7745);
xnor U8452 (N_8452,N_7942,N_7611);
nand U8453 (N_8453,N_7772,N_7671);
and U8454 (N_8454,N_7600,N_7920);
and U8455 (N_8455,N_7760,N_7580);
xnor U8456 (N_8456,N_7848,N_7275);
xnor U8457 (N_8457,N_7730,N_7401);
xnor U8458 (N_8458,N_7664,N_7431);
xnor U8459 (N_8459,N_7261,N_7327);
and U8460 (N_8460,N_7931,N_7628);
or U8461 (N_8461,N_7430,N_7254);
xnor U8462 (N_8462,N_7772,N_7322);
nand U8463 (N_8463,N_7292,N_7975);
and U8464 (N_8464,N_7471,N_7592);
xor U8465 (N_8465,N_7898,N_7627);
nor U8466 (N_8466,N_7667,N_7471);
nand U8467 (N_8467,N_7650,N_7503);
or U8468 (N_8468,N_7302,N_7496);
and U8469 (N_8469,N_7858,N_7208);
nand U8470 (N_8470,N_7739,N_7446);
xor U8471 (N_8471,N_7416,N_7469);
and U8472 (N_8472,N_7410,N_7562);
and U8473 (N_8473,N_7919,N_7565);
nor U8474 (N_8474,N_7983,N_7596);
nand U8475 (N_8475,N_7871,N_7219);
xnor U8476 (N_8476,N_7833,N_7518);
nand U8477 (N_8477,N_7711,N_7772);
xnor U8478 (N_8478,N_7635,N_7423);
nor U8479 (N_8479,N_7891,N_7900);
xnor U8480 (N_8480,N_7789,N_7499);
xnor U8481 (N_8481,N_7335,N_7817);
xor U8482 (N_8482,N_7266,N_7375);
xor U8483 (N_8483,N_7703,N_7996);
xor U8484 (N_8484,N_7789,N_7531);
xor U8485 (N_8485,N_7919,N_7339);
xor U8486 (N_8486,N_7898,N_7992);
nand U8487 (N_8487,N_7648,N_7378);
and U8488 (N_8488,N_7653,N_7671);
nand U8489 (N_8489,N_7959,N_7747);
and U8490 (N_8490,N_7994,N_7667);
nand U8491 (N_8491,N_7800,N_7277);
nor U8492 (N_8492,N_7866,N_7811);
xnor U8493 (N_8493,N_7633,N_7892);
and U8494 (N_8494,N_7563,N_7813);
nand U8495 (N_8495,N_7300,N_7342);
xnor U8496 (N_8496,N_7932,N_7670);
xor U8497 (N_8497,N_7945,N_7260);
nor U8498 (N_8498,N_7463,N_7617);
and U8499 (N_8499,N_7989,N_7528);
nor U8500 (N_8500,N_7706,N_7521);
nand U8501 (N_8501,N_7348,N_7360);
nor U8502 (N_8502,N_7408,N_7659);
nand U8503 (N_8503,N_7980,N_7986);
and U8504 (N_8504,N_7841,N_7412);
xor U8505 (N_8505,N_7792,N_7659);
and U8506 (N_8506,N_7919,N_7642);
nor U8507 (N_8507,N_7823,N_7346);
xor U8508 (N_8508,N_7940,N_7221);
and U8509 (N_8509,N_7808,N_7207);
or U8510 (N_8510,N_7745,N_7777);
nor U8511 (N_8511,N_7428,N_7544);
or U8512 (N_8512,N_7975,N_7781);
xnor U8513 (N_8513,N_7926,N_7540);
nand U8514 (N_8514,N_7978,N_7738);
nor U8515 (N_8515,N_7371,N_7213);
xor U8516 (N_8516,N_7968,N_7570);
or U8517 (N_8517,N_7340,N_7818);
nor U8518 (N_8518,N_7652,N_7314);
or U8519 (N_8519,N_7969,N_7663);
nor U8520 (N_8520,N_7856,N_7839);
xnor U8521 (N_8521,N_7428,N_7954);
nand U8522 (N_8522,N_7487,N_7926);
or U8523 (N_8523,N_7335,N_7529);
and U8524 (N_8524,N_7215,N_7593);
xor U8525 (N_8525,N_7293,N_7248);
nand U8526 (N_8526,N_7716,N_7307);
xnor U8527 (N_8527,N_7897,N_7536);
nor U8528 (N_8528,N_7820,N_7314);
nand U8529 (N_8529,N_7831,N_7962);
xor U8530 (N_8530,N_7873,N_7543);
nand U8531 (N_8531,N_7917,N_7684);
and U8532 (N_8532,N_7954,N_7532);
or U8533 (N_8533,N_7302,N_7846);
nand U8534 (N_8534,N_7637,N_7703);
and U8535 (N_8535,N_7239,N_7717);
xor U8536 (N_8536,N_7815,N_7422);
nor U8537 (N_8537,N_7488,N_7654);
or U8538 (N_8538,N_7232,N_7974);
nand U8539 (N_8539,N_7439,N_7707);
nand U8540 (N_8540,N_7883,N_7343);
nor U8541 (N_8541,N_7407,N_7920);
and U8542 (N_8542,N_7631,N_7555);
and U8543 (N_8543,N_7440,N_7824);
and U8544 (N_8544,N_7604,N_7803);
xnor U8545 (N_8545,N_7880,N_7638);
xnor U8546 (N_8546,N_7609,N_7414);
nand U8547 (N_8547,N_7238,N_7781);
nand U8548 (N_8548,N_7587,N_7418);
xnor U8549 (N_8549,N_7315,N_7557);
xor U8550 (N_8550,N_7516,N_7446);
and U8551 (N_8551,N_7670,N_7994);
xor U8552 (N_8552,N_7888,N_7915);
and U8553 (N_8553,N_7965,N_7734);
nand U8554 (N_8554,N_7666,N_7285);
nand U8555 (N_8555,N_7482,N_7788);
or U8556 (N_8556,N_7506,N_7953);
and U8557 (N_8557,N_7333,N_7246);
xnor U8558 (N_8558,N_7434,N_7379);
or U8559 (N_8559,N_7922,N_7982);
and U8560 (N_8560,N_7642,N_7907);
xor U8561 (N_8561,N_7789,N_7224);
or U8562 (N_8562,N_7839,N_7732);
nor U8563 (N_8563,N_7994,N_7738);
nor U8564 (N_8564,N_7639,N_7769);
nor U8565 (N_8565,N_7414,N_7373);
nand U8566 (N_8566,N_7527,N_7678);
xor U8567 (N_8567,N_7252,N_7501);
nand U8568 (N_8568,N_7844,N_7294);
and U8569 (N_8569,N_7239,N_7549);
nand U8570 (N_8570,N_7726,N_7352);
or U8571 (N_8571,N_7877,N_7329);
nor U8572 (N_8572,N_7363,N_7685);
and U8573 (N_8573,N_7872,N_7451);
or U8574 (N_8574,N_7889,N_7453);
or U8575 (N_8575,N_7808,N_7960);
xor U8576 (N_8576,N_7510,N_7381);
nor U8577 (N_8577,N_7903,N_7969);
nand U8578 (N_8578,N_7385,N_7742);
xnor U8579 (N_8579,N_7322,N_7405);
nor U8580 (N_8580,N_7382,N_7609);
or U8581 (N_8581,N_7681,N_7584);
xnor U8582 (N_8582,N_7657,N_7677);
nor U8583 (N_8583,N_7652,N_7999);
or U8584 (N_8584,N_7728,N_7366);
nor U8585 (N_8585,N_7514,N_7706);
xor U8586 (N_8586,N_7620,N_7270);
nor U8587 (N_8587,N_7879,N_7372);
or U8588 (N_8588,N_7567,N_7864);
nand U8589 (N_8589,N_7567,N_7683);
and U8590 (N_8590,N_7852,N_7634);
and U8591 (N_8591,N_7869,N_7303);
and U8592 (N_8592,N_7977,N_7947);
or U8593 (N_8593,N_7487,N_7785);
nand U8594 (N_8594,N_7374,N_7615);
or U8595 (N_8595,N_7959,N_7856);
nand U8596 (N_8596,N_7600,N_7660);
nand U8597 (N_8597,N_7295,N_7982);
nor U8598 (N_8598,N_7658,N_7263);
or U8599 (N_8599,N_7839,N_7232);
and U8600 (N_8600,N_7642,N_7412);
and U8601 (N_8601,N_7429,N_7532);
and U8602 (N_8602,N_7704,N_7311);
nand U8603 (N_8603,N_7217,N_7898);
nor U8604 (N_8604,N_7521,N_7306);
or U8605 (N_8605,N_7407,N_7837);
or U8606 (N_8606,N_7731,N_7748);
and U8607 (N_8607,N_7202,N_7227);
nor U8608 (N_8608,N_7478,N_7940);
nor U8609 (N_8609,N_7993,N_7994);
or U8610 (N_8610,N_7356,N_7420);
nor U8611 (N_8611,N_7593,N_7628);
nor U8612 (N_8612,N_7743,N_7741);
and U8613 (N_8613,N_7833,N_7357);
nor U8614 (N_8614,N_7700,N_7581);
and U8615 (N_8615,N_7533,N_7355);
nand U8616 (N_8616,N_7894,N_7659);
nor U8617 (N_8617,N_7400,N_7419);
or U8618 (N_8618,N_7973,N_7561);
xor U8619 (N_8619,N_7618,N_7270);
xor U8620 (N_8620,N_7770,N_7549);
or U8621 (N_8621,N_7604,N_7504);
xor U8622 (N_8622,N_7251,N_7273);
nor U8623 (N_8623,N_7991,N_7492);
nand U8624 (N_8624,N_7809,N_7507);
and U8625 (N_8625,N_7446,N_7367);
nand U8626 (N_8626,N_7900,N_7873);
nand U8627 (N_8627,N_7438,N_7255);
nor U8628 (N_8628,N_7402,N_7943);
nor U8629 (N_8629,N_7603,N_7988);
xnor U8630 (N_8630,N_7596,N_7558);
xor U8631 (N_8631,N_7778,N_7600);
and U8632 (N_8632,N_7371,N_7232);
and U8633 (N_8633,N_7878,N_7538);
or U8634 (N_8634,N_7524,N_7889);
or U8635 (N_8635,N_7733,N_7613);
xor U8636 (N_8636,N_7832,N_7856);
xor U8637 (N_8637,N_7398,N_7737);
xor U8638 (N_8638,N_7303,N_7342);
xor U8639 (N_8639,N_7286,N_7669);
xor U8640 (N_8640,N_7884,N_7975);
or U8641 (N_8641,N_7941,N_7386);
nand U8642 (N_8642,N_7270,N_7408);
and U8643 (N_8643,N_7439,N_7589);
and U8644 (N_8644,N_7803,N_7296);
or U8645 (N_8645,N_7212,N_7840);
or U8646 (N_8646,N_7267,N_7255);
or U8647 (N_8647,N_7340,N_7388);
or U8648 (N_8648,N_7409,N_7533);
nor U8649 (N_8649,N_7444,N_7353);
nor U8650 (N_8650,N_7755,N_7301);
and U8651 (N_8651,N_7860,N_7539);
nor U8652 (N_8652,N_7710,N_7397);
or U8653 (N_8653,N_7318,N_7400);
nor U8654 (N_8654,N_7897,N_7736);
nand U8655 (N_8655,N_7987,N_7711);
nand U8656 (N_8656,N_7278,N_7284);
and U8657 (N_8657,N_7291,N_7425);
and U8658 (N_8658,N_7303,N_7475);
and U8659 (N_8659,N_7747,N_7918);
nor U8660 (N_8660,N_7819,N_7812);
or U8661 (N_8661,N_7438,N_7356);
xnor U8662 (N_8662,N_7387,N_7911);
nor U8663 (N_8663,N_7477,N_7657);
nor U8664 (N_8664,N_7791,N_7468);
and U8665 (N_8665,N_7397,N_7310);
nor U8666 (N_8666,N_7987,N_7302);
nand U8667 (N_8667,N_7527,N_7819);
xor U8668 (N_8668,N_7300,N_7907);
nor U8669 (N_8669,N_7780,N_7826);
nand U8670 (N_8670,N_7734,N_7368);
nand U8671 (N_8671,N_7918,N_7489);
nand U8672 (N_8672,N_7462,N_7936);
and U8673 (N_8673,N_7589,N_7383);
nor U8674 (N_8674,N_7896,N_7604);
or U8675 (N_8675,N_7747,N_7652);
or U8676 (N_8676,N_7208,N_7571);
xnor U8677 (N_8677,N_7691,N_7791);
nor U8678 (N_8678,N_7968,N_7627);
xnor U8679 (N_8679,N_7768,N_7982);
and U8680 (N_8680,N_7759,N_7727);
xor U8681 (N_8681,N_7993,N_7277);
nor U8682 (N_8682,N_7561,N_7968);
xor U8683 (N_8683,N_7336,N_7209);
xor U8684 (N_8684,N_7536,N_7803);
xor U8685 (N_8685,N_7623,N_7227);
and U8686 (N_8686,N_7246,N_7386);
xor U8687 (N_8687,N_7204,N_7938);
and U8688 (N_8688,N_7379,N_7889);
xnor U8689 (N_8689,N_7477,N_7993);
and U8690 (N_8690,N_7469,N_7464);
nand U8691 (N_8691,N_7364,N_7298);
and U8692 (N_8692,N_7776,N_7554);
nor U8693 (N_8693,N_7782,N_7669);
and U8694 (N_8694,N_7498,N_7892);
and U8695 (N_8695,N_7665,N_7830);
nor U8696 (N_8696,N_7219,N_7959);
or U8697 (N_8697,N_7445,N_7757);
and U8698 (N_8698,N_7968,N_7582);
or U8699 (N_8699,N_7445,N_7815);
nand U8700 (N_8700,N_7368,N_7282);
and U8701 (N_8701,N_7846,N_7634);
and U8702 (N_8702,N_7264,N_7303);
xor U8703 (N_8703,N_7962,N_7244);
and U8704 (N_8704,N_7577,N_7332);
or U8705 (N_8705,N_7678,N_7955);
xor U8706 (N_8706,N_7987,N_7428);
or U8707 (N_8707,N_7629,N_7630);
or U8708 (N_8708,N_7663,N_7632);
and U8709 (N_8709,N_7221,N_7355);
xnor U8710 (N_8710,N_7760,N_7437);
nor U8711 (N_8711,N_7750,N_7476);
nor U8712 (N_8712,N_7835,N_7366);
nand U8713 (N_8713,N_7510,N_7704);
nand U8714 (N_8714,N_7407,N_7314);
xnor U8715 (N_8715,N_7757,N_7236);
nor U8716 (N_8716,N_7601,N_7382);
and U8717 (N_8717,N_7597,N_7910);
nand U8718 (N_8718,N_7937,N_7977);
or U8719 (N_8719,N_7596,N_7359);
and U8720 (N_8720,N_7882,N_7440);
xor U8721 (N_8721,N_7645,N_7952);
nand U8722 (N_8722,N_7302,N_7995);
or U8723 (N_8723,N_7690,N_7564);
or U8724 (N_8724,N_7360,N_7939);
xnor U8725 (N_8725,N_7499,N_7372);
and U8726 (N_8726,N_7772,N_7514);
xnor U8727 (N_8727,N_7598,N_7389);
nand U8728 (N_8728,N_7204,N_7646);
xnor U8729 (N_8729,N_7695,N_7759);
and U8730 (N_8730,N_7234,N_7621);
nand U8731 (N_8731,N_7804,N_7844);
xnor U8732 (N_8732,N_7279,N_7521);
or U8733 (N_8733,N_7606,N_7526);
and U8734 (N_8734,N_7553,N_7927);
or U8735 (N_8735,N_7647,N_7202);
xnor U8736 (N_8736,N_7707,N_7988);
nor U8737 (N_8737,N_7981,N_7615);
or U8738 (N_8738,N_7567,N_7771);
or U8739 (N_8739,N_7695,N_7334);
nand U8740 (N_8740,N_7631,N_7377);
and U8741 (N_8741,N_7879,N_7839);
nand U8742 (N_8742,N_7337,N_7825);
or U8743 (N_8743,N_7254,N_7547);
nor U8744 (N_8744,N_7734,N_7808);
xor U8745 (N_8745,N_7878,N_7642);
or U8746 (N_8746,N_7967,N_7926);
nand U8747 (N_8747,N_7768,N_7777);
nor U8748 (N_8748,N_7210,N_7703);
nand U8749 (N_8749,N_7920,N_7786);
xor U8750 (N_8750,N_7307,N_7247);
nand U8751 (N_8751,N_7377,N_7438);
and U8752 (N_8752,N_7236,N_7680);
or U8753 (N_8753,N_7826,N_7581);
or U8754 (N_8754,N_7781,N_7900);
nand U8755 (N_8755,N_7452,N_7883);
and U8756 (N_8756,N_7433,N_7851);
nor U8757 (N_8757,N_7822,N_7914);
and U8758 (N_8758,N_7593,N_7812);
or U8759 (N_8759,N_7807,N_7714);
and U8760 (N_8760,N_7237,N_7314);
and U8761 (N_8761,N_7994,N_7611);
xnor U8762 (N_8762,N_7264,N_7973);
nand U8763 (N_8763,N_7556,N_7698);
xor U8764 (N_8764,N_7243,N_7872);
xor U8765 (N_8765,N_7938,N_7549);
nand U8766 (N_8766,N_7969,N_7673);
xor U8767 (N_8767,N_7522,N_7454);
or U8768 (N_8768,N_7495,N_7787);
xnor U8769 (N_8769,N_7513,N_7251);
nor U8770 (N_8770,N_7376,N_7676);
xnor U8771 (N_8771,N_7322,N_7688);
nand U8772 (N_8772,N_7732,N_7378);
xor U8773 (N_8773,N_7544,N_7526);
nor U8774 (N_8774,N_7285,N_7929);
and U8775 (N_8775,N_7344,N_7661);
nor U8776 (N_8776,N_7715,N_7260);
nor U8777 (N_8777,N_7788,N_7585);
or U8778 (N_8778,N_7937,N_7925);
nand U8779 (N_8779,N_7405,N_7852);
nand U8780 (N_8780,N_7561,N_7522);
xnor U8781 (N_8781,N_7958,N_7605);
nor U8782 (N_8782,N_7856,N_7923);
nand U8783 (N_8783,N_7613,N_7546);
nor U8784 (N_8784,N_7651,N_7510);
nor U8785 (N_8785,N_7404,N_7285);
or U8786 (N_8786,N_7441,N_7334);
nand U8787 (N_8787,N_7934,N_7250);
nand U8788 (N_8788,N_7212,N_7479);
nor U8789 (N_8789,N_7790,N_7430);
nor U8790 (N_8790,N_7669,N_7585);
or U8791 (N_8791,N_7248,N_7929);
nand U8792 (N_8792,N_7920,N_7539);
nor U8793 (N_8793,N_7668,N_7956);
xor U8794 (N_8794,N_7906,N_7535);
xnor U8795 (N_8795,N_7656,N_7735);
nand U8796 (N_8796,N_7960,N_7751);
nor U8797 (N_8797,N_7655,N_7785);
nor U8798 (N_8798,N_7835,N_7952);
nand U8799 (N_8799,N_7445,N_7544);
nor U8800 (N_8800,N_8477,N_8324);
or U8801 (N_8801,N_8684,N_8545);
nor U8802 (N_8802,N_8311,N_8694);
nor U8803 (N_8803,N_8372,N_8230);
nor U8804 (N_8804,N_8592,N_8280);
or U8805 (N_8805,N_8681,N_8183);
nand U8806 (N_8806,N_8375,N_8757);
or U8807 (N_8807,N_8362,N_8649);
nor U8808 (N_8808,N_8504,N_8748);
or U8809 (N_8809,N_8431,N_8312);
and U8810 (N_8810,N_8089,N_8038);
xor U8811 (N_8811,N_8162,N_8202);
nor U8812 (N_8812,N_8598,N_8701);
or U8813 (N_8813,N_8692,N_8783);
nand U8814 (N_8814,N_8107,N_8277);
xor U8815 (N_8815,N_8672,N_8423);
nor U8816 (N_8816,N_8747,N_8315);
nor U8817 (N_8817,N_8473,N_8133);
or U8818 (N_8818,N_8779,N_8199);
and U8819 (N_8819,N_8485,N_8191);
nor U8820 (N_8820,N_8009,N_8755);
and U8821 (N_8821,N_8480,N_8627);
nor U8822 (N_8822,N_8554,N_8391);
or U8823 (N_8823,N_8261,N_8765);
xnor U8824 (N_8824,N_8051,N_8588);
xnor U8825 (N_8825,N_8031,N_8101);
and U8826 (N_8826,N_8212,N_8460);
and U8827 (N_8827,N_8023,N_8158);
nand U8828 (N_8828,N_8656,N_8514);
and U8829 (N_8829,N_8319,N_8658);
nor U8830 (N_8830,N_8635,N_8595);
or U8831 (N_8831,N_8087,N_8267);
nor U8832 (N_8832,N_8518,N_8785);
or U8833 (N_8833,N_8169,N_8088);
nor U8834 (N_8834,N_8084,N_8299);
nand U8835 (N_8835,N_8585,N_8578);
nor U8836 (N_8836,N_8249,N_8095);
nor U8837 (N_8837,N_8043,N_8664);
nor U8838 (N_8838,N_8110,N_8078);
nand U8839 (N_8839,N_8502,N_8237);
and U8840 (N_8840,N_8631,N_8003);
and U8841 (N_8841,N_8296,N_8198);
nor U8842 (N_8842,N_8053,N_8390);
xnor U8843 (N_8843,N_8516,N_8062);
xor U8844 (N_8844,N_8234,N_8594);
nor U8845 (N_8845,N_8490,N_8703);
and U8846 (N_8846,N_8400,N_8710);
xnor U8847 (N_8847,N_8056,N_8629);
and U8848 (N_8848,N_8609,N_8732);
nand U8849 (N_8849,N_8175,N_8601);
and U8850 (N_8850,N_8418,N_8626);
nand U8851 (N_8851,N_8569,N_8313);
and U8852 (N_8852,N_8673,N_8690);
or U8853 (N_8853,N_8793,N_8790);
xnor U8854 (N_8854,N_8462,N_8528);
xor U8855 (N_8855,N_8276,N_8714);
xnor U8856 (N_8856,N_8103,N_8674);
nor U8857 (N_8857,N_8695,N_8567);
and U8858 (N_8858,N_8558,N_8345);
nor U8859 (N_8859,N_8069,N_8409);
and U8860 (N_8860,N_8467,N_8449);
and U8861 (N_8861,N_8229,N_8723);
or U8862 (N_8862,N_8144,N_8411);
xnor U8863 (N_8863,N_8041,N_8711);
nor U8864 (N_8864,N_8641,N_8179);
nor U8865 (N_8865,N_8688,N_8314);
nand U8866 (N_8866,N_8549,N_8253);
and U8867 (N_8867,N_8729,N_8301);
and U8868 (N_8868,N_8021,N_8660);
nor U8869 (N_8869,N_8424,N_8376);
nor U8870 (N_8870,N_8553,N_8140);
nand U8871 (N_8871,N_8541,N_8392);
and U8872 (N_8872,N_8282,N_8116);
xor U8873 (N_8873,N_8736,N_8278);
or U8874 (N_8874,N_8515,N_8603);
nor U8875 (N_8875,N_8758,N_8383);
or U8876 (N_8876,N_8086,N_8037);
nor U8877 (N_8877,N_8241,N_8573);
nand U8878 (N_8878,N_8250,N_8117);
xor U8879 (N_8879,N_8568,N_8652);
xnor U8880 (N_8880,N_8364,N_8283);
nand U8881 (N_8881,N_8269,N_8587);
xnor U8882 (N_8882,N_8094,N_8063);
and U8883 (N_8883,N_8483,N_8047);
nor U8884 (N_8884,N_8525,N_8511);
xnor U8885 (N_8885,N_8339,N_8147);
nand U8886 (N_8886,N_8709,N_8610);
xor U8887 (N_8887,N_8772,N_8002);
and U8888 (N_8888,N_8176,N_8687);
xnor U8889 (N_8889,N_8799,N_8746);
xnor U8890 (N_8890,N_8605,N_8228);
xor U8891 (N_8891,N_8427,N_8214);
nor U8892 (N_8892,N_8150,N_8293);
or U8893 (N_8893,N_8120,N_8328);
and U8894 (N_8894,N_8033,N_8520);
or U8895 (N_8895,N_8190,N_8034);
nand U8896 (N_8896,N_8638,N_8481);
or U8897 (N_8897,N_8661,N_8343);
xor U8898 (N_8898,N_8090,N_8264);
xor U8899 (N_8899,N_8721,N_8048);
or U8900 (N_8900,N_8153,N_8497);
xnor U8901 (N_8901,N_8355,N_8239);
nand U8902 (N_8902,N_8042,N_8219);
nor U8903 (N_8903,N_8071,N_8479);
nand U8904 (N_8904,N_8618,N_8671);
xnor U8905 (N_8905,N_8776,N_8039);
and U8906 (N_8906,N_8458,N_8074);
nand U8907 (N_8907,N_8471,N_8001);
or U8908 (N_8908,N_8354,N_8243);
nand U8909 (N_8909,N_8767,N_8226);
nor U8910 (N_8910,N_8489,N_8630);
xor U8911 (N_8911,N_8338,N_8507);
and U8912 (N_8912,N_8075,N_8281);
nor U8913 (N_8913,N_8099,N_8413);
nand U8914 (N_8914,N_8509,N_8579);
and U8915 (N_8915,N_8717,N_8325);
and U8916 (N_8916,N_8559,N_8194);
nand U8917 (N_8917,N_8361,N_8650);
and U8918 (N_8918,N_8719,N_8675);
nor U8919 (N_8919,N_8256,N_8771);
nand U8920 (N_8920,N_8181,N_8255);
nand U8921 (N_8921,N_8538,N_8308);
nand U8922 (N_8922,N_8118,N_8007);
xor U8923 (N_8923,N_8450,N_8220);
or U8924 (N_8924,N_8204,N_8055);
xor U8925 (N_8925,N_8070,N_8533);
nand U8926 (N_8926,N_8059,N_8524);
nand U8927 (N_8927,N_8026,N_8535);
nor U8928 (N_8928,N_8326,N_8552);
nor U8929 (N_8929,N_8546,N_8307);
and U8930 (N_8930,N_8164,N_8182);
nor U8931 (N_8931,N_8309,N_8741);
or U8932 (N_8932,N_8706,N_8344);
nor U8933 (N_8933,N_8446,N_8434);
nand U8934 (N_8934,N_8699,N_8209);
xnor U8935 (N_8935,N_8349,N_8384);
xnor U8936 (N_8936,N_8447,N_8780);
nor U8937 (N_8937,N_8404,N_8396);
nor U8938 (N_8938,N_8642,N_8461);
and U8939 (N_8939,N_8640,N_8334);
and U8940 (N_8940,N_8764,N_8297);
nor U8941 (N_8941,N_8134,N_8245);
nand U8942 (N_8942,N_8288,N_8091);
nand U8943 (N_8943,N_8123,N_8024);
or U8944 (N_8944,N_8527,N_8625);
and U8945 (N_8945,N_8663,N_8646);
nand U8946 (N_8946,N_8213,N_8359);
nor U8947 (N_8947,N_8268,N_8200);
nor U8948 (N_8948,N_8459,N_8797);
nand U8949 (N_8949,N_8718,N_8682);
nor U8950 (N_8950,N_8284,N_8125);
nand U8951 (N_8951,N_8342,N_8734);
xor U8952 (N_8952,N_8006,N_8798);
or U8953 (N_8953,N_8020,N_8348);
and U8954 (N_8954,N_8068,N_8104);
or U8955 (N_8955,N_8464,N_8680);
or U8956 (N_8956,N_8394,N_8218);
and U8957 (N_8957,N_8224,N_8697);
nor U8958 (N_8958,N_8614,N_8337);
or U8959 (N_8959,N_8725,N_8487);
or U8960 (N_8960,N_8557,N_8763);
nand U8961 (N_8961,N_8290,N_8628);
nand U8962 (N_8962,N_8265,N_8122);
or U8963 (N_8963,N_8556,N_8600);
xnor U8964 (N_8964,N_8401,N_8180);
and U8965 (N_8965,N_8724,N_8248);
or U8966 (N_8966,N_8437,N_8433);
or U8967 (N_8967,N_8634,N_8065);
and U8968 (N_8968,N_8367,N_8659);
and U8969 (N_8969,N_8512,N_8072);
nand U8970 (N_8970,N_8292,N_8114);
nand U8971 (N_8971,N_8583,N_8124);
or U8972 (N_8972,N_8206,N_8574);
and U8973 (N_8973,N_8049,N_8111);
nand U8974 (N_8974,N_8470,N_8670);
or U8975 (N_8975,N_8310,N_8686);
xor U8976 (N_8976,N_8782,N_8662);
xnor U8977 (N_8977,N_8531,N_8773);
and U8978 (N_8978,N_8454,N_8227);
xnor U8979 (N_8979,N_8657,N_8542);
nand U8980 (N_8980,N_8073,N_8060);
nand U8981 (N_8981,N_8215,N_8728);
and U8982 (N_8982,N_8366,N_8045);
or U8983 (N_8983,N_8160,N_8781);
nand U8984 (N_8984,N_8128,N_8655);
and U8985 (N_8985,N_8145,N_8014);
and U8986 (N_8986,N_8258,N_8453);
nand U8987 (N_8987,N_8607,N_8193);
nor U8988 (N_8988,N_8373,N_8146);
or U8989 (N_8989,N_8027,N_8572);
nor U8990 (N_8990,N_8010,N_8352);
xor U8991 (N_8991,N_8238,N_8207);
nand U8992 (N_8992,N_8406,N_8496);
or U8993 (N_8993,N_8223,N_8632);
nand U8994 (N_8994,N_8320,N_8331);
or U8995 (N_8995,N_8498,N_8156);
nor U8996 (N_8996,N_8102,N_8571);
nand U8997 (N_8997,N_8189,N_8129);
and U8998 (N_8998,N_8380,N_8251);
nand U8999 (N_8999,N_8653,N_8097);
and U9000 (N_9000,N_8526,N_8197);
and U9001 (N_9001,N_8275,N_8612);
or U9002 (N_9002,N_8475,N_8398);
nand U9003 (N_9003,N_8035,N_8685);
nand U9004 (N_9004,N_8693,N_8623);
xor U9005 (N_9005,N_8420,N_8412);
xnor U9006 (N_9006,N_8445,N_8429);
xor U9007 (N_9007,N_8148,N_8196);
and U9008 (N_9008,N_8472,N_8008);
nor U9009 (N_9009,N_8730,N_8443);
or U9010 (N_9010,N_8536,N_8137);
nand U9011 (N_9011,N_8426,N_8171);
nor U9012 (N_9012,N_8774,N_8727);
nor U9013 (N_9013,N_8419,N_8432);
or U9014 (N_9014,N_8257,N_8108);
nand U9015 (N_9015,N_8058,N_8098);
and U9016 (N_9016,N_8360,N_8388);
nor U9017 (N_9017,N_8708,N_8081);
nor U9018 (N_9018,N_8217,N_8295);
xor U9019 (N_9019,N_8768,N_8287);
nand U9020 (N_9020,N_8486,N_8167);
nor U9021 (N_9021,N_8151,N_8092);
xor U9022 (N_9022,N_8506,N_8441);
and U9023 (N_9023,N_8543,N_8754);
nand U9024 (N_9024,N_8501,N_8503);
nand U9025 (N_9025,N_8435,N_8154);
nor U9026 (N_9026,N_8788,N_8455);
nand U9027 (N_9027,N_8540,N_8247);
nand U9028 (N_9028,N_8560,N_8298);
or U9029 (N_9029,N_8766,N_8096);
and U9030 (N_9030,N_8170,N_8751);
nand U9031 (N_9031,N_8112,N_8580);
xor U9032 (N_9032,N_8522,N_8266);
nand U9033 (N_9033,N_8644,N_8499);
and U9034 (N_9034,N_8517,N_8759);
and U9035 (N_9035,N_8208,N_8225);
or U9036 (N_9036,N_8294,N_8645);
nor U9037 (N_9037,N_8018,N_8451);
or U9038 (N_9038,N_8270,N_8775);
xnor U9039 (N_9039,N_8402,N_8565);
xnor U9040 (N_9040,N_8079,N_8738);
or U9041 (N_9041,N_8510,N_8155);
and U9042 (N_9042,N_8456,N_8356);
xor U9043 (N_9043,N_8109,N_8726);
or U9044 (N_9044,N_8405,N_8582);
xnor U9045 (N_9045,N_8066,N_8149);
nand U9046 (N_9046,N_8274,N_8698);
nand U9047 (N_9047,N_8613,N_8080);
nor U9048 (N_9048,N_8668,N_8654);
and U9049 (N_9049,N_8029,N_8700);
nor U9050 (N_9050,N_8621,N_8608);
xnor U9051 (N_9051,N_8702,N_8369);
or U9052 (N_9052,N_8563,N_8619);
or U9053 (N_9053,N_8286,N_8305);
and U9054 (N_9054,N_8704,N_8539);
nor U9055 (N_9055,N_8067,N_8508);
nand U9056 (N_9056,N_8762,N_8387);
and U9057 (N_9057,N_8306,N_8484);
or U9058 (N_9058,N_8555,N_8615);
and U9059 (N_9059,N_8187,N_8778);
nor U9060 (N_9060,N_8597,N_8291);
xor U9061 (N_9061,N_8532,N_8012);
xnor U9062 (N_9062,N_8259,N_8054);
or U9063 (N_9063,N_8683,N_8519);
and U9064 (N_9064,N_8252,N_8316);
xnor U9065 (N_9065,N_8403,N_8584);
and U9066 (N_9066,N_8386,N_8032);
or U9067 (N_9067,N_8415,N_8581);
nor U9068 (N_9068,N_8794,N_8358);
and U9069 (N_9069,N_8500,N_8246);
nand U9070 (N_9070,N_8365,N_8052);
or U9071 (N_9071,N_8566,N_8061);
nand U9072 (N_9072,N_8669,N_8044);
or U9073 (N_9073,N_8713,N_8017);
or U9074 (N_9074,N_8440,N_8476);
nor U9075 (N_9075,N_8351,N_8211);
nand U9076 (N_9076,N_8036,N_8119);
nand U9077 (N_9077,N_8317,N_8168);
and U9078 (N_9078,N_8136,N_8421);
or U9079 (N_9079,N_8466,N_8389);
xor U9080 (N_9080,N_8363,N_8639);
xnor U9081 (N_9081,N_8166,N_8152);
and U9082 (N_9082,N_8195,N_8106);
or U9083 (N_9083,N_8357,N_8350);
and U9084 (N_9084,N_8633,N_8030);
nor U9085 (N_9085,N_8564,N_8488);
nand U9086 (N_9086,N_8408,N_8273);
or U9087 (N_9087,N_8185,N_8093);
or U9088 (N_9088,N_8374,N_8428);
or U9089 (N_9089,N_8188,N_8752);
and U9090 (N_9090,N_8495,N_8300);
or U9091 (N_9091,N_8620,N_8494);
nand U9092 (N_9092,N_8370,N_8753);
xor U9093 (N_9093,N_8013,N_8530);
and U9094 (N_9094,N_8022,N_8750);
or U9095 (N_9095,N_8648,N_8491);
and U9096 (N_9096,N_8705,N_8667);
xor U9097 (N_9097,N_8015,N_8077);
xor U9098 (N_9098,N_8416,N_8272);
nor U9099 (N_9099,N_8205,N_8792);
nor U9100 (N_9100,N_8335,N_8173);
nor U9101 (N_9101,N_8624,N_8016);
nor U9102 (N_9102,N_8622,N_8371);
or U9103 (N_9103,N_8353,N_8561);
xor U9104 (N_9104,N_8544,N_8178);
xnor U9105 (N_9105,N_8465,N_8184);
or U9106 (N_9106,N_8216,N_8028);
nor U9107 (N_9107,N_8733,N_8547);
nand U9108 (N_9108,N_8329,N_8712);
and U9109 (N_9109,N_8064,N_8126);
or U9110 (N_9110,N_8596,N_8323);
nor U9111 (N_9111,N_8436,N_8019);
nor U9112 (N_9112,N_8760,N_8795);
nand U9113 (N_9113,N_8707,N_8050);
xor U9114 (N_9114,N_8586,N_8637);
and U9115 (N_9115,N_8791,N_8599);
xor U9116 (N_9116,N_8399,N_8469);
and U9117 (N_9117,N_8263,N_8347);
nand U9118 (N_9118,N_8395,N_8749);
and U9119 (N_9119,N_8332,N_8602);
nand U9120 (N_9120,N_8046,N_8005);
nor U9121 (N_9121,N_8716,N_8233);
or U9122 (N_9122,N_8192,N_8529);
nand U9123 (N_9123,N_8210,N_8407);
nor U9124 (N_9124,N_8385,N_8575);
xnor U9125 (N_9125,N_8665,N_8593);
or U9126 (N_9126,N_8444,N_8576);
or U9127 (N_9127,N_8534,N_8004);
xnor U9128 (N_9128,N_8143,N_8770);
nand U9129 (N_9129,N_8172,N_8236);
nand U9130 (N_9130,N_8330,N_8604);
nor U9131 (N_9131,N_8100,N_8523);
or U9132 (N_9132,N_8643,N_8769);
or U9133 (N_9133,N_8333,N_8235);
or U9134 (N_9134,N_8493,N_8651);
and U9135 (N_9135,N_8696,N_8011);
nand U9136 (N_9136,N_8000,N_8589);
xnor U9137 (N_9137,N_8786,N_8425);
and U9138 (N_9138,N_8254,N_8203);
or U9139 (N_9139,N_8744,N_8739);
or U9140 (N_9140,N_8742,N_8452);
nand U9141 (N_9141,N_8082,N_8289);
and U9142 (N_9142,N_8722,N_8478);
and U9143 (N_9143,N_8463,N_8745);
nand U9144 (N_9144,N_8740,N_8302);
xor U9145 (N_9145,N_8131,N_8159);
nand U9146 (N_9146,N_8787,N_8796);
nand U9147 (N_9147,N_8303,N_8177);
nand U9148 (N_9148,N_8468,N_8240);
xnor U9149 (N_9149,N_8393,N_8590);
xnor U9150 (N_9150,N_8570,N_8322);
nand U9151 (N_9151,N_8165,N_8142);
and U9152 (N_9152,N_8677,N_8417);
nand U9153 (N_9153,N_8341,N_8422);
nor U9154 (N_9154,N_8232,N_8410);
nor U9155 (N_9155,N_8378,N_8679);
or U9156 (N_9156,N_8438,N_8231);
xor U9157 (N_9157,N_8548,N_8678);
or U9158 (N_9158,N_8141,N_8121);
or U9159 (N_9159,N_8368,N_8720);
nor U9160 (N_9160,N_8201,N_8244);
nand U9161 (N_9161,N_8691,N_8076);
and U9162 (N_9162,N_8676,N_8381);
nor U9163 (N_9163,N_8221,N_8382);
nand U9164 (N_9164,N_8327,N_8262);
nand U9165 (N_9165,N_8113,N_8439);
nand U9166 (N_9166,N_8457,N_8591);
nand U9167 (N_9167,N_8025,N_8537);
nor U9168 (N_9168,N_8174,N_8737);
xor U9169 (N_9169,N_8222,N_8379);
or U9170 (N_9170,N_8521,N_8397);
and U9171 (N_9171,N_8138,N_8448);
or U9172 (N_9172,N_8130,N_8482);
or U9173 (N_9173,N_8336,N_8304);
or U9174 (N_9174,N_8474,N_8377);
or U9175 (N_9175,N_8606,N_8715);
nor U9176 (N_9176,N_8551,N_8513);
or U9177 (N_9177,N_8777,N_8135);
nor U9178 (N_9178,N_8157,N_8647);
nand U9179 (N_9179,N_8346,N_8085);
or U9180 (N_9180,N_8636,N_8057);
nor U9181 (N_9181,N_8139,N_8279);
xor U9182 (N_9182,N_8242,N_8756);
or U9183 (N_9183,N_8666,N_8689);
and U9184 (N_9184,N_8414,N_8784);
nor U9185 (N_9185,N_8735,N_8321);
and U9186 (N_9186,N_8492,N_8163);
and U9187 (N_9187,N_8430,N_8105);
nor U9188 (N_9188,N_8442,N_8115);
nand U9189 (N_9189,N_8318,N_8577);
nand U9190 (N_9190,N_8550,N_8285);
nor U9191 (N_9191,N_8616,N_8611);
and U9192 (N_9192,N_8731,N_8161);
nor U9193 (N_9193,N_8562,N_8271);
xnor U9194 (N_9194,N_8040,N_8186);
xor U9195 (N_9195,N_8260,N_8617);
xor U9196 (N_9196,N_8132,N_8127);
nor U9197 (N_9197,N_8340,N_8505);
and U9198 (N_9198,N_8761,N_8083);
xor U9199 (N_9199,N_8789,N_8743);
nor U9200 (N_9200,N_8554,N_8086);
nor U9201 (N_9201,N_8498,N_8244);
xor U9202 (N_9202,N_8695,N_8396);
and U9203 (N_9203,N_8718,N_8128);
and U9204 (N_9204,N_8257,N_8228);
nand U9205 (N_9205,N_8385,N_8739);
or U9206 (N_9206,N_8615,N_8542);
and U9207 (N_9207,N_8311,N_8486);
or U9208 (N_9208,N_8658,N_8538);
xor U9209 (N_9209,N_8043,N_8425);
xor U9210 (N_9210,N_8723,N_8557);
nor U9211 (N_9211,N_8097,N_8195);
and U9212 (N_9212,N_8257,N_8131);
xnor U9213 (N_9213,N_8296,N_8081);
nor U9214 (N_9214,N_8477,N_8571);
or U9215 (N_9215,N_8029,N_8095);
or U9216 (N_9216,N_8771,N_8172);
or U9217 (N_9217,N_8724,N_8493);
and U9218 (N_9218,N_8033,N_8205);
and U9219 (N_9219,N_8092,N_8601);
nor U9220 (N_9220,N_8307,N_8478);
and U9221 (N_9221,N_8014,N_8376);
xnor U9222 (N_9222,N_8577,N_8394);
and U9223 (N_9223,N_8390,N_8486);
nor U9224 (N_9224,N_8451,N_8558);
xor U9225 (N_9225,N_8237,N_8325);
and U9226 (N_9226,N_8763,N_8741);
xor U9227 (N_9227,N_8517,N_8133);
nand U9228 (N_9228,N_8428,N_8074);
nand U9229 (N_9229,N_8117,N_8647);
nor U9230 (N_9230,N_8786,N_8474);
and U9231 (N_9231,N_8137,N_8621);
nand U9232 (N_9232,N_8254,N_8210);
nor U9233 (N_9233,N_8008,N_8575);
or U9234 (N_9234,N_8716,N_8720);
xor U9235 (N_9235,N_8658,N_8178);
nand U9236 (N_9236,N_8359,N_8759);
xor U9237 (N_9237,N_8387,N_8517);
nor U9238 (N_9238,N_8585,N_8566);
nand U9239 (N_9239,N_8681,N_8572);
nand U9240 (N_9240,N_8390,N_8779);
or U9241 (N_9241,N_8467,N_8256);
nor U9242 (N_9242,N_8622,N_8537);
nand U9243 (N_9243,N_8506,N_8446);
or U9244 (N_9244,N_8281,N_8794);
nand U9245 (N_9245,N_8543,N_8762);
or U9246 (N_9246,N_8788,N_8660);
nor U9247 (N_9247,N_8521,N_8277);
nor U9248 (N_9248,N_8151,N_8655);
nor U9249 (N_9249,N_8425,N_8486);
nand U9250 (N_9250,N_8222,N_8061);
nor U9251 (N_9251,N_8146,N_8733);
nand U9252 (N_9252,N_8077,N_8694);
nand U9253 (N_9253,N_8770,N_8456);
and U9254 (N_9254,N_8470,N_8127);
or U9255 (N_9255,N_8795,N_8532);
xor U9256 (N_9256,N_8557,N_8075);
nor U9257 (N_9257,N_8617,N_8489);
nor U9258 (N_9258,N_8377,N_8429);
nor U9259 (N_9259,N_8748,N_8639);
xor U9260 (N_9260,N_8727,N_8737);
and U9261 (N_9261,N_8507,N_8042);
and U9262 (N_9262,N_8623,N_8135);
and U9263 (N_9263,N_8393,N_8343);
nand U9264 (N_9264,N_8355,N_8168);
nor U9265 (N_9265,N_8094,N_8702);
xnor U9266 (N_9266,N_8346,N_8127);
nand U9267 (N_9267,N_8796,N_8425);
xnor U9268 (N_9268,N_8278,N_8686);
nand U9269 (N_9269,N_8766,N_8397);
nor U9270 (N_9270,N_8563,N_8250);
nand U9271 (N_9271,N_8708,N_8788);
nor U9272 (N_9272,N_8705,N_8225);
or U9273 (N_9273,N_8789,N_8542);
xnor U9274 (N_9274,N_8510,N_8310);
xnor U9275 (N_9275,N_8223,N_8603);
nor U9276 (N_9276,N_8710,N_8678);
or U9277 (N_9277,N_8487,N_8684);
or U9278 (N_9278,N_8519,N_8516);
or U9279 (N_9279,N_8018,N_8604);
and U9280 (N_9280,N_8059,N_8164);
nor U9281 (N_9281,N_8530,N_8249);
or U9282 (N_9282,N_8396,N_8395);
and U9283 (N_9283,N_8205,N_8259);
xor U9284 (N_9284,N_8265,N_8119);
xor U9285 (N_9285,N_8167,N_8093);
nor U9286 (N_9286,N_8301,N_8078);
nor U9287 (N_9287,N_8774,N_8073);
and U9288 (N_9288,N_8307,N_8083);
xnor U9289 (N_9289,N_8183,N_8254);
and U9290 (N_9290,N_8122,N_8202);
nor U9291 (N_9291,N_8059,N_8207);
nor U9292 (N_9292,N_8309,N_8693);
xor U9293 (N_9293,N_8175,N_8188);
nand U9294 (N_9294,N_8256,N_8308);
and U9295 (N_9295,N_8138,N_8686);
and U9296 (N_9296,N_8151,N_8445);
and U9297 (N_9297,N_8539,N_8109);
and U9298 (N_9298,N_8306,N_8424);
nor U9299 (N_9299,N_8099,N_8486);
nor U9300 (N_9300,N_8359,N_8528);
nand U9301 (N_9301,N_8064,N_8794);
xor U9302 (N_9302,N_8294,N_8113);
and U9303 (N_9303,N_8791,N_8351);
or U9304 (N_9304,N_8310,N_8372);
nand U9305 (N_9305,N_8279,N_8067);
or U9306 (N_9306,N_8113,N_8729);
and U9307 (N_9307,N_8316,N_8226);
xnor U9308 (N_9308,N_8061,N_8031);
nand U9309 (N_9309,N_8395,N_8141);
and U9310 (N_9310,N_8099,N_8606);
nand U9311 (N_9311,N_8728,N_8339);
xnor U9312 (N_9312,N_8440,N_8227);
and U9313 (N_9313,N_8612,N_8478);
xor U9314 (N_9314,N_8638,N_8161);
or U9315 (N_9315,N_8121,N_8678);
or U9316 (N_9316,N_8587,N_8657);
and U9317 (N_9317,N_8194,N_8557);
and U9318 (N_9318,N_8227,N_8093);
nand U9319 (N_9319,N_8175,N_8092);
nor U9320 (N_9320,N_8108,N_8028);
nand U9321 (N_9321,N_8547,N_8226);
and U9322 (N_9322,N_8789,N_8773);
nand U9323 (N_9323,N_8496,N_8420);
and U9324 (N_9324,N_8183,N_8355);
or U9325 (N_9325,N_8165,N_8263);
xnor U9326 (N_9326,N_8436,N_8578);
nand U9327 (N_9327,N_8209,N_8550);
or U9328 (N_9328,N_8481,N_8605);
xor U9329 (N_9329,N_8281,N_8783);
and U9330 (N_9330,N_8509,N_8149);
xor U9331 (N_9331,N_8566,N_8795);
xor U9332 (N_9332,N_8443,N_8088);
and U9333 (N_9333,N_8326,N_8518);
and U9334 (N_9334,N_8215,N_8468);
nand U9335 (N_9335,N_8362,N_8650);
or U9336 (N_9336,N_8074,N_8588);
nand U9337 (N_9337,N_8594,N_8390);
nand U9338 (N_9338,N_8390,N_8666);
nand U9339 (N_9339,N_8219,N_8069);
nor U9340 (N_9340,N_8623,N_8195);
nand U9341 (N_9341,N_8719,N_8170);
and U9342 (N_9342,N_8472,N_8673);
or U9343 (N_9343,N_8799,N_8556);
nor U9344 (N_9344,N_8792,N_8215);
and U9345 (N_9345,N_8004,N_8409);
or U9346 (N_9346,N_8049,N_8025);
and U9347 (N_9347,N_8795,N_8584);
xnor U9348 (N_9348,N_8701,N_8322);
and U9349 (N_9349,N_8164,N_8578);
nor U9350 (N_9350,N_8426,N_8629);
xor U9351 (N_9351,N_8184,N_8062);
and U9352 (N_9352,N_8063,N_8755);
xnor U9353 (N_9353,N_8798,N_8337);
xnor U9354 (N_9354,N_8207,N_8068);
or U9355 (N_9355,N_8596,N_8368);
nand U9356 (N_9356,N_8399,N_8560);
or U9357 (N_9357,N_8328,N_8082);
or U9358 (N_9358,N_8209,N_8774);
nand U9359 (N_9359,N_8499,N_8443);
nand U9360 (N_9360,N_8736,N_8214);
xor U9361 (N_9361,N_8453,N_8590);
or U9362 (N_9362,N_8227,N_8242);
and U9363 (N_9363,N_8763,N_8181);
or U9364 (N_9364,N_8472,N_8410);
and U9365 (N_9365,N_8427,N_8135);
xnor U9366 (N_9366,N_8143,N_8268);
nand U9367 (N_9367,N_8245,N_8531);
and U9368 (N_9368,N_8419,N_8301);
xnor U9369 (N_9369,N_8131,N_8368);
or U9370 (N_9370,N_8075,N_8226);
nand U9371 (N_9371,N_8173,N_8677);
nor U9372 (N_9372,N_8403,N_8772);
nor U9373 (N_9373,N_8145,N_8449);
nand U9374 (N_9374,N_8646,N_8733);
nand U9375 (N_9375,N_8792,N_8542);
xor U9376 (N_9376,N_8278,N_8408);
or U9377 (N_9377,N_8003,N_8747);
and U9378 (N_9378,N_8327,N_8663);
nor U9379 (N_9379,N_8442,N_8586);
and U9380 (N_9380,N_8706,N_8387);
nor U9381 (N_9381,N_8164,N_8070);
or U9382 (N_9382,N_8430,N_8716);
nor U9383 (N_9383,N_8285,N_8499);
nand U9384 (N_9384,N_8735,N_8220);
nor U9385 (N_9385,N_8399,N_8405);
or U9386 (N_9386,N_8386,N_8004);
and U9387 (N_9387,N_8233,N_8331);
nor U9388 (N_9388,N_8514,N_8598);
or U9389 (N_9389,N_8097,N_8153);
and U9390 (N_9390,N_8366,N_8536);
xnor U9391 (N_9391,N_8268,N_8643);
or U9392 (N_9392,N_8073,N_8472);
or U9393 (N_9393,N_8627,N_8198);
and U9394 (N_9394,N_8797,N_8570);
xor U9395 (N_9395,N_8771,N_8138);
and U9396 (N_9396,N_8121,N_8081);
xor U9397 (N_9397,N_8553,N_8127);
and U9398 (N_9398,N_8024,N_8787);
xor U9399 (N_9399,N_8581,N_8503);
and U9400 (N_9400,N_8713,N_8075);
or U9401 (N_9401,N_8119,N_8370);
nand U9402 (N_9402,N_8456,N_8434);
nand U9403 (N_9403,N_8642,N_8128);
nand U9404 (N_9404,N_8334,N_8444);
nor U9405 (N_9405,N_8362,N_8329);
or U9406 (N_9406,N_8203,N_8475);
xnor U9407 (N_9407,N_8058,N_8061);
and U9408 (N_9408,N_8023,N_8774);
nand U9409 (N_9409,N_8496,N_8464);
nand U9410 (N_9410,N_8561,N_8145);
nor U9411 (N_9411,N_8095,N_8134);
xor U9412 (N_9412,N_8701,N_8478);
and U9413 (N_9413,N_8699,N_8694);
xnor U9414 (N_9414,N_8026,N_8507);
or U9415 (N_9415,N_8478,N_8134);
nand U9416 (N_9416,N_8202,N_8150);
and U9417 (N_9417,N_8789,N_8114);
and U9418 (N_9418,N_8554,N_8462);
nor U9419 (N_9419,N_8377,N_8307);
nor U9420 (N_9420,N_8453,N_8579);
and U9421 (N_9421,N_8750,N_8573);
nor U9422 (N_9422,N_8342,N_8670);
nor U9423 (N_9423,N_8367,N_8110);
or U9424 (N_9424,N_8292,N_8795);
and U9425 (N_9425,N_8476,N_8540);
nor U9426 (N_9426,N_8023,N_8682);
xor U9427 (N_9427,N_8441,N_8091);
or U9428 (N_9428,N_8094,N_8738);
nor U9429 (N_9429,N_8458,N_8165);
and U9430 (N_9430,N_8319,N_8431);
or U9431 (N_9431,N_8020,N_8488);
and U9432 (N_9432,N_8584,N_8229);
and U9433 (N_9433,N_8734,N_8103);
or U9434 (N_9434,N_8105,N_8142);
or U9435 (N_9435,N_8114,N_8032);
xnor U9436 (N_9436,N_8471,N_8414);
xnor U9437 (N_9437,N_8057,N_8407);
xor U9438 (N_9438,N_8426,N_8003);
and U9439 (N_9439,N_8222,N_8195);
or U9440 (N_9440,N_8520,N_8009);
xor U9441 (N_9441,N_8515,N_8242);
xor U9442 (N_9442,N_8206,N_8132);
xor U9443 (N_9443,N_8195,N_8780);
or U9444 (N_9444,N_8475,N_8406);
nand U9445 (N_9445,N_8216,N_8588);
or U9446 (N_9446,N_8054,N_8250);
or U9447 (N_9447,N_8119,N_8153);
xnor U9448 (N_9448,N_8589,N_8426);
and U9449 (N_9449,N_8166,N_8487);
nand U9450 (N_9450,N_8389,N_8313);
xor U9451 (N_9451,N_8345,N_8505);
nor U9452 (N_9452,N_8333,N_8373);
nor U9453 (N_9453,N_8273,N_8087);
nor U9454 (N_9454,N_8709,N_8092);
and U9455 (N_9455,N_8772,N_8006);
nand U9456 (N_9456,N_8440,N_8570);
nand U9457 (N_9457,N_8070,N_8598);
and U9458 (N_9458,N_8145,N_8152);
xor U9459 (N_9459,N_8163,N_8222);
or U9460 (N_9460,N_8394,N_8425);
nand U9461 (N_9461,N_8051,N_8336);
nor U9462 (N_9462,N_8057,N_8111);
xnor U9463 (N_9463,N_8209,N_8777);
xnor U9464 (N_9464,N_8250,N_8023);
xor U9465 (N_9465,N_8624,N_8600);
and U9466 (N_9466,N_8222,N_8054);
xnor U9467 (N_9467,N_8659,N_8227);
nor U9468 (N_9468,N_8627,N_8783);
xor U9469 (N_9469,N_8133,N_8597);
nor U9470 (N_9470,N_8715,N_8094);
or U9471 (N_9471,N_8349,N_8655);
nand U9472 (N_9472,N_8130,N_8572);
nand U9473 (N_9473,N_8523,N_8106);
xor U9474 (N_9474,N_8265,N_8597);
or U9475 (N_9475,N_8419,N_8360);
xor U9476 (N_9476,N_8592,N_8193);
nor U9477 (N_9477,N_8432,N_8324);
nand U9478 (N_9478,N_8521,N_8704);
nor U9479 (N_9479,N_8113,N_8678);
and U9480 (N_9480,N_8348,N_8646);
nand U9481 (N_9481,N_8696,N_8369);
and U9482 (N_9482,N_8236,N_8303);
nor U9483 (N_9483,N_8615,N_8116);
nor U9484 (N_9484,N_8465,N_8723);
or U9485 (N_9485,N_8126,N_8523);
or U9486 (N_9486,N_8715,N_8179);
nand U9487 (N_9487,N_8402,N_8791);
or U9488 (N_9488,N_8098,N_8509);
and U9489 (N_9489,N_8314,N_8362);
nor U9490 (N_9490,N_8211,N_8353);
xnor U9491 (N_9491,N_8027,N_8378);
and U9492 (N_9492,N_8545,N_8245);
xnor U9493 (N_9493,N_8694,N_8613);
and U9494 (N_9494,N_8747,N_8378);
nand U9495 (N_9495,N_8703,N_8372);
nand U9496 (N_9496,N_8654,N_8603);
nand U9497 (N_9497,N_8211,N_8136);
and U9498 (N_9498,N_8476,N_8720);
xnor U9499 (N_9499,N_8768,N_8555);
nor U9500 (N_9500,N_8196,N_8382);
xor U9501 (N_9501,N_8618,N_8093);
nand U9502 (N_9502,N_8459,N_8170);
and U9503 (N_9503,N_8542,N_8658);
xor U9504 (N_9504,N_8549,N_8358);
and U9505 (N_9505,N_8696,N_8231);
and U9506 (N_9506,N_8732,N_8124);
or U9507 (N_9507,N_8298,N_8202);
xnor U9508 (N_9508,N_8141,N_8521);
or U9509 (N_9509,N_8000,N_8270);
and U9510 (N_9510,N_8690,N_8497);
nor U9511 (N_9511,N_8121,N_8016);
xnor U9512 (N_9512,N_8064,N_8524);
nor U9513 (N_9513,N_8542,N_8459);
nor U9514 (N_9514,N_8333,N_8606);
and U9515 (N_9515,N_8141,N_8712);
and U9516 (N_9516,N_8723,N_8207);
and U9517 (N_9517,N_8104,N_8161);
nand U9518 (N_9518,N_8206,N_8462);
or U9519 (N_9519,N_8617,N_8187);
and U9520 (N_9520,N_8636,N_8342);
or U9521 (N_9521,N_8212,N_8768);
and U9522 (N_9522,N_8533,N_8252);
nor U9523 (N_9523,N_8730,N_8158);
nand U9524 (N_9524,N_8457,N_8125);
and U9525 (N_9525,N_8260,N_8544);
or U9526 (N_9526,N_8535,N_8136);
and U9527 (N_9527,N_8077,N_8689);
nor U9528 (N_9528,N_8627,N_8692);
and U9529 (N_9529,N_8660,N_8588);
and U9530 (N_9530,N_8715,N_8244);
and U9531 (N_9531,N_8442,N_8229);
or U9532 (N_9532,N_8430,N_8627);
nand U9533 (N_9533,N_8434,N_8193);
nand U9534 (N_9534,N_8481,N_8648);
nand U9535 (N_9535,N_8455,N_8364);
or U9536 (N_9536,N_8618,N_8697);
nor U9537 (N_9537,N_8707,N_8486);
xor U9538 (N_9538,N_8542,N_8683);
nand U9539 (N_9539,N_8659,N_8793);
nor U9540 (N_9540,N_8384,N_8588);
nor U9541 (N_9541,N_8435,N_8567);
or U9542 (N_9542,N_8488,N_8469);
xnor U9543 (N_9543,N_8744,N_8404);
and U9544 (N_9544,N_8477,N_8292);
nor U9545 (N_9545,N_8336,N_8061);
nand U9546 (N_9546,N_8382,N_8593);
or U9547 (N_9547,N_8385,N_8711);
xor U9548 (N_9548,N_8098,N_8029);
and U9549 (N_9549,N_8128,N_8154);
and U9550 (N_9550,N_8526,N_8225);
xor U9551 (N_9551,N_8224,N_8079);
or U9552 (N_9552,N_8699,N_8337);
nor U9553 (N_9553,N_8418,N_8769);
and U9554 (N_9554,N_8591,N_8006);
or U9555 (N_9555,N_8328,N_8199);
nor U9556 (N_9556,N_8272,N_8685);
nand U9557 (N_9557,N_8131,N_8434);
and U9558 (N_9558,N_8780,N_8574);
xnor U9559 (N_9559,N_8145,N_8731);
nand U9560 (N_9560,N_8388,N_8232);
nor U9561 (N_9561,N_8170,N_8599);
nor U9562 (N_9562,N_8101,N_8673);
and U9563 (N_9563,N_8162,N_8675);
nor U9564 (N_9564,N_8505,N_8695);
nor U9565 (N_9565,N_8445,N_8269);
and U9566 (N_9566,N_8798,N_8787);
xor U9567 (N_9567,N_8324,N_8263);
or U9568 (N_9568,N_8431,N_8673);
nand U9569 (N_9569,N_8263,N_8127);
nand U9570 (N_9570,N_8256,N_8500);
nor U9571 (N_9571,N_8664,N_8316);
nor U9572 (N_9572,N_8319,N_8171);
or U9573 (N_9573,N_8706,N_8557);
and U9574 (N_9574,N_8318,N_8540);
or U9575 (N_9575,N_8147,N_8413);
nand U9576 (N_9576,N_8066,N_8318);
or U9577 (N_9577,N_8347,N_8771);
and U9578 (N_9578,N_8539,N_8137);
and U9579 (N_9579,N_8010,N_8492);
nand U9580 (N_9580,N_8191,N_8759);
nand U9581 (N_9581,N_8022,N_8468);
and U9582 (N_9582,N_8638,N_8580);
nand U9583 (N_9583,N_8627,N_8042);
or U9584 (N_9584,N_8652,N_8434);
nor U9585 (N_9585,N_8686,N_8129);
nor U9586 (N_9586,N_8502,N_8567);
and U9587 (N_9587,N_8624,N_8711);
nor U9588 (N_9588,N_8646,N_8202);
nand U9589 (N_9589,N_8721,N_8355);
nor U9590 (N_9590,N_8699,N_8207);
nor U9591 (N_9591,N_8010,N_8638);
or U9592 (N_9592,N_8508,N_8691);
nor U9593 (N_9593,N_8566,N_8767);
and U9594 (N_9594,N_8711,N_8018);
nor U9595 (N_9595,N_8122,N_8551);
xor U9596 (N_9596,N_8787,N_8246);
nor U9597 (N_9597,N_8652,N_8207);
xnor U9598 (N_9598,N_8309,N_8000);
xnor U9599 (N_9599,N_8756,N_8263);
and U9600 (N_9600,N_9264,N_9528);
xor U9601 (N_9601,N_8856,N_9541);
or U9602 (N_9602,N_8937,N_9148);
nor U9603 (N_9603,N_9293,N_9575);
nor U9604 (N_9604,N_8851,N_9563);
nand U9605 (N_9605,N_9046,N_9042);
or U9606 (N_9606,N_8849,N_9223);
nand U9607 (N_9607,N_9292,N_9159);
nand U9608 (N_9608,N_9319,N_9192);
or U9609 (N_9609,N_9572,N_9087);
and U9610 (N_9610,N_9463,N_9442);
and U9611 (N_9611,N_9137,N_8811);
nor U9612 (N_9612,N_9581,N_9305);
nor U9613 (N_9613,N_9418,N_9100);
or U9614 (N_9614,N_8987,N_9451);
nor U9615 (N_9615,N_9150,N_9152);
and U9616 (N_9616,N_9465,N_9124);
and U9617 (N_9617,N_8928,N_9249);
nor U9618 (N_9618,N_9111,N_8879);
nand U9619 (N_9619,N_9332,N_9545);
xor U9620 (N_9620,N_9199,N_9445);
nand U9621 (N_9621,N_8877,N_9509);
nor U9622 (N_9622,N_9547,N_9382);
or U9623 (N_9623,N_8907,N_8920);
nand U9624 (N_9624,N_9561,N_9256);
nand U9625 (N_9625,N_9096,N_9306);
or U9626 (N_9626,N_9439,N_8857);
nand U9627 (N_9627,N_9025,N_9140);
and U9628 (N_9628,N_9379,N_9433);
nand U9629 (N_9629,N_9404,N_8847);
nor U9630 (N_9630,N_9540,N_9432);
xnor U9631 (N_9631,N_8986,N_8927);
or U9632 (N_9632,N_9053,N_9513);
and U9633 (N_9633,N_9403,N_9226);
and U9634 (N_9634,N_9061,N_9551);
or U9635 (N_9635,N_9333,N_9274);
and U9636 (N_9636,N_9119,N_9109);
or U9637 (N_9637,N_9479,N_8959);
and U9638 (N_9638,N_8824,N_8969);
nand U9639 (N_9639,N_9452,N_9268);
nand U9640 (N_9640,N_8974,N_9434);
nor U9641 (N_9641,N_9136,N_9019);
nor U9642 (N_9642,N_9212,N_9207);
and U9643 (N_9643,N_8806,N_9459);
or U9644 (N_9644,N_9000,N_8819);
nor U9645 (N_9645,N_8924,N_9176);
or U9646 (N_9646,N_9084,N_9060);
nand U9647 (N_9647,N_8930,N_9098);
and U9648 (N_9648,N_8809,N_9191);
nand U9649 (N_9649,N_9486,N_8834);
xnor U9650 (N_9650,N_9118,N_9393);
and U9651 (N_9651,N_9255,N_9466);
xnor U9652 (N_9652,N_9353,N_9038);
or U9653 (N_9653,N_9090,N_9067);
xnor U9654 (N_9654,N_8844,N_9056);
xor U9655 (N_9655,N_9591,N_9010);
nor U9656 (N_9656,N_9055,N_9394);
xnor U9657 (N_9657,N_9162,N_8801);
or U9658 (N_9658,N_9088,N_8925);
and U9659 (N_9659,N_9473,N_9033);
nor U9660 (N_9660,N_9361,N_9184);
nor U9661 (N_9661,N_9504,N_8982);
nand U9662 (N_9662,N_9027,N_9216);
and U9663 (N_9663,N_9475,N_8983);
or U9664 (N_9664,N_9105,N_9555);
xnor U9665 (N_9665,N_9230,N_9328);
nor U9666 (N_9666,N_9101,N_9001);
or U9667 (N_9667,N_9064,N_8873);
xor U9668 (N_9668,N_9251,N_8871);
nor U9669 (N_9669,N_8945,N_9126);
or U9670 (N_9670,N_9458,N_9533);
nand U9671 (N_9671,N_9344,N_9596);
xnor U9672 (N_9672,N_9576,N_8971);
xor U9673 (N_9673,N_9558,N_9133);
and U9674 (N_9674,N_9356,N_9171);
xor U9675 (N_9675,N_8966,N_9594);
and U9676 (N_9676,N_9254,N_8999);
or U9677 (N_9677,N_8996,N_9435);
and U9678 (N_9678,N_9303,N_9089);
nor U9679 (N_9679,N_9349,N_9099);
nor U9680 (N_9680,N_9320,N_9343);
or U9681 (N_9681,N_9494,N_8965);
nor U9682 (N_9682,N_9085,N_8916);
and U9683 (N_9683,N_8848,N_9075);
xor U9684 (N_9684,N_8821,N_9104);
nor U9685 (N_9685,N_9235,N_8805);
or U9686 (N_9686,N_9009,N_9302);
and U9687 (N_9687,N_9011,N_9414);
xnor U9688 (N_9688,N_9143,N_9441);
nand U9689 (N_9689,N_9566,N_9386);
xor U9690 (N_9690,N_9492,N_9263);
or U9691 (N_9691,N_9097,N_9059);
or U9692 (N_9692,N_9573,N_9266);
nor U9693 (N_9693,N_9275,N_9321);
nand U9694 (N_9694,N_9290,N_9543);
nor U9695 (N_9695,N_8880,N_9440);
or U9696 (N_9696,N_9447,N_8929);
and U9697 (N_9697,N_8872,N_8894);
xor U9698 (N_9698,N_9122,N_9195);
nand U9699 (N_9699,N_9174,N_8935);
and U9700 (N_9700,N_9093,N_9318);
xor U9701 (N_9701,N_9265,N_9490);
xor U9702 (N_9702,N_8828,N_9311);
nand U9703 (N_9703,N_9175,N_9078);
nor U9704 (N_9704,N_9052,N_9516);
nor U9705 (N_9705,N_8886,N_8903);
xnor U9706 (N_9706,N_9051,N_9366);
and U9707 (N_9707,N_9076,N_9301);
xor U9708 (N_9708,N_9429,N_8957);
xor U9709 (N_9709,N_9242,N_9187);
nand U9710 (N_9710,N_8829,N_9383);
xor U9711 (N_9711,N_9161,N_9388);
nand U9712 (N_9712,N_9233,N_8818);
xnor U9713 (N_9713,N_9347,N_9385);
or U9714 (N_9714,N_8850,N_9431);
nor U9715 (N_9715,N_9471,N_9583);
and U9716 (N_9716,N_9579,N_9172);
nand U9717 (N_9717,N_9125,N_9449);
xnor U9718 (N_9718,N_9525,N_9364);
and U9719 (N_9719,N_9080,N_9548);
nor U9720 (N_9720,N_8901,N_9337);
and U9721 (N_9721,N_9021,N_9428);
nand U9722 (N_9722,N_9163,N_8909);
nand U9723 (N_9723,N_9003,N_9495);
and U9724 (N_9724,N_8897,N_9094);
xnor U9725 (N_9725,N_9367,N_9106);
and U9726 (N_9726,N_8960,N_9308);
nor U9727 (N_9727,N_9049,N_9210);
or U9728 (N_9728,N_9584,N_9063);
nand U9729 (N_9729,N_8963,N_9316);
or U9730 (N_9730,N_8931,N_8970);
xor U9731 (N_9731,N_9557,N_8917);
xor U9732 (N_9732,N_9198,N_8853);
nand U9733 (N_9733,N_9348,N_9299);
and U9734 (N_9734,N_9546,N_8979);
nand U9735 (N_9735,N_9219,N_9443);
xor U9736 (N_9736,N_9240,N_9484);
nand U9737 (N_9737,N_9376,N_9043);
nand U9738 (N_9738,N_8878,N_9598);
nand U9739 (N_9739,N_9149,N_9399);
nor U9740 (N_9740,N_9342,N_9472);
nand U9741 (N_9741,N_8993,N_9352);
nand U9742 (N_9742,N_9208,N_9520);
nor U9743 (N_9743,N_8947,N_9396);
xnor U9744 (N_9744,N_9156,N_9582);
nand U9745 (N_9745,N_9389,N_9327);
nor U9746 (N_9746,N_9325,N_9204);
or U9747 (N_9747,N_9410,N_9196);
nand U9748 (N_9748,N_8890,N_9023);
nor U9749 (N_9749,N_9438,N_9411);
or U9750 (N_9750,N_9006,N_9565);
or U9751 (N_9751,N_9539,N_9496);
nand U9752 (N_9752,N_9017,N_9151);
or U9753 (N_9753,N_9568,N_9331);
and U9754 (N_9754,N_9530,N_8949);
and U9755 (N_9755,N_9298,N_9026);
and U9756 (N_9756,N_9322,N_9483);
and U9757 (N_9757,N_9036,N_8923);
nor U9758 (N_9758,N_9229,N_9368);
or U9759 (N_9759,N_8833,N_9487);
xnor U9760 (N_9760,N_9559,N_9534);
xor U9761 (N_9761,N_8898,N_8817);
nor U9762 (N_9762,N_9564,N_9467);
and U9763 (N_9763,N_8899,N_8842);
nor U9764 (N_9764,N_9423,N_8922);
xnor U9765 (N_9765,N_9135,N_9280);
xnor U9766 (N_9766,N_8865,N_9307);
and U9767 (N_9767,N_9120,N_8938);
nand U9768 (N_9768,N_9228,N_9567);
xnor U9769 (N_9769,N_9419,N_8860);
nor U9770 (N_9770,N_9339,N_9008);
or U9771 (N_9771,N_8889,N_9296);
xor U9772 (N_9772,N_9477,N_9515);
or U9773 (N_9773,N_9340,N_9514);
or U9774 (N_9774,N_9107,N_9247);
or U9775 (N_9775,N_9497,N_9574);
nand U9776 (N_9776,N_9138,N_9358);
nor U9777 (N_9777,N_9044,N_9341);
nor U9778 (N_9778,N_9571,N_9128);
and U9779 (N_9779,N_9217,N_9532);
nor U9780 (N_9780,N_8883,N_9409);
xnor U9781 (N_9781,N_9020,N_8952);
xor U9782 (N_9782,N_9457,N_9529);
xor U9783 (N_9783,N_9164,N_9370);
nor U9784 (N_9784,N_9456,N_8958);
and U9785 (N_9785,N_8837,N_9057);
and U9786 (N_9786,N_9374,N_9271);
nor U9787 (N_9787,N_9500,N_8845);
nor U9788 (N_9788,N_9554,N_8951);
and U9789 (N_9789,N_9170,N_9335);
and U9790 (N_9790,N_8998,N_9489);
or U9791 (N_9791,N_9518,N_9326);
xor U9792 (N_9792,N_9276,N_9593);
xor U9793 (N_9793,N_9365,N_9521);
xnor U9794 (N_9794,N_9315,N_9549);
and U9795 (N_9795,N_9362,N_8825);
nor U9796 (N_9796,N_9082,N_9167);
nand U9797 (N_9797,N_8956,N_9405);
xnor U9798 (N_9798,N_9508,N_8841);
nand U9799 (N_9799,N_8985,N_9194);
or U9800 (N_9800,N_8862,N_9517);
nor U9801 (N_9801,N_9544,N_9536);
xnor U9802 (N_9802,N_9130,N_9157);
and U9803 (N_9803,N_8940,N_9197);
and U9804 (N_9804,N_9113,N_9160);
nand U9805 (N_9805,N_9232,N_9189);
nand U9806 (N_9806,N_9589,N_9039);
nand U9807 (N_9807,N_9373,N_9202);
nand U9808 (N_9808,N_9166,N_9185);
or U9809 (N_9809,N_8968,N_9421);
and U9810 (N_9810,N_8888,N_9338);
nand U9811 (N_9811,N_9372,N_9560);
nor U9812 (N_9812,N_9193,N_9336);
and U9813 (N_9813,N_9453,N_8926);
nand U9814 (N_9814,N_8975,N_9273);
xnor U9815 (N_9815,N_9015,N_8904);
or U9816 (N_9816,N_9597,N_9523);
nand U9817 (N_9817,N_9054,N_8864);
xor U9818 (N_9818,N_9289,N_8911);
nand U9819 (N_9819,N_9464,N_9310);
nand U9820 (N_9820,N_8918,N_9079);
and U9821 (N_9821,N_9115,N_8946);
nor U9822 (N_9822,N_9499,N_9129);
or U9823 (N_9823,N_8830,N_9522);
and U9824 (N_9824,N_9103,N_9121);
or U9825 (N_9825,N_9278,N_9281);
nor U9826 (N_9826,N_9324,N_9218);
and U9827 (N_9827,N_9201,N_9312);
xor U9828 (N_9828,N_9236,N_9144);
or U9829 (N_9829,N_9422,N_9040);
or U9830 (N_9830,N_8870,N_9016);
and U9831 (N_9831,N_8816,N_9070);
nand U9832 (N_9832,N_9114,N_9139);
nor U9833 (N_9833,N_9297,N_9012);
xor U9834 (N_9834,N_9412,N_9200);
nor U9835 (N_9835,N_9165,N_9578);
or U9836 (N_9836,N_9260,N_9291);
and U9837 (N_9837,N_9213,N_9183);
and U9838 (N_9838,N_8984,N_9041);
nor U9839 (N_9839,N_9351,N_8964);
nand U9840 (N_9840,N_8896,N_9110);
and U9841 (N_9841,N_8827,N_9004);
nand U9842 (N_9842,N_8895,N_8990);
and U9843 (N_9843,N_9408,N_9127);
or U9844 (N_9844,N_8912,N_9285);
nand U9845 (N_9845,N_8815,N_9267);
nor U9846 (N_9846,N_9317,N_8954);
xnor U9847 (N_9847,N_9346,N_9030);
nor U9848 (N_9848,N_9224,N_9482);
nor U9849 (N_9849,N_9397,N_9527);
xnor U9850 (N_9850,N_8915,N_9550);
and U9851 (N_9851,N_9182,N_9493);
nor U9852 (N_9852,N_9173,N_9444);
xor U9853 (N_9853,N_8866,N_9415);
and U9854 (N_9854,N_9569,N_9214);
xor U9855 (N_9855,N_9225,N_9014);
nor U9856 (N_9856,N_9243,N_9047);
or U9857 (N_9857,N_9430,N_9398);
or U9858 (N_9858,N_9220,N_8800);
xnor U9859 (N_9859,N_9269,N_9417);
xnor U9860 (N_9860,N_8942,N_8855);
xnor U9861 (N_9861,N_9360,N_9245);
and U9862 (N_9862,N_9154,N_9024);
or U9863 (N_9863,N_8826,N_9425);
and U9864 (N_9864,N_9380,N_9313);
nor U9865 (N_9865,N_9227,N_8835);
or U9866 (N_9866,N_8981,N_8997);
nor U9867 (N_9867,N_9270,N_9186);
nor U9868 (N_9868,N_9553,N_9277);
nand U9869 (N_9869,N_8939,N_8876);
xnor U9870 (N_9870,N_9580,N_8944);
nor U9871 (N_9871,N_9519,N_9446);
nor U9872 (N_9872,N_9588,N_8914);
or U9873 (N_9873,N_9304,N_9436);
or U9874 (N_9874,N_9329,N_9209);
nand U9875 (N_9875,N_9460,N_9145);
xor U9876 (N_9876,N_9205,N_8967);
xnor U9877 (N_9877,N_9034,N_9248);
and U9878 (N_9878,N_9142,N_9424);
or U9879 (N_9879,N_9141,N_9381);
nand U9880 (N_9880,N_9354,N_9116);
nor U9881 (N_9881,N_9112,N_9476);
nor U9882 (N_9882,N_8989,N_9506);
or U9883 (N_9883,N_9037,N_9512);
nand U9884 (N_9884,N_9032,N_9066);
xnor U9885 (N_9885,N_9179,N_8859);
nor U9886 (N_9886,N_9002,N_8995);
nor U9887 (N_9887,N_9158,N_9203);
nor U9888 (N_9888,N_9083,N_8988);
or U9889 (N_9889,N_9045,N_9314);
or U9890 (N_9890,N_8803,N_9524);
xor U9891 (N_9891,N_8980,N_9402);
or U9892 (N_9892,N_9416,N_9287);
and U9893 (N_9893,N_8900,N_9074);
or U9894 (N_9894,N_9180,N_8802);
xnor U9895 (N_9895,N_9284,N_9062);
or U9896 (N_9896,N_9146,N_9468);
nand U9897 (N_9897,N_9065,N_8910);
nor U9898 (N_9898,N_8863,N_9252);
nand U9899 (N_9899,N_9234,N_9272);
xor U9900 (N_9900,N_8955,N_9221);
nand U9901 (N_9901,N_9590,N_9108);
nor U9902 (N_9902,N_9359,N_9369);
nand U9903 (N_9903,N_8902,N_9131);
nor U9904 (N_9904,N_8936,N_9363);
nand U9905 (N_9905,N_9510,N_9309);
and U9906 (N_9906,N_8831,N_9448);
nand U9907 (N_9907,N_9538,N_8961);
nor U9908 (N_9908,N_9502,N_9384);
and U9909 (N_9909,N_8881,N_9022);
nand U9910 (N_9910,N_8932,N_9585);
nor U9911 (N_9911,N_8822,N_9387);
and U9912 (N_9912,N_9237,N_8994);
xor U9913 (N_9913,N_9095,N_9259);
xnor U9914 (N_9914,N_9537,N_8973);
nand U9915 (N_9915,N_9241,N_9029);
or U9916 (N_9916,N_9013,N_9587);
xor U9917 (N_9917,N_9007,N_8823);
nand U9918 (N_9918,N_9406,N_9028);
nor U9919 (N_9919,N_9262,N_8977);
and U9920 (N_9920,N_9031,N_9153);
nor U9921 (N_9921,N_9295,N_9222);
nand U9922 (N_9922,N_9599,N_9050);
nand U9923 (N_9923,N_9155,N_9378);
and U9924 (N_9924,N_8934,N_9211);
xnor U9925 (N_9925,N_8906,N_8852);
nor U9926 (N_9926,N_9392,N_9592);
or U9927 (N_9927,N_9261,N_9371);
nand U9928 (N_9928,N_8813,N_8808);
or U9929 (N_9929,N_8962,N_9117);
and U9930 (N_9930,N_8991,N_9562);
nor U9931 (N_9931,N_8908,N_9058);
or U9932 (N_9932,N_9505,N_9491);
nand U9933 (N_9933,N_9355,N_8885);
and U9934 (N_9934,N_9068,N_8913);
and U9935 (N_9935,N_9407,N_8943);
or U9936 (N_9936,N_9257,N_9420);
or U9937 (N_9937,N_9427,N_9330);
nand U9938 (N_9938,N_9488,N_9102);
nor U9939 (N_9939,N_8804,N_8992);
or U9940 (N_9940,N_9258,N_9570);
nand U9941 (N_9941,N_8814,N_9474);
or U9942 (N_9942,N_9426,N_9526);
nor U9943 (N_9943,N_8868,N_8861);
or U9944 (N_9944,N_9239,N_9511);
nor U9945 (N_9945,N_9461,N_9071);
xor U9946 (N_9946,N_9178,N_9215);
and U9947 (N_9947,N_9577,N_9413);
xor U9948 (N_9948,N_8838,N_8948);
nor U9949 (N_9949,N_9238,N_9470);
nand U9950 (N_9950,N_8846,N_9188);
or U9951 (N_9951,N_9244,N_9134);
nor U9952 (N_9952,N_9345,N_8858);
and U9953 (N_9953,N_9390,N_9231);
or U9954 (N_9954,N_9190,N_9350);
nor U9955 (N_9955,N_8921,N_8869);
or U9956 (N_9956,N_9123,N_9206);
and U9957 (N_9957,N_8953,N_8905);
nor U9958 (N_9958,N_9288,N_8972);
and U9959 (N_9959,N_8887,N_8978);
and U9960 (N_9960,N_8941,N_9503);
nand U9961 (N_9961,N_9253,N_9531);
nand U9962 (N_9962,N_9552,N_9073);
xnor U9963 (N_9963,N_8836,N_9279);
xnor U9964 (N_9964,N_9455,N_8839);
nor U9965 (N_9965,N_8976,N_9294);
and U9966 (N_9966,N_9334,N_8840);
nand U9967 (N_9967,N_8812,N_9454);
or U9968 (N_9968,N_9069,N_8874);
or U9969 (N_9969,N_8882,N_9485);
nand U9970 (N_9970,N_8892,N_9081);
nor U9971 (N_9971,N_9147,N_8807);
and U9972 (N_9972,N_9048,N_8820);
or U9973 (N_9973,N_8933,N_9091);
or U9974 (N_9974,N_9072,N_9556);
nand U9975 (N_9975,N_9168,N_9501);
and U9976 (N_9976,N_9250,N_9498);
nor U9977 (N_9977,N_9450,N_9286);
or U9978 (N_9978,N_9469,N_9086);
and U9979 (N_9979,N_9401,N_9478);
xor U9980 (N_9980,N_8950,N_9375);
nor U9981 (N_9981,N_8893,N_8919);
xor U9982 (N_9982,N_9462,N_8854);
nand U9983 (N_9983,N_9400,N_9391);
nand U9984 (N_9984,N_9507,N_9480);
and U9985 (N_9985,N_9181,N_9092);
xor U9986 (N_9986,N_9357,N_8875);
nand U9987 (N_9987,N_8832,N_9377);
nand U9988 (N_9988,N_8867,N_9323);
xor U9989 (N_9989,N_9246,N_9586);
nor U9990 (N_9990,N_9395,N_8884);
nand U9991 (N_9991,N_8810,N_9300);
nand U9992 (N_9992,N_9283,N_9481);
or U9993 (N_9993,N_9535,N_9132);
or U9994 (N_9994,N_9437,N_9282);
or U9995 (N_9995,N_9542,N_9018);
nand U9996 (N_9996,N_8843,N_9005);
xor U9997 (N_9997,N_9595,N_9169);
nand U9998 (N_9998,N_8891,N_9035);
xor U9999 (N_9999,N_9177,N_9077);
xnor U10000 (N_10000,N_8856,N_8918);
nor U10001 (N_10001,N_9353,N_9348);
nand U10002 (N_10002,N_8855,N_9554);
nor U10003 (N_10003,N_8826,N_9287);
and U10004 (N_10004,N_9519,N_9030);
nand U10005 (N_10005,N_8810,N_8936);
nand U10006 (N_10006,N_8832,N_9219);
or U10007 (N_10007,N_9295,N_9046);
xor U10008 (N_10008,N_9086,N_9529);
xnor U10009 (N_10009,N_8868,N_8836);
or U10010 (N_10010,N_8895,N_8863);
nand U10011 (N_10011,N_9392,N_8893);
xnor U10012 (N_10012,N_9299,N_9088);
nor U10013 (N_10013,N_9276,N_9011);
or U10014 (N_10014,N_9419,N_9398);
nor U10015 (N_10015,N_9540,N_9253);
nand U10016 (N_10016,N_9192,N_8866);
nor U10017 (N_10017,N_9059,N_8937);
nand U10018 (N_10018,N_8833,N_9050);
or U10019 (N_10019,N_9569,N_9196);
xor U10020 (N_10020,N_9179,N_8982);
xor U10021 (N_10021,N_9436,N_9551);
or U10022 (N_10022,N_9146,N_9475);
nand U10023 (N_10023,N_9020,N_8968);
or U10024 (N_10024,N_8991,N_9496);
xnor U10025 (N_10025,N_9421,N_8861);
xor U10026 (N_10026,N_8944,N_9501);
or U10027 (N_10027,N_9263,N_9367);
or U10028 (N_10028,N_9394,N_9595);
nor U10029 (N_10029,N_9236,N_9283);
xnor U10030 (N_10030,N_9237,N_9014);
xnor U10031 (N_10031,N_9212,N_9553);
or U10032 (N_10032,N_9074,N_9372);
xor U10033 (N_10033,N_9399,N_9595);
nor U10034 (N_10034,N_8856,N_9002);
and U10035 (N_10035,N_9590,N_8913);
nand U10036 (N_10036,N_9232,N_9243);
xor U10037 (N_10037,N_8812,N_8816);
nor U10038 (N_10038,N_8953,N_8976);
nand U10039 (N_10039,N_8942,N_9379);
or U10040 (N_10040,N_9292,N_9453);
nor U10041 (N_10041,N_8821,N_9052);
or U10042 (N_10042,N_9075,N_9573);
or U10043 (N_10043,N_8884,N_9382);
xor U10044 (N_10044,N_9188,N_8935);
xor U10045 (N_10045,N_9312,N_9459);
nor U10046 (N_10046,N_9391,N_9219);
and U10047 (N_10047,N_9332,N_9128);
or U10048 (N_10048,N_8807,N_9546);
and U10049 (N_10049,N_8838,N_9241);
nor U10050 (N_10050,N_9375,N_8974);
xor U10051 (N_10051,N_9478,N_9481);
and U10052 (N_10052,N_9035,N_9137);
xnor U10053 (N_10053,N_8983,N_9057);
nand U10054 (N_10054,N_9154,N_9245);
nand U10055 (N_10055,N_8944,N_9378);
xnor U10056 (N_10056,N_9332,N_9483);
nor U10057 (N_10057,N_9143,N_9440);
or U10058 (N_10058,N_8852,N_8994);
and U10059 (N_10059,N_8949,N_9103);
nor U10060 (N_10060,N_9092,N_9207);
nor U10061 (N_10061,N_8909,N_8808);
and U10062 (N_10062,N_8891,N_9256);
nand U10063 (N_10063,N_9578,N_9334);
and U10064 (N_10064,N_9199,N_9186);
and U10065 (N_10065,N_9152,N_8839);
xnor U10066 (N_10066,N_8955,N_9125);
or U10067 (N_10067,N_9058,N_9364);
nor U10068 (N_10068,N_9171,N_9387);
xnor U10069 (N_10069,N_9465,N_9133);
or U10070 (N_10070,N_9083,N_9191);
nor U10071 (N_10071,N_9505,N_9501);
and U10072 (N_10072,N_9492,N_9541);
nand U10073 (N_10073,N_8924,N_8896);
nand U10074 (N_10074,N_9374,N_9097);
xor U10075 (N_10075,N_9557,N_8852);
xnor U10076 (N_10076,N_8906,N_9285);
nor U10077 (N_10077,N_8867,N_8817);
xnor U10078 (N_10078,N_9316,N_8805);
xnor U10079 (N_10079,N_8890,N_8985);
and U10080 (N_10080,N_9296,N_9377);
nor U10081 (N_10081,N_9308,N_9290);
xor U10082 (N_10082,N_8956,N_9080);
xnor U10083 (N_10083,N_9165,N_9256);
or U10084 (N_10084,N_9067,N_9239);
nand U10085 (N_10085,N_9540,N_9493);
nand U10086 (N_10086,N_9227,N_9256);
or U10087 (N_10087,N_9004,N_9528);
nor U10088 (N_10088,N_9064,N_9520);
nor U10089 (N_10089,N_9521,N_9244);
nand U10090 (N_10090,N_9013,N_9280);
nand U10091 (N_10091,N_9079,N_9442);
nand U10092 (N_10092,N_9416,N_9262);
xor U10093 (N_10093,N_8856,N_9214);
and U10094 (N_10094,N_9290,N_9316);
nand U10095 (N_10095,N_9412,N_9474);
nand U10096 (N_10096,N_9308,N_8994);
nor U10097 (N_10097,N_8913,N_9503);
nor U10098 (N_10098,N_8931,N_8897);
nand U10099 (N_10099,N_8921,N_9109);
nand U10100 (N_10100,N_8942,N_9536);
or U10101 (N_10101,N_9371,N_9274);
nor U10102 (N_10102,N_9069,N_9374);
and U10103 (N_10103,N_8945,N_9085);
xnor U10104 (N_10104,N_9376,N_9141);
or U10105 (N_10105,N_9469,N_8827);
nand U10106 (N_10106,N_9090,N_9093);
nand U10107 (N_10107,N_9354,N_9156);
and U10108 (N_10108,N_9126,N_9104);
and U10109 (N_10109,N_9192,N_9142);
nor U10110 (N_10110,N_9337,N_9198);
xnor U10111 (N_10111,N_9440,N_9266);
or U10112 (N_10112,N_9590,N_8982);
nand U10113 (N_10113,N_9310,N_9415);
nand U10114 (N_10114,N_9484,N_9109);
and U10115 (N_10115,N_8868,N_9109);
nor U10116 (N_10116,N_8916,N_9013);
or U10117 (N_10117,N_8844,N_9367);
nand U10118 (N_10118,N_8807,N_9568);
or U10119 (N_10119,N_9510,N_8867);
or U10120 (N_10120,N_9202,N_9307);
or U10121 (N_10121,N_8930,N_9241);
nand U10122 (N_10122,N_9564,N_8963);
xor U10123 (N_10123,N_8930,N_9307);
and U10124 (N_10124,N_9357,N_8887);
and U10125 (N_10125,N_9232,N_9471);
xnor U10126 (N_10126,N_8972,N_8932);
and U10127 (N_10127,N_9241,N_9344);
and U10128 (N_10128,N_8896,N_9433);
and U10129 (N_10129,N_8801,N_8912);
or U10130 (N_10130,N_9549,N_9191);
nor U10131 (N_10131,N_9127,N_9265);
or U10132 (N_10132,N_9385,N_8839);
or U10133 (N_10133,N_9186,N_9334);
nor U10134 (N_10134,N_9508,N_9363);
or U10135 (N_10135,N_9335,N_8995);
and U10136 (N_10136,N_8804,N_8941);
or U10137 (N_10137,N_9427,N_9537);
nand U10138 (N_10138,N_9369,N_8839);
or U10139 (N_10139,N_9045,N_9095);
nand U10140 (N_10140,N_9154,N_9451);
or U10141 (N_10141,N_9015,N_9343);
or U10142 (N_10142,N_9030,N_9003);
nand U10143 (N_10143,N_9044,N_9248);
xnor U10144 (N_10144,N_8806,N_9499);
nand U10145 (N_10145,N_8830,N_9120);
or U10146 (N_10146,N_8902,N_9370);
nand U10147 (N_10147,N_8995,N_8919);
or U10148 (N_10148,N_8931,N_9559);
or U10149 (N_10149,N_8979,N_9228);
xor U10150 (N_10150,N_9395,N_9238);
nand U10151 (N_10151,N_9514,N_9556);
or U10152 (N_10152,N_8859,N_9522);
and U10153 (N_10153,N_9380,N_9278);
nand U10154 (N_10154,N_8953,N_9454);
nand U10155 (N_10155,N_9191,N_8910);
and U10156 (N_10156,N_8944,N_8874);
nor U10157 (N_10157,N_9114,N_8845);
nand U10158 (N_10158,N_9238,N_9498);
nor U10159 (N_10159,N_8974,N_9580);
and U10160 (N_10160,N_8866,N_9425);
and U10161 (N_10161,N_8866,N_9372);
xor U10162 (N_10162,N_9593,N_9233);
xor U10163 (N_10163,N_8929,N_9251);
and U10164 (N_10164,N_9054,N_9334);
and U10165 (N_10165,N_9524,N_8959);
nand U10166 (N_10166,N_8909,N_9593);
and U10167 (N_10167,N_9286,N_9235);
and U10168 (N_10168,N_9424,N_9309);
or U10169 (N_10169,N_9089,N_9033);
nor U10170 (N_10170,N_8888,N_9531);
nor U10171 (N_10171,N_9158,N_8852);
and U10172 (N_10172,N_9111,N_9478);
xor U10173 (N_10173,N_9180,N_9249);
xor U10174 (N_10174,N_9231,N_8885);
nand U10175 (N_10175,N_9266,N_9218);
or U10176 (N_10176,N_9166,N_8804);
nor U10177 (N_10177,N_9015,N_9028);
and U10178 (N_10178,N_9407,N_9306);
nor U10179 (N_10179,N_8802,N_8878);
nand U10180 (N_10180,N_9120,N_9392);
and U10181 (N_10181,N_9278,N_8902);
xnor U10182 (N_10182,N_9408,N_8908);
nand U10183 (N_10183,N_9295,N_9107);
and U10184 (N_10184,N_8931,N_9196);
nand U10185 (N_10185,N_8984,N_8958);
nand U10186 (N_10186,N_9503,N_9080);
and U10187 (N_10187,N_9392,N_9148);
and U10188 (N_10188,N_9242,N_9348);
or U10189 (N_10189,N_9520,N_9561);
and U10190 (N_10190,N_8900,N_8944);
nor U10191 (N_10191,N_9390,N_8953);
xnor U10192 (N_10192,N_9101,N_9471);
xor U10193 (N_10193,N_9275,N_9082);
or U10194 (N_10194,N_8930,N_9591);
xnor U10195 (N_10195,N_9421,N_8940);
xor U10196 (N_10196,N_9306,N_9552);
and U10197 (N_10197,N_9423,N_9385);
or U10198 (N_10198,N_9425,N_8929);
nor U10199 (N_10199,N_9393,N_8979);
xor U10200 (N_10200,N_9205,N_8994);
nand U10201 (N_10201,N_8896,N_9220);
nor U10202 (N_10202,N_9595,N_8890);
nor U10203 (N_10203,N_8909,N_9473);
or U10204 (N_10204,N_9093,N_8881);
or U10205 (N_10205,N_8809,N_9287);
xor U10206 (N_10206,N_9587,N_9453);
nor U10207 (N_10207,N_9221,N_9356);
and U10208 (N_10208,N_9576,N_9580);
nand U10209 (N_10209,N_9245,N_9382);
or U10210 (N_10210,N_8878,N_9361);
nand U10211 (N_10211,N_8993,N_9314);
nor U10212 (N_10212,N_9329,N_9223);
and U10213 (N_10213,N_9176,N_9070);
xor U10214 (N_10214,N_9319,N_8953);
and U10215 (N_10215,N_9228,N_9073);
xnor U10216 (N_10216,N_9133,N_9117);
or U10217 (N_10217,N_9519,N_8981);
nor U10218 (N_10218,N_8868,N_9366);
nor U10219 (N_10219,N_9506,N_8907);
xnor U10220 (N_10220,N_9475,N_9264);
nand U10221 (N_10221,N_8867,N_9388);
nand U10222 (N_10222,N_9083,N_9378);
nor U10223 (N_10223,N_9088,N_9236);
xor U10224 (N_10224,N_9019,N_9527);
and U10225 (N_10225,N_9274,N_8985);
and U10226 (N_10226,N_9244,N_9317);
and U10227 (N_10227,N_9589,N_8982);
and U10228 (N_10228,N_9232,N_9185);
and U10229 (N_10229,N_9293,N_9232);
xor U10230 (N_10230,N_9030,N_8825);
or U10231 (N_10231,N_9447,N_8846);
xor U10232 (N_10232,N_9299,N_9226);
nand U10233 (N_10233,N_8977,N_9299);
nand U10234 (N_10234,N_8907,N_8855);
nor U10235 (N_10235,N_8812,N_9307);
or U10236 (N_10236,N_8982,N_9147);
xor U10237 (N_10237,N_9333,N_9359);
nor U10238 (N_10238,N_9579,N_8960);
nand U10239 (N_10239,N_9032,N_9088);
xor U10240 (N_10240,N_9349,N_9064);
nor U10241 (N_10241,N_8860,N_9286);
nand U10242 (N_10242,N_8886,N_9499);
nor U10243 (N_10243,N_9495,N_8820);
or U10244 (N_10244,N_9487,N_8877);
xnor U10245 (N_10245,N_9327,N_8813);
or U10246 (N_10246,N_9550,N_9576);
nor U10247 (N_10247,N_8809,N_9497);
or U10248 (N_10248,N_9117,N_9034);
or U10249 (N_10249,N_9014,N_9356);
nor U10250 (N_10250,N_9596,N_9027);
and U10251 (N_10251,N_9476,N_9585);
and U10252 (N_10252,N_9392,N_9348);
nand U10253 (N_10253,N_9130,N_9391);
xor U10254 (N_10254,N_8934,N_9158);
and U10255 (N_10255,N_9542,N_9536);
or U10256 (N_10256,N_9514,N_9288);
xor U10257 (N_10257,N_9291,N_9564);
xnor U10258 (N_10258,N_9314,N_9440);
and U10259 (N_10259,N_8937,N_9051);
nand U10260 (N_10260,N_9533,N_8814);
and U10261 (N_10261,N_9181,N_9208);
and U10262 (N_10262,N_9599,N_8821);
or U10263 (N_10263,N_9395,N_9501);
nor U10264 (N_10264,N_9489,N_9054);
nand U10265 (N_10265,N_9427,N_9037);
nand U10266 (N_10266,N_9028,N_9010);
xor U10267 (N_10267,N_9234,N_9226);
xnor U10268 (N_10268,N_9536,N_9114);
xnor U10269 (N_10269,N_9034,N_9050);
and U10270 (N_10270,N_8935,N_9051);
nand U10271 (N_10271,N_9337,N_8929);
xnor U10272 (N_10272,N_8944,N_8975);
nor U10273 (N_10273,N_9316,N_9019);
or U10274 (N_10274,N_9019,N_9108);
and U10275 (N_10275,N_9487,N_9435);
and U10276 (N_10276,N_9464,N_9450);
and U10277 (N_10277,N_9027,N_9533);
xor U10278 (N_10278,N_9465,N_9249);
xnor U10279 (N_10279,N_9147,N_9191);
xor U10280 (N_10280,N_8802,N_9109);
or U10281 (N_10281,N_9381,N_8865);
nand U10282 (N_10282,N_9388,N_9190);
xnor U10283 (N_10283,N_9160,N_9590);
or U10284 (N_10284,N_9183,N_9556);
nor U10285 (N_10285,N_9103,N_9366);
xnor U10286 (N_10286,N_9247,N_8812);
or U10287 (N_10287,N_9059,N_9346);
or U10288 (N_10288,N_8831,N_9465);
xnor U10289 (N_10289,N_8842,N_9087);
nand U10290 (N_10290,N_8954,N_9381);
nor U10291 (N_10291,N_9405,N_9597);
xnor U10292 (N_10292,N_9238,N_9205);
and U10293 (N_10293,N_9268,N_9474);
nor U10294 (N_10294,N_9292,N_9115);
nor U10295 (N_10295,N_8945,N_8994);
and U10296 (N_10296,N_9563,N_9247);
nor U10297 (N_10297,N_9438,N_9266);
and U10298 (N_10298,N_9329,N_9178);
or U10299 (N_10299,N_9156,N_9127);
xnor U10300 (N_10300,N_9375,N_9506);
or U10301 (N_10301,N_8956,N_9510);
xnor U10302 (N_10302,N_9253,N_9405);
or U10303 (N_10303,N_9579,N_8872);
xnor U10304 (N_10304,N_9046,N_9156);
xor U10305 (N_10305,N_9007,N_9369);
nand U10306 (N_10306,N_9431,N_9465);
or U10307 (N_10307,N_9087,N_9129);
nor U10308 (N_10308,N_9519,N_9258);
and U10309 (N_10309,N_9353,N_8884);
nor U10310 (N_10310,N_9395,N_9474);
nor U10311 (N_10311,N_9476,N_9230);
and U10312 (N_10312,N_9557,N_9550);
nand U10313 (N_10313,N_9398,N_8970);
and U10314 (N_10314,N_9456,N_9289);
or U10315 (N_10315,N_9417,N_9411);
xor U10316 (N_10316,N_9385,N_9377);
nand U10317 (N_10317,N_9243,N_8845);
nand U10318 (N_10318,N_8995,N_9304);
or U10319 (N_10319,N_9143,N_8954);
xor U10320 (N_10320,N_9469,N_8866);
nand U10321 (N_10321,N_9023,N_9494);
and U10322 (N_10322,N_8882,N_8811);
and U10323 (N_10323,N_9436,N_8919);
nand U10324 (N_10324,N_9565,N_8925);
xor U10325 (N_10325,N_8970,N_8889);
xor U10326 (N_10326,N_9036,N_9521);
and U10327 (N_10327,N_8913,N_9192);
nor U10328 (N_10328,N_9155,N_9402);
and U10329 (N_10329,N_8943,N_9113);
xor U10330 (N_10330,N_9416,N_8845);
or U10331 (N_10331,N_9234,N_9497);
nor U10332 (N_10332,N_8915,N_9091);
nand U10333 (N_10333,N_9230,N_9209);
nand U10334 (N_10334,N_9480,N_9183);
and U10335 (N_10335,N_9489,N_9473);
and U10336 (N_10336,N_9345,N_9347);
nand U10337 (N_10337,N_9117,N_8900);
xor U10338 (N_10338,N_9229,N_8863);
nand U10339 (N_10339,N_8929,N_8960);
or U10340 (N_10340,N_9467,N_9028);
nor U10341 (N_10341,N_9348,N_9355);
xnor U10342 (N_10342,N_9406,N_9034);
xnor U10343 (N_10343,N_9202,N_9022);
nand U10344 (N_10344,N_9119,N_9244);
xor U10345 (N_10345,N_9035,N_9367);
nor U10346 (N_10346,N_8904,N_9535);
and U10347 (N_10347,N_9547,N_9343);
and U10348 (N_10348,N_9025,N_9314);
nor U10349 (N_10349,N_9301,N_9207);
or U10350 (N_10350,N_9095,N_9502);
xnor U10351 (N_10351,N_9209,N_9211);
nor U10352 (N_10352,N_9304,N_9502);
xnor U10353 (N_10353,N_9165,N_9001);
nand U10354 (N_10354,N_9176,N_9496);
xnor U10355 (N_10355,N_9449,N_9431);
xor U10356 (N_10356,N_8836,N_9209);
nand U10357 (N_10357,N_9298,N_9520);
and U10358 (N_10358,N_9052,N_9117);
or U10359 (N_10359,N_8848,N_9315);
nand U10360 (N_10360,N_8884,N_9415);
or U10361 (N_10361,N_8863,N_9001);
nor U10362 (N_10362,N_9524,N_8940);
or U10363 (N_10363,N_9196,N_9251);
or U10364 (N_10364,N_8917,N_9381);
xnor U10365 (N_10365,N_9455,N_9006);
xor U10366 (N_10366,N_9131,N_9494);
nand U10367 (N_10367,N_9285,N_9470);
xor U10368 (N_10368,N_8835,N_9436);
nor U10369 (N_10369,N_8832,N_9060);
and U10370 (N_10370,N_9413,N_9434);
nand U10371 (N_10371,N_9054,N_9122);
xnor U10372 (N_10372,N_9326,N_8921);
nor U10373 (N_10373,N_9292,N_9567);
nor U10374 (N_10374,N_9370,N_9026);
nor U10375 (N_10375,N_8886,N_8854);
nor U10376 (N_10376,N_9315,N_9083);
and U10377 (N_10377,N_9405,N_9300);
nor U10378 (N_10378,N_9343,N_8954);
xor U10379 (N_10379,N_8814,N_9133);
nand U10380 (N_10380,N_9289,N_9088);
nand U10381 (N_10381,N_8979,N_9466);
and U10382 (N_10382,N_9049,N_8886);
or U10383 (N_10383,N_8862,N_9177);
nand U10384 (N_10384,N_9477,N_9589);
or U10385 (N_10385,N_8863,N_9467);
xnor U10386 (N_10386,N_9252,N_9116);
and U10387 (N_10387,N_9181,N_9001);
xnor U10388 (N_10388,N_8909,N_9556);
xnor U10389 (N_10389,N_9586,N_9176);
nand U10390 (N_10390,N_8954,N_9451);
xnor U10391 (N_10391,N_9377,N_8956);
nand U10392 (N_10392,N_8815,N_9461);
and U10393 (N_10393,N_9421,N_9172);
nand U10394 (N_10394,N_9477,N_9532);
and U10395 (N_10395,N_9564,N_9062);
nand U10396 (N_10396,N_8887,N_9292);
and U10397 (N_10397,N_9135,N_9359);
or U10398 (N_10398,N_9529,N_9169);
xor U10399 (N_10399,N_9215,N_9583);
xor U10400 (N_10400,N_10044,N_10252);
nor U10401 (N_10401,N_9923,N_9955);
or U10402 (N_10402,N_9766,N_10136);
and U10403 (N_10403,N_10265,N_9888);
nand U10404 (N_10404,N_9776,N_9869);
nor U10405 (N_10405,N_9631,N_9607);
xnor U10406 (N_10406,N_9764,N_10125);
nand U10407 (N_10407,N_10114,N_10348);
xor U10408 (N_10408,N_9709,N_10042);
xor U10409 (N_10409,N_10092,N_9903);
or U10410 (N_10410,N_10261,N_9845);
or U10411 (N_10411,N_10315,N_10381);
nor U10412 (N_10412,N_10070,N_10239);
or U10413 (N_10413,N_10144,N_10147);
nor U10414 (N_10414,N_10032,N_9938);
or U10415 (N_10415,N_10049,N_10105);
nand U10416 (N_10416,N_10289,N_10337);
nand U10417 (N_10417,N_10204,N_10072);
nand U10418 (N_10418,N_10215,N_9711);
xor U10419 (N_10419,N_9978,N_10318);
nor U10420 (N_10420,N_10190,N_10104);
xor U10421 (N_10421,N_9696,N_10330);
xor U10422 (N_10422,N_9873,N_10119);
xnor U10423 (N_10423,N_9962,N_9778);
xor U10424 (N_10424,N_9747,N_10058);
or U10425 (N_10425,N_10392,N_9769);
nand U10426 (N_10426,N_9694,N_9918);
nand U10427 (N_10427,N_9810,N_9922);
or U10428 (N_10428,N_10160,N_9628);
nand U10429 (N_10429,N_9894,N_9743);
nand U10430 (N_10430,N_9773,N_10314);
or U10431 (N_10431,N_10222,N_9801);
or U10432 (N_10432,N_10145,N_10101);
nand U10433 (N_10433,N_9952,N_9620);
xnor U10434 (N_10434,N_9805,N_10023);
nand U10435 (N_10435,N_10246,N_9913);
or U10436 (N_10436,N_9970,N_10161);
xor U10437 (N_10437,N_10163,N_9860);
or U10438 (N_10438,N_9725,N_10238);
xor U10439 (N_10439,N_9682,N_9901);
nor U10440 (N_10440,N_9821,N_9670);
nor U10441 (N_10441,N_10243,N_9833);
or U10442 (N_10442,N_9914,N_10322);
xnor U10443 (N_10443,N_10067,N_9878);
and U10444 (N_10444,N_10179,N_9789);
and U10445 (N_10445,N_9794,N_9707);
nand U10446 (N_10446,N_10180,N_9880);
or U10447 (N_10447,N_9720,N_10131);
xnor U10448 (N_10448,N_10078,N_10090);
xnor U10449 (N_10449,N_10361,N_9606);
and U10450 (N_10450,N_9925,N_10003);
or U10451 (N_10451,N_10019,N_9910);
and U10452 (N_10452,N_10077,N_10111);
and U10453 (N_10453,N_10218,N_9884);
nand U10454 (N_10454,N_10065,N_10095);
xnor U10455 (N_10455,N_9994,N_10301);
xor U10456 (N_10456,N_10256,N_9905);
or U10457 (N_10457,N_9784,N_10396);
xor U10458 (N_10458,N_9848,N_10287);
or U10459 (N_10459,N_10312,N_9796);
and U10460 (N_10460,N_9639,N_9678);
nand U10461 (N_10461,N_10217,N_10393);
and U10462 (N_10462,N_9814,N_10296);
xor U10463 (N_10463,N_9812,N_9721);
or U10464 (N_10464,N_9625,N_9636);
xnor U10465 (N_10465,N_9924,N_10043);
nand U10466 (N_10466,N_9985,N_9926);
xnor U10467 (N_10467,N_10225,N_9737);
and U10468 (N_10468,N_10288,N_10235);
or U10469 (N_10469,N_9740,N_10081);
and U10470 (N_10470,N_9763,N_9792);
nor U10471 (N_10471,N_10397,N_10055);
nor U10472 (N_10472,N_9849,N_9852);
and U10473 (N_10473,N_9883,N_10386);
nor U10474 (N_10474,N_9758,N_9948);
nand U10475 (N_10475,N_10024,N_9618);
nand U10476 (N_10476,N_9703,N_10358);
nor U10477 (N_10477,N_10272,N_9647);
and U10478 (N_10478,N_10187,N_9716);
or U10479 (N_10479,N_9917,N_10113);
nand U10480 (N_10480,N_9705,N_9993);
xor U10481 (N_10481,N_10012,N_9783);
nand U10482 (N_10482,N_10008,N_10307);
xor U10483 (N_10483,N_9659,N_10069);
and U10484 (N_10484,N_9717,N_9656);
xnor U10485 (N_10485,N_9959,N_9934);
or U10486 (N_10486,N_10201,N_9602);
and U10487 (N_10487,N_10374,N_10005);
or U10488 (N_10488,N_10368,N_9807);
and U10489 (N_10489,N_10025,N_9729);
xor U10490 (N_10490,N_10011,N_9708);
nand U10491 (N_10491,N_9967,N_9770);
and U10492 (N_10492,N_9835,N_10344);
and U10493 (N_10493,N_9850,N_9988);
xnor U10494 (N_10494,N_10093,N_10399);
nand U10495 (N_10495,N_10297,N_9646);
nor U10496 (N_10496,N_9842,N_9964);
or U10497 (N_10497,N_9838,N_10253);
or U10498 (N_10498,N_10353,N_9634);
nand U10499 (N_10499,N_10142,N_9939);
xor U10500 (N_10500,N_10045,N_9638);
or U10501 (N_10501,N_9754,N_9680);
nand U10502 (N_10502,N_10004,N_10300);
and U10503 (N_10503,N_10341,N_10157);
or U10504 (N_10504,N_9688,N_10202);
nand U10505 (N_10505,N_10317,N_10236);
nor U10506 (N_10506,N_10263,N_9992);
and U10507 (N_10507,N_9665,N_10171);
xor U10508 (N_10508,N_10146,N_10387);
xor U10509 (N_10509,N_9731,N_9775);
and U10510 (N_10510,N_9921,N_9829);
nor U10511 (N_10511,N_9865,N_10098);
or U10512 (N_10512,N_9825,N_9881);
nor U10513 (N_10513,N_10033,N_9661);
nor U10514 (N_10514,N_9834,N_10233);
nor U10515 (N_10515,N_10306,N_10205);
or U10516 (N_10516,N_10010,N_9608);
xor U10517 (N_10517,N_9654,N_9828);
nand U10518 (N_10518,N_10073,N_10380);
xnor U10519 (N_10519,N_9898,N_9809);
nand U10520 (N_10520,N_10237,N_9781);
nand U10521 (N_10521,N_10165,N_10240);
xor U10522 (N_10522,N_9645,N_10195);
xor U10523 (N_10523,N_9946,N_10149);
and U10524 (N_10524,N_9870,N_10308);
nand U10525 (N_10525,N_9757,N_9861);
nor U10526 (N_10526,N_9893,N_9624);
nor U10527 (N_10527,N_9772,N_10298);
or U10528 (N_10528,N_9642,N_10327);
xnor U10529 (N_10529,N_10051,N_9960);
xor U10530 (N_10530,N_10115,N_10310);
nand U10531 (N_10531,N_10151,N_9702);
xnor U10532 (N_10532,N_10385,N_9663);
and U10533 (N_10533,N_9995,N_9627);
nand U10534 (N_10534,N_9673,N_9685);
xor U10535 (N_10535,N_9891,N_10197);
or U10536 (N_10536,N_10020,N_9640);
xor U10537 (N_10537,N_10134,N_10200);
nor U10538 (N_10538,N_10340,N_10026);
xor U10539 (N_10539,N_10159,N_9904);
and U10540 (N_10540,N_10013,N_9683);
or U10541 (N_10541,N_10102,N_10259);
or U10542 (N_10542,N_10103,N_9667);
and U10543 (N_10543,N_10107,N_9936);
xnor U10544 (N_10544,N_10124,N_10099);
or U10545 (N_10545,N_9706,N_10123);
and U10546 (N_10546,N_9859,N_10174);
and U10547 (N_10547,N_10291,N_9786);
xnor U10548 (N_10548,N_10189,N_9611);
xor U10549 (N_10549,N_9609,N_10242);
nand U10550 (N_10550,N_9664,N_9875);
or U10551 (N_10551,N_10338,N_10196);
or U10552 (N_10552,N_10129,N_9980);
and U10553 (N_10553,N_10177,N_10021);
nor U10554 (N_10554,N_10191,N_9735);
and U10555 (N_10555,N_10083,N_10141);
and U10556 (N_10556,N_10370,N_9780);
and U10557 (N_10557,N_10168,N_10009);
nor U10558 (N_10558,N_9687,N_10040);
xnor U10559 (N_10559,N_9882,N_9745);
nor U10560 (N_10560,N_9858,N_10267);
nor U10561 (N_10561,N_10203,N_9698);
and U10562 (N_10562,N_10178,N_10220);
nand U10563 (N_10563,N_10309,N_10332);
nand U10564 (N_10564,N_9866,N_9846);
xnor U10565 (N_10565,N_10313,N_10372);
nor U10566 (N_10566,N_9868,N_10038);
or U10567 (N_10567,N_10278,N_10052);
or U10568 (N_10568,N_9931,N_9957);
or U10569 (N_10569,N_9862,N_9819);
or U10570 (N_10570,N_10356,N_10122);
and U10571 (N_10571,N_9759,N_9623);
and U10572 (N_10572,N_10106,N_10229);
nand U10573 (N_10573,N_10324,N_9847);
nor U10574 (N_10574,N_10050,N_9697);
nand U10575 (N_10575,N_10231,N_9824);
nand U10576 (N_10576,N_9704,N_9765);
xnor U10577 (N_10577,N_10183,N_10373);
xnor U10578 (N_10578,N_10228,N_9864);
and U10579 (N_10579,N_10132,N_10339);
and U10580 (N_10580,N_9614,N_10035);
nand U10581 (N_10581,N_9669,N_10388);
xor U10582 (N_10582,N_10375,N_10234);
or U10583 (N_10583,N_10299,N_10279);
nor U10584 (N_10584,N_10007,N_10295);
nor U10585 (N_10585,N_9774,N_9958);
xor U10586 (N_10586,N_9989,N_10214);
xor U10587 (N_10587,N_9951,N_9818);
or U10588 (N_10588,N_10135,N_10172);
xnor U10589 (N_10589,N_10153,N_9666);
or U10590 (N_10590,N_10328,N_10108);
and U10591 (N_10591,N_10329,N_10367);
and U10592 (N_10592,N_9674,N_10017);
nor U10593 (N_10593,N_9612,N_10275);
and U10594 (N_10594,N_9719,N_9815);
or U10595 (N_10595,N_10212,N_9695);
or U10596 (N_10596,N_10362,N_9996);
xnor U10597 (N_10597,N_9710,N_10192);
nand U10598 (N_10598,N_9643,N_10304);
or U10599 (N_10599,N_9790,N_10232);
xnor U10600 (N_10600,N_10398,N_10254);
or U10601 (N_10601,N_10194,N_9738);
and U10602 (N_10602,N_10096,N_9817);
nor U10603 (N_10603,N_10148,N_10034);
xor U10604 (N_10604,N_9975,N_10321);
and U10605 (N_10605,N_9987,N_9728);
or U10606 (N_10606,N_10053,N_9853);
or U10607 (N_10607,N_9843,N_10193);
and U10608 (N_10608,N_9969,N_10037);
nor U10609 (N_10609,N_10127,N_9981);
and U10610 (N_10610,N_9874,N_9854);
nor U10611 (N_10611,N_10060,N_10366);
xor U10612 (N_10612,N_10303,N_10182);
nand U10613 (N_10613,N_9950,N_9826);
nand U10614 (N_10614,N_10284,N_10320);
and U10615 (N_10615,N_10221,N_9871);
nor U10616 (N_10616,N_9732,N_9616);
nand U10617 (N_10617,N_10150,N_10331);
and U10618 (N_10618,N_10158,N_9672);
or U10619 (N_10619,N_10076,N_9902);
nand U10620 (N_10620,N_10185,N_9648);
nor U10621 (N_10621,N_9644,N_10213);
and U10622 (N_10622,N_9676,N_9653);
or U10623 (N_10623,N_9632,N_10082);
or U10624 (N_10624,N_10226,N_10241);
xnor U10625 (N_10625,N_9726,N_10027);
and U10626 (N_10626,N_10276,N_9605);
and U10627 (N_10627,N_9750,N_9816);
xor U10628 (N_10628,N_9982,N_9649);
and U10629 (N_10629,N_10269,N_9916);
nand U10630 (N_10630,N_10360,N_9851);
nor U10631 (N_10631,N_9813,N_9974);
or U10632 (N_10632,N_9855,N_9953);
nor U10633 (N_10633,N_10006,N_10036);
and U10634 (N_10634,N_9840,N_9797);
nor U10635 (N_10635,N_10068,N_10186);
nand U10636 (N_10636,N_10198,N_9937);
nor U10637 (N_10637,N_10245,N_10209);
and U10638 (N_10638,N_10139,N_9675);
and U10639 (N_10639,N_10002,N_10029);
nand U10640 (N_10640,N_10302,N_10384);
and U10641 (N_10641,N_9771,N_9761);
and U10642 (N_10642,N_9637,N_9929);
and U10643 (N_10643,N_9785,N_9892);
and U10644 (N_10644,N_9979,N_9681);
nand U10645 (N_10645,N_9947,N_10206);
xnor U10646 (N_10646,N_10066,N_9691);
nand U10647 (N_10647,N_9787,N_9793);
nand U10648 (N_10648,N_10211,N_9788);
or U10649 (N_10649,N_10224,N_10248);
nand U10650 (N_10650,N_10271,N_9997);
and U10651 (N_10651,N_10117,N_10173);
and U10652 (N_10652,N_9713,N_10336);
nand U10653 (N_10653,N_10383,N_9718);
xnor U10654 (N_10654,N_9723,N_10347);
nand U10655 (N_10655,N_9885,N_10112);
xnor U10656 (N_10656,N_9863,N_9906);
nand U10657 (N_10657,N_10376,N_9690);
nand U10658 (N_10658,N_9886,N_9782);
or U10659 (N_10659,N_10014,N_10094);
and U10660 (N_10660,N_9744,N_9621);
nand U10661 (N_10661,N_10154,N_9739);
nor U10662 (N_10662,N_9971,N_10118);
xor U10663 (N_10663,N_10349,N_9741);
or U10664 (N_10664,N_9908,N_10063);
xnor U10665 (N_10665,N_9662,N_10273);
xor U10666 (N_10666,N_10333,N_9762);
and U10667 (N_10667,N_9700,N_9617);
nor U10668 (N_10668,N_9613,N_10369);
nand U10669 (N_10669,N_9724,N_10210);
nor U10670 (N_10670,N_9965,N_9999);
xor U10671 (N_10671,N_9601,N_10342);
or U10672 (N_10672,N_10293,N_9689);
xor U10673 (N_10673,N_10137,N_10074);
or U10674 (N_10674,N_10100,N_9748);
and U10675 (N_10675,N_10377,N_9779);
nor U10676 (N_10676,N_10266,N_10316);
nand U10677 (N_10677,N_9635,N_10264);
nor U10678 (N_10678,N_9830,N_10355);
and U10679 (N_10679,N_9808,N_9752);
nand U10680 (N_10680,N_9756,N_9972);
xnor U10681 (N_10681,N_10223,N_10250);
and U10682 (N_10682,N_10109,N_10056);
nand U10683 (N_10683,N_10088,N_9800);
or U10684 (N_10684,N_10001,N_10335);
xor U10685 (N_10685,N_9651,N_9777);
or U10686 (N_10686,N_10345,N_10059);
nor U10687 (N_10687,N_10087,N_9630);
nand U10688 (N_10688,N_10364,N_10323);
and U10689 (N_10689,N_10378,N_10175);
or U10690 (N_10690,N_10062,N_9889);
nor U10691 (N_10691,N_9686,N_10152);
or U10692 (N_10692,N_9734,N_10143);
nor U10693 (N_10693,N_9767,N_9831);
xor U10694 (N_10694,N_9932,N_10294);
xnor U10695 (N_10695,N_10244,N_9629);
xor U10696 (N_10696,N_10389,N_9961);
nor U10697 (N_10697,N_9714,N_9841);
nand U10698 (N_10698,N_10130,N_10311);
xnor U10699 (N_10699,N_9899,N_9890);
nand U10700 (N_10700,N_9896,N_9604);
xnor U10701 (N_10701,N_10110,N_9795);
nor U10702 (N_10702,N_9986,N_9657);
nand U10703 (N_10703,N_10216,N_9920);
or U10704 (N_10704,N_10116,N_9600);
and U10705 (N_10705,N_9911,N_10097);
and U10706 (N_10706,N_10166,N_10274);
xor U10707 (N_10707,N_10054,N_9977);
and U10708 (N_10708,N_9832,N_9768);
or U10709 (N_10709,N_10079,N_9742);
nor U10710 (N_10710,N_10086,N_10155);
xnor U10711 (N_10711,N_9935,N_9879);
and U10712 (N_10712,N_9983,N_9919);
nor U10713 (N_10713,N_10022,N_10075);
or U10714 (N_10714,N_9991,N_10039);
xnor U10715 (N_10715,N_9984,N_10162);
or U10716 (N_10716,N_10080,N_10128);
xor U10717 (N_10717,N_9603,N_9949);
xnor U10718 (N_10718,N_10126,N_10283);
and U10719 (N_10719,N_10249,N_10354);
nor U10720 (N_10720,N_10188,N_10282);
and U10721 (N_10721,N_10395,N_10352);
xor U10722 (N_10722,N_10208,N_9655);
or U10723 (N_10723,N_10091,N_10138);
nand U10724 (N_10724,N_10390,N_9615);
nor U10725 (N_10725,N_9803,N_10285);
or U10726 (N_10726,N_10028,N_10167);
and U10727 (N_10727,N_10319,N_10133);
or U10728 (N_10728,N_9806,N_10262);
xor U10729 (N_10729,N_10057,N_9976);
or U10730 (N_10730,N_10290,N_10030);
nor U10731 (N_10731,N_9956,N_9867);
and U10732 (N_10732,N_9802,N_10334);
nand U10733 (N_10733,N_9684,N_9652);
or U10734 (N_10734,N_10207,N_9973);
nor U10735 (N_10735,N_9900,N_10199);
nor U10736 (N_10736,N_10247,N_9895);
and U10737 (N_10737,N_10346,N_9963);
nand U10738 (N_10738,N_9679,N_9753);
and U10739 (N_10739,N_10120,N_9930);
nand U10740 (N_10740,N_10258,N_9968);
and U10741 (N_10741,N_9954,N_9966);
and U10742 (N_10742,N_9940,N_10140);
xnor U10743 (N_10743,N_10184,N_9733);
or U10744 (N_10744,N_10255,N_9872);
nand U10745 (N_10745,N_9804,N_9799);
and U10746 (N_10746,N_9641,N_9811);
xnor U10747 (N_10747,N_10268,N_9791);
or U10748 (N_10748,N_10363,N_9822);
or U10749 (N_10749,N_10046,N_10292);
and U10750 (N_10750,N_10041,N_10379);
or U10751 (N_10751,N_9856,N_10350);
nor U10752 (N_10752,N_10156,N_10089);
and U10753 (N_10753,N_10280,N_9927);
nand U10754 (N_10754,N_9755,N_10371);
xnor U10755 (N_10755,N_9730,N_9909);
nor U10756 (N_10756,N_10326,N_9827);
and U10757 (N_10757,N_10061,N_9701);
nand U10758 (N_10758,N_10219,N_10176);
nor U10759 (N_10759,N_10343,N_10391);
and U10760 (N_10760,N_9692,N_10359);
xor U10761 (N_10761,N_9844,N_10277);
nand U10762 (N_10762,N_9668,N_10084);
nand U10763 (N_10763,N_9823,N_9736);
and U10764 (N_10764,N_9699,N_10230);
nor U10765 (N_10765,N_9650,N_9712);
nand U10766 (N_10766,N_9837,N_9715);
nor U10767 (N_10767,N_10018,N_10286);
nand U10768 (N_10768,N_9998,N_10181);
xor U10769 (N_10769,N_9933,N_10170);
nand U10770 (N_10770,N_10382,N_9839);
and U10771 (N_10771,N_9746,N_9610);
xnor U10772 (N_10772,N_9677,N_9942);
nor U10773 (N_10773,N_9944,N_9897);
or U10774 (N_10774,N_10048,N_9658);
xnor U10775 (N_10775,N_9749,N_10325);
or U10776 (N_10776,N_9633,N_9820);
nor U10777 (N_10777,N_9877,N_10394);
nor U10778 (N_10778,N_9876,N_10365);
and U10779 (N_10779,N_10164,N_9941);
or U10780 (N_10780,N_9943,N_9619);
and U10781 (N_10781,N_10121,N_9722);
nand U10782 (N_10782,N_10251,N_9751);
xnor U10783 (N_10783,N_9857,N_9990);
or U10784 (N_10784,N_10031,N_10064);
nor U10785 (N_10785,N_10260,N_10000);
or U10786 (N_10786,N_10357,N_9626);
and U10787 (N_10787,N_9945,N_10169);
nand U10788 (N_10788,N_10351,N_9798);
and U10789 (N_10789,N_9622,N_10016);
and U10790 (N_10790,N_9836,N_10047);
nand U10791 (N_10791,N_9760,N_9693);
xnor U10792 (N_10792,N_9915,N_9907);
or U10793 (N_10793,N_10071,N_9928);
nand U10794 (N_10794,N_10305,N_10227);
nand U10795 (N_10795,N_9912,N_10281);
nor U10796 (N_10796,N_9727,N_9671);
and U10797 (N_10797,N_9660,N_10015);
xor U10798 (N_10798,N_9887,N_10257);
nand U10799 (N_10799,N_10270,N_10085);
nand U10800 (N_10800,N_10025,N_10303);
and U10801 (N_10801,N_9760,N_9739);
nand U10802 (N_10802,N_9936,N_9990);
nor U10803 (N_10803,N_10331,N_9944);
and U10804 (N_10804,N_9977,N_10114);
xor U10805 (N_10805,N_9737,N_10105);
and U10806 (N_10806,N_10114,N_9695);
xor U10807 (N_10807,N_9641,N_10113);
nand U10808 (N_10808,N_10230,N_10003);
nor U10809 (N_10809,N_10016,N_9935);
nor U10810 (N_10810,N_9907,N_10240);
or U10811 (N_10811,N_9833,N_10324);
xor U10812 (N_10812,N_10094,N_9745);
nand U10813 (N_10813,N_10234,N_9946);
nor U10814 (N_10814,N_9719,N_10296);
or U10815 (N_10815,N_10358,N_9931);
nor U10816 (N_10816,N_9773,N_10085);
xnor U10817 (N_10817,N_10368,N_10096);
xnor U10818 (N_10818,N_10002,N_10325);
xor U10819 (N_10819,N_10356,N_10164);
xnor U10820 (N_10820,N_9830,N_9790);
xnor U10821 (N_10821,N_10181,N_10052);
and U10822 (N_10822,N_9980,N_9792);
nand U10823 (N_10823,N_9617,N_9937);
nand U10824 (N_10824,N_10058,N_9869);
nor U10825 (N_10825,N_10397,N_9876);
or U10826 (N_10826,N_10089,N_9647);
xnor U10827 (N_10827,N_9984,N_9778);
and U10828 (N_10828,N_10301,N_10294);
nand U10829 (N_10829,N_10343,N_9673);
nor U10830 (N_10830,N_10392,N_9665);
xnor U10831 (N_10831,N_10205,N_9995);
nor U10832 (N_10832,N_9795,N_9611);
or U10833 (N_10833,N_9712,N_10281);
or U10834 (N_10834,N_10168,N_9994);
or U10835 (N_10835,N_10318,N_9768);
nand U10836 (N_10836,N_10035,N_9686);
nand U10837 (N_10837,N_9972,N_9797);
or U10838 (N_10838,N_10139,N_9677);
nor U10839 (N_10839,N_9840,N_10339);
and U10840 (N_10840,N_10094,N_9729);
nor U10841 (N_10841,N_10147,N_9949);
or U10842 (N_10842,N_10107,N_9806);
nor U10843 (N_10843,N_10058,N_9626);
nor U10844 (N_10844,N_10378,N_10036);
nand U10845 (N_10845,N_9730,N_9808);
nor U10846 (N_10846,N_10289,N_10162);
and U10847 (N_10847,N_10198,N_10159);
nand U10848 (N_10848,N_9762,N_9721);
nor U10849 (N_10849,N_9824,N_10221);
and U10850 (N_10850,N_9994,N_9933);
or U10851 (N_10851,N_9774,N_10357);
nor U10852 (N_10852,N_9846,N_9880);
nor U10853 (N_10853,N_9765,N_9713);
or U10854 (N_10854,N_9758,N_9618);
nand U10855 (N_10855,N_9601,N_10357);
or U10856 (N_10856,N_10217,N_9860);
or U10857 (N_10857,N_9921,N_10250);
and U10858 (N_10858,N_9807,N_10079);
or U10859 (N_10859,N_9697,N_10339);
xor U10860 (N_10860,N_9621,N_9933);
xnor U10861 (N_10861,N_10106,N_10193);
xnor U10862 (N_10862,N_10169,N_10373);
and U10863 (N_10863,N_9874,N_10002);
nand U10864 (N_10864,N_10163,N_10204);
and U10865 (N_10865,N_9724,N_9769);
or U10866 (N_10866,N_9631,N_9816);
nand U10867 (N_10867,N_10129,N_9618);
or U10868 (N_10868,N_10184,N_10158);
and U10869 (N_10869,N_9945,N_9849);
and U10870 (N_10870,N_9771,N_9916);
or U10871 (N_10871,N_10250,N_10221);
xnor U10872 (N_10872,N_9926,N_10088);
nor U10873 (N_10873,N_10339,N_10273);
nor U10874 (N_10874,N_10333,N_10340);
or U10875 (N_10875,N_10229,N_10005);
nand U10876 (N_10876,N_10046,N_10339);
xor U10877 (N_10877,N_9860,N_10306);
nand U10878 (N_10878,N_10033,N_9876);
nand U10879 (N_10879,N_10025,N_10202);
nand U10880 (N_10880,N_10143,N_10067);
nor U10881 (N_10881,N_9929,N_9753);
and U10882 (N_10882,N_10023,N_9822);
nand U10883 (N_10883,N_9922,N_10002);
or U10884 (N_10884,N_9760,N_10247);
nor U10885 (N_10885,N_10225,N_9864);
or U10886 (N_10886,N_10061,N_10371);
xor U10887 (N_10887,N_10277,N_10130);
or U10888 (N_10888,N_9690,N_9930);
or U10889 (N_10889,N_10376,N_10237);
or U10890 (N_10890,N_10140,N_9930);
nor U10891 (N_10891,N_9962,N_9843);
nor U10892 (N_10892,N_9806,N_10013);
nor U10893 (N_10893,N_9729,N_9609);
nand U10894 (N_10894,N_10233,N_9860);
nor U10895 (N_10895,N_9937,N_9728);
nand U10896 (N_10896,N_10249,N_10206);
nand U10897 (N_10897,N_10182,N_9888);
or U10898 (N_10898,N_10118,N_9629);
xor U10899 (N_10899,N_9622,N_9882);
nor U10900 (N_10900,N_10054,N_9957);
or U10901 (N_10901,N_10202,N_10392);
or U10902 (N_10902,N_9737,N_9726);
and U10903 (N_10903,N_10045,N_10293);
and U10904 (N_10904,N_9856,N_10105);
xor U10905 (N_10905,N_10214,N_10199);
or U10906 (N_10906,N_9626,N_10196);
and U10907 (N_10907,N_10043,N_10102);
nand U10908 (N_10908,N_9679,N_9831);
or U10909 (N_10909,N_9940,N_10044);
xor U10910 (N_10910,N_10275,N_10193);
nand U10911 (N_10911,N_10301,N_9961);
or U10912 (N_10912,N_10080,N_10024);
nand U10913 (N_10913,N_10399,N_10007);
nor U10914 (N_10914,N_9999,N_9938);
xnor U10915 (N_10915,N_9636,N_9960);
xor U10916 (N_10916,N_10063,N_10073);
or U10917 (N_10917,N_10071,N_10181);
or U10918 (N_10918,N_10369,N_9779);
nor U10919 (N_10919,N_9737,N_10127);
nor U10920 (N_10920,N_10008,N_9872);
nor U10921 (N_10921,N_9984,N_9642);
and U10922 (N_10922,N_9744,N_9793);
or U10923 (N_10923,N_10047,N_10312);
xor U10924 (N_10924,N_10143,N_10204);
or U10925 (N_10925,N_10131,N_9978);
or U10926 (N_10926,N_9634,N_9872);
or U10927 (N_10927,N_10337,N_10152);
and U10928 (N_10928,N_10157,N_10079);
nor U10929 (N_10929,N_10227,N_10066);
xnor U10930 (N_10930,N_10260,N_9981);
nor U10931 (N_10931,N_9977,N_9906);
nor U10932 (N_10932,N_9876,N_9962);
and U10933 (N_10933,N_9621,N_9756);
nand U10934 (N_10934,N_10265,N_10087);
nand U10935 (N_10935,N_10344,N_10037);
nor U10936 (N_10936,N_9917,N_9601);
xor U10937 (N_10937,N_9708,N_9906);
nand U10938 (N_10938,N_10310,N_9963);
and U10939 (N_10939,N_9998,N_10065);
or U10940 (N_10940,N_10288,N_10050);
and U10941 (N_10941,N_10240,N_10376);
or U10942 (N_10942,N_9996,N_10314);
or U10943 (N_10943,N_9718,N_10379);
or U10944 (N_10944,N_9791,N_10245);
or U10945 (N_10945,N_10047,N_10179);
xnor U10946 (N_10946,N_10248,N_9640);
and U10947 (N_10947,N_9743,N_9745);
and U10948 (N_10948,N_10232,N_10067);
and U10949 (N_10949,N_10284,N_10100);
and U10950 (N_10950,N_10283,N_9931);
nor U10951 (N_10951,N_10149,N_9823);
xnor U10952 (N_10952,N_10023,N_9895);
or U10953 (N_10953,N_10358,N_9669);
and U10954 (N_10954,N_10070,N_9698);
nor U10955 (N_10955,N_10380,N_9774);
nor U10956 (N_10956,N_9836,N_9785);
or U10957 (N_10957,N_9625,N_10043);
nor U10958 (N_10958,N_10317,N_9712);
nor U10959 (N_10959,N_9815,N_10355);
and U10960 (N_10960,N_9739,N_10223);
or U10961 (N_10961,N_10241,N_10265);
nand U10962 (N_10962,N_10015,N_9611);
or U10963 (N_10963,N_10168,N_10013);
xnor U10964 (N_10964,N_9746,N_9787);
nand U10965 (N_10965,N_9724,N_9928);
or U10966 (N_10966,N_9725,N_9888);
and U10967 (N_10967,N_10326,N_9865);
nand U10968 (N_10968,N_10187,N_10070);
xor U10969 (N_10969,N_9864,N_9764);
xnor U10970 (N_10970,N_9714,N_9709);
nand U10971 (N_10971,N_10236,N_10148);
nor U10972 (N_10972,N_9973,N_9682);
nand U10973 (N_10973,N_9756,N_10090);
xnor U10974 (N_10974,N_9671,N_10008);
or U10975 (N_10975,N_9813,N_10054);
nor U10976 (N_10976,N_10202,N_10163);
nand U10977 (N_10977,N_10156,N_9984);
or U10978 (N_10978,N_10012,N_10298);
nor U10979 (N_10979,N_9882,N_9869);
nand U10980 (N_10980,N_10020,N_10119);
xnor U10981 (N_10981,N_9961,N_9632);
nor U10982 (N_10982,N_9774,N_10074);
nor U10983 (N_10983,N_10117,N_10207);
and U10984 (N_10984,N_9949,N_9729);
nand U10985 (N_10985,N_10218,N_10173);
and U10986 (N_10986,N_10009,N_9875);
and U10987 (N_10987,N_10100,N_9757);
nor U10988 (N_10988,N_9998,N_9667);
nand U10989 (N_10989,N_10363,N_9606);
nand U10990 (N_10990,N_10356,N_10298);
and U10991 (N_10991,N_10272,N_9967);
or U10992 (N_10992,N_9830,N_9941);
nor U10993 (N_10993,N_10001,N_10187);
and U10994 (N_10994,N_10117,N_9628);
xnor U10995 (N_10995,N_10342,N_9758);
and U10996 (N_10996,N_10167,N_9754);
nor U10997 (N_10997,N_10104,N_9988);
nor U10998 (N_10998,N_10176,N_10328);
xnor U10999 (N_10999,N_9834,N_9988);
and U11000 (N_11000,N_10047,N_10363);
nor U11001 (N_11001,N_10139,N_10181);
nand U11002 (N_11002,N_10289,N_9659);
nand U11003 (N_11003,N_9698,N_10212);
or U11004 (N_11004,N_9654,N_10012);
and U11005 (N_11005,N_9610,N_10363);
nor U11006 (N_11006,N_10312,N_9845);
or U11007 (N_11007,N_9652,N_9727);
nor U11008 (N_11008,N_9993,N_10061);
xnor U11009 (N_11009,N_10395,N_10201);
or U11010 (N_11010,N_10132,N_10133);
nor U11011 (N_11011,N_10234,N_9973);
xor U11012 (N_11012,N_10095,N_9907);
or U11013 (N_11013,N_9698,N_10320);
and U11014 (N_11014,N_9907,N_9621);
xor U11015 (N_11015,N_10089,N_9948);
and U11016 (N_11016,N_9776,N_9937);
or U11017 (N_11017,N_9694,N_10349);
or U11018 (N_11018,N_9926,N_10138);
or U11019 (N_11019,N_10144,N_9837);
and U11020 (N_11020,N_9912,N_9642);
xor U11021 (N_11021,N_10267,N_10065);
nand U11022 (N_11022,N_10357,N_10130);
nor U11023 (N_11023,N_9605,N_10356);
nand U11024 (N_11024,N_10186,N_10122);
xnor U11025 (N_11025,N_10012,N_9764);
nor U11026 (N_11026,N_9611,N_10179);
nand U11027 (N_11027,N_9922,N_10395);
nand U11028 (N_11028,N_9678,N_9906);
and U11029 (N_11029,N_10156,N_9792);
nor U11030 (N_11030,N_9752,N_9634);
nor U11031 (N_11031,N_9867,N_9951);
nor U11032 (N_11032,N_9930,N_9770);
or U11033 (N_11033,N_10016,N_10369);
xnor U11034 (N_11034,N_10241,N_10198);
or U11035 (N_11035,N_9631,N_10309);
or U11036 (N_11036,N_9967,N_9980);
and U11037 (N_11037,N_9808,N_10068);
or U11038 (N_11038,N_9701,N_10217);
nor U11039 (N_11039,N_9649,N_9644);
nand U11040 (N_11040,N_10132,N_9798);
and U11041 (N_11041,N_9986,N_9983);
nand U11042 (N_11042,N_10203,N_10299);
or U11043 (N_11043,N_10260,N_10314);
nor U11044 (N_11044,N_9617,N_10001);
nand U11045 (N_11045,N_9863,N_10112);
nand U11046 (N_11046,N_10008,N_9690);
or U11047 (N_11047,N_10308,N_10258);
xor U11048 (N_11048,N_10059,N_9811);
nand U11049 (N_11049,N_10324,N_10093);
nand U11050 (N_11050,N_9776,N_10065);
xnor U11051 (N_11051,N_10089,N_9881);
nand U11052 (N_11052,N_9978,N_9665);
xor U11053 (N_11053,N_9768,N_9632);
nor U11054 (N_11054,N_9895,N_10186);
nand U11055 (N_11055,N_10357,N_9671);
nand U11056 (N_11056,N_9993,N_9873);
nor U11057 (N_11057,N_9802,N_9864);
nand U11058 (N_11058,N_10124,N_9989);
xnor U11059 (N_11059,N_10308,N_10292);
or U11060 (N_11060,N_10214,N_9937);
and U11061 (N_11061,N_9656,N_10289);
xnor U11062 (N_11062,N_10395,N_9639);
and U11063 (N_11063,N_9857,N_10005);
and U11064 (N_11064,N_10001,N_10231);
nor U11065 (N_11065,N_9713,N_9690);
xor U11066 (N_11066,N_10333,N_10354);
xor U11067 (N_11067,N_10106,N_9723);
xnor U11068 (N_11068,N_10262,N_9867);
nor U11069 (N_11069,N_10149,N_9703);
nand U11070 (N_11070,N_10026,N_10180);
nand U11071 (N_11071,N_10291,N_10355);
xnor U11072 (N_11072,N_9764,N_9834);
xor U11073 (N_11073,N_9808,N_10149);
or U11074 (N_11074,N_9759,N_10047);
nand U11075 (N_11075,N_9802,N_9875);
or U11076 (N_11076,N_10082,N_9673);
and U11077 (N_11077,N_9608,N_10190);
xnor U11078 (N_11078,N_9847,N_9809);
xnor U11079 (N_11079,N_9902,N_10058);
or U11080 (N_11080,N_9642,N_10344);
nand U11081 (N_11081,N_9749,N_10035);
nand U11082 (N_11082,N_10292,N_10372);
nand U11083 (N_11083,N_10100,N_10240);
nor U11084 (N_11084,N_10195,N_10125);
and U11085 (N_11085,N_9985,N_10124);
and U11086 (N_11086,N_9867,N_9815);
nand U11087 (N_11087,N_10027,N_9696);
nand U11088 (N_11088,N_10264,N_10169);
nor U11089 (N_11089,N_9791,N_9792);
or U11090 (N_11090,N_9976,N_9995);
or U11091 (N_11091,N_10052,N_9977);
and U11092 (N_11092,N_10193,N_9696);
and U11093 (N_11093,N_9683,N_9750);
nor U11094 (N_11094,N_9605,N_10046);
nand U11095 (N_11095,N_10178,N_9913);
or U11096 (N_11096,N_9996,N_9620);
nor U11097 (N_11097,N_9639,N_10109);
nand U11098 (N_11098,N_9964,N_10001);
nand U11099 (N_11099,N_10176,N_9865);
and U11100 (N_11100,N_9672,N_10022);
nor U11101 (N_11101,N_9927,N_9774);
and U11102 (N_11102,N_9979,N_10035);
xor U11103 (N_11103,N_9971,N_9670);
nand U11104 (N_11104,N_10265,N_10297);
or U11105 (N_11105,N_10006,N_10079);
nand U11106 (N_11106,N_9652,N_10284);
and U11107 (N_11107,N_10244,N_10310);
or U11108 (N_11108,N_10128,N_9994);
xnor U11109 (N_11109,N_9649,N_9765);
nor U11110 (N_11110,N_9954,N_9922);
and U11111 (N_11111,N_10198,N_9836);
or U11112 (N_11112,N_9886,N_10216);
nor U11113 (N_11113,N_10147,N_10156);
nor U11114 (N_11114,N_10131,N_9772);
nand U11115 (N_11115,N_9992,N_9830);
xnor U11116 (N_11116,N_10158,N_9820);
xor U11117 (N_11117,N_10292,N_10064);
or U11118 (N_11118,N_9804,N_10365);
and U11119 (N_11119,N_10211,N_10188);
nand U11120 (N_11120,N_10269,N_9967);
or U11121 (N_11121,N_9891,N_10101);
xor U11122 (N_11122,N_9679,N_10152);
xor U11123 (N_11123,N_10014,N_10225);
or U11124 (N_11124,N_9707,N_9752);
nor U11125 (N_11125,N_10316,N_10093);
nor U11126 (N_11126,N_10393,N_9670);
or U11127 (N_11127,N_10020,N_10283);
nand U11128 (N_11128,N_10339,N_9633);
or U11129 (N_11129,N_10073,N_10228);
and U11130 (N_11130,N_9649,N_10024);
xnor U11131 (N_11131,N_10154,N_9918);
or U11132 (N_11132,N_10226,N_10095);
nand U11133 (N_11133,N_10186,N_9629);
nand U11134 (N_11134,N_10123,N_9960);
or U11135 (N_11135,N_9847,N_10183);
nand U11136 (N_11136,N_9815,N_9792);
nand U11137 (N_11137,N_10084,N_9866);
nand U11138 (N_11138,N_9678,N_10299);
nand U11139 (N_11139,N_9601,N_10146);
nor U11140 (N_11140,N_10043,N_10056);
or U11141 (N_11141,N_10235,N_10119);
nor U11142 (N_11142,N_9770,N_10368);
or U11143 (N_11143,N_10308,N_10219);
nor U11144 (N_11144,N_9675,N_10356);
nand U11145 (N_11145,N_9762,N_10153);
nand U11146 (N_11146,N_9603,N_10200);
nand U11147 (N_11147,N_10293,N_9936);
nor U11148 (N_11148,N_10059,N_9878);
and U11149 (N_11149,N_9903,N_9642);
xor U11150 (N_11150,N_9734,N_9869);
xnor U11151 (N_11151,N_9752,N_9870);
or U11152 (N_11152,N_9620,N_10138);
and U11153 (N_11153,N_9851,N_9783);
nor U11154 (N_11154,N_10261,N_9876);
nand U11155 (N_11155,N_10014,N_9791);
nor U11156 (N_11156,N_9930,N_10260);
and U11157 (N_11157,N_10045,N_10010);
or U11158 (N_11158,N_9781,N_10251);
nand U11159 (N_11159,N_9890,N_9740);
or U11160 (N_11160,N_10351,N_10277);
and U11161 (N_11161,N_9647,N_9600);
nor U11162 (N_11162,N_9928,N_9989);
nand U11163 (N_11163,N_10219,N_10303);
and U11164 (N_11164,N_10283,N_10336);
xnor U11165 (N_11165,N_9615,N_10283);
nand U11166 (N_11166,N_9625,N_9760);
and U11167 (N_11167,N_10387,N_9766);
nor U11168 (N_11168,N_9807,N_9997);
and U11169 (N_11169,N_10320,N_9843);
nor U11170 (N_11170,N_10376,N_10100);
or U11171 (N_11171,N_9606,N_10048);
nand U11172 (N_11172,N_10105,N_10156);
and U11173 (N_11173,N_10146,N_10313);
or U11174 (N_11174,N_10057,N_10318);
nor U11175 (N_11175,N_9718,N_9711);
or U11176 (N_11176,N_9700,N_10390);
nand U11177 (N_11177,N_10168,N_10270);
and U11178 (N_11178,N_10078,N_10059);
or U11179 (N_11179,N_9932,N_9629);
nor U11180 (N_11180,N_9764,N_9688);
xor U11181 (N_11181,N_9936,N_10153);
nor U11182 (N_11182,N_9660,N_9799);
nand U11183 (N_11183,N_10198,N_10146);
xnor U11184 (N_11184,N_9711,N_10003);
nor U11185 (N_11185,N_9988,N_10275);
xor U11186 (N_11186,N_9772,N_9836);
nand U11187 (N_11187,N_9610,N_9924);
or U11188 (N_11188,N_9657,N_10023);
nand U11189 (N_11189,N_9920,N_9872);
or U11190 (N_11190,N_9859,N_10085);
xor U11191 (N_11191,N_9942,N_9823);
and U11192 (N_11192,N_9694,N_10020);
nor U11193 (N_11193,N_10028,N_10094);
and U11194 (N_11194,N_10381,N_9917);
nand U11195 (N_11195,N_10300,N_10185);
and U11196 (N_11196,N_9725,N_10056);
xnor U11197 (N_11197,N_9901,N_10119);
nand U11198 (N_11198,N_10163,N_9622);
or U11199 (N_11199,N_10250,N_9805);
nor U11200 (N_11200,N_11098,N_11081);
and U11201 (N_11201,N_11167,N_10679);
xor U11202 (N_11202,N_10880,N_10758);
or U11203 (N_11203,N_10937,N_10546);
xnor U11204 (N_11204,N_10452,N_10939);
or U11205 (N_11205,N_10798,N_10716);
nand U11206 (N_11206,N_11134,N_10478);
nor U11207 (N_11207,N_11046,N_11130);
xor U11208 (N_11208,N_10988,N_10487);
nor U11209 (N_11209,N_10582,N_11023);
nand U11210 (N_11210,N_10741,N_11156);
or U11211 (N_11211,N_11002,N_10540);
nand U11212 (N_11212,N_10753,N_10914);
nor U11213 (N_11213,N_11153,N_11168);
and U11214 (N_11214,N_11032,N_11048);
and U11215 (N_11215,N_10594,N_11113);
or U11216 (N_11216,N_10477,N_11013);
nand U11217 (N_11217,N_10521,N_10512);
nor U11218 (N_11218,N_10772,N_10488);
nand U11219 (N_11219,N_10974,N_10782);
or U11220 (N_11220,N_11196,N_11014);
nand U11221 (N_11221,N_10891,N_10998);
or U11222 (N_11222,N_10777,N_10976);
nor U11223 (N_11223,N_11079,N_10622);
or U11224 (N_11224,N_10514,N_10639);
nand U11225 (N_11225,N_11049,N_10474);
nand U11226 (N_11226,N_11179,N_10461);
xor U11227 (N_11227,N_10678,N_10931);
or U11228 (N_11228,N_11063,N_10444);
or U11229 (N_11229,N_10970,N_10655);
nand U11230 (N_11230,N_10971,N_10841);
nand U11231 (N_11231,N_10710,N_10797);
nand U11232 (N_11232,N_11111,N_10405);
or U11233 (N_11233,N_11084,N_11089);
or U11234 (N_11234,N_10996,N_10942);
and U11235 (N_11235,N_11067,N_11024);
or U11236 (N_11236,N_10447,N_11021);
or U11237 (N_11237,N_11030,N_10550);
nor U11238 (N_11238,N_11095,N_10602);
nor U11239 (N_11239,N_11136,N_10689);
xor U11240 (N_11240,N_10849,N_10975);
and U11241 (N_11241,N_10936,N_10822);
and U11242 (N_11242,N_10432,N_11012);
xnor U11243 (N_11243,N_10862,N_10744);
and U11244 (N_11244,N_10613,N_11114);
nor U11245 (N_11245,N_10544,N_10493);
and U11246 (N_11246,N_10462,N_10445);
or U11247 (N_11247,N_10569,N_10532);
xor U11248 (N_11248,N_10652,N_10811);
nand U11249 (N_11249,N_10497,N_11164);
nor U11250 (N_11250,N_10788,N_11019);
and U11251 (N_11251,N_11078,N_10981);
nand U11252 (N_11252,N_10732,N_10993);
and U11253 (N_11253,N_10752,N_10802);
or U11254 (N_11254,N_10449,N_10943);
nand U11255 (N_11255,N_11142,N_11007);
xor U11256 (N_11256,N_10940,N_10759);
nor U11257 (N_11257,N_10948,N_10906);
nor U11258 (N_11258,N_10623,N_10778);
and U11259 (N_11259,N_10875,N_10784);
and U11260 (N_11260,N_10792,N_10572);
or U11261 (N_11261,N_10756,N_10883);
nor U11262 (N_11262,N_10536,N_10677);
nand U11263 (N_11263,N_10469,N_10437);
nand U11264 (N_11264,N_11198,N_11151);
nand U11265 (N_11265,N_11141,N_11105);
nor U11266 (N_11266,N_11072,N_10593);
or U11267 (N_11267,N_10838,N_10787);
nor U11268 (N_11268,N_11120,N_11004);
or U11269 (N_11269,N_11177,N_10992);
and U11270 (N_11270,N_10507,N_11090);
and U11271 (N_11271,N_10921,N_10872);
nor U11272 (N_11272,N_10825,N_11119);
or U11273 (N_11273,N_11034,N_10610);
xor U11274 (N_11274,N_10587,N_10923);
and U11275 (N_11275,N_10706,N_10588);
nand U11276 (N_11276,N_10633,N_11045);
or U11277 (N_11277,N_11029,N_10694);
xnor U11278 (N_11278,N_10952,N_10486);
nor U11279 (N_11279,N_10728,N_11133);
nor U11280 (N_11280,N_10676,N_10684);
xnor U11281 (N_11281,N_10877,N_10799);
or U11282 (N_11282,N_10714,N_10554);
nand U11283 (N_11283,N_10808,N_10551);
nand U11284 (N_11284,N_10903,N_10769);
and U11285 (N_11285,N_10969,N_10928);
nor U11286 (N_11286,N_10977,N_11092);
xor U11287 (N_11287,N_10630,N_10905);
or U11288 (N_11288,N_10423,N_10803);
xor U11289 (N_11289,N_10505,N_10421);
or U11290 (N_11290,N_10909,N_10407);
nor U11291 (N_11291,N_10660,N_11188);
nand U11292 (N_11292,N_10653,N_11195);
or U11293 (N_11293,N_11077,N_10878);
and U11294 (N_11294,N_11165,N_10829);
or U11295 (N_11295,N_10763,N_10579);
xor U11296 (N_11296,N_11117,N_10483);
xnor U11297 (N_11297,N_10615,N_10597);
and U11298 (N_11298,N_11194,N_10738);
and U11299 (N_11299,N_10916,N_10501);
xor U11300 (N_11300,N_10583,N_10847);
or U11301 (N_11301,N_10665,N_11197);
or U11302 (N_11302,N_10561,N_10791);
nand U11303 (N_11303,N_10658,N_11093);
xnor U11304 (N_11304,N_11182,N_10956);
or U11305 (N_11305,N_10785,N_10637);
nor U11306 (N_11306,N_10767,N_11064);
xnor U11307 (N_11307,N_10672,N_10851);
nand U11308 (N_11308,N_10990,N_11010);
xnor U11309 (N_11309,N_11148,N_10754);
and U11310 (N_11310,N_11056,N_10688);
xor U11311 (N_11311,N_10635,N_10946);
or U11312 (N_11312,N_10647,N_10793);
or U11313 (N_11313,N_10446,N_10729);
nor U11314 (N_11314,N_10826,N_10901);
xnor U11315 (N_11315,N_10559,N_10605);
or U11316 (N_11316,N_11132,N_11037);
or U11317 (N_11317,N_10520,N_10962);
nand U11318 (N_11318,N_10629,N_10750);
xnor U11319 (N_11319,N_10814,N_11094);
and U11320 (N_11320,N_10459,N_11083);
nor U11321 (N_11321,N_10417,N_10831);
and U11322 (N_11322,N_10454,N_10641);
nand U11323 (N_11323,N_11074,N_10666);
and U11324 (N_11324,N_10453,N_11028);
xor U11325 (N_11325,N_10836,N_10620);
and U11326 (N_11326,N_10834,N_10489);
or U11327 (N_11327,N_10929,N_10595);
nand U11328 (N_11328,N_10618,N_10468);
nand U11329 (N_11329,N_10762,N_10567);
or U11330 (N_11330,N_10954,N_10542);
xnor U11331 (N_11331,N_11001,N_10528);
and U11332 (N_11332,N_11121,N_11144);
nor U11333 (N_11333,N_10959,N_10824);
nor U11334 (N_11334,N_10757,N_10693);
or U11335 (N_11335,N_10671,N_10917);
and U11336 (N_11336,N_10720,N_11099);
nor U11337 (N_11337,N_10853,N_10715);
nor U11338 (N_11338,N_10815,N_11088);
xnor U11339 (N_11339,N_11062,N_11190);
xor U11340 (N_11340,N_11073,N_11175);
nand U11341 (N_11341,N_10433,N_10403);
nor U11342 (N_11342,N_10661,N_10723);
nand U11343 (N_11343,N_10945,N_10491);
and U11344 (N_11344,N_10589,N_10857);
nor U11345 (N_11345,N_10850,N_10492);
and U11346 (N_11346,N_11000,N_11068);
nor U11347 (N_11347,N_10402,N_10794);
and U11348 (N_11348,N_10513,N_11086);
nand U11349 (N_11349,N_11158,N_10889);
and U11350 (N_11350,N_10702,N_10817);
or U11351 (N_11351,N_10746,N_11071);
and U11352 (N_11352,N_10899,N_10420);
or U11353 (N_11353,N_10621,N_11199);
xnor U11354 (N_11354,N_10854,N_10632);
xnor U11355 (N_11355,N_11127,N_10484);
nor U11356 (N_11356,N_10781,N_10460);
nand U11357 (N_11357,N_10575,N_11076);
nor U11358 (N_11358,N_10852,N_10692);
or U11359 (N_11359,N_10424,N_11118);
nand U11360 (N_11360,N_10504,N_10960);
xor U11361 (N_11361,N_10418,N_10711);
and U11362 (N_11362,N_10590,N_10966);
and U11363 (N_11363,N_10869,N_10830);
or U11364 (N_11364,N_10846,N_10570);
and U11365 (N_11365,N_11183,N_10411);
nor U11366 (N_11366,N_10519,N_10624);
and U11367 (N_11367,N_10807,N_10419);
nand U11368 (N_11368,N_10464,N_10922);
nor U11369 (N_11369,N_10832,N_11103);
and U11370 (N_11370,N_11091,N_10731);
nor U11371 (N_11371,N_10518,N_10596);
or U11372 (N_11372,N_10842,N_10691);
xor U11373 (N_11373,N_10481,N_10675);
and U11374 (N_11374,N_11069,N_11140);
xnor U11375 (N_11375,N_10627,N_10991);
nand U11376 (N_11376,N_11059,N_10743);
nor U11377 (N_11377,N_11128,N_10871);
xnor U11378 (N_11378,N_10810,N_10776);
and U11379 (N_11379,N_10455,N_10934);
xnor U11380 (N_11380,N_10896,N_10888);
nor U11381 (N_11381,N_10848,N_10668);
and U11382 (N_11382,N_10480,N_10973);
xor U11383 (N_11383,N_10450,N_10664);
nor U11384 (N_11384,N_11057,N_11163);
nor U11385 (N_11385,N_11184,N_11058);
xnor U11386 (N_11386,N_10577,N_10586);
nor U11387 (N_11387,N_11087,N_10795);
xnor U11388 (N_11388,N_11172,N_10547);
xor U11389 (N_11389,N_10773,N_10548);
or U11390 (N_11390,N_11160,N_10638);
nand U11391 (N_11391,N_10713,N_10642);
nor U11392 (N_11392,N_10409,N_11109);
xnor U11393 (N_11393,N_10584,N_11174);
nand U11394 (N_11394,N_10534,N_10733);
and U11395 (N_11395,N_10573,N_10765);
xnor U11396 (N_11396,N_10443,N_10428);
xnor U11397 (N_11397,N_10475,N_11041);
nor U11398 (N_11398,N_11112,N_10885);
nand U11399 (N_11399,N_11038,N_11003);
or U11400 (N_11400,N_10845,N_10541);
nor U11401 (N_11401,N_10707,N_10646);
nand U11402 (N_11402,N_11051,N_10574);
or U11403 (N_11403,N_11106,N_10495);
and U11404 (N_11404,N_11005,N_10631);
or U11405 (N_11405,N_11129,N_10525);
xor U11406 (N_11406,N_11047,N_10760);
and U11407 (N_11407,N_11017,N_10783);
nand U11408 (N_11408,N_11018,N_10537);
or U11409 (N_11409,N_10435,N_10912);
and U11410 (N_11410,N_10603,N_11027);
xnor U11411 (N_11411,N_10709,N_10606);
or U11412 (N_11412,N_10400,N_10681);
nor U11413 (N_11413,N_10961,N_10697);
or U11414 (N_11414,N_11178,N_10686);
nand U11415 (N_11415,N_11082,N_10699);
xnor U11416 (N_11416,N_10774,N_10545);
and U11417 (N_11417,N_10436,N_10565);
xor U11418 (N_11418,N_10724,N_11009);
nand U11419 (N_11419,N_10585,N_10751);
or U11420 (N_11420,N_10745,N_10806);
nand U11421 (N_11421,N_10893,N_10979);
xor U11422 (N_11422,N_10987,N_10401);
nor U11423 (N_11423,N_10619,N_10964);
nor U11424 (N_11424,N_10485,N_10986);
or U11425 (N_11425,N_10911,N_10951);
nand U11426 (N_11426,N_11025,N_10674);
and U11427 (N_11427,N_10415,N_10482);
and U11428 (N_11428,N_10616,N_10978);
and U11429 (N_11429,N_10566,N_11070);
nor U11430 (N_11430,N_10670,N_10982);
or U11431 (N_11431,N_10685,N_10790);
or U11432 (N_11432,N_10448,N_10835);
xnor U11433 (N_11433,N_11131,N_10989);
nand U11434 (N_11434,N_11169,N_10683);
or U11435 (N_11435,N_10673,N_10650);
and U11436 (N_11436,N_11191,N_10458);
xnor U11437 (N_11437,N_10933,N_11126);
nand U11438 (N_11438,N_10412,N_11102);
xnor U11439 (N_11439,N_11033,N_10500);
and U11440 (N_11440,N_10578,N_11139);
nand U11441 (N_11441,N_10898,N_10479);
nor U11442 (N_11442,N_11043,N_11104);
nor U11443 (N_11443,N_10434,N_10530);
nor U11444 (N_11444,N_10581,N_10611);
and U11445 (N_11445,N_10999,N_11040);
nand U11446 (N_11446,N_11185,N_10768);
nor U11447 (N_11447,N_10608,N_10995);
nand U11448 (N_11448,N_10737,N_10522);
nor U11449 (N_11449,N_10747,N_10703);
xor U11450 (N_11450,N_11044,N_10704);
and U11451 (N_11451,N_10859,N_10502);
nand U11452 (N_11452,N_10947,N_10749);
or U11453 (N_11453,N_10498,N_10687);
nand U11454 (N_11454,N_10680,N_11180);
and U11455 (N_11455,N_10963,N_10913);
nand U11456 (N_11456,N_10718,N_10531);
nand U11457 (N_11457,N_10427,N_11124);
or U11458 (N_11458,N_10628,N_10965);
nand U11459 (N_11459,N_10466,N_10843);
nand U11460 (N_11460,N_10508,N_10552);
xnor U11461 (N_11461,N_10667,N_10726);
and U11462 (N_11462,N_11036,N_10819);
and U11463 (N_11463,N_10614,N_11031);
nor U11464 (N_11464,N_10950,N_10844);
nand U11465 (N_11465,N_10972,N_10696);
and U11466 (N_11466,N_10556,N_10983);
xor U11467 (N_11467,N_10467,N_11149);
or U11468 (N_11468,N_10721,N_10980);
xor U11469 (N_11469,N_11054,N_10563);
nor U11470 (N_11470,N_10698,N_10509);
xor U11471 (N_11471,N_10821,N_10471);
and U11472 (N_11472,N_11015,N_10775);
and U11473 (N_11473,N_11186,N_10957);
or U11474 (N_11474,N_10408,N_10780);
xnor U11475 (N_11475,N_11161,N_10740);
and U11476 (N_11476,N_10813,N_10742);
and U11477 (N_11477,N_10555,N_11193);
or U11478 (N_11478,N_10727,N_10429);
and U11479 (N_11479,N_11125,N_10470);
xor U11480 (N_11480,N_11052,N_11006);
nor U11481 (N_11481,N_11022,N_10656);
and U11482 (N_11482,N_10890,N_10915);
nor U11483 (N_11483,N_11143,N_11181);
and U11484 (N_11484,N_10499,N_11173);
nand U11485 (N_11485,N_10410,N_11053);
nand U11486 (N_11486,N_10543,N_10626);
nand U11487 (N_11487,N_11110,N_10553);
xnor U11488 (N_11488,N_11116,N_11085);
and U11489 (N_11489,N_11026,N_10538);
and U11490 (N_11490,N_10604,N_10406);
nor U11491 (N_11491,N_10643,N_10907);
nor U11492 (N_11492,N_10918,N_10725);
nor U11493 (N_11493,N_10700,N_10645);
or U11494 (N_11494,N_11189,N_10837);
and U11495 (N_11495,N_10764,N_10796);
and U11496 (N_11496,N_10657,N_10465);
and U11497 (N_11497,N_11147,N_10490);
nor U11498 (N_11498,N_10695,N_10562);
and U11499 (N_11499,N_10456,N_10935);
and U11500 (N_11500,N_10730,N_10955);
nand U11501 (N_11501,N_10828,N_10904);
nor U11502 (N_11502,N_10708,N_10868);
or U11503 (N_11503,N_10476,N_10924);
or U11504 (N_11504,N_10812,N_10533);
or U11505 (N_11505,N_10870,N_10617);
or U11506 (N_11506,N_11080,N_10866);
xnor U11507 (N_11507,N_10422,N_10771);
and U11508 (N_11508,N_10598,N_10414);
nand U11509 (N_11509,N_10580,N_10425);
or U11510 (N_11510,N_11157,N_10515);
nand U11511 (N_11511,N_10413,N_11100);
or U11512 (N_11512,N_10734,N_10855);
nand U11513 (N_11513,N_11122,N_10997);
nand U11514 (N_11514,N_10705,N_10430);
and U11515 (N_11515,N_11039,N_10722);
or U11516 (N_11516,N_10517,N_10881);
or U11517 (N_11517,N_10920,N_11066);
and U11518 (N_11518,N_10431,N_10927);
nand U11519 (N_11519,N_10770,N_11060);
and U11520 (N_11520,N_11146,N_10600);
nor U11521 (N_11521,N_10930,N_10503);
nand U11522 (N_11522,N_10820,N_10659);
nand U11523 (N_11523,N_10669,N_11050);
nand U11524 (N_11524,N_11020,N_10644);
or U11525 (N_11525,N_11154,N_10463);
nor U11526 (N_11526,N_10856,N_10897);
and U11527 (N_11527,N_10648,N_10539);
xnor U11528 (N_11528,N_11171,N_10779);
xnor U11529 (N_11529,N_10416,N_10887);
nand U11530 (N_11530,N_10494,N_11137);
or U11531 (N_11531,N_10958,N_11166);
xor U11532 (N_11532,N_10506,N_10809);
or U11533 (N_11533,N_10524,N_11096);
xnor U11534 (N_11534,N_10404,N_10549);
and U11535 (N_11535,N_10527,N_10442);
or U11536 (N_11536,N_10892,N_10441);
xor U11537 (N_11537,N_10867,N_11176);
and U11538 (N_11538,N_11107,N_11152);
nor U11539 (N_11539,N_10900,N_10860);
nor U11540 (N_11540,N_10874,N_10560);
and U11541 (N_11541,N_10755,N_10879);
or U11542 (N_11542,N_10876,N_10861);
xnor U11543 (N_11543,N_10440,N_10649);
and U11544 (N_11544,N_10526,N_11008);
xor U11545 (N_11545,N_10511,N_10944);
nor U11546 (N_11546,N_10919,N_11145);
nor U11547 (N_11547,N_10523,N_10651);
nor U11548 (N_11548,N_10926,N_10805);
or U11549 (N_11549,N_11159,N_10910);
nand U11550 (N_11550,N_10558,N_10863);
nand U11551 (N_11551,N_11162,N_10748);
and U11552 (N_11552,N_11187,N_10908);
xor U11553 (N_11553,N_10865,N_11138);
nor U11554 (N_11554,N_10801,N_10636);
or U11555 (N_11555,N_10967,N_10858);
xor U11556 (N_11556,N_10496,N_10438);
xnor U11557 (N_11557,N_10833,N_11101);
nand U11558 (N_11558,N_10719,N_10557);
nor U11559 (N_11559,N_10457,N_11016);
xor U11560 (N_11560,N_10535,N_10902);
nor U11561 (N_11561,N_10564,N_10662);
or U11562 (N_11562,N_10607,N_10529);
nor U11563 (N_11563,N_10592,N_11055);
or U11564 (N_11564,N_11061,N_11075);
and U11565 (N_11565,N_10625,N_11135);
nand U11566 (N_11566,N_10968,N_10576);
and U11567 (N_11567,N_11155,N_10882);
and U11568 (N_11568,N_10766,N_10640);
nor U11569 (N_11569,N_10634,N_11011);
nor U11570 (N_11570,N_10816,N_11065);
xnor U11571 (N_11571,N_10886,N_11108);
xor U11572 (N_11572,N_11150,N_10839);
or U11573 (N_11573,N_10601,N_10571);
xnor U11574 (N_11574,N_10654,N_10823);
nand U11575 (N_11575,N_10932,N_10804);
or U11576 (N_11576,N_10840,N_10516);
nand U11577 (N_11577,N_11170,N_10473);
nor U11578 (N_11578,N_11115,N_10818);
and U11579 (N_11579,N_10712,N_10938);
and U11580 (N_11580,N_10472,N_10591);
xnor U11581 (N_11581,N_10735,N_10736);
or U11582 (N_11582,N_11123,N_10690);
nand U11583 (N_11583,N_10994,N_10827);
nor U11584 (N_11584,N_10786,N_10599);
or U11585 (N_11585,N_10800,N_10884);
and U11586 (N_11586,N_11192,N_10612);
or U11587 (N_11587,N_10761,N_10663);
xnor U11588 (N_11588,N_10426,N_11035);
xnor U11589 (N_11589,N_10451,N_10717);
nand U11590 (N_11590,N_10873,N_10439);
nand U11591 (N_11591,N_10568,N_10953);
nor U11592 (N_11592,N_10609,N_11097);
and U11593 (N_11593,N_10941,N_10701);
nand U11594 (N_11594,N_10739,N_11042);
and U11595 (N_11595,N_10895,N_10864);
or U11596 (N_11596,N_10510,N_10894);
xnor U11597 (N_11597,N_10949,N_10789);
nand U11598 (N_11598,N_10984,N_10985);
xnor U11599 (N_11599,N_10682,N_10925);
nor U11600 (N_11600,N_11119,N_10640);
or U11601 (N_11601,N_10465,N_10509);
xor U11602 (N_11602,N_10939,N_10803);
and U11603 (N_11603,N_11122,N_10559);
and U11604 (N_11604,N_10699,N_10718);
xnor U11605 (N_11605,N_11035,N_10831);
nand U11606 (N_11606,N_10780,N_11195);
nand U11607 (N_11607,N_10448,N_10655);
and U11608 (N_11608,N_10588,N_10895);
or U11609 (N_11609,N_10676,N_10434);
and U11610 (N_11610,N_10751,N_10425);
or U11611 (N_11611,N_10563,N_10814);
xor U11612 (N_11612,N_10621,N_10935);
nand U11613 (N_11613,N_10935,N_11099);
nor U11614 (N_11614,N_11024,N_10871);
and U11615 (N_11615,N_10443,N_10567);
nand U11616 (N_11616,N_10986,N_10974);
nand U11617 (N_11617,N_10752,N_11086);
xor U11618 (N_11618,N_10617,N_11118);
or U11619 (N_11619,N_10691,N_10904);
nand U11620 (N_11620,N_10790,N_11031);
nand U11621 (N_11621,N_10658,N_10474);
xnor U11622 (N_11622,N_10865,N_10980);
or U11623 (N_11623,N_10801,N_10672);
and U11624 (N_11624,N_10963,N_10862);
nand U11625 (N_11625,N_10698,N_11044);
xnor U11626 (N_11626,N_11023,N_10606);
nand U11627 (N_11627,N_10709,N_10833);
xnor U11628 (N_11628,N_10727,N_11058);
or U11629 (N_11629,N_10881,N_10833);
xor U11630 (N_11630,N_11103,N_10435);
and U11631 (N_11631,N_10925,N_10837);
and U11632 (N_11632,N_10403,N_10840);
nor U11633 (N_11633,N_10856,N_10682);
nor U11634 (N_11634,N_10926,N_11037);
and U11635 (N_11635,N_11147,N_10712);
nand U11636 (N_11636,N_10597,N_10541);
nand U11637 (N_11637,N_11137,N_10585);
xnor U11638 (N_11638,N_10752,N_10417);
nand U11639 (N_11639,N_11080,N_10562);
nor U11640 (N_11640,N_10827,N_10558);
xnor U11641 (N_11641,N_10823,N_10819);
nor U11642 (N_11642,N_10527,N_10675);
xnor U11643 (N_11643,N_10473,N_10921);
nor U11644 (N_11644,N_11017,N_11193);
xor U11645 (N_11645,N_11113,N_10612);
xnor U11646 (N_11646,N_10927,N_11041);
and U11647 (N_11647,N_10502,N_10858);
nor U11648 (N_11648,N_10604,N_10568);
and U11649 (N_11649,N_10778,N_11034);
nand U11650 (N_11650,N_11035,N_10796);
or U11651 (N_11651,N_10894,N_10670);
and U11652 (N_11652,N_10659,N_11091);
xnor U11653 (N_11653,N_10867,N_11023);
nand U11654 (N_11654,N_10700,N_11060);
nand U11655 (N_11655,N_10644,N_11087);
and U11656 (N_11656,N_10582,N_10566);
and U11657 (N_11657,N_10724,N_10514);
nand U11658 (N_11658,N_11069,N_10937);
or U11659 (N_11659,N_11117,N_11116);
nand U11660 (N_11660,N_10522,N_10955);
or U11661 (N_11661,N_10923,N_11013);
or U11662 (N_11662,N_11136,N_11188);
nor U11663 (N_11663,N_11002,N_11196);
xor U11664 (N_11664,N_10403,N_11126);
and U11665 (N_11665,N_10997,N_11114);
or U11666 (N_11666,N_10539,N_10644);
or U11667 (N_11667,N_10579,N_11048);
nor U11668 (N_11668,N_10409,N_10655);
xnor U11669 (N_11669,N_10800,N_10968);
xnor U11670 (N_11670,N_10429,N_10832);
or U11671 (N_11671,N_10586,N_10528);
nor U11672 (N_11672,N_10417,N_11149);
and U11673 (N_11673,N_10565,N_11046);
nor U11674 (N_11674,N_10607,N_11066);
nand U11675 (N_11675,N_10714,N_10568);
or U11676 (N_11676,N_10671,N_10582);
nand U11677 (N_11677,N_10830,N_11125);
nor U11678 (N_11678,N_10990,N_10844);
or U11679 (N_11679,N_10908,N_10731);
xnor U11680 (N_11680,N_10674,N_10532);
nand U11681 (N_11681,N_11040,N_11026);
and U11682 (N_11682,N_10641,N_10511);
or U11683 (N_11683,N_11001,N_10864);
and U11684 (N_11684,N_10539,N_10846);
xnor U11685 (N_11685,N_10423,N_10886);
or U11686 (N_11686,N_10858,N_10814);
xor U11687 (N_11687,N_10642,N_10967);
nor U11688 (N_11688,N_10730,N_11113);
and U11689 (N_11689,N_10667,N_10717);
xnor U11690 (N_11690,N_10603,N_11058);
nand U11691 (N_11691,N_10457,N_10608);
nand U11692 (N_11692,N_10737,N_10787);
xnor U11693 (N_11693,N_10843,N_10434);
nor U11694 (N_11694,N_11099,N_10628);
xnor U11695 (N_11695,N_10893,N_11192);
nand U11696 (N_11696,N_10490,N_11148);
nand U11697 (N_11697,N_10680,N_11099);
xnor U11698 (N_11698,N_10851,N_10922);
and U11699 (N_11699,N_10686,N_10413);
nand U11700 (N_11700,N_10863,N_10925);
and U11701 (N_11701,N_10418,N_10864);
xnor U11702 (N_11702,N_10484,N_10894);
or U11703 (N_11703,N_10480,N_10921);
or U11704 (N_11704,N_10768,N_10840);
or U11705 (N_11705,N_10916,N_10409);
nand U11706 (N_11706,N_10993,N_11103);
or U11707 (N_11707,N_10786,N_11079);
nand U11708 (N_11708,N_10730,N_10819);
nor U11709 (N_11709,N_10548,N_10787);
xor U11710 (N_11710,N_11138,N_11178);
xnor U11711 (N_11711,N_10523,N_11194);
or U11712 (N_11712,N_10899,N_11140);
nor U11713 (N_11713,N_10843,N_11159);
nand U11714 (N_11714,N_10567,N_10452);
and U11715 (N_11715,N_10784,N_11175);
nor U11716 (N_11716,N_10436,N_11137);
nand U11717 (N_11717,N_11019,N_10595);
xnor U11718 (N_11718,N_11087,N_10553);
and U11719 (N_11719,N_10800,N_10644);
nor U11720 (N_11720,N_10591,N_10507);
xor U11721 (N_11721,N_10929,N_10746);
nand U11722 (N_11722,N_10619,N_10925);
xnor U11723 (N_11723,N_11029,N_10627);
nor U11724 (N_11724,N_10903,N_10415);
and U11725 (N_11725,N_10874,N_10721);
nand U11726 (N_11726,N_10498,N_11140);
nand U11727 (N_11727,N_10992,N_10647);
nor U11728 (N_11728,N_11181,N_10582);
nand U11729 (N_11729,N_10641,N_10440);
nor U11730 (N_11730,N_10752,N_10708);
xnor U11731 (N_11731,N_11007,N_10717);
nand U11732 (N_11732,N_10486,N_10604);
and U11733 (N_11733,N_10531,N_10474);
nor U11734 (N_11734,N_10523,N_10971);
xor U11735 (N_11735,N_11153,N_11121);
or U11736 (N_11736,N_10844,N_10487);
nor U11737 (N_11737,N_11191,N_10564);
and U11738 (N_11738,N_10449,N_11062);
xor U11739 (N_11739,N_10720,N_10551);
or U11740 (N_11740,N_10719,N_11021);
nand U11741 (N_11741,N_10675,N_10410);
nand U11742 (N_11742,N_11160,N_10739);
nor U11743 (N_11743,N_11054,N_10941);
nand U11744 (N_11744,N_10910,N_10848);
xnor U11745 (N_11745,N_10778,N_10747);
xnor U11746 (N_11746,N_11138,N_10649);
nand U11747 (N_11747,N_10975,N_10969);
nand U11748 (N_11748,N_11035,N_10422);
and U11749 (N_11749,N_10607,N_11133);
nor U11750 (N_11750,N_10954,N_11026);
nand U11751 (N_11751,N_11119,N_10943);
and U11752 (N_11752,N_10644,N_10534);
or U11753 (N_11753,N_10998,N_10627);
or U11754 (N_11754,N_10723,N_11178);
nand U11755 (N_11755,N_10842,N_10674);
or U11756 (N_11756,N_11064,N_10649);
or U11757 (N_11757,N_10530,N_10494);
xnor U11758 (N_11758,N_10840,N_11179);
nand U11759 (N_11759,N_10860,N_10569);
and U11760 (N_11760,N_10964,N_10884);
and U11761 (N_11761,N_10750,N_10495);
and U11762 (N_11762,N_10936,N_10782);
xnor U11763 (N_11763,N_10530,N_11119);
and U11764 (N_11764,N_10703,N_10725);
xor U11765 (N_11765,N_11057,N_10461);
nand U11766 (N_11766,N_10656,N_10698);
nor U11767 (N_11767,N_11112,N_11123);
and U11768 (N_11768,N_11097,N_10830);
and U11769 (N_11769,N_10966,N_11135);
nor U11770 (N_11770,N_11195,N_11121);
xor U11771 (N_11771,N_11089,N_10811);
nor U11772 (N_11772,N_10541,N_11143);
nand U11773 (N_11773,N_11037,N_10624);
xor U11774 (N_11774,N_10963,N_10569);
or U11775 (N_11775,N_11033,N_10912);
nand U11776 (N_11776,N_10427,N_10866);
nand U11777 (N_11777,N_10937,N_11022);
nand U11778 (N_11778,N_10639,N_11015);
and U11779 (N_11779,N_10542,N_10826);
or U11780 (N_11780,N_10698,N_10568);
or U11781 (N_11781,N_10642,N_10411);
nor U11782 (N_11782,N_10713,N_10884);
xor U11783 (N_11783,N_10593,N_10899);
and U11784 (N_11784,N_11196,N_10840);
xnor U11785 (N_11785,N_10992,N_10786);
nand U11786 (N_11786,N_10520,N_11096);
xor U11787 (N_11787,N_10715,N_10881);
or U11788 (N_11788,N_10939,N_10923);
and U11789 (N_11789,N_11047,N_10764);
or U11790 (N_11790,N_10604,N_11135);
nor U11791 (N_11791,N_10643,N_11166);
xnor U11792 (N_11792,N_11197,N_10564);
xor U11793 (N_11793,N_10918,N_10547);
and U11794 (N_11794,N_10892,N_10673);
or U11795 (N_11795,N_10592,N_11195);
xnor U11796 (N_11796,N_11037,N_11048);
xor U11797 (N_11797,N_10902,N_10585);
or U11798 (N_11798,N_10612,N_11072);
or U11799 (N_11799,N_11131,N_10503);
nor U11800 (N_11800,N_10739,N_10765);
nand U11801 (N_11801,N_10646,N_10924);
nand U11802 (N_11802,N_10955,N_10509);
nand U11803 (N_11803,N_10903,N_11027);
or U11804 (N_11804,N_11123,N_11023);
and U11805 (N_11805,N_10798,N_10595);
and U11806 (N_11806,N_10778,N_10940);
and U11807 (N_11807,N_10861,N_10612);
xnor U11808 (N_11808,N_10586,N_10841);
xor U11809 (N_11809,N_10630,N_10514);
or U11810 (N_11810,N_10497,N_10695);
xor U11811 (N_11811,N_11137,N_10758);
and U11812 (N_11812,N_10610,N_10462);
nor U11813 (N_11813,N_10635,N_10928);
and U11814 (N_11814,N_10722,N_10830);
and U11815 (N_11815,N_10556,N_10531);
or U11816 (N_11816,N_10705,N_11157);
xor U11817 (N_11817,N_10957,N_11137);
xor U11818 (N_11818,N_10840,N_10681);
and U11819 (N_11819,N_11078,N_11156);
nor U11820 (N_11820,N_10818,N_10629);
or U11821 (N_11821,N_10540,N_10929);
and U11822 (N_11822,N_11115,N_10616);
or U11823 (N_11823,N_10949,N_11118);
xnor U11824 (N_11824,N_11010,N_10446);
nor U11825 (N_11825,N_11194,N_10965);
nor U11826 (N_11826,N_11073,N_10906);
and U11827 (N_11827,N_10842,N_10802);
nor U11828 (N_11828,N_10765,N_11031);
and U11829 (N_11829,N_10792,N_10695);
or U11830 (N_11830,N_11142,N_10791);
nor U11831 (N_11831,N_10987,N_10843);
nor U11832 (N_11832,N_10463,N_11036);
nand U11833 (N_11833,N_10626,N_10618);
or U11834 (N_11834,N_10649,N_10504);
nor U11835 (N_11835,N_10991,N_10704);
nand U11836 (N_11836,N_10761,N_11022);
or U11837 (N_11837,N_11187,N_10539);
and U11838 (N_11838,N_10956,N_10991);
nand U11839 (N_11839,N_11153,N_11199);
and U11840 (N_11840,N_11104,N_10484);
xor U11841 (N_11841,N_10667,N_11122);
and U11842 (N_11842,N_10869,N_10505);
nor U11843 (N_11843,N_10861,N_10661);
nand U11844 (N_11844,N_10987,N_11175);
nand U11845 (N_11845,N_11165,N_10841);
or U11846 (N_11846,N_10539,N_10826);
or U11847 (N_11847,N_10543,N_10562);
or U11848 (N_11848,N_10959,N_11172);
or U11849 (N_11849,N_10641,N_10522);
or U11850 (N_11850,N_10676,N_10726);
nor U11851 (N_11851,N_11134,N_10572);
xnor U11852 (N_11852,N_10923,N_11042);
xor U11853 (N_11853,N_10820,N_11014);
nor U11854 (N_11854,N_10715,N_11004);
nor U11855 (N_11855,N_10837,N_10828);
nand U11856 (N_11856,N_11167,N_11129);
nor U11857 (N_11857,N_10587,N_11001);
nand U11858 (N_11858,N_10708,N_10825);
or U11859 (N_11859,N_11157,N_11062);
nand U11860 (N_11860,N_10544,N_10632);
xnor U11861 (N_11861,N_10871,N_10755);
and U11862 (N_11862,N_10448,N_10577);
nand U11863 (N_11863,N_10406,N_10997);
or U11864 (N_11864,N_10835,N_10681);
and U11865 (N_11865,N_10515,N_10627);
xnor U11866 (N_11866,N_10580,N_10459);
nor U11867 (N_11867,N_10865,N_10756);
and U11868 (N_11868,N_10630,N_10834);
or U11869 (N_11869,N_10667,N_11015);
nor U11870 (N_11870,N_10428,N_10920);
xor U11871 (N_11871,N_10471,N_10968);
nand U11872 (N_11872,N_10996,N_10921);
nand U11873 (N_11873,N_10537,N_10694);
or U11874 (N_11874,N_10571,N_10407);
xor U11875 (N_11875,N_10952,N_10471);
xnor U11876 (N_11876,N_10533,N_10866);
nor U11877 (N_11877,N_10661,N_10959);
and U11878 (N_11878,N_10480,N_11158);
xnor U11879 (N_11879,N_10472,N_10690);
and U11880 (N_11880,N_10868,N_10455);
and U11881 (N_11881,N_10861,N_10564);
nor U11882 (N_11882,N_10451,N_10843);
xnor U11883 (N_11883,N_10489,N_10873);
and U11884 (N_11884,N_11094,N_11162);
or U11885 (N_11885,N_10691,N_10454);
nor U11886 (N_11886,N_10912,N_10920);
or U11887 (N_11887,N_11018,N_10738);
nor U11888 (N_11888,N_10862,N_10616);
nand U11889 (N_11889,N_10769,N_11183);
and U11890 (N_11890,N_10446,N_10438);
xor U11891 (N_11891,N_10577,N_10754);
nand U11892 (N_11892,N_11151,N_10796);
and U11893 (N_11893,N_10734,N_10675);
or U11894 (N_11894,N_11154,N_10613);
xnor U11895 (N_11895,N_10705,N_10684);
or U11896 (N_11896,N_11096,N_11126);
xor U11897 (N_11897,N_10968,N_10678);
nor U11898 (N_11898,N_11053,N_11106);
or U11899 (N_11899,N_10767,N_10769);
or U11900 (N_11900,N_11191,N_10732);
nor U11901 (N_11901,N_10829,N_11117);
or U11902 (N_11902,N_11102,N_10595);
and U11903 (N_11903,N_11014,N_11051);
or U11904 (N_11904,N_10486,N_10534);
nand U11905 (N_11905,N_10773,N_11025);
xor U11906 (N_11906,N_10617,N_10417);
and U11907 (N_11907,N_10952,N_10624);
nor U11908 (N_11908,N_10441,N_10422);
and U11909 (N_11909,N_10700,N_10670);
or U11910 (N_11910,N_10729,N_10669);
nor U11911 (N_11911,N_11093,N_10521);
nand U11912 (N_11912,N_10641,N_10689);
and U11913 (N_11913,N_10550,N_10994);
xnor U11914 (N_11914,N_10570,N_10787);
or U11915 (N_11915,N_10555,N_10680);
or U11916 (N_11916,N_11119,N_10874);
xor U11917 (N_11917,N_10868,N_11083);
and U11918 (N_11918,N_10713,N_10931);
nand U11919 (N_11919,N_10901,N_10505);
xnor U11920 (N_11920,N_10925,N_11114);
or U11921 (N_11921,N_11150,N_10589);
or U11922 (N_11922,N_10726,N_11172);
nand U11923 (N_11923,N_10669,N_10862);
nand U11924 (N_11924,N_10839,N_10972);
and U11925 (N_11925,N_10651,N_10491);
nand U11926 (N_11926,N_10905,N_11157);
nor U11927 (N_11927,N_10531,N_10511);
xnor U11928 (N_11928,N_10949,N_10682);
and U11929 (N_11929,N_10719,N_10564);
nand U11930 (N_11930,N_10874,N_10782);
or U11931 (N_11931,N_10505,N_10590);
or U11932 (N_11932,N_11016,N_10671);
and U11933 (N_11933,N_10578,N_11113);
or U11934 (N_11934,N_11095,N_10937);
xnor U11935 (N_11935,N_10924,N_10526);
xor U11936 (N_11936,N_10838,N_10613);
and U11937 (N_11937,N_10905,N_10412);
nand U11938 (N_11938,N_10877,N_11094);
nand U11939 (N_11939,N_11066,N_10662);
nand U11940 (N_11940,N_11143,N_10730);
nor U11941 (N_11941,N_10810,N_10959);
nand U11942 (N_11942,N_10953,N_10669);
nand U11943 (N_11943,N_11019,N_11145);
or U11944 (N_11944,N_10955,N_11021);
nor U11945 (N_11945,N_10846,N_10727);
xor U11946 (N_11946,N_10680,N_10617);
xnor U11947 (N_11947,N_10440,N_11072);
or U11948 (N_11948,N_10544,N_10893);
nor U11949 (N_11949,N_10549,N_11113);
or U11950 (N_11950,N_10494,N_10413);
xor U11951 (N_11951,N_11144,N_10894);
nor U11952 (N_11952,N_10714,N_10652);
and U11953 (N_11953,N_10891,N_10968);
nand U11954 (N_11954,N_10724,N_10473);
and U11955 (N_11955,N_10993,N_10789);
xnor U11956 (N_11956,N_10900,N_10471);
or U11957 (N_11957,N_10566,N_10449);
or U11958 (N_11958,N_11157,N_10808);
xnor U11959 (N_11959,N_11170,N_10487);
xor U11960 (N_11960,N_10765,N_10525);
and U11961 (N_11961,N_10606,N_10640);
and U11962 (N_11962,N_10731,N_10838);
and U11963 (N_11963,N_10729,N_10442);
or U11964 (N_11964,N_10998,N_10747);
xnor U11965 (N_11965,N_11087,N_10787);
nand U11966 (N_11966,N_11110,N_10561);
or U11967 (N_11967,N_11160,N_10528);
and U11968 (N_11968,N_10796,N_11162);
xor U11969 (N_11969,N_10431,N_10675);
xor U11970 (N_11970,N_10679,N_11093);
and U11971 (N_11971,N_10960,N_10822);
xor U11972 (N_11972,N_10466,N_10784);
nand U11973 (N_11973,N_10429,N_10427);
nor U11974 (N_11974,N_11009,N_10969);
xnor U11975 (N_11975,N_11158,N_11168);
and U11976 (N_11976,N_10795,N_10512);
nor U11977 (N_11977,N_10828,N_10818);
nor U11978 (N_11978,N_10415,N_10660);
or U11979 (N_11979,N_11198,N_10879);
xor U11980 (N_11980,N_10974,N_10466);
or U11981 (N_11981,N_10982,N_10737);
or U11982 (N_11982,N_11046,N_10477);
nor U11983 (N_11983,N_11052,N_10839);
nor U11984 (N_11984,N_10438,N_11025);
and U11985 (N_11985,N_10687,N_10650);
and U11986 (N_11986,N_10571,N_10995);
nor U11987 (N_11987,N_10875,N_10661);
or U11988 (N_11988,N_11029,N_11020);
nor U11989 (N_11989,N_11082,N_10783);
or U11990 (N_11990,N_10829,N_10759);
nor U11991 (N_11991,N_10816,N_10927);
and U11992 (N_11992,N_10421,N_10609);
and U11993 (N_11993,N_10912,N_10456);
xor U11994 (N_11994,N_10559,N_10908);
and U11995 (N_11995,N_11093,N_10836);
nand U11996 (N_11996,N_10511,N_10425);
xor U11997 (N_11997,N_11101,N_10959);
nor U11998 (N_11998,N_10464,N_10953);
xor U11999 (N_11999,N_10699,N_10803);
xnor U12000 (N_12000,N_11467,N_11595);
or U12001 (N_12001,N_11934,N_11399);
or U12002 (N_12002,N_11861,N_11333);
nor U12003 (N_12003,N_11327,N_11297);
nor U12004 (N_12004,N_11310,N_11279);
or U12005 (N_12005,N_11375,N_11920);
nand U12006 (N_12006,N_11721,N_11306);
nor U12007 (N_12007,N_11845,N_11982);
nor U12008 (N_12008,N_11722,N_11970);
xor U12009 (N_12009,N_11303,N_11283);
nand U12010 (N_12010,N_11864,N_11299);
xnor U12011 (N_12011,N_11581,N_11538);
nand U12012 (N_12012,N_11727,N_11505);
and U12013 (N_12013,N_11342,N_11256);
xor U12014 (N_12014,N_11961,N_11205);
nand U12015 (N_12015,N_11824,N_11856);
nor U12016 (N_12016,N_11708,N_11573);
xnor U12017 (N_12017,N_11387,N_11849);
nor U12018 (N_12018,N_11648,N_11755);
or U12019 (N_12019,N_11221,N_11971);
xor U12020 (N_12020,N_11656,N_11707);
nand U12021 (N_12021,N_11698,N_11880);
or U12022 (N_12022,N_11913,N_11560);
nor U12023 (N_12023,N_11989,N_11368);
nor U12024 (N_12024,N_11705,N_11300);
nand U12025 (N_12025,N_11572,N_11816);
nand U12026 (N_12026,N_11246,N_11808);
nand U12027 (N_12027,N_11544,N_11263);
or U12028 (N_12028,N_11392,N_11959);
or U12029 (N_12029,N_11833,N_11967);
or U12030 (N_12030,N_11366,N_11529);
and U12031 (N_12031,N_11703,N_11650);
and U12032 (N_12032,N_11582,N_11556);
or U12033 (N_12033,N_11753,N_11957);
nand U12034 (N_12034,N_11424,N_11740);
nand U12035 (N_12035,N_11397,N_11302);
nor U12036 (N_12036,N_11615,N_11713);
xor U12037 (N_12037,N_11429,N_11382);
nand U12038 (N_12038,N_11769,N_11752);
and U12039 (N_12039,N_11576,N_11909);
xnor U12040 (N_12040,N_11348,N_11594);
nand U12041 (N_12041,N_11364,N_11887);
nand U12042 (N_12042,N_11886,N_11749);
and U12043 (N_12043,N_11642,N_11453);
nand U12044 (N_12044,N_11519,N_11501);
and U12045 (N_12045,N_11676,N_11285);
or U12046 (N_12046,N_11686,N_11253);
nand U12047 (N_12047,N_11267,N_11475);
nand U12048 (N_12048,N_11549,N_11380);
or U12049 (N_12049,N_11464,N_11811);
or U12050 (N_12050,N_11893,N_11930);
xnor U12051 (N_12051,N_11292,N_11684);
nor U12052 (N_12052,N_11803,N_11349);
nor U12053 (N_12053,N_11953,N_11454);
nor U12054 (N_12054,N_11580,N_11249);
or U12055 (N_12055,N_11428,N_11626);
nand U12056 (N_12056,N_11491,N_11559);
nand U12057 (N_12057,N_11487,N_11513);
nand U12058 (N_12058,N_11717,N_11350);
nand U12059 (N_12059,N_11590,N_11683);
nor U12060 (N_12060,N_11810,N_11432);
nand U12061 (N_12061,N_11696,N_11881);
or U12062 (N_12062,N_11756,N_11272);
and U12063 (N_12063,N_11919,N_11438);
nand U12064 (N_12064,N_11217,N_11578);
nor U12065 (N_12065,N_11984,N_11687);
or U12066 (N_12066,N_11660,N_11916);
xnor U12067 (N_12067,N_11227,N_11782);
nand U12068 (N_12068,N_11914,N_11830);
and U12069 (N_12069,N_11295,N_11461);
or U12070 (N_12070,N_11284,N_11935);
xor U12071 (N_12071,N_11895,N_11430);
and U12072 (N_12072,N_11431,N_11484);
nand U12073 (N_12073,N_11635,N_11439);
nand U12074 (N_12074,N_11710,N_11558);
or U12075 (N_12075,N_11613,N_11821);
xor U12076 (N_12076,N_11609,N_11669);
nor U12077 (N_12077,N_11465,N_11264);
xnor U12078 (N_12078,N_11663,N_11321);
and U12079 (N_12079,N_11328,N_11606);
and U12080 (N_12080,N_11618,N_11335);
nand U12081 (N_12081,N_11904,N_11602);
nor U12082 (N_12082,N_11421,N_11346);
nor U12083 (N_12083,N_11975,N_11992);
or U12084 (N_12084,N_11825,N_11437);
nand U12085 (N_12085,N_11241,N_11879);
nor U12086 (N_12086,N_11492,N_11416);
nand U12087 (N_12087,N_11462,N_11860);
or U12088 (N_12088,N_11472,N_11903);
and U12089 (N_12089,N_11608,N_11712);
nor U12090 (N_12090,N_11983,N_11890);
or U12091 (N_12091,N_11786,N_11770);
nand U12092 (N_12092,N_11807,N_11456);
or U12093 (N_12093,N_11357,N_11406);
nand U12094 (N_12094,N_11469,N_11912);
and U12095 (N_12095,N_11885,N_11535);
and U12096 (N_12096,N_11367,N_11981);
nand U12097 (N_12097,N_11665,N_11378);
or U12098 (N_12098,N_11802,N_11353);
xnor U12099 (N_12099,N_11514,N_11381);
nand U12100 (N_12100,N_11557,N_11979);
or U12101 (N_12101,N_11204,N_11837);
or U12102 (N_12102,N_11695,N_11471);
or U12103 (N_12103,N_11385,N_11488);
xnor U12104 (N_12104,N_11985,N_11443);
or U12105 (N_12105,N_11815,N_11685);
and U12106 (N_12106,N_11497,N_11702);
and U12107 (N_12107,N_11878,N_11835);
nand U12108 (N_12108,N_11675,N_11628);
nor U12109 (N_12109,N_11719,N_11948);
xnor U12110 (N_12110,N_11334,N_11208);
and U12111 (N_12111,N_11804,N_11638);
nand U12112 (N_12112,N_11330,N_11842);
and U12113 (N_12113,N_11575,N_11289);
or U12114 (N_12114,N_11248,N_11616);
nor U12115 (N_12115,N_11261,N_11737);
xnor U12116 (N_12116,N_11760,N_11372);
nand U12117 (N_12117,N_11963,N_11525);
xnor U12118 (N_12118,N_11344,N_11460);
and U12119 (N_12119,N_11901,N_11278);
nand U12120 (N_12120,N_11945,N_11444);
and U12121 (N_12121,N_11990,N_11257);
nand U12122 (N_12122,N_11796,N_11401);
nor U12123 (N_12123,N_11447,N_11341);
xnor U12124 (N_12124,N_11569,N_11723);
nor U12125 (N_12125,N_11458,N_11924);
xnor U12126 (N_12126,N_11792,N_11817);
or U12127 (N_12127,N_11550,N_11907);
nand U12128 (N_12128,N_11905,N_11286);
nand U12129 (N_12129,N_11840,N_11280);
nand U12130 (N_12130,N_11900,N_11269);
nor U12131 (N_12131,N_11388,N_11528);
nor U12132 (N_12132,N_11258,N_11250);
xnor U12133 (N_12133,N_11800,N_11345);
nor U12134 (N_12134,N_11466,N_11522);
and U12135 (N_12135,N_11584,N_11474);
xnor U12136 (N_12136,N_11697,N_11997);
nand U12137 (N_12137,N_11718,N_11586);
and U12138 (N_12138,N_11503,N_11694);
xnor U12139 (N_12139,N_11340,N_11892);
nand U12140 (N_12140,N_11242,N_11754);
or U12141 (N_12141,N_11910,N_11894);
and U12142 (N_12142,N_11667,N_11527);
xor U12143 (N_12143,N_11778,N_11658);
or U12144 (N_12144,N_11511,N_11724);
nand U12145 (N_12145,N_11938,N_11852);
xor U12146 (N_12146,N_11974,N_11479);
and U12147 (N_12147,N_11746,N_11361);
and U12148 (N_12148,N_11932,N_11728);
and U12149 (N_12149,N_11906,N_11631);
and U12150 (N_12150,N_11747,N_11379);
xor U12151 (N_12151,N_11795,N_11603);
nor U12152 (N_12152,N_11352,N_11389);
and U12153 (N_12153,N_11681,N_11855);
nor U12154 (N_12154,N_11636,N_11598);
nand U12155 (N_12155,N_11709,N_11275);
nand U12156 (N_12156,N_11309,N_11790);
nand U12157 (N_12157,N_11794,N_11551);
and U12158 (N_12158,N_11831,N_11536);
nand U12159 (N_12159,N_11733,N_11741);
nand U12160 (N_12160,N_11415,N_11599);
xnor U12161 (N_12161,N_11771,N_11926);
nor U12162 (N_12162,N_11617,N_11827);
nand U12163 (N_12163,N_11254,N_11597);
and U12164 (N_12164,N_11287,N_11570);
or U12165 (N_12165,N_11425,N_11200);
and U12166 (N_12166,N_11374,N_11412);
nand U12167 (N_12167,N_11515,N_11748);
nand U12168 (N_12168,N_11918,N_11772);
xnor U12169 (N_12169,N_11784,N_11470);
or U12170 (N_12170,N_11496,N_11214);
nor U12171 (N_12171,N_11689,N_11644);
nor U12172 (N_12172,N_11371,N_11478);
nand U12173 (N_12173,N_11777,N_11414);
nand U12174 (N_12174,N_11859,N_11632);
nor U12175 (N_12175,N_11629,N_11716);
or U12176 (N_12176,N_11941,N_11902);
nor U12177 (N_12177,N_11206,N_11678);
nor U12178 (N_12178,N_11925,N_11779);
or U12179 (N_12179,N_11620,N_11441);
nand U12180 (N_12180,N_11383,N_11884);
nor U12181 (N_12181,N_11624,N_11225);
nand U12182 (N_12182,N_11301,N_11543);
or U12183 (N_12183,N_11435,N_11585);
or U12184 (N_12184,N_11679,N_11991);
or U12185 (N_12185,N_11823,N_11498);
or U12186 (N_12186,N_11502,N_11715);
xor U12187 (N_12187,N_11818,N_11596);
nand U12188 (N_12188,N_11838,N_11661);
and U12189 (N_12189,N_11673,N_11555);
xor U12190 (N_12190,N_11314,N_11493);
or U12191 (N_12191,N_11672,N_11373);
or U12192 (N_12192,N_11571,N_11944);
xor U12193 (N_12193,N_11420,N_11977);
and U12194 (N_12194,N_11291,N_11995);
xor U12195 (N_12195,N_11362,N_11922);
nor U12196 (N_12196,N_11547,N_11757);
nand U12197 (N_12197,N_11858,N_11523);
and U12198 (N_12198,N_11394,N_11245);
nor U12199 (N_12199,N_11896,N_11288);
nor U12200 (N_12200,N_11232,N_11294);
nor U12201 (N_12201,N_11876,N_11481);
xnor U12202 (N_12202,N_11230,N_11396);
or U12203 (N_12203,N_11325,N_11561);
or U12204 (N_12204,N_11812,N_11468);
xnor U12205 (N_12205,N_11237,N_11736);
xor U12206 (N_12206,N_11316,N_11434);
xnor U12207 (N_12207,N_11423,N_11231);
nand U12208 (N_12208,N_11480,N_11775);
nand U12209 (N_12209,N_11908,N_11391);
nand U12210 (N_12210,N_11994,N_11298);
nand U12211 (N_12211,N_11701,N_11645);
xor U12212 (N_12212,N_11273,N_11593);
nand U12213 (N_12213,N_11854,N_11542);
nand U12214 (N_12214,N_11395,N_11370);
or U12215 (N_12215,N_11730,N_11870);
nand U12216 (N_12216,N_11869,N_11268);
nand U12217 (N_12217,N_11336,N_11962);
xor U12218 (N_12218,N_11212,N_11442);
xor U12219 (N_12219,N_11448,N_11940);
nand U12220 (N_12220,N_11220,N_11873);
and U12221 (N_12221,N_11343,N_11518);
nor U12222 (N_12222,N_11836,N_11201);
or U12223 (N_12223,N_11332,N_11408);
nor U12224 (N_12224,N_11911,N_11766);
or U12225 (N_12225,N_11634,N_11751);
nand U12226 (N_12226,N_11577,N_11347);
or U12227 (N_12227,N_11931,N_11304);
and U12228 (N_12228,N_11937,N_11251);
nor U12229 (N_12229,N_11600,N_11972);
and U12230 (N_12230,N_11773,N_11252);
or U12231 (N_12231,N_11489,N_11574);
or U12232 (N_12232,N_11563,N_11623);
or U12233 (N_12233,N_11376,N_11764);
and U12234 (N_12234,N_11483,N_11318);
nor U12235 (N_12235,N_11791,N_11998);
nor U12236 (N_12236,N_11568,N_11240);
or U12237 (N_12237,N_11589,N_11671);
or U12238 (N_12238,N_11988,N_11567);
xor U12239 (N_12239,N_11915,N_11674);
and U12240 (N_12240,N_11726,N_11356);
nand U12241 (N_12241,N_11780,N_11761);
nand U12242 (N_12242,N_11459,N_11649);
and U12243 (N_12243,N_11311,N_11235);
xor U12244 (N_12244,N_11476,N_11954);
and U12245 (N_12245,N_11734,N_11512);
nand U12246 (N_12246,N_11882,N_11946);
nand U12247 (N_12247,N_11765,N_11211);
nor U12248 (N_12248,N_11405,N_11739);
xnor U12249 (N_12249,N_11517,N_11844);
or U12250 (N_12250,N_11260,N_11643);
nor U12251 (N_12251,N_11565,N_11612);
nand U12252 (N_12252,N_11704,N_11693);
xor U12253 (N_12253,N_11729,N_11244);
xor U12254 (N_12254,N_11411,N_11947);
or U12255 (N_12255,N_11863,N_11768);
xnor U12256 (N_12256,N_11843,N_11516);
or U12257 (N_12257,N_11452,N_11339);
and U12258 (N_12258,N_11851,N_11744);
and U12259 (N_12259,N_11323,N_11846);
nor U12260 (N_12260,N_11419,N_11714);
xor U12261 (N_12261,N_11814,N_11952);
and U12262 (N_12262,N_11546,N_11207);
xnor U12263 (N_12263,N_11797,N_11731);
and U12264 (N_12264,N_11641,N_11363);
nand U12265 (N_12265,N_11742,N_11354);
or U12266 (N_12266,N_11446,N_11545);
nand U12267 (N_12267,N_11562,N_11874);
nor U12268 (N_12268,N_11664,N_11520);
xor U12269 (N_12269,N_11451,N_11706);
and U12270 (N_12270,N_11993,N_11725);
xor U12271 (N_12271,N_11233,N_11588);
or U12272 (N_12272,N_11677,N_11711);
or U12273 (N_12273,N_11923,N_11688);
nor U12274 (N_12274,N_11738,N_11322);
xor U12275 (N_12275,N_11243,N_11999);
and U12276 (N_12276,N_11450,N_11331);
nor U12277 (N_12277,N_11276,N_11506);
or U12278 (N_12278,N_11407,N_11533);
and U12279 (N_12279,N_11592,N_11477);
nand U12280 (N_12280,N_11619,N_11317);
nor U12281 (N_12281,N_11942,N_11690);
nand U12282 (N_12282,N_11427,N_11889);
nor U12283 (N_12283,N_11866,N_11789);
nor U12284 (N_12284,N_11735,N_11899);
xor U12285 (N_12285,N_11313,N_11202);
or U12286 (N_12286,N_11762,N_11891);
and U12287 (N_12287,N_11282,N_11819);
nor U12288 (N_12288,N_11591,N_11554);
nor U12289 (N_12289,N_11255,N_11524);
xnor U12290 (N_12290,N_11871,N_11670);
and U12291 (N_12291,N_11607,N_11351);
nor U12292 (N_12292,N_11720,N_11743);
and U12293 (N_12293,N_11308,N_11978);
or U12294 (N_12294,N_11965,N_11783);
xnor U12295 (N_12295,N_11700,N_11320);
nand U12296 (N_12296,N_11312,N_11358);
nor U12297 (N_12297,N_11949,N_11950);
xor U12298 (N_12298,N_11605,N_11865);
nand U12299 (N_12299,N_11500,N_11763);
xnor U12300 (N_12300,N_11622,N_11386);
xor U12301 (N_12301,N_11987,N_11247);
nand U12302 (N_12302,N_11234,N_11929);
nand U12303 (N_12303,N_11531,N_11402);
nand U12304 (N_12304,N_11315,N_11759);
nand U12305 (N_12305,N_11504,N_11410);
nand U12306 (N_12306,N_11973,N_11359);
or U12307 (N_12307,N_11485,N_11223);
nand U12308 (N_12308,N_11583,N_11473);
or U12309 (N_12309,N_11651,N_11564);
nand U12310 (N_12310,N_11440,N_11787);
nor U12311 (N_12311,N_11621,N_11839);
nand U12312 (N_12312,N_11270,N_11857);
and U12313 (N_12313,N_11262,N_11828);
nor U12314 (N_12314,N_11933,N_11449);
and U12315 (N_12315,N_11625,N_11548);
or U12316 (N_12316,N_11463,N_11976);
xor U12317 (N_12317,N_11939,N_11307);
nand U12318 (N_12318,N_11680,N_11521);
xnor U12319 (N_12319,N_11541,N_11426);
or U12320 (N_12320,N_11277,N_11875);
and U12321 (N_12321,N_11652,N_11668);
and U12322 (N_12322,N_11526,N_11611);
xor U12323 (N_12323,N_11691,N_11537);
nor U12324 (N_12324,N_11850,N_11457);
nor U12325 (N_12325,N_11682,N_11813);
nand U12326 (N_12326,N_11219,N_11337);
nor U12327 (N_12327,N_11785,N_11964);
or U12328 (N_12328,N_11960,N_11360);
xnor U12329 (N_12329,N_11654,N_11579);
or U12330 (N_12330,N_11210,N_11610);
and U12331 (N_12331,N_11822,N_11883);
nor U12332 (N_12332,N_11601,N_11482);
or U12333 (N_12333,N_11627,N_11888);
or U12334 (N_12334,N_11490,N_11239);
nand U12335 (N_12335,N_11951,N_11820);
or U12336 (N_12336,N_11653,N_11226);
nor U12337 (N_12337,N_11774,N_11604);
nor U12338 (N_12338,N_11928,N_11418);
nor U12339 (N_12339,N_11848,N_11867);
nand U12340 (N_12340,N_11305,N_11216);
xor U12341 (N_12341,N_11955,N_11637);
or U12342 (N_12342,N_11417,N_11980);
nor U12343 (N_12343,N_11877,N_11324);
nand U12344 (N_12344,N_11403,N_11445);
nand U12345 (N_12345,N_11495,N_11228);
xnor U12346 (N_12346,N_11968,N_11898);
nor U12347 (N_12347,N_11218,N_11647);
and U12348 (N_12348,N_11338,N_11969);
or U12349 (N_12349,N_11433,N_11390);
and U12350 (N_12350,N_11587,N_11566);
xnor U12351 (N_12351,N_11832,N_11532);
nand U12352 (N_12352,N_11266,N_11767);
nand U12353 (N_12353,N_11826,N_11238);
xor U12354 (N_12354,N_11404,N_11805);
nand U12355 (N_12355,N_11326,N_11509);
nand U12356 (N_12356,N_11732,N_11921);
or U12357 (N_12357,N_11369,N_11209);
xnor U12358 (N_12358,N_11927,N_11868);
and U12359 (N_12359,N_11862,N_11499);
nand U12360 (N_12360,N_11966,N_11274);
or U12361 (N_12361,N_11986,N_11943);
or U12362 (N_12362,N_11553,N_11917);
nor U12363 (N_12363,N_11809,N_11409);
nand U12364 (N_12364,N_11692,N_11265);
and U12365 (N_12365,N_11224,N_11666);
nand U12366 (N_12366,N_11834,N_11958);
nor U12367 (N_12367,N_11781,N_11776);
xnor U12368 (N_12368,N_11281,N_11793);
xnor U12369 (N_12369,N_11398,N_11841);
and U12370 (N_12370,N_11847,N_11897);
or U12371 (N_12371,N_11853,N_11639);
xnor U12372 (N_12372,N_11745,N_11633);
and U12373 (N_12373,N_11540,N_11799);
and U12374 (N_12374,N_11494,N_11455);
xor U12375 (N_12375,N_11229,N_11215);
and U12376 (N_12376,N_11662,N_11659);
or U12377 (N_12377,N_11655,N_11872);
or U12378 (N_12378,N_11750,N_11507);
nor U12379 (N_12379,N_11806,N_11319);
xnor U12380 (N_12380,N_11956,N_11436);
or U12381 (N_12381,N_11801,N_11699);
xnor U12382 (N_12382,N_11222,N_11614);
or U12383 (N_12383,N_11377,N_11422);
nand U12384 (N_12384,N_11508,N_11630);
or U12385 (N_12385,N_11530,N_11290);
xnor U12386 (N_12386,N_11646,N_11384);
and U12387 (N_12387,N_11829,N_11640);
or U12388 (N_12388,N_11203,N_11329);
nor U12389 (N_12389,N_11259,N_11510);
xnor U12390 (N_12390,N_11293,N_11552);
xnor U12391 (N_12391,N_11355,N_11996);
nand U12392 (N_12392,N_11413,N_11539);
and U12393 (N_12393,N_11393,N_11788);
or U12394 (N_12394,N_11213,N_11400);
nor U12395 (N_12395,N_11798,N_11296);
nand U12396 (N_12396,N_11936,N_11657);
nor U12397 (N_12397,N_11486,N_11236);
nand U12398 (N_12398,N_11365,N_11271);
nand U12399 (N_12399,N_11758,N_11534);
nand U12400 (N_12400,N_11556,N_11647);
nand U12401 (N_12401,N_11928,N_11925);
nand U12402 (N_12402,N_11762,N_11237);
xor U12403 (N_12403,N_11541,N_11564);
nand U12404 (N_12404,N_11828,N_11490);
xnor U12405 (N_12405,N_11322,N_11572);
nand U12406 (N_12406,N_11878,N_11791);
nor U12407 (N_12407,N_11952,N_11369);
nor U12408 (N_12408,N_11732,N_11745);
and U12409 (N_12409,N_11273,N_11284);
nand U12410 (N_12410,N_11397,N_11547);
or U12411 (N_12411,N_11638,N_11239);
nor U12412 (N_12412,N_11501,N_11413);
nand U12413 (N_12413,N_11355,N_11790);
nor U12414 (N_12414,N_11614,N_11674);
or U12415 (N_12415,N_11878,N_11739);
or U12416 (N_12416,N_11437,N_11664);
nor U12417 (N_12417,N_11503,N_11233);
or U12418 (N_12418,N_11547,N_11253);
nor U12419 (N_12419,N_11791,N_11618);
and U12420 (N_12420,N_11372,N_11683);
and U12421 (N_12421,N_11499,N_11637);
and U12422 (N_12422,N_11627,N_11834);
nor U12423 (N_12423,N_11275,N_11284);
nand U12424 (N_12424,N_11566,N_11792);
nand U12425 (N_12425,N_11383,N_11342);
and U12426 (N_12426,N_11934,N_11259);
or U12427 (N_12427,N_11616,N_11218);
or U12428 (N_12428,N_11835,N_11501);
or U12429 (N_12429,N_11413,N_11287);
nor U12430 (N_12430,N_11724,N_11911);
xor U12431 (N_12431,N_11543,N_11286);
nor U12432 (N_12432,N_11732,N_11354);
xnor U12433 (N_12433,N_11746,N_11809);
and U12434 (N_12434,N_11580,N_11611);
xor U12435 (N_12435,N_11699,N_11966);
and U12436 (N_12436,N_11425,N_11475);
or U12437 (N_12437,N_11494,N_11667);
nand U12438 (N_12438,N_11221,N_11623);
nor U12439 (N_12439,N_11628,N_11298);
nand U12440 (N_12440,N_11399,N_11686);
and U12441 (N_12441,N_11412,N_11982);
xnor U12442 (N_12442,N_11965,N_11648);
or U12443 (N_12443,N_11226,N_11495);
or U12444 (N_12444,N_11389,N_11468);
and U12445 (N_12445,N_11874,N_11808);
xnor U12446 (N_12446,N_11387,N_11937);
nand U12447 (N_12447,N_11726,N_11556);
nand U12448 (N_12448,N_11978,N_11924);
or U12449 (N_12449,N_11985,N_11982);
and U12450 (N_12450,N_11629,N_11347);
xor U12451 (N_12451,N_11253,N_11379);
and U12452 (N_12452,N_11618,N_11716);
and U12453 (N_12453,N_11621,N_11803);
or U12454 (N_12454,N_11804,N_11878);
nand U12455 (N_12455,N_11491,N_11881);
nor U12456 (N_12456,N_11262,N_11737);
nor U12457 (N_12457,N_11212,N_11673);
and U12458 (N_12458,N_11877,N_11859);
or U12459 (N_12459,N_11691,N_11456);
nand U12460 (N_12460,N_11403,N_11831);
xnor U12461 (N_12461,N_11259,N_11808);
nor U12462 (N_12462,N_11871,N_11843);
or U12463 (N_12463,N_11979,N_11951);
nor U12464 (N_12464,N_11255,N_11940);
and U12465 (N_12465,N_11372,N_11409);
nor U12466 (N_12466,N_11507,N_11634);
nor U12467 (N_12467,N_11206,N_11380);
nor U12468 (N_12468,N_11662,N_11813);
or U12469 (N_12469,N_11949,N_11538);
or U12470 (N_12470,N_11496,N_11478);
xnor U12471 (N_12471,N_11238,N_11737);
nand U12472 (N_12472,N_11560,N_11380);
nand U12473 (N_12473,N_11894,N_11380);
or U12474 (N_12474,N_11481,N_11688);
and U12475 (N_12475,N_11957,N_11509);
nor U12476 (N_12476,N_11510,N_11389);
nor U12477 (N_12477,N_11946,N_11724);
nand U12478 (N_12478,N_11480,N_11487);
nand U12479 (N_12479,N_11761,N_11478);
and U12480 (N_12480,N_11703,N_11880);
nor U12481 (N_12481,N_11817,N_11293);
nor U12482 (N_12482,N_11209,N_11380);
or U12483 (N_12483,N_11600,N_11925);
nand U12484 (N_12484,N_11880,N_11241);
xor U12485 (N_12485,N_11767,N_11328);
nor U12486 (N_12486,N_11393,N_11751);
and U12487 (N_12487,N_11387,N_11229);
or U12488 (N_12488,N_11676,N_11862);
and U12489 (N_12489,N_11717,N_11404);
and U12490 (N_12490,N_11626,N_11989);
or U12491 (N_12491,N_11903,N_11337);
xor U12492 (N_12492,N_11916,N_11766);
nand U12493 (N_12493,N_11652,N_11346);
and U12494 (N_12494,N_11612,N_11726);
or U12495 (N_12495,N_11714,N_11773);
and U12496 (N_12496,N_11304,N_11240);
nand U12497 (N_12497,N_11968,N_11315);
nand U12498 (N_12498,N_11651,N_11383);
xnor U12499 (N_12499,N_11738,N_11705);
or U12500 (N_12500,N_11377,N_11489);
nand U12501 (N_12501,N_11265,N_11375);
xnor U12502 (N_12502,N_11961,N_11539);
or U12503 (N_12503,N_11988,N_11744);
nor U12504 (N_12504,N_11745,N_11940);
xor U12505 (N_12505,N_11779,N_11888);
nand U12506 (N_12506,N_11470,N_11788);
nor U12507 (N_12507,N_11350,N_11788);
nor U12508 (N_12508,N_11508,N_11800);
nor U12509 (N_12509,N_11637,N_11736);
and U12510 (N_12510,N_11957,N_11436);
xnor U12511 (N_12511,N_11284,N_11807);
and U12512 (N_12512,N_11261,N_11406);
nand U12513 (N_12513,N_11260,N_11649);
xor U12514 (N_12514,N_11953,N_11751);
nand U12515 (N_12515,N_11537,N_11479);
nor U12516 (N_12516,N_11605,N_11890);
nand U12517 (N_12517,N_11407,N_11928);
or U12518 (N_12518,N_11637,N_11445);
nand U12519 (N_12519,N_11254,N_11321);
or U12520 (N_12520,N_11734,N_11947);
nand U12521 (N_12521,N_11272,N_11505);
xor U12522 (N_12522,N_11541,N_11620);
or U12523 (N_12523,N_11237,N_11971);
nand U12524 (N_12524,N_11839,N_11971);
nor U12525 (N_12525,N_11823,N_11831);
nand U12526 (N_12526,N_11304,N_11846);
and U12527 (N_12527,N_11791,N_11940);
nand U12528 (N_12528,N_11944,N_11669);
and U12529 (N_12529,N_11227,N_11365);
or U12530 (N_12530,N_11751,N_11786);
or U12531 (N_12531,N_11950,N_11297);
nor U12532 (N_12532,N_11268,N_11262);
nand U12533 (N_12533,N_11605,N_11455);
nor U12534 (N_12534,N_11284,N_11334);
xor U12535 (N_12535,N_11240,N_11499);
xor U12536 (N_12536,N_11459,N_11475);
xnor U12537 (N_12537,N_11818,N_11771);
xnor U12538 (N_12538,N_11807,N_11569);
or U12539 (N_12539,N_11780,N_11326);
nand U12540 (N_12540,N_11483,N_11607);
nor U12541 (N_12541,N_11481,N_11924);
or U12542 (N_12542,N_11235,N_11718);
or U12543 (N_12543,N_11487,N_11908);
or U12544 (N_12544,N_11251,N_11844);
and U12545 (N_12545,N_11903,N_11831);
and U12546 (N_12546,N_11697,N_11234);
nor U12547 (N_12547,N_11513,N_11509);
and U12548 (N_12548,N_11309,N_11641);
xor U12549 (N_12549,N_11616,N_11942);
or U12550 (N_12550,N_11646,N_11677);
nor U12551 (N_12551,N_11704,N_11370);
xor U12552 (N_12552,N_11875,N_11354);
or U12553 (N_12553,N_11597,N_11336);
nor U12554 (N_12554,N_11675,N_11379);
xor U12555 (N_12555,N_11360,N_11385);
nor U12556 (N_12556,N_11611,N_11901);
nor U12557 (N_12557,N_11994,N_11202);
or U12558 (N_12558,N_11604,N_11380);
xnor U12559 (N_12559,N_11869,N_11502);
xor U12560 (N_12560,N_11760,N_11610);
nand U12561 (N_12561,N_11994,N_11557);
or U12562 (N_12562,N_11548,N_11938);
xor U12563 (N_12563,N_11334,N_11312);
nor U12564 (N_12564,N_11767,N_11987);
xor U12565 (N_12565,N_11838,N_11268);
or U12566 (N_12566,N_11755,N_11845);
nor U12567 (N_12567,N_11266,N_11369);
xnor U12568 (N_12568,N_11574,N_11495);
nand U12569 (N_12569,N_11955,N_11513);
nor U12570 (N_12570,N_11460,N_11473);
and U12571 (N_12571,N_11926,N_11367);
nor U12572 (N_12572,N_11733,N_11813);
nor U12573 (N_12573,N_11902,N_11258);
nand U12574 (N_12574,N_11677,N_11602);
and U12575 (N_12575,N_11437,N_11569);
or U12576 (N_12576,N_11682,N_11981);
nor U12577 (N_12577,N_11674,N_11798);
xor U12578 (N_12578,N_11961,N_11951);
nand U12579 (N_12579,N_11351,N_11709);
and U12580 (N_12580,N_11275,N_11521);
xnor U12581 (N_12581,N_11492,N_11502);
or U12582 (N_12582,N_11964,N_11617);
xnor U12583 (N_12583,N_11590,N_11893);
nor U12584 (N_12584,N_11379,N_11986);
nand U12585 (N_12585,N_11406,N_11909);
or U12586 (N_12586,N_11676,N_11236);
and U12587 (N_12587,N_11510,N_11644);
xor U12588 (N_12588,N_11620,N_11424);
or U12589 (N_12589,N_11314,N_11566);
and U12590 (N_12590,N_11395,N_11622);
nor U12591 (N_12591,N_11909,N_11850);
and U12592 (N_12592,N_11623,N_11993);
or U12593 (N_12593,N_11252,N_11983);
nand U12594 (N_12594,N_11376,N_11771);
xnor U12595 (N_12595,N_11943,N_11660);
xor U12596 (N_12596,N_11797,N_11538);
or U12597 (N_12597,N_11328,N_11995);
and U12598 (N_12598,N_11826,N_11344);
or U12599 (N_12599,N_11576,N_11265);
or U12600 (N_12600,N_11438,N_11772);
and U12601 (N_12601,N_11916,N_11902);
nand U12602 (N_12602,N_11265,N_11867);
and U12603 (N_12603,N_11970,N_11765);
nand U12604 (N_12604,N_11263,N_11221);
nand U12605 (N_12605,N_11803,N_11431);
or U12606 (N_12606,N_11624,N_11686);
xor U12607 (N_12607,N_11571,N_11226);
xnor U12608 (N_12608,N_11506,N_11519);
nand U12609 (N_12609,N_11993,N_11374);
xor U12610 (N_12610,N_11322,N_11937);
nor U12611 (N_12611,N_11603,N_11387);
and U12612 (N_12612,N_11579,N_11806);
nand U12613 (N_12613,N_11957,N_11479);
and U12614 (N_12614,N_11976,N_11863);
xnor U12615 (N_12615,N_11669,N_11217);
nor U12616 (N_12616,N_11596,N_11557);
or U12617 (N_12617,N_11404,N_11541);
and U12618 (N_12618,N_11469,N_11301);
or U12619 (N_12619,N_11266,N_11683);
or U12620 (N_12620,N_11326,N_11463);
or U12621 (N_12621,N_11885,N_11583);
and U12622 (N_12622,N_11240,N_11610);
or U12623 (N_12623,N_11696,N_11681);
xnor U12624 (N_12624,N_11868,N_11781);
nand U12625 (N_12625,N_11377,N_11319);
xnor U12626 (N_12626,N_11645,N_11472);
nand U12627 (N_12627,N_11476,N_11625);
xor U12628 (N_12628,N_11794,N_11580);
or U12629 (N_12629,N_11355,N_11803);
or U12630 (N_12630,N_11418,N_11806);
nor U12631 (N_12631,N_11498,N_11474);
nand U12632 (N_12632,N_11219,N_11368);
xnor U12633 (N_12633,N_11728,N_11513);
and U12634 (N_12634,N_11310,N_11907);
and U12635 (N_12635,N_11844,N_11869);
nand U12636 (N_12636,N_11285,N_11839);
nor U12637 (N_12637,N_11744,N_11424);
nor U12638 (N_12638,N_11290,N_11985);
xnor U12639 (N_12639,N_11765,N_11647);
xor U12640 (N_12640,N_11807,N_11766);
nor U12641 (N_12641,N_11730,N_11812);
nor U12642 (N_12642,N_11495,N_11504);
or U12643 (N_12643,N_11572,N_11658);
xnor U12644 (N_12644,N_11690,N_11213);
and U12645 (N_12645,N_11232,N_11235);
xor U12646 (N_12646,N_11624,N_11655);
nand U12647 (N_12647,N_11745,N_11207);
or U12648 (N_12648,N_11998,N_11697);
xor U12649 (N_12649,N_11972,N_11459);
and U12650 (N_12650,N_11202,N_11688);
or U12651 (N_12651,N_11631,N_11301);
and U12652 (N_12652,N_11932,N_11976);
xor U12653 (N_12653,N_11495,N_11761);
and U12654 (N_12654,N_11755,N_11350);
nor U12655 (N_12655,N_11589,N_11748);
or U12656 (N_12656,N_11249,N_11844);
or U12657 (N_12657,N_11890,N_11641);
and U12658 (N_12658,N_11847,N_11891);
nand U12659 (N_12659,N_11622,N_11886);
and U12660 (N_12660,N_11267,N_11791);
xor U12661 (N_12661,N_11371,N_11750);
and U12662 (N_12662,N_11214,N_11450);
and U12663 (N_12663,N_11334,N_11733);
nor U12664 (N_12664,N_11412,N_11678);
nor U12665 (N_12665,N_11594,N_11211);
nand U12666 (N_12666,N_11940,N_11871);
or U12667 (N_12667,N_11780,N_11654);
or U12668 (N_12668,N_11457,N_11475);
nor U12669 (N_12669,N_11900,N_11263);
xnor U12670 (N_12670,N_11577,N_11225);
or U12671 (N_12671,N_11415,N_11930);
xor U12672 (N_12672,N_11759,N_11838);
and U12673 (N_12673,N_11483,N_11875);
nand U12674 (N_12674,N_11418,N_11465);
xnor U12675 (N_12675,N_11408,N_11569);
and U12676 (N_12676,N_11503,N_11229);
nand U12677 (N_12677,N_11368,N_11642);
nor U12678 (N_12678,N_11487,N_11200);
or U12679 (N_12679,N_11866,N_11878);
or U12680 (N_12680,N_11579,N_11285);
nor U12681 (N_12681,N_11227,N_11688);
nor U12682 (N_12682,N_11730,N_11549);
or U12683 (N_12683,N_11317,N_11668);
xnor U12684 (N_12684,N_11685,N_11622);
nor U12685 (N_12685,N_11880,N_11261);
nand U12686 (N_12686,N_11967,N_11838);
and U12687 (N_12687,N_11344,N_11884);
xnor U12688 (N_12688,N_11595,N_11686);
nand U12689 (N_12689,N_11513,N_11420);
xnor U12690 (N_12690,N_11244,N_11341);
and U12691 (N_12691,N_11440,N_11690);
nor U12692 (N_12692,N_11575,N_11210);
nand U12693 (N_12693,N_11925,N_11881);
xnor U12694 (N_12694,N_11902,N_11869);
nor U12695 (N_12695,N_11910,N_11301);
xor U12696 (N_12696,N_11663,N_11200);
nor U12697 (N_12697,N_11848,N_11341);
nand U12698 (N_12698,N_11799,N_11319);
or U12699 (N_12699,N_11690,N_11640);
nor U12700 (N_12700,N_11435,N_11724);
or U12701 (N_12701,N_11737,N_11376);
nor U12702 (N_12702,N_11949,N_11704);
or U12703 (N_12703,N_11359,N_11464);
nor U12704 (N_12704,N_11858,N_11333);
nand U12705 (N_12705,N_11324,N_11912);
and U12706 (N_12706,N_11938,N_11475);
or U12707 (N_12707,N_11901,N_11875);
and U12708 (N_12708,N_11273,N_11405);
and U12709 (N_12709,N_11380,N_11734);
nand U12710 (N_12710,N_11757,N_11420);
xnor U12711 (N_12711,N_11473,N_11663);
and U12712 (N_12712,N_11737,N_11966);
nand U12713 (N_12713,N_11376,N_11832);
nor U12714 (N_12714,N_11568,N_11859);
and U12715 (N_12715,N_11702,N_11901);
xor U12716 (N_12716,N_11335,N_11388);
or U12717 (N_12717,N_11888,N_11575);
nor U12718 (N_12718,N_11607,N_11583);
nor U12719 (N_12719,N_11919,N_11636);
or U12720 (N_12720,N_11203,N_11482);
or U12721 (N_12721,N_11812,N_11943);
nand U12722 (N_12722,N_11656,N_11599);
nand U12723 (N_12723,N_11768,N_11711);
and U12724 (N_12724,N_11691,N_11558);
nor U12725 (N_12725,N_11284,N_11756);
xnor U12726 (N_12726,N_11439,N_11337);
nor U12727 (N_12727,N_11251,N_11653);
nor U12728 (N_12728,N_11604,N_11660);
nand U12729 (N_12729,N_11462,N_11716);
and U12730 (N_12730,N_11372,N_11483);
or U12731 (N_12731,N_11943,N_11729);
nand U12732 (N_12732,N_11609,N_11625);
nand U12733 (N_12733,N_11409,N_11290);
or U12734 (N_12734,N_11221,N_11838);
xor U12735 (N_12735,N_11244,N_11330);
xor U12736 (N_12736,N_11644,N_11654);
or U12737 (N_12737,N_11739,N_11642);
nand U12738 (N_12738,N_11925,N_11510);
xor U12739 (N_12739,N_11748,N_11829);
and U12740 (N_12740,N_11421,N_11547);
or U12741 (N_12741,N_11745,N_11484);
and U12742 (N_12742,N_11612,N_11678);
nand U12743 (N_12743,N_11305,N_11561);
and U12744 (N_12744,N_11641,N_11683);
and U12745 (N_12745,N_11898,N_11274);
and U12746 (N_12746,N_11991,N_11832);
or U12747 (N_12747,N_11560,N_11661);
xnor U12748 (N_12748,N_11323,N_11768);
nor U12749 (N_12749,N_11593,N_11403);
or U12750 (N_12750,N_11752,N_11401);
or U12751 (N_12751,N_11641,N_11478);
xor U12752 (N_12752,N_11574,N_11490);
nor U12753 (N_12753,N_11869,N_11953);
xor U12754 (N_12754,N_11518,N_11945);
xor U12755 (N_12755,N_11481,N_11941);
and U12756 (N_12756,N_11660,N_11987);
and U12757 (N_12757,N_11853,N_11612);
and U12758 (N_12758,N_11286,N_11890);
nand U12759 (N_12759,N_11453,N_11683);
xor U12760 (N_12760,N_11898,N_11903);
nand U12761 (N_12761,N_11643,N_11825);
nand U12762 (N_12762,N_11328,N_11354);
xor U12763 (N_12763,N_11895,N_11857);
xor U12764 (N_12764,N_11737,N_11792);
nand U12765 (N_12765,N_11845,N_11745);
or U12766 (N_12766,N_11231,N_11714);
xor U12767 (N_12767,N_11557,N_11995);
xnor U12768 (N_12768,N_11494,N_11599);
xor U12769 (N_12769,N_11342,N_11740);
and U12770 (N_12770,N_11650,N_11448);
and U12771 (N_12771,N_11600,N_11446);
nand U12772 (N_12772,N_11852,N_11685);
nor U12773 (N_12773,N_11627,N_11217);
and U12774 (N_12774,N_11644,N_11448);
xor U12775 (N_12775,N_11620,N_11913);
xor U12776 (N_12776,N_11812,N_11507);
or U12777 (N_12777,N_11974,N_11556);
xnor U12778 (N_12778,N_11936,N_11274);
nand U12779 (N_12779,N_11663,N_11890);
xnor U12780 (N_12780,N_11693,N_11845);
or U12781 (N_12781,N_11347,N_11345);
nand U12782 (N_12782,N_11467,N_11880);
nor U12783 (N_12783,N_11418,N_11776);
nand U12784 (N_12784,N_11868,N_11879);
or U12785 (N_12785,N_11343,N_11317);
or U12786 (N_12786,N_11970,N_11640);
and U12787 (N_12787,N_11321,N_11593);
and U12788 (N_12788,N_11517,N_11581);
nor U12789 (N_12789,N_11746,N_11530);
or U12790 (N_12790,N_11659,N_11405);
or U12791 (N_12791,N_11435,N_11220);
xnor U12792 (N_12792,N_11845,N_11522);
xor U12793 (N_12793,N_11953,N_11569);
or U12794 (N_12794,N_11790,N_11327);
xnor U12795 (N_12795,N_11310,N_11557);
or U12796 (N_12796,N_11579,N_11670);
nand U12797 (N_12797,N_11427,N_11881);
nand U12798 (N_12798,N_11361,N_11696);
and U12799 (N_12799,N_11939,N_11576);
and U12800 (N_12800,N_12473,N_12307);
xor U12801 (N_12801,N_12434,N_12276);
nor U12802 (N_12802,N_12526,N_12103);
nand U12803 (N_12803,N_12183,N_12179);
nor U12804 (N_12804,N_12743,N_12447);
nand U12805 (N_12805,N_12204,N_12602);
or U12806 (N_12806,N_12421,N_12363);
and U12807 (N_12807,N_12060,N_12286);
and U12808 (N_12808,N_12778,N_12340);
xor U12809 (N_12809,N_12016,N_12043);
or U12810 (N_12810,N_12501,N_12796);
and U12811 (N_12811,N_12719,N_12351);
nand U12812 (N_12812,N_12359,N_12372);
or U12813 (N_12813,N_12677,N_12456);
xnor U12814 (N_12814,N_12328,N_12226);
or U12815 (N_12815,N_12138,N_12534);
and U12816 (N_12816,N_12504,N_12232);
nand U12817 (N_12817,N_12026,N_12066);
nand U12818 (N_12818,N_12166,N_12368);
and U12819 (N_12819,N_12735,N_12281);
nand U12820 (N_12820,N_12107,N_12694);
and U12821 (N_12821,N_12762,N_12393);
or U12822 (N_12822,N_12094,N_12667);
nand U12823 (N_12823,N_12300,N_12295);
xor U12824 (N_12824,N_12680,N_12317);
xnor U12825 (N_12825,N_12203,N_12745);
xnor U12826 (N_12826,N_12779,N_12112);
nand U12827 (N_12827,N_12303,N_12180);
or U12828 (N_12828,N_12387,N_12342);
nor U12829 (N_12829,N_12047,N_12427);
or U12830 (N_12830,N_12323,N_12588);
and U12831 (N_12831,N_12057,N_12210);
xor U12832 (N_12832,N_12321,N_12253);
nor U12833 (N_12833,N_12123,N_12111);
nor U12834 (N_12834,N_12242,N_12348);
or U12835 (N_12835,N_12108,N_12480);
nand U12836 (N_12836,N_12669,N_12791);
nor U12837 (N_12837,N_12464,N_12632);
or U12838 (N_12838,N_12320,N_12326);
or U12839 (N_12839,N_12079,N_12714);
or U12840 (N_12840,N_12312,N_12246);
and U12841 (N_12841,N_12515,N_12338);
xnor U12842 (N_12842,N_12064,N_12491);
and U12843 (N_12843,N_12214,N_12760);
nor U12844 (N_12844,N_12751,N_12020);
or U12845 (N_12845,N_12655,N_12593);
or U12846 (N_12846,N_12578,N_12285);
nand U12847 (N_12847,N_12229,N_12185);
and U12848 (N_12848,N_12598,N_12708);
nor U12849 (N_12849,N_12182,N_12054);
and U12850 (N_12850,N_12622,N_12362);
xor U12851 (N_12851,N_12579,N_12380);
nand U12852 (N_12852,N_12699,N_12412);
and U12853 (N_12853,N_12014,N_12547);
or U12854 (N_12854,N_12440,N_12799);
and U12855 (N_12855,N_12413,N_12153);
nand U12856 (N_12856,N_12116,N_12687);
or U12857 (N_12857,N_12083,N_12013);
nand U12858 (N_12858,N_12592,N_12557);
nor U12859 (N_12859,N_12068,N_12136);
nand U12860 (N_12860,N_12336,N_12065);
nor U12861 (N_12861,N_12788,N_12268);
xnor U12862 (N_12862,N_12710,N_12439);
or U12863 (N_12863,N_12221,N_12192);
xor U12864 (N_12864,N_12178,N_12304);
xor U12865 (N_12865,N_12048,N_12584);
or U12866 (N_12866,N_12776,N_12543);
nor U12867 (N_12867,N_12332,N_12702);
nand U12868 (N_12868,N_12305,N_12518);
nand U12869 (N_12869,N_12442,N_12104);
nand U12870 (N_12870,N_12205,N_12199);
nand U12871 (N_12871,N_12759,N_12154);
nand U12872 (N_12872,N_12683,N_12436);
and U12873 (N_12873,N_12503,N_12318);
nand U12874 (N_12874,N_12748,N_12451);
and U12875 (N_12875,N_12089,N_12511);
or U12876 (N_12876,N_12084,N_12675);
xor U12877 (N_12877,N_12597,N_12209);
nor U12878 (N_12878,N_12656,N_12635);
nand U12879 (N_12879,N_12376,N_12438);
nand U12880 (N_12880,N_12015,N_12149);
nor U12881 (N_12881,N_12409,N_12659);
xnor U12882 (N_12882,N_12789,N_12604);
or U12883 (N_12883,N_12525,N_12755);
xnor U12884 (N_12884,N_12522,N_12494);
nor U12885 (N_12885,N_12040,N_12255);
nand U12886 (N_12886,N_12408,N_12781);
xor U12887 (N_12887,N_12704,N_12074);
nand U12888 (N_12888,N_12093,N_12249);
or U12889 (N_12889,N_12512,N_12402);
and U12890 (N_12890,N_12572,N_12390);
and U12891 (N_12891,N_12453,N_12388);
nand U12892 (N_12892,N_12010,N_12155);
and U12893 (N_12893,N_12398,N_12533);
and U12894 (N_12894,N_12437,N_12175);
and U12895 (N_12895,N_12186,N_12033);
and U12896 (N_12896,N_12037,N_12661);
xnor U12897 (N_12897,N_12580,N_12654);
nor U12898 (N_12898,N_12097,N_12234);
nor U12899 (N_12899,N_12308,N_12457);
nor U12900 (N_12900,N_12141,N_12469);
nor U12901 (N_12901,N_12044,N_12200);
xor U12902 (N_12902,N_12615,N_12206);
nand U12903 (N_12903,N_12552,N_12029);
and U12904 (N_12904,N_12299,N_12628);
or U12905 (N_12905,N_12637,N_12264);
nand U12906 (N_12906,N_12091,N_12092);
xor U12907 (N_12907,N_12128,N_12244);
or U12908 (N_12908,N_12401,N_12273);
nand U12909 (N_12909,N_12489,N_12617);
nor U12910 (N_12910,N_12441,N_12536);
and U12911 (N_12911,N_12275,N_12395);
or U12912 (N_12912,N_12056,N_12310);
xnor U12913 (N_12913,N_12577,N_12196);
or U12914 (N_12914,N_12734,N_12647);
or U12915 (N_12915,N_12757,N_12357);
xor U12916 (N_12916,N_12478,N_12425);
nor U12917 (N_12917,N_12158,N_12718);
and U12918 (N_12918,N_12375,N_12430);
xor U12919 (N_12919,N_12007,N_12365);
xor U12920 (N_12920,N_12233,N_12608);
nor U12921 (N_12921,N_12260,N_12293);
xor U12922 (N_12922,N_12361,N_12679);
xor U12923 (N_12923,N_12201,N_12638);
nand U12924 (N_12924,N_12493,N_12674);
nor U12925 (N_12925,N_12207,N_12258);
or U12926 (N_12926,N_12100,N_12383);
and U12927 (N_12927,N_12370,N_12730);
or U12928 (N_12928,N_12485,N_12591);
xnor U12929 (N_12929,N_12018,N_12227);
nor U12930 (N_12930,N_12055,N_12171);
nor U12931 (N_12931,N_12551,N_12521);
nand U12932 (N_12932,N_12746,N_12549);
or U12933 (N_12933,N_12771,N_12753);
nand U12934 (N_12934,N_12049,N_12486);
and U12935 (N_12935,N_12392,N_12382);
nand U12936 (N_12936,N_12193,N_12184);
xnor U12937 (N_12937,N_12125,N_12477);
xor U12938 (N_12938,N_12252,N_12793);
and U12939 (N_12939,N_12137,N_12174);
nor U12940 (N_12940,N_12432,N_12532);
nor U12941 (N_12941,N_12053,N_12524);
and U12942 (N_12942,N_12262,N_12768);
or U12943 (N_12943,N_12554,N_12523);
and U12944 (N_12944,N_12645,N_12662);
nor U12945 (N_12945,N_12220,N_12565);
nor U12946 (N_12946,N_12405,N_12767);
or U12947 (N_12947,N_12646,N_12649);
xor U12948 (N_12948,N_12298,N_12225);
and U12949 (N_12949,N_12017,N_12752);
or U12950 (N_12950,N_12177,N_12140);
or U12951 (N_12951,N_12292,N_12240);
and U12952 (N_12952,N_12777,N_12082);
nor U12953 (N_12953,N_12720,N_12563);
or U12954 (N_12954,N_12119,N_12665);
nand U12955 (N_12955,N_12217,N_12463);
nor U12956 (N_12956,N_12198,N_12411);
nor U12957 (N_12957,N_12620,N_12231);
nand U12958 (N_12958,N_12098,N_12230);
nand U12959 (N_12959,N_12465,N_12250);
xor U12960 (N_12960,N_12725,N_12676);
or U12961 (N_12961,N_12459,N_12556);
nor U12962 (N_12962,N_12423,N_12626);
nor U12963 (N_12963,N_12723,N_12036);
xnor U12964 (N_12964,N_12245,N_12187);
xor U12965 (N_12965,N_12352,N_12701);
nand U12966 (N_12966,N_12132,N_12527);
nor U12967 (N_12967,N_12564,N_12021);
nor U12968 (N_12968,N_12085,N_12031);
nor U12969 (N_12969,N_12668,N_12163);
nor U12970 (N_12970,N_12347,N_12650);
nand U12971 (N_12971,N_12594,N_12756);
and U12972 (N_12972,N_12311,N_12228);
or U12973 (N_12973,N_12490,N_12173);
and U12974 (N_12974,N_12416,N_12507);
or U12975 (N_12975,N_12775,N_12455);
xor U12976 (N_12976,N_12574,N_12386);
or U12977 (N_12977,N_12280,N_12337);
xor U12978 (N_12978,N_12052,N_12707);
nor U12979 (N_12979,N_12785,N_12329);
xnor U12980 (N_12980,N_12619,N_12706);
or U12981 (N_12981,N_12681,N_12474);
and U12982 (N_12982,N_12333,N_12600);
or U12983 (N_12983,N_12302,N_12695);
and U12984 (N_12984,N_12639,N_12058);
and U12985 (N_12985,N_12691,N_12120);
nor U12986 (N_12986,N_12195,N_12061);
nor U12987 (N_12987,N_12324,N_12479);
and U12988 (N_12988,N_12063,N_12703);
nand U12989 (N_12989,N_12030,N_12548);
and U12990 (N_12990,N_12167,N_12261);
nor U12991 (N_12991,N_12599,N_12028);
nand U12992 (N_12992,N_12164,N_12389);
and U12993 (N_12993,N_12350,N_12290);
and U12994 (N_12994,N_12287,N_12127);
and U12995 (N_12995,N_12378,N_12259);
nand U12996 (N_12996,N_12143,N_12651);
nor U12997 (N_12997,N_12722,N_12513);
nor U12998 (N_12998,N_12219,N_12309);
nor U12999 (N_12999,N_12297,N_12355);
and U13000 (N_13000,N_12101,N_12783);
xor U13001 (N_13001,N_12222,N_12535);
nand U13002 (N_13002,N_12254,N_12315);
nor U13003 (N_13003,N_12571,N_12476);
or U13004 (N_13004,N_12733,N_12467);
nand U13005 (N_13005,N_12160,N_12062);
nand U13006 (N_13006,N_12142,N_12197);
or U13007 (N_13007,N_12553,N_12462);
nand U13008 (N_13008,N_12582,N_12397);
nand U13009 (N_13009,N_12696,N_12454);
xor U13010 (N_13010,N_12624,N_12514);
xnor U13011 (N_13011,N_12537,N_12585);
and U13012 (N_13012,N_12096,N_12658);
and U13013 (N_13013,N_12000,N_12327);
or U13014 (N_13014,N_12575,N_12446);
and U13015 (N_13015,N_12090,N_12247);
xor U13016 (N_13016,N_12278,N_12224);
and U13017 (N_13017,N_12152,N_12769);
xor U13018 (N_13018,N_12277,N_12288);
nor U13019 (N_13019,N_12106,N_12406);
nand U13020 (N_13020,N_12157,N_12099);
nand U13021 (N_13021,N_12148,N_12741);
xnor U13022 (N_13022,N_12761,N_12188);
and U13023 (N_13023,N_12773,N_12241);
xor U13024 (N_13024,N_12528,N_12698);
nor U13025 (N_13025,N_12122,N_12519);
nand U13026 (N_13026,N_12283,N_12110);
nand U13027 (N_13027,N_12322,N_12483);
xnor U13028 (N_13028,N_12077,N_12400);
and U13029 (N_13029,N_12343,N_12069);
and U13030 (N_13030,N_12130,N_12611);
xnor U13031 (N_13031,N_12381,N_12417);
nand U13032 (N_13032,N_12024,N_12023);
nand U13033 (N_13033,N_12566,N_12294);
xnor U13034 (N_13034,N_12335,N_12448);
or U13035 (N_13035,N_12095,N_12027);
and U13036 (N_13036,N_12129,N_12118);
and U13037 (N_13037,N_12570,N_12139);
and U13038 (N_13038,N_12341,N_12510);
or U13039 (N_13039,N_12728,N_12282);
nor U13040 (N_13040,N_12629,N_12078);
and U13041 (N_13041,N_12742,N_12444);
nor U13042 (N_13042,N_12251,N_12606);
nand U13043 (N_13043,N_12727,N_12265);
xnor U13044 (N_13044,N_12612,N_12487);
and U13045 (N_13045,N_12272,N_12731);
and U13046 (N_13046,N_12555,N_12428);
and U13047 (N_13047,N_12765,N_12750);
or U13048 (N_13048,N_12325,N_12663);
nand U13049 (N_13049,N_12419,N_12542);
and U13050 (N_13050,N_12189,N_12072);
or U13051 (N_13051,N_12770,N_12424);
nand U13052 (N_13052,N_12156,N_12685);
or U13053 (N_13053,N_12377,N_12460);
and U13054 (N_13054,N_12481,N_12729);
nand U13055 (N_13055,N_12509,N_12739);
and U13056 (N_13056,N_12712,N_12236);
nor U13057 (N_13057,N_12059,N_12697);
or U13058 (N_13058,N_12505,N_12529);
nand U13059 (N_13059,N_12172,N_12468);
xnor U13060 (N_13060,N_12114,N_12051);
nand U13061 (N_13061,N_12373,N_12634);
nor U13062 (N_13062,N_12794,N_12216);
and U13063 (N_13063,N_12354,N_12589);
nand U13064 (N_13064,N_12609,N_12466);
nor U13065 (N_13065,N_12786,N_12168);
xor U13066 (N_13066,N_12191,N_12176);
nor U13067 (N_13067,N_12420,N_12145);
xnor U13068 (N_13068,N_12330,N_12569);
nand U13069 (N_13069,N_12603,N_12670);
xor U13070 (N_13070,N_12688,N_12508);
xnor U13071 (N_13071,N_12223,N_12539);
xor U13072 (N_13072,N_12218,N_12492);
and U13073 (N_13073,N_12117,N_12445);
or U13074 (N_13074,N_12429,N_12008);
and U13075 (N_13075,N_12339,N_12657);
or U13076 (N_13076,N_12541,N_12644);
nand U13077 (N_13077,N_12652,N_12763);
nor U13078 (N_13078,N_12019,N_12738);
and U13079 (N_13079,N_12671,N_12484);
nor U13080 (N_13080,N_12621,N_12009);
and U13081 (N_13081,N_12418,N_12345);
and U13082 (N_13082,N_12431,N_12291);
or U13083 (N_13083,N_12165,N_12653);
nor U13084 (N_13084,N_12666,N_12296);
nand U13085 (N_13085,N_12784,N_12081);
nand U13086 (N_13086,N_12737,N_12006);
nor U13087 (N_13087,N_12035,N_12792);
or U13088 (N_13088,N_12237,N_12627);
nor U13089 (N_13089,N_12371,N_12147);
xor U13090 (N_13090,N_12146,N_12516);
xor U13091 (N_13091,N_12071,N_12497);
xor U13092 (N_13092,N_12686,N_12313);
xnor U13093 (N_13093,N_12590,N_12011);
and U13094 (N_13094,N_12374,N_12538);
or U13095 (N_13095,N_12520,N_12289);
xor U13096 (N_13096,N_12369,N_12349);
xor U13097 (N_13097,N_12475,N_12159);
and U13098 (N_13098,N_12780,N_12001);
nor U13099 (N_13099,N_12126,N_12134);
nand U13100 (N_13100,N_12102,N_12530);
nand U13101 (N_13101,N_12625,N_12266);
nand U13102 (N_13102,N_12208,N_12076);
nand U13103 (N_13103,N_12144,N_12631);
xor U13104 (N_13104,N_12170,N_12782);
and U13105 (N_13105,N_12070,N_12150);
xor U13106 (N_13106,N_12744,N_12169);
or U13107 (N_13107,N_12726,N_12559);
nand U13108 (N_13108,N_12435,N_12581);
or U13109 (N_13109,N_12614,N_12573);
nor U13110 (N_13110,N_12787,N_12716);
nor U13111 (N_13111,N_12568,N_12038);
xnor U13112 (N_13112,N_12798,N_12640);
xnor U13113 (N_13113,N_12472,N_12391);
nor U13114 (N_13114,N_12396,N_12238);
xor U13115 (N_13115,N_12764,N_12692);
nand U13116 (N_13116,N_12364,N_12039);
nor U13117 (N_13117,N_12732,N_12041);
nor U13118 (N_13118,N_12181,N_12190);
xor U13119 (N_13119,N_12660,N_12358);
or U13120 (N_13120,N_12724,N_12133);
xor U13121 (N_13121,N_12747,N_12613);
and U13122 (N_13122,N_12766,N_12705);
nor U13123 (N_13123,N_12002,N_12558);
and U13124 (N_13124,N_12689,N_12506);
xnor U13125 (N_13125,N_12003,N_12601);
xor U13126 (N_13126,N_12105,N_12540);
or U13127 (N_13127,N_12618,N_12546);
and U13128 (N_13128,N_12749,N_12673);
or U13129 (N_13129,N_12215,N_12005);
or U13130 (N_13130,N_12496,N_12693);
nand U13131 (N_13131,N_12790,N_12162);
or U13132 (N_13132,N_12360,N_12797);
nor U13133 (N_13133,N_12595,N_12113);
nor U13134 (N_13134,N_12279,N_12004);
xnor U13135 (N_13135,N_12353,N_12334);
or U13136 (N_13136,N_12124,N_12471);
or U13137 (N_13137,N_12517,N_12499);
nor U13138 (N_13138,N_12239,N_12795);
nand U13139 (N_13139,N_12306,N_12356);
or U13140 (N_13140,N_12717,N_12086);
and U13141 (N_13141,N_12022,N_12678);
or U13142 (N_13142,N_12045,N_12422);
nand U13143 (N_13143,N_12560,N_12032);
xor U13144 (N_13144,N_12256,N_12407);
and U13145 (N_13145,N_12450,N_12012);
and U13146 (N_13146,N_12270,N_12586);
and U13147 (N_13147,N_12034,N_12088);
xnor U13148 (N_13148,N_12690,N_12495);
or U13149 (N_13149,N_12274,N_12684);
and U13150 (N_13150,N_12443,N_12587);
nand U13151 (N_13151,N_12050,N_12319);
xnor U13152 (N_13152,N_12080,N_12458);
nor U13153 (N_13153,N_12774,N_12500);
nand U13154 (N_13154,N_12067,N_12046);
xor U13155 (N_13155,N_12550,N_12583);
nand U13156 (N_13156,N_12452,N_12561);
nor U13157 (N_13157,N_12721,N_12284);
xnor U13158 (N_13158,N_12202,N_12610);
and U13159 (N_13159,N_12161,N_12502);
or U13160 (N_13160,N_12344,N_12404);
or U13161 (N_13161,N_12562,N_12121);
or U13162 (N_13162,N_12544,N_12498);
and U13163 (N_13163,N_12042,N_12385);
nor U13164 (N_13164,N_12384,N_12664);
nor U13165 (N_13165,N_12025,N_12367);
nor U13166 (N_13166,N_12648,N_12772);
nand U13167 (N_13167,N_12087,N_12403);
and U13168 (N_13168,N_12672,N_12331);
nor U13169 (N_13169,N_12641,N_12643);
or U13170 (N_13170,N_12596,N_12109);
xnor U13171 (N_13171,N_12482,N_12700);
or U13172 (N_13172,N_12567,N_12607);
nand U13173 (N_13173,N_12616,N_12713);
xor U13174 (N_13174,N_12316,N_12715);
nand U13175 (N_13175,N_12426,N_12488);
xor U13176 (N_13176,N_12151,N_12257);
nand U13177 (N_13177,N_12709,N_12605);
xor U13178 (N_13178,N_12682,N_12531);
nand U13179 (N_13179,N_12346,N_12379);
nor U13180 (N_13180,N_12075,N_12248);
xnor U13181 (N_13181,N_12213,N_12433);
xnor U13182 (N_13182,N_12135,N_12711);
nor U13183 (N_13183,N_12267,N_12211);
nor U13184 (N_13184,N_12269,N_12399);
nand U13185 (N_13185,N_12263,N_12194);
xnor U13186 (N_13186,N_12576,N_12271);
or U13187 (N_13187,N_12131,N_12470);
or U13188 (N_13188,N_12758,N_12754);
xnor U13189 (N_13189,N_12410,N_12449);
nor U13190 (N_13190,N_12461,N_12243);
xnor U13191 (N_13191,N_12073,N_12623);
nor U13192 (N_13192,N_12301,N_12366);
or U13193 (N_13193,N_12235,N_12642);
nand U13194 (N_13194,N_12636,N_12740);
nand U13195 (N_13195,N_12630,N_12736);
nor U13196 (N_13196,N_12115,N_12314);
nand U13197 (N_13197,N_12633,N_12414);
and U13198 (N_13198,N_12415,N_12394);
and U13199 (N_13199,N_12212,N_12545);
or U13200 (N_13200,N_12002,N_12062);
or U13201 (N_13201,N_12192,N_12718);
xor U13202 (N_13202,N_12317,N_12645);
nor U13203 (N_13203,N_12363,N_12440);
nor U13204 (N_13204,N_12361,N_12709);
xnor U13205 (N_13205,N_12674,N_12189);
xnor U13206 (N_13206,N_12789,N_12477);
or U13207 (N_13207,N_12053,N_12761);
and U13208 (N_13208,N_12533,N_12059);
or U13209 (N_13209,N_12088,N_12668);
and U13210 (N_13210,N_12470,N_12673);
xor U13211 (N_13211,N_12390,N_12450);
and U13212 (N_13212,N_12063,N_12164);
nor U13213 (N_13213,N_12346,N_12334);
or U13214 (N_13214,N_12791,N_12402);
nand U13215 (N_13215,N_12746,N_12574);
xnor U13216 (N_13216,N_12407,N_12682);
and U13217 (N_13217,N_12133,N_12094);
nand U13218 (N_13218,N_12438,N_12531);
and U13219 (N_13219,N_12170,N_12155);
xnor U13220 (N_13220,N_12733,N_12648);
xnor U13221 (N_13221,N_12088,N_12084);
or U13222 (N_13222,N_12511,N_12069);
xnor U13223 (N_13223,N_12072,N_12279);
and U13224 (N_13224,N_12679,N_12715);
nand U13225 (N_13225,N_12513,N_12666);
nor U13226 (N_13226,N_12178,N_12149);
nor U13227 (N_13227,N_12702,N_12581);
nor U13228 (N_13228,N_12527,N_12598);
nor U13229 (N_13229,N_12498,N_12637);
and U13230 (N_13230,N_12001,N_12235);
or U13231 (N_13231,N_12121,N_12585);
nand U13232 (N_13232,N_12576,N_12086);
nand U13233 (N_13233,N_12355,N_12740);
or U13234 (N_13234,N_12122,N_12241);
or U13235 (N_13235,N_12575,N_12643);
nor U13236 (N_13236,N_12607,N_12110);
or U13237 (N_13237,N_12131,N_12556);
xnor U13238 (N_13238,N_12221,N_12677);
or U13239 (N_13239,N_12399,N_12464);
nand U13240 (N_13240,N_12236,N_12340);
nor U13241 (N_13241,N_12625,N_12050);
xor U13242 (N_13242,N_12239,N_12211);
xnor U13243 (N_13243,N_12116,N_12361);
nor U13244 (N_13244,N_12544,N_12647);
xor U13245 (N_13245,N_12241,N_12205);
xnor U13246 (N_13246,N_12361,N_12103);
nand U13247 (N_13247,N_12569,N_12219);
and U13248 (N_13248,N_12093,N_12003);
nand U13249 (N_13249,N_12484,N_12103);
nor U13250 (N_13250,N_12698,N_12462);
xnor U13251 (N_13251,N_12794,N_12669);
and U13252 (N_13252,N_12522,N_12223);
nor U13253 (N_13253,N_12774,N_12347);
or U13254 (N_13254,N_12034,N_12120);
and U13255 (N_13255,N_12351,N_12238);
and U13256 (N_13256,N_12602,N_12108);
or U13257 (N_13257,N_12110,N_12729);
or U13258 (N_13258,N_12017,N_12562);
and U13259 (N_13259,N_12142,N_12075);
and U13260 (N_13260,N_12272,N_12205);
xnor U13261 (N_13261,N_12592,N_12056);
and U13262 (N_13262,N_12671,N_12002);
nand U13263 (N_13263,N_12684,N_12601);
and U13264 (N_13264,N_12142,N_12192);
or U13265 (N_13265,N_12382,N_12312);
or U13266 (N_13266,N_12532,N_12158);
or U13267 (N_13267,N_12643,N_12408);
or U13268 (N_13268,N_12412,N_12773);
nand U13269 (N_13269,N_12374,N_12196);
xor U13270 (N_13270,N_12577,N_12614);
xnor U13271 (N_13271,N_12283,N_12490);
nor U13272 (N_13272,N_12127,N_12569);
nand U13273 (N_13273,N_12036,N_12179);
or U13274 (N_13274,N_12755,N_12372);
or U13275 (N_13275,N_12713,N_12046);
nor U13276 (N_13276,N_12603,N_12083);
or U13277 (N_13277,N_12208,N_12359);
and U13278 (N_13278,N_12140,N_12585);
nand U13279 (N_13279,N_12755,N_12748);
and U13280 (N_13280,N_12786,N_12631);
xnor U13281 (N_13281,N_12297,N_12198);
nand U13282 (N_13282,N_12467,N_12168);
nand U13283 (N_13283,N_12226,N_12153);
and U13284 (N_13284,N_12179,N_12322);
xnor U13285 (N_13285,N_12339,N_12515);
and U13286 (N_13286,N_12504,N_12771);
xor U13287 (N_13287,N_12357,N_12465);
nand U13288 (N_13288,N_12331,N_12218);
nand U13289 (N_13289,N_12715,N_12002);
xnor U13290 (N_13290,N_12044,N_12421);
nand U13291 (N_13291,N_12339,N_12567);
and U13292 (N_13292,N_12208,N_12064);
xor U13293 (N_13293,N_12030,N_12697);
nand U13294 (N_13294,N_12226,N_12437);
and U13295 (N_13295,N_12772,N_12466);
xnor U13296 (N_13296,N_12089,N_12120);
nor U13297 (N_13297,N_12092,N_12680);
xor U13298 (N_13298,N_12125,N_12025);
or U13299 (N_13299,N_12264,N_12621);
nor U13300 (N_13300,N_12433,N_12604);
xor U13301 (N_13301,N_12562,N_12186);
or U13302 (N_13302,N_12538,N_12744);
and U13303 (N_13303,N_12756,N_12672);
or U13304 (N_13304,N_12091,N_12738);
and U13305 (N_13305,N_12084,N_12510);
xnor U13306 (N_13306,N_12268,N_12093);
xnor U13307 (N_13307,N_12299,N_12304);
xor U13308 (N_13308,N_12062,N_12672);
nor U13309 (N_13309,N_12068,N_12242);
nor U13310 (N_13310,N_12718,N_12062);
or U13311 (N_13311,N_12361,N_12556);
or U13312 (N_13312,N_12202,N_12461);
nor U13313 (N_13313,N_12365,N_12164);
and U13314 (N_13314,N_12457,N_12215);
nand U13315 (N_13315,N_12399,N_12450);
nor U13316 (N_13316,N_12523,N_12753);
nand U13317 (N_13317,N_12357,N_12510);
and U13318 (N_13318,N_12675,N_12746);
xor U13319 (N_13319,N_12156,N_12469);
and U13320 (N_13320,N_12388,N_12117);
or U13321 (N_13321,N_12187,N_12578);
or U13322 (N_13322,N_12329,N_12246);
nand U13323 (N_13323,N_12120,N_12160);
and U13324 (N_13324,N_12203,N_12351);
nor U13325 (N_13325,N_12090,N_12060);
xnor U13326 (N_13326,N_12789,N_12687);
and U13327 (N_13327,N_12692,N_12309);
nand U13328 (N_13328,N_12279,N_12564);
nand U13329 (N_13329,N_12775,N_12447);
and U13330 (N_13330,N_12538,N_12363);
nor U13331 (N_13331,N_12501,N_12587);
nor U13332 (N_13332,N_12018,N_12702);
nor U13333 (N_13333,N_12774,N_12272);
and U13334 (N_13334,N_12384,N_12435);
and U13335 (N_13335,N_12570,N_12372);
nand U13336 (N_13336,N_12497,N_12171);
or U13337 (N_13337,N_12588,N_12115);
nand U13338 (N_13338,N_12508,N_12156);
nand U13339 (N_13339,N_12375,N_12709);
nand U13340 (N_13340,N_12399,N_12703);
nor U13341 (N_13341,N_12699,N_12315);
or U13342 (N_13342,N_12158,N_12001);
and U13343 (N_13343,N_12759,N_12677);
xnor U13344 (N_13344,N_12113,N_12121);
and U13345 (N_13345,N_12135,N_12592);
nor U13346 (N_13346,N_12797,N_12606);
and U13347 (N_13347,N_12146,N_12439);
xnor U13348 (N_13348,N_12604,N_12439);
nor U13349 (N_13349,N_12428,N_12519);
xnor U13350 (N_13350,N_12518,N_12629);
nor U13351 (N_13351,N_12627,N_12208);
and U13352 (N_13352,N_12341,N_12732);
and U13353 (N_13353,N_12287,N_12422);
nor U13354 (N_13354,N_12524,N_12495);
nand U13355 (N_13355,N_12558,N_12149);
and U13356 (N_13356,N_12662,N_12305);
nand U13357 (N_13357,N_12464,N_12345);
nor U13358 (N_13358,N_12687,N_12422);
nor U13359 (N_13359,N_12270,N_12205);
xnor U13360 (N_13360,N_12097,N_12608);
xnor U13361 (N_13361,N_12393,N_12292);
xor U13362 (N_13362,N_12630,N_12100);
nand U13363 (N_13363,N_12503,N_12099);
nor U13364 (N_13364,N_12710,N_12784);
nand U13365 (N_13365,N_12102,N_12628);
and U13366 (N_13366,N_12547,N_12325);
xor U13367 (N_13367,N_12467,N_12770);
nor U13368 (N_13368,N_12379,N_12262);
nor U13369 (N_13369,N_12694,N_12020);
nor U13370 (N_13370,N_12577,N_12367);
nor U13371 (N_13371,N_12037,N_12340);
and U13372 (N_13372,N_12192,N_12535);
nand U13373 (N_13373,N_12190,N_12623);
nor U13374 (N_13374,N_12448,N_12469);
or U13375 (N_13375,N_12580,N_12505);
xor U13376 (N_13376,N_12324,N_12613);
xor U13377 (N_13377,N_12074,N_12541);
xnor U13378 (N_13378,N_12181,N_12593);
xnor U13379 (N_13379,N_12050,N_12161);
or U13380 (N_13380,N_12266,N_12729);
nor U13381 (N_13381,N_12396,N_12173);
xnor U13382 (N_13382,N_12177,N_12491);
or U13383 (N_13383,N_12070,N_12343);
xnor U13384 (N_13384,N_12589,N_12739);
nor U13385 (N_13385,N_12122,N_12699);
xnor U13386 (N_13386,N_12321,N_12032);
or U13387 (N_13387,N_12411,N_12087);
and U13388 (N_13388,N_12515,N_12558);
xor U13389 (N_13389,N_12342,N_12233);
or U13390 (N_13390,N_12289,N_12775);
nand U13391 (N_13391,N_12233,N_12259);
xnor U13392 (N_13392,N_12230,N_12245);
xor U13393 (N_13393,N_12385,N_12154);
or U13394 (N_13394,N_12755,N_12185);
nor U13395 (N_13395,N_12631,N_12475);
nor U13396 (N_13396,N_12629,N_12693);
nand U13397 (N_13397,N_12208,N_12263);
xnor U13398 (N_13398,N_12543,N_12165);
nor U13399 (N_13399,N_12591,N_12498);
nand U13400 (N_13400,N_12702,N_12645);
xnor U13401 (N_13401,N_12410,N_12529);
nor U13402 (N_13402,N_12254,N_12033);
nor U13403 (N_13403,N_12041,N_12613);
xnor U13404 (N_13404,N_12231,N_12282);
or U13405 (N_13405,N_12209,N_12091);
and U13406 (N_13406,N_12151,N_12224);
or U13407 (N_13407,N_12296,N_12586);
or U13408 (N_13408,N_12669,N_12491);
or U13409 (N_13409,N_12003,N_12546);
nor U13410 (N_13410,N_12119,N_12677);
nand U13411 (N_13411,N_12442,N_12249);
and U13412 (N_13412,N_12194,N_12667);
xor U13413 (N_13413,N_12488,N_12584);
or U13414 (N_13414,N_12630,N_12131);
and U13415 (N_13415,N_12217,N_12258);
nand U13416 (N_13416,N_12145,N_12765);
nor U13417 (N_13417,N_12619,N_12197);
xnor U13418 (N_13418,N_12596,N_12262);
and U13419 (N_13419,N_12317,N_12305);
nor U13420 (N_13420,N_12326,N_12347);
xnor U13421 (N_13421,N_12511,N_12007);
nor U13422 (N_13422,N_12214,N_12145);
or U13423 (N_13423,N_12079,N_12035);
or U13424 (N_13424,N_12011,N_12080);
xor U13425 (N_13425,N_12725,N_12478);
nand U13426 (N_13426,N_12793,N_12123);
and U13427 (N_13427,N_12051,N_12432);
xnor U13428 (N_13428,N_12140,N_12099);
and U13429 (N_13429,N_12336,N_12072);
nand U13430 (N_13430,N_12179,N_12379);
or U13431 (N_13431,N_12623,N_12193);
or U13432 (N_13432,N_12703,N_12529);
nor U13433 (N_13433,N_12258,N_12023);
and U13434 (N_13434,N_12043,N_12169);
and U13435 (N_13435,N_12251,N_12680);
nand U13436 (N_13436,N_12300,N_12749);
nand U13437 (N_13437,N_12491,N_12000);
xor U13438 (N_13438,N_12618,N_12460);
xor U13439 (N_13439,N_12207,N_12694);
and U13440 (N_13440,N_12339,N_12108);
xnor U13441 (N_13441,N_12791,N_12727);
or U13442 (N_13442,N_12373,N_12561);
and U13443 (N_13443,N_12657,N_12327);
xor U13444 (N_13444,N_12326,N_12133);
and U13445 (N_13445,N_12430,N_12797);
nand U13446 (N_13446,N_12147,N_12669);
xor U13447 (N_13447,N_12224,N_12249);
nor U13448 (N_13448,N_12200,N_12790);
and U13449 (N_13449,N_12475,N_12227);
and U13450 (N_13450,N_12119,N_12162);
xnor U13451 (N_13451,N_12453,N_12161);
xnor U13452 (N_13452,N_12078,N_12120);
nor U13453 (N_13453,N_12000,N_12287);
nand U13454 (N_13454,N_12439,N_12236);
nand U13455 (N_13455,N_12145,N_12665);
nor U13456 (N_13456,N_12348,N_12373);
nor U13457 (N_13457,N_12334,N_12438);
nand U13458 (N_13458,N_12318,N_12522);
nor U13459 (N_13459,N_12604,N_12213);
or U13460 (N_13460,N_12543,N_12595);
and U13461 (N_13461,N_12031,N_12442);
nor U13462 (N_13462,N_12622,N_12665);
and U13463 (N_13463,N_12378,N_12379);
nor U13464 (N_13464,N_12366,N_12141);
or U13465 (N_13465,N_12662,N_12546);
or U13466 (N_13466,N_12042,N_12789);
nand U13467 (N_13467,N_12651,N_12003);
nand U13468 (N_13468,N_12786,N_12666);
or U13469 (N_13469,N_12719,N_12461);
nor U13470 (N_13470,N_12414,N_12508);
and U13471 (N_13471,N_12001,N_12310);
xor U13472 (N_13472,N_12337,N_12015);
or U13473 (N_13473,N_12290,N_12363);
nand U13474 (N_13474,N_12727,N_12193);
nand U13475 (N_13475,N_12502,N_12197);
xor U13476 (N_13476,N_12150,N_12045);
and U13477 (N_13477,N_12144,N_12566);
and U13478 (N_13478,N_12740,N_12202);
nor U13479 (N_13479,N_12770,N_12058);
nor U13480 (N_13480,N_12550,N_12124);
nand U13481 (N_13481,N_12541,N_12450);
nand U13482 (N_13482,N_12281,N_12479);
nand U13483 (N_13483,N_12795,N_12701);
nor U13484 (N_13484,N_12653,N_12015);
or U13485 (N_13485,N_12589,N_12213);
xor U13486 (N_13486,N_12163,N_12678);
nand U13487 (N_13487,N_12306,N_12683);
and U13488 (N_13488,N_12658,N_12054);
and U13489 (N_13489,N_12406,N_12280);
and U13490 (N_13490,N_12643,N_12789);
nor U13491 (N_13491,N_12152,N_12342);
or U13492 (N_13492,N_12122,N_12280);
xor U13493 (N_13493,N_12096,N_12591);
nor U13494 (N_13494,N_12397,N_12744);
or U13495 (N_13495,N_12170,N_12000);
nand U13496 (N_13496,N_12155,N_12711);
nand U13497 (N_13497,N_12667,N_12674);
nor U13498 (N_13498,N_12148,N_12636);
and U13499 (N_13499,N_12556,N_12757);
nand U13500 (N_13500,N_12393,N_12633);
nand U13501 (N_13501,N_12115,N_12127);
and U13502 (N_13502,N_12605,N_12571);
nand U13503 (N_13503,N_12143,N_12575);
nand U13504 (N_13504,N_12352,N_12026);
and U13505 (N_13505,N_12235,N_12189);
nand U13506 (N_13506,N_12321,N_12324);
or U13507 (N_13507,N_12317,N_12613);
xnor U13508 (N_13508,N_12056,N_12094);
nor U13509 (N_13509,N_12715,N_12041);
xnor U13510 (N_13510,N_12524,N_12037);
or U13511 (N_13511,N_12212,N_12432);
and U13512 (N_13512,N_12701,N_12757);
nor U13513 (N_13513,N_12764,N_12637);
nor U13514 (N_13514,N_12585,N_12213);
or U13515 (N_13515,N_12201,N_12210);
nand U13516 (N_13516,N_12057,N_12657);
nor U13517 (N_13517,N_12244,N_12621);
nand U13518 (N_13518,N_12053,N_12074);
xor U13519 (N_13519,N_12126,N_12231);
and U13520 (N_13520,N_12557,N_12753);
and U13521 (N_13521,N_12236,N_12341);
or U13522 (N_13522,N_12736,N_12059);
and U13523 (N_13523,N_12725,N_12074);
or U13524 (N_13524,N_12550,N_12691);
nand U13525 (N_13525,N_12033,N_12197);
xor U13526 (N_13526,N_12631,N_12392);
nor U13527 (N_13527,N_12161,N_12304);
xor U13528 (N_13528,N_12758,N_12155);
nor U13529 (N_13529,N_12551,N_12327);
and U13530 (N_13530,N_12751,N_12451);
nand U13531 (N_13531,N_12264,N_12016);
nor U13532 (N_13532,N_12214,N_12558);
nand U13533 (N_13533,N_12137,N_12071);
and U13534 (N_13534,N_12288,N_12368);
nand U13535 (N_13535,N_12782,N_12772);
or U13536 (N_13536,N_12282,N_12312);
xnor U13537 (N_13537,N_12638,N_12196);
xor U13538 (N_13538,N_12785,N_12042);
nor U13539 (N_13539,N_12220,N_12202);
xnor U13540 (N_13540,N_12529,N_12797);
nor U13541 (N_13541,N_12293,N_12655);
xnor U13542 (N_13542,N_12307,N_12617);
nor U13543 (N_13543,N_12405,N_12385);
xor U13544 (N_13544,N_12736,N_12717);
nand U13545 (N_13545,N_12778,N_12672);
and U13546 (N_13546,N_12241,N_12511);
and U13547 (N_13547,N_12770,N_12265);
nand U13548 (N_13548,N_12544,N_12725);
nand U13549 (N_13549,N_12514,N_12384);
and U13550 (N_13550,N_12553,N_12486);
nor U13551 (N_13551,N_12622,N_12573);
and U13552 (N_13552,N_12453,N_12793);
nand U13553 (N_13553,N_12109,N_12125);
nand U13554 (N_13554,N_12573,N_12535);
nand U13555 (N_13555,N_12354,N_12232);
nand U13556 (N_13556,N_12038,N_12535);
nand U13557 (N_13557,N_12348,N_12371);
or U13558 (N_13558,N_12716,N_12109);
xnor U13559 (N_13559,N_12300,N_12788);
xnor U13560 (N_13560,N_12508,N_12661);
xor U13561 (N_13561,N_12458,N_12482);
and U13562 (N_13562,N_12483,N_12109);
nand U13563 (N_13563,N_12139,N_12082);
and U13564 (N_13564,N_12556,N_12746);
xor U13565 (N_13565,N_12300,N_12746);
or U13566 (N_13566,N_12564,N_12348);
and U13567 (N_13567,N_12335,N_12596);
xnor U13568 (N_13568,N_12462,N_12229);
nor U13569 (N_13569,N_12334,N_12487);
or U13570 (N_13570,N_12139,N_12324);
and U13571 (N_13571,N_12791,N_12585);
nand U13572 (N_13572,N_12759,N_12465);
nand U13573 (N_13573,N_12631,N_12300);
or U13574 (N_13574,N_12532,N_12087);
and U13575 (N_13575,N_12766,N_12241);
and U13576 (N_13576,N_12105,N_12013);
or U13577 (N_13577,N_12538,N_12065);
and U13578 (N_13578,N_12090,N_12034);
or U13579 (N_13579,N_12675,N_12416);
nor U13580 (N_13580,N_12303,N_12179);
nand U13581 (N_13581,N_12404,N_12111);
nor U13582 (N_13582,N_12646,N_12253);
nor U13583 (N_13583,N_12660,N_12778);
nand U13584 (N_13584,N_12767,N_12427);
nand U13585 (N_13585,N_12437,N_12692);
or U13586 (N_13586,N_12735,N_12333);
nor U13587 (N_13587,N_12528,N_12286);
xnor U13588 (N_13588,N_12215,N_12316);
xor U13589 (N_13589,N_12585,N_12142);
xnor U13590 (N_13590,N_12570,N_12422);
and U13591 (N_13591,N_12121,N_12502);
xnor U13592 (N_13592,N_12769,N_12608);
xnor U13593 (N_13593,N_12332,N_12039);
and U13594 (N_13594,N_12161,N_12206);
or U13595 (N_13595,N_12364,N_12276);
nor U13596 (N_13596,N_12734,N_12021);
xor U13597 (N_13597,N_12797,N_12349);
nor U13598 (N_13598,N_12240,N_12534);
or U13599 (N_13599,N_12571,N_12780);
and U13600 (N_13600,N_13534,N_13581);
nor U13601 (N_13601,N_13026,N_13542);
and U13602 (N_13602,N_13508,N_13246);
and U13603 (N_13603,N_12940,N_13171);
xor U13604 (N_13604,N_12901,N_13566);
xor U13605 (N_13605,N_13206,N_13055);
or U13606 (N_13606,N_13091,N_13428);
xnor U13607 (N_13607,N_12995,N_12977);
and U13608 (N_13608,N_12947,N_13022);
nand U13609 (N_13609,N_13072,N_13362);
nand U13610 (N_13610,N_13369,N_13045);
xnor U13611 (N_13611,N_13105,N_13284);
xnor U13612 (N_13612,N_13180,N_13108);
nand U13613 (N_13613,N_13219,N_13495);
nand U13614 (N_13614,N_13043,N_13253);
xnor U13615 (N_13615,N_13133,N_13558);
and U13616 (N_13616,N_13524,N_13194);
and U13617 (N_13617,N_13032,N_12954);
nor U13618 (N_13618,N_13274,N_13373);
and U13619 (N_13619,N_13443,N_12882);
and U13620 (N_13620,N_12819,N_13233);
and U13621 (N_13621,N_13323,N_13367);
and U13622 (N_13622,N_13132,N_13299);
and U13623 (N_13623,N_13537,N_13068);
xor U13624 (N_13624,N_12859,N_12806);
or U13625 (N_13625,N_13058,N_13151);
or U13626 (N_13626,N_13097,N_13118);
nor U13627 (N_13627,N_13391,N_12937);
or U13628 (N_13628,N_13498,N_12847);
and U13629 (N_13629,N_13135,N_13479);
or U13630 (N_13630,N_13520,N_13444);
xor U13631 (N_13631,N_12986,N_12851);
nor U13632 (N_13632,N_13514,N_12969);
and U13633 (N_13633,N_13150,N_12918);
and U13634 (N_13634,N_13156,N_12934);
xnor U13635 (N_13635,N_13185,N_13557);
and U13636 (N_13636,N_12990,N_13110);
nand U13637 (N_13637,N_13376,N_13510);
and U13638 (N_13638,N_13139,N_13169);
nand U13639 (N_13639,N_12822,N_12867);
or U13640 (N_13640,N_13241,N_13073);
or U13641 (N_13641,N_12972,N_12820);
xnor U13642 (N_13642,N_13315,N_13014);
xnor U13643 (N_13643,N_13506,N_13075);
and U13644 (N_13644,N_13485,N_13296);
nand U13645 (N_13645,N_13387,N_13287);
or U13646 (N_13646,N_13399,N_12854);
xnor U13647 (N_13647,N_13433,N_12996);
and U13648 (N_13648,N_13006,N_13407);
and U13649 (N_13649,N_13061,N_12805);
or U13650 (N_13650,N_13504,N_13278);
xor U13651 (N_13651,N_13333,N_13039);
nor U13652 (N_13652,N_13568,N_13594);
or U13653 (N_13653,N_13567,N_13402);
or U13654 (N_13654,N_12932,N_13067);
xnor U13655 (N_13655,N_12965,N_13466);
or U13656 (N_13656,N_13128,N_13578);
nor U13657 (N_13657,N_13442,N_12912);
and U13658 (N_13658,N_13228,N_12823);
xnor U13659 (N_13659,N_13462,N_12998);
nand U13660 (N_13660,N_13174,N_13147);
nor U13661 (N_13661,N_13168,N_13280);
nand U13662 (N_13662,N_12983,N_13413);
or U13663 (N_13663,N_13213,N_13234);
nand U13664 (N_13664,N_12804,N_13307);
nor U13665 (N_13665,N_12922,N_13175);
xnor U13666 (N_13666,N_13124,N_13029);
nor U13667 (N_13667,N_13321,N_13334);
nand U13668 (N_13668,N_12833,N_13145);
nor U13669 (N_13669,N_12840,N_13205);
or U13670 (N_13670,N_13208,N_12900);
or U13671 (N_13671,N_13358,N_13488);
xor U13672 (N_13672,N_12881,N_13515);
and U13673 (N_13673,N_12907,N_13183);
and U13674 (N_13674,N_13117,N_13056);
or U13675 (N_13675,N_13503,N_12930);
nand U13676 (N_13676,N_13035,N_13390);
nand U13677 (N_13677,N_13393,N_13003);
and U13678 (N_13678,N_13597,N_13409);
or U13679 (N_13679,N_12843,N_13497);
and U13680 (N_13680,N_13541,N_13474);
nor U13681 (N_13681,N_13157,N_13562);
or U13682 (N_13682,N_12814,N_12908);
xor U13683 (N_13683,N_12803,N_12878);
xnor U13684 (N_13684,N_12890,N_13395);
nand U13685 (N_13685,N_12839,N_13220);
xor U13686 (N_13686,N_13312,N_13001);
or U13687 (N_13687,N_12862,N_13554);
nand U13688 (N_13688,N_13584,N_12999);
and U13689 (N_13689,N_12910,N_13215);
xor U13690 (N_13690,N_12821,N_13107);
xnor U13691 (N_13691,N_13187,N_12985);
nand U13692 (N_13692,N_12923,N_13109);
nand U13693 (N_13693,N_13300,N_13364);
xor U13694 (N_13694,N_13487,N_13521);
xor U13695 (N_13695,N_13222,N_13533);
nand U13696 (N_13696,N_13027,N_13350);
nand U13697 (N_13697,N_13465,N_13528);
nand U13698 (N_13698,N_13481,N_13502);
nand U13699 (N_13699,N_13083,N_13327);
and U13700 (N_13700,N_13282,N_12898);
and U13701 (N_13701,N_13539,N_13448);
nor U13702 (N_13702,N_13404,N_13293);
or U13703 (N_13703,N_12921,N_12861);
nor U13704 (N_13704,N_13527,N_12849);
nor U13705 (N_13705,N_12993,N_13082);
and U13706 (N_13706,N_13152,N_12809);
nand U13707 (N_13707,N_13181,N_13231);
nor U13708 (N_13708,N_13057,N_13200);
nor U13709 (N_13709,N_13306,N_13529);
or U13710 (N_13710,N_13530,N_13144);
nor U13711 (N_13711,N_13400,N_12870);
and U13712 (N_13712,N_13389,N_13463);
xnor U13713 (N_13713,N_13033,N_13450);
nor U13714 (N_13714,N_13211,N_13326);
nor U13715 (N_13715,N_13071,N_13398);
or U13716 (N_13716,N_12869,N_13113);
xnor U13717 (N_13717,N_12879,N_13344);
xnor U13718 (N_13718,N_13551,N_13210);
nand U13719 (N_13719,N_12962,N_13297);
nand U13720 (N_13720,N_13374,N_13491);
and U13721 (N_13721,N_13511,N_13453);
nand U13722 (N_13722,N_13002,N_13074);
xnor U13723 (N_13723,N_13254,N_13161);
or U13724 (N_13724,N_13204,N_13189);
nand U13725 (N_13725,N_13346,N_12974);
and U13726 (N_13726,N_13456,N_13249);
or U13727 (N_13727,N_12987,N_13019);
or U13728 (N_13728,N_13199,N_13025);
nor U13729 (N_13729,N_13090,N_12812);
nand U13730 (N_13730,N_13532,N_13207);
nor U13731 (N_13731,N_13264,N_12897);
xnor U13732 (N_13732,N_12975,N_13375);
nand U13733 (N_13733,N_13218,N_13190);
nand U13734 (N_13734,N_13182,N_13084);
or U13735 (N_13735,N_13353,N_13011);
nor U13736 (N_13736,N_12831,N_13329);
nand U13737 (N_13737,N_13094,N_12951);
nand U13738 (N_13738,N_13411,N_13243);
and U13739 (N_13739,N_12845,N_13010);
nand U13740 (N_13740,N_12802,N_12844);
nor U13741 (N_13741,N_13425,N_12949);
or U13742 (N_13742,N_12846,N_12832);
nand U13743 (N_13743,N_12935,N_13272);
or U13744 (N_13744,N_13547,N_13403);
nand U13745 (N_13745,N_13309,N_13553);
and U13746 (N_13746,N_12991,N_13357);
or U13747 (N_13747,N_13436,N_13359);
xnor U13748 (N_13748,N_13085,N_13125);
nand U13749 (N_13749,N_13447,N_13098);
and U13750 (N_13750,N_13494,N_13081);
or U13751 (N_13751,N_13561,N_13038);
and U13752 (N_13752,N_12971,N_13062);
nor U13753 (N_13753,N_13483,N_12834);
or U13754 (N_13754,N_13324,N_12958);
nand U13755 (N_13755,N_12904,N_13516);
nor U13756 (N_13756,N_13020,N_13470);
and U13757 (N_13757,N_13066,N_13192);
and U13758 (N_13758,N_13418,N_12984);
and U13759 (N_13759,N_12945,N_13587);
nand U13760 (N_13760,N_13155,N_13088);
or U13761 (N_13761,N_13341,N_13355);
nand U13762 (N_13762,N_13103,N_13500);
nand U13763 (N_13763,N_13356,N_13507);
xor U13764 (N_13764,N_13560,N_12929);
or U13765 (N_13765,N_13401,N_13040);
and U13766 (N_13766,N_13240,N_12810);
nor U13767 (N_13767,N_13165,N_12813);
xor U13768 (N_13768,N_13096,N_13095);
and U13769 (N_13769,N_13188,N_13009);
xnor U13770 (N_13770,N_12961,N_13477);
nand U13771 (N_13771,N_13114,N_12976);
nor U13772 (N_13772,N_13381,N_13251);
xnor U13773 (N_13773,N_13505,N_13415);
nand U13774 (N_13774,N_12902,N_13538);
and U13775 (N_13775,N_13454,N_13386);
nor U13776 (N_13776,N_13338,N_13260);
nand U13777 (N_13777,N_13340,N_13146);
nor U13778 (N_13778,N_13476,N_12994);
and U13779 (N_13779,N_13288,N_12919);
nor U13780 (N_13780,N_13173,N_13069);
and U13781 (N_13781,N_13252,N_12928);
and U13782 (N_13782,N_12926,N_12948);
and U13783 (N_13783,N_12939,N_13596);
nor U13784 (N_13784,N_13179,N_13053);
nand U13785 (N_13785,N_12876,N_13544);
or U13786 (N_13786,N_13130,N_13232);
or U13787 (N_13787,N_13408,N_13255);
and U13788 (N_13788,N_13429,N_13149);
or U13789 (N_13789,N_13570,N_13384);
and U13790 (N_13790,N_13380,N_13250);
or U13791 (N_13791,N_12953,N_12905);
nand U13792 (N_13792,N_13064,N_13572);
nor U13793 (N_13793,N_12992,N_13079);
or U13794 (N_13794,N_13267,N_13410);
or U13795 (N_13795,N_13115,N_13354);
or U13796 (N_13796,N_13298,N_13431);
nand U13797 (N_13797,N_13414,N_12946);
xor U13798 (N_13798,N_13184,N_12891);
or U13799 (N_13799,N_13478,N_13311);
or U13800 (N_13800,N_13087,N_13080);
or U13801 (N_13801,N_13049,N_13577);
xor U13802 (N_13802,N_13259,N_12981);
or U13803 (N_13803,N_13592,N_12887);
or U13804 (N_13804,N_12927,N_12880);
nor U13805 (N_13805,N_13116,N_12853);
nand U13806 (N_13806,N_13154,N_12857);
nand U13807 (N_13807,N_13522,N_13366);
nor U13808 (N_13808,N_13123,N_13129);
or U13809 (N_13809,N_13590,N_13256);
nor U13810 (N_13810,N_13370,N_13313);
or U13811 (N_13811,N_12864,N_13261);
nand U13812 (N_13812,N_13037,N_13330);
and U13813 (N_13813,N_13159,N_13092);
nor U13814 (N_13814,N_13316,N_12877);
and U13815 (N_13815,N_13000,N_13583);
nand U13816 (N_13816,N_13588,N_13172);
nor U13817 (N_13817,N_12875,N_13054);
xnor U13818 (N_13818,N_13435,N_13238);
xor U13819 (N_13819,N_12850,N_13441);
nor U13820 (N_13820,N_12873,N_12826);
or U13821 (N_13821,N_12944,N_13556);
nand U13822 (N_13822,N_13106,N_13430);
or U13823 (N_13823,N_13289,N_13266);
nor U13824 (N_13824,N_13127,N_13499);
and U13825 (N_13825,N_12842,N_12988);
nand U13826 (N_13826,N_12906,N_13265);
and U13827 (N_13827,N_12896,N_12943);
and U13828 (N_13828,N_13276,N_12893);
or U13829 (N_13829,N_13439,N_13004);
nand U13830 (N_13830,N_13385,N_12848);
xor U13831 (N_13831,N_13216,N_13427);
or U13832 (N_13832,N_13093,N_13416);
and U13833 (N_13833,N_13575,N_13305);
nand U13834 (N_13834,N_12825,N_13349);
and U13835 (N_13835,N_13531,N_13193);
nor U13836 (N_13836,N_13226,N_13047);
xnor U13837 (N_13837,N_12978,N_13018);
xor U13838 (N_13838,N_13153,N_13164);
nor U13839 (N_13839,N_13290,N_13351);
or U13840 (N_13840,N_13482,N_13457);
xnor U13841 (N_13841,N_12933,N_13424);
nor U13842 (N_13842,N_12916,N_13143);
and U13843 (N_13843,N_13475,N_13163);
or U13844 (N_13844,N_12889,N_13137);
nand U13845 (N_13845,N_12852,N_13519);
nor U13846 (N_13846,N_13569,N_12966);
nand U13847 (N_13847,N_12968,N_13052);
nand U13848 (N_13848,N_13270,N_12980);
xnor U13849 (N_13849,N_13166,N_12835);
nand U13850 (N_13850,N_13335,N_13523);
nand U13851 (N_13851,N_13046,N_12957);
xnor U13852 (N_13852,N_13438,N_13455);
nor U13853 (N_13853,N_13573,N_13574);
nand U13854 (N_13854,N_12963,N_12816);
and U13855 (N_13855,N_13480,N_13065);
nand U13856 (N_13856,N_12829,N_13247);
nor U13857 (N_13857,N_13236,N_13513);
nor U13858 (N_13858,N_13191,N_12911);
nand U13859 (N_13859,N_13360,N_13445);
nand U13860 (N_13860,N_13227,N_13034);
xor U13861 (N_13861,N_13509,N_13501);
and U13862 (N_13862,N_13012,N_13229);
and U13863 (N_13863,N_13593,N_12950);
nor U13864 (N_13864,N_13013,N_13294);
and U13865 (N_13865,N_13469,N_13176);
xor U13866 (N_13866,N_13464,N_13459);
nor U13867 (N_13867,N_13365,N_12863);
nand U13868 (N_13868,N_12903,N_13111);
nand U13869 (N_13869,N_13060,N_12885);
or U13870 (N_13870,N_13239,N_12925);
and U13871 (N_13871,N_13201,N_13277);
or U13872 (N_13872,N_13015,N_13472);
nand U13873 (N_13873,N_13031,N_13248);
or U13874 (N_13874,N_12913,N_13197);
or U13875 (N_13875,N_13467,N_13526);
xor U13876 (N_13876,N_13304,N_13394);
xnor U13877 (N_13877,N_13063,N_12868);
nor U13878 (N_13878,N_13451,N_12828);
or U13879 (N_13879,N_13432,N_13372);
and U13880 (N_13880,N_13285,N_12872);
nand U13881 (N_13881,N_13078,N_13552);
and U13882 (N_13882,N_13468,N_13262);
nand U13883 (N_13883,N_13412,N_13382);
and U13884 (N_13884,N_12827,N_13217);
nor U13885 (N_13885,N_13490,N_13585);
and U13886 (N_13886,N_13126,N_13017);
and U13887 (N_13887,N_13405,N_13050);
and U13888 (N_13888,N_13122,N_12955);
or U13889 (N_13889,N_13271,N_13279);
xnor U13890 (N_13890,N_13048,N_12973);
and U13891 (N_13891,N_13203,N_13377);
and U13892 (N_13892,N_13589,N_13540);
and U13893 (N_13893,N_12895,N_13437);
or U13894 (N_13894,N_12979,N_13212);
xor U13895 (N_13895,N_13317,N_13582);
or U13896 (N_13896,N_12915,N_13286);
xnor U13897 (N_13897,N_13347,N_12960);
or U13898 (N_13898,N_12837,N_13077);
nand U13899 (N_13899,N_12914,N_13564);
xor U13900 (N_13900,N_13016,N_12811);
and U13901 (N_13901,N_13028,N_13244);
nand U13902 (N_13902,N_13426,N_12856);
and U13903 (N_13903,N_13120,N_13396);
xor U13904 (N_13904,N_13224,N_13059);
nor U13905 (N_13905,N_13104,N_13195);
and U13906 (N_13906,N_13517,N_13525);
xnor U13907 (N_13907,N_13337,N_13598);
xnor U13908 (N_13908,N_13548,N_12836);
nor U13909 (N_13909,N_13140,N_13202);
and U13910 (N_13910,N_13257,N_13101);
xor U13911 (N_13911,N_13167,N_13361);
nor U13912 (N_13912,N_13258,N_13342);
nor U13913 (N_13913,N_13158,N_13245);
or U13914 (N_13914,N_13112,N_12807);
and U13915 (N_13915,N_12884,N_12941);
xnor U13916 (N_13916,N_13417,N_13141);
nor U13917 (N_13917,N_13392,N_13269);
xor U13918 (N_13918,N_13230,N_13089);
nor U13919 (N_13919,N_13328,N_13492);
nand U13920 (N_13920,N_13363,N_12967);
xor U13921 (N_13921,N_13545,N_12841);
or U13922 (N_13922,N_12959,N_13136);
xor U13923 (N_13923,N_12970,N_13580);
nand U13924 (N_13924,N_12838,N_13586);
nand U13925 (N_13925,N_13452,N_13100);
or U13926 (N_13926,N_13295,N_13461);
xor U13927 (N_13927,N_13599,N_12815);
xor U13928 (N_13928,N_13565,N_13419);
xor U13929 (N_13929,N_13378,N_13237);
xor U13930 (N_13930,N_13449,N_13024);
nand U13931 (N_13931,N_12997,N_13302);
nor U13932 (N_13932,N_12855,N_12909);
and U13933 (N_13933,N_13331,N_12989);
xnor U13934 (N_13934,N_13005,N_13235);
xnor U13935 (N_13935,N_13422,N_13446);
and U13936 (N_13936,N_13379,N_13512);
nor U13937 (N_13937,N_13555,N_13579);
or U13938 (N_13938,N_13162,N_13352);
nand U13939 (N_13939,N_12894,N_13322);
xor U13940 (N_13940,N_12800,N_13339);
nor U13941 (N_13941,N_13423,N_12871);
and U13942 (N_13942,N_13051,N_13198);
and U13943 (N_13943,N_12860,N_12892);
nand U13944 (N_13944,N_13223,N_12952);
nor U13945 (N_13945,N_13186,N_13397);
nor U13946 (N_13946,N_13308,N_13434);
xnor U13947 (N_13947,N_13268,N_12917);
or U13948 (N_13948,N_13310,N_13242);
nor U13949 (N_13949,N_13042,N_13460);
or U13950 (N_13950,N_13160,N_13292);
nor U13951 (N_13951,N_13214,N_13543);
nor U13952 (N_13952,N_13225,N_13086);
nand U13953 (N_13953,N_13371,N_13021);
nand U13954 (N_13954,N_13489,N_12801);
nor U13955 (N_13955,N_13406,N_13332);
xor U13956 (N_13956,N_13099,N_12924);
nor U13957 (N_13957,N_13576,N_12942);
or U13958 (N_13958,N_13076,N_13134);
and U13959 (N_13959,N_13170,N_13301);
nand U13960 (N_13960,N_12938,N_13007);
nand U13961 (N_13961,N_13440,N_13023);
and U13962 (N_13962,N_13473,N_12936);
nand U13963 (N_13963,N_13549,N_13142);
xnor U13964 (N_13964,N_12920,N_12817);
xor U13965 (N_13965,N_13036,N_12865);
or U13966 (N_13966,N_12888,N_13421);
or U13967 (N_13967,N_13131,N_13383);
nor U13968 (N_13968,N_12883,N_13221);
and U13969 (N_13969,N_13044,N_13177);
xor U13970 (N_13970,N_13291,N_13420);
nand U13971 (N_13971,N_13283,N_12886);
and U13972 (N_13972,N_13121,N_13041);
nor U13973 (N_13973,N_13348,N_13550);
and U13974 (N_13974,N_13546,N_12931);
nor U13975 (N_13975,N_13102,N_13536);
xnor U13976 (N_13976,N_13535,N_13320);
nor U13977 (N_13977,N_12899,N_13281);
or U13978 (N_13978,N_13325,N_12808);
nor U13979 (N_13979,N_12830,N_13008);
and U13980 (N_13980,N_13319,N_13070);
or U13981 (N_13981,N_13318,N_13343);
or U13982 (N_13982,N_12964,N_13119);
nand U13983 (N_13983,N_13496,N_13196);
or U13984 (N_13984,N_13314,N_13518);
or U13985 (N_13985,N_13563,N_13471);
nand U13986 (N_13986,N_12956,N_13571);
or U13987 (N_13987,N_13484,N_13486);
xor U13988 (N_13988,N_12858,N_13030);
and U13989 (N_13989,N_13493,N_13138);
or U13990 (N_13990,N_13591,N_13345);
and U13991 (N_13991,N_13559,N_12982);
nand U13992 (N_13992,N_13458,N_13275);
nand U13993 (N_13993,N_13595,N_12824);
or U13994 (N_13994,N_13209,N_12818);
nor U13995 (N_13995,N_13303,N_13148);
xor U13996 (N_13996,N_13178,N_13263);
nor U13997 (N_13997,N_13273,N_13368);
xor U13998 (N_13998,N_13336,N_12874);
nand U13999 (N_13999,N_12866,N_13388);
nor U14000 (N_14000,N_13500,N_13027);
nor U14001 (N_14001,N_12955,N_13136);
xnor U14002 (N_14002,N_13074,N_13344);
and U14003 (N_14003,N_12860,N_13572);
nor U14004 (N_14004,N_12805,N_13251);
nand U14005 (N_14005,N_13096,N_12833);
nor U14006 (N_14006,N_13107,N_13465);
nor U14007 (N_14007,N_13228,N_13168);
xor U14008 (N_14008,N_13251,N_13178);
or U14009 (N_14009,N_12816,N_13260);
nand U14010 (N_14010,N_13243,N_12887);
nor U14011 (N_14011,N_13441,N_13484);
and U14012 (N_14012,N_13483,N_13427);
xor U14013 (N_14013,N_13036,N_13392);
xor U14014 (N_14014,N_12912,N_13261);
xnor U14015 (N_14015,N_12976,N_13344);
or U14016 (N_14016,N_13286,N_13110);
nand U14017 (N_14017,N_13088,N_13288);
nor U14018 (N_14018,N_13068,N_13309);
and U14019 (N_14019,N_13314,N_12957);
and U14020 (N_14020,N_12926,N_13224);
xnor U14021 (N_14021,N_12932,N_13199);
xor U14022 (N_14022,N_13157,N_13331);
nand U14023 (N_14023,N_13057,N_13216);
nand U14024 (N_14024,N_12896,N_13108);
xnor U14025 (N_14025,N_13381,N_13197);
or U14026 (N_14026,N_12874,N_12885);
or U14027 (N_14027,N_13394,N_13495);
xnor U14028 (N_14028,N_13326,N_13434);
xnor U14029 (N_14029,N_13422,N_12802);
and U14030 (N_14030,N_12897,N_13105);
and U14031 (N_14031,N_13345,N_13050);
nor U14032 (N_14032,N_13320,N_12930);
and U14033 (N_14033,N_13082,N_12848);
nand U14034 (N_14034,N_12866,N_12830);
or U14035 (N_14035,N_13370,N_13288);
nand U14036 (N_14036,N_12896,N_12941);
nor U14037 (N_14037,N_13449,N_13109);
nand U14038 (N_14038,N_13011,N_13306);
nor U14039 (N_14039,N_13594,N_13550);
xnor U14040 (N_14040,N_13190,N_13050);
nand U14041 (N_14041,N_13459,N_13335);
xor U14042 (N_14042,N_13030,N_12911);
xor U14043 (N_14043,N_12843,N_12943);
and U14044 (N_14044,N_13575,N_13197);
nand U14045 (N_14045,N_13434,N_13227);
nor U14046 (N_14046,N_13160,N_12977);
or U14047 (N_14047,N_13467,N_13045);
nor U14048 (N_14048,N_12998,N_13137);
xnor U14049 (N_14049,N_13435,N_13523);
nor U14050 (N_14050,N_13068,N_13576);
nor U14051 (N_14051,N_13595,N_13323);
xnor U14052 (N_14052,N_13202,N_13034);
nand U14053 (N_14053,N_13234,N_13475);
nand U14054 (N_14054,N_13164,N_13007);
xor U14055 (N_14055,N_13579,N_12962);
and U14056 (N_14056,N_13257,N_13258);
xor U14057 (N_14057,N_12916,N_13199);
nand U14058 (N_14058,N_12939,N_13543);
nand U14059 (N_14059,N_12927,N_13378);
xor U14060 (N_14060,N_13376,N_13584);
or U14061 (N_14061,N_13412,N_13078);
nand U14062 (N_14062,N_13183,N_12956);
xnor U14063 (N_14063,N_13240,N_13542);
nor U14064 (N_14064,N_13217,N_12980);
nor U14065 (N_14065,N_13000,N_12984);
nor U14066 (N_14066,N_13201,N_13147);
xnor U14067 (N_14067,N_13102,N_13448);
nor U14068 (N_14068,N_13069,N_13298);
or U14069 (N_14069,N_13199,N_12837);
and U14070 (N_14070,N_13220,N_12876);
and U14071 (N_14071,N_13547,N_13204);
and U14072 (N_14072,N_13333,N_13511);
or U14073 (N_14073,N_13580,N_12800);
nand U14074 (N_14074,N_13114,N_13251);
and U14075 (N_14075,N_13021,N_13154);
nand U14076 (N_14076,N_13196,N_12924);
or U14077 (N_14077,N_12972,N_12814);
or U14078 (N_14078,N_12854,N_12814);
or U14079 (N_14079,N_13490,N_13267);
and U14080 (N_14080,N_13164,N_13360);
xor U14081 (N_14081,N_13598,N_12809);
nand U14082 (N_14082,N_13237,N_13593);
nor U14083 (N_14083,N_13155,N_13413);
or U14084 (N_14084,N_13357,N_13176);
nand U14085 (N_14085,N_12904,N_13545);
xor U14086 (N_14086,N_13268,N_12993);
nand U14087 (N_14087,N_12999,N_13173);
nor U14088 (N_14088,N_13572,N_13217);
and U14089 (N_14089,N_12860,N_13381);
xor U14090 (N_14090,N_13032,N_13380);
nand U14091 (N_14091,N_13509,N_12858);
nor U14092 (N_14092,N_13210,N_13521);
nor U14093 (N_14093,N_13400,N_13467);
nor U14094 (N_14094,N_13547,N_13146);
nand U14095 (N_14095,N_12922,N_12916);
nand U14096 (N_14096,N_13515,N_12863);
xnor U14097 (N_14097,N_12829,N_13399);
nand U14098 (N_14098,N_13212,N_13076);
xnor U14099 (N_14099,N_12930,N_13479);
and U14100 (N_14100,N_13489,N_13102);
nand U14101 (N_14101,N_12960,N_12986);
and U14102 (N_14102,N_13133,N_13323);
nor U14103 (N_14103,N_13302,N_13335);
nand U14104 (N_14104,N_13562,N_12942);
or U14105 (N_14105,N_13233,N_13270);
nand U14106 (N_14106,N_13594,N_12915);
or U14107 (N_14107,N_13125,N_12874);
and U14108 (N_14108,N_12970,N_13335);
nor U14109 (N_14109,N_13414,N_13366);
nand U14110 (N_14110,N_13071,N_13544);
and U14111 (N_14111,N_13222,N_12907);
xor U14112 (N_14112,N_12933,N_12879);
and U14113 (N_14113,N_12994,N_13056);
or U14114 (N_14114,N_13128,N_13426);
nor U14115 (N_14115,N_13537,N_13219);
and U14116 (N_14116,N_12937,N_13145);
nor U14117 (N_14117,N_12952,N_13199);
nand U14118 (N_14118,N_13547,N_12847);
nor U14119 (N_14119,N_13175,N_13123);
xnor U14120 (N_14120,N_13231,N_13538);
and U14121 (N_14121,N_13055,N_13368);
and U14122 (N_14122,N_13244,N_13187);
nand U14123 (N_14123,N_13073,N_13101);
or U14124 (N_14124,N_13003,N_13227);
nor U14125 (N_14125,N_13439,N_12869);
xnor U14126 (N_14126,N_13094,N_13284);
nor U14127 (N_14127,N_13091,N_13346);
or U14128 (N_14128,N_13483,N_13055);
nand U14129 (N_14129,N_13232,N_12826);
or U14130 (N_14130,N_13552,N_12953);
xnor U14131 (N_14131,N_13005,N_13480);
nand U14132 (N_14132,N_13133,N_12886);
nor U14133 (N_14133,N_13258,N_13420);
nand U14134 (N_14134,N_12834,N_12957);
and U14135 (N_14135,N_13107,N_12974);
or U14136 (N_14136,N_13246,N_13424);
xnor U14137 (N_14137,N_13180,N_13456);
and U14138 (N_14138,N_12928,N_13424);
nand U14139 (N_14139,N_13296,N_13546);
nor U14140 (N_14140,N_12977,N_13162);
or U14141 (N_14141,N_12948,N_13194);
nor U14142 (N_14142,N_13550,N_13181);
nor U14143 (N_14143,N_13587,N_12880);
nand U14144 (N_14144,N_13066,N_13416);
nand U14145 (N_14145,N_13577,N_13357);
xnor U14146 (N_14146,N_13085,N_12874);
xor U14147 (N_14147,N_13319,N_13512);
and U14148 (N_14148,N_13227,N_13194);
nand U14149 (N_14149,N_12911,N_12849);
nand U14150 (N_14150,N_12822,N_13442);
xor U14151 (N_14151,N_12885,N_13302);
nor U14152 (N_14152,N_12857,N_12897);
xor U14153 (N_14153,N_13107,N_12916);
or U14154 (N_14154,N_13161,N_13246);
nor U14155 (N_14155,N_13387,N_13480);
nor U14156 (N_14156,N_13437,N_13531);
nor U14157 (N_14157,N_13016,N_13300);
and U14158 (N_14158,N_13062,N_13123);
or U14159 (N_14159,N_13035,N_13334);
and U14160 (N_14160,N_13421,N_13265);
or U14161 (N_14161,N_13175,N_13419);
nand U14162 (N_14162,N_12901,N_13159);
nand U14163 (N_14163,N_12883,N_13218);
or U14164 (N_14164,N_13318,N_13402);
nand U14165 (N_14165,N_13504,N_13310);
nand U14166 (N_14166,N_13177,N_12996);
and U14167 (N_14167,N_13326,N_13515);
nor U14168 (N_14168,N_12928,N_13477);
or U14169 (N_14169,N_13395,N_12854);
xor U14170 (N_14170,N_12951,N_13223);
nand U14171 (N_14171,N_13291,N_13320);
and U14172 (N_14172,N_13010,N_13125);
and U14173 (N_14173,N_13356,N_13581);
and U14174 (N_14174,N_13103,N_12982);
and U14175 (N_14175,N_13462,N_12824);
xnor U14176 (N_14176,N_13446,N_13171);
and U14177 (N_14177,N_12983,N_13055);
xnor U14178 (N_14178,N_13170,N_12927);
nor U14179 (N_14179,N_13077,N_12832);
nor U14180 (N_14180,N_12905,N_12893);
nor U14181 (N_14181,N_13572,N_12975);
nor U14182 (N_14182,N_12884,N_13163);
and U14183 (N_14183,N_13536,N_12959);
nand U14184 (N_14184,N_13533,N_12888);
or U14185 (N_14185,N_12990,N_13026);
nor U14186 (N_14186,N_13270,N_13021);
nor U14187 (N_14187,N_13436,N_12837);
xnor U14188 (N_14188,N_13091,N_13086);
or U14189 (N_14189,N_13572,N_12855);
and U14190 (N_14190,N_12914,N_13495);
nand U14191 (N_14191,N_12823,N_13520);
nor U14192 (N_14192,N_13556,N_12948);
nor U14193 (N_14193,N_13263,N_13209);
and U14194 (N_14194,N_13074,N_13368);
xor U14195 (N_14195,N_13581,N_12946);
xor U14196 (N_14196,N_12943,N_12915);
or U14197 (N_14197,N_12810,N_12869);
nand U14198 (N_14198,N_13509,N_13196);
nor U14199 (N_14199,N_13376,N_13185);
or U14200 (N_14200,N_13511,N_13110);
nand U14201 (N_14201,N_13592,N_13004);
and U14202 (N_14202,N_12932,N_13292);
nor U14203 (N_14203,N_13555,N_13128);
nand U14204 (N_14204,N_13281,N_13258);
or U14205 (N_14205,N_13281,N_12898);
nor U14206 (N_14206,N_13093,N_13229);
nor U14207 (N_14207,N_13015,N_13115);
xor U14208 (N_14208,N_13062,N_13498);
and U14209 (N_14209,N_13097,N_13351);
or U14210 (N_14210,N_13582,N_13236);
nand U14211 (N_14211,N_13219,N_13542);
nand U14212 (N_14212,N_13532,N_12971);
and U14213 (N_14213,N_13227,N_12962);
nand U14214 (N_14214,N_13524,N_13124);
and U14215 (N_14215,N_13447,N_13436);
and U14216 (N_14216,N_12896,N_13265);
or U14217 (N_14217,N_13299,N_13144);
nand U14218 (N_14218,N_13117,N_13100);
nand U14219 (N_14219,N_13357,N_13425);
or U14220 (N_14220,N_13141,N_13491);
nand U14221 (N_14221,N_12862,N_13166);
nor U14222 (N_14222,N_13560,N_13107);
nand U14223 (N_14223,N_13162,N_13401);
nand U14224 (N_14224,N_12852,N_12940);
and U14225 (N_14225,N_12967,N_12989);
nor U14226 (N_14226,N_13194,N_13371);
or U14227 (N_14227,N_13397,N_13006);
or U14228 (N_14228,N_12939,N_12859);
nor U14229 (N_14229,N_13468,N_13188);
xnor U14230 (N_14230,N_13165,N_13321);
or U14231 (N_14231,N_13025,N_13137);
and U14232 (N_14232,N_13104,N_13556);
xor U14233 (N_14233,N_13463,N_13255);
and U14234 (N_14234,N_13083,N_13261);
xnor U14235 (N_14235,N_13103,N_13321);
and U14236 (N_14236,N_13482,N_12901);
nand U14237 (N_14237,N_13027,N_13228);
nor U14238 (N_14238,N_13021,N_12820);
nand U14239 (N_14239,N_12812,N_13453);
nand U14240 (N_14240,N_13374,N_13585);
nand U14241 (N_14241,N_13070,N_13322);
nor U14242 (N_14242,N_13501,N_13599);
nand U14243 (N_14243,N_13491,N_13132);
and U14244 (N_14244,N_12817,N_13113);
xnor U14245 (N_14245,N_13231,N_12907);
or U14246 (N_14246,N_13059,N_12811);
or U14247 (N_14247,N_12875,N_13324);
nor U14248 (N_14248,N_13321,N_13149);
and U14249 (N_14249,N_13541,N_13063);
and U14250 (N_14250,N_12967,N_13312);
and U14251 (N_14251,N_13256,N_13546);
and U14252 (N_14252,N_13188,N_13333);
or U14253 (N_14253,N_13082,N_12878);
nand U14254 (N_14254,N_13234,N_13535);
nor U14255 (N_14255,N_13085,N_13315);
nand U14256 (N_14256,N_13248,N_13294);
and U14257 (N_14257,N_13550,N_13327);
nand U14258 (N_14258,N_13537,N_13291);
xor U14259 (N_14259,N_12991,N_13527);
nand U14260 (N_14260,N_13214,N_12864);
nor U14261 (N_14261,N_12802,N_13244);
nor U14262 (N_14262,N_12930,N_13023);
nand U14263 (N_14263,N_12810,N_12802);
and U14264 (N_14264,N_13299,N_13589);
nor U14265 (N_14265,N_13468,N_13421);
nand U14266 (N_14266,N_13357,N_13053);
nand U14267 (N_14267,N_13507,N_13554);
and U14268 (N_14268,N_12889,N_13124);
and U14269 (N_14269,N_13009,N_13343);
or U14270 (N_14270,N_13326,N_13113);
nand U14271 (N_14271,N_13227,N_13430);
or U14272 (N_14272,N_13077,N_13022);
nand U14273 (N_14273,N_13433,N_12913);
xor U14274 (N_14274,N_12817,N_13445);
and U14275 (N_14275,N_12814,N_13352);
and U14276 (N_14276,N_13362,N_13093);
xnor U14277 (N_14277,N_13086,N_13503);
nor U14278 (N_14278,N_12986,N_12896);
nand U14279 (N_14279,N_13122,N_13495);
or U14280 (N_14280,N_13373,N_13106);
or U14281 (N_14281,N_13419,N_13280);
nand U14282 (N_14282,N_12832,N_12953);
nor U14283 (N_14283,N_13547,N_13128);
or U14284 (N_14284,N_12863,N_12954);
nor U14285 (N_14285,N_13468,N_12924);
xnor U14286 (N_14286,N_13080,N_12984);
nand U14287 (N_14287,N_12927,N_13146);
xnor U14288 (N_14288,N_13018,N_13400);
nand U14289 (N_14289,N_13369,N_13514);
nand U14290 (N_14290,N_13592,N_13154);
or U14291 (N_14291,N_13394,N_13583);
nand U14292 (N_14292,N_13155,N_13337);
nand U14293 (N_14293,N_12911,N_13141);
xnor U14294 (N_14294,N_12993,N_13071);
or U14295 (N_14295,N_13091,N_13388);
xnor U14296 (N_14296,N_13226,N_12908);
nand U14297 (N_14297,N_12904,N_12839);
nand U14298 (N_14298,N_13022,N_13320);
xnor U14299 (N_14299,N_13593,N_13506);
nor U14300 (N_14300,N_12946,N_12872);
or U14301 (N_14301,N_12953,N_13457);
nand U14302 (N_14302,N_12800,N_13512);
xnor U14303 (N_14303,N_13486,N_13125);
xnor U14304 (N_14304,N_13458,N_13442);
and U14305 (N_14305,N_13349,N_13023);
nand U14306 (N_14306,N_12940,N_12976);
nand U14307 (N_14307,N_12990,N_13579);
and U14308 (N_14308,N_13405,N_13534);
nor U14309 (N_14309,N_13466,N_12816);
and U14310 (N_14310,N_13586,N_12844);
and U14311 (N_14311,N_13065,N_13165);
nand U14312 (N_14312,N_13071,N_13140);
or U14313 (N_14313,N_13385,N_13559);
and U14314 (N_14314,N_13470,N_13303);
or U14315 (N_14315,N_13357,N_13265);
or U14316 (N_14316,N_13471,N_13250);
nor U14317 (N_14317,N_13159,N_13464);
nor U14318 (N_14318,N_13409,N_12928);
and U14319 (N_14319,N_13471,N_13117);
and U14320 (N_14320,N_13578,N_13397);
xnor U14321 (N_14321,N_12927,N_13227);
nand U14322 (N_14322,N_12900,N_13225);
or U14323 (N_14323,N_13040,N_13017);
or U14324 (N_14324,N_12951,N_13504);
nor U14325 (N_14325,N_13141,N_13517);
nor U14326 (N_14326,N_13002,N_13151);
nor U14327 (N_14327,N_13512,N_13025);
nor U14328 (N_14328,N_13286,N_13349);
and U14329 (N_14329,N_12807,N_12948);
nand U14330 (N_14330,N_13466,N_13346);
or U14331 (N_14331,N_13472,N_13115);
xnor U14332 (N_14332,N_12875,N_13164);
nor U14333 (N_14333,N_13461,N_12998);
nor U14334 (N_14334,N_12856,N_12848);
nand U14335 (N_14335,N_13529,N_13566);
nor U14336 (N_14336,N_13391,N_13302);
nor U14337 (N_14337,N_12981,N_13421);
xnor U14338 (N_14338,N_13127,N_12825);
xor U14339 (N_14339,N_13290,N_13532);
xor U14340 (N_14340,N_13356,N_13264);
nand U14341 (N_14341,N_12910,N_12994);
or U14342 (N_14342,N_13496,N_13123);
or U14343 (N_14343,N_12900,N_12825);
nand U14344 (N_14344,N_12863,N_13513);
or U14345 (N_14345,N_12845,N_13500);
or U14346 (N_14346,N_13369,N_13433);
nand U14347 (N_14347,N_13488,N_12936);
nand U14348 (N_14348,N_13397,N_12991);
nand U14349 (N_14349,N_13283,N_13144);
xor U14350 (N_14350,N_12932,N_13226);
xor U14351 (N_14351,N_12816,N_13450);
xnor U14352 (N_14352,N_12963,N_13119);
or U14353 (N_14353,N_12948,N_12804);
nand U14354 (N_14354,N_13131,N_13312);
nand U14355 (N_14355,N_13405,N_12869);
xnor U14356 (N_14356,N_13530,N_13485);
or U14357 (N_14357,N_13316,N_13073);
and U14358 (N_14358,N_13258,N_12892);
nor U14359 (N_14359,N_13550,N_13575);
nand U14360 (N_14360,N_13211,N_13187);
or U14361 (N_14361,N_12833,N_13549);
nand U14362 (N_14362,N_12959,N_12848);
xnor U14363 (N_14363,N_13124,N_13028);
xor U14364 (N_14364,N_13362,N_13044);
xor U14365 (N_14365,N_13349,N_13488);
and U14366 (N_14366,N_13572,N_13171);
and U14367 (N_14367,N_13199,N_13019);
xnor U14368 (N_14368,N_12849,N_13331);
and U14369 (N_14369,N_13583,N_12810);
and U14370 (N_14370,N_13380,N_13346);
or U14371 (N_14371,N_12976,N_12887);
xor U14372 (N_14372,N_13497,N_13433);
nor U14373 (N_14373,N_13197,N_13565);
nand U14374 (N_14374,N_13494,N_13135);
nand U14375 (N_14375,N_13384,N_13477);
xnor U14376 (N_14376,N_13492,N_12904);
or U14377 (N_14377,N_12805,N_12860);
and U14378 (N_14378,N_13428,N_12945);
xor U14379 (N_14379,N_13356,N_13328);
nor U14380 (N_14380,N_13035,N_13366);
nand U14381 (N_14381,N_13072,N_13112);
nand U14382 (N_14382,N_13260,N_13176);
nor U14383 (N_14383,N_13427,N_13359);
nor U14384 (N_14384,N_13096,N_12817);
xor U14385 (N_14385,N_13384,N_13237);
or U14386 (N_14386,N_13336,N_13331);
and U14387 (N_14387,N_13379,N_13103);
nor U14388 (N_14388,N_12931,N_13533);
or U14389 (N_14389,N_13303,N_12994);
and U14390 (N_14390,N_12857,N_13272);
xor U14391 (N_14391,N_13159,N_13376);
xnor U14392 (N_14392,N_13381,N_12872);
xor U14393 (N_14393,N_13278,N_13543);
or U14394 (N_14394,N_12841,N_12804);
or U14395 (N_14395,N_12972,N_13140);
and U14396 (N_14396,N_13525,N_13224);
or U14397 (N_14397,N_13288,N_13569);
nor U14398 (N_14398,N_13264,N_13222);
and U14399 (N_14399,N_13185,N_13175);
xnor U14400 (N_14400,N_13866,N_14319);
or U14401 (N_14401,N_13835,N_14064);
xnor U14402 (N_14402,N_13873,N_13877);
nand U14403 (N_14403,N_14133,N_14134);
nor U14404 (N_14404,N_13646,N_14283);
xor U14405 (N_14405,N_13737,N_14177);
or U14406 (N_14406,N_13939,N_14334);
and U14407 (N_14407,N_14073,N_13688);
and U14408 (N_14408,N_14137,N_13639);
xor U14409 (N_14409,N_13611,N_13643);
or U14410 (N_14410,N_14171,N_13677);
and U14411 (N_14411,N_14119,N_14333);
xnor U14412 (N_14412,N_14196,N_14385);
nand U14413 (N_14413,N_13744,N_13924);
nand U14414 (N_14414,N_14352,N_13789);
and U14415 (N_14415,N_13684,N_13862);
or U14416 (N_14416,N_14114,N_14041);
or U14417 (N_14417,N_14144,N_13809);
and U14418 (N_14418,N_14237,N_13794);
xnor U14419 (N_14419,N_13977,N_13651);
nand U14420 (N_14420,N_13991,N_14243);
nand U14421 (N_14421,N_14005,N_13722);
nor U14422 (N_14422,N_14354,N_14106);
nand U14423 (N_14423,N_14088,N_13997);
and U14424 (N_14424,N_13755,N_13878);
xor U14425 (N_14425,N_14032,N_14065);
nand U14426 (N_14426,N_14249,N_14317);
xor U14427 (N_14427,N_14301,N_13821);
and U14428 (N_14428,N_13847,N_14049);
or U14429 (N_14429,N_14351,N_13950);
and U14430 (N_14430,N_14014,N_13990);
nand U14431 (N_14431,N_13669,N_14099);
or U14432 (N_14432,N_13691,N_14257);
xor U14433 (N_14433,N_14310,N_14348);
xor U14434 (N_14434,N_14029,N_13813);
nor U14435 (N_14435,N_14213,N_14173);
nand U14436 (N_14436,N_13870,N_14080);
nand U14437 (N_14437,N_13674,N_14265);
nand U14438 (N_14438,N_14353,N_13909);
xor U14439 (N_14439,N_14185,N_14377);
or U14440 (N_14440,N_14231,N_13826);
nor U14441 (N_14441,N_14392,N_13750);
nand U14442 (N_14442,N_13682,N_13773);
xnor U14443 (N_14443,N_13978,N_13683);
and U14444 (N_14444,N_14107,N_14108);
xor U14445 (N_14445,N_14054,N_14262);
xor U14446 (N_14446,N_14274,N_14003);
xor U14447 (N_14447,N_13928,N_13786);
and U14448 (N_14448,N_13752,N_13719);
and U14449 (N_14449,N_14182,N_13687);
nor U14450 (N_14450,N_14258,N_13917);
nand U14451 (N_14451,N_13896,N_14176);
xnor U14452 (N_14452,N_14184,N_14271);
or U14453 (N_14453,N_13738,N_13717);
nor U14454 (N_14454,N_14150,N_13779);
nand U14455 (N_14455,N_14223,N_13884);
or U14456 (N_14456,N_14035,N_14021);
nand U14457 (N_14457,N_14376,N_14395);
nand U14458 (N_14458,N_14285,N_13985);
nand U14459 (N_14459,N_13706,N_13655);
and U14460 (N_14460,N_13681,N_14207);
and U14461 (N_14461,N_13972,N_14039);
xnor U14462 (N_14462,N_14228,N_13998);
nand U14463 (N_14463,N_13751,N_13652);
xor U14464 (N_14464,N_14240,N_13852);
and U14465 (N_14465,N_14360,N_14323);
xor U14466 (N_14466,N_14277,N_13937);
and U14467 (N_14467,N_13995,N_14188);
or U14468 (N_14468,N_13795,N_14076);
nand U14469 (N_14469,N_14209,N_13949);
nand U14470 (N_14470,N_13802,N_14020);
nor U14471 (N_14471,N_13665,N_14379);
nor U14472 (N_14472,N_13837,N_13758);
nand U14473 (N_14473,N_13904,N_13634);
xnor U14474 (N_14474,N_13938,N_14071);
nand U14475 (N_14475,N_14215,N_14284);
nor U14476 (N_14476,N_14342,N_13854);
xnor U14477 (N_14477,N_13858,N_14236);
nand U14478 (N_14478,N_13960,N_14357);
nor U14479 (N_14479,N_13720,N_13881);
xor U14480 (N_14480,N_13935,N_13603);
and U14481 (N_14481,N_13976,N_14368);
nand U14482 (N_14482,N_13782,N_14307);
nand U14483 (N_14483,N_13828,N_13705);
or U14484 (N_14484,N_13628,N_14104);
xor U14485 (N_14485,N_14063,N_13894);
or U14486 (N_14486,N_14186,N_14100);
xnor U14487 (N_14487,N_14110,N_14252);
or U14488 (N_14488,N_13733,N_14273);
or U14489 (N_14489,N_13983,N_14141);
nand U14490 (N_14490,N_13908,N_14127);
and U14491 (N_14491,N_14227,N_14168);
or U14492 (N_14492,N_14151,N_14335);
nor U14493 (N_14493,N_14372,N_13624);
xor U14494 (N_14494,N_14361,N_13606);
nor U14495 (N_14495,N_13732,N_13885);
xor U14496 (N_14496,N_14004,N_13996);
nor U14497 (N_14497,N_13914,N_13815);
nand U14498 (N_14498,N_14200,N_14089);
xnor U14499 (N_14499,N_13934,N_14198);
nand U14500 (N_14500,N_13820,N_13667);
xor U14501 (N_14501,N_14346,N_13848);
xor U14502 (N_14502,N_14128,N_13798);
nand U14503 (N_14503,N_13975,N_13644);
nand U14504 (N_14504,N_13658,N_14025);
nor U14505 (N_14505,N_13875,N_13863);
and U14506 (N_14506,N_14092,N_14316);
nand U14507 (N_14507,N_13657,N_14381);
nand U14508 (N_14508,N_14009,N_14396);
and U14509 (N_14509,N_13776,N_14298);
nor U14510 (N_14510,N_13855,N_13953);
nand U14511 (N_14511,N_14102,N_14072);
xnor U14512 (N_14512,N_13856,N_13636);
or U14513 (N_14513,N_13721,N_13845);
nor U14514 (N_14514,N_13696,N_14261);
or U14515 (N_14515,N_14197,N_13713);
nor U14516 (N_14516,N_14299,N_13715);
or U14517 (N_14517,N_14061,N_13754);
nand U14518 (N_14518,N_14083,N_13723);
nand U14519 (N_14519,N_14275,N_14024);
nor U14520 (N_14520,N_13936,N_13625);
nor U14521 (N_14521,N_13673,N_14218);
nor U14522 (N_14522,N_14135,N_13927);
or U14523 (N_14523,N_14362,N_14159);
and U14524 (N_14524,N_14060,N_14044);
nand U14525 (N_14525,N_13966,N_14081);
nand U14526 (N_14526,N_14205,N_14389);
nand U14527 (N_14527,N_13641,N_13796);
xor U14528 (N_14528,N_14382,N_13906);
nor U14529 (N_14529,N_13648,N_14355);
and U14530 (N_14530,N_14272,N_14253);
nand U14531 (N_14531,N_13618,N_13818);
nand U14532 (N_14532,N_14096,N_14047);
or U14533 (N_14533,N_14082,N_13695);
and U14534 (N_14534,N_13843,N_14331);
nor U14535 (N_14535,N_14328,N_13942);
xor U14536 (N_14536,N_13635,N_13853);
nand U14537 (N_14537,N_14312,N_13808);
nor U14538 (N_14538,N_13787,N_14219);
and U14539 (N_14539,N_13613,N_14350);
and U14540 (N_14540,N_14022,N_14152);
nor U14541 (N_14541,N_13816,N_13701);
nand U14542 (N_14542,N_13697,N_13740);
nand U14543 (N_14543,N_13882,N_13822);
or U14544 (N_14544,N_14117,N_13790);
and U14545 (N_14545,N_14214,N_13982);
nand U14546 (N_14546,N_14130,N_14378);
xnor U14547 (N_14547,N_13708,N_14387);
or U14548 (N_14548,N_14212,N_13788);
or U14549 (N_14549,N_14181,N_13860);
or U14550 (N_14550,N_13833,N_13910);
and U14551 (N_14551,N_14220,N_14279);
and U14552 (N_14552,N_14070,N_14023);
or U14553 (N_14553,N_13670,N_14393);
xnor U14554 (N_14554,N_14129,N_14146);
nand U14555 (N_14555,N_14260,N_14246);
or U14556 (N_14556,N_13785,N_14050);
nand U14557 (N_14557,N_13830,N_13619);
or U14558 (N_14558,N_14305,N_14345);
or U14559 (N_14559,N_14148,N_14195);
and U14560 (N_14560,N_13711,N_13944);
nand U14561 (N_14561,N_14291,N_13955);
or U14562 (N_14562,N_14040,N_13887);
and U14563 (N_14563,N_13956,N_14097);
nand U14564 (N_14564,N_14391,N_13913);
or U14565 (N_14565,N_13760,N_13897);
or U14566 (N_14566,N_13609,N_14031);
nor U14567 (N_14567,N_13659,N_14235);
or U14568 (N_14568,N_14225,N_13844);
xor U14569 (N_14569,N_14363,N_13879);
or U14570 (N_14570,N_14303,N_13849);
or U14571 (N_14571,N_13840,N_14203);
xor U14572 (N_14572,N_14158,N_14139);
or U14573 (N_14573,N_14090,N_14086);
nand U14574 (N_14574,N_14125,N_14233);
nand U14575 (N_14575,N_14098,N_13948);
and U14576 (N_14576,N_14344,N_14375);
nor U14577 (N_14577,N_14057,N_13645);
or U14578 (N_14578,N_14264,N_14247);
nor U14579 (N_14579,N_13861,N_13797);
nand U14580 (N_14580,N_13661,N_13959);
nand U14581 (N_14581,N_14068,N_14315);
nor U14582 (N_14582,N_13640,N_13889);
nand U14583 (N_14583,N_13685,N_13911);
xor U14584 (N_14584,N_14033,N_13679);
and U14585 (N_14585,N_13805,N_13838);
or U14586 (N_14586,N_14145,N_13704);
and U14587 (N_14587,N_13756,N_13698);
nand U14588 (N_14588,N_13608,N_14314);
or U14589 (N_14589,N_13933,N_14101);
or U14590 (N_14590,N_14138,N_13841);
nor U14591 (N_14591,N_13890,N_13918);
and U14592 (N_14592,N_13872,N_13689);
nand U14593 (N_14593,N_13614,N_14142);
nor U14594 (N_14594,N_13999,N_14380);
or U14595 (N_14595,N_14045,N_13626);
and U14596 (N_14596,N_13926,N_13675);
nand U14597 (N_14597,N_14322,N_13662);
nor U14598 (N_14598,N_14241,N_13987);
and U14599 (N_14599,N_14111,N_13943);
or U14600 (N_14600,N_13731,N_13857);
nand U14601 (N_14601,N_14122,N_14294);
nor U14602 (N_14602,N_13989,N_13791);
xnor U14603 (N_14603,N_14201,N_14276);
nor U14604 (N_14604,N_13690,N_14311);
or U14605 (N_14605,N_13746,N_14232);
or U14606 (N_14606,N_14077,N_13869);
or U14607 (N_14607,N_14154,N_13768);
nor U14608 (N_14608,N_14297,N_13814);
and U14609 (N_14609,N_14131,N_14170);
and U14610 (N_14610,N_14229,N_14193);
or U14611 (N_14611,N_13629,N_13678);
and U14612 (N_14612,N_14079,N_14055);
nand U14613 (N_14613,N_13647,N_14325);
and U14614 (N_14614,N_14046,N_13880);
nand U14615 (N_14615,N_14339,N_13851);
nand U14616 (N_14616,N_13901,N_13601);
xnor U14617 (N_14617,N_13770,N_13792);
or U14618 (N_14618,N_14194,N_13783);
or U14619 (N_14619,N_14290,N_13620);
and U14620 (N_14620,N_14058,N_14292);
or U14621 (N_14621,N_14118,N_13915);
nor U14622 (N_14622,N_13902,N_13734);
nor U14623 (N_14623,N_14069,N_13958);
and U14624 (N_14624,N_13693,N_13931);
xnor U14625 (N_14625,N_13699,N_14308);
and U14626 (N_14626,N_14282,N_14289);
or U14627 (N_14627,N_14051,N_13947);
and U14628 (N_14628,N_14109,N_13672);
or U14629 (N_14629,N_14084,N_14062);
or U14630 (N_14630,N_13799,N_13607);
xor U14631 (N_14631,N_13850,N_14397);
and U14632 (N_14632,N_13812,N_13747);
or U14633 (N_14633,N_13718,N_13759);
and U14634 (N_14634,N_13874,N_14187);
xor U14635 (N_14635,N_13605,N_13804);
nand U14636 (N_14636,N_13832,N_13839);
and U14637 (N_14637,N_14037,N_14105);
nor U14638 (N_14638,N_13656,N_13970);
nand U14639 (N_14639,N_13666,N_14006);
or U14640 (N_14640,N_14116,N_14390);
and U14641 (N_14641,N_13604,N_14075);
nand U14642 (N_14642,N_13771,N_14126);
xnor U14643 (N_14643,N_13967,N_13980);
or U14644 (N_14644,N_14293,N_13765);
or U14645 (N_14645,N_13781,N_13710);
nand U14646 (N_14646,N_13957,N_14269);
and U14647 (N_14647,N_14002,N_14113);
and U14648 (N_14648,N_13649,N_14162);
xnor U14649 (N_14649,N_13981,N_14026);
xor U14650 (N_14650,N_13653,N_13676);
nor U14651 (N_14651,N_13663,N_14036);
xor U14652 (N_14652,N_13994,N_14165);
or U14653 (N_14653,N_13757,N_14222);
nor U14654 (N_14654,N_14038,N_13753);
and U14655 (N_14655,N_13846,N_13964);
or U14656 (N_14656,N_13775,N_14224);
or U14657 (N_14657,N_13993,N_13630);
xnor U14658 (N_14658,N_13824,N_13724);
and U14659 (N_14659,N_14366,N_14093);
nor U14660 (N_14660,N_13617,N_14370);
nor U14661 (N_14661,N_13974,N_13986);
nand U14662 (N_14662,N_13600,N_14123);
nor U14663 (N_14663,N_13965,N_14164);
and U14664 (N_14664,N_14163,N_13712);
or U14665 (N_14665,N_13725,N_14302);
or U14666 (N_14666,N_13660,N_14210);
xnor U14667 (N_14667,N_14327,N_13622);
xor U14668 (N_14668,N_13899,N_14191);
and U14669 (N_14669,N_13859,N_13612);
xor U14670 (N_14670,N_13766,N_13883);
or U14671 (N_14671,N_13616,N_14178);
nand U14672 (N_14672,N_14248,N_13803);
nor U14673 (N_14673,N_14027,N_14156);
nand U14674 (N_14674,N_14018,N_13893);
nand U14675 (N_14675,N_13726,N_14115);
xnor U14676 (N_14676,N_14221,N_14140);
or U14677 (N_14677,N_14367,N_13664);
nand U14678 (N_14678,N_13971,N_13778);
xnor U14679 (N_14679,N_13735,N_13898);
and U14680 (N_14680,N_14371,N_13727);
nand U14681 (N_14681,N_14239,N_14216);
or U14682 (N_14682,N_14365,N_14028);
or U14683 (N_14683,N_14016,N_13992);
or U14684 (N_14684,N_14034,N_14288);
nand U14685 (N_14685,N_13919,N_14008);
xnor U14686 (N_14686,N_13864,N_13702);
xnor U14687 (N_14687,N_14043,N_14091);
xnor U14688 (N_14688,N_13736,N_14208);
and U14689 (N_14689,N_13749,N_14394);
nor U14690 (N_14690,N_13742,N_13984);
or U14691 (N_14691,N_14112,N_13627);
nor U14692 (N_14692,N_14374,N_14256);
nand U14693 (N_14693,N_14384,N_14007);
and U14694 (N_14694,N_13793,N_13784);
nand U14695 (N_14695,N_13829,N_14373);
nor U14696 (N_14696,N_14226,N_14217);
nand U14697 (N_14697,N_14179,N_14242);
or U14698 (N_14698,N_14296,N_14001);
nor U14699 (N_14699,N_14267,N_13900);
or U14700 (N_14700,N_14358,N_13767);
or U14701 (N_14701,N_13806,N_14048);
nor U14702 (N_14702,N_13707,N_13637);
nand U14703 (N_14703,N_14143,N_13623);
xnor U14704 (N_14704,N_13969,N_14341);
or U14705 (N_14705,N_13741,N_14304);
or U14706 (N_14706,N_13774,N_14052);
nor U14707 (N_14707,N_13811,N_14281);
nand U14708 (N_14708,N_14244,N_13729);
and U14709 (N_14709,N_13642,N_14155);
nor U14710 (N_14710,N_14320,N_13867);
nor U14711 (N_14711,N_13876,N_13945);
xnor U14712 (N_14712,N_13777,N_13823);
nor U14713 (N_14713,N_13946,N_13920);
or U14714 (N_14714,N_14019,N_13951);
nor U14715 (N_14715,N_14012,N_14309);
xor U14716 (N_14716,N_13800,N_14347);
nand U14717 (N_14717,N_14103,N_14192);
or U14718 (N_14718,N_13961,N_14202);
nand U14719 (N_14719,N_13772,N_13871);
or U14720 (N_14720,N_14337,N_14078);
or U14721 (N_14721,N_14017,N_14167);
nand U14722 (N_14722,N_14153,N_14147);
and U14723 (N_14723,N_13739,N_13761);
nand U14724 (N_14724,N_13610,N_14332);
and U14725 (N_14725,N_14356,N_13745);
or U14726 (N_14726,N_14399,N_14330);
nand U14727 (N_14727,N_13615,N_14259);
nor U14728 (N_14728,N_14169,N_13892);
and U14729 (N_14729,N_14204,N_13671);
nand U14730 (N_14730,N_13932,N_14053);
xor U14731 (N_14731,N_13668,N_13905);
nand U14732 (N_14732,N_14326,N_14295);
nand U14733 (N_14733,N_14287,N_13602);
or U14734 (N_14734,N_13728,N_13836);
xor U14735 (N_14735,N_13633,N_14199);
nor U14736 (N_14736,N_14183,N_14254);
and U14737 (N_14737,N_14336,N_14306);
and U14738 (N_14738,N_13891,N_13952);
nor U14739 (N_14739,N_14270,N_13963);
and U14740 (N_14740,N_14056,N_14059);
xnor U14741 (N_14741,N_14388,N_14338);
nand U14742 (N_14742,N_14120,N_13930);
xnor U14743 (N_14743,N_13621,N_13631);
or U14744 (N_14744,N_13940,N_14364);
or U14745 (N_14745,N_13780,N_13810);
and U14746 (N_14746,N_14015,N_14250);
nand U14747 (N_14747,N_14010,N_13831);
xnor U14748 (N_14748,N_13886,N_14085);
nand U14749 (N_14749,N_13834,N_14074);
nor U14750 (N_14750,N_13686,N_13923);
xor U14751 (N_14751,N_14398,N_14013);
and U14752 (N_14752,N_13888,N_13954);
nor U14753 (N_14753,N_14180,N_14174);
nor U14754 (N_14754,N_13916,N_13716);
nor U14755 (N_14755,N_14166,N_13807);
and U14756 (N_14756,N_14087,N_14268);
and U14757 (N_14757,N_14030,N_14280);
and U14758 (N_14758,N_13842,N_13692);
xor U14759 (N_14759,N_14318,N_13764);
nor U14760 (N_14760,N_13865,N_13769);
nor U14761 (N_14761,N_13748,N_14245);
and U14762 (N_14762,N_14000,N_13925);
or U14763 (N_14763,N_14324,N_14313);
or U14764 (N_14764,N_13801,N_14095);
and U14765 (N_14765,N_13912,N_13962);
nand U14766 (N_14766,N_13650,N_14161);
nor U14767 (N_14767,N_14343,N_14121);
and U14768 (N_14768,N_14251,N_14160);
or U14769 (N_14769,N_14149,N_14266);
nor U14770 (N_14770,N_13654,N_14190);
or U14771 (N_14771,N_13680,N_13694);
or U14772 (N_14772,N_13929,N_14132);
nand U14773 (N_14773,N_14386,N_13632);
or U14774 (N_14774,N_14211,N_14255);
nor U14775 (N_14775,N_14157,N_13968);
and U14776 (N_14776,N_13827,N_14011);
xor U14777 (N_14777,N_14136,N_14340);
nor U14778 (N_14778,N_13895,N_14124);
or U14779 (N_14779,N_13743,N_13922);
xor U14780 (N_14780,N_13921,N_14238);
nand U14781 (N_14781,N_13941,N_13700);
nor U14782 (N_14782,N_13638,N_13763);
and U14783 (N_14783,N_13988,N_14383);
xor U14784 (N_14784,N_13714,N_13819);
nor U14785 (N_14785,N_14329,N_14094);
nor U14786 (N_14786,N_13703,N_14286);
nor U14787 (N_14787,N_13973,N_14066);
or U14788 (N_14788,N_14067,N_13730);
and U14789 (N_14789,N_14189,N_13979);
or U14790 (N_14790,N_14042,N_13868);
or U14791 (N_14791,N_14278,N_14172);
and U14792 (N_14792,N_13903,N_14300);
xnor U14793 (N_14793,N_14359,N_14349);
or U14794 (N_14794,N_14234,N_14230);
nand U14795 (N_14795,N_14206,N_13762);
nor U14796 (N_14796,N_13709,N_14263);
xnor U14797 (N_14797,N_14369,N_13825);
and U14798 (N_14798,N_13907,N_14175);
and U14799 (N_14799,N_14321,N_13817);
nor U14800 (N_14800,N_13984,N_14266);
nand U14801 (N_14801,N_14149,N_14273);
and U14802 (N_14802,N_13663,N_14191);
nor U14803 (N_14803,N_14134,N_14103);
xor U14804 (N_14804,N_13882,N_14127);
nand U14805 (N_14805,N_14213,N_14372);
nor U14806 (N_14806,N_14105,N_14119);
and U14807 (N_14807,N_14203,N_14068);
and U14808 (N_14808,N_13640,N_14040);
nand U14809 (N_14809,N_14115,N_14250);
xnor U14810 (N_14810,N_13892,N_13740);
nand U14811 (N_14811,N_13689,N_13828);
or U14812 (N_14812,N_14123,N_14260);
or U14813 (N_14813,N_14032,N_13930);
xor U14814 (N_14814,N_14270,N_14100);
nor U14815 (N_14815,N_14251,N_14077);
and U14816 (N_14816,N_14316,N_13975);
or U14817 (N_14817,N_13694,N_13700);
nor U14818 (N_14818,N_14204,N_14371);
nand U14819 (N_14819,N_13648,N_13604);
xor U14820 (N_14820,N_13908,N_13614);
or U14821 (N_14821,N_13618,N_13785);
nor U14822 (N_14822,N_13759,N_13659);
and U14823 (N_14823,N_13614,N_14299);
nor U14824 (N_14824,N_13923,N_13600);
nand U14825 (N_14825,N_14205,N_14322);
nor U14826 (N_14826,N_14367,N_13655);
and U14827 (N_14827,N_14036,N_13803);
xor U14828 (N_14828,N_14231,N_14084);
nand U14829 (N_14829,N_13901,N_14296);
nand U14830 (N_14830,N_14021,N_13920);
xnor U14831 (N_14831,N_13759,N_14034);
xnor U14832 (N_14832,N_13619,N_14014);
and U14833 (N_14833,N_13832,N_14038);
xor U14834 (N_14834,N_13922,N_13868);
xnor U14835 (N_14835,N_13962,N_14012);
xnor U14836 (N_14836,N_14144,N_14222);
nand U14837 (N_14837,N_14359,N_14322);
or U14838 (N_14838,N_14380,N_13653);
nor U14839 (N_14839,N_13627,N_14255);
and U14840 (N_14840,N_13609,N_13898);
and U14841 (N_14841,N_13677,N_13929);
and U14842 (N_14842,N_13745,N_14307);
nand U14843 (N_14843,N_13697,N_14046);
and U14844 (N_14844,N_13602,N_13848);
or U14845 (N_14845,N_13667,N_14133);
nor U14846 (N_14846,N_13958,N_14174);
xnor U14847 (N_14847,N_13810,N_14075);
xnor U14848 (N_14848,N_13729,N_13605);
nand U14849 (N_14849,N_14095,N_13854);
and U14850 (N_14850,N_14050,N_13921);
xnor U14851 (N_14851,N_14042,N_14158);
and U14852 (N_14852,N_14113,N_13804);
nand U14853 (N_14853,N_14008,N_13656);
or U14854 (N_14854,N_14225,N_14152);
nor U14855 (N_14855,N_14242,N_13843);
xnor U14856 (N_14856,N_14304,N_14158);
nand U14857 (N_14857,N_14182,N_13998);
and U14858 (N_14858,N_14256,N_14161);
xor U14859 (N_14859,N_14044,N_14190);
or U14860 (N_14860,N_13975,N_13984);
nor U14861 (N_14861,N_14181,N_14193);
nor U14862 (N_14862,N_14264,N_14025);
nand U14863 (N_14863,N_13844,N_13714);
and U14864 (N_14864,N_13813,N_13863);
and U14865 (N_14865,N_13930,N_14123);
or U14866 (N_14866,N_13729,N_14341);
and U14867 (N_14867,N_14259,N_14269);
and U14868 (N_14868,N_13664,N_14288);
and U14869 (N_14869,N_14046,N_13614);
or U14870 (N_14870,N_13628,N_14049);
and U14871 (N_14871,N_14236,N_14201);
xnor U14872 (N_14872,N_13884,N_13747);
or U14873 (N_14873,N_14309,N_14028);
and U14874 (N_14874,N_13659,N_14327);
nand U14875 (N_14875,N_13654,N_13839);
and U14876 (N_14876,N_14083,N_13810);
or U14877 (N_14877,N_13996,N_13784);
xnor U14878 (N_14878,N_14039,N_13853);
nand U14879 (N_14879,N_14160,N_14313);
nand U14880 (N_14880,N_14372,N_14203);
xnor U14881 (N_14881,N_13892,N_14377);
or U14882 (N_14882,N_13657,N_14097);
xor U14883 (N_14883,N_13692,N_13709);
nand U14884 (N_14884,N_13603,N_13909);
nand U14885 (N_14885,N_13978,N_14194);
nor U14886 (N_14886,N_13773,N_13713);
nor U14887 (N_14887,N_13968,N_13915);
nand U14888 (N_14888,N_13938,N_13871);
nor U14889 (N_14889,N_14001,N_14346);
nand U14890 (N_14890,N_14075,N_13638);
nand U14891 (N_14891,N_14240,N_14014);
nand U14892 (N_14892,N_14268,N_13968);
xnor U14893 (N_14893,N_13882,N_14148);
or U14894 (N_14894,N_14035,N_14258);
xnor U14895 (N_14895,N_13752,N_13896);
xnor U14896 (N_14896,N_13675,N_13787);
nor U14897 (N_14897,N_14247,N_14307);
or U14898 (N_14898,N_14218,N_13921);
nor U14899 (N_14899,N_14389,N_13838);
and U14900 (N_14900,N_13914,N_13946);
or U14901 (N_14901,N_14134,N_14258);
or U14902 (N_14902,N_14337,N_14039);
nor U14903 (N_14903,N_14206,N_13857);
and U14904 (N_14904,N_14195,N_13843);
xnor U14905 (N_14905,N_14256,N_13768);
and U14906 (N_14906,N_14107,N_14367);
xnor U14907 (N_14907,N_14263,N_14063);
and U14908 (N_14908,N_13801,N_13903);
nand U14909 (N_14909,N_14022,N_13936);
nand U14910 (N_14910,N_13864,N_13752);
or U14911 (N_14911,N_14268,N_14322);
nand U14912 (N_14912,N_14197,N_13926);
nand U14913 (N_14913,N_13952,N_14319);
nor U14914 (N_14914,N_13940,N_13821);
nand U14915 (N_14915,N_13923,N_14213);
and U14916 (N_14916,N_14141,N_13653);
or U14917 (N_14917,N_14166,N_14332);
nand U14918 (N_14918,N_13630,N_14296);
xor U14919 (N_14919,N_14028,N_14109);
nand U14920 (N_14920,N_13964,N_13700);
and U14921 (N_14921,N_14266,N_14175);
or U14922 (N_14922,N_14277,N_13792);
xnor U14923 (N_14923,N_13822,N_14186);
nor U14924 (N_14924,N_14382,N_13629);
or U14925 (N_14925,N_14375,N_14332);
xor U14926 (N_14926,N_13834,N_13666);
and U14927 (N_14927,N_13737,N_14366);
xor U14928 (N_14928,N_14242,N_13906);
nor U14929 (N_14929,N_13777,N_13645);
or U14930 (N_14930,N_14199,N_14291);
or U14931 (N_14931,N_13888,N_14240);
or U14932 (N_14932,N_13710,N_14202);
xor U14933 (N_14933,N_14243,N_13714);
or U14934 (N_14934,N_13809,N_13971);
or U14935 (N_14935,N_14266,N_14287);
or U14936 (N_14936,N_14378,N_14153);
and U14937 (N_14937,N_14046,N_14026);
nor U14938 (N_14938,N_14019,N_13904);
or U14939 (N_14939,N_13666,N_13820);
nor U14940 (N_14940,N_13972,N_14257);
and U14941 (N_14941,N_14389,N_13855);
nand U14942 (N_14942,N_14147,N_14161);
nand U14943 (N_14943,N_14143,N_14197);
nand U14944 (N_14944,N_13807,N_13995);
nand U14945 (N_14945,N_13632,N_13770);
and U14946 (N_14946,N_14138,N_14071);
nor U14947 (N_14947,N_14259,N_13680);
or U14948 (N_14948,N_13830,N_14311);
or U14949 (N_14949,N_14205,N_14118);
nand U14950 (N_14950,N_14070,N_13686);
or U14951 (N_14951,N_14121,N_14230);
and U14952 (N_14952,N_13703,N_13933);
or U14953 (N_14953,N_13990,N_13696);
nor U14954 (N_14954,N_13901,N_13680);
nand U14955 (N_14955,N_14155,N_13626);
and U14956 (N_14956,N_13630,N_13806);
or U14957 (N_14957,N_14178,N_14111);
and U14958 (N_14958,N_14116,N_13976);
nand U14959 (N_14959,N_14006,N_13978);
or U14960 (N_14960,N_14314,N_13638);
or U14961 (N_14961,N_14188,N_14159);
or U14962 (N_14962,N_14389,N_14327);
nor U14963 (N_14963,N_13889,N_14021);
nor U14964 (N_14964,N_14245,N_13613);
nand U14965 (N_14965,N_13883,N_13669);
or U14966 (N_14966,N_13765,N_13703);
or U14967 (N_14967,N_14062,N_13715);
nand U14968 (N_14968,N_13861,N_14243);
xor U14969 (N_14969,N_13727,N_13900);
and U14970 (N_14970,N_14101,N_14072);
or U14971 (N_14971,N_14334,N_13776);
and U14972 (N_14972,N_14284,N_14119);
and U14973 (N_14973,N_14287,N_14121);
or U14974 (N_14974,N_14144,N_14100);
xor U14975 (N_14975,N_14021,N_13656);
nor U14976 (N_14976,N_13907,N_14281);
nor U14977 (N_14977,N_13706,N_14207);
nand U14978 (N_14978,N_14344,N_13718);
or U14979 (N_14979,N_14190,N_13729);
or U14980 (N_14980,N_14397,N_14015);
nand U14981 (N_14981,N_13784,N_14220);
nor U14982 (N_14982,N_14179,N_13927);
nor U14983 (N_14983,N_14312,N_14160);
and U14984 (N_14984,N_14201,N_13682);
or U14985 (N_14985,N_14245,N_13721);
nor U14986 (N_14986,N_13709,N_14392);
nor U14987 (N_14987,N_14133,N_14300);
or U14988 (N_14988,N_14399,N_13705);
nand U14989 (N_14989,N_13976,N_13643);
nor U14990 (N_14990,N_13854,N_13909);
and U14991 (N_14991,N_14343,N_13912);
xor U14992 (N_14992,N_14279,N_14186);
and U14993 (N_14993,N_14007,N_14012);
xnor U14994 (N_14994,N_13699,N_14276);
and U14995 (N_14995,N_13613,N_13714);
nand U14996 (N_14996,N_14132,N_14123);
xor U14997 (N_14997,N_13685,N_13857);
xor U14998 (N_14998,N_14190,N_14176);
xor U14999 (N_14999,N_13714,N_14053);
or U15000 (N_15000,N_13621,N_13704);
and U15001 (N_15001,N_14132,N_13905);
nor U15002 (N_15002,N_14132,N_14275);
nor U15003 (N_15003,N_13809,N_14145);
or U15004 (N_15004,N_14166,N_13653);
and U15005 (N_15005,N_13871,N_13627);
nand U15006 (N_15006,N_14216,N_14286);
nor U15007 (N_15007,N_14166,N_14274);
xor U15008 (N_15008,N_14066,N_13800);
nor U15009 (N_15009,N_14177,N_13797);
xor U15010 (N_15010,N_13944,N_14059);
nor U15011 (N_15011,N_13872,N_13603);
nor U15012 (N_15012,N_14036,N_14395);
xor U15013 (N_15013,N_14011,N_14213);
nor U15014 (N_15014,N_13921,N_13830);
xnor U15015 (N_15015,N_13844,N_14354);
nor U15016 (N_15016,N_14076,N_14301);
or U15017 (N_15017,N_13890,N_14353);
and U15018 (N_15018,N_13902,N_14327);
nand U15019 (N_15019,N_14386,N_14000);
and U15020 (N_15020,N_14174,N_13799);
nor U15021 (N_15021,N_14393,N_13934);
or U15022 (N_15022,N_13837,N_14285);
and U15023 (N_15023,N_14029,N_13616);
xor U15024 (N_15024,N_13940,N_14363);
or U15025 (N_15025,N_13624,N_13985);
nand U15026 (N_15026,N_13851,N_13889);
nor U15027 (N_15027,N_13835,N_14005);
nand U15028 (N_15028,N_14052,N_13613);
xnor U15029 (N_15029,N_13623,N_13640);
xnor U15030 (N_15030,N_13912,N_13836);
and U15031 (N_15031,N_14105,N_14036);
and U15032 (N_15032,N_14379,N_14255);
or U15033 (N_15033,N_14101,N_14168);
and U15034 (N_15034,N_14166,N_14244);
or U15035 (N_15035,N_14005,N_13651);
nor U15036 (N_15036,N_14015,N_13695);
nor U15037 (N_15037,N_14035,N_14208);
nor U15038 (N_15038,N_13773,N_14159);
xnor U15039 (N_15039,N_14287,N_13739);
xnor U15040 (N_15040,N_14116,N_13715);
and U15041 (N_15041,N_14164,N_14220);
xor U15042 (N_15042,N_14013,N_13952);
xnor U15043 (N_15043,N_14154,N_14086);
nand U15044 (N_15044,N_13637,N_14153);
and U15045 (N_15045,N_13945,N_13819);
xnor U15046 (N_15046,N_13718,N_13674);
nor U15047 (N_15047,N_14141,N_14330);
and U15048 (N_15048,N_14072,N_14176);
nand U15049 (N_15049,N_13652,N_14193);
nor U15050 (N_15050,N_14373,N_13869);
or U15051 (N_15051,N_14086,N_14163);
or U15052 (N_15052,N_14222,N_14293);
xnor U15053 (N_15053,N_13771,N_13866);
nor U15054 (N_15054,N_14320,N_13834);
nor U15055 (N_15055,N_14175,N_13890);
and U15056 (N_15056,N_13963,N_13900);
xor U15057 (N_15057,N_14063,N_13839);
or U15058 (N_15058,N_13882,N_14008);
xnor U15059 (N_15059,N_13736,N_13793);
nand U15060 (N_15060,N_13690,N_13956);
or U15061 (N_15061,N_14316,N_14034);
nand U15062 (N_15062,N_14385,N_14325);
or U15063 (N_15063,N_13975,N_13631);
or U15064 (N_15064,N_14243,N_13938);
or U15065 (N_15065,N_14199,N_13739);
nor U15066 (N_15066,N_13679,N_14244);
nand U15067 (N_15067,N_13961,N_13651);
or U15068 (N_15068,N_14278,N_14271);
nand U15069 (N_15069,N_14302,N_13791);
nor U15070 (N_15070,N_14390,N_13716);
nor U15071 (N_15071,N_14374,N_13806);
nand U15072 (N_15072,N_14027,N_14385);
xnor U15073 (N_15073,N_14117,N_14337);
nor U15074 (N_15074,N_13812,N_13603);
nor U15075 (N_15075,N_13884,N_14104);
and U15076 (N_15076,N_14170,N_14055);
or U15077 (N_15077,N_14235,N_13719);
xor U15078 (N_15078,N_13792,N_13665);
and U15079 (N_15079,N_13931,N_14231);
and U15080 (N_15080,N_13742,N_13730);
nand U15081 (N_15081,N_14256,N_13798);
xor U15082 (N_15082,N_14071,N_14397);
and U15083 (N_15083,N_14293,N_14079);
and U15084 (N_15084,N_13805,N_14084);
and U15085 (N_15085,N_14220,N_14154);
nand U15086 (N_15086,N_14365,N_13819);
nor U15087 (N_15087,N_13707,N_14095);
nor U15088 (N_15088,N_13602,N_14362);
nor U15089 (N_15089,N_13763,N_13751);
and U15090 (N_15090,N_13876,N_14359);
nand U15091 (N_15091,N_14170,N_13958);
and U15092 (N_15092,N_13902,N_14171);
nor U15093 (N_15093,N_14193,N_13880);
nor U15094 (N_15094,N_13765,N_14066);
or U15095 (N_15095,N_14375,N_13862);
nor U15096 (N_15096,N_13694,N_14132);
nor U15097 (N_15097,N_14310,N_14376);
and U15098 (N_15098,N_13979,N_13930);
nor U15099 (N_15099,N_14309,N_13698);
and U15100 (N_15100,N_13939,N_14131);
nor U15101 (N_15101,N_13890,N_14388);
nand U15102 (N_15102,N_14248,N_13642);
xnor U15103 (N_15103,N_13700,N_13883);
nor U15104 (N_15104,N_14396,N_13994);
nor U15105 (N_15105,N_14175,N_13735);
or U15106 (N_15106,N_14010,N_13686);
nand U15107 (N_15107,N_13964,N_13678);
or U15108 (N_15108,N_14076,N_13693);
xnor U15109 (N_15109,N_13867,N_14269);
or U15110 (N_15110,N_13860,N_13612);
nor U15111 (N_15111,N_14352,N_14203);
or U15112 (N_15112,N_14367,N_13753);
nor U15113 (N_15113,N_13630,N_13986);
nor U15114 (N_15114,N_14119,N_14260);
nor U15115 (N_15115,N_13782,N_14015);
nor U15116 (N_15116,N_13601,N_13784);
nor U15117 (N_15117,N_13907,N_14337);
nand U15118 (N_15118,N_13603,N_14046);
or U15119 (N_15119,N_14174,N_14060);
nand U15120 (N_15120,N_13622,N_14383);
or U15121 (N_15121,N_13989,N_14388);
or U15122 (N_15122,N_13609,N_14204);
nand U15123 (N_15123,N_13803,N_14153);
nand U15124 (N_15124,N_14216,N_13921);
and U15125 (N_15125,N_13877,N_14397);
or U15126 (N_15126,N_13950,N_13767);
and U15127 (N_15127,N_13857,N_14366);
and U15128 (N_15128,N_14093,N_14189);
nor U15129 (N_15129,N_13739,N_13813);
or U15130 (N_15130,N_13969,N_13717);
or U15131 (N_15131,N_13654,N_14300);
nand U15132 (N_15132,N_14362,N_14033);
nand U15133 (N_15133,N_13962,N_13769);
nand U15134 (N_15134,N_14046,N_13763);
or U15135 (N_15135,N_14189,N_13795);
nor U15136 (N_15136,N_13755,N_13676);
nor U15137 (N_15137,N_13975,N_13608);
or U15138 (N_15138,N_14242,N_14144);
nand U15139 (N_15139,N_14303,N_14219);
xor U15140 (N_15140,N_13817,N_14229);
nand U15141 (N_15141,N_13679,N_14230);
and U15142 (N_15142,N_14001,N_13940);
or U15143 (N_15143,N_14160,N_13665);
xnor U15144 (N_15144,N_13649,N_13936);
and U15145 (N_15145,N_14287,N_14002);
or U15146 (N_15146,N_13663,N_14213);
nand U15147 (N_15147,N_14294,N_13992);
nand U15148 (N_15148,N_13864,N_13609);
nor U15149 (N_15149,N_14352,N_13902);
nand U15150 (N_15150,N_13711,N_13902);
and U15151 (N_15151,N_14084,N_14359);
and U15152 (N_15152,N_13682,N_14073);
and U15153 (N_15153,N_14316,N_14156);
and U15154 (N_15154,N_14086,N_14185);
or U15155 (N_15155,N_13922,N_13697);
nor U15156 (N_15156,N_13690,N_14134);
nand U15157 (N_15157,N_14187,N_14376);
and U15158 (N_15158,N_14003,N_14218);
nor U15159 (N_15159,N_13754,N_13949);
and U15160 (N_15160,N_14184,N_14196);
nor U15161 (N_15161,N_13982,N_14221);
nand U15162 (N_15162,N_14234,N_13726);
nor U15163 (N_15163,N_13827,N_14237);
xnor U15164 (N_15164,N_14304,N_14058);
nor U15165 (N_15165,N_13850,N_13709);
and U15166 (N_15166,N_14042,N_14348);
or U15167 (N_15167,N_13760,N_14038);
nand U15168 (N_15168,N_14149,N_13648);
xor U15169 (N_15169,N_13602,N_13768);
nand U15170 (N_15170,N_14334,N_13682);
nor U15171 (N_15171,N_13740,N_14334);
xnor U15172 (N_15172,N_14292,N_13640);
and U15173 (N_15173,N_13694,N_13856);
nand U15174 (N_15174,N_14002,N_14232);
or U15175 (N_15175,N_14085,N_14237);
xor U15176 (N_15176,N_14148,N_13669);
nand U15177 (N_15177,N_13914,N_14334);
or U15178 (N_15178,N_13932,N_14097);
and U15179 (N_15179,N_14118,N_14283);
nand U15180 (N_15180,N_14187,N_13977);
xor U15181 (N_15181,N_13628,N_13639);
and U15182 (N_15182,N_13666,N_13614);
nor U15183 (N_15183,N_13687,N_13969);
nor U15184 (N_15184,N_13918,N_14318);
nand U15185 (N_15185,N_14222,N_13994);
or U15186 (N_15186,N_14243,N_14272);
xor U15187 (N_15187,N_14115,N_13642);
nand U15188 (N_15188,N_14278,N_14205);
and U15189 (N_15189,N_14265,N_14060);
or U15190 (N_15190,N_13818,N_13826);
nor U15191 (N_15191,N_14138,N_13901);
and U15192 (N_15192,N_13990,N_13754);
and U15193 (N_15193,N_14228,N_14193);
xor U15194 (N_15194,N_13801,N_14053);
nor U15195 (N_15195,N_14332,N_13904);
or U15196 (N_15196,N_13611,N_14245);
or U15197 (N_15197,N_14146,N_14046);
and U15198 (N_15198,N_14380,N_14279);
or U15199 (N_15199,N_13816,N_14317);
nor U15200 (N_15200,N_14847,N_14613);
nor U15201 (N_15201,N_14544,N_14895);
and U15202 (N_15202,N_14804,N_14590);
and U15203 (N_15203,N_14499,N_15015);
nor U15204 (N_15204,N_14797,N_14416);
xnor U15205 (N_15205,N_14548,N_15139);
xor U15206 (N_15206,N_14795,N_14607);
nor U15207 (N_15207,N_15108,N_14939);
nand U15208 (N_15208,N_14932,N_14681);
or U15209 (N_15209,N_14423,N_14755);
nor U15210 (N_15210,N_14532,N_14641);
nand U15211 (N_15211,N_14835,N_15002);
nand U15212 (N_15212,N_14771,N_15112);
nor U15213 (N_15213,N_14820,N_14821);
nand U15214 (N_15214,N_15173,N_15022);
xor U15215 (N_15215,N_14807,N_14500);
nand U15216 (N_15216,N_14968,N_14488);
or U15217 (N_15217,N_15097,N_15012);
and U15218 (N_15218,N_14661,N_14603);
nand U15219 (N_15219,N_14749,N_14440);
nor U15220 (N_15220,N_14586,N_14974);
nor U15221 (N_15221,N_15105,N_15035);
nor U15222 (N_15222,N_14766,N_14930);
nand U15223 (N_15223,N_15116,N_14549);
nand U15224 (N_15224,N_14752,N_14600);
nor U15225 (N_15225,N_14863,N_14868);
nor U15226 (N_15226,N_14840,N_14563);
xor U15227 (N_15227,N_14450,N_15111);
nor U15228 (N_15228,N_14561,N_15059);
nor U15229 (N_15229,N_14492,N_14806);
or U15230 (N_15230,N_14478,N_14577);
or U15231 (N_15231,N_14616,N_14683);
xor U15232 (N_15232,N_14833,N_15092);
nor U15233 (N_15233,N_15102,N_14426);
and U15234 (N_15234,N_14550,N_14822);
xor U15235 (N_15235,N_14839,N_15080);
or U15236 (N_15236,N_14486,N_14865);
or U15237 (N_15237,N_15136,N_14893);
nor U15238 (N_15238,N_14668,N_15174);
nor U15239 (N_15239,N_14900,N_14575);
and U15240 (N_15240,N_14536,N_14658);
and U15241 (N_15241,N_14962,N_14652);
and U15242 (N_15242,N_15129,N_15011);
and U15243 (N_15243,N_14773,N_14653);
or U15244 (N_15244,N_15055,N_14958);
and U15245 (N_15245,N_14869,N_14497);
nor U15246 (N_15246,N_14988,N_15188);
nand U15247 (N_15247,N_14506,N_14754);
and U15248 (N_15248,N_14467,N_14911);
or U15249 (N_15249,N_14963,N_14526);
xor U15250 (N_15250,N_14543,N_14503);
xnor U15251 (N_15251,N_15017,N_14626);
nor U15252 (N_15252,N_14477,N_14717);
and U15253 (N_15253,N_15029,N_14464);
nand U15254 (N_15254,N_15166,N_14924);
nand U15255 (N_15255,N_14485,N_14579);
nand U15256 (N_15256,N_14929,N_14961);
xor U15257 (N_15257,N_14859,N_14995);
and U15258 (N_15258,N_14815,N_14636);
or U15259 (N_15259,N_15197,N_15145);
nor U15260 (N_15260,N_15077,N_14838);
xnor U15261 (N_15261,N_14711,N_14928);
nor U15262 (N_15262,N_14894,N_15070);
or U15263 (N_15263,N_15090,N_15170);
nand U15264 (N_15264,N_15052,N_15041);
and U15265 (N_15265,N_15098,N_15143);
xor U15266 (N_15266,N_14659,N_14825);
nor U15267 (N_15267,N_14511,N_14702);
or U15268 (N_15268,N_14745,N_14734);
and U15269 (N_15269,N_14850,N_14610);
nand U15270 (N_15270,N_14562,N_15156);
and U15271 (N_15271,N_15152,N_14743);
and U15272 (N_15272,N_15127,N_14912);
xor U15273 (N_15273,N_14685,N_15162);
xor U15274 (N_15274,N_15151,N_15083);
nor U15275 (N_15275,N_15199,N_14976);
nor U15276 (N_15276,N_14405,N_14713);
or U15277 (N_15277,N_14934,N_15008);
xor U15278 (N_15278,N_14760,N_15050);
xor U15279 (N_15279,N_14637,N_15118);
nand U15280 (N_15280,N_14774,N_14978);
or U15281 (N_15281,N_14722,N_15007);
or U15282 (N_15282,N_15176,N_15086);
nand U15283 (N_15283,N_14617,N_14646);
nand U15284 (N_15284,N_14400,N_15043);
xor U15285 (N_15285,N_14759,N_15138);
or U15286 (N_15286,N_14878,N_15082);
nor U15287 (N_15287,N_14629,N_14425);
nor U15288 (N_15288,N_15184,N_15177);
and U15289 (N_15289,N_15028,N_14901);
and U15290 (N_15290,N_14744,N_14857);
nand U15291 (N_15291,N_14446,N_15103);
and U15292 (N_15292,N_14468,N_14430);
nor U15293 (N_15293,N_14474,N_14566);
xnor U15294 (N_15294,N_15181,N_14622);
and U15295 (N_15295,N_15040,N_15042);
nand U15296 (N_15296,N_14625,N_14973);
xnor U15297 (N_15297,N_14747,N_15126);
xnor U15298 (N_15298,N_15065,N_15114);
xnor U15299 (N_15299,N_14966,N_14419);
nand U15300 (N_15300,N_14854,N_14777);
xor U15301 (N_15301,N_14905,N_14670);
nor U15302 (N_15302,N_14620,N_14699);
or U15303 (N_15303,N_15071,N_14953);
and U15304 (N_15304,N_14782,N_15193);
xnor U15305 (N_15305,N_15067,N_14783);
or U15306 (N_15306,N_15066,N_15119);
and U15307 (N_15307,N_14791,N_15146);
nand U15308 (N_15308,N_14509,N_15075);
nand U15309 (N_15309,N_14634,N_14411);
nand U15310 (N_15310,N_15115,N_14708);
and U15311 (N_15311,N_14612,N_15099);
nand U15312 (N_15312,N_14457,N_14580);
xor U15313 (N_15313,N_14873,N_14551);
nor U15314 (N_15314,N_14794,N_15140);
or U15315 (N_15315,N_15117,N_15198);
xnor U15316 (N_15316,N_14919,N_14843);
and U15317 (N_15317,N_14409,N_14557);
and U15318 (N_15318,N_15123,N_14648);
nor U15319 (N_15319,N_15034,N_14552);
xnor U15320 (N_15320,N_14948,N_14951);
nand U15321 (N_15321,N_14647,N_14619);
and U15322 (N_15322,N_14990,N_14437);
nor U15323 (N_15323,N_15100,N_14585);
or U15324 (N_15324,N_14584,N_14707);
xnor U15325 (N_15325,N_14882,N_14639);
nor U15326 (N_15326,N_14917,N_15125);
or U15327 (N_15327,N_14694,N_14808);
and U15328 (N_15328,N_15060,N_14864);
or U15329 (N_15329,N_14518,N_15027);
nor U15330 (N_15330,N_15026,N_14984);
nand U15331 (N_15331,N_14714,N_14650);
or U15332 (N_15332,N_14505,N_15120);
or U15333 (N_15333,N_15164,N_14877);
and U15334 (N_15334,N_14989,N_14792);
or U15335 (N_15335,N_14471,N_14898);
or U15336 (N_15336,N_14902,N_15044);
and U15337 (N_15337,N_14727,N_15049);
nor U15338 (N_15338,N_14768,N_14805);
nor U15339 (N_15339,N_14621,N_14483);
and U15340 (N_15340,N_14753,N_14906);
and U15341 (N_15341,N_15093,N_14860);
and U15342 (N_15342,N_14945,N_14655);
xor U15343 (N_15343,N_14671,N_14779);
nor U15344 (N_15344,N_14539,N_14537);
nand U15345 (N_15345,N_14632,N_15079);
or U15346 (N_15346,N_14582,N_14447);
xnor U15347 (N_15347,N_14677,N_14710);
or U15348 (N_15348,N_14516,N_14459);
and U15349 (N_15349,N_14569,N_14880);
xnor U15350 (N_15350,N_14605,N_14846);
xnor U15351 (N_15351,N_14871,N_14700);
or U15352 (N_15352,N_14684,N_15048);
xor U15353 (N_15353,N_14461,N_14431);
nor U15354 (N_15354,N_15095,N_14834);
and U15355 (N_15355,N_14523,N_15054);
and U15356 (N_15356,N_14975,N_15068);
and U15357 (N_15357,N_14925,N_15134);
and U15358 (N_15358,N_14570,N_15155);
nor U15359 (N_15359,N_14682,N_14916);
nand U15360 (N_15360,N_14842,N_15069);
xor U15361 (N_15361,N_14407,N_15063);
nand U15362 (N_15362,N_14798,N_14933);
nand U15363 (N_15363,N_15175,N_14410);
nor U15364 (N_15364,N_14444,N_14765);
and U15365 (N_15365,N_14980,N_14418);
or U15366 (N_15366,N_14730,N_15089);
and U15367 (N_15367,N_14421,N_15109);
or U15368 (N_15368,N_14855,N_14493);
nor U15369 (N_15369,N_14540,N_15169);
nor U15370 (N_15370,N_14827,N_14631);
or U15371 (N_15371,N_14908,N_14413);
nor U15372 (N_15372,N_14719,N_14504);
or U15373 (N_15373,N_14851,N_14524);
and U15374 (N_15374,N_14720,N_14718);
nand U15375 (N_15375,N_15045,N_14427);
nand U15376 (N_15376,N_14609,N_15194);
nand U15377 (N_15377,N_14952,N_14599);
or U15378 (N_15378,N_14433,N_14740);
xnor U15379 (N_15379,N_14983,N_14424);
or U15380 (N_15380,N_14943,N_14748);
or U15381 (N_15381,N_14941,N_14614);
nor U15382 (N_15382,N_14417,N_14482);
nor U15383 (N_15383,N_14695,N_14936);
nand U15384 (N_15384,N_15178,N_15073);
xnor U15385 (N_15385,N_15171,N_14964);
nor U15386 (N_15386,N_14669,N_14826);
and U15387 (N_15387,N_15147,N_14432);
nor U15388 (N_15388,N_14802,N_14615);
nor U15389 (N_15389,N_14588,N_14829);
or U15390 (N_15390,N_14831,N_14776);
nand U15391 (N_15391,N_14487,N_15160);
xor U15392 (N_15392,N_14534,N_14462);
nor U15393 (N_15393,N_14852,N_15107);
nor U15394 (N_15394,N_14618,N_14675);
xnor U15395 (N_15395,N_14491,N_14848);
or U15396 (N_15396,N_14866,N_14883);
and U15397 (N_15397,N_14856,N_14502);
or U15398 (N_15398,N_14520,N_14667);
xor U15399 (N_15399,N_14688,N_14571);
or U15400 (N_15400,N_15006,N_14602);
or U15401 (N_15401,N_15154,N_14415);
xor U15402 (N_15402,N_15031,N_14959);
nor U15403 (N_15403,N_14796,N_15110);
and U15404 (N_15404,N_14756,N_15137);
or U15405 (N_15405,N_14507,N_15039);
and U15406 (N_15406,N_14674,N_14956);
or U15407 (N_15407,N_14788,N_14531);
xnor U15408 (N_15408,N_15016,N_14456);
and U15409 (N_15409,N_14982,N_15096);
xnor U15410 (N_15410,N_14698,N_14994);
xor U15411 (N_15411,N_14598,N_14554);
xor U15412 (N_15412,N_14793,N_14750);
and U15413 (N_15413,N_14801,N_14723);
nand U15414 (N_15414,N_15158,N_15128);
xnor U15415 (N_15415,N_14741,N_15051);
nor U15416 (N_15416,N_15009,N_14998);
and U15417 (N_15417,N_14763,N_15148);
xor U15418 (N_15418,N_14960,N_14451);
or U15419 (N_15419,N_14784,N_14897);
or U15420 (N_15420,N_14828,N_14965);
nand U15421 (N_15421,N_15056,N_14676);
xor U15422 (N_15422,N_14538,N_14697);
nand U15423 (N_15423,N_14780,N_14654);
or U15424 (N_15424,N_14448,N_14672);
nand U15425 (N_15425,N_14525,N_14689);
nand U15426 (N_15426,N_14412,N_14957);
or U15427 (N_15427,N_14484,N_14886);
nor U15428 (N_15428,N_14559,N_14583);
or U15429 (N_15429,N_15150,N_14594);
or U15430 (N_15430,N_15182,N_14910);
nand U15431 (N_15431,N_14824,N_14899);
or U15432 (N_15432,N_14611,N_14515);
or U15433 (N_15433,N_14705,N_14696);
xor U15434 (N_15434,N_14977,N_14832);
xnor U15435 (N_15435,N_14633,N_14731);
nand U15436 (N_15436,N_15161,N_14439);
nor U15437 (N_15437,N_14687,N_14738);
xnor U15438 (N_15438,N_15000,N_14606);
nor U15439 (N_15439,N_14940,N_15192);
nor U15440 (N_15440,N_14885,N_14666);
and U15441 (N_15441,N_14533,N_14937);
nand U15442 (N_15442,N_14429,N_14879);
nor U15443 (N_15443,N_14589,N_14909);
nor U15444 (N_15444,N_14896,N_14830);
nand U15445 (N_15445,N_14420,N_14690);
or U15446 (N_15446,N_14887,N_14819);
nand U15447 (N_15447,N_15132,N_14403);
nor U15448 (N_15448,N_15047,N_14872);
nand U15449 (N_15449,N_14649,N_14442);
nand U15450 (N_15450,N_14874,N_15130);
and U15451 (N_15451,N_14498,N_14469);
nor U15452 (N_15452,N_14949,N_14709);
nor U15453 (N_15453,N_14761,N_14679);
nand U15454 (N_15454,N_15004,N_14913);
xnor U15455 (N_15455,N_15032,N_14642);
nor U15456 (N_15456,N_14853,N_15179);
nand U15457 (N_15457,N_15001,N_15183);
nand U15458 (N_15458,N_14657,N_15122);
or U15459 (N_15459,N_14817,N_14915);
or U15460 (N_15460,N_14422,N_15195);
xnor U15461 (N_15461,N_14903,N_14472);
xor U15462 (N_15462,N_14733,N_14428);
xnor U15463 (N_15463,N_14553,N_14522);
xor U15464 (N_15464,N_14724,N_15030);
or U15465 (N_15465,N_14568,N_14463);
nand U15466 (N_15466,N_14979,N_14596);
and U15467 (N_15467,N_14489,N_14920);
or U15468 (N_15468,N_15036,N_14786);
or U15469 (N_15469,N_14762,N_14728);
xnor U15470 (N_15470,N_14861,N_15037);
nand U15471 (N_15471,N_14567,N_14452);
nand U15472 (N_15472,N_15159,N_14862);
and U15473 (N_15473,N_14944,N_15106);
xor U15474 (N_15474,N_15020,N_15180);
xor U15475 (N_15475,N_14578,N_14758);
xnor U15476 (N_15476,N_14624,N_14816);
xnor U15477 (N_15477,N_14954,N_14673);
nand U15478 (N_15478,N_15064,N_14781);
xnor U15479 (N_15479,N_14889,N_15131);
xnor U15480 (N_15480,N_15072,N_14875);
and U15481 (N_15481,N_15010,N_14986);
or U15482 (N_15482,N_14775,N_14926);
nor U15483 (N_15483,N_14528,N_15057);
and U15484 (N_15484,N_14560,N_14595);
and U15485 (N_15485,N_15168,N_14996);
and U15486 (N_15486,N_14455,N_14541);
nand U15487 (N_15487,N_15144,N_14546);
nor U15488 (N_15488,N_15153,N_14521);
and U15489 (N_15489,N_15088,N_14927);
and U15490 (N_15490,N_14529,N_15005);
xor U15491 (N_15491,N_14814,N_14712);
nand U15492 (N_15492,N_14601,N_14985);
nand U15493 (N_15493,N_14971,N_14757);
nor U15494 (N_15494,N_14867,N_14818);
and U15495 (N_15495,N_15172,N_15046);
or U15496 (N_15496,N_15163,N_15091);
or U15497 (N_15497,N_14701,N_14969);
nor U15498 (N_15498,N_14408,N_15058);
nand U15499 (N_15499,N_14716,N_14630);
xor U15500 (N_15500,N_15121,N_14772);
nand U15501 (N_15501,N_14942,N_14458);
or U15502 (N_15502,N_14514,N_15142);
xor U15503 (N_15503,N_14907,N_14729);
or U15504 (N_15504,N_14535,N_14921);
xor U15505 (N_15505,N_14627,N_14592);
nor U15506 (N_15506,N_15024,N_14591);
and U15507 (N_15507,N_14558,N_14643);
and U15508 (N_15508,N_14555,N_14803);
nand U15509 (N_15509,N_15190,N_15094);
and U15510 (N_15510,N_14742,N_14715);
and U15511 (N_15511,N_14576,N_15013);
nor U15512 (N_15512,N_14800,N_14645);
nand U15513 (N_15513,N_14811,N_14809);
or U15514 (N_15514,N_14767,N_15165);
nand U15515 (N_15515,N_14946,N_14573);
or U15516 (N_15516,N_15133,N_14406);
xor U15517 (N_15517,N_14764,N_14787);
or U15518 (N_15518,N_14884,N_14950);
nor U15519 (N_15519,N_14736,N_14845);
nor U15520 (N_15520,N_14836,N_14680);
nand U15521 (N_15521,N_14438,N_15014);
or U15522 (N_15522,N_15196,N_15135);
and U15523 (N_15523,N_14527,N_14635);
and U15524 (N_15524,N_14545,N_15061);
nor U15525 (N_15525,N_14918,N_14693);
nand U15526 (N_15526,N_14678,N_14725);
xnor U15527 (N_15527,N_14453,N_14692);
and U15528 (N_15528,N_14512,N_14481);
nand U15529 (N_15529,N_15167,N_14993);
and U15530 (N_15530,N_14997,N_14651);
xor U15531 (N_15531,N_14475,N_14770);
or U15532 (N_15532,N_14501,N_15038);
and U15533 (N_15533,N_14991,N_14510);
nand U15534 (N_15534,N_14769,N_14849);
and U15535 (N_15535,N_14890,N_14445);
nand U15536 (N_15536,N_15021,N_14876);
nand U15537 (N_15537,N_15019,N_14914);
and U15538 (N_15538,N_14799,N_14881);
nor U15539 (N_15539,N_14608,N_14443);
xnor U15540 (N_15540,N_14746,N_14858);
xnor U15541 (N_15541,N_14970,N_14530);
nor U15542 (N_15542,N_15157,N_14479);
and U15543 (N_15543,N_14656,N_14581);
xnor U15544 (N_15544,N_14737,N_14449);
nand U15545 (N_15545,N_14542,N_14721);
xnor U15546 (N_15546,N_14992,N_15053);
nor U15547 (N_15547,N_15085,N_15074);
and U15548 (N_15548,N_14810,N_14703);
xnor U15549 (N_15549,N_14644,N_14460);
and U15550 (N_15550,N_14891,N_14789);
nor U15551 (N_15551,N_15189,N_14841);
or U15552 (N_15552,N_14434,N_15124);
and U15553 (N_15553,N_15078,N_14663);
nand U15554 (N_15554,N_14726,N_14465);
and U15555 (N_15555,N_14436,N_14935);
xor U15556 (N_15556,N_15018,N_14490);
xor U15557 (N_15557,N_14967,N_15087);
xnor U15558 (N_15558,N_14564,N_14547);
nor U15559 (N_15559,N_14414,N_14473);
and U15560 (N_15560,N_15062,N_14972);
xnor U15561 (N_15561,N_14454,N_14441);
and U15562 (N_15562,N_14470,N_14587);
and U15563 (N_15563,N_14597,N_14999);
or U15564 (N_15564,N_14593,N_14844);
nor U15565 (N_15565,N_14823,N_14638);
and U15566 (N_15566,N_14665,N_14778);
nand U15567 (N_15567,N_14495,N_14466);
nand U15568 (N_15568,N_15033,N_14660);
or U15569 (N_15569,N_14664,N_14623);
nand U15570 (N_15570,N_14888,N_14947);
nor U15571 (N_15571,N_14494,N_15191);
nor U15572 (N_15572,N_14496,N_14981);
xor U15573 (N_15573,N_15081,N_14640);
or U15574 (N_15574,N_14556,N_14691);
xor U15575 (N_15575,N_14739,N_14751);
and U15576 (N_15576,N_14785,N_14955);
or U15577 (N_15577,N_14938,N_14837);
nand U15578 (N_15578,N_14790,N_14519);
or U15579 (N_15579,N_15186,N_14480);
or U15580 (N_15580,N_14565,N_14402);
or U15581 (N_15581,N_14732,N_14735);
nand U15582 (N_15582,N_15185,N_15025);
xor U15583 (N_15583,N_15101,N_14628);
nand U15584 (N_15584,N_14574,N_14435);
nor U15585 (N_15585,N_14508,N_14476);
or U15586 (N_15586,N_14870,N_14662);
and U15587 (N_15587,N_14517,N_14572);
nand U15588 (N_15588,N_14604,N_14904);
or U15589 (N_15589,N_14987,N_15003);
nor U15590 (N_15590,N_15187,N_14812);
or U15591 (N_15591,N_15076,N_14513);
and U15592 (N_15592,N_14813,N_14923);
nor U15593 (N_15593,N_15141,N_15023);
nor U15594 (N_15594,N_14892,N_14931);
nor U15595 (N_15595,N_14401,N_14706);
nand U15596 (N_15596,N_14704,N_15084);
and U15597 (N_15597,N_14404,N_14686);
xor U15598 (N_15598,N_15149,N_15104);
xnor U15599 (N_15599,N_14922,N_15113);
nand U15600 (N_15600,N_15100,N_15077);
nand U15601 (N_15601,N_14951,N_14536);
xnor U15602 (N_15602,N_15157,N_14528);
nor U15603 (N_15603,N_15113,N_14792);
and U15604 (N_15604,N_14751,N_14418);
nand U15605 (N_15605,N_14464,N_14862);
nor U15606 (N_15606,N_15027,N_14424);
xnor U15607 (N_15607,N_14630,N_14553);
nor U15608 (N_15608,N_14748,N_14738);
xor U15609 (N_15609,N_14404,N_15112);
xor U15610 (N_15610,N_15150,N_14537);
nand U15611 (N_15611,N_14430,N_14653);
xnor U15612 (N_15612,N_14473,N_15151);
or U15613 (N_15613,N_14736,N_14687);
xor U15614 (N_15614,N_14761,N_15099);
xnor U15615 (N_15615,N_14970,N_14870);
nand U15616 (N_15616,N_14594,N_14885);
and U15617 (N_15617,N_14932,N_14836);
nand U15618 (N_15618,N_14947,N_14521);
nor U15619 (N_15619,N_14746,N_14645);
or U15620 (N_15620,N_14571,N_15170);
and U15621 (N_15621,N_14467,N_14632);
or U15622 (N_15622,N_14703,N_14525);
nor U15623 (N_15623,N_15038,N_14993);
or U15624 (N_15624,N_14918,N_14793);
or U15625 (N_15625,N_14457,N_15190);
and U15626 (N_15626,N_15179,N_14976);
nand U15627 (N_15627,N_14636,N_14637);
nor U15628 (N_15628,N_14653,N_15151);
nor U15629 (N_15629,N_14657,N_14768);
or U15630 (N_15630,N_14627,N_14848);
xor U15631 (N_15631,N_14694,N_15099);
nor U15632 (N_15632,N_15003,N_15174);
nand U15633 (N_15633,N_15098,N_14620);
or U15634 (N_15634,N_14920,N_15123);
nor U15635 (N_15635,N_14601,N_15197);
or U15636 (N_15636,N_15021,N_15156);
nand U15637 (N_15637,N_15041,N_14482);
xor U15638 (N_15638,N_14573,N_14695);
nand U15639 (N_15639,N_15110,N_15002);
xor U15640 (N_15640,N_14681,N_14478);
or U15641 (N_15641,N_14506,N_15087);
or U15642 (N_15642,N_14424,N_15136);
nand U15643 (N_15643,N_14691,N_14713);
nor U15644 (N_15644,N_14722,N_14716);
and U15645 (N_15645,N_15024,N_14764);
nand U15646 (N_15646,N_14923,N_15119);
nand U15647 (N_15647,N_14653,N_15158);
xor U15648 (N_15648,N_15196,N_15123);
nor U15649 (N_15649,N_14862,N_14951);
nand U15650 (N_15650,N_14618,N_14494);
and U15651 (N_15651,N_14789,N_14953);
or U15652 (N_15652,N_15016,N_14979);
xor U15653 (N_15653,N_14493,N_14590);
and U15654 (N_15654,N_14425,N_15186);
nor U15655 (N_15655,N_14621,N_14462);
or U15656 (N_15656,N_15030,N_14652);
nor U15657 (N_15657,N_15175,N_14878);
and U15658 (N_15658,N_15130,N_14759);
xor U15659 (N_15659,N_14786,N_14907);
nand U15660 (N_15660,N_14632,N_14866);
xor U15661 (N_15661,N_14969,N_14654);
nor U15662 (N_15662,N_14577,N_15061);
and U15663 (N_15663,N_14415,N_14544);
nor U15664 (N_15664,N_15129,N_15041);
xnor U15665 (N_15665,N_14753,N_14514);
xor U15666 (N_15666,N_14712,N_14473);
xnor U15667 (N_15667,N_14651,N_14820);
and U15668 (N_15668,N_15034,N_15117);
nor U15669 (N_15669,N_14724,N_15113);
and U15670 (N_15670,N_15036,N_14469);
or U15671 (N_15671,N_14412,N_14784);
nand U15672 (N_15672,N_14569,N_14654);
and U15673 (N_15673,N_14698,N_14565);
or U15674 (N_15674,N_15191,N_14496);
or U15675 (N_15675,N_15142,N_14724);
xnor U15676 (N_15676,N_15196,N_14616);
or U15677 (N_15677,N_15041,N_14527);
or U15678 (N_15678,N_14493,N_15141);
or U15679 (N_15679,N_14790,N_15030);
or U15680 (N_15680,N_14956,N_15105);
xor U15681 (N_15681,N_14775,N_15051);
and U15682 (N_15682,N_14422,N_15078);
nor U15683 (N_15683,N_14412,N_15084);
nand U15684 (N_15684,N_15154,N_14958);
or U15685 (N_15685,N_14671,N_14620);
and U15686 (N_15686,N_14435,N_14825);
and U15687 (N_15687,N_15196,N_15036);
and U15688 (N_15688,N_14732,N_14686);
xor U15689 (N_15689,N_15063,N_14572);
or U15690 (N_15690,N_14875,N_14884);
nor U15691 (N_15691,N_14733,N_14667);
xor U15692 (N_15692,N_14428,N_14582);
nand U15693 (N_15693,N_14535,N_14796);
nor U15694 (N_15694,N_14784,N_14872);
nor U15695 (N_15695,N_14438,N_14484);
or U15696 (N_15696,N_14776,N_14585);
and U15697 (N_15697,N_14719,N_15169);
nand U15698 (N_15698,N_14740,N_15104);
and U15699 (N_15699,N_14619,N_14815);
xor U15700 (N_15700,N_14890,N_14403);
xnor U15701 (N_15701,N_14441,N_14983);
nand U15702 (N_15702,N_15088,N_14499);
and U15703 (N_15703,N_14896,N_14978);
and U15704 (N_15704,N_14617,N_15062);
xor U15705 (N_15705,N_14527,N_14586);
and U15706 (N_15706,N_15177,N_14970);
nand U15707 (N_15707,N_14995,N_14894);
nor U15708 (N_15708,N_14901,N_14439);
or U15709 (N_15709,N_14763,N_14587);
or U15710 (N_15710,N_14472,N_14943);
and U15711 (N_15711,N_14824,N_14494);
nand U15712 (N_15712,N_14480,N_14567);
nand U15713 (N_15713,N_14728,N_14684);
nand U15714 (N_15714,N_15129,N_14510);
nor U15715 (N_15715,N_14830,N_15158);
nand U15716 (N_15716,N_14544,N_14618);
or U15717 (N_15717,N_14963,N_14722);
or U15718 (N_15718,N_14977,N_14960);
or U15719 (N_15719,N_15096,N_14423);
nor U15720 (N_15720,N_14927,N_14970);
nand U15721 (N_15721,N_14527,N_14989);
and U15722 (N_15722,N_15136,N_14533);
nand U15723 (N_15723,N_14618,N_14879);
or U15724 (N_15724,N_14768,N_14786);
and U15725 (N_15725,N_14491,N_15026);
nor U15726 (N_15726,N_14854,N_14889);
and U15727 (N_15727,N_14797,N_14501);
or U15728 (N_15728,N_14776,N_14711);
xnor U15729 (N_15729,N_15189,N_15002);
xnor U15730 (N_15730,N_15198,N_14882);
xnor U15731 (N_15731,N_15162,N_14663);
nor U15732 (N_15732,N_14518,N_14582);
xor U15733 (N_15733,N_14857,N_14442);
xnor U15734 (N_15734,N_14879,N_15196);
nor U15735 (N_15735,N_14579,N_15006);
nor U15736 (N_15736,N_14921,N_15164);
nor U15737 (N_15737,N_14512,N_14665);
nand U15738 (N_15738,N_14594,N_14535);
or U15739 (N_15739,N_14758,N_14434);
and U15740 (N_15740,N_14666,N_14453);
or U15741 (N_15741,N_14991,N_14484);
xnor U15742 (N_15742,N_14535,N_14494);
nand U15743 (N_15743,N_14746,N_15097);
nand U15744 (N_15744,N_14516,N_14923);
nor U15745 (N_15745,N_14662,N_15016);
nand U15746 (N_15746,N_15106,N_15182);
nor U15747 (N_15747,N_14561,N_14729);
and U15748 (N_15748,N_15099,N_14627);
and U15749 (N_15749,N_14504,N_15053);
xnor U15750 (N_15750,N_14782,N_14952);
nor U15751 (N_15751,N_15082,N_15009);
nand U15752 (N_15752,N_14854,N_14698);
nor U15753 (N_15753,N_15004,N_14987);
or U15754 (N_15754,N_14698,N_14595);
and U15755 (N_15755,N_14764,N_14848);
or U15756 (N_15756,N_14866,N_14767);
or U15757 (N_15757,N_14843,N_14675);
and U15758 (N_15758,N_14820,N_14879);
or U15759 (N_15759,N_14570,N_14965);
and U15760 (N_15760,N_15005,N_15058);
nand U15761 (N_15761,N_14784,N_14728);
and U15762 (N_15762,N_14839,N_14498);
and U15763 (N_15763,N_14637,N_14742);
xor U15764 (N_15764,N_14470,N_14626);
nor U15765 (N_15765,N_14904,N_14462);
and U15766 (N_15766,N_14911,N_14881);
or U15767 (N_15767,N_15050,N_14799);
xor U15768 (N_15768,N_14790,N_14737);
nor U15769 (N_15769,N_15096,N_14977);
xnor U15770 (N_15770,N_14744,N_14602);
or U15771 (N_15771,N_14605,N_14820);
or U15772 (N_15772,N_14668,N_15126);
or U15773 (N_15773,N_14570,N_15098);
or U15774 (N_15774,N_14773,N_14607);
nand U15775 (N_15775,N_14709,N_14723);
xor U15776 (N_15776,N_14752,N_14491);
xnor U15777 (N_15777,N_15088,N_14871);
xnor U15778 (N_15778,N_14400,N_14878);
xor U15779 (N_15779,N_14526,N_14973);
nor U15780 (N_15780,N_15004,N_15007);
nand U15781 (N_15781,N_14917,N_14831);
nand U15782 (N_15782,N_14517,N_14501);
nand U15783 (N_15783,N_14699,N_14916);
and U15784 (N_15784,N_15174,N_14430);
and U15785 (N_15785,N_14852,N_15105);
nand U15786 (N_15786,N_14651,N_15123);
or U15787 (N_15787,N_14848,N_14581);
nand U15788 (N_15788,N_15150,N_14706);
xnor U15789 (N_15789,N_14750,N_14505);
nand U15790 (N_15790,N_15071,N_14900);
nand U15791 (N_15791,N_14678,N_14676);
nor U15792 (N_15792,N_14667,N_14415);
xor U15793 (N_15793,N_14619,N_14930);
nor U15794 (N_15794,N_14859,N_14782);
and U15795 (N_15795,N_15125,N_14937);
and U15796 (N_15796,N_14960,N_14760);
nand U15797 (N_15797,N_14809,N_15176);
nand U15798 (N_15798,N_14561,N_14417);
or U15799 (N_15799,N_14435,N_14992);
xnor U15800 (N_15800,N_14858,N_14979);
xor U15801 (N_15801,N_14482,N_14872);
and U15802 (N_15802,N_14680,N_15032);
nand U15803 (N_15803,N_14407,N_14842);
or U15804 (N_15804,N_14742,N_14601);
nand U15805 (N_15805,N_14920,N_15071);
or U15806 (N_15806,N_14734,N_15034);
and U15807 (N_15807,N_14513,N_14992);
and U15808 (N_15808,N_14824,N_14647);
nor U15809 (N_15809,N_14585,N_14745);
xnor U15810 (N_15810,N_14624,N_14942);
nor U15811 (N_15811,N_15022,N_14662);
nand U15812 (N_15812,N_15151,N_14513);
xor U15813 (N_15813,N_15015,N_14761);
nor U15814 (N_15814,N_14919,N_14777);
or U15815 (N_15815,N_14459,N_14750);
nor U15816 (N_15816,N_14780,N_14670);
xnor U15817 (N_15817,N_14531,N_14824);
xnor U15818 (N_15818,N_14906,N_14523);
or U15819 (N_15819,N_14514,N_14846);
or U15820 (N_15820,N_14851,N_14418);
nor U15821 (N_15821,N_14756,N_14572);
xnor U15822 (N_15822,N_14918,N_15045);
nor U15823 (N_15823,N_15039,N_14855);
nand U15824 (N_15824,N_15148,N_14406);
nand U15825 (N_15825,N_14438,N_14493);
or U15826 (N_15826,N_14870,N_14592);
or U15827 (N_15827,N_14845,N_14541);
xor U15828 (N_15828,N_14413,N_15045);
and U15829 (N_15829,N_14562,N_14449);
or U15830 (N_15830,N_14489,N_14455);
nand U15831 (N_15831,N_14870,N_15070);
or U15832 (N_15832,N_14946,N_14462);
nand U15833 (N_15833,N_14843,N_14748);
or U15834 (N_15834,N_15086,N_14749);
and U15835 (N_15835,N_14760,N_14608);
nor U15836 (N_15836,N_14586,N_15051);
nand U15837 (N_15837,N_15118,N_14880);
nor U15838 (N_15838,N_14886,N_14493);
or U15839 (N_15839,N_14433,N_14880);
nor U15840 (N_15840,N_15101,N_14686);
nand U15841 (N_15841,N_14495,N_14507);
nor U15842 (N_15842,N_14772,N_15104);
nand U15843 (N_15843,N_14500,N_14576);
xnor U15844 (N_15844,N_14422,N_14785);
and U15845 (N_15845,N_14508,N_15191);
nor U15846 (N_15846,N_14902,N_14423);
or U15847 (N_15847,N_14700,N_14932);
and U15848 (N_15848,N_15072,N_14741);
or U15849 (N_15849,N_14422,N_14973);
and U15850 (N_15850,N_14442,N_14847);
nand U15851 (N_15851,N_15034,N_14692);
xor U15852 (N_15852,N_15112,N_15080);
nand U15853 (N_15853,N_15017,N_15154);
nor U15854 (N_15854,N_14791,N_15079);
nor U15855 (N_15855,N_15150,N_15130);
nand U15856 (N_15856,N_14562,N_14740);
and U15857 (N_15857,N_14498,N_15144);
nor U15858 (N_15858,N_14593,N_14972);
or U15859 (N_15859,N_14717,N_14484);
and U15860 (N_15860,N_15092,N_15035);
xnor U15861 (N_15861,N_15070,N_14903);
and U15862 (N_15862,N_14504,N_14654);
nor U15863 (N_15863,N_15174,N_14408);
xnor U15864 (N_15864,N_14405,N_15086);
or U15865 (N_15865,N_14594,N_14581);
and U15866 (N_15866,N_14933,N_15191);
and U15867 (N_15867,N_14668,N_14860);
nand U15868 (N_15868,N_14649,N_14636);
nand U15869 (N_15869,N_14881,N_15142);
nand U15870 (N_15870,N_14718,N_14839);
and U15871 (N_15871,N_14857,N_15076);
nor U15872 (N_15872,N_14440,N_14831);
xor U15873 (N_15873,N_14960,N_14970);
or U15874 (N_15874,N_15147,N_14420);
and U15875 (N_15875,N_14617,N_14588);
or U15876 (N_15876,N_14874,N_15049);
nor U15877 (N_15877,N_14521,N_14801);
or U15878 (N_15878,N_14869,N_14685);
xnor U15879 (N_15879,N_14796,N_15037);
and U15880 (N_15880,N_14608,N_14877);
xor U15881 (N_15881,N_15004,N_14782);
xnor U15882 (N_15882,N_15063,N_14603);
and U15883 (N_15883,N_14640,N_14694);
nand U15884 (N_15884,N_14861,N_15157);
and U15885 (N_15885,N_14569,N_14784);
and U15886 (N_15886,N_14618,N_14807);
nand U15887 (N_15887,N_14840,N_14905);
nand U15888 (N_15888,N_14529,N_14856);
or U15889 (N_15889,N_14839,N_14663);
or U15890 (N_15890,N_15043,N_14749);
and U15891 (N_15891,N_15111,N_14795);
and U15892 (N_15892,N_15153,N_15063);
or U15893 (N_15893,N_14889,N_14751);
nand U15894 (N_15894,N_14969,N_14937);
and U15895 (N_15895,N_15094,N_14547);
or U15896 (N_15896,N_14937,N_14964);
or U15897 (N_15897,N_15095,N_14880);
xor U15898 (N_15898,N_14772,N_14808);
nand U15899 (N_15899,N_14844,N_14726);
nand U15900 (N_15900,N_15132,N_15191);
and U15901 (N_15901,N_14977,N_14490);
and U15902 (N_15902,N_14959,N_14781);
nor U15903 (N_15903,N_14865,N_14881);
or U15904 (N_15904,N_14714,N_15124);
and U15905 (N_15905,N_15075,N_14891);
and U15906 (N_15906,N_14633,N_14850);
nor U15907 (N_15907,N_14817,N_14477);
and U15908 (N_15908,N_14753,N_15188);
and U15909 (N_15909,N_14910,N_14565);
and U15910 (N_15910,N_14436,N_14467);
nand U15911 (N_15911,N_14487,N_14879);
nor U15912 (N_15912,N_15078,N_14836);
xnor U15913 (N_15913,N_15089,N_14882);
nand U15914 (N_15914,N_15076,N_14538);
xnor U15915 (N_15915,N_15126,N_14657);
nor U15916 (N_15916,N_15195,N_14908);
or U15917 (N_15917,N_15077,N_15184);
or U15918 (N_15918,N_15045,N_14403);
nor U15919 (N_15919,N_14811,N_14719);
nor U15920 (N_15920,N_15124,N_14646);
xnor U15921 (N_15921,N_14598,N_14582);
xor U15922 (N_15922,N_14446,N_14440);
xor U15923 (N_15923,N_14496,N_14652);
or U15924 (N_15924,N_14837,N_14511);
nor U15925 (N_15925,N_14863,N_15174);
xor U15926 (N_15926,N_15135,N_14610);
xor U15927 (N_15927,N_14937,N_14755);
or U15928 (N_15928,N_14917,N_14926);
nor U15929 (N_15929,N_14971,N_15166);
and U15930 (N_15930,N_14798,N_14550);
nor U15931 (N_15931,N_14960,N_14408);
nor U15932 (N_15932,N_14916,N_14461);
xnor U15933 (N_15933,N_15056,N_14407);
xor U15934 (N_15934,N_14648,N_14405);
or U15935 (N_15935,N_14899,N_14660);
nor U15936 (N_15936,N_15087,N_14653);
nor U15937 (N_15937,N_15199,N_14596);
and U15938 (N_15938,N_14873,N_15169);
and U15939 (N_15939,N_14852,N_14814);
or U15940 (N_15940,N_15019,N_15149);
nor U15941 (N_15941,N_14419,N_15078);
or U15942 (N_15942,N_15115,N_15162);
or U15943 (N_15943,N_14623,N_14699);
nor U15944 (N_15944,N_14808,N_14437);
xnor U15945 (N_15945,N_15067,N_14494);
and U15946 (N_15946,N_14866,N_14872);
nand U15947 (N_15947,N_15166,N_14440);
xor U15948 (N_15948,N_14526,N_14577);
nand U15949 (N_15949,N_15045,N_15178);
nand U15950 (N_15950,N_15101,N_14561);
or U15951 (N_15951,N_14724,N_14774);
xnor U15952 (N_15952,N_14588,N_14789);
or U15953 (N_15953,N_15002,N_14537);
or U15954 (N_15954,N_15042,N_14733);
xor U15955 (N_15955,N_14721,N_15005);
xor U15956 (N_15956,N_14597,N_15122);
or U15957 (N_15957,N_14930,N_14651);
nor U15958 (N_15958,N_14621,N_14777);
and U15959 (N_15959,N_14477,N_14966);
or U15960 (N_15960,N_14801,N_14522);
or U15961 (N_15961,N_14914,N_15152);
nor U15962 (N_15962,N_14777,N_15163);
and U15963 (N_15963,N_14787,N_14869);
nand U15964 (N_15964,N_14748,N_15199);
and U15965 (N_15965,N_14557,N_14601);
and U15966 (N_15966,N_14605,N_15130);
xor U15967 (N_15967,N_14891,N_14957);
and U15968 (N_15968,N_14450,N_14987);
and U15969 (N_15969,N_14690,N_14499);
xor U15970 (N_15970,N_14442,N_14656);
and U15971 (N_15971,N_14680,N_14645);
nand U15972 (N_15972,N_14676,N_15002);
or U15973 (N_15973,N_14956,N_15123);
nand U15974 (N_15974,N_14723,N_14402);
and U15975 (N_15975,N_14473,N_14898);
and U15976 (N_15976,N_14748,N_14823);
xnor U15977 (N_15977,N_15055,N_14402);
xnor U15978 (N_15978,N_14601,N_15098);
nor U15979 (N_15979,N_14527,N_14403);
or U15980 (N_15980,N_15072,N_14443);
nor U15981 (N_15981,N_14842,N_14421);
nand U15982 (N_15982,N_15005,N_14729);
xnor U15983 (N_15983,N_14501,N_14677);
xnor U15984 (N_15984,N_14620,N_15169);
nand U15985 (N_15985,N_15153,N_14620);
nand U15986 (N_15986,N_14953,N_15055);
nand U15987 (N_15987,N_14864,N_15068);
nand U15988 (N_15988,N_14940,N_14652);
nor U15989 (N_15989,N_15091,N_15109);
xor U15990 (N_15990,N_14430,N_14621);
xnor U15991 (N_15991,N_14439,N_15112);
and U15992 (N_15992,N_14798,N_15048);
and U15993 (N_15993,N_14991,N_14734);
xnor U15994 (N_15994,N_14957,N_15103);
and U15995 (N_15995,N_14470,N_14842);
and U15996 (N_15996,N_14918,N_14794);
xor U15997 (N_15997,N_14588,N_14984);
or U15998 (N_15998,N_14466,N_14577);
and U15999 (N_15999,N_14521,N_14900);
or U16000 (N_16000,N_15713,N_15782);
nand U16001 (N_16001,N_15656,N_15666);
nor U16002 (N_16002,N_15881,N_15882);
and U16003 (N_16003,N_15488,N_15496);
nand U16004 (N_16004,N_15264,N_15277);
or U16005 (N_16005,N_15221,N_15256);
and U16006 (N_16006,N_15268,N_15891);
and U16007 (N_16007,N_15467,N_15573);
or U16008 (N_16008,N_15314,N_15602);
nand U16009 (N_16009,N_15451,N_15466);
and U16010 (N_16010,N_15606,N_15286);
xor U16011 (N_16011,N_15671,N_15381);
xor U16012 (N_16012,N_15851,N_15417);
nand U16013 (N_16013,N_15492,N_15691);
and U16014 (N_16014,N_15215,N_15257);
nand U16015 (N_16015,N_15910,N_15677);
or U16016 (N_16016,N_15911,N_15325);
nor U16017 (N_16017,N_15478,N_15834);
or U16018 (N_16018,N_15355,N_15883);
xnor U16019 (N_16019,N_15448,N_15892);
and U16020 (N_16020,N_15217,N_15820);
and U16021 (N_16021,N_15561,N_15824);
or U16022 (N_16022,N_15937,N_15383);
or U16023 (N_16023,N_15522,N_15864);
nor U16024 (N_16024,N_15955,N_15704);
xnor U16025 (N_16025,N_15690,N_15698);
nand U16026 (N_16026,N_15990,N_15896);
nand U16027 (N_16027,N_15791,N_15238);
nor U16028 (N_16028,N_15976,N_15970);
or U16029 (N_16029,N_15661,N_15736);
nand U16030 (N_16030,N_15761,N_15668);
xnor U16031 (N_16031,N_15768,N_15873);
xor U16032 (N_16032,N_15719,N_15356);
nand U16033 (N_16033,N_15537,N_15751);
and U16034 (N_16034,N_15614,N_15211);
nand U16035 (N_16035,N_15619,N_15425);
or U16036 (N_16036,N_15793,N_15795);
and U16037 (N_16037,N_15835,N_15624);
nand U16038 (N_16038,N_15975,N_15214);
nor U16039 (N_16039,N_15401,N_15311);
and U16040 (N_16040,N_15797,N_15641);
nand U16041 (N_16041,N_15905,N_15426);
or U16042 (N_16042,N_15716,N_15718);
nor U16043 (N_16043,N_15227,N_15755);
nor U16044 (N_16044,N_15515,N_15954);
nor U16045 (N_16045,N_15702,N_15309);
nor U16046 (N_16046,N_15407,N_15458);
xnor U16047 (N_16047,N_15323,N_15574);
or U16048 (N_16048,N_15950,N_15708);
nand U16049 (N_16049,N_15419,N_15831);
xnor U16050 (N_16050,N_15998,N_15326);
nand U16051 (N_16051,N_15732,N_15897);
and U16052 (N_16052,N_15332,N_15748);
nand U16053 (N_16053,N_15530,N_15610);
and U16054 (N_16054,N_15428,N_15622);
xnor U16055 (N_16055,N_15234,N_15995);
and U16056 (N_16056,N_15673,N_15549);
nor U16057 (N_16057,N_15945,N_15813);
or U16058 (N_16058,N_15894,N_15380);
nand U16059 (N_16059,N_15988,N_15302);
xnor U16060 (N_16060,N_15292,N_15633);
and U16061 (N_16061,N_15908,N_15457);
nor U16062 (N_16062,N_15735,N_15301);
xor U16063 (N_16063,N_15699,N_15915);
nand U16064 (N_16064,N_15391,N_15526);
xor U16065 (N_16065,N_15801,N_15336);
nand U16066 (N_16066,N_15290,N_15878);
nand U16067 (N_16067,N_15230,N_15559);
nor U16068 (N_16068,N_15340,N_15613);
and U16069 (N_16069,N_15552,N_15544);
xnor U16070 (N_16070,N_15934,N_15972);
nand U16071 (N_16071,N_15480,N_15463);
or U16072 (N_16072,N_15536,N_15501);
or U16073 (N_16073,N_15365,N_15600);
xnor U16074 (N_16074,N_15649,N_15669);
or U16075 (N_16075,N_15684,N_15477);
or U16076 (N_16076,N_15228,N_15476);
xor U16077 (N_16077,N_15351,N_15992);
xnor U16078 (N_16078,N_15395,N_15339);
and U16079 (N_16079,N_15293,N_15278);
nor U16080 (N_16080,N_15766,N_15361);
xnor U16081 (N_16081,N_15858,N_15479);
nand U16082 (N_16082,N_15590,N_15660);
nand U16083 (N_16083,N_15495,N_15201);
nor U16084 (N_16084,N_15728,N_15814);
xnor U16085 (N_16085,N_15281,N_15960);
nor U16086 (N_16086,N_15403,N_15371);
or U16087 (N_16087,N_15884,N_15280);
xnor U16088 (N_16088,N_15743,N_15631);
or U16089 (N_16089,N_15429,N_15289);
or U16090 (N_16090,N_15266,N_15304);
nand U16091 (N_16091,N_15294,N_15275);
nor U16092 (N_16092,N_15416,N_15785);
or U16093 (N_16093,N_15822,N_15946);
and U16094 (N_16094,N_15222,N_15672);
xnor U16095 (N_16095,N_15879,N_15978);
and U16096 (N_16096,N_15890,N_15734);
xor U16097 (N_16097,N_15900,N_15723);
or U16098 (N_16098,N_15930,N_15678);
or U16099 (N_16099,N_15907,N_15469);
and U16100 (N_16100,N_15848,N_15993);
nand U16101 (N_16101,N_15508,N_15385);
and U16102 (N_16102,N_15249,N_15541);
nor U16103 (N_16103,N_15529,N_15303);
or U16104 (N_16104,N_15453,N_15759);
xnor U16105 (N_16105,N_15717,N_15772);
xnor U16106 (N_16106,N_15564,N_15424);
nor U16107 (N_16107,N_15373,N_15260);
xnor U16108 (N_16108,N_15465,N_15956);
nor U16109 (N_16109,N_15406,N_15650);
or U16110 (N_16110,N_15977,N_15237);
or U16111 (N_16111,N_15951,N_15343);
nor U16112 (N_16112,N_15534,N_15593);
and U16113 (N_16113,N_15957,N_15357);
or U16114 (N_16114,N_15511,N_15405);
or U16115 (N_16115,N_15913,N_15812);
or U16116 (N_16116,N_15524,N_15577);
or U16117 (N_16117,N_15432,N_15438);
or U16118 (N_16118,N_15575,N_15571);
or U16119 (N_16119,N_15986,N_15832);
xor U16120 (N_16120,N_15262,N_15589);
and U16121 (N_16121,N_15692,N_15363);
and U16122 (N_16122,N_15845,N_15244);
or U16123 (N_16123,N_15578,N_15710);
and U16124 (N_16124,N_15546,N_15358);
or U16125 (N_16125,N_15909,N_15248);
nand U16126 (N_16126,N_15830,N_15700);
xnor U16127 (N_16127,N_15450,N_15617);
xnor U16128 (N_16128,N_15885,N_15291);
nand U16129 (N_16129,N_15595,N_15877);
and U16130 (N_16130,N_15826,N_15798);
or U16131 (N_16131,N_15642,N_15558);
xor U16132 (N_16132,N_15846,N_15362);
xor U16133 (N_16133,N_15963,N_15553);
nor U16134 (N_16134,N_15611,N_15923);
nand U16135 (N_16135,N_15521,N_15348);
and U16136 (N_16136,N_15654,N_15706);
or U16137 (N_16137,N_15922,N_15212);
and U16138 (N_16138,N_15647,N_15608);
nand U16139 (N_16139,N_15418,N_15497);
or U16140 (N_16140,N_15758,N_15346);
nor U16141 (N_16141,N_15844,N_15780);
and U16142 (N_16142,N_15247,N_15685);
nor U16143 (N_16143,N_15800,N_15863);
or U16144 (N_16144,N_15322,N_15338);
xor U16145 (N_16145,N_15352,N_15958);
nor U16146 (N_16146,N_15724,N_15973);
nand U16147 (N_16147,N_15505,N_15714);
nand U16148 (N_16148,N_15532,N_15583);
xnor U16149 (N_16149,N_15490,N_15412);
xor U16150 (N_16150,N_15806,N_15274);
nor U16151 (N_16151,N_15756,N_15369);
nor U16152 (N_16152,N_15841,N_15962);
or U16153 (N_16153,N_15808,N_15632);
nor U16154 (N_16154,N_15431,N_15754);
nor U16155 (N_16155,N_15737,N_15202);
or U16156 (N_16156,N_15636,N_15368);
or U16157 (N_16157,N_15967,N_15738);
xor U16158 (N_16158,N_15994,N_15764);
or U16159 (N_16159,N_15538,N_15648);
and U16160 (N_16160,N_15435,N_15367);
and U16161 (N_16161,N_15635,N_15924);
xnor U16162 (N_16162,N_15252,N_15441);
and U16163 (N_16163,N_15607,N_15439);
nor U16164 (N_16164,N_15341,N_15572);
or U16165 (N_16165,N_15484,N_15250);
nor U16166 (N_16166,N_15839,N_15686);
or U16167 (N_16167,N_15520,N_15491);
nand U16168 (N_16168,N_15517,N_15295);
xor U16169 (N_16169,N_15207,N_15833);
nand U16170 (N_16170,N_15398,N_15790);
xor U16171 (N_16171,N_15639,N_15903);
or U16172 (N_16172,N_15390,N_15442);
and U16173 (N_16173,N_15475,N_15246);
nor U16174 (N_16174,N_15665,N_15688);
or U16175 (N_16175,N_15447,N_15512);
xor U16176 (N_16176,N_15792,N_15560);
xor U16177 (N_16177,N_15499,N_15667);
and U16178 (N_16178,N_15218,N_15209);
or U16179 (N_16179,N_15916,N_15964);
and U16180 (N_16180,N_15267,N_15263);
nand U16181 (N_16181,N_15997,N_15787);
nand U16182 (N_16182,N_15444,N_15638);
xor U16183 (N_16183,N_15411,N_15461);
nand U16184 (N_16184,N_15454,N_15825);
nor U16185 (N_16185,N_15781,N_15337);
or U16186 (N_16186,N_15752,N_15370);
xor U16187 (N_16187,N_15771,N_15605);
nor U16188 (N_16188,N_15640,N_15926);
xor U16189 (N_16189,N_15456,N_15705);
nor U16190 (N_16190,N_15655,N_15566);
nand U16191 (N_16191,N_15902,N_15345);
xor U16192 (N_16192,N_15644,N_15305);
and U16193 (N_16193,N_15446,N_15927);
xnor U16194 (N_16194,N_15939,N_15270);
or U16195 (N_16195,N_15220,N_15949);
nor U16196 (N_16196,N_15223,N_15504);
nand U16197 (N_16197,N_15837,N_15464);
xnor U16198 (N_16198,N_15971,N_15414);
xor U16199 (N_16199,N_15612,N_15865);
nand U16200 (N_16200,N_15422,N_15819);
nand U16201 (N_16201,N_15952,N_15366);
xor U16202 (N_16202,N_15396,N_15204);
xnor U16203 (N_16203,N_15308,N_15265);
nand U16204 (N_16204,N_15855,N_15778);
or U16205 (N_16205,N_15460,N_15674);
nand U16206 (N_16206,N_15682,N_15298);
nand U16207 (N_16207,N_15402,N_15836);
nand U16208 (N_16208,N_15486,N_15707);
or U16209 (N_16209,N_15860,N_15443);
nand U16210 (N_16210,N_15319,N_15856);
or U16211 (N_16211,N_15662,N_15509);
or U16212 (N_16212,N_15557,N_15914);
or U16213 (N_16213,N_15585,N_15984);
xor U16214 (N_16214,N_15240,N_15519);
nor U16215 (N_16215,N_15804,N_15777);
xor U16216 (N_16216,N_15898,N_15763);
or U16217 (N_16217,N_15510,N_15818);
xor U16218 (N_16218,N_15940,N_15675);
and U16219 (N_16219,N_15842,N_15353);
and U16220 (N_16220,N_15576,N_15276);
nor U16221 (N_16221,N_15296,N_15239);
nor U16222 (N_16222,N_15592,N_15528);
and U16223 (N_16223,N_15554,N_15944);
or U16224 (N_16224,N_15929,N_15551);
xor U16225 (N_16225,N_15979,N_15947);
or U16226 (N_16226,N_15843,N_15948);
or U16227 (N_16227,N_15899,N_15657);
nand U16228 (N_16228,N_15333,N_15556);
nor U16229 (N_16229,N_15205,N_15703);
and U16230 (N_16230,N_15821,N_15874);
nor U16231 (N_16231,N_15773,N_15436);
xor U16232 (N_16232,N_15623,N_15601);
xnor U16233 (N_16233,N_15745,N_15941);
xor U16234 (N_16234,N_15387,N_15696);
xnor U16235 (N_16235,N_15681,N_15261);
or U16236 (N_16236,N_15313,N_15889);
nor U16237 (N_16237,N_15410,N_15329);
or U16238 (N_16238,N_15862,N_15533);
and U16239 (N_16239,N_15518,N_15615);
and U16240 (N_16240,N_15604,N_15854);
nor U16241 (N_16241,N_15985,N_15627);
nand U16242 (N_16242,N_15853,N_15965);
or U16243 (N_16243,N_15350,N_15769);
or U16244 (N_16244,N_15372,N_15796);
nor U16245 (N_16245,N_15581,N_15969);
and U16246 (N_16246,N_15770,N_15729);
or U16247 (N_16247,N_15720,N_15750);
nand U16248 (N_16248,N_15507,N_15200);
nor U16249 (N_16249,N_15543,N_15482);
and U16250 (N_16250,N_15774,N_15999);
nand U16251 (N_16251,N_15628,N_15321);
xor U16252 (N_16252,N_15349,N_15282);
or U16253 (N_16253,N_15550,N_15235);
or U16254 (N_16254,N_15584,N_15394);
nand U16255 (N_16255,N_15794,N_15474);
and U16256 (N_16256,N_15535,N_15823);
xnor U16257 (N_16257,N_15746,N_15680);
or U16258 (N_16258,N_15502,N_15437);
nand U16259 (N_16259,N_15503,N_15388);
nand U16260 (N_16260,N_15868,N_15386);
xor U16261 (N_16261,N_15799,N_15231);
and U16262 (N_16262,N_15376,N_15434);
or U16263 (N_16263,N_15875,N_15493);
xor U16264 (N_16264,N_15827,N_15664);
xnor U16265 (N_16265,N_15241,N_15870);
xnor U16266 (N_16266,N_15472,N_15328);
nor U16267 (N_16267,N_15789,N_15547);
nand U16268 (N_16268,N_15229,N_15727);
nand U16269 (N_16269,N_15701,N_15471);
nand U16270 (N_16270,N_15725,N_15609);
and U16271 (N_16271,N_15440,N_15857);
xor U16272 (N_16272,N_15288,N_15243);
or U16273 (N_16273,N_15829,N_15974);
or U16274 (N_16274,N_15494,N_15637);
xnor U16275 (N_16275,N_15539,N_15959);
and U16276 (N_16276,N_15562,N_15786);
or U16277 (N_16277,N_15374,N_15413);
nand U16278 (N_16278,N_15880,N_15625);
nor U16279 (N_16279,N_15310,N_15255);
nor U16280 (N_16280,N_15749,N_15359);
or U16281 (N_16281,N_15726,N_15807);
or U16282 (N_16282,N_15760,N_15579);
and U16283 (N_16283,N_15500,N_15683);
xor U16284 (N_16284,N_15315,N_15225);
xnor U16285 (N_16285,N_15563,N_15616);
nor U16286 (N_16286,N_15330,N_15936);
or U16287 (N_16287,N_15485,N_15815);
nand U16288 (N_16288,N_15364,N_15514);
or U16289 (N_16289,N_15271,N_15695);
nor U16290 (N_16290,N_15802,N_15906);
and U16291 (N_16291,N_15487,N_15320);
nor U16292 (N_16292,N_15966,N_15596);
nor U16293 (N_16293,N_15226,N_15213);
nor U16294 (N_16294,N_15850,N_15462);
nor U16295 (N_16295,N_15981,N_15810);
nor U16296 (N_16296,N_15379,N_15312);
nor U16297 (N_16297,N_15693,N_15287);
or U16298 (N_16298,N_15525,N_15459);
and U16299 (N_16299,N_15621,N_15506);
nand U16300 (N_16300,N_15811,N_15297);
nand U16301 (N_16301,N_15327,N_15569);
nand U16302 (N_16302,N_15378,N_15757);
and U16303 (N_16303,N_15861,N_15646);
or U16304 (N_16304,N_15919,N_15630);
xnor U16305 (N_16305,N_15620,N_15285);
xor U16306 (N_16306,N_15921,N_15730);
xnor U16307 (N_16307,N_15470,N_15901);
or U16308 (N_16308,N_15481,N_15817);
or U16309 (N_16309,N_15587,N_15886);
nand U16310 (N_16310,N_15849,N_15283);
nor U16311 (N_16311,N_15389,N_15382);
or U16312 (N_16312,N_15259,N_15455);
nand U16313 (N_16313,N_15876,N_15567);
or U16314 (N_16314,N_15676,N_15258);
or U16315 (N_16315,N_15603,N_15568);
nand U16316 (N_16316,N_15427,N_15887);
or U16317 (N_16317,N_15742,N_15384);
nor U16318 (N_16318,N_15762,N_15731);
nand U16319 (N_16319,N_15232,N_15210);
and U16320 (N_16320,N_15206,N_15912);
or U16321 (N_16321,N_15659,N_15473);
or U16322 (N_16322,N_15893,N_15334);
nor U16323 (N_16323,N_15803,N_15933);
and U16324 (N_16324,N_15709,N_15273);
or U16325 (N_16325,N_15580,N_15867);
or U16326 (N_16326,N_15599,N_15423);
nand U16327 (N_16327,N_15753,N_15306);
nand U16328 (N_16328,N_15242,N_15449);
xor U16329 (N_16329,N_15445,N_15219);
nor U16330 (N_16330,N_15816,N_15739);
and U16331 (N_16331,N_15740,N_15318);
or U16332 (N_16332,N_15360,N_15747);
nor U16333 (N_16333,N_15216,N_15586);
or U16334 (N_16334,N_15961,N_15943);
nor U16335 (N_16335,N_15697,N_15545);
and U16336 (N_16336,N_15653,N_15859);
nand U16337 (N_16337,N_15931,N_15775);
and U16338 (N_16338,N_15253,N_15344);
or U16339 (N_16339,N_15269,N_15399);
or U16340 (N_16340,N_15765,N_15783);
nor U16341 (N_16341,N_15408,N_15629);
nor U16342 (N_16342,N_15203,N_15430);
nand U16343 (N_16343,N_15744,N_15393);
and U16344 (N_16344,N_15987,N_15542);
and U16345 (N_16345,N_15645,N_15523);
or U16346 (N_16346,N_15888,N_15254);
or U16347 (N_16347,N_15400,N_15392);
and U16348 (N_16348,N_15869,N_15626);
or U16349 (N_16349,N_15866,N_15224);
xnor U16350 (N_16350,N_15871,N_15989);
nor U16351 (N_16351,N_15722,N_15489);
and U16352 (N_16352,N_15980,N_15307);
and U16353 (N_16353,N_15982,N_15208);
nand U16354 (N_16354,N_15588,N_15548);
nor U16355 (N_16355,N_15513,N_15925);
nand U16356 (N_16356,N_15983,N_15694);
nor U16357 (N_16357,N_15767,N_15872);
nor U16358 (N_16358,N_15643,N_15375);
xor U16359 (N_16359,N_15928,N_15377);
nand U16360 (N_16360,N_15618,N_15316);
nand U16361 (N_16361,N_15409,N_15597);
nand U16362 (N_16362,N_15299,N_15555);
and U16363 (N_16363,N_15935,N_15300);
or U16364 (N_16364,N_15942,N_15397);
xor U16365 (N_16365,N_15712,N_15779);
or U16366 (N_16366,N_15415,N_15663);
nand U16367 (N_16367,N_15452,N_15570);
nand U16368 (N_16368,N_15324,N_15828);
nand U16369 (N_16369,N_15651,N_15658);
xor U16370 (N_16370,N_15634,N_15516);
nor U16371 (N_16371,N_15582,N_15531);
nor U16372 (N_16372,N_15991,N_15904);
nand U16373 (N_16373,N_15233,N_15918);
nand U16374 (N_16374,N_15838,N_15565);
and U16375 (N_16375,N_15540,N_15968);
and U16376 (N_16376,N_15953,N_15917);
nand U16377 (N_16377,N_15687,N_15404);
xnor U16378 (N_16378,N_15784,N_15272);
xor U16379 (N_16379,N_15468,N_15805);
nand U16380 (N_16380,N_15895,N_15594);
and U16381 (N_16381,N_15421,N_15284);
nand U16382 (N_16382,N_15733,N_15741);
and U16383 (N_16383,N_15679,N_15840);
xor U16384 (N_16384,N_15347,N_15420);
or U16385 (N_16385,N_15245,N_15354);
or U16386 (N_16386,N_15996,N_15317);
or U16387 (N_16387,N_15670,N_15433);
nand U16388 (N_16388,N_15279,N_15591);
or U16389 (N_16389,N_15652,N_15711);
and U16390 (N_16390,N_15721,N_15483);
nand U16391 (N_16391,N_15920,N_15527);
or U16392 (N_16392,N_15852,N_15788);
xnor U16393 (N_16393,N_15847,N_15938);
nor U16394 (N_16394,N_15342,N_15689);
or U16395 (N_16395,N_15331,N_15932);
nor U16396 (N_16396,N_15598,N_15715);
xor U16397 (N_16397,N_15251,N_15498);
nor U16398 (N_16398,N_15236,N_15776);
and U16399 (N_16399,N_15809,N_15335);
and U16400 (N_16400,N_15887,N_15496);
nor U16401 (N_16401,N_15261,N_15371);
and U16402 (N_16402,N_15381,N_15436);
or U16403 (N_16403,N_15881,N_15696);
and U16404 (N_16404,N_15274,N_15352);
and U16405 (N_16405,N_15203,N_15494);
nand U16406 (N_16406,N_15461,N_15813);
xor U16407 (N_16407,N_15241,N_15896);
or U16408 (N_16408,N_15761,N_15363);
or U16409 (N_16409,N_15363,N_15895);
xnor U16410 (N_16410,N_15318,N_15495);
nor U16411 (N_16411,N_15486,N_15204);
nor U16412 (N_16412,N_15930,N_15300);
or U16413 (N_16413,N_15647,N_15858);
and U16414 (N_16414,N_15596,N_15970);
and U16415 (N_16415,N_15427,N_15947);
or U16416 (N_16416,N_15482,N_15985);
nor U16417 (N_16417,N_15865,N_15464);
and U16418 (N_16418,N_15552,N_15851);
nor U16419 (N_16419,N_15713,N_15840);
nand U16420 (N_16420,N_15939,N_15472);
nor U16421 (N_16421,N_15688,N_15498);
and U16422 (N_16422,N_15231,N_15801);
nor U16423 (N_16423,N_15370,N_15947);
xnor U16424 (N_16424,N_15229,N_15356);
nor U16425 (N_16425,N_15499,N_15441);
nand U16426 (N_16426,N_15399,N_15756);
xor U16427 (N_16427,N_15497,N_15436);
nor U16428 (N_16428,N_15829,N_15822);
nand U16429 (N_16429,N_15539,N_15535);
xnor U16430 (N_16430,N_15760,N_15400);
or U16431 (N_16431,N_15719,N_15692);
nor U16432 (N_16432,N_15469,N_15451);
nor U16433 (N_16433,N_15352,N_15417);
nor U16434 (N_16434,N_15455,N_15552);
or U16435 (N_16435,N_15587,N_15858);
xnor U16436 (N_16436,N_15290,N_15335);
xnor U16437 (N_16437,N_15702,N_15708);
nor U16438 (N_16438,N_15531,N_15732);
xnor U16439 (N_16439,N_15638,N_15791);
xnor U16440 (N_16440,N_15320,N_15260);
or U16441 (N_16441,N_15475,N_15356);
xnor U16442 (N_16442,N_15362,N_15826);
nand U16443 (N_16443,N_15230,N_15364);
nand U16444 (N_16444,N_15510,N_15728);
xor U16445 (N_16445,N_15322,N_15877);
nand U16446 (N_16446,N_15943,N_15259);
or U16447 (N_16447,N_15352,N_15251);
xor U16448 (N_16448,N_15787,N_15629);
xor U16449 (N_16449,N_15595,N_15254);
nor U16450 (N_16450,N_15542,N_15812);
and U16451 (N_16451,N_15273,N_15869);
nand U16452 (N_16452,N_15385,N_15461);
nand U16453 (N_16453,N_15648,N_15383);
nor U16454 (N_16454,N_15356,N_15703);
xor U16455 (N_16455,N_15744,N_15606);
nor U16456 (N_16456,N_15639,N_15517);
or U16457 (N_16457,N_15412,N_15686);
xnor U16458 (N_16458,N_15950,N_15816);
nand U16459 (N_16459,N_15477,N_15332);
xnor U16460 (N_16460,N_15538,N_15837);
xor U16461 (N_16461,N_15836,N_15604);
nand U16462 (N_16462,N_15805,N_15753);
xnor U16463 (N_16463,N_15945,N_15650);
nor U16464 (N_16464,N_15262,N_15767);
xor U16465 (N_16465,N_15361,N_15843);
xor U16466 (N_16466,N_15851,N_15218);
xor U16467 (N_16467,N_15276,N_15358);
nand U16468 (N_16468,N_15849,N_15723);
and U16469 (N_16469,N_15821,N_15545);
or U16470 (N_16470,N_15431,N_15222);
nand U16471 (N_16471,N_15612,N_15526);
nand U16472 (N_16472,N_15802,N_15890);
nor U16473 (N_16473,N_15468,N_15957);
or U16474 (N_16474,N_15524,N_15581);
and U16475 (N_16475,N_15812,N_15363);
nand U16476 (N_16476,N_15663,N_15969);
or U16477 (N_16477,N_15209,N_15742);
nor U16478 (N_16478,N_15810,N_15467);
nand U16479 (N_16479,N_15475,N_15223);
and U16480 (N_16480,N_15540,N_15988);
and U16481 (N_16481,N_15528,N_15672);
xnor U16482 (N_16482,N_15248,N_15702);
nor U16483 (N_16483,N_15946,N_15609);
and U16484 (N_16484,N_15791,N_15682);
and U16485 (N_16485,N_15452,N_15547);
xnor U16486 (N_16486,N_15615,N_15669);
nor U16487 (N_16487,N_15749,N_15881);
nand U16488 (N_16488,N_15815,N_15629);
nand U16489 (N_16489,N_15586,N_15334);
xnor U16490 (N_16490,N_15211,N_15577);
nand U16491 (N_16491,N_15488,N_15770);
xor U16492 (N_16492,N_15900,N_15752);
and U16493 (N_16493,N_15925,N_15597);
and U16494 (N_16494,N_15915,N_15393);
and U16495 (N_16495,N_15357,N_15602);
or U16496 (N_16496,N_15572,N_15994);
or U16497 (N_16497,N_15638,N_15304);
xor U16498 (N_16498,N_15802,N_15577);
nor U16499 (N_16499,N_15482,N_15939);
and U16500 (N_16500,N_15517,N_15383);
xnor U16501 (N_16501,N_15223,N_15744);
and U16502 (N_16502,N_15366,N_15662);
and U16503 (N_16503,N_15957,N_15396);
nand U16504 (N_16504,N_15635,N_15710);
xnor U16505 (N_16505,N_15963,N_15465);
nor U16506 (N_16506,N_15256,N_15969);
nor U16507 (N_16507,N_15563,N_15209);
nand U16508 (N_16508,N_15214,N_15501);
nand U16509 (N_16509,N_15299,N_15396);
nand U16510 (N_16510,N_15360,N_15824);
and U16511 (N_16511,N_15840,N_15644);
and U16512 (N_16512,N_15954,N_15945);
and U16513 (N_16513,N_15212,N_15664);
nor U16514 (N_16514,N_15990,N_15327);
nor U16515 (N_16515,N_15355,N_15632);
nor U16516 (N_16516,N_15242,N_15947);
xnor U16517 (N_16517,N_15908,N_15848);
or U16518 (N_16518,N_15424,N_15396);
xor U16519 (N_16519,N_15990,N_15223);
or U16520 (N_16520,N_15303,N_15575);
xnor U16521 (N_16521,N_15515,N_15872);
xnor U16522 (N_16522,N_15864,N_15671);
or U16523 (N_16523,N_15512,N_15682);
or U16524 (N_16524,N_15760,N_15446);
nand U16525 (N_16525,N_15302,N_15881);
nor U16526 (N_16526,N_15373,N_15570);
nand U16527 (N_16527,N_15880,N_15624);
nand U16528 (N_16528,N_15466,N_15205);
nand U16529 (N_16529,N_15735,N_15458);
and U16530 (N_16530,N_15595,N_15553);
nand U16531 (N_16531,N_15626,N_15944);
or U16532 (N_16532,N_15474,N_15966);
and U16533 (N_16533,N_15979,N_15608);
nor U16534 (N_16534,N_15931,N_15246);
nand U16535 (N_16535,N_15931,N_15971);
and U16536 (N_16536,N_15911,N_15966);
nor U16537 (N_16537,N_15227,N_15887);
and U16538 (N_16538,N_15808,N_15996);
xnor U16539 (N_16539,N_15488,N_15344);
and U16540 (N_16540,N_15322,N_15567);
nand U16541 (N_16541,N_15374,N_15629);
xor U16542 (N_16542,N_15421,N_15691);
or U16543 (N_16543,N_15717,N_15787);
and U16544 (N_16544,N_15445,N_15639);
and U16545 (N_16545,N_15231,N_15904);
and U16546 (N_16546,N_15893,N_15947);
nor U16547 (N_16547,N_15853,N_15209);
and U16548 (N_16548,N_15321,N_15347);
or U16549 (N_16549,N_15488,N_15495);
nand U16550 (N_16550,N_15250,N_15837);
and U16551 (N_16551,N_15881,N_15522);
xor U16552 (N_16552,N_15361,N_15387);
or U16553 (N_16553,N_15981,N_15270);
xnor U16554 (N_16554,N_15888,N_15390);
or U16555 (N_16555,N_15639,N_15418);
and U16556 (N_16556,N_15956,N_15757);
nand U16557 (N_16557,N_15622,N_15748);
and U16558 (N_16558,N_15220,N_15568);
and U16559 (N_16559,N_15606,N_15435);
nand U16560 (N_16560,N_15859,N_15482);
nor U16561 (N_16561,N_15279,N_15837);
or U16562 (N_16562,N_15233,N_15514);
xnor U16563 (N_16563,N_15573,N_15774);
nand U16564 (N_16564,N_15287,N_15542);
or U16565 (N_16565,N_15235,N_15267);
nor U16566 (N_16566,N_15759,N_15569);
or U16567 (N_16567,N_15663,N_15579);
and U16568 (N_16568,N_15948,N_15559);
nor U16569 (N_16569,N_15791,N_15878);
xor U16570 (N_16570,N_15539,N_15804);
nand U16571 (N_16571,N_15986,N_15331);
and U16572 (N_16572,N_15565,N_15361);
and U16573 (N_16573,N_15440,N_15603);
xnor U16574 (N_16574,N_15640,N_15747);
xor U16575 (N_16575,N_15369,N_15319);
nand U16576 (N_16576,N_15334,N_15955);
xor U16577 (N_16577,N_15312,N_15650);
xor U16578 (N_16578,N_15657,N_15422);
xnor U16579 (N_16579,N_15327,N_15543);
and U16580 (N_16580,N_15828,N_15462);
and U16581 (N_16581,N_15699,N_15331);
nand U16582 (N_16582,N_15412,N_15311);
xor U16583 (N_16583,N_15657,N_15247);
nand U16584 (N_16584,N_15853,N_15654);
xnor U16585 (N_16585,N_15550,N_15476);
nand U16586 (N_16586,N_15378,N_15836);
or U16587 (N_16587,N_15712,N_15687);
or U16588 (N_16588,N_15651,N_15462);
or U16589 (N_16589,N_15770,N_15907);
nand U16590 (N_16590,N_15631,N_15739);
or U16591 (N_16591,N_15432,N_15677);
nor U16592 (N_16592,N_15463,N_15985);
nor U16593 (N_16593,N_15723,N_15267);
or U16594 (N_16594,N_15315,N_15770);
xnor U16595 (N_16595,N_15999,N_15718);
nor U16596 (N_16596,N_15257,N_15823);
xor U16597 (N_16597,N_15304,N_15308);
or U16598 (N_16598,N_15645,N_15962);
nand U16599 (N_16599,N_15813,N_15561);
or U16600 (N_16600,N_15394,N_15467);
nand U16601 (N_16601,N_15491,N_15747);
xor U16602 (N_16602,N_15695,N_15503);
xor U16603 (N_16603,N_15203,N_15719);
nand U16604 (N_16604,N_15950,N_15778);
xnor U16605 (N_16605,N_15515,N_15800);
and U16606 (N_16606,N_15339,N_15582);
nor U16607 (N_16607,N_15916,N_15212);
xnor U16608 (N_16608,N_15660,N_15213);
and U16609 (N_16609,N_15931,N_15585);
nand U16610 (N_16610,N_15274,N_15646);
nand U16611 (N_16611,N_15412,N_15809);
and U16612 (N_16612,N_15854,N_15718);
or U16613 (N_16613,N_15320,N_15947);
xnor U16614 (N_16614,N_15727,N_15906);
nand U16615 (N_16615,N_15231,N_15657);
and U16616 (N_16616,N_15384,N_15915);
or U16617 (N_16617,N_15608,N_15308);
nand U16618 (N_16618,N_15841,N_15864);
or U16619 (N_16619,N_15668,N_15312);
or U16620 (N_16620,N_15507,N_15564);
nand U16621 (N_16621,N_15498,N_15449);
nor U16622 (N_16622,N_15433,N_15300);
nor U16623 (N_16623,N_15502,N_15358);
nand U16624 (N_16624,N_15373,N_15823);
nand U16625 (N_16625,N_15646,N_15605);
xor U16626 (N_16626,N_15654,N_15301);
nand U16627 (N_16627,N_15703,N_15665);
xor U16628 (N_16628,N_15728,N_15370);
or U16629 (N_16629,N_15686,N_15712);
and U16630 (N_16630,N_15582,N_15355);
or U16631 (N_16631,N_15579,N_15795);
nor U16632 (N_16632,N_15228,N_15423);
and U16633 (N_16633,N_15375,N_15698);
or U16634 (N_16634,N_15672,N_15596);
nor U16635 (N_16635,N_15473,N_15437);
or U16636 (N_16636,N_15545,N_15426);
and U16637 (N_16637,N_15242,N_15244);
and U16638 (N_16638,N_15940,N_15723);
or U16639 (N_16639,N_15274,N_15210);
nand U16640 (N_16640,N_15678,N_15366);
nor U16641 (N_16641,N_15239,N_15371);
nor U16642 (N_16642,N_15780,N_15517);
nor U16643 (N_16643,N_15389,N_15719);
nor U16644 (N_16644,N_15709,N_15521);
xor U16645 (N_16645,N_15484,N_15202);
xnor U16646 (N_16646,N_15873,N_15265);
nor U16647 (N_16647,N_15919,N_15575);
or U16648 (N_16648,N_15581,N_15415);
or U16649 (N_16649,N_15485,N_15311);
nand U16650 (N_16650,N_15605,N_15285);
and U16651 (N_16651,N_15899,N_15369);
xor U16652 (N_16652,N_15893,N_15802);
nor U16653 (N_16653,N_15283,N_15965);
and U16654 (N_16654,N_15508,N_15491);
and U16655 (N_16655,N_15640,N_15612);
nand U16656 (N_16656,N_15925,N_15731);
xor U16657 (N_16657,N_15520,N_15420);
xnor U16658 (N_16658,N_15394,N_15809);
xor U16659 (N_16659,N_15725,N_15239);
xor U16660 (N_16660,N_15607,N_15824);
xor U16661 (N_16661,N_15635,N_15409);
nor U16662 (N_16662,N_15473,N_15555);
or U16663 (N_16663,N_15766,N_15672);
nand U16664 (N_16664,N_15752,N_15799);
and U16665 (N_16665,N_15246,N_15940);
nor U16666 (N_16666,N_15703,N_15487);
xor U16667 (N_16667,N_15542,N_15303);
xor U16668 (N_16668,N_15900,N_15470);
and U16669 (N_16669,N_15328,N_15557);
nor U16670 (N_16670,N_15434,N_15785);
and U16671 (N_16671,N_15845,N_15771);
nand U16672 (N_16672,N_15686,N_15471);
and U16673 (N_16673,N_15662,N_15969);
and U16674 (N_16674,N_15714,N_15459);
xnor U16675 (N_16675,N_15650,N_15936);
xor U16676 (N_16676,N_15503,N_15721);
and U16677 (N_16677,N_15818,N_15236);
xor U16678 (N_16678,N_15789,N_15493);
nand U16679 (N_16679,N_15807,N_15437);
or U16680 (N_16680,N_15872,N_15816);
xnor U16681 (N_16681,N_15558,N_15330);
xor U16682 (N_16682,N_15943,N_15859);
or U16683 (N_16683,N_15750,N_15805);
and U16684 (N_16684,N_15589,N_15446);
nor U16685 (N_16685,N_15536,N_15720);
nand U16686 (N_16686,N_15950,N_15571);
nand U16687 (N_16687,N_15815,N_15769);
and U16688 (N_16688,N_15354,N_15791);
nor U16689 (N_16689,N_15513,N_15322);
or U16690 (N_16690,N_15415,N_15387);
nor U16691 (N_16691,N_15298,N_15530);
and U16692 (N_16692,N_15413,N_15608);
xor U16693 (N_16693,N_15848,N_15702);
xnor U16694 (N_16694,N_15536,N_15422);
and U16695 (N_16695,N_15930,N_15937);
and U16696 (N_16696,N_15954,N_15594);
or U16697 (N_16697,N_15384,N_15875);
xor U16698 (N_16698,N_15600,N_15472);
nor U16699 (N_16699,N_15723,N_15868);
nor U16700 (N_16700,N_15917,N_15384);
nand U16701 (N_16701,N_15564,N_15820);
nand U16702 (N_16702,N_15949,N_15491);
nor U16703 (N_16703,N_15200,N_15609);
nand U16704 (N_16704,N_15277,N_15984);
nor U16705 (N_16705,N_15472,N_15418);
and U16706 (N_16706,N_15257,N_15335);
or U16707 (N_16707,N_15460,N_15410);
nand U16708 (N_16708,N_15206,N_15770);
nand U16709 (N_16709,N_15265,N_15651);
and U16710 (N_16710,N_15240,N_15593);
nand U16711 (N_16711,N_15690,N_15314);
xor U16712 (N_16712,N_15641,N_15453);
nor U16713 (N_16713,N_15386,N_15655);
nor U16714 (N_16714,N_15811,N_15875);
xnor U16715 (N_16715,N_15812,N_15227);
or U16716 (N_16716,N_15401,N_15861);
nand U16717 (N_16717,N_15870,N_15467);
or U16718 (N_16718,N_15306,N_15777);
or U16719 (N_16719,N_15301,N_15878);
and U16720 (N_16720,N_15485,N_15700);
nor U16721 (N_16721,N_15654,N_15916);
nor U16722 (N_16722,N_15205,N_15983);
and U16723 (N_16723,N_15936,N_15646);
or U16724 (N_16724,N_15624,N_15860);
nand U16725 (N_16725,N_15757,N_15607);
xor U16726 (N_16726,N_15395,N_15437);
and U16727 (N_16727,N_15874,N_15836);
nand U16728 (N_16728,N_15594,N_15682);
or U16729 (N_16729,N_15550,N_15314);
and U16730 (N_16730,N_15738,N_15837);
nand U16731 (N_16731,N_15627,N_15673);
or U16732 (N_16732,N_15251,N_15843);
xnor U16733 (N_16733,N_15949,N_15294);
nor U16734 (N_16734,N_15862,N_15207);
or U16735 (N_16735,N_15362,N_15257);
xor U16736 (N_16736,N_15932,N_15980);
and U16737 (N_16737,N_15789,N_15373);
xor U16738 (N_16738,N_15802,N_15209);
nor U16739 (N_16739,N_15568,N_15243);
nand U16740 (N_16740,N_15718,N_15434);
nand U16741 (N_16741,N_15239,N_15600);
and U16742 (N_16742,N_15263,N_15672);
and U16743 (N_16743,N_15414,N_15359);
nand U16744 (N_16744,N_15249,N_15880);
and U16745 (N_16745,N_15283,N_15415);
and U16746 (N_16746,N_15843,N_15220);
and U16747 (N_16747,N_15848,N_15377);
xor U16748 (N_16748,N_15202,N_15207);
and U16749 (N_16749,N_15377,N_15281);
and U16750 (N_16750,N_15547,N_15258);
nor U16751 (N_16751,N_15854,N_15957);
nor U16752 (N_16752,N_15213,N_15558);
and U16753 (N_16753,N_15410,N_15708);
or U16754 (N_16754,N_15718,N_15857);
nand U16755 (N_16755,N_15643,N_15302);
nand U16756 (N_16756,N_15472,N_15288);
xnor U16757 (N_16757,N_15656,N_15348);
xnor U16758 (N_16758,N_15522,N_15746);
nand U16759 (N_16759,N_15678,N_15857);
xor U16760 (N_16760,N_15549,N_15465);
or U16761 (N_16761,N_15836,N_15321);
or U16762 (N_16762,N_15468,N_15930);
xnor U16763 (N_16763,N_15244,N_15924);
and U16764 (N_16764,N_15452,N_15881);
and U16765 (N_16765,N_15232,N_15203);
xor U16766 (N_16766,N_15667,N_15318);
or U16767 (N_16767,N_15597,N_15682);
nand U16768 (N_16768,N_15222,N_15456);
and U16769 (N_16769,N_15496,N_15970);
nor U16770 (N_16770,N_15266,N_15791);
and U16771 (N_16771,N_15379,N_15219);
xnor U16772 (N_16772,N_15416,N_15304);
and U16773 (N_16773,N_15818,N_15979);
nand U16774 (N_16774,N_15457,N_15946);
and U16775 (N_16775,N_15314,N_15834);
or U16776 (N_16776,N_15652,N_15498);
and U16777 (N_16777,N_15550,N_15302);
nor U16778 (N_16778,N_15314,N_15303);
nand U16779 (N_16779,N_15644,N_15972);
and U16780 (N_16780,N_15424,N_15823);
nand U16781 (N_16781,N_15452,N_15815);
and U16782 (N_16782,N_15219,N_15503);
xnor U16783 (N_16783,N_15905,N_15520);
and U16784 (N_16784,N_15365,N_15428);
nand U16785 (N_16785,N_15339,N_15551);
nor U16786 (N_16786,N_15407,N_15201);
nand U16787 (N_16787,N_15962,N_15304);
and U16788 (N_16788,N_15420,N_15397);
or U16789 (N_16789,N_15544,N_15642);
and U16790 (N_16790,N_15397,N_15240);
xnor U16791 (N_16791,N_15407,N_15781);
or U16792 (N_16792,N_15343,N_15547);
and U16793 (N_16793,N_15400,N_15271);
nor U16794 (N_16794,N_15702,N_15726);
xnor U16795 (N_16795,N_15967,N_15673);
or U16796 (N_16796,N_15761,N_15406);
xnor U16797 (N_16797,N_15762,N_15252);
xnor U16798 (N_16798,N_15386,N_15599);
xnor U16799 (N_16799,N_15559,N_15637);
nor U16800 (N_16800,N_16712,N_16685);
nor U16801 (N_16801,N_16124,N_16045);
nor U16802 (N_16802,N_16311,N_16738);
xnor U16803 (N_16803,N_16742,N_16037);
xor U16804 (N_16804,N_16617,N_16403);
nor U16805 (N_16805,N_16533,N_16273);
or U16806 (N_16806,N_16492,N_16352);
and U16807 (N_16807,N_16391,N_16298);
or U16808 (N_16808,N_16219,N_16699);
and U16809 (N_16809,N_16146,N_16212);
nor U16810 (N_16810,N_16556,N_16017);
xor U16811 (N_16811,N_16153,N_16511);
nor U16812 (N_16812,N_16449,N_16107);
nand U16813 (N_16813,N_16325,N_16058);
and U16814 (N_16814,N_16784,N_16084);
or U16815 (N_16815,N_16276,N_16326);
xnor U16816 (N_16816,N_16248,N_16178);
nor U16817 (N_16817,N_16207,N_16719);
or U16818 (N_16818,N_16134,N_16695);
and U16819 (N_16819,N_16039,N_16554);
and U16820 (N_16820,N_16289,N_16531);
nor U16821 (N_16821,N_16680,N_16229);
xnor U16822 (N_16822,N_16164,N_16597);
and U16823 (N_16823,N_16372,N_16615);
xor U16824 (N_16824,N_16484,N_16553);
and U16825 (N_16825,N_16452,N_16131);
and U16826 (N_16826,N_16038,N_16413);
nand U16827 (N_16827,N_16123,N_16566);
and U16828 (N_16828,N_16697,N_16135);
nand U16829 (N_16829,N_16540,N_16555);
nand U16830 (N_16830,N_16429,N_16430);
nand U16831 (N_16831,N_16184,N_16225);
or U16832 (N_16832,N_16376,N_16684);
and U16833 (N_16833,N_16522,N_16646);
nand U16834 (N_16834,N_16573,N_16033);
nand U16835 (N_16835,N_16424,N_16661);
nor U16836 (N_16836,N_16381,N_16499);
and U16837 (N_16837,N_16004,N_16655);
and U16838 (N_16838,N_16741,N_16223);
and U16839 (N_16839,N_16643,N_16454);
or U16840 (N_16840,N_16075,N_16588);
or U16841 (N_16841,N_16116,N_16503);
xor U16842 (N_16842,N_16176,N_16189);
or U16843 (N_16843,N_16027,N_16118);
xnor U16844 (N_16844,N_16291,N_16609);
nor U16845 (N_16845,N_16431,N_16122);
or U16846 (N_16846,N_16532,N_16401);
and U16847 (N_16847,N_16305,N_16638);
nand U16848 (N_16848,N_16036,N_16493);
nor U16849 (N_16849,N_16689,N_16177);
or U16850 (N_16850,N_16256,N_16001);
xor U16851 (N_16851,N_16120,N_16307);
xor U16852 (N_16852,N_16789,N_16716);
and U16853 (N_16853,N_16147,N_16560);
nand U16854 (N_16854,N_16386,N_16073);
xor U16855 (N_16855,N_16010,N_16018);
and U16856 (N_16856,N_16347,N_16142);
and U16857 (N_16857,N_16420,N_16589);
or U16858 (N_16858,N_16415,N_16734);
nor U16859 (N_16859,N_16737,N_16568);
xor U16860 (N_16860,N_16149,N_16151);
nand U16861 (N_16861,N_16557,N_16337);
nor U16862 (N_16862,N_16214,N_16119);
nor U16863 (N_16863,N_16239,N_16731);
nor U16864 (N_16864,N_16726,N_16714);
xnor U16865 (N_16865,N_16088,N_16282);
and U16866 (N_16866,N_16315,N_16414);
xor U16867 (N_16867,N_16012,N_16361);
or U16868 (N_16868,N_16469,N_16693);
xor U16869 (N_16869,N_16482,N_16561);
or U16870 (N_16870,N_16312,N_16495);
and U16871 (N_16871,N_16517,N_16261);
nor U16872 (N_16872,N_16764,N_16270);
and U16873 (N_16873,N_16190,N_16504);
xnor U16874 (N_16874,N_16290,N_16095);
xnor U16875 (N_16875,N_16127,N_16034);
or U16876 (N_16876,N_16096,N_16254);
xnor U16877 (N_16877,N_16098,N_16519);
xnor U16878 (N_16878,N_16623,N_16668);
nor U16879 (N_16879,N_16777,N_16404);
and U16880 (N_16880,N_16303,N_16411);
or U16881 (N_16881,N_16093,N_16494);
or U16882 (N_16882,N_16729,N_16071);
and U16883 (N_16883,N_16160,N_16125);
xnor U16884 (N_16884,N_16245,N_16000);
and U16885 (N_16885,N_16199,N_16152);
or U16886 (N_16886,N_16306,N_16733);
or U16887 (N_16887,N_16537,N_16259);
and U16888 (N_16888,N_16175,N_16479);
nor U16889 (N_16889,N_16687,N_16209);
nor U16890 (N_16890,N_16294,N_16456);
xor U16891 (N_16891,N_16678,N_16062);
and U16892 (N_16892,N_16525,N_16637);
or U16893 (N_16893,N_16535,N_16630);
nor U16894 (N_16894,N_16044,N_16309);
or U16895 (N_16895,N_16483,N_16410);
nor U16896 (N_16896,N_16222,N_16613);
xor U16897 (N_16897,N_16193,N_16496);
and U16898 (N_16898,N_16536,N_16473);
or U16899 (N_16899,N_16766,N_16300);
or U16900 (N_16900,N_16232,N_16057);
or U16901 (N_16901,N_16752,N_16360);
and U16902 (N_16902,N_16331,N_16648);
nand U16903 (N_16903,N_16626,N_16156);
nand U16904 (N_16904,N_16007,N_16663);
or U16905 (N_16905,N_16115,N_16770);
or U16906 (N_16906,N_16409,N_16612);
nor U16907 (N_16907,N_16500,N_16709);
xnor U16908 (N_16908,N_16130,N_16246);
or U16909 (N_16909,N_16757,N_16754);
or U16910 (N_16910,N_16335,N_16328);
xnor U16911 (N_16911,N_16079,N_16393);
xnor U16912 (N_16912,N_16200,N_16489);
and U16913 (N_16913,N_16744,N_16475);
nor U16914 (N_16914,N_16605,N_16608);
or U16915 (N_16915,N_16275,N_16435);
and U16916 (N_16916,N_16002,N_16292);
and U16917 (N_16917,N_16128,N_16715);
nor U16918 (N_16918,N_16213,N_16692);
nand U16919 (N_16919,N_16284,N_16451);
xor U16920 (N_16920,N_16694,N_16308);
and U16921 (N_16921,N_16750,N_16669);
nand U16922 (N_16922,N_16696,N_16793);
or U16923 (N_16923,N_16481,N_16534);
or U16924 (N_16924,N_16163,N_16286);
nor U16925 (N_16925,N_16129,N_16285);
nor U16926 (N_16926,N_16183,N_16139);
nor U16927 (N_16927,N_16353,N_16601);
nor U16928 (N_16928,N_16249,N_16218);
or U16929 (N_16929,N_16400,N_16264);
xor U16930 (N_16930,N_16477,N_16405);
or U16931 (N_16931,N_16437,N_16610);
nor U16932 (N_16932,N_16216,N_16467);
nand U16933 (N_16933,N_16108,N_16649);
xnor U16934 (N_16934,N_16448,N_16572);
nor U16935 (N_16935,N_16329,N_16665);
nand U16936 (N_16936,N_16583,N_16418);
or U16937 (N_16937,N_16730,N_16580);
or U16938 (N_16938,N_16510,N_16453);
nand U16939 (N_16939,N_16136,N_16625);
nor U16940 (N_16940,N_16322,N_16528);
or U16941 (N_16941,N_16594,N_16578);
nand U16942 (N_16942,N_16640,N_16090);
xor U16943 (N_16943,N_16769,N_16094);
and U16944 (N_16944,N_16539,N_16201);
or U16945 (N_16945,N_16546,N_16547);
and U16946 (N_16946,N_16097,N_16584);
and U16947 (N_16947,N_16611,N_16382);
or U16948 (N_16948,N_16622,N_16564);
xnor U16949 (N_16949,N_16652,N_16518);
or U16950 (N_16950,N_16049,N_16502);
nand U16951 (N_16951,N_16604,N_16362);
xnor U16952 (N_16952,N_16722,N_16272);
nor U16953 (N_16953,N_16340,N_16215);
or U16954 (N_16954,N_16258,N_16042);
xor U16955 (N_16955,N_16498,N_16639);
and U16956 (N_16956,N_16055,N_16641);
and U16957 (N_16957,N_16569,N_16582);
nor U16958 (N_16958,N_16188,N_16666);
nand U16959 (N_16959,N_16278,N_16544);
and U16960 (N_16960,N_16732,N_16185);
nor U16961 (N_16961,N_16776,N_16645);
xor U16962 (N_16962,N_16579,N_16542);
nand U16963 (N_16963,N_16713,N_16304);
or U16964 (N_16964,N_16792,N_16236);
nand U16965 (N_16965,N_16231,N_16054);
xor U16966 (N_16966,N_16059,N_16791);
nor U16967 (N_16967,N_16591,N_16174);
nor U16968 (N_16968,N_16786,N_16047);
or U16969 (N_16969,N_16455,N_16636);
or U16970 (N_16970,N_16653,N_16723);
or U16971 (N_16971,N_16150,N_16364);
xor U16972 (N_16972,N_16756,N_16026);
nand U16973 (N_16973,N_16576,N_16602);
and U16974 (N_16974,N_16395,N_16682);
and U16975 (N_16975,N_16771,N_16702);
or U16976 (N_16976,N_16043,N_16006);
nor U16977 (N_16977,N_16182,N_16552);
or U16978 (N_16978,N_16755,N_16472);
or U16979 (N_16979,N_16747,N_16488);
xor U16980 (N_16980,N_16787,N_16132);
xor U16981 (N_16981,N_16072,N_16330);
nor U16982 (N_16982,N_16657,N_16767);
nand U16983 (N_16983,N_16367,N_16628);
xnor U16984 (N_16984,N_16436,N_16562);
nand U16985 (N_16985,N_16461,N_16110);
or U16986 (N_16986,N_16425,N_16344);
nand U16987 (N_16987,N_16061,N_16359);
nor U16988 (N_16988,N_16357,N_16619);
xor U16989 (N_16989,N_16016,N_16363);
nor U16990 (N_16990,N_16217,N_16234);
nand U16991 (N_16991,N_16111,N_16023);
and U16992 (N_16992,N_16796,N_16099);
xnor U16993 (N_16993,N_16237,N_16720);
nand U16994 (N_16994,N_16512,N_16463);
nand U16995 (N_16995,N_16013,N_16358);
or U16996 (N_16996,N_16029,N_16240);
or U16997 (N_16997,N_16567,N_16066);
xnor U16998 (N_16998,N_16736,N_16080);
and U16999 (N_16999,N_16667,N_16725);
xor U17000 (N_17000,N_16250,N_16423);
or U17001 (N_17001,N_16140,N_16670);
nor U17002 (N_17002,N_16799,N_16197);
and U17003 (N_17003,N_16334,N_16025);
or U17004 (N_17004,N_16050,N_16078);
xor U17005 (N_17005,N_16592,N_16775);
nand U17006 (N_17006,N_16320,N_16024);
xor U17007 (N_17007,N_16447,N_16076);
nor U17008 (N_17008,N_16144,N_16549);
or U17009 (N_17009,N_16032,N_16356);
nor U17010 (N_17010,N_16260,N_16263);
or U17011 (N_17011,N_16656,N_16782);
and U17012 (N_17012,N_16779,N_16465);
and U17013 (N_17013,N_16265,N_16206);
or U17014 (N_17014,N_16087,N_16082);
nand U17015 (N_17015,N_16471,N_16121);
xor U17016 (N_17016,N_16745,N_16527);
xnor U17017 (N_17017,N_16041,N_16476);
xor U17018 (N_17018,N_16717,N_16487);
nor U17019 (N_17019,N_16235,N_16545);
xor U17020 (N_17020,N_16468,N_16179);
xor U17021 (N_17021,N_16407,N_16438);
or U17022 (N_17022,N_16154,N_16421);
and U17023 (N_17023,N_16574,N_16040);
or U17024 (N_17024,N_16313,N_16633);
nor U17025 (N_17025,N_16297,N_16681);
nor U17026 (N_17026,N_16384,N_16180);
nand U17027 (N_17027,N_16171,N_16718);
and U17028 (N_17028,N_16051,N_16432);
xor U17029 (N_17029,N_16046,N_16759);
or U17030 (N_17030,N_16672,N_16052);
and U17031 (N_17031,N_16513,N_16145);
or U17032 (N_17032,N_16346,N_16683);
xor U17033 (N_17033,N_16104,N_16283);
xnor U17034 (N_17034,N_16708,N_16618);
or U17035 (N_17035,N_16318,N_16571);
nor U17036 (N_17036,N_16005,N_16558);
nor U17037 (N_17037,N_16203,N_16761);
and U17038 (N_17038,N_16100,N_16398);
or U17039 (N_17039,N_16490,N_16048);
or U17040 (N_17040,N_16390,N_16768);
xor U17041 (N_17041,N_16575,N_16676);
or U17042 (N_17042,N_16780,N_16157);
and U17043 (N_17043,N_16243,N_16763);
or U17044 (N_17044,N_16370,N_16614);
or U17045 (N_17045,N_16508,N_16607);
and U17046 (N_17046,N_16762,N_16365);
and U17047 (N_17047,N_16711,N_16267);
nand U17048 (N_17048,N_16765,N_16773);
nor U17049 (N_17049,N_16426,N_16748);
xnor U17050 (N_17050,N_16143,N_16368);
or U17051 (N_17051,N_16620,N_16529);
nand U17052 (N_17052,N_16538,N_16374);
nand U17053 (N_17053,N_16408,N_16380);
or U17054 (N_17054,N_16478,N_16541);
or U17055 (N_17055,N_16590,N_16659);
xor U17056 (N_17056,N_16596,N_16443);
nor U17057 (N_17057,N_16551,N_16707);
nand U17058 (N_17058,N_16230,N_16686);
nor U17059 (N_17059,N_16226,N_16795);
and U17060 (N_17060,N_16210,N_16585);
or U17061 (N_17061,N_16507,N_16383);
and U17062 (N_17062,N_16158,N_16774);
and U17063 (N_17063,N_16599,N_16621);
nand U17064 (N_17064,N_16654,N_16092);
nand U17065 (N_17065,N_16205,N_16195);
nor U17066 (N_17066,N_16375,N_16412);
xnor U17067 (N_17067,N_16251,N_16015);
nand U17068 (N_17068,N_16349,N_16089);
nand U17069 (N_17069,N_16606,N_16269);
xnor U17070 (N_17070,N_16598,N_16371);
nand U17071 (N_17071,N_16319,N_16137);
nor U17072 (N_17072,N_16586,N_16563);
and U17073 (N_17073,N_16063,N_16113);
nor U17074 (N_17074,N_16753,N_16740);
xnor U17075 (N_17075,N_16422,N_16470);
xnor U17076 (N_17076,N_16444,N_16194);
or U17077 (N_17077,N_16701,N_16397);
nor U17078 (N_17078,N_16523,N_16280);
and U17079 (N_17079,N_16650,N_16241);
nand U17080 (N_17080,N_16068,N_16354);
and U17081 (N_17081,N_16760,N_16069);
and U17082 (N_17082,N_16279,N_16735);
and U17083 (N_17083,N_16281,N_16434);
or U17084 (N_17084,N_16081,N_16746);
or U17085 (N_17085,N_16227,N_16021);
xnor U17086 (N_17086,N_16662,N_16106);
or U17087 (N_17087,N_16783,N_16343);
nor U17088 (N_17088,N_16515,N_16797);
or U17089 (N_17089,N_16440,N_16242);
nor U17090 (N_17090,N_16060,N_16141);
and U17091 (N_17091,N_16366,N_16521);
xnor U17092 (N_17092,N_16168,N_16014);
nor U17093 (N_17093,N_16394,N_16244);
nor U17094 (N_17094,N_16446,N_16170);
or U17095 (N_17095,N_16565,N_16067);
and U17096 (N_17096,N_16458,N_16065);
and U17097 (N_17097,N_16327,N_16387);
and U17098 (N_17098,N_16671,N_16406);
nor U17099 (N_17099,N_16530,N_16083);
nand U17100 (N_17100,N_16520,N_16485);
or U17101 (N_17101,N_16674,N_16003);
and U17102 (N_17102,N_16442,N_16101);
and U17103 (N_17103,N_16064,N_16202);
or U17104 (N_17104,N_16192,N_16798);
xor U17105 (N_17105,N_16324,N_16457);
nor U17106 (N_17106,N_16155,N_16355);
and U17107 (N_17107,N_16651,N_16186);
and U17108 (N_17108,N_16271,N_16758);
or U17109 (N_17109,N_16332,N_16388);
xor U17110 (N_17110,N_16698,N_16439);
or U17111 (N_17111,N_16728,N_16166);
nor U17112 (N_17112,N_16486,N_16316);
or U17113 (N_17113,N_16196,N_16516);
and U17114 (N_17114,N_16600,N_16379);
or U17115 (N_17115,N_16691,N_16314);
and U17116 (N_17116,N_16373,N_16474);
and U17117 (N_17117,N_16342,N_16233);
nor U17118 (N_17118,N_16008,N_16570);
and U17119 (N_17119,N_16739,N_16399);
and U17120 (N_17120,N_16109,N_16743);
nor U17121 (N_17121,N_16724,N_16165);
nor U17122 (N_17122,N_16338,N_16028);
or U17123 (N_17123,N_16035,N_16169);
nor U17124 (N_17124,N_16255,N_16339);
nor U17125 (N_17125,N_16056,N_16117);
or U17126 (N_17126,N_16198,N_16514);
or U17127 (N_17127,N_16632,N_16491);
xnor U17128 (N_17128,N_16257,N_16268);
nand U17129 (N_17129,N_16505,N_16660);
nand U17130 (N_17130,N_16497,N_16710);
nor U17131 (N_17131,N_16595,N_16385);
nand U17132 (N_17132,N_16704,N_16204);
and U17133 (N_17133,N_16091,N_16070);
nand U17134 (N_17134,N_16266,N_16428);
xnor U17135 (N_17135,N_16159,N_16301);
nor U17136 (N_17136,N_16794,N_16550);
xor U17137 (N_17137,N_16296,N_16627);
xor U17138 (N_17138,N_16220,N_16228);
xnor U17139 (N_17139,N_16103,N_16524);
nand U17140 (N_17140,N_16624,N_16333);
or U17141 (N_17141,N_16378,N_16173);
or U17142 (N_17142,N_16350,N_16105);
xor U17143 (N_17143,N_16679,N_16148);
or U17144 (N_17144,N_16790,N_16074);
or U17145 (N_17145,N_16441,N_16020);
xor U17146 (N_17146,N_16114,N_16011);
and U17147 (N_17147,N_16433,N_16019);
and U17148 (N_17148,N_16543,N_16673);
nand U17149 (N_17149,N_16721,N_16022);
and U17150 (N_17150,N_16252,N_16727);
or U17151 (N_17151,N_16288,N_16581);
nand U17152 (N_17152,N_16772,N_16277);
nand U17153 (N_17153,N_16647,N_16295);
nor U17154 (N_17154,N_16077,N_16253);
and U17155 (N_17155,N_16187,N_16167);
or U17156 (N_17156,N_16642,N_16688);
or U17157 (N_17157,N_16238,N_16402);
nor U17158 (N_17158,N_16593,N_16459);
or U17159 (N_17159,N_16631,N_16191);
or U17160 (N_17160,N_16427,N_16785);
nand U17161 (N_17161,N_16526,N_16161);
or U17162 (N_17162,N_16392,N_16788);
or U17163 (N_17163,N_16247,N_16085);
nor U17164 (N_17164,N_16112,N_16172);
xor U17165 (N_17165,N_16506,N_16287);
and U17166 (N_17166,N_16703,N_16480);
or U17167 (N_17167,N_16181,N_16417);
xnor U17168 (N_17168,N_16781,N_16224);
xor U17169 (N_17169,N_16030,N_16749);
xor U17170 (N_17170,N_16644,N_16445);
xor U17171 (N_17171,N_16658,N_16664);
nor U17172 (N_17172,N_16321,N_16396);
nor U17173 (N_17173,N_16462,N_16501);
nand U17174 (N_17174,N_16336,N_16706);
and U17175 (N_17175,N_16629,N_16126);
or U17176 (N_17176,N_16675,N_16419);
nand U17177 (N_17177,N_16031,N_16345);
xnor U17178 (N_17178,N_16450,N_16138);
nand U17179 (N_17179,N_16262,N_16466);
nand U17180 (N_17180,N_16208,N_16548);
nand U17181 (N_17181,N_16369,N_16133);
xnor U17182 (N_17182,N_16690,N_16700);
xor U17183 (N_17183,N_16603,N_16635);
nor U17184 (N_17184,N_16211,N_16377);
or U17185 (N_17185,N_16351,N_16416);
xnor U17186 (N_17186,N_16341,N_16634);
and U17187 (N_17187,N_16274,N_16317);
nand U17188 (N_17188,N_16348,N_16778);
nor U17189 (N_17189,N_16299,N_16705);
or U17190 (N_17190,N_16221,N_16293);
or U17191 (N_17191,N_16464,N_16751);
and U17192 (N_17192,N_16389,N_16559);
nor U17193 (N_17193,N_16302,N_16509);
nand U17194 (N_17194,N_16587,N_16310);
or U17195 (N_17195,N_16577,N_16460);
nor U17196 (N_17196,N_16677,N_16102);
nor U17197 (N_17197,N_16616,N_16009);
and U17198 (N_17198,N_16323,N_16086);
nor U17199 (N_17199,N_16053,N_16162);
and U17200 (N_17200,N_16464,N_16369);
nand U17201 (N_17201,N_16398,N_16585);
and U17202 (N_17202,N_16753,N_16727);
nand U17203 (N_17203,N_16122,N_16121);
or U17204 (N_17204,N_16512,N_16700);
xor U17205 (N_17205,N_16760,N_16470);
nand U17206 (N_17206,N_16042,N_16163);
nand U17207 (N_17207,N_16068,N_16795);
and U17208 (N_17208,N_16607,N_16429);
xnor U17209 (N_17209,N_16031,N_16142);
or U17210 (N_17210,N_16554,N_16396);
xnor U17211 (N_17211,N_16477,N_16655);
xnor U17212 (N_17212,N_16622,N_16359);
and U17213 (N_17213,N_16257,N_16536);
and U17214 (N_17214,N_16080,N_16501);
and U17215 (N_17215,N_16045,N_16642);
nor U17216 (N_17216,N_16054,N_16245);
nor U17217 (N_17217,N_16581,N_16478);
nand U17218 (N_17218,N_16063,N_16789);
or U17219 (N_17219,N_16480,N_16376);
or U17220 (N_17220,N_16386,N_16506);
nor U17221 (N_17221,N_16514,N_16637);
nor U17222 (N_17222,N_16298,N_16790);
nor U17223 (N_17223,N_16591,N_16669);
nand U17224 (N_17224,N_16111,N_16798);
and U17225 (N_17225,N_16635,N_16699);
or U17226 (N_17226,N_16706,N_16393);
and U17227 (N_17227,N_16684,N_16754);
xnor U17228 (N_17228,N_16750,N_16128);
nand U17229 (N_17229,N_16421,N_16780);
nand U17230 (N_17230,N_16671,N_16312);
xnor U17231 (N_17231,N_16153,N_16689);
and U17232 (N_17232,N_16189,N_16033);
xor U17233 (N_17233,N_16205,N_16389);
nor U17234 (N_17234,N_16073,N_16378);
nand U17235 (N_17235,N_16457,N_16739);
and U17236 (N_17236,N_16537,N_16557);
xnor U17237 (N_17237,N_16554,N_16707);
xor U17238 (N_17238,N_16090,N_16104);
nor U17239 (N_17239,N_16543,N_16390);
or U17240 (N_17240,N_16245,N_16585);
xor U17241 (N_17241,N_16375,N_16775);
xnor U17242 (N_17242,N_16110,N_16386);
nand U17243 (N_17243,N_16431,N_16721);
and U17244 (N_17244,N_16197,N_16435);
or U17245 (N_17245,N_16211,N_16420);
and U17246 (N_17246,N_16310,N_16406);
or U17247 (N_17247,N_16426,N_16339);
nand U17248 (N_17248,N_16712,N_16470);
nor U17249 (N_17249,N_16661,N_16708);
xor U17250 (N_17250,N_16651,N_16069);
or U17251 (N_17251,N_16284,N_16399);
nor U17252 (N_17252,N_16030,N_16025);
and U17253 (N_17253,N_16139,N_16526);
xor U17254 (N_17254,N_16604,N_16676);
xnor U17255 (N_17255,N_16327,N_16058);
nand U17256 (N_17256,N_16384,N_16342);
nand U17257 (N_17257,N_16240,N_16583);
and U17258 (N_17258,N_16534,N_16170);
nor U17259 (N_17259,N_16757,N_16328);
nand U17260 (N_17260,N_16749,N_16248);
nor U17261 (N_17261,N_16158,N_16790);
or U17262 (N_17262,N_16546,N_16109);
nand U17263 (N_17263,N_16358,N_16778);
nand U17264 (N_17264,N_16022,N_16663);
or U17265 (N_17265,N_16716,N_16667);
nand U17266 (N_17266,N_16284,N_16015);
nand U17267 (N_17267,N_16674,N_16058);
xnor U17268 (N_17268,N_16176,N_16709);
nand U17269 (N_17269,N_16422,N_16493);
nor U17270 (N_17270,N_16006,N_16441);
nor U17271 (N_17271,N_16315,N_16186);
nor U17272 (N_17272,N_16514,N_16144);
nor U17273 (N_17273,N_16727,N_16108);
nor U17274 (N_17274,N_16733,N_16305);
xor U17275 (N_17275,N_16736,N_16669);
and U17276 (N_17276,N_16727,N_16766);
nand U17277 (N_17277,N_16245,N_16697);
xnor U17278 (N_17278,N_16225,N_16272);
or U17279 (N_17279,N_16486,N_16491);
or U17280 (N_17280,N_16669,N_16675);
nand U17281 (N_17281,N_16608,N_16553);
and U17282 (N_17282,N_16237,N_16680);
nor U17283 (N_17283,N_16759,N_16262);
nand U17284 (N_17284,N_16479,N_16754);
xnor U17285 (N_17285,N_16768,N_16446);
xor U17286 (N_17286,N_16680,N_16486);
xor U17287 (N_17287,N_16713,N_16430);
xnor U17288 (N_17288,N_16172,N_16008);
nor U17289 (N_17289,N_16296,N_16282);
nor U17290 (N_17290,N_16715,N_16655);
or U17291 (N_17291,N_16718,N_16232);
nand U17292 (N_17292,N_16660,N_16515);
or U17293 (N_17293,N_16360,N_16011);
nand U17294 (N_17294,N_16202,N_16368);
and U17295 (N_17295,N_16709,N_16457);
nand U17296 (N_17296,N_16304,N_16655);
and U17297 (N_17297,N_16704,N_16778);
and U17298 (N_17298,N_16222,N_16644);
xnor U17299 (N_17299,N_16731,N_16566);
and U17300 (N_17300,N_16785,N_16452);
nor U17301 (N_17301,N_16278,N_16796);
xor U17302 (N_17302,N_16020,N_16620);
nand U17303 (N_17303,N_16388,N_16172);
nand U17304 (N_17304,N_16187,N_16135);
or U17305 (N_17305,N_16388,N_16319);
nor U17306 (N_17306,N_16657,N_16323);
xnor U17307 (N_17307,N_16625,N_16422);
and U17308 (N_17308,N_16020,N_16159);
or U17309 (N_17309,N_16715,N_16709);
xnor U17310 (N_17310,N_16706,N_16760);
nand U17311 (N_17311,N_16102,N_16494);
and U17312 (N_17312,N_16224,N_16262);
xor U17313 (N_17313,N_16595,N_16419);
and U17314 (N_17314,N_16495,N_16118);
nand U17315 (N_17315,N_16487,N_16265);
or U17316 (N_17316,N_16012,N_16559);
or U17317 (N_17317,N_16170,N_16613);
and U17318 (N_17318,N_16054,N_16633);
and U17319 (N_17319,N_16562,N_16186);
and U17320 (N_17320,N_16654,N_16139);
or U17321 (N_17321,N_16362,N_16566);
xnor U17322 (N_17322,N_16132,N_16228);
and U17323 (N_17323,N_16623,N_16410);
and U17324 (N_17324,N_16722,N_16448);
xor U17325 (N_17325,N_16464,N_16259);
nor U17326 (N_17326,N_16227,N_16372);
nand U17327 (N_17327,N_16788,N_16165);
and U17328 (N_17328,N_16050,N_16199);
nor U17329 (N_17329,N_16590,N_16277);
xor U17330 (N_17330,N_16537,N_16233);
nand U17331 (N_17331,N_16203,N_16660);
xor U17332 (N_17332,N_16067,N_16722);
and U17333 (N_17333,N_16131,N_16048);
or U17334 (N_17334,N_16567,N_16584);
nor U17335 (N_17335,N_16746,N_16773);
or U17336 (N_17336,N_16234,N_16058);
or U17337 (N_17337,N_16252,N_16090);
or U17338 (N_17338,N_16799,N_16645);
or U17339 (N_17339,N_16230,N_16284);
nor U17340 (N_17340,N_16402,N_16572);
and U17341 (N_17341,N_16700,N_16470);
or U17342 (N_17342,N_16397,N_16754);
nand U17343 (N_17343,N_16642,N_16040);
xnor U17344 (N_17344,N_16545,N_16679);
xnor U17345 (N_17345,N_16671,N_16418);
and U17346 (N_17346,N_16529,N_16191);
or U17347 (N_17347,N_16533,N_16622);
and U17348 (N_17348,N_16155,N_16445);
nand U17349 (N_17349,N_16657,N_16102);
and U17350 (N_17350,N_16352,N_16563);
nand U17351 (N_17351,N_16163,N_16500);
and U17352 (N_17352,N_16212,N_16578);
xor U17353 (N_17353,N_16603,N_16659);
xor U17354 (N_17354,N_16429,N_16788);
xor U17355 (N_17355,N_16753,N_16630);
or U17356 (N_17356,N_16086,N_16035);
xnor U17357 (N_17357,N_16435,N_16492);
nor U17358 (N_17358,N_16700,N_16238);
xnor U17359 (N_17359,N_16129,N_16798);
xnor U17360 (N_17360,N_16391,N_16271);
nand U17361 (N_17361,N_16352,N_16626);
and U17362 (N_17362,N_16289,N_16177);
nand U17363 (N_17363,N_16596,N_16041);
nor U17364 (N_17364,N_16400,N_16365);
or U17365 (N_17365,N_16467,N_16594);
nor U17366 (N_17366,N_16783,N_16095);
or U17367 (N_17367,N_16330,N_16796);
or U17368 (N_17368,N_16004,N_16192);
and U17369 (N_17369,N_16385,N_16555);
xnor U17370 (N_17370,N_16587,N_16650);
nand U17371 (N_17371,N_16736,N_16462);
nand U17372 (N_17372,N_16014,N_16401);
xor U17373 (N_17373,N_16408,N_16403);
xor U17374 (N_17374,N_16472,N_16336);
nand U17375 (N_17375,N_16413,N_16765);
nand U17376 (N_17376,N_16364,N_16494);
xnor U17377 (N_17377,N_16104,N_16293);
nand U17378 (N_17378,N_16754,N_16203);
xor U17379 (N_17379,N_16248,N_16538);
xnor U17380 (N_17380,N_16255,N_16301);
or U17381 (N_17381,N_16788,N_16075);
or U17382 (N_17382,N_16632,N_16397);
and U17383 (N_17383,N_16439,N_16108);
or U17384 (N_17384,N_16699,N_16611);
nor U17385 (N_17385,N_16265,N_16361);
nand U17386 (N_17386,N_16386,N_16077);
or U17387 (N_17387,N_16491,N_16701);
nor U17388 (N_17388,N_16174,N_16018);
and U17389 (N_17389,N_16156,N_16767);
nand U17390 (N_17390,N_16521,N_16210);
and U17391 (N_17391,N_16540,N_16045);
and U17392 (N_17392,N_16546,N_16469);
or U17393 (N_17393,N_16131,N_16664);
xnor U17394 (N_17394,N_16459,N_16336);
and U17395 (N_17395,N_16070,N_16313);
xnor U17396 (N_17396,N_16156,N_16320);
and U17397 (N_17397,N_16535,N_16079);
or U17398 (N_17398,N_16387,N_16758);
nand U17399 (N_17399,N_16467,N_16391);
or U17400 (N_17400,N_16285,N_16567);
nor U17401 (N_17401,N_16703,N_16059);
or U17402 (N_17402,N_16531,N_16553);
or U17403 (N_17403,N_16229,N_16244);
nor U17404 (N_17404,N_16432,N_16402);
xor U17405 (N_17405,N_16697,N_16567);
or U17406 (N_17406,N_16498,N_16021);
and U17407 (N_17407,N_16503,N_16681);
nor U17408 (N_17408,N_16676,N_16532);
nor U17409 (N_17409,N_16136,N_16229);
and U17410 (N_17410,N_16316,N_16475);
xnor U17411 (N_17411,N_16583,N_16747);
xnor U17412 (N_17412,N_16471,N_16784);
or U17413 (N_17413,N_16520,N_16359);
xnor U17414 (N_17414,N_16466,N_16291);
or U17415 (N_17415,N_16108,N_16531);
nor U17416 (N_17416,N_16704,N_16421);
nand U17417 (N_17417,N_16553,N_16413);
and U17418 (N_17418,N_16524,N_16711);
nand U17419 (N_17419,N_16495,N_16509);
and U17420 (N_17420,N_16094,N_16100);
nor U17421 (N_17421,N_16184,N_16375);
and U17422 (N_17422,N_16376,N_16588);
nand U17423 (N_17423,N_16294,N_16684);
nor U17424 (N_17424,N_16369,N_16306);
nand U17425 (N_17425,N_16278,N_16742);
nand U17426 (N_17426,N_16234,N_16630);
xor U17427 (N_17427,N_16425,N_16729);
nand U17428 (N_17428,N_16528,N_16135);
xnor U17429 (N_17429,N_16317,N_16671);
nand U17430 (N_17430,N_16543,N_16080);
nand U17431 (N_17431,N_16517,N_16467);
or U17432 (N_17432,N_16574,N_16092);
xor U17433 (N_17433,N_16292,N_16023);
nor U17434 (N_17434,N_16553,N_16208);
nor U17435 (N_17435,N_16179,N_16052);
and U17436 (N_17436,N_16585,N_16195);
nand U17437 (N_17437,N_16051,N_16455);
nand U17438 (N_17438,N_16399,N_16101);
and U17439 (N_17439,N_16603,N_16672);
nand U17440 (N_17440,N_16731,N_16205);
xor U17441 (N_17441,N_16197,N_16235);
and U17442 (N_17442,N_16754,N_16109);
xnor U17443 (N_17443,N_16026,N_16301);
nand U17444 (N_17444,N_16004,N_16557);
or U17445 (N_17445,N_16094,N_16289);
nand U17446 (N_17446,N_16030,N_16620);
nor U17447 (N_17447,N_16114,N_16786);
nor U17448 (N_17448,N_16733,N_16302);
nor U17449 (N_17449,N_16761,N_16742);
xnor U17450 (N_17450,N_16234,N_16442);
nor U17451 (N_17451,N_16259,N_16388);
or U17452 (N_17452,N_16178,N_16525);
nor U17453 (N_17453,N_16771,N_16779);
nor U17454 (N_17454,N_16452,N_16289);
and U17455 (N_17455,N_16534,N_16781);
nand U17456 (N_17456,N_16271,N_16411);
and U17457 (N_17457,N_16596,N_16482);
or U17458 (N_17458,N_16222,N_16404);
nor U17459 (N_17459,N_16433,N_16635);
and U17460 (N_17460,N_16108,N_16513);
nor U17461 (N_17461,N_16107,N_16783);
xor U17462 (N_17462,N_16075,N_16579);
and U17463 (N_17463,N_16222,N_16349);
nand U17464 (N_17464,N_16251,N_16072);
nand U17465 (N_17465,N_16119,N_16345);
nand U17466 (N_17466,N_16661,N_16422);
nand U17467 (N_17467,N_16721,N_16172);
and U17468 (N_17468,N_16337,N_16765);
nor U17469 (N_17469,N_16075,N_16409);
nor U17470 (N_17470,N_16473,N_16794);
and U17471 (N_17471,N_16254,N_16026);
nand U17472 (N_17472,N_16245,N_16411);
xnor U17473 (N_17473,N_16112,N_16052);
and U17474 (N_17474,N_16365,N_16649);
and U17475 (N_17475,N_16478,N_16302);
nand U17476 (N_17476,N_16263,N_16383);
nor U17477 (N_17477,N_16092,N_16624);
and U17478 (N_17478,N_16571,N_16255);
or U17479 (N_17479,N_16647,N_16497);
nor U17480 (N_17480,N_16338,N_16763);
nand U17481 (N_17481,N_16798,N_16450);
and U17482 (N_17482,N_16655,N_16337);
and U17483 (N_17483,N_16270,N_16485);
xor U17484 (N_17484,N_16600,N_16052);
xor U17485 (N_17485,N_16293,N_16727);
or U17486 (N_17486,N_16167,N_16543);
nor U17487 (N_17487,N_16586,N_16238);
and U17488 (N_17488,N_16263,N_16066);
xnor U17489 (N_17489,N_16745,N_16162);
and U17490 (N_17490,N_16080,N_16607);
xor U17491 (N_17491,N_16024,N_16754);
or U17492 (N_17492,N_16715,N_16662);
nand U17493 (N_17493,N_16121,N_16779);
xnor U17494 (N_17494,N_16348,N_16599);
xor U17495 (N_17495,N_16614,N_16003);
nand U17496 (N_17496,N_16478,N_16343);
or U17497 (N_17497,N_16469,N_16528);
nor U17498 (N_17498,N_16157,N_16336);
nor U17499 (N_17499,N_16650,N_16696);
nor U17500 (N_17500,N_16547,N_16393);
xnor U17501 (N_17501,N_16085,N_16199);
nor U17502 (N_17502,N_16474,N_16174);
and U17503 (N_17503,N_16072,N_16215);
and U17504 (N_17504,N_16326,N_16539);
nor U17505 (N_17505,N_16197,N_16103);
or U17506 (N_17506,N_16639,N_16655);
and U17507 (N_17507,N_16280,N_16014);
and U17508 (N_17508,N_16704,N_16774);
nor U17509 (N_17509,N_16625,N_16705);
nand U17510 (N_17510,N_16720,N_16786);
nor U17511 (N_17511,N_16217,N_16568);
xnor U17512 (N_17512,N_16542,N_16241);
and U17513 (N_17513,N_16656,N_16170);
or U17514 (N_17514,N_16039,N_16178);
nand U17515 (N_17515,N_16616,N_16085);
and U17516 (N_17516,N_16663,N_16305);
xnor U17517 (N_17517,N_16731,N_16290);
nand U17518 (N_17518,N_16356,N_16263);
nand U17519 (N_17519,N_16232,N_16787);
or U17520 (N_17520,N_16197,N_16132);
nand U17521 (N_17521,N_16167,N_16648);
and U17522 (N_17522,N_16169,N_16637);
xor U17523 (N_17523,N_16510,N_16102);
xnor U17524 (N_17524,N_16748,N_16666);
nand U17525 (N_17525,N_16189,N_16107);
and U17526 (N_17526,N_16511,N_16230);
xor U17527 (N_17527,N_16200,N_16541);
and U17528 (N_17528,N_16657,N_16554);
nor U17529 (N_17529,N_16167,N_16281);
nor U17530 (N_17530,N_16109,N_16612);
nand U17531 (N_17531,N_16335,N_16346);
xnor U17532 (N_17532,N_16465,N_16159);
xor U17533 (N_17533,N_16665,N_16681);
nor U17534 (N_17534,N_16466,N_16449);
nor U17535 (N_17535,N_16133,N_16787);
nand U17536 (N_17536,N_16787,N_16087);
xor U17537 (N_17537,N_16582,N_16418);
nor U17538 (N_17538,N_16542,N_16453);
xor U17539 (N_17539,N_16140,N_16381);
xnor U17540 (N_17540,N_16441,N_16577);
and U17541 (N_17541,N_16382,N_16650);
and U17542 (N_17542,N_16562,N_16534);
and U17543 (N_17543,N_16149,N_16597);
nor U17544 (N_17544,N_16767,N_16659);
and U17545 (N_17545,N_16687,N_16576);
and U17546 (N_17546,N_16077,N_16123);
or U17547 (N_17547,N_16225,N_16283);
nand U17548 (N_17548,N_16306,N_16401);
and U17549 (N_17549,N_16791,N_16400);
xor U17550 (N_17550,N_16674,N_16139);
xnor U17551 (N_17551,N_16112,N_16762);
xnor U17552 (N_17552,N_16080,N_16756);
nand U17553 (N_17553,N_16708,N_16009);
xor U17554 (N_17554,N_16268,N_16350);
xnor U17555 (N_17555,N_16479,N_16425);
nor U17556 (N_17556,N_16523,N_16487);
xnor U17557 (N_17557,N_16054,N_16109);
or U17558 (N_17558,N_16777,N_16532);
nor U17559 (N_17559,N_16085,N_16293);
and U17560 (N_17560,N_16328,N_16771);
nand U17561 (N_17561,N_16771,N_16729);
or U17562 (N_17562,N_16639,N_16288);
nor U17563 (N_17563,N_16487,N_16473);
or U17564 (N_17564,N_16343,N_16701);
nor U17565 (N_17565,N_16574,N_16202);
nand U17566 (N_17566,N_16277,N_16232);
and U17567 (N_17567,N_16575,N_16693);
xor U17568 (N_17568,N_16401,N_16342);
nand U17569 (N_17569,N_16693,N_16269);
or U17570 (N_17570,N_16371,N_16277);
or U17571 (N_17571,N_16084,N_16023);
or U17572 (N_17572,N_16387,N_16521);
nand U17573 (N_17573,N_16702,N_16700);
or U17574 (N_17574,N_16380,N_16144);
xnor U17575 (N_17575,N_16610,N_16138);
xor U17576 (N_17576,N_16447,N_16104);
and U17577 (N_17577,N_16085,N_16452);
or U17578 (N_17578,N_16181,N_16232);
and U17579 (N_17579,N_16481,N_16078);
nor U17580 (N_17580,N_16529,N_16430);
or U17581 (N_17581,N_16000,N_16361);
xnor U17582 (N_17582,N_16692,N_16248);
xnor U17583 (N_17583,N_16737,N_16743);
and U17584 (N_17584,N_16065,N_16344);
or U17585 (N_17585,N_16504,N_16668);
and U17586 (N_17586,N_16294,N_16364);
nor U17587 (N_17587,N_16274,N_16625);
and U17588 (N_17588,N_16576,N_16028);
and U17589 (N_17589,N_16395,N_16229);
nand U17590 (N_17590,N_16246,N_16639);
xor U17591 (N_17591,N_16209,N_16393);
nor U17592 (N_17592,N_16653,N_16227);
or U17593 (N_17593,N_16781,N_16064);
nor U17594 (N_17594,N_16534,N_16417);
nand U17595 (N_17595,N_16683,N_16126);
or U17596 (N_17596,N_16074,N_16745);
and U17597 (N_17597,N_16225,N_16304);
nand U17598 (N_17598,N_16588,N_16690);
nor U17599 (N_17599,N_16684,N_16062);
xnor U17600 (N_17600,N_16973,N_17173);
and U17601 (N_17601,N_17271,N_16972);
nor U17602 (N_17602,N_17163,N_17264);
or U17603 (N_17603,N_16872,N_17144);
xnor U17604 (N_17604,N_17090,N_17463);
nand U17605 (N_17605,N_17046,N_17143);
xnor U17606 (N_17606,N_17358,N_16804);
or U17607 (N_17607,N_17482,N_16809);
xnor U17608 (N_17608,N_17304,N_16948);
nand U17609 (N_17609,N_17330,N_17287);
nor U17610 (N_17610,N_17540,N_17479);
xnor U17611 (N_17611,N_16834,N_16824);
nor U17612 (N_17612,N_17322,N_17373);
or U17613 (N_17613,N_17275,N_16810);
and U17614 (N_17614,N_17132,N_16895);
nor U17615 (N_17615,N_17489,N_17177);
nand U17616 (N_17616,N_17546,N_17403);
nand U17617 (N_17617,N_17074,N_17566);
nand U17618 (N_17618,N_17051,N_17478);
and U17619 (N_17619,N_16969,N_16861);
nand U17620 (N_17620,N_17258,N_16996);
nor U17621 (N_17621,N_17099,N_16954);
and U17622 (N_17622,N_17563,N_17541);
xnor U17623 (N_17623,N_17102,N_17551);
xnor U17624 (N_17624,N_17187,N_17195);
nor U17625 (N_17625,N_17574,N_17005);
or U17626 (N_17626,N_17101,N_16800);
or U17627 (N_17627,N_17336,N_17146);
nand U17628 (N_17628,N_17383,N_17462);
nand U17629 (N_17629,N_17255,N_16841);
and U17630 (N_17630,N_17172,N_17218);
nand U17631 (N_17631,N_16874,N_16913);
and U17632 (N_17632,N_17485,N_16934);
or U17633 (N_17633,N_17039,N_17060);
nor U17634 (N_17634,N_17480,N_17184);
xor U17635 (N_17635,N_16967,N_17596);
xnor U17636 (N_17636,N_17130,N_17022);
xnor U17637 (N_17637,N_17376,N_17585);
nand U17638 (N_17638,N_17451,N_17023);
and U17639 (N_17639,N_17449,N_17538);
or U17640 (N_17640,N_16924,N_16981);
nand U17641 (N_17641,N_17424,N_17435);
nor U17642 (N_17642,N_17355,N_16887);
nand U17643 (N_17643,N_17512,N_17350);
or U17644 (N_17644,N_17242,N_17379);
or U17645 (N_17645,N_17018,N_16971);
nand U17646 (N_17646,N_17511,N_17515);
nor U17647 (N_17647,N_16878,N_16807);
or U17648 (N_17648,N_16937,N_17374);
nor U17649 (N_17649,N_17473,N_17138);
nand U17650 (N_17650,N_16905,N_17565);
and U17651 (N_17651,N_17158,N_17477);
xnor U17652 (N_17652,N_17085,N_17548);
and U17653 (N_17653,N_16904,N_16906);
xnor U17654 (N_17654,N_17237,N_17148);
or U17655 (N_17655,N_16833,N_17091);
nand U17656 (N_17656,N_17497,N_17211);
xnor U17657 (N_17657,N_17009,N_16994);
or U17658 (N_17658,N_16876,N_17442);
or U17659 (N_17659,N_16822,N_17028);
and U17660 (N_17660,N_17307,N_17153);
xnor U17661 (N_17661,N_17007,N_17209);
and U17662 (N_17662,N_17127,N_17407);
nor U17663 (N_17663,N_16858,N_17069);
or U17664 (N_17664,N_17554,N_17289);
and U17665 (N_17665,N_16916,N_17315);
or U17666 (N_17666,N_16839,N_17006);
nor U17667 (N_17667,N_17397,N_16982);
xnor U17668 (N_17668,N_16953,N_17351);
nand U17669 (N_17669,N_17308,N_16859);
nor U17670 (N_17670,N_16910,N_16952);
nor U17671 (N_17671,N_17096,N_17500);
nor U17672 (N_17672,N_17295,N_16988);
or U17673 (N_17673,N_17152,N_17254);
and U17674 (N_17674,N_16832,N_17415);
xnor U17675 (N_17675,N_16831,N_17530);
nor U17676 (N_17676,N_17243,N_17557);
and U17677 (N_17677,N_16873,N_17579);
xor U17678 (N_17678,N_17213,N_17589);
nand U17679 (N_17679,N_16976,N_17320);
and U17680 (N_17680,N_17398,N_16815);
nor U17681 (N_17681,N_17492,N_17290);
or U17682 (N_17682,N_17133,N_17265);
nor U17683 (N_17683,N_17468,N_17079);
nand U17684 (N_17684,N_17576,N_17520);
and U17685 (N_17685,N_17142,N_16984);
xor U17686 (N_17686,N_16880,N_16978);
nor U17687 (N_17687,N_17252,N_16902);
nor U17688 (N_17688,N_16914,N_17278);
nor U17689 (N_17689,N_17418,N_16957);
nor U17690 (N_17690,N_17454,N_17444);
and U17691 (N_17691,N_16935,N_17274);
or U17692 (N_17692,N_17529,N_17334);
xnor U17693 (N_17693,N_17422,N_17168);
or U17694 (N_17694,N_17131,N_16977);
nand U17695 (N_17695,N_17030,N_16899);
and U17696 (N_17696,N_17077,N_17537);
and U17697 (N_17697,N_17333,N_16802);
nor U17698 (N_17698,N_17120,N_17081);
xnor U17699 (N_17699,N_17276,N_17447);
nor U17700 (N_17700,N_16854,N_16888);
xor U17701 (N_17701,N_17460,N_17450);
and U17702 (N_17702,N_17321,N_16927);
nand U17703 (N_17703,N_16845,N_17409);
nor U17704 (N_17704,N_17327,N_17516);
and U17705 (N_17705,N_17441,N_17391);
xor U17706 (N_17706,N_17001,N_17395);
and U17707 (N_17707,N_16816,N_17000);
or U17708 (N_17708,N_17103,N_16860);
nor U17709 (N_17709,N_17393,N_17134);
nand U17710 (N_17710,N_17509,N_17584);
or U17711 (N_17711,N_16985,N_16947);
and U17712 (N_17712,N_17228,N_17093);
xnor U17713 (N_17713,N_17065,N_16817);
or U17714 (N_17714,N_16922,N_17588);
and U17715 (N_17715,N_17371,N_17408);
or U17716 (N_17716,N_17021,N_17149);
nand U17717 (N_17717,N_17410,N_17340);
nor U17718 (N_17718,N_16979,N_17201);
nand U17719 (N_17719,N_16882,N_17224);
and U17720 (N_17720,N_17019,N_16930);
and U17721 (N_17721,N_16938,N_17517);
and U17722 (N_17722,N_17439,N_17121);
and U17723 (N_17723,N_17286,N_16819);
nand U17724 (N_17724,N_17270,N_17108);
or U17725 (N_17725,N_16852,N_17285);
and U17726 (N_17726,N_17034,N_16875);
and U17727 (N_17727,N_16912,N_17191);
nand U17728 (N_17728,N_17421,N_17216);
or U17729 (N_17729,N_17481,N_16945);
nor U17730 (N_17730,N_17362,N_17543);
and U17731 (N_17731,N_16950,N_17032);
nor U17732 (N_17732,N_17491,N_17200);
and U17733 (N_17733,N_16961,N_17110);
nor U17734 (N_17734,N_16885,N_17113);
or U17735 (N_17735,N_17140,N_17125);
nand U17736 (N_17736,N_16840,N_16964);
or U17737 (N_17737,N_16829,N_17573);
nand U17738 (N_17738,N_17331,N_17488);
xnor U17739 (N_17739,N_17292,N_17220);
and U17740 (N_17740,N_17354,N_17202);
nor U17741 (N_17741,N_17236,N_16806);
or U17742 (N_17742,N_17135,N_17183);
xnor U17743 (N_17743,N_17305,N_17267);
nand U17744 (N_17744,N_17319,N_17083);
xnor U17745 (N_17745,N_17159,N_17377);
nor U17746 (N_17746,N_17461,N_16986);
or U17747 (N_17747,N_17426,N_16932);
nor U17748 (N_17748,N_17370,N_17024);
and U17749 (N_17749,N_16907,N_17219);
and U17750 (N_17750,N_17229,N_17094);
or U17751 (N_17751,N_17151,N_17343);
nand U17752 (N_17752,N_17273,N_16863);
nor U17753 (N_17753,N_17555,N_17561);
nand U17754 (N_17754,N_17298,N_17569);
nor U17755 (N_17755,N_16818,N_17396);
xor U17756 (N_17756,N_16987,N_16933);
or U17757 (N_17757,N_17437,N_17082);
or U17758 (N_17758,N_16812,N_17367);
xor U17759 (N_17759,N_17232,N_16866);
nor U17760 (N_17760,N_17076,N_16893);
nor U17761 (N_17761,N_17198,N_17595);
nand U17762 (N_17762,N_17197,N_17507);
or U17763 (N_17763,N_17423,N_17339);
xnor U17764 (N_17764,N_17075,N_17325);
and U17765 (N_17765,N_17095,N_17414);
nor U17766 (N_17766,N_17510,N_17235);
nor U17767 (N_17767,N_17549,N_17189);
nor U17768 (N_17768,N_17136,N_16856);
xor U17769 (N_17769,N_17092,N_17524);
and U17770 (N_17770,N_16993,N_17050);
or U17771 (N_17771,N_16843,N_16963);
xnor U17772 (N_17772,N_17059,N_16917);
or U17773 (N_17773,N_17470,N_16825);
and U17774 (N_17774,N_17513,N_17244);
nor U17775 (N_17775,N_17313,N_17472);
or U17776 (N_17776,N_17361,N_17378);
nor U17777 (N_17777,N_17227,N_17586);
xnor U17778 (N_17778,N_17086,N_17073);
xnor U17779 (N_17779,N_17487,N_16920);
xnor U17780 (N_17780,N_17057,N_17544);
nand U17781 (N_17781,N_16915,N_17126);
nor U17782 (N_17782,N_17432,N_17049);
nor U17783 (N_17783,N_17160,N_17128);
or U17784 (N_17784,N_17257,N_16928);
and U17785 (N_17785,N_17471,N_17453);
and U17786 (N_17786,N_17337,N_17411);
nor U17787 (N_17787,N_17031,N_16966);
nand U17788 (N_17788,N_16814,N_17518);
and U17789 (N_17789,N_17154,N_17427);
nand U17790 (N_17790,N_17003,N_17545);
nand U17791 (N_17791,N_17014,N_17053);
xor U17792 (N_17792,N_17192,N_17582);
xor U17793 (N_17793,N_17210,N_17259);
or U17794 (N_17794,N_16997,N_16908);
xor U17795 (N_17795,N_17416,N_17360);
xor U17796 (N_17796,N_17583,N_17266);
or U17797 (N_17797,N_17328,N_16879);
xor U17798 (N_17798,N_16853,N_16886);
and U17799 (N_17799,N_17332,N_17015);
xor U17800 (N_17800,N_16965,N_17147);
nor U17801 (N_17801,N_17483,N_16921);
nor U17802 (N_17802,N_17277,N_17250);
and U17803 (N_17803,N_17348,N_17498);
or U17804 (N_17804,N_17240,N_17591);
or U17805 (N_17805,N_16869,N_17139);
xnor U17806 (N_17806,N_17346,N_17458);
nor U17807 (N_17807,N_17186,N_16944);
or U17808 (N_17808,N_17193,N_17314);
and U17809 (N_17809,N_17288,N_17533);
and U17810 (N_17810,N_17041,N_16865);
and U17811 (N_17811,N_17245,N_17317);
and U17812 (N_17812,N_16942,N_17100);
nand U17813 (N_17813,N_16889,N_17388);
xor U17814 (N_17814,N_17519,N_16868);
nand U17815 (N_17815,N_17112,N_17026);
xnor U17816 (N_17816,N_17114,N_17347);
xor U17817 (N_17817,N_17047,N_17523);
and U17818 (N_17818,N_17353,N_16951);
nor U17819 (N_17819,N_17419,N_17587);
and U17820 (N_17820,N_17067,N_17299);
nor U17821 (N_17821,N_17206,N_17562);
and U17822 (N_17822,N_17029,N_17556);
or U17823 (N_17823,N_17056,N_17020);
nor U17824 (N_17824,N_17011,N_17558);
or U17825 (N_17825,N_17063,N_17469);
nand U17826 (N_17826,N_17098,N_17078);
and U17827 (N_17827,N_17045,N_17580);
and U17828 (N_17828,N_17542,N_17165);
or U17829 (N_17829,N_16890,N_17593);
or U17830 (N_17830,N_17180,N_17399);
nor U17831 (N_17831,N_16960,N_17522);
xnor U17832 (N_17832,N_17214,N_17311);
and U17833 (N_17833,N_17465,N_17107);
xor U17834 (N_17834,N_17207,N_16884);
or U17835 (N_17835,N_17221,N_17064);
or U17836 (N_17836,N_17428,N_17035);
nor U17837 (N_17837,N_17440,N_17089);
nand U17838 (N_17838,N_17294,N_16980);
nor U17839 (N_17839,N_17455,N_17230);
or U17840 (N_17840,N_17404,N_17043);
and U17841 (N_17841,N_16974,N_16999);
xor U17842 (N_17842,N_17446,N_16983);
nor U17843 (N_17843,N_17166,N_16862);
xor U17844 (N_17844,N_17156,N_17246);
xor U17845 (N_17845,N_17306,N_17284);
nor U17846 (N_17846,N_16801,N_17526);
or U17847 (N_17847,N_16842,N_17002);
and U17848 (N_17848,N_16990,N_17162);
and U17849 (N_17849,N_17592,N_17316);
or U17850 (N_17850,N_17429,N_17532);
nor U17851 (N_17851,N_17194,N_16975);
nand U17852 (N_17852,N_16992,N_17417);
and U17853 (N_17853,N_17301,N_17369);
and U17854 (N_17854,N_17217,N_17155);
and U17855 (N_17855,N_17495,N_17326);
xor U17856 (N_17856,N_17502,N_17575);
or U17857 (N_17857,N_17445,N_17400);
and U17858 (N_17858,N_17312,N_17384);
nor U17859 (N_17859,N_17234,N_17071);
nor U17860 (N_17860,N_17072,N_17375);
or U17861 (N_17861,N_17190,N_17027);
nand U17862 (N_17862,N_17150,N_16837);
xnor U17863 (N_17863,N_17486,N_17534);
or U17864 (N_17864,N_17256,N_17042);
xnor U17865 (N_17865,N_17356,N_17223);
xor U17866 (N_17866,N_16813,N_16919);
nor U17867 (N_17867,N_17084,N_17282);
xnor U17868 (N_17868,N_17323,N_16939);
and U17869 (N_17869,N_17283,N_16943);
nand U17870 (N_17870,N_16958,N_17341);
and U17871 (N_17871,N_17061,N_17318);
nor U17872 (N_17872,N_17268,N_16898);
or U17873 (N_17873,N_16956,N_16826);
nand U17874 (N_17874,N_17203,N_16864);
and U17875 (N_17875,N_17413,N_16896);
and U17876 (N_17876,N_17436,N_16883);
or U17877 (N_17877,N_16946,N_17357);
or U17878 (N_17878,N_17590,N_17233);
and U17879 (N_17879,N_17247,N_16835);
xor U17880 (N_17880,N_17279,N_17122);
xor U17881 (N_17881,N_17116,N_17037);
nor U17882 (N_17882,N_17205,N_17179);
and U17883 (N_17883,N_17297,N_17597);
or U17884 (N_17884,N_17238,N_17044);
and U17885 (N_17885,N_17560,N_17559);
xor U17886 (N_17886,N_17536,N_17004);
nor U17887 (N_17887,N_16929,N_17598);
and U17888 (N_17888,N_17309,N_17188);
xor U17889 (N_17889,N_17387,N_17010);
xor U17890 (N_17890,N_17302,N_17364);
nand U17891 (N_17891,N_17109,N_17017);
and U17892 (N_17892,N_17503,N_17484);
nand U17893 (N_17893,N_17070,N_17272);
nor U17894 (N_17894,N_17553,N_17514);
xor U17895 (N_17895,N_16998,N_17452);
or U17896 (N_17896,N_17296,N_17448);
or U17897 (N_17897,N_16830,N_16836);
nor U17898 (N_17898,N_17363,N_16847);
nor U17899 (N_17899,N_16846,N_17300);
nor U17900 (N_17900,N_16897,N_17594);
or U17901 (N_17901,N_16891,N_17506);
nand U17902 (N_17902,N_17199,N_17171);
nor U17903 (N_17903,N_16970,N_17459);
nand U17904 (N_17904,N_17547,N_16991);
xor U17905 (N_17905,N_16808,N_17366);
and U17906 (N_17906,N_17124,N_17345);
nand U17907 (N_17907,N_16940,N_17161);
nand U17908 (N_17908,N_17251,N_17389);
nand U17909 (N_17909,N_17344,N_16962);
or U17910 (N_17910,N_16941,N_17476);
and U17911 (N_17911,N_16949,N_17496);
nor U17912 (N_17912,N_17467,N_17386);
and U17913 (N_17913,N_17040,N_17572);
nor U17914 (N_17914,N_17392,N_16838);
nand U17915 (N_17915,N_17382,N_17385);
and U17916 (N_17916,N_17182,N_17204);
nor U17917 (N_17917,N_16823,N_17381);
xor U17918 (N_17918,N_17303,N_17431);
or U17919 (N_17919,N_16857,N_17550);
and U17920 (N_17920,N_17349,N_17434);
and U17921 (N_17921,N_17280,N_16894);
nand U17922 (N_17922,N_17525,N_17420);
or U17923 (N_17923,N_16881,N_17401);
nand U17924 (N_17924,N_17490,N_17062);
nand U17925 (N_17925,N_17215,N_16892);
and U17926 (N_17926,N_17038,N_16820);
and U17927 (N_17927,N_17260,N_16900);
and U17928 (N_17928,N_17170,N_17008);
xor U17929 (N_17929,N_17066,N_17368);
nor U17930 (N_17930,N_17338,N_17464);
xor U17931 (N_17931,N_17164,N_17571);
or U17932 (N_17932,N_17552,N_17406);
nor U17933 (N_17933,N_17352,N_17058);
nor U17934 (N_17934,N_16821,N_16870);
xnor U17935 (N_17935,N_17225,N_17466);
xor U17936 (N_17936,N_17111,N_16968);
and U17937 (N_17937,N_17178,N_16803);
nor U17938 (N_17938,N_17068,N_17438);
nand U17939 (N_17939,N_16959,N_17145);
nor U17940 (N_17940,N_16855,N_17539);
and U17941 (N_17941,N_17527,N_17425);
nand U17942 (N_17942,N_16931,N_17174);
nand U17943 (N_17943,N_16877,N_17185);
xor U17944 (N_17944,N_17493,N_17141);
or U17945 (N_17945,N_17097,N_17106);
xnor U17946 (N_17946,N_17105,N_16995);
and U17947 (N_17947,N_17248,N_17036);
or U17948 (N_17948,N_17504,N_17016);
nor U17949 (N_17949,N_17167,N_17335);
nor U17950 (N_17950,N_17531,N_16936);
and U17951 (N_17951,N_17430,N_17443);
xnor U17952 (N_17952,N_17117,N_17054);
nor U17953 (N_17953,N_17499,N_17599);
nand U17954 (N_17954,N_17013,N_17380);
or U17955 (N_17955,N_17433,N_17474);
and U17956 (N_17956,N_17261,N_17521);
or U17957 (N_17957,N_17025,N_17269);
and U17958 (N_17958,N_16909,N_17329);
and U17959 (N_17959,N_17342,N_17087);
and U17960 (N_17960,N_17157,N_16903);
nor U17961 (N_17961,N_17222,N_17281);
nor U17962 (N_17962,N_17055,N_17115);
xor U17963 (N_17963,N_16805,N_17196);
and U17964 (N_17964,N_17372,N_17365);
xnor U17965 (N_17965,N_17263,N_16851);
xnor U17966 (N_17966,N_17475,N_17457);
nor U17967 (N_17967,N_16871,N_17505);
nor U17968 (N_17968,N_17137,N_17119);
nand U17969 (N_17969,N_16925,N_17048);
and U17970 (N_17970,N_17129,N_17412);
nand U17971 (N_17971,N_17359,N_17567);
nor U17972 (N_17972,N_16955,N_17528);
or U17973 (N_17973,N_16848,N_17262);
and U17974 (N_17974,N_17581,N_17231);
nor U17975 (N_17975,N_16811,N_17176);
and U17976 (N_17976,N_16918,N_17578);
xnor U17977 (N_17977,N_17104,N_17570);
and U17978 (N_17978,N_17175,N_16901);
nand U17979 (N_17979,N_17501,N_17181);
or U17980 (N_17980,N_16850,N_17249);
xor U17981 (N_17981,N_17402,N_17118);
or U17982 (N_17982,N_17293,N_17088);
nor U17983 (N_17983,N_17208,N_16911);
nand U17984 (N_17984,N_16828,N_17212);
nor U17985 (N_17985,N_17123,N_16867);
nor U17986 (N_17986,N_17405,N_17239);
nor U17987 (N_17987,N_17012,N_16849);
and U17988 (N_17988,N_16989,N_17535);
xnor U17989 (N_17989,N_17394,N_17253);
or U17990 (N_17990,N_17324,N_17456);
xnor U17991 (N_17991,N_17033,N_16827);
nor U17992 (N_17992,N_17226,N_16926);
or U17993 (N_17993,N_17291,N_17080);
nand U17994 (N_17994,N_17577,N_17169);
xor U17995 (N_17995,N_17568,N_17494);
or U17996 (N_17996,N_16844,N_16923);
xnor U17997 (N_17997,N_17564,N_17241);
nor U17998 (N_17998,N_17052,N_17508);
xnor U17999 (N_17999,N_17310,N_17390);
nor U18000 (N_18000,N_17323,N_17322);
and U18001 (N_18001,N_17053,N_16886);
or U18002 (N_18002,N_17438,N_16844);
nor U18003 (N_18003,N_17022,N_16911);
nor U18004 (N_18004,N_16993,N_17051);
or U18005 (N_18005,N_17364,N_17159);
nand U18006 (N_18006,N_17333,N_17296);
nor U18007 (N_18007,N_16849,N_16888);
nor U18008 (N_18008,N_17310,N_17108);
xnor U18009 (N_18009,N_16805,N_17198);
or U18010 (N_18010,N_16981,N_16827);
and U18011 (N_18011,N_17047,N_17073);
or U18012 (N_18012,N_17135,N_16869);
xnor U18013 (N_18013,N_16851,N_17415);
or U18014 (N_18014,N_16848,N_17364);
nor U18015 (N_18015,N_16885,N_17203);
or U18016 (N_18016,N_17445,N_17279);
and U18017 (N_18017,N_17043,N_16997);
nor U18018 (N_18018,N_17393,N_17213);
and U18019 (N_18019,N_17077,N_17040);
xnor U18020 (N_18020,N_17504,N_17385);
nor U18021 (N_18021,N_17191,N_16875);
nand U18022 (N_18022,N_17411,N_16912);
and U18023 (N_18023,N_17127,N_17463);
and U18024 (N_18024,N_17074,N_17184);
or U18025 (N_18025,N_16876,N_16861);
xor U18026 (N_18026,N_17370,N_17571);
nand U18027 (N_18027,N_17332,N_17132);
or U18028 (N_18028,N_16957,N_16803);
xnor U18029 (N_18029,N_16984,N_17478);
nor U18030 (N_18030,N_17156,N_17371);
nor U18031 (N_18031,N_16852,N_17500);
nor U18032 (N_18032,N_17277,N_16863);
and U18033 (N_18033,N_16974,N_17036);
nand U18034 (N_18034,N_16992,N_16800);
xnor U18035 (N_18035,N_17336,N_16861);
nand U18036 (N_18036,N_16830,N_16947);
xnor U18037 (N_18037,N_17532,N_17370);
xnor U18038 (N_18038,N_17373,N_17501);
or U18039 (N_18039,N_17090,N_16914);
xor U18040 (N_18040,N_17415,N_17109);
and U18041 (N_18041,N_17373,N_17090);
xor U18042 (N_18042,N_17368,N_17400);
or U18043 (N_18043,N_17536,N_17455);
and U18044 (N_18044,N_17283,N_17085);
nand U18045 (N_18045,N_16878,N_17430);
or U18046 (N_18046,N_16865,N_17465);
and U18047 (N_18047,N_17282,N_17395);
nor U18048 (N_18048,N_17087,N_16896);
nand U18049 (N_18049,N_17491,N_17097);
nand U18050 (N_18050,N_17253,N_17166);
or U18051 (N_18051,N_17116,N_17007);
xor U18052 (N_18052,N_16913,N_17024);
or U18053 (N_18053,N_16903,N_17207);
nor U18054 (N_18054,N_17441,N_16870);
or U18055 (N_18055,N_17112,N_17246);
and U18056 (N_18056,N_17102,N_16813);
and U18057 (N_18057,N_17162,N_17543);
xor U18058 (N_18058,N_17596,N_16970);
or U18059 (N_18059,N_17423,N_17455);
and U18060 (N_18060,N_17340,N_17393);
nand U18061 (N_18061,N_17550,N_16890);
nor U18062 (N_18062,N_16819,N_17579);
or U18063 (N_18063,N_17345,N_17293);
nand U18064 (N_18064,N_17218,N_16935);
or U18065 (N_18065,N_16882,N_17385);
nand U18066 (N_18066,N_17000,N_17370);
and U18067 (N_18067,N_17262,N_16985);
and U18068 (N_18068,N_17518,N_17323);
and U18069 (N_18069,N_16898,N_16889);
nor U18070 (N_18070,N_17231,N_16996);
nor U18071 (N_18071,N_17205,N_17326);
xor U18072 (N_18072,N_17555,N_17061);
or U18073 (N_18073,N_16988,N_16803);
and U18074 (N_18074,N_17437,N_17025);
and U18075 (N_18075,N_17447,N_16888);
and U18076 (N_18076,N_16800,N_16933);
or U18077 (N_18077,N_16852,N_16933);
nor U18078 (N_18078,N_17152,N_17104);
and U18079 (N_18079,N_17365,N_17345);
nand U18080 (N_18080,N_17065,N_16953);
xor U18081 (N_18081,N_17091,N_17505);
and U18082 (N_18082,N_16936,N_17227);
xor U18083 (N_18083,N_17016,N_16866);
or U18084 (N_18084,N_16919,N_17394);
nor U18085 (N_18085,N_17376,N_17225);
nor U18086 (N_18086,N_16881,N_17010);
nor U18087 (N_18087,N_17561,N_17129);
nand U18088 (N_18088,N_17203,N_17092);
nand U18089 (N_18089,N_17434,N_16994);
and U18090 (N_18090,N_17469,N_16825);
xor U18091 (N_18091,N_17276,N_17485);
and U18092 (N_18092,N_16993,N_17059);
nor U18093 (N_18093,N_17046,N_17544);
xnor U18094 (N_18094,N_17077,N_17129);
and U18095 (N_18095,N_17533,N_17391);
and U18096 (N_18096,N_17022,N_17209);
nand U18097 (N_18097,N_16821,N_17584);
nand U18098 (N_18098,N_17518,N_17006);
or U18099 (N_18099,N_17234,N_16904);
nor U18100 (N_18100,N_17230,N_17277);
nor U18101 (N_18101,N_17395,N_17440);
nor U18102 (N_18102,N_17135,N_17031);
nor U18103 (N_18103,N_16804,N_17167);
or U18104 (N_18104,N_17501,N_17334);
xnor U18105 (N_18105,N_16823,N_16990);
nand U18106 (N_18106,N_17235,N_17098);
and U18107 (N_18107,N_17214,N_16935);
xnor U18108 (N_18108,N_17177,N_17317);
nor U18109 (N_18109,N_17539,N_17052);
nor U18110 (N_18110,N_16849,N_17376);
or U18111 (N_18111,N_17299,N_17208);
and U18112 (N_18112,N_17044,N_17069);
or U18113 (N_18113,N_16823,N_17033);
or U18114 (N_18114,N_16917,N_17052);
nor U18115 (N_18115,N_17015,N_16972);
nor U18116 (N_18116,N_17132,N_16815);
nand U18117 (N_18117,N_17478,N_17277);
nand U18118 (N_18118,N_17040,N_17317);
nand U18119 (N_18119,N_17556,N_17067);
or U18120 (N_18120,N_17551,N_16907);
nand U18121 (N_18121,N_16922,N_17462);
xnor U18122 (N_18122,N_17189,N_16968);
and U18123 (N_18123,N_17456,N_17552);
nor U18124 (N_18124,N_17470,N_17209);
nand U18125 (N_18125,N_16930,N_16813);
and U18126 (N_18126,N_17493,N_16855);
nor U18127 (N_18127,N_17226,N_17139);
xnor U18128 (N_18128,N_17209,N_16879);
xor U18129 (N_18129,N_16921,N_17175);
or U18130 (N_18130,N_17457,N_16986);
or U18131 (N_18131,N_17477,N_16958);
and U18132 (N_18132,N_16834,N_16958);
and U18133 (N_18133,N_17302,N_17374);
nor U18134 (N_18134,N_17201,N_17574);
and U18135 (N_18135,N_16868,N_17213);
or U18136 (N_18136,N_17179,N_17599);
nor U18137 (N_18137,N_17456,N_16803);
and U18138 (N_18138,N_17112,N_17015);
and U18139 (N_18139,N_17298,N_17567);
nor U18140 (N_18140,N_17471,N_17555);
nand U18141 (N_18141,N_16826,N_16965);
nor U18142 (N_18142,N_17298,N_17419);
xnor U18143 (N_18143,N_17328,N_17134);
nor U18144 (N_18144,N_17518,N_17587);
nor U18145 (N_18145,N_16865,N_16873);
nand U18146 (N_18146,N_16980,N_17014);
nand U18147 (N_18147,N_17005,N_17111);
nand U18148 (N_18148,N_17026,N_17362);
nand U18149 (N_18149,N_17100,N_16873);
and U18150 (N_18150,N_17422,N_17033);
nand U18151 (N_18151,N_16933,N_16937);
and U18152 (N_18152,N_17195,N_17212);
xnor U18153 (N_18153,N_16805,N_16933);
nor U18154 (N_18154,N_17017,N_17521);
xnor U18155 (N_18155,N_17410,N_17543);
nand U18156 (N_18156,N_17302,N_17585);
xor U18157 (N_18157,N_16952,N_17127);
nand U18158 (N_18158,N_17335,N_17018);
nor U18159 (N_18159,N_17214,N_17370);
and U18160 (N_18160,N_17501,N_16981);
xnor U18161 (N_18161,N_17326,N_17150);
xor U18162 (N_18162,N_17038,N_17103);
nor U18163 (N_18163,N_17027,N_16985);
nor U18164 (N_18164,N_17503,N_17575);
nor U18165 (N_18165,N_17349,N_16815);
or U18166 (N_18166,N_17104,N_17463);
or U18167 (N_18167,N_16900,N_17266);
nor U18168 (N_18168,N_17026,N_17352);
and U18169 (N_18169,N_17327,N_16844);
nor U18170 (N_18170,N_17285,N_16975);
and U18171 (N_18171,N_17086,N_17112);
nand U18172 (N_18172,N_17401,N_17317);
nor U18173 (N_18173,N_17097,N_17129);
nand U18174 (N_18174,N_17312,N_17499);
and U18175 (N_18175,N_17052,N_17116);
and U18176 (N_18176,N_17104,N_17473);
xor U18177 (N_18177,N_17401,N_16924);
xor U18178 (N_18178,N_17574,N_17247);
or U18179 (N_18179,N_16970,N_17351);
nand U18180 (N_18180,N_17080,N_17501);
nand U18181 (N_18181,N_17360,N_16825);
and U18182 (N_18182,N_17377,N_17417);
nand U18183 (N_18183,N_16869,N_17045);
nand U18184 (N_18184,N_17234,N_17331);
nand U18185 (N_18185,N_16835,N_17179);
nor U18186 (N_18186,N_17261,N_17523);
and U18187 (N_18187,N_17575,N_17441);
xnor U18188 (N_18188,N_17218,N_17052);
xnor U18189 (N_18189,N_16819,N_17435);
or U18190 (N_18190,N_17513,N_17460);
nor U18191 (N_18191,N_17228,N_17213);
and U18192 (N_18192,N_16949,N_17071);
nor U18193 (N_18193,N_17384,N_17445);
or U18194 (N_18194,N_17047,N_17170);
nor U18195 (N_18195,N_17514,N_16996);
or U18196 (N_18196,N_17330,N_16828);
nor U18197 (N_18197,N_17210,N_17052);
or U18198 (N_18198,N_17267,N_17087);
nor U18199 (N_18199,N_17526,N_16968);
nand U18200 (N_18200,N_16879,N_17313);
and U18201 (N_18201,N_16823,N_17149);
and U18202 (N_18202,N_17053,N_17123);
or U18203 (N_18203,N_16952,N_16875);
nor U18204 (N_18204,N_17113,N_17531);
xor U18205 (N_18205,N_17268,N_17249);
nand U18206 (N_18206,N_17133,N_16994);
xor U18207 (N_18207,N_16873,N_17176);
or U18208 (N_18208,N_16963,N_16807);
nand U18209 (N_18209,N_17549,N_17236);
nand U18210 (N_18210,N_17434,N_17353);
nor U18211 (N_18211,N_16896,N_17381);
and U18212 (N_18212,N_17547,N_16988);
xor U18213 (N_18213,N_16889,N_16952);
nand U18214 (N_18214,N_17097,N_17130);
or U18215 (N_18215,N_17368,N_16996);
xor U18216 (N_18216,N_17401,N_16883);
or U18217 (N_18217,N_17146,N_17541);
or U18218 (N_18218,N_16869,N_17452);
and U18219 (N_18219,N_17243,N_17163);
nor U18220 (N_18220,N_17069,N_16978);
nor U18221 (N_18221,N_17006,N_17572);
nor U18222 (N_18222,N_16988,N_17501);
nor U18223 (N_18223,N_17146,N_17097);
xor U18224 (N_18224,N_17577,N_16982);
nor U18225 (N_18225,N_16963,N_17192);
or U18226 (N_18226,N_16818,N_16935);
nand U18227 (N_18227,N_17564,N_17263);
nand U18228 (N_18228,N_17535,N_17346);
nor U18229 (N_18229,N_17513,N_17387);
nor U18230 (N_18230,N_16947,N_17039);
and U18231 (N_18231,N_17518,N_17059);
xor U18232 (N_18232,N_17335,N_17340);
nor U18233 (N_18233,N_16912,N_17383);
nor U18234 (N_18234,N_17195,N_16982);
and U18235 (N_18235,N_17412,N_16927);
and U18236 (N_18236,N_17211,N_17116);
xnor U18237 (N_18237,N_17578,N_17328);
or U18238 (N_18238,N_17337,N_17540);
nor U18239 (N_18239,N_17395,N_16805);
nor U18240 (N_18240,N_17557,N_17260);
or U18241 (N_18241,N_17531,N_16975);
or U18242 (N_18242,N_17043,N_16934);
xnor U18243 (N_18243,N_17180,N_17148);
or U18244 (N_18244,N_16895,N_16890);
or U18245 (N_18245,N_17353,N_17264);
or U18246 (N_18246,N_17293,N_17538);
and U18247 (N_18247,N_17066,N_17173);
nand U18248 (N_18248,N_17208,N_16949);
nor U18249 (N_18249,N_16865,N_17116);
nand U18250 (N_18250,N_17578,N_17275);
and U18251 (N_18251,N_17410,N_17425);
xnor U18252 (N_18252,N_17257,N_16890);
nor U18253 (N_18253,N_17033,N_17301);
or U18254 (N_18254,N_16977,N_17183);
nand U18255 (N_18255,N_17103,N_17338);
xor U18256 (N_18256,N_17180,N_17104);
or U18257 (N_18257,N_16933,N_16801);
and U18258 (N_18258,N_17411,N_16838);
nor U18259 (N_18259,N_17137,N_17179);
and U18260 (N_18260,N_17016,N_17014);
and U18261 (N_18261,N_17388,N_17281);
xor U18262 (N_18262,N_17421,N_17109);
xor U18263 (N_18263,N_16917,N_17160);
nand U18264 (N_18264,N_16859,N_17169);
nand U18265 (N_18265,N_16888,N_17192);
xnor U18266 (N_18266,N_16834,N_17027);
xnor U18267 (N_18267,N_17063,N_16864);
or U18268 (N_18268,N_16969,N_16999);
and U18269 (N_18269,N_17037,N_17561);
or U18270 (N_18270,N_17581,N_17161);
and U18271 (N_18271,N_17271,N_16873);
and U18272 (N_18272,N_17318,N_17052);
or U18273 (N_18273,N_16931,N_17378);
or U18274 (N_18274,N_17186,N_17125);
xor U18275 (N_18275,N_16909,N_17444);
or U18276 (N_18276,N_17439,N_17365);
nand U18277 (N_18277,N_16856,N_17322);
xnor U18278 (N_18278,N_17144,N_17563);
or U18279 (N_18279,N_16947,N_17017);
nand U18280 (N_18280,N_17579,N_17450);
nor U18281 (N_18281,N_17101,N_17053);
nand U18282 (N_18282,N_17254,N_17083);
or U18283 (N_18283,N_17303,N_16902);
xnor U18284 (N_18284,N_17004,N_17141);
and U18285 (N_18285,N_16959,N_17165);
nor U18286 (N_18286,N_17129,N_17192);
or U18287 (N_18287,N_17212,N_17583);
nor U18288 (N_18288,N_17384,N_17299);
nand U18289 (N_18289,N_16902,N_16917);
or U18290 (N_18290,N_16859,N_17149);
and U18291 (N_18291,N_17397,N_16933);
xnor U18292 (N_18292,N_16909,N_17486);
xnor U18293 (N_18293,N_17017,N_17270);
and U18294 (N_18294,N_17487,N_17261);
or U18295 (N_18295,N_16897,N_17570);
and U18296 (N_18296,N_17158,N_17390);
nor U18297 (N_18297,N_16835,N_17281);
nand U18298 (N_18298,N_16912,N_16853);
nand U18299 (N_18299,N_17206,N_16807);
xnor U18300 (N_18300,N_17365,N_17352);
and U18301 (N_18301,N_16881,N_17295);
nand U18302 (N_18302,N_16951,N_17277);
nand U18303 (N_18303,N_17090,N_17065);
or U18304 (N_18304,N_17552,N_17277);
and U18305 (N_18305,N_17245,N_17365);
xor U18306 (N_18306,N_17434,N_17559);
and U18307 (N_18307,N_17382,N_17422);
xnor U18308 (N_18308,N_17441,N_17539);
xnor U18309 (N_18309,N_17447,N_17576);
nand U18310 (N_18310,N_17418,N_17156);
nor U18311 (N_18311,N_17161,N_16938);
nor U18312 (N_18312,N_17117,N_17139);
or U18313 (N_18313,N_16875,N_16909);
nand U18314 (N_18314,N_17010,N_17511);
and U18315 (N_18315,N_16918,N_16953);
nand U18316 (N_18316,N_17261,N_17060);
nor U18317 (N_18317,N_17459,N_16911);
and U18318 (N_18318,N_17098,N_17219);
or U18319 (N_18319,N_16872,N_16965);
nand U18320 (N_18320,N_17517,N_17143);
nand U18321 (N_18321,N_16821,N_17060);
xor U18322 (N_18322,N_16959,N_17060);
and U18323 (N_18323,N_17039,N_16930);
xnor U18324 (N_18324,N_17295,N_16980);
nor U18325 (N_18325,N_17103,N_17284);
xnor U18326 (N_18326,N_17113,N_17416);
xor U18327 (N_18327,N_17242,N_17517);
nor U18328 (N_18328,N_17320,N_17546);
or U18329 (N_18329,N_17246,N_17175);
nand U18330 (N_18330,N_17046,N_17368);
nor U18331 (N_18331,N_16908,N_17469);
and U18332 (N_18332,N_16815,N_17081);
xnor U18333 (N_18333,N_17403,N_17533);
nor U18334 (N_18334,N_17138,N_17381);
and U18335 (N_18335,N_17005,N_17476);
nand U18336 (N_18336,N_17531,N_16858);
or U18337 (N_18337,N_16974,N_17370);
nor U18338 (N_18338,N_17069,N_17462);
or U18339 (N_18339,N_16903,N_17260);
xnor U18340 (N_18340,N_17046,N_17454);
nand U18341 (N_18341,N_16848,N_17050);
xnor U18342 (N_18342,N_17324,N_17566);
nor U18343 (N_18343,N_17015,N_17049);
nand U18344 (N_18344,N_17471,N_17392);
or U18345 (N_18345,N_17124,N_17238);
and U18346 (N_18346,N_17235,N_16900);
and U18347 (N_18347,N_17179,N_16942);
nor U18348 (N_18348,N_17537,N_17084);
or U18349 (N_18349,N_17447,N_16951);
nand U18350 (N_18350,N_16948,N_16998);
and U18351 (N_18351,N_17332,N_16807);
xnor U18352 (N_18352,N_17267,N_17054);
or U18353 (N_18353,N_16828,N_16884);
xnor U18354 (N_18354,N_17588,N_17144);
and U18355 (N_18355,N_16845,N_17065);
nand U18356 (N_18356,N_17359,N_17045);
nor U18357 (N_18357,N_17291,N_17236);
or U18358 (N_18358,N_17187,N_16855);
nand U18359 (N_18359,N_16812,N_16968);
and U18360 (N_18360,N_17043,N_17568);
and U18361 (N_18361,N_17386,N_17027);
nand U18362 (N_18362,N_17242,N_17587);
or U18363 (N_18363,N_17269,N_16827);
or U18364 (N_18364,N_16854,N_17550);
xnor U18365 (N_18365,N_16946,N_17325);
and U18366 (N_18366,N_17028,N_16944);
xnor U18367 (N_18367,N_17257,N_17340);
nor U18368 (N_18368,N_17115,N_16905);
and U18369 (N_18369,N_16847,N_17471);
or U18370 (N_18370,N_17495,N_17215);
nor U18371 (N_18371,N_17313,N_17325);
nand U18372 (N_18372,N_17059,N_17184);
or U18373 (N_18373,N_17035,N_17300);
xor U18374 (N_18374,N_16875,N_16855);
nor U18375 (N_18375,N_17057,N_17005);
and U18376 (N_18376,N_17282,N_17071);
xor U18377 (N_18377,N_17015,N_17016);
xor U18378 (N_18378,N_16914,N_17449);
or U18379 (N_18379,N_17431,N_17203);
xor U18380 (N_18380,N_17476,N_16879);
nand U18381 (N_18381,N_17048,N_16815);
or U18382 (N_18382,N_17202,N_16958);
and U18383 (N_18383,N_16926,N_17365);
nand U18384 (N_18384,N_17536,N_16944);
xnor U18385 (N_18385,N_17220,N_16930);
xor U18386 (N_18386,N_17020,N_17396);
xor U18387 (N_18387,N_17511,N_16854);
nand U18388 (N_18388,N_17329,N_17598);
and U18389 (N_18389,N_17109,N_16963);
nor U18390 (N_18390,N_17092,N_17277);
or U18391 (N_18391,N_17081,N_17492);
or U18392 (N_18392,N_17325,N_17017);
nand U18393 (N_18393,N_17556,N_17429);
and U18394 (N_18394,N_17421,N_17171);
nor U18395 (N_18395,N_16899,N_16826);
and U18396 (N_18396,N_17064,N_17428);
and U18397 (N_18397,N_17283,N_16929);
nand U18398 (N_18398,N_17204,N_16890);
or U18399 (N_18399,N_17189,N_17432);
nor U18400 (N_18400,N_17864,N_18044);
nor U18401 (N_18401,N_18234,N_17721);
and U18402 (N_18402,N_18298,N_18276);
nor U18403 (N_18403,N_18398,N_17895);
nand U18404 (N_18404,N_17905,N_17964);
and U18405 (N_18405,N_17619,N_17917);
nor U18406 (N_18406,N_17691,N_18356);
nand U18407 (N_18407,N_17996,N_18272);
nand U18408 (N_18408,N_18079,N_17612);
xnor U18409 (N_18409,N_18278,N_18053);
nand U18410 (N_18410,N_18026,N_18149);
or U18411 (N_18411,N_18048,N_18258);
nand U18412 (N_18412,N_18254,N_18023);
or U18413 (N_18413,N_18319,N_18144);
xnor U18414 (N_18414,N_17773,N_18037);
and U18415 (N_18415,N_17933,N_18176);
nor U18416 (N_18416,N_18020,N_18185);
nand U18417 (N_18417,N_17757,N_17650);
nor U18418 (N_18418,N_17784,N_17990);
and U18419 (N_18419,N_18046,N_18374);
nor U18420 (N_18420,N_18324,N_18248);
and U18421 (N_18421,N_17720,N_17700);
or U18422 (N_18422,N_17663,N_18004);
xor U18423 (N_18423,N_17787,N_18148);
xor U18424 (N_18424,N_18315,N_18120);
or U18425 (N_18425,N_18098,N_17714);
nand U18426 (N_18426,N_18121,N_18204);
nor U18427 (N_18427,N_18198,N_17742);
xor U18428 (N_18428,N_17897,N_18213);
xnor U18429 (N_18429,N_17927,N_17708);
nand U18430 (N_18430,N_18240,N_18360);
xor U18431 (N_18431,N_17608,N_17791);
xor U18432 (N_18432,N_17898,N_18289);
or U18433 (N_18433,N_18009,N_17849);
and U18434 (N_18434,N_18231,N_18348);
and U18435 (N_18435,N_18122,N_18218);
xnor U18436 (N_18436,N_17821,N_18101);
or U18437 (N_18437,N_17661,N_18192);
and U18438 (N_18438,N_17886,N_18080);
and U18439 (N_18439,N_17688,N_18001);
nand U18440 (N_18440,N_17916,N_18264);
and U18441 (N_18441,N_18334,N_17869);
xor U18442 (N_18442,N_17843,N_17769);
and U18443 (N_18443,N_17948,N_17777);
and U18444 (N_18444,N_17651,N_17707);
nand U18445 (N_18445,N_17960,N_18395);
and U18446 (N_18446,N_18022,N_18104);
and U18447 (N_18447,N_17803,N_17918);
nand U18448 (N_18448,N_18214,N_17727);
or U18449 (N_18449,N_17736,N_17965);
nor U18450 (N_18450,N_17852,N_17765);
xor U18451 (N_18451,N_17672,N_17915);
nand U18452 (N_18452,N_18019,N_18327);
nand U18453 (N_18453,N_17702,N_17668);
nand U18454 (N_18454,N_17794,N_17810);
and U18455 (N_18455,N_18367,N_17719);
and U18456 (N_18456,N_17871,N_18156);
and U18457 (N_18457,N_17985,N_17799);
and U18458 (N_18458,N_17621,N_17838);
and U18459 (N_18459,N_17633,N_18372);
xor U18460 (N_18460,N_17999,N_18394);
nand U18461 (N_18461,N_17988,N_18293);
nand U18462 (N_18462,N_17970,N_18181);
and U18463 (N_18463,N_17882,N_18270);
nand U18464 (N_18464,N_18010,N_17713);
nor U18465 (N_18465,N_17923,N_17796);
nand U18466 (N_18466,N_18034,N_17690);
and U18467 (N_18467,N_17639,N_17634);
or U18468 (N_18468,N_17807,N_18112);
and U18469 (N_18469,N_17903,N_17795);
and U18470 (N_18470,N_18136,N_17913);
or U18471 (N_18471,N_18283,N_17695);
or U18472 (N_18472,N_17630,N_17977);
nand U18473 (N_18473,N_17962,N_17831);
or U18474 (N_18474,N_17804,N_18035);
or U18475 (N_18475,N_17674,N_17638);
or U18476 (N_18476,N_17855,N_18145);
nand U18477 (N_18477,N_17701,N_17772);
nor U18478 (N_18478,N_18342,N_17780);
and U18479 (N_18479,N_18199,N_18141);
nor U18480 (N_18480,N_18369,N_18197);
nor U18481 (N_18481,N_18297,N_17739);
xnor U18482 (N_18482,N_18377,N_17826);
and U18483 (N_18483,N_17767,N_17665);
xor U18484 (N_18484,N_17854,N_18201);
or U18485 (N_18485,N_17866,N_18209);
nor U18486 (N_18486,N_18376,N_18060);
nor U18487 (N_18487,N_18094,N_18280);
xnor U18488 (N_18488,N_18368,N_18143);
xnor U18489 (N_18489,N_18396,N_18229);
nand U18490 (N_18490,N_18294,N_17881);
nor U18491 (N_18491,N_18353,N_18050);
xnor U18492 (N_18492,N_17825,N_17997);
xnor U18493 (N_18493,N_17954,N_17685);
or U18494 (N_18494,N_17762,N_17697);
nand U18495 (N_18495,N_18308,N_18277);
nor U18496 (N_18496,N_18390,N_18203);
nand U18497 (N_18497,N_18347,N_17818);
or U18498 (N_18498,N_18027,N_18383);
nor U18499 (N_18499,N_17649,N_18116);
or U18500 (N_18500,N_18132,N_18117);
and U18501 (N_18501,N_17643,N_18256);
nor U18502 (N_18502,N_17752,N_17790);
and U18503 (N_18503,N_17993,N_17816);
xnor U18504 (N_18504,N_17693,N_18051);
xor U18505 (N_18505,N_17932,N_17968);
or U18506 (N_18506,N_17912,N_18239);
nand U18507 (N_18507,N_17950,N_18165);
and U18508 (N_18508,N_18296,N_17830);
nor U18509 (N_18509,N_18205,N_17856);
nand U18510 (N_18510,N_18320,N_17722);
nand U18511 (N_18511,N_17694,N_18263);
xor U18512 (N_18512,N_18028,N_18069);
and U18513 (N_18513,N_17822,N_18261);
or U18514 (N_18514,N_18118,N_17944);
and U18515 (N_18515,N_18386,N_18110);
and U18516 (N_18516,N_17745,N_17610);
nor U18517 (N_18517,N_18077,N_18056);
nand U18518 (N_18518,N_17675,N_18091);
or U18519 (N_18519,N_17711,N_18179);
xnor U18520 (N_18520,N_18066,N_18173);
or U18521 (N_18521,N_17874,N_18333);
nor U18522 (N_18522,N_17737,N_18139);
xnor U18523 (N_18523,N_17924,N_18178);
and U18524 (N_18524,N_18221,N_17802);
and U18525 (N_18525,N_17601,N_17836);
nor U18526 (N_18526,N_17979,N_17963);
nor U18527 (N_18527,N_18232,N_17622);
nor U18528 (N_18528,N_18155,N_18375);
xor U18529 (N_18529,N_18206,N_17880);
nor U18530 (N_18530,N_17914,N_17906);
xor U18531 (N_18531,N_17641,N_18302);
nor U18532 (N_18532,N_17760,N_17605);
nor U18533 (N_18533,N_18182,N_17656);
nor U18534 (N_18534,N_17770,N_17861);
xor U18535 (N_18535,N_17961,N_17792);
nor U18536 (N_18536,N_17788,N_18236);
nor U18537 (N_18537,N_17669,N_17890);
nor U18538 (N_18538,N_17683,N_17659);
nand U18539 (N_18539,N_18049,N_17910);
xnor U18540 (N_18540,N_17805,N_18247);
and U18541 (N_18541,N_18194,N_18012);
nand U18542 (N_18542,N_18140,N_17718);
or U18543 (N_18543,N_17764,N_18275);
or U18544 (N_18544,N_18024,N_18337);
and U18545 (N_18545,N_17726,N_18159);
nor U18546 (N_18546,N_18115,N_17870);
or U18547 (N_18547,N_18260,N_18305);
or U18548 (N_18548,N_17715,N_17603);
or U18549 (N_18549,N_18371,N_18146);
nor U18550 (N_18550,N_18288,N_17824);
and U18551 (N_18551,N_18067,N_17834);
nand U18552 (N_18552,N_17637,N_18029);
and U18553 (N_18553,N_17751,N_18335);
nand U18554 (N_18554,N_17823,N_18059);
xor U18555 (N_18555,N_17863,N_18061);
nor U18556 (N_18556,N_17686,N_18107);
nor U18557 (N_18557,N_17640,N_17820);
or U18558 (N_18558,N_17952,N_17666);
or U18559 (N_18559,N_18161,N_17862);
nand U18560 (N_18560,N_18190,N_17936);
or U18561 (N_18561,N_17889,N_18138);
xnor U18562 (N_18562,N_17837,N_17934);
nand U18563 (N_18563,N_18030,N_18290);
nor U18564 (N_18564,N_17884,N_17632);
nor U18565 (N_18565,N_18378,N_17725);
nor U18566 (N_18566,N_18226,N_17776);
or U18567 (N_18567,N_17723,N_17983);
nor U18568 (N_18568,N_18108,N_18040);
nor U18569 (N_18569,N_18154,N_17626);
and U18570 (N_18570,N_18129,N_17867);
nand U18571 (N_18571,N_18325,N_18249);
or U18572 (N_18572,N_17828,N_18245);
or U18573 (N_18573,N_17853,N_17696);
or U18574 (N_18574,N_17717,N_18151);
nand U18575 (N_18575,N_18097,N_17989);
xnor U18576 (N_18576,N_18338,N_17966);
or U18577 (N_18577,N_18153,N_17972);
or U18578 (N_18578,N_17710,N_18281);
xnor U18579 (N_18579,N_18031,N_18211);
or U18580 (N_18580,N_17938,N_17677);
and U18581 (N_18581,N_17931,N_18177);
xnor U18582 (N_18582,N_17763,N_17833);
nor U18583 (N_18583,N_17967,N_17782);
nand U18584 (N_18584,N_18253,N_17607);
nand U18585 (N_18585,N_17613,N_17892);
or U18586 (N_18586,N_17857,N_17749);
xor U18587 (N_18587,N_18262,N_18220);
or U18588 (N_18588,N_18219,N_17879);
and U18589 (N_18589,N_17644,N_18358);
nor U18590 (N_18590,N_17609,N_18180);
or U18591 (N_18591,N_18343,N_18168);
nand U18592 (N_18592,N_18064,N_17980);
or U18593 (N_18593,N_17744,N_18167);
nor U18594 (N_18594,N_18244,N_17768);
and U18595 (N_18595,N_18332,N_17635);
nor U18596 (N_18596,N_17998,N_17671);
xnor U18597 (N_18597,N_18126,N_17922);
nor U18598 (N_18598,N_18299,N_18225);
nand U18599 (N_18599,N_17908,N_18307);
or U18600 (N_18600,N_18076,N_17646);
nand U18601 (N_18601,N_18391,N_17684);
and U18602 (N_18602,N_17682,N_18216);
nand U18603 (N_18603,N_17887,N_18123);
xnor U18604 (N_18604,N_18323,N_17786);
xnor U18605 (N_18605,N_18235,N_17800);
nor U18606 (N_18606,N_17740,N_18025);
xnor U18607 (N_18607,N_18152,N_18088);
xor U18608 (N_18608,N_18354,N_18033);
xor U18609 (N_18609,N_18243,N_17900);
or U18610 (N_18610,N_17883,N_18363);
xor U18611 (N_18611,N_17653,N_18212);
nand U18612 (N_18612,N_17629,N_18352);
and U18613 (N_18613,N_18252,N_18114);
xnor U18614 (N_18614,N_18350,N_18142);
and U18615 (N_18615,N_18196,N_18399);
xnor U18616 (N_18616,N_17835,N_18286);
xor U18617 (N_18617,N_17919,N_18063);
and U18618 (N_18618,N_17705,N_18224);
or U18619 (N_18619,N_18238,N_18357);
nor U18620 (N_18620,N_18015,N_17746);
or U18621 (N_18621,N_17812,N_18021);
and U18622 (N_18622,N_17687,N_17808);
xnor U18623 (N_18623,N_18379,N_17928);
or U18624 (N_18624,N_18300,N_18246);
nor U18625 (N_18625,N_18113,N_17730);
or U18626 (N_18626,N_17814,N_18385);
and U18627 (N_18627,N_18392,N_18295);
or U18628 (N_18628,N_18380,N_18047);
nor U18629 (N_18629,N_17941,N_17991);
xnor U18630 (N_18630,N_18070,N_18166);
nor U18631 (N_18631,N_17827,N_18092);
nor U18632 (N_18632,N_17628,N_17907);
nand U18633 (N_18633,N_18073,N_17606);
or U18634 (N_18634,N_18018,N_18291);
or U18635 (N_18635,N_17655,N_17951);
nor U18636 (N_18636,N_18075,N_17945);
nand U18637 (N_18637,N_17847,N_18174);
xnor U18638 (N_18638,N_18084,N_17832);
or U18639 (N_18639,N_17728,N_18128);
nor U18640 (N_18640,N_18125,N_17899);
xnor U18641 (N_18641,N_18169,N_17955);
and U18642 (N_18642,N_17636,N_18388);
and U18643 (N_18643,N_17648,N_18311);
xnor U18644 (N_18644,N_18314,N_17733);
xor U18645 (N_18645,N_18267,N_17995);
xor U18646 (N_18646,N_17809,N_17738);
or U18647 (N_18647,N_18002,N_17771);
and U18648 (N_18648,N_17747,N_18111);
nor U18649 (N_18649,N_17706,N_17766);
nor U18650 (N_18650,N_17842,N_17971);
or U18651 (N_18651,N_17986,N_18147);
nand U18652 (N_18652,N_17750,N_17698);
and U18653 (N_18653,N_18036,N_18131);
nand U18654 (N_18654,N_18109,N_17623);
nand U18655 (N_18655,N_17819,N_18191);
or U18656 (N_18656,N_17981,N_18105);
xnor U18657 (N_18657,N_18043,N_18103);
xor U18658 (N_18658,N_17678,N_17743);
nor U18659 (N_18659,N_17627,N_18086);
nor U18660 (N_18660,N_18382,N_17896);
xor U18661 (N_18661,N_17956,N_18310);
xnor U18662 (N_18662,N_18208,N_17615);
xor U18663 (N_18663,N_18013,N_17958);
nor U18664 (N_18664,N_17909,N_18393);
or U18665 (N_18665,N_17920,N_18119);
xnor U18666 (N_18666,N_18257,N_18366);
and U18667 (N_18667,N_18329,N_17673);
xnor U18668 (N_18668,N_17959,N_17875);
or U18669 (N_18669,N_17729,N_18309);
or U18670 (N_18670,N_17850,N_17873);
xnor U18671 (N_18671,N_17600,N_18389);
nor U18672 (N_18672,N_18135,N_17930);
or U18673 (N_18673,N_18215,N_17617);
and U18674 (N_18674,N_18273,N_18162);
or U18675 (N_18675,N_18274,N_17785);
nor U18676 (N_18676,N_18362,N_17779);
xor U18677 (N_18677,N_18222,N_18137);
and U18678 (N_18678,N_17789,N_17647);
or U18679 (N_18679,N_17878,N_17676);
nand U18680 (N_18680,N_17953,N_17658);
and U18681 (N_18681,N_17741,N_18359);
nand U18682 (N_18682,N_18387,N_17929);
or U18683 (N_18683,N_17811,N_17815);
nand U18684 (N_18684,N_17652,N_18345);
and U18685 (N_18685,N_17716,N_17664);
or U18686 (N_18686,N_17885,N_18330);
and U18687 (N_18687,N_18200,N_18187);
or U18688 (N_18688,N_18188,N_17943);
and U18689 (N_18689,N_18316,N_18202);
or U18690 (N_18690,N_17775,N_18365);
or U18691 (N_18691,N_18102,N_18301);
xnor U18692 (N_18692,N_18172,N_17798);
nor U18693 (N_18693,N_18336,N_17982);
or U18694 (N_18694,N_18279,N_17625);
xor U18695 (N_18695,N_18065,N_17654);
or U18696 (N_18696,N_18082,N_18326);
xor U18697 (N_18697,N_18157,N_18317);
nor U18698 (N_18698,N_17860,N_17872);
xnor U18699 (N_18699,N_17865,N_17797);
nand U18700 (N_18700,N_17957,N_18087);
and U18701 (N_18701,N_17748,N_18361);
or U18702 (N_18702,N_17921,N_17731);
and U18703 (N_18703,N_18133,N_18341);
and U18704 (N_18704,N_18313,N_17926);
nor U18705 (N_18705,N_17829,N_17774);
xnor U18706 (N_18706,N_17734,N_18014);
or U18707 (N_18707,N_17781,N_18071);
xor U18708 (N_18708,N_18042,N_18106);
and U18709 (N_18709,N_18318,N_17709);
xnor U18710 (N_18710,N_18008,N_18349);
nor U18711 (N_18711,N_17868,N_18269);
or U18712 (N_18712,N_17806,N_17624);
xor U18713 (N_18713,N_17946,N_17891);
nor U18714 (N_18714,N_17620,N_17969);
and U18715 (N_18715,N_18062,N_18304);
xor U18716 (N_18716,N_18292,N_17901);
and U18717 (N_18717,N_18081,N_17949);
nor U18718 (N_18718,N_18045,N_17732);
nor U18719 (N_18719,N_18007,N_18321);
nor U18720 (N_18720,N_17976,N_17618);
or U18721 (N_18721,N_18237,N_17937);
or U18722 (N_18722,N_17611,N_17848);
nor U18723 (N_18723,N_18207,N_18100);
nor U18724 (N_18724,N_17801,N_17679);
or U18725 (N_18725,N_18055,N_18052);
or U18726 (N_18726,N_17973,N_18384);
nand U18727 (N_18727,N_18250,N_17778);
nand U18728 (N_18728,N_18090,N_17680);
nand U18729 (N_18729,N_17783,N_18268);
xor U18730 (N_18730,N_17851,N_17940);
xor U18731 (N_18731,N_18000,N_17793);
and U18732 (N_18732,N_17935,N_18150);
xnor U18733 (N_18733,N_18340,N_18282);
and U18734 (N_18734,N_18210,N_18266);
and U18735 (N_18735,N_18355,N_17692);
xnor U18736 (N_18736,N_17662,N_17689);
xnor U18737 (N_18737,N_17844,N_17876);
nand U18738 (N_18738,N_17753,N_18072);
nand U18739 (N_18739,N_18085,N_18160);
xor U18740 (N_18740,N_18285,N_17939);
nor U18741 (N_18741,N_17987,N_18093);
xnor U18742 (N_18742,N_18171,N_18364);
nand U18743 (N_18743,N_18095,N_18223);
and U18744 (N_18744,N_17994,N_17902);
nor U18745 (N_18745,N_18054,N_18303);
or U18746 (N_18746,N_18328,N_18175);
or U18747 (N_18747,N_18074,N_18344);
xor U18748 (N_18748,N_17754,N_18339);
xnor U18749 (N_18749,N_18078,N_18312);
or U18750 (N_18750,N_18242,N_18038);
or U18751 (N_18751,N_17681,N_18005);
or U18752 (N_18752,N_17660,N_18370);
xnor U18753 (N_18753,N_17893,N_17759);
or U18754 (N_18754,N_18351,N_17703);
nand U18755 (N_18755,N_18183,N_17817);
nor U18756 (N_18756,N_18124,N_18306);
xor U18757 (N_18757,N_18259,N_17631);
nand U18758 (N_18758,N_17925,N_17667);
nand U18759 (N_18759,N_17616,N_18158);
nand U18760 (N_18760,N_18096,N_18241);
and U18761 (N_18761,N_18041,N_17845);
xor U18762 (N_18762,N_17704,N_18271);
xor U18763 (N_18763,N_18184,N_18265);
or U18764 (N_18764,N_18381,N_18057);
or U18765 (N_18765,N_17841,N_17992);
nor U18766 (N_18766,N_18251,N_17813);
or U18767 (N_18767,N_18287,N_17877);
and U18768 (N_18768,N_18230,N_18130);
and U18769 (N_18769,N_18193,N_17755);
and U18770 (N_18770,N_17984,N_18032);
xnor U18771 (N_18771,N_18127,N_18331);
and U18772 (N_18772,N_17859,N_18164);
or U18773 (N_18773,N_18170,N_18039);
and U18774 (N_18774,N_18006,N_17974);
nand U18775 (N_18775,N_17642,N_17839);
nor U18776 (N_18776,N_17894,N_17657);
and U18777 (N_18777,N_18284,N_17724);
xnor U18778 (N_18778,N_18099,N_18083);
nor U18779 (N_18779,N_18003,N_18089);
nor U18780 (N_18780,N_18189,N_17645);
and U18781 (N_18781,N_18163,N_17858);
nand U18782 (N_18782,N_18228,N_18195);
nand U18783 (N_18783,N_18016,N_17602);
nor U18784 (N_18784,N_17735,N_18186);
xor U18785 (N_18785,N_17942,N_17888);
nor U18786 (N_18786,N_18227,N_17670);
nor U18787 (N_18787,N_18134,N_18017);
and U18788 (N_18788,N_17846,N_17978);
nor U18789 (N_18789,N_18373,N_17947);
nand U18790 (N_18790,N_17604,N_18058);
nand U18791 (N_18791,N_18255,N_17975);
or U18792 (N_18792,N_18322,N_18233);
xor U18793 (N_18793,N_18346,N_17712);
nor U18794 (N_18794,N_18217,N_17614);
and U18795 (N_18795,N_18397,N_17904);
xor U18796 (N_18796,N_17756,N_17840);
and U18797 (N_18797,N_17761,N_18068);
and U18798 (N_18798,N_17911,N_17699);
nand U18799 (N_18799,N_18011,N_17758);
and U18800 (N_18800,N_17830,N_18312);
xnor U18801 (N_18801,N_18128,N_17942);
or U18802 (N_18802,N_18268,N_17803);
xnor U18803 (N_18803,N_18347,N_17676);
xnor U18804 (N_18804,N_17737,N_17645);
nor U18805 (N_18805,N_17630,N_18068);
nand U18806 (N_18806,N_18370,N_18098);
xnor U18807 (N_18807,N_17984,N_17857);
xnor U18808 (N_18808,N_18250,N_18170);
nand U18809 (N_18809,N_18311,N_17884);
nand U18810 (N_18810,N_17804,N_17736);
nand U18811 (N_18811,N_17928,N_18021);
xor U18812 (N_18812,N_18152,N_18384);
or U18813 (N_18813,N_17867,N_17820);
nor U18814 (N_18814,N_17801,N_18298);
or U18815 (N_18815,N_17796,N_17843);
and U18816 (N_18816,N_17882,N_18147);
and U18817 (N_18817,N_17704,N_18287);
and U18818 (N_18818,N_17753,N_18175);
nand U18819 (N_18819,N_18067,N_17937);
nor U18820 (N_18820,N_17718,N_18395);
and U18821 (N_18821,N_17615,N_18235);
and U18822 (N_18822,N_17800,N_18293);
nand U18823 (N_18823,N_18218,N_18191);
and U18824 (N_18824,N_17779,N_18012);
xor U18825 (N_18825,N_17674,N_17636);
or U18826 (N_18826,N_17870,N_18358);
xnor U18827 (N_18827,N_17881,N_18071);
nand U18828 (N_18828,N_17656,N_17623);
nand U18829 (N_18829,N_17792,N_18207);
nand U18830 (N_18830,N_18396,N_18133);
nor U18831 (N_18831,N_17920,N_18388);
xnor U18832 (N_18832,N_17746,N_17651);
nand U18833 (N_18833,N_18172,N_18315);
xnor U18834 (N_18834,N_17784,N_17795);
xnor U18835 (N_18835,N_18335,N_17928);
nand U18836 (N_18836,N_17819,N_17692);
nand U18837 (N_18837,N_18325,N_18293);
nand U18838 (N_18838,N_18262,N_18291);
xnor U18839 (N_18839,N_17684,N_17755);
and U18840 (N_18840,N_18386,N_18322);
nor U18841 (N_18841,N_18353,N_17775);
nor U18842 (N_18842,N_18268,N_17841);
xnor U18843 (N_18843,N_18277,N_18357);
nor U18844 (N_18844,N_18276,N_18087);
and U18845 (N_18845,N_18231,N_17930);
xnor U18846 (N_18846,N_18318,N_18215);
xor U18847 (N_18847,N_18365,N_17987);
or U18848 (N_18848,N_17974,N_18090);
nor U18849 (N_18849,N_18025,N_17828);
nand U18850 (N_18850,N_17696,N_18260);
or U18851 (N_18851,N_17947,N_17995);
nor U18852 (N_18852,N_17711,N_17953);
nor U18853 (N_18853,N_18191,N_18023);
nand U18854 (N_18854,N_18326,N_18119);
or U18855 (N_18855,N_18077,N_17794);
and U18856 (N_18856,N_17632,N_18226);
nand U18857 (N_18857,N_18036,N_18057);
nand U18858 (N_18858,N_17838,N_17850);
nor U18859 (N_18859,N_18059,N_18306);
or U18860 (N_18860,N_17606,N_18059);
and U18861 (N_18861,N_17918,N_18216);
nor U18862 (N_18862,N_17787,N_17997);
nor U18863 (N_18863,N_18106,N_17764);
nand U18864 (N_18864,N_17915,N_18357);
nor U18865 (N_18865,N_17964,N_18229);
nand U18866 (N_18866,N_17981,N_17633);
and U18867 (N_18867,N_18142,N_18162);
xor U18868 (N_18868,N_18077,N_18071);
and U18869 (N_18869,N_17672,N_18178);
nor U18870 (N_18870,N_18042,N_18370);
nand U18871 (N_18871,N_18046,N_17644);
nor U18872 (N_18872,N_18058,N_17872);
or U18873 (N_18873,N_17694,N_18205);
and U18874 (N_18874,N_17872,N_18339);
xor U18875 (N_18875,N_18215,N_18392);
nand U18876 (N_18876,N_17731,N_18168);
xor U18877 (N_18877,N_18386,N_18323);
nand U18878 (N_18878,N_17906,N_17605);
or U18879 (N_18879,N_18082,N_18052);
or U18880 (N_18880,N_17620,N_17640);
nor U18881 (N_18881,N_17928,N_18123);
xnor U18882 (N_18882,N_17883,N_17669);
and U18883 (N_18883,N_18258,N_18282);
and U18884 (N_18884,N_17851,N_17991);
nor U18885 (N_18885,N_18077,N_18194);
and U18886 (N_18886,N_17929,N_17761);
xor U18887 (N_18887,N_18276,N_18139);
and U18888 (N_18888,N_17806,N_18013);
or U18889 (N_18889,N_18278,N_17994);
and U18890 (N_18890,N_18271,N_17883);
xnor U18891 (N_18891,N_18274,N_18053);
xor U18892 (N_18892,N_17632,N_17842);
nand U18893 (N_18893,N_17966,N_18315);
nand U18894 (N_18894,N_17729,N_18251);
and U18895 (N_18895,N_17884,N_18377);
nand U18896 (N_18896,N_17939,N_18045);
and U18897 (N_18897,N_17691,N_17876);
xor U18898 (N_18898,N_17723,N_17986);
or U18899 (N_18899,N_17741,N_18381);
and U18900 (N_18900,N_18040,N_18038);
or U18901 (N_18901,N_17971,N_17826);
nor U18902 (N_18902,N_17828,N_17793);
and U18903 (N_18903,N_18260,N_18265);
or U18904 (N_18904,N_18093,N_17949);
xnor U18905 (N_18905,N_18084,N_18130);
nand U18906 (N_18906,N_17955,N_18080);
nor U18907 (N_18907,N_18155,N_18376);
nor U18908 (N_18908,N_17763,N_18183);
nor U18909 (N_18909,N_18011,N_18386);
xnor U18910 (N_18910,N_18299,N_17671);
nand U18911 (N_18911,N_18131,N_18339);
nor U18912 (N_18912,N_17800,N_17941);
and U18913 (N_18913,N_17689,N_18222);
and U18914 (N_18914,N_17884,N_18313);
or U18915 (N_18915,N_17799,N_17631);
xor U18916 (N_18916,N_17990,N_18314);
and U18917 (N_18917,N_17862,N_17660);
or U18918 (N_18918,N_17888,N_17980);
nor U18919 (N_18919,N_17955,N_18001);
xor U18920 (N_18920,N_18399,N_17843);
or U18921 (N_18921,N_18240,N_18302);
and U18922 (N_18922,N_18272,N_18166);
xor U18923 (N_18923,N_17674,N_17725);
nor U18924 (N_18924,N_18133,N_18382);
nand U18925 (N_18925,N_18380,N_17895);
and U18926 (N_18926,N_17945,N_18042);
and U18927 (N_18927,N_17727,N_17654);
and U18928 (N_18928,N_18302,N_18176);
and U18929 (N_18929,N_18136,N_17801);
xor U18930 (N_18930,N_18076,N_18173);
xor U18931 (N_18931,N_18392,N_17683);
nor U18932 (N_18932,N_17994,N_17820);
and U18933 (N_18933,N_17674,N_17955);
nor U18934 (N_18934,N_17838,N_18201);
or U18935 (N_18935,N_17722,N_18358);
nor U18936 (N_18936,N_17705,N_18348);
and U18937 (N_18937,N_18166,N_17677);
nand U18938 (N_18938,N_18058,N_17790);
or U18939 (N_18939,N_17865,N_17756);
and U18940 (N_18940,N_17983,N_18186);
xor U18941 (N_18941,N_17934,N_17786);
nand U18942 (N_18942,N_17985,N_18161);
and U18943 (N_18943,N_18127,N_17896);
xor U18944 (N_18944,N_18105,N_17902);
nor U18945 (N_18945,N_18265,N_18001);
or U18946 (N_18946,N_17638,N_18031);
nand U18947 (N_18947,N_18303,N_17842);
xor U18948 (N_18948,N_17888,N_18015);
xor U18949 (N_18949,N_17940,N_18178);
nor U18950 (N_18950,N_17760,N_17951);
or U18951 (N_18951,N_17892,N_18256);
xnor U18952 (N_18952,N_18131,N_18362);
and U18953 (N_18953,N_18206,N_17693);
or U18954 (N_18954,N_18382,N_18383);
and U18955 (N_18955,N_18274,N_18145);
or U18956 (N_18956,N_17834,N_18385);
nor U18957 (N_18957,N_18002,N_18094);
and U18958 (N_18958,N_17864,N_17601);
nor U18959 (N_18959,N_18186,N_17972);
or U18960 (N_18960,N_17851,N_18242);
nand U18961 (N_18961,N_18204,N_18356);
and U18962 (N_18962,N_18030,N_17609);
nor U18963 (N_18963,N_18278,N_17607);
or U18964 (N_18964,N_17670,N_18136);
nor U18965 (N_18965,N_17783,N_17856);
nand U18966 (N_18966,N_18273,N_17787);
or U18967 (N_18967,N_17913,N_18188);
nand U18968 (N_18968,N_18376,N_18255);
nand U18969 (N_18969,N_17853,N_17941);
nor U18970 (N_18970,N_17692,N_18094);
or U18971 (N_18971,N_17773,N_18164);
nand U18972 (N_18972,N_17853,N_17970);
nor U18973 (N_18973,N_17800,N_17965);
nand U18974 (N_18974,N_17845,N_17858);
and U18975 (N_18975,N_17780,N_17791);
and U18976 (N_18976,N_18122,N_18380);
xor U18977 (N_18977,N_17879,N_18138);
or U18978 (N_18978,N_17604,N_18068);
nand U18979 (N_18979,N_18121,N_18279);
or U18980 (N_18980,N_17645,N_18263);
xor U18981 (N_18981,N_18202,N_17721);
nor U18982 (N_18982,N_17948,N_18191);
nand U18983 (N_18983,N_18150,N_18278);
xor U18984 (N_18984,N_17738,N_18286);
nor U18985 (N_18985,N_17624,N_18299);
nand U18986 (N_18986,N_17808,N_18228);
or U18987 (N_18987,N_18338,N_17834);
and U18988 (N_18988,N_18350,N_17702);
or U18989 (N_18989,N_17939,N_18293);
nand U18990 (N_18990,N_17769,N_17947);
and U18991 (N_18991,N_18151,N_17781);
nor U18992 (N_18992,N_17922,N_17633);
xnor U18993 (N_18993,N_17712,N_17786);
nand U18994 (N_18994,N_18033,N_17701);
and U18995 (N_18995,N_17784,N_17628);
nor U18996 (N_18996,N_17815,N_17778);
and U18997 (N_18997,N_18138,N_17929);
nor U18998 (N_18998,N_17886,N_18143);
or U18999 (N_18999,N_18163,N_17794);
nand U19000 (N_19000,N_18087,N_18266);
nand U19001 (N_19001,N_17862,N_18033);
nand U19002 (N_19002,N_18086,N_17678);
or U19003 (N_19003,N_17919,N_17845);
nor U19004 (N_19004,N_18108,N_18170);
or U19005 (N_19005,N_17643,N_18232);
nand U19006 (N_19006,N_18170,N_17656);
nand U19007 (N_19007,N_17858,N_17721);
xor U19008 (N_19008,N_18035,N_18224);
nand U19009 (N_19009,N_17673,N_18105);
nor U19010 (N_19010,N_17641,N_18272);
and U19011 (N_19011,N_17842,N_17624);
xor U19012 (N_19012,N_17931,N_18237);
nand U19013 (N_19013,N_17743,N_18346);
nor U19014 (N_19014,N_17950,N_17999);
or U19015 (N_19015,N_18391,N_18062);
and U19016 (N_19016,N_18261,N_17665);
and U19017 (N_19017,N_17661,N_17616);
or U19018 (N_19018,N_18271,N_17828);
and U19019 (N_19019,N_18010,N_17866);
and U19020 (N_19020,N_18112,N_17863);
nor U19021 (N_19021,N_17807,N_18012);
and U19022 (N_19022,N_18285,N_17721);
nor U19023 (N_19023,N_18387,N_18358);
and U19024 (N_19024,N_18073,N_18319);
or U19025 (N_19025,N_17742,N_18030);
nand U19026 (N_19026,N_18294,N_17622);
nand U19027 (N_19027,N_18064,N_17707);
nand U19028 (N_19028,N_17823,N_18073);
xor U19029 (N_19029,N_17991,N_17875);
nand U19030 (N_19030,N_18024,N_18369);
xor U19031 (N_19031,N_18352,N_17880);
or U19032 (N_19032,N_18269,N_17605);
nand U19033 (N_19033,N_18004,N_17601);
xor U19034 (N_19034,N_18095,N_18331);
nor U19035 (N_19035,N_17971,N_17878);
and U19036 (N_19036,N_18175,N_17760);
nand U19037 (N_19037,N_18021,N_18206);
nand U19038 (N_19038,N_18096,N_18108);
xor U19039 (N_19039,N_17943,N_17955);
xnor U19040 (N_19040,N_17972,N_18102);
and U19041 (N_19041,N_18326,N_17611);
and U19042 (N_19042,N_18135,N_17967);
or U19043 (N_19043,N_18095,N_18382);
nor U19044 (N_19044,N_17998,N_18351);
nand U19045 (N_19045,N_17618,N_17950);
nand U19046 (N_19046,N_18359,N_17925);
nor U19047 (N_19047,N_17962,N_17721);
xor U19048 (N_19048,N_17638,N_17851);
xor U19049 (N_19049,N_17832,N_17610);
nand U19050 (N_19050,N_18399,N_18126);
or U19051 (N_19051,N_17633,N_18209);
xnor U19052 (N_19052,N_18371,N_17806);
nor U19053 (N_19053,N_17619,N_17959);
nand U19054 (N_19054,N_17777,N_17713);
or U19055 (N_19055,N_17953,N_17921);
or U19056 (N_19056,N_17845,N_18120);
and U19057 (N_19057,N_18217,N_17942);
and U19058 (N_19058,N_18395,N_18387);
nand U19059 (N_19059,N_17915,N_18072);
nor U19060 (N_19060,N_17745,N_17834);
or U19061 (N_19061,N_17619,N_17766);
nand U19062 (N_19062,N_17784,N_18308);
or U19063 (N_19063,N_17637,N_18040);
xnor U19064 (N_19064,N_18171,N_18118);
or U19065 (N_19065,N_18324,N_18047);
or U19066 (N_19066,N_17875,N_18330);
or U19067 (N_19067,N_17879,N_18013);
or U19068 (N_19068,N_18102,N_17827);
and U19069 (N_19069,N_17658,N_17781);
nand U19070 (N_19070,N_18144,N_18067);
nor U19071 (N_19071,N_17865,N_17723);
or U19072 (N_19072,N_17886,N_17925);
nand U19073 (N_19073,N_17704,N_17616);
or U19074 (N_19074,N_17797,N_18387);
or U19075 (N_19075,N_18068,N_17895);
nor U19076 (N_19076,N_17878,N_18141);
and U19077 (N_19077,N_17624,N_17923);
nor U19078 (N_19078,N_18064,N_18043);
or U19079 (N_19079,N_18344,N_18121);
xnor U19080 (N_19080,N_17698,N_17860);
nand U19081 (N_19081,N_18128,N_17784);
or U19082 (N_19082,N_17973,N_17662);
and U19083 (N_19083,N_18181,N_17987);
xnor U19084 (N_19084,N_17959,N_17602);
nand U19085 (N_19085,N_18302,N_17919);
xor U19086 (N_19086,N_18257,N_17807);
xor U19087 (N_19087,N_18374,N_18078);
and U19088 (N_19088,N_17738,N_18183);
nor U19089 (N_19089,N_18303,N_17955);
xnor U19090 (N_19090,N_17649,N_18397);
nand U19091 (N_19091,N_18218,N_18223);
nand U19092 (N_19092,N_18085,N_17960);
and U19093 (N_19093,N_17737,N_17876);
nand U19094 (N_19094,N_17697,N_18072);
nand U19095 (N_19095,N_18115,N_17638);
or U19096 (N_19096,N_17619,N_17845);
and U19097 (N_19097,N_17783,N_18053);
nand U19098 (N_19098,N_17934,N_17877);
or U19099 (N_19099,N_17748,N_18395);
nor U19100 (N_19100,N_18167,N_18035);
xnor U19101 (N_19101,N_17937,N_18226);
nor U19102 (N_19102,N_17815,N_17608);
xnor U19103 (N_19103,N_18168,N_18374);
xor U19104 (N_19104,N_18040,N_17866);
or U19105 (N_19105,N_18239,N_18307);
xnor U19106 (N_19106,N_18090,N_18145);
and U19107 (N_19107,N_17955,N_17786);
nor U19108 (N_19108,N_17923,N_18165);
or U19109 (N_19109,N_18242,N_18334);
nor U19110 (N_19110,N_18069,N_17902);
nand U19111 (N_19111,N_17677,N_18116);
nor U19112 (N_19112,N_18258,N_17764);
and U19113 (N_19113,N_18350,N_17844);
nor U19114 (N_19114,N_17613,N_18221);
or U19115 (N_19115,N_18204,N_17940);
xnor U19116 (N_19116,N_17967,N_17653);
and U19117 (N_19117,N_18164,N_18001);
nand U19118 (N_19118,N_17696,N_18175);
and U19119 (N_19119,N_18266,N_18369);
xnor U19120 (N_19120,N_18394,N_18213);
xnor U19121 (N_19121,N_18242,N_18165);
and U19122 (N_19122,N_18080,N_18113);
and U19123 (N_19123,N_18059,N_17773);
and U19124 (N_19124,N_18106,N_18184);
or U19125 (N_19125,N_17970,N_18186);
or U19126 (N_19126,N_17811,N_18139);
or U19127 (N_19127,N_17821,N_18294);
nand U19128 (N_19128,N_18194,N_18299);
xnor U19129 (N_19129,N_18177,N_17904);
nor U19130 (N_19130,N_18130,N_18273);
nor U19131 (N_19131,N_18312,N_17697);
or U19132 (N_19132,N_17615,N_17979);
xor U19133 (N_19133,N_17802,N_18140);
or U19134 (N_19134,N_18346,N_17637);
and U19135 (N_19135,N_17678,N_18399);
nand U19136 (N_19136,N_17946,N_17667);
or U19137 (N_19137,N_18055,N_17681);
nand U19138 (N_19138,N_17904,N_18135);
nor U19139 (N_19139,N_17780,N_18350);
xor U19140 (N_19140,N_17630,N_17965);
nor U19141 (N_19141,N_17741,N_17750);
or U19142 (N_19142,N_17964,N_17704);
or U19143 (N_19143,N_17955,N_18000);
or U19144 (N_19144,N_18245,N_18033);
nand U19145 (N_19145,N_17808,N_18164);
nand U19146 (N_19146,N_18298,N_18181);
nand U19147 (N_19147,N_17923,N_18049);
or U19148 (N_19148,N_17768,N_17802);
xnor U19149 (N_19149,N_18108,N_18292);
and U19150 (N_19150,N_18093,N_17649);
and U19151 (N_19151,N_17809,N_17821);
or U19152 (N_19152,N_18349,N_17903);
nand U19153 (N_19153,N_17668,N_18162);
nor U19154 (N_19154,N_18047,N_18181);
xor U19155 (N_19155,N_17688,N_18358);
xor U19156 (N_19156,N_18342,N_17719);
nor U19157 (N_19157,N_17902,N_18379);
or U19158 (N_19158,N_18015,N_17864);
or U19159 (N_19159,N_18005,N_18129);
nor U19160 (N_19160,N_17906,N_18340);
xnor U19161 (N_19161,N_18197,N_17879);
xor U19162 (N_19162,N_18013,N_18262);
nor U19163 (N_19163,N_18379,N_17804);
nor U19164 (N_19164,N_18128,N_18348);
nor U19165 (N_19165,N_18231,N_17987);
nor U19166 (N_19166,N_17840,N_17656);
nand U19167 (N_19167,N_17813,N_17714);
xor U19168 (N_19168,N_17954,N_18221);
nand U19169 (N_19169,N_18112,N_17720);
and U19170 (N_19170,N_17938,N_17914);
or U19171 (N_19171,N_18234,N_17996);
or U19172 (N_19172,N_18376,N_18303);
or U19173 (N_19173,N_17901,N_17851);
and U19174 (N_19174,N_18006,N_17889);
and U19175 (N_19175,N_17853,N_17625);
nor U19176 (N_19176,N_18171,N_17798);
or U19177 (N_19177,N_17612,N_17788);
nand U19178 (N_19178,N_18144,N_17851);
nand U19179 (N_19179,N_17689,N_17813);
and U19180 (N_19180,N_18333,N_18315);
or U19181 (N_19181,N_17759,N_18094);
and U19182 (N_19182,N_17821,N_17627);
nand U19183 (N_19183,N_17989,N_18223);
nor U19184 (N_19184,N_17897,N_17679);
nand U19185 (N_19185,N_17992,N_18243);
xnor U19186 (N_19186,N_17739,N_18296);
nor U19187 (N_19187,N_17913,N_17726);
or U19188 (N_19188,N_17747,N_18314);
nor U19189 (N_19189,N_17689,N_17922);
and U19190 (N_19190,N_17809,N_17611);
or U19191 (N_19191,N_17921,N_18365);
xnor U19192 (N_19192,N_18059,N_17746);
xor U19193 (N_19193,N_17755,N_17692);
or U19194 (N_19194,N_17819,N_17704);
and U19195 (N_19195,N_18277,N_17711);
nor U19196 (N_19196,N_18318,N_18221);
nor U19197 (N_19197,N_18013,N_17892);
or U19198 (N_19198,N_18159,N_17928);
nor U19199 (N_19199,N_17746,N_17601);
and U19200 (N_19200,N_19178,N_18702);
or U19201 (N_19201,N_18804,N_18657);
nand U19202 (N_19202,N_18487,N_18472);
nor U19203 (N_19203,N_19199,N_19085);
and U19204 (N_19204,N_18890,N_19133);
and U19205 (N_19205,N_18835,N_18427);
nor U19206 (N_19206,N_18827,N_18496);
and U19207 (N_19207,N_18900,N_18676);
nand U19208 (N_19208,N_18565,N_18765);
and U19209 (N_19209,N_19196,N_19067);
nor U19210 (N_19210,N_18432,N_18972);
and U19211 (N_19211,N_18756,N_19155);
or U19212 (N_19212,N_18936,N_18534);
nand U19213 (N_19213,N_18442,N_18692);
or U19214 (N_19214,N_18548,N_18797);
or U19215 (N_19215,N_18624,N_19059);
xnor U19216 (N_19216,N_18982,N_18974);
xnor U19217 (N_19217,N_19076,N_18810);
xor U19218 (N_19218,N_18887,N_19061);
nand U19219 (N_19219,N_19037,N_19197);
or U19220 (N_19220,N_18991,N_18540);
xor U19221 (N_19221,N_18598,N_18531);
nand U19222 (N_19222,N_18473,N_18669);
or U19223 (N_19223,N_18866,N_18717);
or U19224 (N_19224,N_19122,N_19152);
nand U19225 (N_19225,N_18787,N_18819);
and U19226 (N_19226,N_18532,N_18821);
nand U19227 (N_19227,N_19169,N_19089);
nand U19228 (N_19228,N_18646,N_18783);
and U19229 (N_19229,N_19106,N_19144);
and U19230 (N_19230,N_18450,N_18460);
xor U19231 (N_19231,N_18652,N_18840);
nor U19232 (N_19232,N_19098,N_19002);
or U19233 (N_19233,N_18731,N_18685);
or U19234 (N_19234,N_18599,N_18988);
and U19235 (N_19235,N_19170,N_18916);
or U19236 (N_19236,N_18666,N_18788);
nand U19237 (N_19237,N_18488,N_18923);
or U19238 (N_19238,N_18612,N_18556);
and U19239 (N_19239,N_19014,N_18857);
or U19240 (N_19240,N_18814,N_18751);
or U19241 (N_19241,N_18523,N_18679);
nor U19242 (N_19242,N_18885,N_18808);
nor U19243 (N_19243,N_18406,N_19032);
or U19244 (N_19244,N_18914,N_18910);
and U19245 (N_19245,N_18800,N_19154);
and U19246 (N_19246,N_18948,N_18525);
or U19247 (N_19247,N_18956,N_19131);
and U19248 (N_19248,N_18513,N_18530);
nor U19249 (N_19249,N_18457,N_18941);
nor U19250 (N_19250,N_18898,N_18480);
and U19251 (N_19251,N_18594,N_19072);
nor U19252 (N_19252,N_19146,N_18777);
nor U19253 (N_19253,N_19175,N_19115);
nand U19254 (N_19254,N_19016,N_18851);
nand U19255 (N_19255,N_18820,N_18665);
xnor U19256 (N_19256,N_18932,N_18508);
xor U19257 (N_19257,N_18414,N_18909);
and U19258 (N_19258,N_18620,N_18522);
and U19259 (N_19259,N_18836,N_18673);
xnor U19260 (N_19260,N_18786,N_18763);
xnor U19261 (N_19261,N_18650,N_18767);
nand U19262 (N_19262,N_19010,N_19025);
and U19263 (N_19263,N_19086,N_18600);
xor U19264 (N_19264,N_18644,N_18519);
xnor U19265 (N_19265,N_18856,N_19109);
nor U19266 (N_19266,N_18882,N_18733);
nor U19267 (N_19267,N_18928,N_19176);
nor U19268 (N_19268,N_19100,N_19172);
xnor U19269 (N_19269,N_18430,N_19052);
and U19270 (N_19270,N_18538,N_18520);
nor U19271 (N_19271,N_19057,N_18682);
and U19272 (N_19272,N_18805,N_19163);
and U19273 (N_19273,N_19117,N_18608);
nor U19274 (N_19274,N_18455,N_18759);
nor U19275 (N_19275,N_19042,N_18554);
nor U19276 (N_19276,N_18843,N_18683);
and U19277 (N_19277,N_18438,N_18962);
and U19278 (N_19278,N_19026,N_19005);
or U19279 (N_19279,N_19049,N_18604);
and U19280 (N_19280,N_19004,N_18413);
or U19281 (N_19281,N_18785,N_18552);
nand U19282 (N_19282,N_18541,N_19195);
nor U19283 (N_19283,N_18634,N_18780);
and U19284 (N_19284,N_18891,N_18415);
xnor U19285 (N_19285,N_18636,N_18892);
xnor U19286 (N_19286,N_18574,N_19080);
nor U19287 (N_19287,N_18828,N_18509);
or U19288 (N_19288,N_19066,N_18566);
and U19289 (N_19289,N_18689,N_19095);
or U19290 (N_19290,N_18870,N_18663);
nand U19291 (N_19291,N_18605,N_18811);
or U19292 (N_19292,N_18424,N_18493);
or U19293 (N_19293,N_18651,N_19064);
nand U19294 (N_19294,N_18654,N_18755);
and U19295 (N_19295,N_18422,N_18467);
or U19296 (N_19296,N_18999,N_19027);
nand U19297 (N_19297,N_18831,N_18917);
nor U19298 (N_19298,N_19093,N_18770);
xor U19299 (N_19299,N_18497,N_18960);
xnor U19300 (N_19300,N_18639,N_18647);
or U19301 (N_19301,N_18838,N_18724);
nand U19302 (N_19302,N_18859,N_18946);
and U19303 (N_19303,N_18727,N_18533);
and U19304 (N_19304,N_18921,N_18579);
nor U19305 (N_19305,N_18589,N_18494);
and U19306 (N_19306,N_18617,N_19103);
and U19307 (N_19307,N_18485,N_18464);
and U19308 (N_19308,N_19055,N_18483);
and U19309 (N_19309,N_19185,N_19160);
nand U19310 (N_19310,N_19036,N_18908);
or U19311 (N_19311,N_18661,N_18878);
or U19312 (N_19312,N_18638,N_18569);
or U19313 (N_19313,N_18526,N_18906);
or U19314 (N_19314,N_18515,N_18436);
nor U19315 (N_19315,N_18815,N_18521);
nor U19316 (N_19316,N_18510,N_18627);
nor U19317 (N_19317,N_18401,N_18626);
nor U19318 (N_19318,N_18593,N_18935);
or U19319 (N_19319,N_18420,N_18700);
and U19320 (N_19320,N_18729,N_18897);
xnor U19321 (N_19321,N_18894,N_18772);
nand U19322 (N_19322,N_18454,N_18907);
nor U19323 (N_19323,N_18499,N_18874);
and U19324 (N_19324,N_18869,N_18789);
xnor U19325 (N_19325,N_18660,N_18730);
or U19326 (N_19326,N_19166,N_18684);
xnor U19327 (N_19327,N_18477,N_18518);
nand U19328 (N_19328,N_18681,N_18484);
and U19329 (N_19329,N_19090,N_18686);
or U19330 (N_19330,N_18744,N_18572);
nor U19331 (N_19331,N_18867,N_18606);
nand U19332 (N_19332,N_19077,N_18402);
nor U19333 (N_19333,N_18864,N_18816);
xor U19334 (N_19334,N_18969,N_19142);
xnor U19335 (N_19335,N_18721,N_18877);
nor U19336 (N_19336,N_18977,N_18975);
or U19337 (N_19337,N_18954,N_18839);
and U19338 (N_19338,N_18580,N_18938);
xor U19339 (N_19339,N_19024,N_18535);
or U19340 (N_19340,N_18913,N_18778);
nand U19341 (N_19341,N_18983,N_18451);
and U19342 (N_19342,N_18698,N_19031);
nand U19343 (N_19343,N_18970,N_18813);
or U19344 (N_19344,N_19143,N_18461);
and U19345 (N_19345,N_18668,N_18826);
and U19346 (N_19346,N_19137,N_18409);
nor U19347 (N_19347,N_18735,N_19149);
nor U19348 (N_19348,N_18746,N_18711);
xnor U19349 (N_19349,N_18794,N_18537);
nand U19350 (N_19350,N_19074,N_18680);
or U19351 (N_19351,N_18421,N_19111);
nand U19352 (N_19352,N_19132,N_18806);
or U19353 (N_19353,N_18918,N_18904);
nand U19354 (N_19354,N_18630,N_18903);
and U19355 (N_19355,N_18973,N_18996);
xor U19356 (N_19356,N_18911,N_19073);
xnor U19357 (N_19357,N_18926,N_18832);
nand U19358 (N_19358,N_18656,N_18516);
nor U19359 (N_19359,N_19127,N_18400);
nor U19360 (N_19360,N_18905,N_18912);
nor U19361 (N_19361,N_18985,N_19051);
or U19362 (N_19362,N_18490,N_18631);
nor U19363 (N_19363,N_19088,N_18582);
nor U19364 (N_19364,N_18691,N_18678);
xor U19365 (N_19365,N_18837,N_18628);
or U19366 (N_19366,N_18435,N_18674);
nand U19367 (N_19367,N_18899,N_19147);
nor U19368 (N_19368,N_18449,N_19009);
and U19369 (N_19369,N_18830,N_18703);
xor U19370 (N_19370,N_18934,N_19023);
and U19371 (N_19371,N_18944,N_18726);
and U19372 (N_19372,N_19116,N_18699);
xor U19373 (N_19373,N_18544,N_19041);
or U19374 (N_19374,N_18584,N_18774);
xnor U19375 (N_19375,N_18677,N_18981);
nand U19376 (N_19376,N_18919,N_18475);
nor U19377 (N_19377,N_18775,N_18790);
and U19378 (N_19378,N_18635,N_19112);
or U19379 (N_19379,N_18539,N_18862);
or U19380 (N_19380,N_19135,N_18971);
nor U19381 (N_19381,N_19186,N_19007);
nor U19382 (N_19382,N_18514,N_18842);
or U19383 (N_19383,N_18434,N_18920);
xor U19384 (N_19384,N_18924,N_18701);
xnor U19385 (N_19385,N_18896,N_18511);
and U19386 (N_19386,N_18459,N_18466);
and U19387 (N_19387,N_18613,N_18564);
and U19388 (N_19388,N_18667,N_19013);
nor U19389 (N_19389,N_18637,N_18444);
nand U19390 (N_19390,N_19015,N_18953);
and U19391 (N_19391,N_19164,N_19124);
nor U19392 (N_19392,N_18798,N_18633);
nand U19393 (N_19393,N_18949,N_18796);
or U19394 (N_19394,N_18618,N_18771);
and U19395 (N_19395,N_18687,N_18641);
xnor U19396 (N_19396,N_18433,N_18855);
nor U19397 (N_19397,N_18714,N_18925);
xnor U19398 (N_19398,N_19028,N_18748);
nand U19399 (N_19399,N_18448,N_18592);
nand U19400 (N_19400,N_19045,N_18712);
or U19401 (N_19401,N_19139,N_18588);
nor U19402 (N_19402,N_18583,N_18443);
nor U19403 (N_19403,N_18852,N_19012);
nor U19404 (N_19404,N_18986,N_19044);
nand U19405 (N_19405,N_18615,N_19091);
nor U19406 (N_19406,N_19017,N_18562);
nor U19407 (N_19407,N_18495,N_18884);
nand U19408 (N_19408,N_18547,N_18622);
xnor U19409 (N_19409,N_18945,N_18845);
xnor U19410 (N_19410,N_19162,N_18428);
and U19411 (N_19411,N_19157,N_19128);
nor U19412 (N_19412,N_19130,N_18479);
xor U19413 (N_19413,N_18966,N_18648);
and U19414 (N_19414,N_19123,N_18426);
nand U19415 (N_19415,N_19003,N_18690);
nand U19416 (N_19416,N_19081,N_18875);
and U19417 (N_19417,N_19168,N_18411);
and U19418 (N_19418,N_18528,N_18629);
or U19419 (N_19419,N_18792,N_19187);
and U19420 (N_19420,N_18740,N_18546);
and U19421 (N_19421,N_18706,N_18833);
xnor U19422 (N_19422,N_18964,N_18801);
or U19423 (N_19423,N_18482,N_18841);
nand U19424 (N_19424,N_19094,N_18876);
nand U19425 (N_19425,N_18848,N_18718);
xor U19426 (N_19426,N_18880,N_18616);
nand U19427 (N_19427,N_19190,N_18872);
nor U19428 (N_19428,N_19177,N_18715);
or U19429 (N_19429,N_18764,N_18462);
or U19430 (N_19430,N_18555,N_18560);
or U19431 (N_19431,N_19141,N_18978);
xnor U19432 (N_19432,N_18614,N_18559);
xnor U19433 (N_19433,N_18858,N_19110);
nand U19434 (N_19434,N_19113,N_18854);
xnor U19435 (N_19435,N_18930,N_18441);
and U19436 (N_19436,N_19039,N_18722);
xnor U19437 (N_19437,N_18591,N_19079);
xnor U19438 (N_19438,N_19034,N_18976);
xnor U19439 (N_19439,N_19192,N_18807);
and U19440 (N_19440,N_18959,N_18517);
xnor U19441 (N_19441,N_19134,N_19071);
nand U19442 (N_19442,N_18829,N_18557);
nand U19443 (N_19443,N_18824,N_18643);
nor U19444 (N_19444,N_18550,N_18809);
xnor U19445 (N_19445,N_18961,N_18445);
xnor U19446 (N_19446,N_18942,N_18645);
xor U19447 (N_19447,N_18586,N_18542);
nor U19448 (N_19448,N_19058,N_18470);
xor U19449 (N_19449,N_18403,N_18995);
and U19450 (N_19450,N_19108,N_18965);
and U19451 (N_19451,N_19158,N_18659);
nor U19452 (N_19452,N_18716,N_18781);
nand U19453 (N_19453,N_18784,N_18597);
or U19454 (N_19454,N_18407,N_18453);
and U19455 (N_19455,N_18750,N_18704);
nand U19456 (N_19456,N_18581,N_18737);
nor U19457 (N_19457,N_18883,N_19092);
xnor U19458 (N_19458,N_18922,N_18446);
and U19459 (N_19459,N_18863,N_18492);
and U19460 (N_19460,N_18505,N_18697);
and U19461 (N_19461,N_18931,N_18670);
nand U19462 (N_19462,N_19065,N_19107);
and U19463 (N_19463,N_18527,N_18452);
nand U19464 (N_19464,N_19087,N_18571);
or U19465 (N_19465,N_18768,N_18895);
nand U19466 (N_19466,N_18739,N_18871);
or U19467 (N_19467,N_19148,N_18958);
nand U19468 (N_19468,N_18500,N_18990);
or U19469 (N_19469,N_19048,N_18447);
and U19470 (N_19470,N_18861,N_19145);
xor U19471 (N_19471,N_19138,N_18947);
nand U19472 (N_19472,N_18933,N_19029);
xor U19473 (N_19473,N_18632,N_19040);
and U19474 (N_19474,N_18955,N_19000);
xnor U19475 (N_19475,N_19118,N_18927);
nand U19476 (N_19476,N_19019,N_18762);
xor U19477 (N_19477,N_18543,N_18723);
nor U19478 (N_19478,N_18468,N_19129);
nand U19479 (N_19479,N_18465,N_19191);
or U19480 (N_19480,N_18980,N_18879);
nor U19481 (N_19481,N_18760,N_19083);
nand U19482 (N_19482,N_18893,N_19193);
or U19483 (N_19483,N_18671,N_19161);
and U19484 (N_19484,N_18619,N_18553);
nand U19485 (N_19485,N_18968,N_19104);
and U19486 (N_19486,N_19022,N_18549);
or U19487 (N_19487,N_18440,N_19001);
nor U19488 (N_19488,N_18489,N_18967);
nand U19489 (N_19489,N_19174,N_19060);
nand U19490 (N_19490,N_18719,N_18749);
and U19491 (N_19491,N_18688,N_18507);
xnor U19492 (N_19492,N_18707,N_19018);
xor U19493 (N_19493,N_18994,N_18607);
xor U19494 (N_19494,N_18766,N_19078);
xor U19495 (N_19495,N_19062,N_18463);
nand U19496 (N_19496,N_19069,N_18818);
and U19497 (N_19497,N_18417,N_18412);
nor U19498 (N_19498,N_18963,N_18725);
or U19499 (N_19499,N_19167,N_19020);
and U19500 (N_19500,N_19030,N_18476);
nor U19501 (N_19501,N_18623,N_18585);
or U19502 (N_19502,N_18649,N_18405);
xor U19503 (N_19503,N_18992,N_19179);
and U19504 (N_19504,N_18577,N_18653);
nand U19505 (N_19505,N_19035,N_19084);
nor U19506 (N_19506,N_18743,N_19097);
nand U19507 (N_19507,N_19183,N_18951);
nand U19508 (N_19508,N_18793,N_19159);
xnor U19509 (N_19509,N_19038,N_19198);
and U19510 (N_19510,N_18503,N_18901);
nor U19511 (N_19511,N_18728,N_19075);
nand U19512 (N_19512,N_18950,N_19043);
xnor U19513 (N_19513,N_18802,N_18847);
or U19514 (N_19514,N_18524,N_18710);
nor U19515 (N_19515,N_18989,N_19033);
and U19516 (N_19516,N_18478,N_18757);
xor U19517 (N_19517,N_18664,N_18590);
and U19518 (N_19518,N_18803,N_19047);
xnor U19519 (N_19519,N_18625,N_18439);
xor U19520 (N_19520,N_18779,N_19194);
and U19521 (N_19521,N_18611,N_19126);
xor U19522 (N_19522,N_18957,N_18570);
and U19523 (N_19523,N_18987,N_19068);
nand U19524 (N_19524,N_19125,N_18609);
and U19525 (N_19525,N_18425,N_19165);
xor U19526 (N_19526,N_19173,N_18881);
nor U19527 (N_19527,N_19063,N_18741);
nand U19528 (N_19528,N_18596,N_18929);
or U19529 (N_19529,N_18709,N_18658);
and U19530 (N_19530,N_18695,N_18773);
nor U19531 (N_19531,N_18846,N_18745);
nand U19532 (N_19532,N_18868,N_18742);
nand U19533 (N_19533,N_19150,N_19082);
and U19534 (N_19534,N_18575,N_18886);
and U19535 (N_19535,N_18713,N_18825);
and U19536 (N_19536,N_18937,N_18416);
or U19537 (N_19537,N_18491,N_18860);
and U19538 (N_19538,N_19054,N_18782);
nand U19539 (N_19539,N_18823,N_18834);
and U19540 (N_19540,N_18952,N_18429);
nand U19541 (N_19541,N_18799,N_18850);
nor U19542 (N_19542,N_18915,N_19156);
nor U19543 (N_19543,N_18997,N_18419);
and U19544 (N_19544,N_18734,N_18993);
nor U19545 (N_19545,N_18761,N_18705);
and U19546 (N_19546,N_18979,N_18563);
or U19547 (N_19547,N_19140,N_18431);
and U19548 (N_19548,N_18754,N_18601);
or U19549 (N_19549,N_18849,N_19053);
nand U19550 (N_19550,N_18640,N_18561);
or U19551 (N_19551,N_19136,N_18873);
or U19552 (N_19552,N_18498,N_19189);
nand U19553 (N_19553,N_18418,N_18943);
nand U19554 (N_19554,N_18529,N_19151);
and U19555 (N_19555,N_19056,N_18512);
xnor U19556 (N_19556,N_19099,N_18568);
xor U19557 (N_19557,N_19006,N_19011);
nor U19558 (N_19558,N_19046,N_18736);
or U19559 (N_19559,N_18998,N_18889);
nand U19560 (N_19560,N_18693,N_18747);
xor U19561 (N_19561,N_18458,N_18939);
xor U19562 (N_19562,N_18708,N_18822);
or U19563 (N_19563,N_18456,N_18853);
nor U19564 (N_19564,N_18844,N_18642);
xor U19565 (N_19565,N_19188,N_19021);
or U19566 (N_19566,N_18481,N_18769);
and U19567 (N_19567,N_18791,N_19008);
nand U19568 (N_19568,N_18603,N_18696);
xnor U19569 (N_19569,N_19180,N_18408);
xor U19570 (N_19570,N_18984,N_18504);
and U19571 (N_19571,N_19184,N_18410);
xor U19572 (N_19572,N_19102,N_18812);
nor U19573 (N_19573,N_18423,N_18506);
or U19574 (N_19574,N_19070,N_18471);
or U19575 (N_19575,N_18587,N_19171);
xor U19576 (N_19576,N_18486,N_18758);
and U19577 (N_19577,N_18469,N_18576);
or U19578 (N_19578,N_18595,N_18437);
nand U19579 (N_19579,N_18551,N_18672);
xor U19580 (N_19580,N_19120,N_18610);
nor U19581 (N_19581,N_18776,N_18720);
nand U19582 (N_19582,N_18732,N_19153);
and U19583 (N_19583,N_18573,N_18558);
or U19584 (N_19584,N_19050,N_19121);
nand U19585 (N_19585,N_18738,N_18753);
and U19586 (N_19586,N_19114,N_19181);
and U19587 (N_19587,N_18621,N_18502);
xor U19588 (N_19588,N_18567,N_18817);
and U19589 (N_19589,N_18536,N_18675);
nand U19590 (N_19590,N_19182,N_18888);
nand U19591 (N_19591,N_19096,N_18694);
and U19592 (N_19592,N_19119,N_18404);
or U19593 (N_19593,N_18474,N_19101);
and U19594 (N_19594,N_18662,N_18655);
nand U19595 (N_19595,N_18795,N_18578);
or U19596 (N_19596,N_18940,N_18752);
nand U19597 (N_19597,N_18501,N_18602);
nor U19598 (N_19598,N_19105,N_18902);
and U19599 (N_19599,N_18545,N_18865);
nor U19600 (N_19600,N_18484,N_18444);
or U19601 (N_19601,N_18954,N_18703);
and U19602 (N_19602,N_18469,N_19190);
or U19603 (N_19603,N_18486,N_18542);
or U19604 (N_19604,N_18914,N_18887);
or U19605 (N_19605,N_19009,N_18696);
or U19606 (N_19606,N_18532,N_18924);
nand U19607 (N_19607,N_19188,N_18750);
nor U19608 (N_19608,N_18659,N_18900);
xor U19609 (N_19609,N_19165,N_18660);
xor U19610 (N_19610,N_19164,N_19020);
nor U19611 (N_19611,N_18624,N_18507);
nand U19612 (N_19612,N_18762,N_18977);
nor U19613 (N_19613,N_18565,N_18994);
xor U19614 (N_19614,N_18788,N_18731);
nor U19615 (N_19615,N_18878,N_18717);
nand U19616 (N_19616,N_18788,N_18645);
and U19617 (N_19617,N_18924,N_18822);
or U19618 (N_19618,N_18452,N_19074);
xor U19619 (N_19619,N_18602,N_18820);
nor U19620 (N_19620,N_19040,N_18834);
nand U19621 (N_19621,N_19179,N_19036);
nand U19622 (N_19622,N_18609,N_18467);
nand U19623 (N_19623,N_19198,N_18534);
xnor U19624 (N_19624,N_19023,N_18619);
and U19625 (N_19625,N_19059,N_18689);
and U19626 (N_19626,N_18989,N_18706);
and U19627 (N_19627,N_18436,N_18621);
nand U19628 (N_19628,N_19088,N_19089);
and U19629 (N_19629,N_18531,N_18492);
nor U19630 (N_19630,N_19076,N_19155);
nand U19631 (N_19631,N_18644,N_18503);
or U19632 (N_19632,N_18528,N_18720);
or U19633 (N_19633,N_18783,N_18531);
and U19634 (N_19634,N_18638,N_18508);
or U19635 (N_19635,N_18424,N_18639);
xnor U19636 (N_19636,N_18619,N_18879);
nor U19637 (N_19637,N_18416,N_19167);
nand U19638 (N_19638,N_18709,N_18578);
or U19639 (N_19639,N_18569,N_18644);
nand U19640 (N_19640,N_18604,N_18942);
xor U19641 (N_19641,N_18673,N_18501);
nand U19642 (N_19642,N_18962,N_18745);
xnor U19643 (N_19643,N_18456,N_19134);
and U19644 (N_19644,N_18882,N_19186);
and U19645 (N_19645,N_19197,N_19075);
nand U19646 (N_19646,N_18792,N_19170);
xnor U19647 (N_19647,N_18486,N_19065);
nand U19648 (N_19648,N_18748,N_19141);
xnor U19649 (N_19649,N_18508,N_18816);
or U19650 (N_19650,N_19170,N_18458);
nor U19651 (N_19651,N_19163,N_18824);
and U19652 (N_19652,N_18792,N_18975);
or U19653 (N_19653,N_18754,N_18706);
xor U19654 (N_19654,N_18679,N_19006);
nor U19655 (N_19655,N_18412,N_18658);
or U19656 (N_19656,N_19090,N_19032);
xor U19657 (N_19657,N_19034,N_18956);
and U19658 (N_19658,N_18634,N_18836);
nor U19659 (N_19659,N_18417,N_18952);
xnor U19660 (N_19660,N_18491,N_18634);
nor U19661 (N_19661,N_19114,N_18466);
or U19662 (N_19662,N_19147,N_18803);
nor U19663 (N_19663,N_19029,N_18544);
or U19664 (N_19664,N_18829,N_18816);
nor U19665 (N_19665,N_18689,N_19063);
and U19666 (N_19666,N_19165,N_18536);
nor U19667 (N_19667,N_18439,N_18556);
nand U19668 (N_19668,N_19081,N_18678);
nor U19669 (N_19669,N_19010,N_18822);
xnor U19670 (N_19670,N_18656,N_19102);
and U19671 (N_19671,N_18564,N_18512);
or U19672 (N_19672,N_18995,N_19091);
and U19673 (N_19673,N_18794,N_18605);
nand U19674 (N_19674,N_18929,N_18419);
or U19675 (N_19675,N_19029,N_19056);
nand U19676 (N_19676,N_18809,N_18600);
and U19677 (N_19677,N_19054,N_19111);
nand U19678 (N_19678,N_18695,N_19039);
nor U19679 (N_19679,N_18551,N_18901);
or U19680 (N_19680,N_18849,N_19151);
xor U19681 (N_19681,N_18443,N_18546);
nor U19682 (N_19682,N_18819,N_18633);
nor U19683 (N_19683,N_18908,N_18759);
and U19684 (N_19684,N_18823,N_18748);
and U19685 (N_19685,N_19011,N_18875);
xnor U19686 (N_19686,N_19076,N_19045);
and U19687 (N_19687,N_18487,N_18589);
or U19688 (N_19688,N_18460,N_18566);
and U19689 (N_19689,N_18894,N_18839);
or U19690 (N_19690,N_18929,N_18702);
nor U19691 (N_19691,N_19093,N_18842);
and U19692 (N_19692,N_18856,N_18567);
or U19693 (N_19693,N_19080,N_18775);
nand U19694 (N_19694,N_18754,N_18404);
and U19695 (N_19695,N_19061,N_19011);
or U19696 (N_19696,N_19085,N_18692);
and U19697 (N_19697,N_18573,N_18832);
nand U19698 (N_19698,N_19065,N_18894);
or U19699 (N_19699,N_18640,N_18694);
and U19700 (N_19700,N_18616,N_18477);
nand U19701 (N_19701,N_19028,N_18854);
xnor U19702 (N_19702,N_18784,N_19147);
nor U19703 (N_19703,N_18990,N_18594);
nor U19704 (N_19704,N_18751,N_18957);
or U19705 (N_19705,N_18960,N_18440);
xnor U19706 (N_19706,N_18561,N_19105);
xor U19707 (N_19707,N_18758,N_19047);
or U19708 (N_19708,N_19114,N_19005);
nor U19709 (N_19709,N_18420,N_18566);
xor U19710 (N_19710,N_18994,N_19123);
nand U19711 (N_19711,N_18536,N_18725);
and U19712 (N_19712,N_18615,N_19095);
nor U19713 (N_19713,N_19011,N_18848);
and U19714 (N_19714,N_19092,N_18991);
nand U19715 (N_19715,N_19012,N_18663);
or U19716 (N_19716,N_18408,N_18575);
nand U19717 (N_19717,N_19037,N_18721);
nand U19718 (N_19718,N_18421,N_18569);
nor U19719 (N_19719,N_18664,N_18848);
and U19720 (N_19720,N_18493,N_19132);
nor U19721 (N_19721,N_18977,N_18919);
or U19722 (N_19722,N_19041,N_18883);
and U19723 (N_19723,N_18868,N_19106);
nand U19724 (N_19724,N_18579,N_19083);
nor U19725 (N_19725,N_18643,N_18541);
or U19726 (N_19726,N_18936,N_18563);
nand U19727 (N_19727,N_19050,N_18550);
nor U19728 (N_19728,N_18437,N_18867);
nor U19729 (N_19729,N_19168,N_19099);
nor U19730 (N_19730,N_18954,N_18530);
and U19731 (N_19731,N_18947,N_19068);
and U19732 (N_19732,N_18906,N_19154);
and U19733 (N_19733,N_18420,N_18699);
nor U19734 (N_19734,N_19070,N_18621);
nand U19735 (N_19735,N_19047,N_18551);
xor U19736 (N_19736,N_18842,N_18455);
xor U19737 (N_19737,N_19092,N_18870);
and U19738 (N_19738,N_19024,N_18687);
xor U19739 (N_19739,N_18499,N_18611);
or U19740 (N_19740,N_18616,N_18580);
and U19741 (N_19741,N_18471,N_19098);
or U19742 (N_19742,N_19114,N_18862);
xnor U19743 (N_19743,N_18743,N_18778);
nand U19744 (N_19744,N_19175,N_19070);
nor U19745 (N_19745,N_18734,N_19168);
nand U19746 (N_19746,N_18620,N_19094);
nor U19747 (N_19747,N_19186,N_19013);
nand U19748 (N_19748,N_18936,N_19142);
and U19749 (N_19749,N_18847,N_18481);
or U19750 (N_19750,N_19033,N_18521);
nor U19751 (N_19751,N_18507,N_18825);
and U19752 (N_19752,N_19107,N_18442);
and U19753 (N_19753,N_18549,N_18412);
or U19754 (N_19754,N_18500,N_18510);
and U19755 (N_19755,N_18788,N_18496);
xor U19756 (N_19756,N_18649,N_19188);
xor U19757 (N_19757,N_19142,N_18896);
and U19758 (N_19758,N_19009,N_18514);
xor U19759 (N_19759,N_19116,N_18599);
or U19760 (N_19760,N_18618,N_19192);
or U19761 (N_19761,N_18850,N_18597);
or U19762 (N_19762,N_18810,N_18498);
nor U19763 (N_19763,N_18644,N_18937);
nand U19764 (N_19764,N_19062,N_18944);
and U19765 (N_19765,N_18466,N_18893);
nand U19766 (N_19766,N_18927,N_18571);
nand U19767 (N_19767,N_18843,N_19065);
nand U19768 (N_19768,N_18895,N_19117);
nor U19769 (N_19769,N_18731,N_19016);
nand U19770 (N_19770,N_18488,N_19125);
xor U19771 (N_19771,N_18826,N_18576);
xnor U19772 (N_19772,N_19138,N_18671);
nand U19773 (N_19773,N_18949,N_18975);
nand U19774 (N_19774,N_18430,N_19029);
nor U19775 (N_19775,N_19110,N_19001);
nor U19776 (N_19776,N_18985,N_18813);
nor U19777 (N_19777,N_18565,N_18768);
nand U19778 (N_19778,N_18882,N_18931);
xnor U19779 (N_19779,N_18704,N_18621);
xor U19780 (N_19780,N_18931,N_18754);
or U19781 (N_19781,N_18832,N_18949);
or U19782 (N_19782,N_18769,N_18535);
nand U19783 (N_19783,N_19112,N_19120);
and U19784 (N_19784,N_18861,N_18440);
and U19785 (N_19785,N_18922,N_18564);
nand U19786 (N_19786,N_19176,N_19172);
nor U19787 (N_19787,N_19009,N_18791);
nand U19788 (N_19788,N_18774,N_18882);
nor U19789 (N_19789,N_18521,N_18948);
and U19790 (N_19790,N_18559,N_18528);
nor U19791 (N_19791,N_18539,N_18418);
or U19792 (N_19792,N_18794,N_18416);
and U19793 (N_19793,N_18772,N_18736);
or U19794 (N_19794,N_18896,N_18833);
nor U19795 (N_19795,N_18671,N_18405);
and U19796 (N_19796,N_18920,N_18575);
nand U19797 (N_19797,N_19192,N_19067);
xor U19798 (N_19798,N_18830,N_18970);
and U19799 (N_19799,N_18717,N_18545);
nor U19800 (N_19800,N_18645,N_18561);
nand U19801 (N_19801,N_19107,N_19087);
nor U19802 (N_19802,N_18963,N_18459);
xor U19803 (N_19803,N_18793,N_18644);
nand U19804 (N_19804,N_19132,N_18999);
nor U19805 (N_19805,N_19021,N_18698);
and U19806 (N_19806,N_19144,N_19025);
nand U19807 (N_19807,N_18566,N_18873);
and U19808 (N_19808,N_19176,N_18748);
xnor U19809 (N_19809,N_18785,N_19194);
or U19810 (N_19810,N_18971,N_18470);
and U19811 (N_19811,N_18759,N_18510);
nand U19812 (N_19812,N_18527,N_18886);
xor U19813 (N_19813,N_18575,N_18472);
or U19814 (N_19814,N_18693,N_18460);
nor U19815 (N_19815,N_18635,N_18845);
or U19816 (N_19816,N_18639,N_18791);
or U19817 (N_19817,N_18900,N_18434);
nand U19818 (N_19818,N_18946,N_18593);
xor U19819 (N_19819,N_18964,N_18979);
and U19820 (N_19820,N_18772,N_18870);
or U19821 (N_19821,N_18521,N_18863);
and U19822 (N_19822,N_18496,N_18481);
nand U19823 (N_19823,N_18588,N_18622);
nor U19824 (N_19824,N_18501,N_19182);
xnor U19825 (N_19825,N_19091,N_18631);
nor U19826 (N_19826,N_18627,N_18615);
xnor U19827 (N_19827,N_19028,N_19041);
and U19828 (N_19828,N_18413,N_18409);
nor U19829 (N_19829,N_18575,N_18740);
xnor U19830 (N_19830,N_18862,N_18555);
nand U19831 (N_19831,N_18838,N_18914);
nor U19832 (N_19832,N_18543,N_19014);
and U19833 (N_19833,N_18835,N_18767);
nand U19834 (N_19834,N_18471,N_18560);
and U19835 (N_19835,N_18717,N_18972);
or U19836 (N_19836,N_18787,N_18546);
nor U19837 (N_19837,N_18855,N_18574);
nor U19838 (N_19838,N_18483,N_18558);
nor U19839 (N_19839,N_18506,N_18490);
nand U19840 (N_19840,N_18970,N_18853);
or U19841 (N_19841,N_19178,N_19104);
nor U19842 (N_19842,N_18723,N_18457);
and U19843 (N_19843,N_18914,N_19046);
or U19844 (N_19844,N_18677,N_18838);
xor U19845 (N_19845,N_18794,N_18739);
nand U19846 (N_19846,N_18655,N_18899);
or U19847 (N_19847,N_18619,N_18909);
and U19848 (N_19848,N_18650,N_18499);
and U19849 (N_19849,N_18831,N_19012);
or U19850 (N_19850,N_18683,N_19143);
nor U19851 (N_19851,N_18474,N_19084);
nand U19852 (N_19852,N_18711,N_18406);
and U19853 (N_19853,N_19180,N_18547);
or U19854 (N_19854,N_19088,N_18557);
nor U19855 (N_19855,N_18783,N_19017);
or U19856 (N_19856,N_18672,N_19125);
or U19857 (N_19857,N_18981,N_18691);
or U19858 (N_19858,N_19113,N_19185);
xor U19859 (N_19859,N_18627,N_18961);
or U19860 (N_19860,N_18405,N_18461);
nand U19861 (N_19861,N_18755,N_18737);
nand U19862 (N_19862,N_19078,N_18723);
xor U19863 (N_19863,N_18511,N_19117);
or U19864 (N_19864,N_19126,N_18987);
nor U19865 (N_19865,N_19136,N_18578);
or U19866 (N_19866,N_18493,N_18952);
xor U19867 (N_19867,N_18482,N_18917);
or U19868 (N_19868,N_19132,N_18866);
nand U19869 (N_19869,N_19012,N_18640);
and U19870 (N_19870,N_18843,N_18438);
or U19871 (N_19871,N_19190,N_18506);
nand U19872 (N_19872,N_18462,N_18713);
xor U19873 (N_19873,N_18516,N_18770);
xor U19874 (N_19874,N_18686,N_19081);
xor U19875 (N_19875,N_19113,N_18967);
or U19876 (N_19876,N_18622,N_18729);
nor U19877 (N_19877,N_19007,N_18699);
nand U19878 (N_19878,N_18528,N_18448);
xor U19879 (N_19879,N_18725,N_18851);
nand U19880 (N_19880,N_18808,N_18497);
nand U19881 (N_19881,N_18669,N_18807);
nand U19882 (N_19882,N_18733,N_18665);
or U19883 (N_19883,N_18558,N_18930);
nor U19884 (N_19884,N_18520,N_18418);
and U19885 (N_19885,N_18452,N_18570);
and U19886 (N_19886,N_19192,N_19032);
nand U19887 (N_19887,N_18662,N_18444);
nand U19888 (N_19888,N_18868,N_19061);
or U19889 (N_19889,N_18625,N_18507);
nor U19890 (N_19890,N_18976,N_18895);
xor U19891 (N_19891,N_18909,N_18561);
and U19892 (N_19892,N_18669,N_18868);
and U19893 (N_19893,N_18769,N_18774);
nand U19894 (N_19894,N_19175,N_19191);
or U19895 (N_19895,N_18774,N_18792);
xnor U19896 (N_19896,N_18544,N_18449);
nor U19897 (N_19897,N_18526,N_18657);
and U19898 (N_19898,N_18674,N_18990);
xnor U19899 (N_19899,N_18551,N_18502);
or U19900 (N_19900,N_19033,N_19051);
or U19901 (N_19901,N_18463,N_18497);
nor U19902 (N_19902,N_18884,N_18923);
xor U19903 (N_19903,N_18674,N_19056);
nor U19904 (N_19904,N_18532,N_18431);
or U19905 (N_19905,N_18579,N_18751);
xnor U19906 (N_19906,N_19158,N_18472);
or U19907 (N_19907,N_18799,N_18832);
or U19908 (N_19908,N_19095,N_19122);
xnor U19909 (N_19909,N_19036,N_18609);
and U19910 (N_19910,N_19164,N_18670);
or U19911 (N_19911,N_18549,N_18955);
and U19912 (N_19912,N_18893,N_18440);
nor U19913 (N_19913,N_18972,N_18981);
and U19914 (N_19914,N_18514,N_18439);
nand U19915 (N_19915,N_18502,N_18701);
nand U19916 (N_19916,N_18421,N_18872);
nor U19917 (N_19917,N_18617,N_19163);
nand U19918 (N_19918,N_18417,N_19029);
nor U19919 (N_19919,N_19014,N_18578);
nor U19920 (N_19920,N_19014,N_18549);
xor U19921 (N_19921,N_18625,N_19096);
nand U19922 (N_19922,N_18634,N_18921);
and U19923 (N_19923,N_18612,N_18598);
or U19924 (N_19924,N_19127,N_18966);
nor U19925 (N_19925,N_18653,N_18840);
nand U19926 (N_19926,N_18743,N_18537);
nor U19927 (N_19927,N_19143,N_18978);
or U19928 (N_19928,N_18907,N_18408);
nand U19929 (N_19929,N_18491,N_18432);
or U19930 (N_19930,N_18917,N_19186);
nand U19931 (N_19931,N_18742,N_18622);
xnor U19932 (N_19932,N_18584,N_18529);
xnor U19933 (N_19933,N_19140,N_18705);
and U19934 (N_19934,N_19138,N_18926);
nand U19935 (N_19935,N_19053,N_18555);
or U19936 (N_19936,N_18881,N_18923);
xnor U19937 (N_19937,N_18890,N_19139);
xor U19938 (N_19938,N_18696,N_18565);
xor U19939 (N_19939,N_18730,N_18835);
and U19940 (N_19940,N_18760,N_18521);
xor U19941 (N_19941,N_18711,N_19080);
nand U19942 (N_19942,N_18780,N_18502);
or U19943 (N_19943,N_18843,N_18961);
or U19944 (N_19944,N_18891,N_18713);
nor U19945 (N_19945,N_18724,N_18888);
xnor U19946 (N_19946,N_18657,N_18954);
nand U19947 (N_19947,N_18577,N_18918);
xor U19948 (N_19948,N_18718,N_18424);
nor U19949 (N_19949,N_18613,N_18860);
and U19950 (N_19950,N_19054,N_18644);
and U19951 (N_19951,N_19105,N_18924);
and U19952 (N_19952,N_18701,N_18932);
xnor U19953 (N_19953,N_19051,N_18974);
xnor U19954 (N_19954,N_19028,N_18784);
nand U19955 (N_19955,N_18809,N_18721);
xnor U19956 (N_19956,N_18735,N_18930);
or U19957 (N_19957,N_18830,N_18710);
and U19958 (N_19958,N_18998,N_18785);
or U19959 (N_19959,N_18746,N_19021);
nor U19960 (N_19960,N_18735,N_18999);
and U19961 (N_19961,N_18935,N_18774);
xor U19962 (N_19962,N_18745,N_18667);
or U19963 (N_19963,N_18540,N_19108);
xor U19964 (N_19964,N_18904,N_18403);
and U19965 (N_19965,N_18644,N_18877);
or U19966 (N_19966,N_18663,N_18628);
nand U19967 (N_19967,N_19189,N_18652);
or U19968 (N_19968,N_18924,N_18642);
or U19969 (N_19969,N_18617,N_18772);
or U19970 (N_19970,N_18558,N_18920);
or U19971 (N_19971,N_18766,N_18793);
xor U19972 (N_19972,N_18578,N_18608);
and U19973 (N_19973,N_18493,N_18569);
nand U19974 (N_19974,N_18605,N_18504);
xnor U19975 (N_19975,N_18778,N_18439);
nor U19976 (N_19976,N_19025,N_19066);
nor U19977 (N_19977,N_18567,N_18711);
and U19978 (N_19978,N_18878,N_19188);
and U19979 (N_19979,N_19024,N_18799);
nor U19980 (N_19980,N_18977,N_18695);
and U19981 (N_19981,N_19009,N_19022);
nand U19982 (N_19982,N_18985,N_18493);
nand U19983 (N_19983,N_18772,N_19078);
and U19984 (N_19984,N_19020,N_18457);
and U19985 (N_19985,N_19147,N_18638);
or U19986 (N_19986,N_19185,N_18641);
nand U19987 (N_19987,N_18615,N_18481);
or U19988 (N_19988,N_18643,N_18901);
nor U19989 (N_19989,N_19194,N_19131);
nand U19990 (N_19990,N_18797,N_18749);
and U19991 (N_19991,N_19166,N_19103);
and U19992 (N_19992,N_18824,N_18613);
and U19993 (N_19993,N_18608,N_18563);
nand U19994 (N_19994,N_18674,N_18903);
and U19995 (N_19995,N_18883,N_18752);
nand U19996 (N_19996,N_19043,N_19158);
nor U19997 (N_19997,N_18984,N_19087);
nand U19998 (N_19998,N_19059,N_19067);
nand U19999 (N_19999,N_18645,N_18659);
or UO_0 (O_0,N_19469,N_19844);
nand UO_1 (O_1,N_19712,N_19432);
and UO_2 (O_2,N_19471,N_19453);
or UO_3 (O_3,N_19731,N_19276);
nor UO_4 (O_4,N_19609,N_19880);
nand UO_5 (O_5,N_19689,N_19327);
nor UO_6 (O_6,N_19328,N_19672);
or UO_7 (O_7,N_19636,N_19948);
nand UO_8 (O_8,N_19785,N_19748);
nor UO_9 (O_9,N_19598,N_19778);
xor UO_10 (O_10,N_19898,N_19299);
nand UO_11 (O_11,N_19373,N_19938);
nor UO_12 (O_12,N_19615,N_19631);
and UO_13 (O_13,N_19370,N_19462);
nor UO_14 (O_14,N_19901,N_19539);
or UO_15 (O_15,N_19547,N_19380);
and UO_16 (O_16,N_19679,N_19542);
nand UO_17 (O_17,N_19915,N_19703);
nand UO_18 (O_18,N_19757,N_19916);
xnor UO_19 (O_19,N_19979,N_19805);
nand UO_20 (O_20,N_19696,N_19570);
nand UO_21 (O_21,N_19217,N_19945);
or UO_22 (O_22,N_19498,N_19552);
or UO_23 (O_23,N_19999,N_19486);
and UO_24 (O_24,N_19518,N_19808);
nor UO_25 (O_25,N_19993,N_19905);
nand UO_26 (O_26,N_19566,N_19933);
nand UO_27 (O_27,N_19378,N_19216);
or UO_28 (O_28,N_19337,N_19209);
nand UO_29 (O_29,N_19681,N_19253);
and UO_30 (O_30,N_19887,N_19418);
and UO_31 (O_31,N_19258,N_19387);
nand UO_32 (O_32,N_19761,N_19798);
xor UO_33 (O_33,N_19569,N_19245);
xnor UO_34 (O_34,N_19708,N_19357);
and UO_35 (O_35,N_19336,N_19807);
xnor UO_36 (O_36,N_19751,N_19333);
nor UO_37 (O_37,N_19838,N_19830);
nor UO_38 (O_38,N_19316,N_19446);
nor UO_39 (O_39,N_19958,N_19946);
and UO_40 (O_40,N_19727,N_19740);
or UO_41 (O_41,N_19802,N_19300);
nor UO_42 (O_42,N_19558,N_19226);
nand UO_43 (O_43,N_19580,N_19416);
nor UO_44 (O_44,N_19579,N_19350);
or UO_45 (O_45,N_19991,N_19629);
and UO_46 (O_46,N_19725,N_19526);
nand UO_47 (O_47,N_19787,N_19275);
and UO_48 (O_48,N_19829,N_19438);
or UO_49 (O_49,N_19487,N_19235);
nand UO_50 (O_50,N_19595,N_19641);
or UO_51 (O_51,N_19674,N_19866);
nand UO_52 (O_52,N_19967,N_19291);
nand UO_53 (O_53,N_19450,N_19826);
or UO_54 (O_54,N_19252,N_19698);
and UO_55 (O_55,N_19667,N_19799);
and UO_56 (O_56,N_19415,N_19989);
xnor UO_57 (O_57,N_19367,N_19458);
or UO_58 (O_58,N_19496,N_19995);
nor UO_59 (O_59,N_19814,N_19369);
or UO_60 (O_60,N_19335,N_19825);
or UO_61 (O_61,N_19861,N_19356);
and UO_62 (O_62,N_19746,N_19288);
and UO_63 (O_63,N_19535,N_19957);
xnor UO_64 (O_64,N_19943,N_19326);
or UO_65 (O_65,N_19764,N_19540);
or UO_66 (O_66,N_19640,N_19318);
nor UO_67 (O_67,N_19922,N_19550);
nand UO_68 (O_68,N_19665,N_19472);
xor UO_69 (O_69,N_19319,N_19914);
or UO_70 (O_70,N_19515,N_19308);
xnor UO_71 (O_71,N_19225,N_19243);
xnor UO_72 (O_72,N_19514,N_19315);
nand UO_73 (O_73,N_19573,N_19788);
nand UO_74 (O_74,N_19634,N_19488);
and UO_75 (O_75,N_19295,N_19951);
xnor UO_76 (O_76,N_19375,N_19613);
nand UO_77 (O_77,N_19544,N_19855);
xnor UO_78 (O_78,N_19507,N_19841);
nand UO_79 (O_79,N_19200,N_19256);
and UO_80 (O_80,N_19289,N_19988);
xor UO_81 (O_81,N_19931,N_19668);
xnor UO_82 (O_82,N_19351,N_19242);
nand UO_83 (O_83,N_19965,N_19831);
xor UO_84 (O_84,N_19341,N_19459);
xnor UO_85 (O_85,N_19846,N_19893);
nor UO_86 (O_86,N_19571,N_19647);
and UO_87 (O_87,N_19497,N_19524);
nor UO_88 (O_88,N_19810,N_19714);
and UO_89 (O_89,N_19403,N_19968);
or UO_90 (O_90,N_19690,N_19301);
nand UO_91 (O_91,N_19833,N_19424);
nand UO_92 (O_92,N_19221,N_19870);
and UO_93 (O_93,N_19441,N_19924);
xnor UO_94 (O_94,N_19549,N_19456);
or UO_95 (O_95,N_19448,N_19440);
nor UO_96 (O_96,N_19952,N_19412);
nor UO_97 (O_97,N_19966,N_19695);
nand UO_98 (O_98,N_19207,N_19425);
and UO_99 (O_99,N_19774,N_19651);
nor UO_100 (O_100,N_19240,N_19919);
and UO_101 (O_101,N_19331,N_19669);
or UO_102 (O_102,N_19902,N_19590);
nand UO_103 (O_103,N_19710,N_19345);
nand UO_104 (O_104,N_19869,N_19232);
or UO_105 (O_105,N_19509,N_19859);
or UO_106 (O_106,N_19494,N_19280);
xor UO_107 (O_107,N_19892,N_19974);
nand UO_108 (O_108,N_19700,N_19447);
or UO_109 (O_109,N_19852,N_19972);
or UO_110 (O_110,N_19863,N_19652);
nor UO_111 (O_111,N_19741,N_19281);
nor UO_112 (O_112,N_19950,N_19692);
and UO_113 (O_113,N_19560,N_19675);
or UO_114 (O_114,N_19660,N_19398);
and UO_115 (O_115,N_19793,N_19208);
or UO_116 (O_116,N_19728,N_19546);
nand UO_117 (O_117,N_19928,N_19682);
or UO_118 (O_118,N_19865,N_19934);
xor UO_119 (O_119,N_19603,N_19791);
xor UO_120 (O_120,N_19231,N_19278);
nand UO_121 (O_121,N_19997,N_19267);
xor UO_122 (O_122,N_19873,N_19426);
or UO_123 (O_123,N_19666,N_19658);
or UO_124 (O_124,N_19474,N_19437);
and UO_125 (O_125,N_19739,N_19930);
and UO_126 (O_126,N_19586,N_19720);
and UO_127 (O_127,N_19929,N_19954);
nor UO_128 (O_128,N_19904,N_19449);
xnor UO_129 (O_129,N_19320,N_19639);
and UO_130 (O_130,N_19685,N_19721);
nor UO_131 (O_131,N_19860,N_19342);
nor UO_132 (O_132,N_19747,N_19955);
or UO_133 (O_133,N_19628,N_19877);
or UO_134 (O_134,N_19619,N_19274);
or UO_135 (O_135,N_19532,N_19935);
and UO_136 (O_136,N_19287,N_19352);
nor UO_137 (O_137,N_19214,N_19963);
xor UO_138 (O_138,N_19385,N_19557);
nor UO_139 (O_139,N_19769,N_19349);
and UO_140 (O_140,N_19980,N_19466);
and UO_141 (O_141,N_19545,N_19875);
nor UO_142 (O_142,N_19597,N_19277);
and UO_143 (O_143,N_19358,N_19238);
nor UO_144 (O_144,N_19390,N_19325);
nand UO_145 (O_145,N_19523,N_19971);
nand UO_146 (O_146,N_19854,N_19874);
nor UO_147 (O_147,N_19835,N_19562);
and UO_148 (O_148,N_19427,N_19491);
nand UO_149 (O_149,N_19251,N_19864);
nand UO_150 (O_150,N_19484,N_19400);
nand UO_151 (O_151,N_19576,N_19306);
or UO_152 (O_152,N_19797,N_19789);
nor UO_153 (O_153,N_19722,N_19563);
nor UO_154 (O_154,N_19559,N_19848);
nor UO_155 (O_155,N_19286,N_19699);
or UO_156 (O_156,N_19229,N_19502);
nor UO_157 (O_157,N_19812,N_19673);
or UO_158 (O_158,N_19436,N_19405);
and UO_159 (O_159,N_19719,N_19978);
and UO_160 (O_160,N_19511,N_19371);
or UO_161 (O_161,N_19409,N_19305);
nor UO_162 (O_162,N_19269,N_19454);
nor UO_163 (O_163,N_19606,N_19917);
nor UO_164 (O_164,N_19994,N_19876);
or UO_165 (O_165,N_19953,N_19885);
xnor UO_166 (O_166,N_19733,N_19348);
or UO_167 (O_167,N_19813,N_19768);
xnor UO_168 (O_168,N_19470,N_19536);
nor UO_169 (O_169,N_19605,N_19364);
xnor UO_170 (O_170,N_19617,N_19816);
nand UO_171 (O_171,N_19961,N_19399);
or UO_172 (O_172,N_19483,N_19604);
nor UO_173 (O_173,N_19265,N_19411);
xor UO_174 (O_174,N_19384,N_19332);
or UO_175 (O_175,N_19659,N_19250);
or UO_176 (O_176,N_19975,N_19766);
and UO_177 (O_177,N_19827,N_19244);
xor UO_178 (O_178,N_19255,N_19910);
and UO_179 (O_179,N_19777,N_19479);
nand UO_180 (O_180,N_19588,N_19693);
nor UO_181 (O_181,N_19611,N_19804);
nor UO_182 (O_182,N_19969,N_19402);
nand UO_183 (O_183,N_19589,N_19849);
and UO_184 (O_184,N_19445,N_19435);
xor UO_185 (O_185,N_19422,N_19803);
or UO_186 (O_186,N_19581,N_19260);
nand UO_187 (O_187,N_19460,N_19656);
or UO_188 (O_188,N_19261,N_19688);
nor UO_189 (O_189,N_19944,N_19836);
nor UO_190 (O_190,N_19763,N_19233);
xor UO_191 (O_191,N_19664,N_19346);
nor UO_192 (O_192,N_19821,N_19879);
nor UO_193 (O_193,N_19900,N_19554);
xnor UO_194 (O_194,N_19284,N_19780);
and UO_195 (O_195,N_19420,N_19537);
nand UO_196 (O_196,N_19354,N_19285);
xnor UO_197 (O_197,N_19556,N_19670);
xnor UO_198 (O_198,N_19775,N_19361);
nor UO_199 (O_199,N_19294,N_19249);
nor UO_200 (O_200,N_19809,N_19851);
or UO_201 (O_201,N_19223,N_19247);
or UO_202 (O_202,N_19272,N_19429);
or UO_203 (O_203,N_19266,N_19213);
and UO_204 (O_204,N_19646,N_19786);
nor UO_205 (O_205,N_19417,N_19467);
nor UO_206 (O_206,N_19206,N_19282);
nor UO_207 (O_207,N_19947,N_19228);
nor UO_208 (O_208,N_19843,N_19800);
xnor UO_209 (O_209,N_19921,N_19822);
nand UO_210 (O_210,N_19618,N_19414);
nand UO_211 (O_211,N_19531,N_19239);
nor UO_212 (O_212,N_19762,N_19505);
xnor UO_213 (O_213,N_19686,N_19891);
or UO_214 (O_214,N_19745,N_19736);
nor UO_215 (O_215,N_19510,N_19599);
xnor UO_216 (O_216,N_19959,N_19362);
xor UO_217 (O_217,N_19401,N_19704);
and UO_218 (O_218,N_19729,N_19625);
nand UO_219 (O_219,N_19302,N_19832);
nor UO_220 (O_220,N_19663,N_19324);
or UO_221 (O_221,N_19476,N_19592);
xor UO_222 (O_222,N_19464,N_19273);
xnor UO_223 (O_223,N_19713,N_19224);
or UO_224 (O_224,N_19311,N_19339);
or UO_225 (O_225,N_19886,N_19477);
or UO_226 (O_226,N_19584,N_19899);
nor UO_227 (O_227,N_19754,N_19998);
or UO_228 (O_228,N_19270,N_19632);
nand UO_229 (O_229,N_19527,N_19386);
and UO_230 (O_230,N_19205,N_19372);
and UO_231 (O_231,N_19977,N_19796);
and UO_232 (O_232,N_19428,N_19707);
xnor UO_233 (O_233,N_19530,N_19680);
xnor UO_234 (O_234,N_19872,N_19819);
nand UO_235 (O_235,N_19926,N_19219);
and UO_236 (O_236,N_19858,N_19338);
nor UO_237 (O_237,N_19795,N_19732);
nor UO_238 (O_238,N_19406,N_19726);
xnor UO_239 (O_239,N_19622,N_19254);
and UO_240 (O_240,N_19212,N_19443);
xor UO_241 (O_241,N_19347,N_19577);
nor UO_242 (O_242,N_19633,N_19455);
and UO_243 (O_243,N_19236,N_19382);
xnor UO_244 (O_244,N_19850,N_19987);
nand UO_245 (O_245,N_19936,N_19723);
and UO_246 (O_246,N_19779,N_19594);
nand UO_247 (O_247,N_19653,N_19990);
nor UO_248 (O_248,N_19635,N_19313);
and UO_249 (O_249,N_19396,N_19508);
or UO_250 (O_250,N_19730,N_19837);
or UO_251 (O_251,N_19734,N_19492);
nand UO_252 (O_252,N_19890,N_19574);
nor UO_253 (O_253,N_19434,N_19564);
xor UO_254 (O_254,N_19490,N_19596);
or UO_255 (O_255,N_19587,N_19343);
nor UO_256 (O_256,N_19442,N_19627);
nand UO_257 (O_257,N_19363,N_19772);
nand UO_258 (O_258,N_19478,N_19237);
xor UO_259 (O_259,N_19909,N_19908);
and UO_260 (O_260,N_19828,N_19701);
xor UO_261 (O_261,N_19355,N_19533);
nor UO_262 (O_262,N_19374,N_19475);
and UO_263 (O_263,N_19495,N_19612);
xnor UO_264 (O_264,N_19662,N_19884);
nor UO_265 (O_265,N_19623,N_19691);
xor UO_266 (O_266,N_19842,N_19578);
nand UO_267 (O_267,N_19702,N_19918);
and UO_268 (O_268,N_19461,N_19824);
xnor UO_269 (O_269,N_19407,N_19624);
nor UO_270 (O_270,N_19867,N_19290);
and UO_271 (O_271,N_19368,N_19257);
nor UO_272 (O_272,N_19776,N_19894);
xor UO_273 (O_273,N_19329,N_19655);
xor UO_274 (O_274,N_19616,N_19585);
or UO_275 (O_275,N_19684,N_19735);
or UO_276 (O_276,N_19521,N_19310);
and UO_277 (O_277,N_19984,N_19847);
or UO_278 (O_278,N_19561,N_19264);
and UO_279 (O_279,N_19465,N_19283);
nor UO_280 (O_280,N_19481,N_19431);
nor UO_281 (O_281,N_19293,N_19397);
nor UO_282 (O_282,N_19230,N_19582);
nand UO_283 (O_283,N_19503,N_19755);
and UO_284 (O_284,N_19985,N_19365);
nand UO_285 (O_285,N_19381,N_19962);
xor UO_286 (O_286,N_19608,N_19697);
and UO_287 (O_287,N_19379,N_19304);
nand UO_288 (O_288,N_19419,N_19642);
nand UO_289 (O_289,N_19408,N_19742);
and UO_290 (O_290,N_19519,N_19897);
nor UO_291 (O_291,N_19705,N_19648);
xor UO_292 (O_292,N_19782,N_19234);
and UO_293 (O_293,N_19210,N_19413);
and UO_294 (O_294,N_19610,N_19303);
nor UO_295 (O_295,N_19575,N_19359);
xnor UO_296 (O_296,N_19657,N_19949);
and UO_297 (O_297,N_19394,N_19340);
or UO_298 (O_298,N_19218,N_19932);
and UO_299 (O_299,N_19840,N_19759);
nand UO_300 (O_300,N_19906,N_19683);
xnor UO_301 (O_301,N_19749,N_19551);
or UO_302 (O_302,N_19202,N_19907);
xnor UO_303 (O_303,N_19925,N_19882);
nand UO_304 (O_304,N_19553,N_19353);
nand UO_305 (O_305,N_19499,N_19312);
or UO_306 (O_306,N_19555,N_19687);
and UO_307 (O_307,N_19820,N_19806);
nand UO_308 (O_308,N_19856,N_19493);
xnor UO_309 (O_309,N_19377,N_19716);
xor UO_310 (O_310,N_19942,N_19473);
and UO_311 (O_311,N_19292,N_19981);
xnor UO_312 (O_312,N_19970,N_19996);
xnor UO_313 (O_313,N_19637,N_19323);
nand UO_314 (O_314,N_19792,N_19896);
or UO_315 (O_315,N_19489,N_19259);
nand UO_316 (O_316,N_19204,N_19548);
and UO_317 (O_317,N_19522,N_19423);
or UO_318 (O_318,N_19817,N_19534);
nand UO_319 (O_319,N_19927,N_19645);
or UO_320 (O_320,N_19528,N_19621);
xor UO_321 (O_321,N_19334,N_19601);
xor UO_322 (O_322,N_19773,N_19767);
xor UO_323 (O_323,N_19889,N_19392);
or UO_324 (O_324,N_19433,N_19718);
or UO_325 (O_325,N_19878,N_19868);
nor UO_326 (O_326,N_19593,N_19976);
or UO_327 (O_327,N_19992,N_19451);
and UO_328 (O_328,N_19818,N_19983);
nor UO_329 (O_329,N_19541,N_19602);
and UO_330 (O_330,N_19706,N_19485);
nor UO_331 (O_331,N_19583,N_19752);
nor UO_332 (O_332,N_19794,N_19643);
and UO_333 (O_333,N_19895,N_19383);
and UO_334 (O_334,N_19737,N_19463);
and UO_335 (O_335,N_19600,N_19750);
nand UO_336 (O_336,N_19517,N_19516);
xor UO_337 (O_337,N_19314,N_19421);
and UO_338 (O_338,N_19614,N_19676);
xnor UO_339 (O_339,N_19650,N_19939);
nor UO_340 (O_340,N_19709,N_19630);
nand UO_341 (O_341,N_19543,N_19538);
nand UO_342 (O_342,N_19638,N_19201);
or UO_343 (O_343,N_19694,N_19724);
or UO_344 (O_344,N_19923,N_19279);
nand UO_345 (O_345,N_19626,N_19760);
nand UO_346 (O_346,N_19388,N_19321);
or UO_347 (O_347,N_19389,N_19771);
xnor UO_348 (O_348,N_19513,N_19940);
nor UO_349 (O_349,N_19986,N_19317);
xnor UO_350 (O_350,N_19956,N_19607);
and UO_351 (O_351,N_19360,N_19964);
nand UO_352 (O_352,N_19220,N_19911);
xor UO_353 (O_353,N_19262,N_19444);
xnor UO_354 (O_354,N_19823,N_19883);
nor UO_355 (O_355,N_19982,N_19565);
nand UO_356 (O_356,N_19529,N_19717);
or UO_357 (O_357,N_19888,N_19756);
nor UO_358 (O_358,N_19765,N_19430);
or UO_359 (O_359,N_19834,N_19500);
nor UO_360 (O_360,N_19227,N_19410);
and UO_361 (O_361,N_19248,N_19960);
nand UO_362 (O_362,N_19322,N_19298);
nor UO_363 (O_363,N_19661,N_19591);
nand UO_364 (O_364,N_19912,N_19457);
and UO_365 (O_365,N_19480,N_19404);
xor UO_366 (O_366,N_19941,N_19862);
nor UO_367 (O_367,N_19715,N_19738);
or UO_368 (O_368,N_19620,N_19811);
xor UO_369 (O_369,N_19781,N_19395);
nand UO_370 (O_370,N_19853,N_19330);
and UO_371 (O_371,N_19770,N_19203);
nor UO_372 (O_372,N_19263,N_19296);
or UO_373 (O_373,N_19366,N_19654);
or UO_374 (O_374,N_19344,N_19845);
or UO_375 (O_375,N_19309,N_19211);
nor UO_376 (O_376,N_19758,N_19525);
or UO_377 (O_377,N_19506,N_19391);
or UO_378 (O_378,N_19572,N_19937);
or UO_379 (O_379,N_19482,N_19504);
and UO_380 (O_380,N_19512,N_19468);
nand UO_381 (O_381,N_19393,N_19567);
xor UO_382 (O_382,N_19246,N_19678);
nor UO_383 (O_383,N_19753,N_19297);
nand UO_384 (O_384,N_19903,N_19920);
nand UO_385 (O_385,N_19644,N_19215);
nand UO_386 (O_386,N_19815,N_19271);
or UO_387 (O_387,N_19913,N_19783);
xnor UO_388 (O_388,N_19222,N_19743);
nor UO_389 (O_389,N_19439,N_19857);
or UO_390 (O_390,N_19784,N_19452);
and UO_391 (O_391,N_19839,N_19677);
or UO_392 (O_392,N_19871,N_19307);
nor UO_393 (O_393,N_19671,N_19520);
nor UO_394 (O_394,N_19744,N_19711);
or UO_395 (O_395,N_19568,N_19649);
xor UO_396 (O_396,N_19801,N_19973);
xor UO_397 (O_397,N_19241,N_19501);
xor UO_398 (O_398,N_19268,N_19376);
xnor UO_399 (O_399,N_19790,N_19881);
and UO_400 (O_400,N_19286,N_19810);
nor UO_401 (O_401,N_19585,N_19345);
nor UO_402 (O_402,N_19692,N_19280);
or UO_403 (O_403,N_19315,N_19255);
nand UO_404 (O_404,N_19560,N_19667);
and UO_405 (O_405,N_19241,N_19672);
xor UO_406 (O_406,N_19376,N_19535);
or UO_407 (O_407,N_19897,N_19799);
nor UO_408 (O_408,N_19233,N_19505);
or UO_409 (O_409,N_19913,N_19969);
or UO_410 (O_410,N_19735,N_19644);
or UO_411 (O_411,N_19732,N_19770);
or UO_412 (O_412,N_19307,N_19546);
xor UO_413 (O_413,N_19280,N_19371);
and UO_414 (O_414,N_19890,N_19553);
nand UO_415 (O_415,N_19412,N_19891);
and UO_416 (O_416,N_19338,N_19760);
xor UO_417 (O_417,N_19206,N_19510);
xor UO_418 (O_418,N_19386,N_19789);
or UO_419 (O_419,N_19723,N_19385);
xor UO_420 (O_420,N_19896,N_19456);
nand UO_421 (O_421,N_19768,N_19458);
and UO_422 (O_422,N_19569,N_19634);
nor UO_423 (O_423,N_19429,N_19810);
and UO_424 (O_424,N_19766,N_19912);
nor UO_425 (O_425,N_19590,N_19204);
nor UO_426 (O_426,N_19737,N_19279);
and UO_427 (O_427,N_19620,N_19694);
and UO_428 (O_428,N_19739,N_19853);
or UO_429 (O_429,N_19404,N_19687);
xor UO_430 (O_430,N_19351,N_19618);
or UO_431 (O_431,N_19545,N_19547);
or UO_432 (O_432,N_19956,N_19216);
nor UO_433 (O_433,N_19592,N_19824);
nand UO_434 (O_434,N_19506,N_19819);
nand UO_435 (O_435,N_19970,N_19659);
nand UO_436 (O_436,N_19411,N_19601);
or UO_437 (O_437,N_19691,N_19549);
nor UO_438 (O_438,N_19903,N_19748);
and UO_439 (O_439,N_19896,N_19772);
and UO_440 (O_440,N_19329,N_19462);
xor UO_441 (O_441,N_19809,N_19623);
xor UO_442 (O_442,N_19678,N_19267);
and UO_443 (O_443,N_19420,N_19251);
or UO_444 (O_444,N_19848,N_19545);
and UO_445 (O_445,N_19524,N_19416);
or UO_446 (O_446,N_19348,N_19556);
and UO_447 (O_447,N_19645,N_19514);
and UO_448 (O_448,N_19371,N_19738);
or UO_449 (O_449,N_19302,N_19872);
nor UO_450 (O_450,N_19685,N_19797);
nor UO_451 (O_451,N_19470,N_19225);
and UO_452 (O_452,N_19867,N_19689);
nand UO_453 (O_453,N_19516,N_19218);
nand UO_454 (O_454,N_19296,N_19838);
nand UO_455 (O_455,N_19710,N_19512);
nand UO_456 (O_456,N_19259,N_19898);
nand UO_457 (O_457,N_19959,N_19438);
or UO_458 (O_458,N_19495,N_19607);
xor UO_459 (O_459,N_19221,N_19664);
and UO_460 (O_460,N_19903,N_19780);
nor UO_461 (O_461,N_19503,N_19385);
and UO_462 (O_462,N_19799,N_19780);
xnor UO_463 (O_463,N_19657,N_19610);
and UO_464 (O_464,N_19363,N_19753);
and UO_465 (O_465,N_19405,N_19308);
nand UO_466 (O_466,N_19685,N_19990);
nor UO_467 (O_467,N_19264,N_19365);
nor UO_468 (O_468,N_19219,N_19782);
or UO_469 (O_469,N_19739,N_19985);
nor UO_470 (O_470,N_19827,N_19795);
nand UO_471 (O_471,N_19483,N_19631);
and UO_472 (O_472,N_19570,N_19606);
or UO_473 (O_473,N_19325,N_19749);
xor UO_474 (O_474,N_19997,N_19772);
and UO_475 (O_475,N_19317,N_19333);
or UO_476 (O_476,N_19311,N_19941);
or UO_477 (O_477,N_19825,N_19607);
and UO_478 (O_478,N_19516,N_19778);
nor UO_479 (O_479,N_19819,N_19726);
nor UO_480 (O_480,N_19546,N_19605);
or UO_481 (O_481,N_19937,N_19202);
and UO_482 (O_482,N_19347,N_19254);
nand UO_483 (O_483,N_19687,N_19633);
nand UO_484 (O_484,N_19466,N_19618);
xor UO_485 (O_485,N_19479,N_19354);
or UO_486 (O_486,N_19632,N_19300);
nand UO_487 (O_487,N_19362,N_19696);
and UO_488 (O_488,N_19525,N_19863);
nor UO_489 (O_489,N_19440,N_19323);
xnor UO_490 (O_490,N_19982,N_19728);
nor UO_491 (O_491,N_19910,N_19885);
nor UO_492 (O_492,N_19812,N_19685);
and UO_493 (O_493,N_19514,N_19423);
nor UO_494 (O_494,N_19931,N_19634);
nor UO_495 (O_495,N_19573,N_19896);
and UO_496 (O_496,N_19973,N_19850);
or UO_497 (O_497,N_19796,N_19952);
and UO_498 (O_498,N_19664,N_19569);
xor UO_499 (O_499,N_19678,N_19321);
nand UO_500 (O_500,N_19876,N_19332);
and UO_501 (O_501,N_19265,N_19590);
or UO_502 (O_502,N_19745,N_19448);
nor UO_503 (O_503,N_19221,N_19931);
and UO_504 (O_504,N_19306,N_19908);
or UO_505 (O_505,N_19453,N_19482);
and UO_506 (O_506,N_19474,N_19362);
nand UO_507 (O_507,N_19994,N_19700);
or UO_508 (O_508,N_19420,N_19939);
nor UO_509 (O_509,N_19422,N_19424);
nor UO_510 (O_510,N_19851,N_19831);
nand UO_511 (O_511,N_19694,N_19415);
nand UO_512 (O_512,N_19637,N_19447);
xor UO_513 (O_513,N_19392,N_19282);
or UO_514 (O_514,N_19862,N_19472);
nand UO_515 (O_515,N_19479,N_19663);
nand UO_516 (O_516,N_19257,N_19765);
or UO_517 (O_517,N_19873,N_19450);
nand UO_518 (O_518,N_19229,N_19355);
nor UO_519 (O_519,N_19573,N_19677);
nand UO_520 (O_520,N_19733,N_19799);
nand UO_521 (O_521,N_19232,N_19954);
and UO_522 (O_522,N_19654,N_19402);
and UO_523 (O_523,N_19473,N_19608);
or UO_524 (O_524,N_19837,N_19699);
or UO_525 (O_525,N_19235,N_19919);
and UO_526 (O_526,N_19511,N_19715);
nor UO_527 (O_527,N_19341,N_19975);
or UO_528 (O_528,N_19852,N_19204);
xor UO_529 (O_529,N_19758,N_19400);
nand UO_530 (O_530,N_19995,N_19235);
or UO_531 (O_531,N_19793,N_19754);
or UO_532 (O_532,N_19339,N_19911);
nand UO_533 (O_533,N_19739,N_19745);
or UO_534 (O_534,N_19306,N_19975);
and UO_535 (O_535,N_19410,N_19998);
xnor UO_536 (O_536,N_19565,N_19499);
and UO_537 (O_537,N_19483,N_19841);
or UO_538 (O_538,N_19592,N_19734);
or UO_539 (O_539,N_19385,N_19786);
xor UO_540 (O_540,N_19472,N_19411);
and UO_541 (O_541,N_19322,N_19771);
or UO_542 (O_542,N_19717,N_19757);
or UO_543 (O_543,N_19504,N_19505);
and UO_544 (O_544,N_19378,N_19363);
and UO_545 (O_545,N_19290,N_19372);
xnor UO_546 (O_546,N_19644,N_19495);
or UO_547 (O_547,N_19312,N_19221);
or UO_548 (O_548,N_19417,N_19334);
and UO_549 (O_549,N_19484,N_19937);
and UO_550 (O_550,N_19828,N_19620);
nor UO_551 (O_551,N_19244,N_19234);
and UO_552 (O_552,N_19894,N_19441);
nor UO_553 (O_553,N_19267,N_19801);
or UO_554 (O_554,N_19550,N_19485);
nand UO_555 (O_555,N_19228,N_19215);
nand UO_556 (O_556,N_19479,N_19666);
xor UO_557 (O_557,N_19609,N_19520);
and UO_558 (O_558,N_19698,N_19678);
nand UO_559 (O_559,N_19708,N_19596);
and UO_560 (O_560,N_19482,N_19322);
xor UO_561 (O_561,N_19896,N_19999);
and UO_562 (O_562,N_19949,N_19206);
and UO_563 (O_563,N_19921,N_19286);
and UO_564 (O_564,N_19477,N_19384);
nand UO_565 (O_565,N_19664,N_19255);
nor UO_566 (O_566,N_19372,N_19882);
and UO_567 (O_567,N_19654,N_19637);
nor UO_568 (O_568,N_19829,N_19234);
nor UO_569 (O_569,N_19650,N_19402);
or UO_570 (O_570,N_19520,N_19705);
and UO_571 (O_571,N_19756,N_19510);
nor UO_572 (O_572,N_19824,N_19580);
xnor UO_573 (O_573,N_19682,N_19921);
nand UO_574 (O_574,N_19886,N_19601);
or UO_575 (O_575,N_19293,N_19228);
or UO_576 (O_576,N_19534,N_19763);
and UO_577 (O_577,N_19526,N_19481);
or UO_578 (O_578,N_19472,N_19516);
or UO_579 (O_579,N_19644,N_19747);
nand UO_580 (O_580,N_19984,N_19710);
or UO_581 (O_581,N_19863,N_19935);
nand UO_582 (O_582,N_19320,N_19310);
nor UO_583 (O_583,N_19534,N_19603);
nand UO_584 (O_584,N_19273,N_19349);
and UO_585 (O_585,N_19491,N_19627);
and UO_586 (O_586,N_19961,N_19369);
nand UO_587 (O_587,N_19797,N_19902);
nand UO_588 (O_588,N_19401,N_19715);
or UO_589 (O_589,N_19755,N_19959);
and UO_590 (O_590,N_19445,N_19740);
or UO_591 (O_591,N_19720,N_19983);
nor UO_592 (O_592,N_19237,N_19705);
xor UO_593 (O_593,N_19334,N_19884);
nand UO_594 (O_594,N_19813,N_19370);
nor UO_595 (O_595,N_19479,N_19674);
xnor UO_596 (O_596,N_19301,N_19705);
xnor UO_597 (O_597,N_19402,N_19533);
nor UO_598 (O_598,N_19745,N_19231);
nor UO_599 (O_599,N_19443,N_19682);
nor UO_600 (O_600,N_19509,N_19510);
and UO_601 (O_601,N_19667,N_19519);
nand UO_602 (O_602,N_19826,N_19301);
xor UO_603 (O_603,N_19250,N_19879);
nor UO_604 (O_604,N_19811,N_19838);
nor UO_605 (O_605,N_19820,N_19819);
nor UO_606 (O_606,N_19555,N_19794);
and UO_607 (O_607,N_19318,N_19882);
xor UO_608 (O_608,N_19967,N_19662);
xor UO_609 (O_609,N_19589,N_19330);
xor UO_610 (O_610,N_19609,N_19577);
or UO_611 (O_611,N_19493,N_19998);
nor UO_612 (O_612,N_19525,N_19900);
and UO_613 (O_613,N_19366,N_19811);
nand UO_614 (O_614,N_19722,N_19289);
nand UO_615 (O_615,N_19880,N_19444);
xor UO_616 (O_616,N_19759,N_19494);
nor UO_617 (O_617,N_19911,N_19483);
and UO_618 (O_618,N_19281,N_19341);
xnor UO_619 (O_619,N_19518,N_19761);
and UO_620 (O_620,N_19250,N_19429);
nor UO_621 (O_621,N_19758,N_19994);
and UO_622 (O_622,N_19463,N_19538);
nor UO_623 (O_623,N_19906,N_19277);
nor UO_624 (O_624,N_19886,N_19317);
or UO_625 (O_625,N_19883,N_19853);
and UO_626 (O_626,N_19214,N_19441);
and UO_627 (O_627,N_19728,N_19511);
and UO_628 (O_628,N_19831,N_19296);
or UO_629 (O_629,N_19300,N_19595);
or UO_630 (O_630,N_19372,N_19855);
and UO_631 (O_631,N_19582,N_19965);
nand UO_632 (O_632,N_19676,N_19479);
xor UO_633 (O_633,N_19515,N_19599);
nor UO_634 (O_634,N_19555,N_19621);
nand UO_635 (O_635,N_19322,N_19445);
nand UO_636 (O_636,N_19921,N_19242);
or UO_637 (O_637,N_19383,N_19999);
nor UO_638 (O_638,N_19595,N_19861);
nand UO_639 (O_639,N_19607,N_19856);
xor UO_640 (O_640,N_19477,N_19432);
nor UO_641 (O_641,N_19554,N_19752);
or UO_642 (O_642,N_19820,N_19417);
and UO_643 (O_643,N_19286,N_19363);
nand UO_644 (O_644,N_19434,N_19722);
and UO_645 (O_645,N_19567,N_19482);
nor UO_646 (O_646,N_19572,N_19751);
or UO_647 (O_647,N_19706,N_19430);
nand UO_648 (O_648,N_19655,N_19743);
xnor UO_649 (O_649,N_19804,N_19956);
or UO_650 (O_650,N_19757,N_19523);
nand UO_651 (O_651,N_19888,N_19330);
and UO_652 (O_652,N_19426,N_19328);
and UO_653 (O_653,N_19614,N_19965);
nand UO_654 (O_654,N_19317,N_19462);
and UO_655 (O_655,N_19894,N_19318);
nor UO_656 (O_656,N_19909,N_19809);
or UO_657 (O_657,N_19253,N_19493);
and UO_658 (O_658,N_19827,N_19934);
and UO_659 (O_659,N_19382,N_19940);
or UO_660 (O_660,N_19745,N_19542);
nand UO_661 (O_661,N_19236,N_19862);
and UO_662 (O_662,N_19771,N_19440);
and UO_663 (O_663,N_19926,N_19773);
and UO_664 (O_664,N_19319,N_19333);
and UO_665 (O_665,N_19260,N_19482);
xnor UO_666 (O_666,N_19870,N_19765);
xnor UO_667 (O_667,N_19230,N_19442);
and UO_668 (O_668,N_19399,N_19624);
nand UO_669 (O_669,N_19932,N_19369);
and UO_670 (O_670,N_19785,N_19814);
nand UO_671 (O_671,N_19628,N_19746);
or UO_672 (O_672,N_19435,N_19499);
or UO_673 (O_673,N_19978,N_19420);
or UO_674 (O_674,N_19599,N_19539);
xnor UO_675 (O_675,N_19313,N_19636);
nor UO_676 (O_676,N_19598,N_19449);
nor UO_677 (O_677,N_19983,N_19994);
nor UO_678 (O_678,N_19989,N_19790);
xor UO_679 (O_679,N_19474,N_19331);
xor UO_680 (O_680,N_19319,N_19723);
nor UO_681 (O_681,N_19286,N_19783);
or UO_682 (O_682,N_19491,N_19473);
and UO_683 (O_683,N_19283,N_19297);
or UO_684 (O_684,N_19915,N_19528);
and UO_685 (O_685,N_19423,N_19855);
nor UO_686 (O_686,N_19892,N_19330);
or UO_687 (O_687,N_19275,N_19200);
nand UO_688 (O_688,N_19363,N_19984);
nor UO_689 (O_689,N_19881,N_19413);
or UO_690 (O_690,N_19381,N_19647);
nand UO_691 (O_691,N_19269,N_19590);
nor UO_692 (O_692,N_19467,N_19865);
nand UO_693 (O_693,N_19726,N_19427);
xnor UO_694 (O_694,N_19981,N_19302);
xnor UO_695 (O_695,N_19692,N_19691);
nor UO_696 (O_696,N_19236,N_19668);
and UO_697 (O_697,N_19583,N_19466);
xnor UO_698 (O_698,N_19505,N_19242);
or UO_699 (O_699,N_19950,N_19569);
nor UO_700 (O_700,N_19608,N_19861);
xor UO_701 (O_701,N_19428,N_19334);
nor UO_702 (O_702,N_19707,N_19439);
xor UO_703 (O_703,N_19495,N_19339);
and UO_704 (O_704,N_19248,N_19959);
xor UO_705 (O_705,N_19252,N_19970);
xor UO_706 (O_706,N_19283,N_19399);
xor UO_707 (O_707,N_19911,N_19487);
nor UO_708 (O_708,N_19481,N_19798);
and UO_709 (O_709,N_19368,N_19790);
or UO_710 (O_710,N_19280,N_19402);
and UO_711 (O_711,N_19442,N_19758);
nor UO_712 (O_712,N_19786,N_19347);
nor UO_713 (O_713,N_19541,N_19813);
and UO_714 (O_714,N_19972,N_19363);
nor UO_715 (O_715,N_19973,N_19659);
xnor UO_716 (O_716,N_19859,N_19882);
nor UO_717 (O_717,N_19670,N_19652);
nor UO_718 (O_718,N_19331,N_19323);
xor UO_719 (O_719,N_19681,N_19323);
nand UO_720 (O_720,N_19518,N_19635);
or UO_721 (O_721,N_19729,N_19811);
nand UO_722 (O_722,N_19264,N_19238);
and UO_723 (O_723,N_19441,N_19430);
xnor UO_724 (O_724,N_19801,N_19695);
or UO_725 (O_725,N_19447,N_19312);
nand UO_726 (O_726,N_19203,N_19243);
xor UO_727 (O_727,N_19445,N_19667);
and UO_728 (O_728,N_19255,N_19495);
nand UO_729 (O_729,N_19503,N_19432);
nor UO_730 (O_730,N_19596,N_19394);
nand UO_731 (O_731,N_19372,N_19611);
or UO_732 (O_732,N_19544,N_19717);
nand UO_733 (O_733,N_19498,N_19698);
and UO_734 (O_734,N_19301,N_19874);
or UO_735 (O_735,N_19227,N_19748);
and UO_736 (O_736,N_19699,N_19929);
xnor UO_737 (O_737,N_19556,N_19905);
and UO_738 (O_738,N_19604,N_19973);
nand UO_739 (O_739,N_19357,N_19633);
or UO_740 (O_740,N_19401,N_19723);
or UO_741 (O_741,N_19907,N_19442);
or UO_742 (O_742,N_19591,N_19204);
nand UO_743 (O_743,N_19873,N_19574);
nand UO_744 (O_744,N_19458,N_19434);
xnor UO_745 (O_745,N_19931,N_19356);
and UO_746 (O_746,N_19349,N_19675);
nand UO_747 (O_747,N_19344,N_19643);
and UO_748 (O_748,N_19489,N_19872);
xnor UO_749 (O_749,N_19637,N_19325);
nand UO_750 (O_750,N_19938,N_19883);
xnor UO_751 (O_751,N_19651,N_19720);
nand UO_752 (O_752,N_19209,N_19891);
or UO_753 (O_753,N_19391,N_19768);
and UO_754 (O_754,N_19305,N_19481);
xnor UO_755 (O_755,N_19540,N_19942);
xor UO_756 (O_756,N_19462,N_19976);
or UO_757 (O_757,N_19366,N_19925);
xnor UO_758 (O_758,N_19830,N_19588);
nor UO_759 (O_759,N_19203,N_19789);
and UO_760 (O_760,N_19979,N_19719);
or UO_761 (O_761,N_19469,N_19442);
nand UO_762 (O_762,N_19733,N_19467);
nand UO_763 (O_763,N_19869,N_19822);
xnor UO_764 (O_764,N_19272,N_19641);
or UO_765 (O_765,N_19965,N_19545);
nand UO_766 (O_766,N_19223,N_19257);
nand UO_767 (O_767,N_19976,N_19800);
or UO_768 (O_768,N_19878,N_19649);
nand UO_769 (O_769,N_19243,N_19478);
xnor UO_770 (O_770,N_19454,N_19413);
or UO_771 (O_771,N_19361,N_19979);
and UO_772 (O_772,N_19552,N_19774);
nor UO_773 (O_773,N_19754,N_19268);
nor UO_774 (O_774,N_19461,N_19918);
or UO_775 (O_775,N_19236,N_19595);
nor UO_776 (O_776,N_19234,N_19798);
nor UO_777 (O_777,N_19211,N_19327);
nand UO_778 (O_778,N_19523,N_19678);
nand UO_779 (O_779,N_19707,N_19599);
nand UO_780 (O_780,N_19770,N_19259);
nand UO_781 (O_781,N_19823,N_19776);
xnor UO_782 (O_782,N_19945,N_19706);
nor UO_783 (O_783,N_19303,N_19915);
nor UO_784 (O_784,N_19345,N_19738);
and UO_785 (O_785,N_19368,N_19608);
nand UO_786 (O_786,N_19434,N_19767);
nor UO_787 (O_787,N_19711,N_19794);
and UO_788 (O_788,N_19278,N_19824);
and UO_789 (O_789,N_19939,N_19879);
xor UO_790 (O_790,N_19636,N_19393);
nand UO_791 (O_791,N_19470,N_19994);
nand UO_792 (O_792,N_19919,N_19361);
nor UO_793 (O_793,N_19342,N_19500);
and UO_794 (O_794,N_19917,N_19584);
or UO_795 (O_795,N_19401,N_19579);
and UO_796 (O_796,N_19902,N_19376);
and UO_797 (O_797,N_19952,N_19410);
xnor UO_798 (O_798,N_19759,N_19440);
nor UO_799 (O_799,N_19233,N_19967);
and UO_800 (O_800,N_19363,N_19433);
and UO_801 (O_801,N_19859,N_19444);
nand UO_802 (O_802,N_19730,N_19504);
nor UO_803 (O_803,N_19273,N_19481);
and UO_804 (O_804,N_19809,N_19512);
nor UO_805 (O_805,N_19581,N_19247);
nand UO_806 (O_806,N_19215,N_19661);
and UO_807 (O_807,N_19769,N_19514);
nand UO_808 (O_808,N_19398,N_19931);
and UO_809 (O_809,N_19727,N_19667);
or UO_810 (O_810,N_19800,N_19713);
xnor UO_811 (O_811,N_19508,N_19316);
xor UO_812 (O_812,N_19700,N_19249);
or UO_813 (O_813,N_19557,N_19995);
nor UO_814 (O_814,N_19593,N_19473);
and UO_815 (O_815,N_19385,N_19747);
nand UO_816 (O_816,N_19881,N_19972);
xnor UO_817 (O_817,N_19213,N_19291);
or UO_818 (O_818,N_19303,N_19939);
xnor UO_819 (O_819,N_19626,N_19684);
nor UO_820 (O_820,N_19241,N_19340);
or UO_821 (O_821,N_19767,N_19216);
and UO_822 (O_822,N_19399,N_19877);
nand UO_823 (O_823,N_19850,N_19505);
nor UO_824 (O_824,N_19653,N_19740);
xor UO_825 (O_825,N_19745,N_19271);
xor UO_826 (O_826,N_19295,N_19820);
nand UO_827 (O_827,N_19575,N_19741);
and UO_828 (O_828,N_19363,N_19953);
or UO_829 (O_829,N_19712,N_19710);
or UO_830 (O_830,N_19982,N_19797);
nor UO_831 (O_831,N_19365,N_19557);
and UO_832 (O_832,N_19311,N_19832);
nor UO_833 (O_833,N_19659,N_19872);
xor UO_834 (O_834,N_19849,N_19236);
nor UO_835 (O_835,N_19440,N_19333);
xnor UO_836 (O_836,N_19841,N_19482);
or UO_837 (O_837,N_19478,N_19323);
nand UO_838 (O_838,N_19279,N_19557);
or UO_839 (O_839,N_19482,N_19264);
xor UO_840 (O_840,N_19716,N_19991);
nand UO_841 (O_841,N_19321,N_19692);
xor UO_842 (O_842,N_19970,N_19528);
nand UO_843 (O_843,N_19961,N_19215);
and UO_844 (O_844,N_19673,N_19633);
and UO_845 (O_845,N_19400,N_19591);
nor UO_846 (O_846,N_19644,N_19582);
nand UO_847 (O_847,N_19957,N_19207);
or UO_848 (O_848,N_19455,N_19438);
nor UO_849 (O_849,N_19278,N_19405);
or UO_850 (O_850,N_19203,N_19468);
and UO_851 (O_851,N_19595,N_19560);
xor UO_852 (O_852,N_19661,N_19603);
nand UO_853 (O_853,N_19980,N_19673);
xnor UO_854 (O_854,N_19373,N_19368);
nor UO_855 (O_855,N_19268,N_19252);
nor UO_856 (O_856,N_19584,N_19496);
and UO_857 (O_857,N_19449,N_19357);
nand UO_858 (O_858,N_19335,N_19984);
nor UO_859 (O_859,N_19526,N_19216);
or UO_860 (O_860,N_19858,N_19588);
or UO_861 (O_861,N_19862,N_19392);
xor UO_862 (O_862,N_19892,N_19967);
or UO_863 (O_863,N_19878,N_19286);
xnor UO_864 (O_864,N_19495,N_19920);
or UO_865 (O_865,N_19474,N_19294);
and UO_866 (O_866,N_19886,N_19925);
nor UO_867 (O_867,N_19226,N_19432);
nor UO_868 (O_868,N_19295,N_19663);
and UO_869 (O_869,N_19966,N_19357);
and UO_870 (O_870,N_19832,N_19403);
and UO_871 (O_871,N_19608,N_19691);
nand UO_872 (O_872,N_19354,N_19496);
nand UO_873 (O_873,N_19418,N_19953);
and UO_874 (O_874,N_19561,N_19698);
nand UO_875 (O_875,N_19529,N_19492);
and UO_876 (O_876,N_19895,N_19851);
and UO_877 (O_877,N_19702,N_19609);
nor UO_878 (O_878,N_19537,N_19772);
nand UO_879 (O_879,N_19819,N_19790);
nand UO_880 (O_880,N_19216,N_19437);
or UO_881 (O_881,N_19719,N_19531);
nand UO_882 (O_882,N_19917,N_19240);
xnor UO_883 (O_883,N_19531,N_19500);
nand UO_884 (O_884,N_19411,N_19416);
nor UO_885 (O_885,N_19644,N_19660);
nand UO_886 (O_886,N_19702,N_19929);
nand UO_887 (O_887,N_19532,N_19551);
or UO_888 (O_888,N_19825,N_19880);
nor UO_889 (O_889,N_19436,N_19940);
and UO_890 (O_890,N_19679,N_19518);
and UO_891 (O_891,N_19844,N_19617);
or UO_892 (O_892,N_19297,N_19524);
nand UO_893 (O_893,N_19623,N_19902);
xnor UO_894 (O_894,N_19810,N_19997);
and UO_895 (O_895,N_19920,N_19215);
or UO_896 (O_896,N_19328,N_19223);
nor UO_897 (O_897,N_19280,N_19923);
nand UO_898 (O_898,N_19554,N_19805);
and UO_899 (O_899,N_19708,N_19360);
and UO_900 (O_900,N_19217,N_19854);
and UO_901 (O_901,N_19279,N_19238);
and UO_902 (O_902,N_19390,N_19582);
nor UO_903 (O_903,N_19894,N_19505);
xor UO_904 (O_904,N_19643,N_19717);
and UO_905 (O_905,N_19872,N_19263);
nand UO_906 (O_906,N_19845,N_19612);
xor UO_907 (O_907,N_19289,N_19526);
xor UO_908 (O_908,N_19371,N_19878);
and UO_909 (O_909,N_19515,N_19796);
nor UO_910 (O_910,N_19313,N_19267);
or UO_911 (O_911,N_19425,N_19306);
or UO_912 (O_912,N_19545,N_19550);
xor UO_913 (O_913,N_19207,N_19824);
nand UO_914 (O_914,N_19626,N_19938);
nor UO_915 (O_915,N_19511,N_19342);
nand UO_916 (O_916,N_19937,N_19712);
xor UO_917 (O_917,N_19880,N_19703);
or UO_918 (O_918,N_19211,N_19563);
or UO_919 (O_919,N_19226,N_19621);
xor UO_920 (O_920,N_19844,N_19808);
nor UO_921 (O_921,N_19342,N_19374);
or UO_922 (O_922,N_19438,N_19964);
nor UO_923 (O_923,N_19741,N_19787);
or UO_924 (O_924,N_19998,N_19686);
or UO_925 (O_925,N_19758,N_19391);
nand UO_926 (O_926,N_19817,N_19487);
xor UO_927 (O_927,N_19330,N_19555);
xnor UO_928 (O_928,N_19387,N_19485);
xnor UO_929 (O_929,N_19286,N_19611);
nor UO_930 (O_930,N_19742,N_19465);
and UO_931 (O_931,N_19760,N_19443);
or UO_932 (O_932,N_19595,N_19782);
xnor UO_933 (O_933,N_19261,N_19568);
xnor UO_934 (O_934,N_19441,N_19428);
nand UO_935 (O_935,N_19595,N_19593);
or UO_936 (O_936,N_19265,N_19363);
or UO_937 (O_937,N_19521,N_19584);
nand UO_938 (O_938,N_19977,N_19936);
nand UO_939 (O_939,N_19426,N_19757);
and UO_940 (O_940,N_19657,N_19276);
nand UO_941 (O_941,N_19590,N_19625);
nor UO_942 (O_942,N_19537,N_19492);
nand UO_943 (O_943,N_19605,N_19734);
xnor UO_944 (O_944,N_19383,N_19543);
or UO_945 (O_945,N_19258,N_19791);
or UO_946 (O_946,N_19728,N_19273);
nand UO_947 (O_947,N_19462,N_19326);
xnor UO_948 (O_948,N_19938,N_19482);
xor UO_949 (O_949,N_19930,N_19428);
or UO_950 (O_950,N_19723,N_19972);
or UO_951 (O_951,N_19662,N_19875);
nand UO_952 (O_952,N_19528,N_19894);
and UO_953 (O_953,N_19317,N_19961);
xor UO_954 (O_954,N_19282,N_19878);
or UO_955 (O_955,N_19520,N_19222);
nor UO_956 (O_956,N_19391,N_19863);
nand UO_957 (O_957,N_19530,N_19216);
xnor UO_958 (O_958,N_19280,N_19200);
or UO_959 (O_959,N_19844,N_19839);
and UO_960 (O_960,N_19964,N_19900);
nor UO_961 (O_961,N_19203,N_19751);
nand UO_962 (O_962,N_19704,N_19630);
nor UO_963 (O_963,N_19799,N_19857);
xor UO_964 (O_964,N_19622,N_19726);
and UO_965 (O_965,N_19827,N_19779);
or UO_966 (O_966,N_19314,N_19402);
and UO_967 (O_967,N_19803,N_19719);
nand UO_968 (O_968,N_19270,N_19668);
xor UO_969 (O_969,N_19672,N_19475);
and UO_970 (O_970,N_19285,N_19827);
xor UO_971 (O_971,N_19915,N_19859);
xor UO_972 (O_972,N_19988,N_19599);
xnor UO_973 (O_973,N_19558,N_19314);
xnor UO_974 (O_974,N_19350,N_19964);
and UO_975 (O_975,N_19282,N_19761);
and UO_976 (O_976,N_19659,N_19694);
or UO_977 (O_977,N_19911,N_19729);
nor UO_978 (O_978,N_19322,N_19282);
nand UO_979 (O_979,N_19392,N_19278);
xor UO_980 (O_980,N_19716,N_19338);
or UO_981 (O_981,N_19327,N_19548);
or UO_982 (O_982,N_19448,N_19351);
nand UO_983 (O_983,N_19855,N_19633);
nand UO_984 (O_984,N_19684,N_19739);
or UO_985 (O_985,N_19618,N_19407);
or UO_986 (O_986,N_19552,N_19424);
xor UO_987 (O_987,N_19666,N_19766);
nand UO_988 (O_988,N_19437,N_19818);
nor UO_989 (O_989,N_19228,N_19420);
nor UO_990 (O_990,N_19388,N_19282);
nand UO_991 (O_991,N_19335,N_19439);
xnor UO_992 (O_992,N_19926,N_19651);
or UO_993 (O_993,N_19854,N_19698);
xor UO_994 (O_994,N_19948,N_19686);
and UO_995 (O_995,N_19974,N_19238);
xnor UO_996 (O_996,N_19227,N_19511);
xor UO_997 (O_997,N_19795,N_19907);
and UO_998 (O_998,N_19575,N_19552);
nand UO_999 (O_999,N_19225,N_19907);
nand UO_1000 (O_1000,N_19790,N_19844);
xor UO_1001 (O_1001,N_19299,N_19291);
xnor UO_1002 (O_1002,N_19962,N_19640);
and UO_1003 (O_1003,N_19638,N_19267);
and UO_1004 (O_1004,N_19464,N_19208);
nor UO_1005 (O_1005,N_19547,N_19759);
nor UO_1006 (O_1006,N_19444,N_19634);
xnor UO_1007 (O_1007,N_19693,N_19893);
nand UO_1008 (O_1008,N_19287,N_19674);
nand UO_1009 (O_1009,N_19724,N_19398);
and UO_1010 (O_1010,N_19757,N_19705);
nor UO_1011 (O_1011,N_19905,N_19335);
nor UO_1012 (O_1012,N_19356,N_19638);
or UO_1013 (O_1013,N_19776,N_19276);
and UO_1014 (O_1014,N_19996,N_19259);
and UO_1015 (O_1015,N_19975,N_19478);
nor UO_1016 (O_1016,N_19271,N_19429);
and UO_1017 (O_1017,N_19594,N_19658);
nand UO_1018 (O_1018,N_19500,N_19363);
and UO_1019 (O_1019,N_19811,N_19732);
or UO_1020 (O_1020,N_19416,N_19329);
nand UO_1021 (O_1021,N_19332,N_19319);
and UO_1022 (O_1022,N_19657,N_19583);
or UO_1023 (O_1023,N_19598,N_19909);
or UO_1024 (O_1024,N_19327,N_19478);
nor UO_1025 (O_1025,N_19976,N_19989);
and UO_1026 (O_1026,N_19513,N_19933);
nand UO_1027 (O_1027,N_19599,N_19752);
nand UO_1028 (O_1028,N_19334,N_19313);
xor UO_1029 (O_1029,N_19326,N_19794);
and UO_1030 (O_1030,N_19937,N_19298);
xnor UO_1031 (O_1031,N_19229,N_19774);
nand UO_1032 (O_1032,N_19923,N_19297);
or UO_1033 (O_1033,N_19793,N_19427);
nand UO_1034 (O_1034,N_19576,N_19376);
nand UO_1035 (O_1035,N_19925,N_19365);
or UO_1036 (O_1036,N_19715,N_19301);
xor UO_1037 (O_1037,N_19818,N_19334);
xor UO_1038 (O_1038,N_19854,N_19892);
nor UO_1039 (O_1039,N_19607,N_19947);
xnor UO_1040 (O_1040,N_19658,N_19744);
or UO_1041 (O_1041,N_19229,N_19446);
or UO_1042 (O_1042,N_19523,N_19935);
nor UO_1043 (O_1043,N_19416,N_19239);
nor UO_1044 (O_1044,N_19266,N_19944);
nand UO_1045 (O_1045,N_19990,N_19325);
and UO_1046 (O_1046,N_19410,N_19894);
and UO_1047 (O_1047,N_19858,N_19266);
or UO_1048 (O_1048,N_19936,N_19236);
nor UO_1049 (O_1049,N_19954,N_19588);
xnor UO_1050 (O_1050,N_19620,N_19497);
xor UO_1051 (O_1051,N_19897,N_19809);
and UO_1052 (O_1052,N_19392,N_19891);
nor UO_1053 (O_1053,N_19224,N_19511);
nor UO_1054 (O_1054,N_19475,N_19647);
xnor UO_1055 (O_1055,N_19229,N_19512);
nand UO_1056 (O_1056,N_19246,N_19688);
nor UO_1057 (O_1057,N_19536,N_19849);
xor UO_1058 (O_1058,N_19688,N_19464);
nor UO_1059 (O_1059,N_19270,N_19476);
and UO_1060 (O_1060,N_19618,N_19867);
xor UO_1061 (O_1061,N_19726,N_19559);
xor UO_1062 (O_1062,N_19792,N_19328);
nor UO_1063 (O_1063,N_19686,N_19738);
or UO_1064 (O_1064,N_19434,N_19883);
nor UO_1065 (O_1065,N_19263,N_19370);
or UO_1066 (O_1066,N_19338,N_19423);
nand UO_1067 (O_1067,N_19282,N_19466);
nand UO_1068 (O_1068,N_19294,N_19348);
nand UO_1069 (O_1069,N_19677,N_19384);
and UO_1070 (O_1070,N_19769,N_19466);
and UO_1071 (O_1071,N_19504,N_19404);
nand UO_1072 (O_1072,N_19614,N_19574);
or UO_1073 (O_1073,N_19996,N_19635);
nor UO_1074 (O_1074,N_19574,N_19830);
nor UO_1075 (O_1075,N_19912,N_19211);
and UO_1076 (O_1076,N_19687,N_19966);
and UO_1077 (O_1077,N_19522,N_19691);
nand UO_1078 (O_1078,N_19795,N_19538);
or UO_1079 (O_1079,N_19348,N_19876);
xnor UO_1080 (O_1080,N_19606,N_19947);
nand UO_1081 (O_1081,N_19353,N_19242);
xor UO_1082 (O_1082,N_19358,N_19637);
nor UO_1083 (O_1083,N_19457,N_19960);
or UO_1084 (O_1084,N_19451,N_19292);
nor UO_1085 (O_1085,N_19713,N_19731);
nand UO_1086 (O_1086,N_19365,N_19895);
nor UO_1087 (O_1087,N_19758,N_19792);
and UO_1088 (O_1088,N_19860,N_19970);
and UO_1089 (O_1089,N_19973,N_19829);
xnor UO_1090 (O_1090,N_19817,N_19792);
nor UO_1091 (O_1091,N_19803,N_19552);
nand UO_1092 (O_1092,N_19443,N_19806);
or UO_1093 (O_1093,N_19970,N_19446);
xnor UO_1094 (O_1094,N_19280,N_19572);
xor UO_1095 (O_1095,N_19569,N_19815);
or UO_1096 (O_1096,N_19630,N_19694);
xor UO_1097 (O_1097,N_19715,N_19394);
or UO_1098 (O_1098,N_19674,N_19971);
nand UO_1099 (O_1099,N_19559,N_19992);
and UO_1100 (O_1100,N_19801,N_19821);
xnor UO_1101 (O_1101,N_19618,N_19611);
and UO_1102 (O_1102,N_19542,N_19736);
nand UO_1103 (O_1103,N_19689,N_19593);
and UO_1104 (O_1104,N_19503,N_19838);
xor UO_1105 (O_1105,N_19361,N_19266);
nor UO_1106 (O_1106,N_19491,N_19740);
and UO_1107 (O_1107,N_19622,N_19716);
nand UO_1108 (O_1108,N_19428,N_19611);
xnor UO_1109 (O_1109,N_19883,N_19289);
xor UO_1110 (O_1110,N_19393,N_19955);
or UO_1111 (O_1111,N_19917,N_19248);
nand UO_1112 (O_1112,N_19768,N_19961);
or UO_1113 (O_1113,N_19377,N_19284);
or UO_1114 (O_1114,N_19686,N_19464);
or UO_1115 (O_1115,N_19806,N_19389);
and UO_1116 (O_1116,N_19847,N_19782);
nand UO_1117 (O_1117,N_19742,N_19627);
and UO_1118 (O_1118,N_19535,N_19825);
nor UO_1119 (O_1119,N_19773,N_19893);
nand UO_1120 (O_1120,N_19750,N_19760);
xnor UO_1121 (O_1121,N_19799,N_19480);
or UO_1122 (O_1122,N_19743,N_19366);
nor UO_1123 (O_1123,N_19818,N_19745);
or UO_1124 (O_1124,N_19378,N_19260);
nand UO_1125 (O_1125,N_19455,N_19327);
and UO_1126 (O_1126,N_19984,N_19933);
or UO_1127 (O_1127,N_19414,N_19314);
and UO_1128 (O_1128,N_19439,N_19964);
and UO_1129 (O_1129,N_19263,N_19617);
nor UO_1130 (O_1130,N_19634,N_19219);
nor UO_1131 (O_1131,N_19292,N_19628);
xor UO_1132 (O_1132,N_19754,N_19777);
nand UO_1133 (O_1133,N_19277,N_19537);
nand UO_1134 (O_1134,N_19505,N_19383);
nor UO_1135 (O_1135,N_19917,N_19901);
nor UO_1136 (O_1136,N_19792,N_19265);
xnor UO_1137 (O_1137,N_19431,N_19535);
or UO_1138 (O_1138,N_19984,N_19441);
or UO_1139 (O_1139,N_19621,N_19347);
xor UO_1140 (O_1140,N_19603,N_19346);
xnor UO_1141 (O_1141,N_19359,N_19667);
nor UO_1142 (O_1142,N_19261,N_19452);
and UO_1143 (O_1143,N_19510,N_19251);
nand UO_1144 (O_1144,N_19237,N_19331);
xor UO_1145 (O_1145,N_19635,N_19610);
nor UO_1146 (O_1146,N_19920,N_19751);
nor UO_1147 (O_1147,N_19437,N_19529);
and UO_1148 (O_1148,N_19699,N_19405);
and UO_1149 (O_1149,N_19684,N_19258);
nand UO_1150 (O_1150,N_19735,N_19789);
or UO_1151 (O_1151,N_19738,N_19963);
and UO_1152 (O_1152,N_19665,N_19457);
nor UO_1153 (O_1153,N_19244,N_19465);
xnor UO_1154 (O_1154,N_19841,N_19423);
xor UO_1155 (O_1155,N_19734,N_19601);
nor UO_1156 (O_1156,N_19376,N_19989);
or UO_1157 (O_1157,N_19562,N_19462);
nor UO_1158 (O_1158,N_19480,N_19832);
and UO_1159 (O_1159,N_19675,N_19810);
nor UO_1160 (O_1160,N_19409,N_19483);
and UO_1161 (O_1161,N_19212,N_19935);
and UO_1162 (O_1162,N_19752,N_19809);
and UO_1163 (O_1163,N_19732,N_19374);
or UO_1164 (O_1164,N_19903,N_19586);
nor UO_1165 (O_1165,N_19666,N_19312);
nand UO_1166 (O_1166,N_19539,N_19584);
or UO_1167 (O_1167,N_19983,N_19387);
xnor UO_1168 (O_1168,N_19327,N_19541);
or UO_1169 (O_1169,N_19712,N_19225);
and UO_1170 (O_1170,N_19708,N_19492);
nand UO_1171 (O_1171,N_19591,N_19495);
nor UO_1172 (O_1172,N_19261,N_19966);
nor UO_1173 (O_1173,N_19471,N_19528);
and UO_1174 (O_1174,N_19341,N_19773);
xor UO_1175 (O_1175,N_19358,N_19472);
or UO_1176 (O_1176,N_19650,N_19964);
nor UO_1177 (O_1177,N_19963,N_19819);
nor UO_1178 (O_1178,N_19382,N_19700);
nand UO_1179 (O_1179,N_19433,N_19838);
xor UO_1180 (O_1180,N_19671,N_19843);
nor UO_1181 (O_1181,N_19774,N_19590);
or UO_1182 (O_1182,N_19964,N_19494);
nand UO_1183 (O_1183,N_19959,N_19636);
or UO_1184 (O_1184,N_19614,N_19856);
nand UO_1185 (O_1185,N_19260,N_19445);
or UO_1186 (O_1186,N_19804,N_19228);
nand UO_1187 (O_1187,N_19538,N_19898);
nor UO_1188 (O_1188,N_19467,N_19298);
or UO_1189 (O_1189,N_19803,N_19766);
nor UO_1190 (O_1190,N_19783,N_19538);
and UO_1191 (O_1191,N_19281,N_19860);
nor UO_1192 (O_1192,N_19244,N_19968);
nand UO_1193 (O_1193,N_19291,N_19870);
or UO_1194 (O_1194,N_19919,N_19949);
and UO_1195 (O_1195,N_19588,N_19217);
or UO_1196 (O_1196,N_19805,N_19702);
or UO_1197 (O_1197,N_19765,N_19307);
xnor UO_1198 (O_1198,N_19745,N_19440);
and UO_1199 (O_1199,N_19632,N_19315);
xnor UO_1200 (O_1200,N_19280,N_19315);
and UO_1201 (O_1201,N_19708,N_19367);
xnor UO_1202 (O_1202,N_19427,N_19443);
and UO_1203 (O_1203,N_19296,N_19627);
nand UO_1204 (O_1204,N_19928,N_19276);
xor UO_1205 (O_1205,N_19880,N_19683);
xnor UO_1206 (O_1206,N_19750,N_19300);
xnor UO_1207 (O_1207,N_19388,N_19687);
nand UO_1208 (O_1208,N_19629,N_19616);
or UO_1209 (O_1209,N_19541,N_19227);
xnor UO_1210 (O_1210,N_19939,N_19812);
xnor UO_1211 (O_1211,N_19721,N_19320);
nand UO_1212 (O_1212,N_19550,N_19476);
nor UO_1213 (O_1213,N_19565,N_19702);
nand UO_1214 (O_1214,N_19800,N_19335);
xor UO_1215 (O_1215,N_19745,N_19608);
nor UO_1216 (O_1216,N_19363,N_19310);
nor UO_1217 (O_1217,N_19589,N_19591);
and UO_1218 (O_1218,N_19505,N_19778);
nand UO_1219 (O_1219,N_19886,N_19605);
xor UO_1220 (O_1220,N_19817,N_19335);
and UO_1221 (O_1221,N_19824,N_19397);
nor UO_1222 (O_1222,N_19678,N_19562);
nand UO_1223 (O_1223,N_19804,N_19952);
nor UO_1224 (O_1224,N_19624,N_19696);
nor UO_1225 (O_1225,N_19318,N_19734);
and UO_1226 (O_1226,N_19484,N_19952);
nand UO_1227 (O_1227,N_19343,N_19943);
nor UO_1228 (O_1228,N_19282,N_19877);
nor UO_1229 (O_1229,N_19449,N_19320);
or UO_1230 (O_1230,N_19379,N_19615);
nand UO_1231 (O_1231,N_19697,N_19550);
xnor UO_1232 (O_1232,N_19212,N_19333);
and UO_1233 (O_1233,N_19212,N_19848);
and UO_1234 (O_1234,N_19962,N_19234);
or UO_1235 (O_1235,N_19298,N_19821);
or UO_1236 (O_1236,N_19639,N_19698);
xor UO_1237 (O_1237,N_19877,N_19885);
nand UO_1238 (O_1238,N_19662,N_19677);
and UO_1239 (O_1239,N_19559,N_19708);
nand UO_1240 (O_1240,N_19982,N_19382);
nor UO_1241 (O_1241,N_19541,N_19912);
and UO_1242 (O_1242,N_19540,N_19557);
and UO_1243 (O_1243,N_19961,N_19830);
nor UO_1244 (O_1244,N_19240,N_19677);
and UO_1245 (O_1245,N_19452,N_19695);
and UO_1246 (O_1246,N_19399,N_19833);
or UO_1247 (O_1247,N_19904,N_19200);
nand UO_1248 (O_1248,N_19556,N_19530);
and UO_1249 (O_1249,N_19793,N_19773);
and UO_1250 (O_1250,N_19224,N_19263);
xnor UO_1251 (O_1251,N_19403,N_19564);
xor UO_1252 (O_1252,N_19273,N_19847);
or UO_1253 (O_1253,N_19989,N_19917);
xor UO_1254 (O_1254,N_19809,N_19443);
nor UO_1255 (O_1255,N_19332,N_19291);
nand UO_1256 (O_1256,N_19592,N_19473);
and UO_1257 (O_1257,N_19643,N_19919);
xnor UO_1258 (O_1258,N_19233,N_19469);
and UO_1259 (O_1259,N_19612,N_19607);
xnor UO_1260 (O_1260,N_19704,N_19725);
nor UO_1261 (O_1261,N_19394,N_19213);
xnor UO_1262 (O_1262,N_19214,N_19408);
or UO_1263 (O_1263,N_19783,N_19587);
xnor UO_1264 (O_1264,N_19276,N_19974);
nor UO_1265 (O_1265,N_19350,N_19801);
and UO_1266 (O_1266,N_19699,N_19390);
nor UO_1267 (O_1267,N_19880,N_19565);
nor UO_1268 (O_1268,N_19489,N_19927);
nor UO_1269 (O_1269,N_19599,N_19535);
or UO_1270 (O_1270,N_19758,N_19553);
nand UO_1271 (O_1271,N_19329,N_19972);
nor UO_1272 (O_1272,N_19807,N_19975);
nand UO_1273 (O_1273,N_19743,N_19312);
and UO_1274 (O_1274,N_19768,N_19278);
nand UO_1275 (O_1275,N_19423,N_19366);
xnor UO_1276 (O_1276,N_19472,N_19914);
nand UO_1277 (O_1277,N_19299,N_19499);
xnor UO_1278 (O_1278,N_19540,N_19325);
or UO_1279 (O_1279,N_19499,N_19634);
nand UO_1280 (O_1280,N_19841,N_19403);
and UO_1281 (O_1281,N_19455,N_19207);
and UO_1282 (O_1282,N_19831,N_19812);
nand UO_1283 (O_1283,N_19253,N_19318);
or UO_1284 (O_1284,N_19624,N_19294);
and UO_1285 (O_1285,N_19728,N_19694);
nand UO_1286 (O_1286,N_19527,N_19714);
nor UO_1287 (O_1287,N_19307,N_19264);
and UO_1288 (O_1288,N_19762,N_19724);
and UO_1289 (O_1289,N_19982,N_19680);
nand UO_1290 (O_1290,N_19763,N_19368);
nor UO_1291 (O_1291,N_19894,N_19331);
xor UO_1292 (O_1292,N_19375,N_19316);
and UO_1293 (O_1293,N_19395,N_19213);
nand UO_1294 (O_1294,N_19771,N_19519);
and UO_1295 (O_1295,N_19718,N_19412);
or UO_1296 (O_1296,N_19766,N_19997);
or UO_1297 (O_1297,N_19274,N_19546);
xnor UO_1298 (O_1298,N_19474,N_19805);
or UO_1299 (O_1299,N_19425,N_19416);
nor UO_1300 (O_1300,N_19663,N_19475);
and UO_1301 (O_1301,N_19286,N_19733);
xor UO_1302 (O_1302,N_19282,N_19319);
nand UO_1303 (O_1303,N_19405,N_19298);
nor UO_1304 (O_1304,N_19914,N_19418);
or UO_1305 (O_1305,N_19215,N_19574);
or UO_1306 (O_1306,N_19654,N_19633);
or UO_1307 (O_1307,N_19378,N_19822);
or UO_1308 (O_1308,N_19410,N_19428);
nand UO_1309 (O_1309,N_19894,N_19958);
nand UO_1310 (O_1310,N_19861,N_19822);
xnor UO_1311 (O_1311,N_19851,N_19217);
xor UO_1312 (O_1312,N_19553,N_19240);
xor UO_1313 (O_1313,N_19303,N_19311);
or UO_1314 (O_1314,N_19903,N_19312);
and UO_1315 (O_1315,N_19904,N_19787);
or UO_1316 (O_1316,N_19421,N_19637);
xnor UO_1317 (O_1317,N_19367,N_19228);
nand UO_1318 (O_1318,N_19924,N_19868);
xor UO_1319 (O_1319,N_19655,N_19919);
and UO_1320 (O_1320,N_19863,N_19452);
and UO_1321 (O_1321,N_19243,N_19936);
and UO_1322 (O_1322,N_19890,N_19676);
nor UO_1323 (O_1323,N_19403,N_19571);
and UO_1324 (O_1324,N_19791,N_19879);
nand UO_1325 (O_1325,N_19207,N_19670);
nor UO_1326 (O_1326,N_19302,N_19972);
nor UO_1327 (O_1327,N_19309,N_19236);
or UO_1328 (O_1328,N_19479,N_19317);
and UO_1329 (O_1329,N_19460,N_19369);
nand UO_1330 (O_1330,N_19604,N_19256);
and UO_1331 (O_1331,N_19305,N_19745);
and UO_1332 (O_1332,N_19573,N_19411);
nor UO_1333 (O_1333,N_19530,N_19851);
and UO_1334 (O_1334,N_19278,N_19348);
and UO_1335 (O_1335,N_19711,N_19753);
xor UO_1336 (O_1336,N_19857,N_19626);
xnor UO_1337 (O_1337,N_19476,N_19289);
or UO_1338 (O_1338,N_19241,N_19420);
xor UO_1339 (O_1339,N_19420,N_19400);
xor UO_1340 (O_1340,N_19516,N_19685);
or UO_1341 (O_1341,N_19710,N_19908);
nand UO_1342 (O_1342,N_19373,N_19869);
or UO_1343 (O_1343,N_19612,N_19715);
or UO_1344 (O_1344,N_19266,N_19947);
nand UO_1345 (O_1345,N_19726,N_19571);
and UO_1346 (O_1346,N_19291,N_19285);
or UO_1347 (O_1347,N_19936,N_19945);
and UO_1348 (O_1348,N_19869,N_19481);
or UO_1349 (O_1349,N_19300,N_19614);
or UO_1350 (O_1350,N_19301,N_19210);
xor UO_1351 (O_1351,N_19560,N_19377);
or UO_1352 (O_1352,N_19491,N_19263);
and UO_1353 (O_1353,N_19205,N_19903);
nand UO_1354 (O_1354,N_19735,N_19505);
xnor UO_1355 (O_1355,N_19407,N_19354);
nand UO_1356 (O_1356,N_19784,N_19662);
and UO_1357 (O_1357,N_19542,N_19732);
and UO_1358 (O_1358,N_19701,N_19953);
xor UO_1359 (O_1359,N_19871,N_19922);
nand UO_1360 (O_1360,N_19444,N_19388);
nor UO_1361 (O_1361,N_19201,N_19252);
or UO_1362 (O_1362,N_19568,N_19601);
nand UO_1363 (O_1363,N_19642,N_19452);
and UO_1364 (O_1364,N_19856,N_19340);
nand UO_1365 (O_1365,N_19827,N_19437);
nor UO_1366 (O_1366,N_19507,N_19304);
nand UO_1367 (O_1367,N_19716,N_19765);
xor UO_1368 (O_1368,N_19777,N_19487);
xor UO_1369 (O_1369,N_19879,N_19403);
nor UO_1370 (O_1370,N_19597,N_19893);
xnor UO_1371 (O_1371,N_19754,N_19670);
nand UO_1372 (O_1372,N_19615,N_19241);
or UO_1373 (O_1373,N_19767,N_19502);
nor UO_1374 (O_1374,N_19532,N_19263);
or UO_1375 (O_1375,N_19716,N_19704);
nand UO_1376 (O_1376,N_19549,N_19293);
xnor UO_1377 (O_1377,N_19412,N_19586);
and UO_1378 (O_1378,N_19626,N_19952);
nand UO_1379 (O_1379,N_19404,N_19991);
nand UO_1380 (O_1380,N_19351,N_19239);
nand UO_1381 (O_1381,N_19377,N_19675);
xor UO_1382 (O_1382,N_19821,N_19320);
xnor UO_1383 (O_1383,N_19987,N_19305);
xnor UO_1384 (O_1384,N_19580,N_19273);
or UO_1385 (O_1385,N_19863,N_19666);
nor UO_1386 (O_1386,N_19848,N_19776);
and UO_1387 (O_1387,N_19412,N_19969);
nand UO_1388 (O_1388,N_19558,N_19628);
nand UO_1389 (O_1389,N_19624,N_19219);
or UO_1390 (O_1390,N_19436,N_19437);
nand UO_1391 (O_1391,N_19722,N_19475);
and UO_1392 (O_1392,N_19723,N_19837);
or UO_1393 (O_1393,N_19215,N_19962);
xor UO_1394 (O_1394,N_19702,N_19600);
and UO_1395 (O_1395,N_19413,N_19537);
nand UO_1396 (O_1396,N_19360,N_19882);
nor UO_1397 (O_1397,N_19680,N_19799);
nand UO_1398 (O_1398,N_19218,N_19738);
xnor UO_1399 (O_1399,N_19978,N_19570);
or UO_1400 (O_1400,N_19673,N_19599);
and UO_1401 (O_1401,N_19598,N_19409);
or UO_1402 (O_1402,N_19399,N_19264);
and UO_1403 (O_1403,N_19315,N_19760);
or UO_1404 (O_1404,N_19273,N_19659);
nor UO_1405 (O_1405,N_19412,N_19514);
or UO_1406 (O_1406,N_19785,N_19847);
nand UO_1407 (O_1407,N_19867,N_19667);
or UO_1408 (O_1408,N_19348,N_19856);
and UO_1409 (O_1409,N_19711,N_19285);
nand UO_1410 (O_1410,N_19220,N_19464);
xor UO_1411 (O_1411,N_19407,N_19619);
or UO_1412 (O_1412,N_19732,N_19755);
or UO_1413 (O_1413,N_19652,N_19454);
xor UO_1414 (O_1414,N_19873,N_19631);
xnor UO_1415 (O_1415,N_19303,N_19556);
nor UO_1416 (O_1416,N_19249,N_19680);
or UO_1417 (O_1417,N_19290,N_19840);
and UO_1418 (O_1418,N_19248,N_19441);
or UO_1419 (O_1419,N_19640,N_19960);
and UO_1420 (O_1420,N_19361,N_19378);
nand UO_1421 (O_1421,N_19209,N_19234);
nand UO_1422 (O_1422,N_19470,N_19696);
nor UO_1423 (O_1423,N_19575,N_19707);
or UO_1424 (O_1424,N_19635,N_19962);
and UO_1425 (O_1425,N_19801,N_19502);
nor UO_1426 (O_1426,N_19554,N_19367);
nand UO_1427 (O_1427,N_19472,N_19495);
and UO_1428 (O_1428,N_19357,N_19566);
nor UO_1429 (O_1429,N_19734,N_19342);
xor UO_1430 (O_1430,N_19836,N_19521);
nand UO_1431 (O_1431,N_19547,N_19920);
or UO_1432 (O_1432,N_19549,N_19361);
and UO_1433 (O_1433,N_19309,N_19484);
nand UO_1434 (O_1434,N_19725,N_19504);
or UO_1435 (O_1435,N_19924,N_19509);
and UO_1436 (O_1436,N_19776,N_19245);
and UO_1437 (O_1437,N_19408,N_19993);
nand UO_1438 (O_1438,N_19627,N_19671);
nor UO_1439 (O_1439,N_19788,N_19422);
nor UO_1440 (O_1440,N_19816,N_19278);
nand UO_1441 (O_1441,N_19691,N_19277);
nand UO_1442 (O_1442,N_19748,N_19494);
and UO_1443 (O_1443,N_19262,N_19731);
xor UO_1444 (O_1444,N_19816,N_19651);
nor UO_1445 (O_1445,N_19252,N_19334);
xor UO_1446 (O_1446,N_19791,N_19510);
nor UO_1447 (O_1447,N_19539,N_19519);
nor UO_1448 (O_1448,N_19686,N_19592);
nand UO_1449 (O_1449,N_19938,N_19301);
xor UO_1450 (O_1450,N_19917,N_19200);
xnor UO_1451 (O_1451,N_19814,N_19830);
and UO_1452 (O_1452,N_19202,N_19526);
nand UO_1453 (O_1453,N_19417,N_19231);
nand UO_1454 (O_1454,N_19658,N_19268);
xor UO_1455 (O_1455,N_19559,N_19464);
nor UO_1456 (O_1456,N_19804,N_19794);
nor UO_1457 (O_1457,N_19279,N_19928);
xnor UO_1458 (O_1458,N_19448,N_19240);
nand UO_1459 (O_1459,N_19494,N_19446);
nor UO_1460 (O_1460,N_19725,N_19669);
xor UO_1461 (O_1461,N_19626,N_19740);
and UO_1462 (O_1462,N_19240,N_19862);
nor UO_1463 (O_1463,N_19395,N_19892);
xnor UO_1464 (O_1464,N_19745,N_19348);
and UO_1465 (O_1465,N_19261,N_19669);
nand UO_1466 (O_1466,N_19762,N_19694);
or UO_1467 (O_1467,N_19325,N_19509);
xor UO_1468 (O_1468,N_19958,N_19842);
or UO_1469 (O_1469,N_19216,N_19611);
or UO_1470 (O_1470,N_19760,N_19939);
and UO_1471 (O_1471,N_19791,N_19961);
nand UO_1472 (O_1472,N_19385,N_19268);
or UO_1473 (O_1473,N_19801,N_19244);
nor UO_1474 (O_1474,N_19738,N_19526);
nor UO_1475 (O_1475,N_19897,N_19560);
xnor UO_1476 (O_1476,N_19313,N_19455);
or UO_1477 (O_1477,N_19205,N_19281);
xor UO_1478 (O_1478,N_19328,N_19873);
nand UO_1479 (O_1479,N_19735,N_19562);
nor UO_1480 (O_1480,N_19503,N_19213);
xor UO_1481 (O_1481,N_19976,N_19745);
or UO_1482 (O_1482,N_19388,N_19723);
nor UO_1483 (O_1483,N_19815,N_19427);
xor UO_1484 (O_1484,N_19677,N_19539);
and UO_1485 (O_1485,N_19600,N_19591);
nand UO_1486 (O_1486,N_19997,N_19876);
and UO_1487 (O_1487,N_19324,N_19307);
and UO_1488 (O_1488,N_19922,N_19633);
or UO_1489 (O_1489,N_19369,N_19569);
and UO_1490 (O_1490,N_19568,N_19417);
nand UO_1491 (O_1491,N_19367,N_19978);
nand UO_1492 (O_1492,N_19260,N_19553);
xor UO_1493 (O_1493,N_19274,N_19442);
and UO_1494 (O_1494,N_19931,N_19324);
or UO_1495 (O_1495,N_19891,N_19501);
and UO_1496 (O_1496,N_19509,N_19350);
or UO_1497 (O_1497,N_19949,N_19487);
or UO_1498 (O_1498,N_19780,N_19840);
or UO_1499 (O_1499,N_19258,N_19452);
or UO_1500 (O_1500,N_19351,N_19223);
and UO_1501 (O_1501,N_19954,N_19343);
or UO_1502 (O_1502,N_19904,N_19749);
xnor UO_1503 (O_1503,N_19714,N_19356);
or UO_1504 (O_1504,N_19770,N_19939);
nor UO_1505 (O_1505,N_19809,N_19452);
and UO_1506 (O_1506,N_19489,N_19347);
nor UO_1507 (O_1507,N_19908,N_19557);
nor UO_1508 (O_1508,N_19681,N_19728);
and UO_1509 (O_1509,N_19547,N_19756);
xnor UO_1510 (O_1510,N_19956,N_19455);
and UO_1511 (O_1511,N_19561,N_19891);
xnor UO_1512 (O_1512,N_19564,N_19332);
xnor UO_1513 (O_1513,N_19990,N_19895);
nand UO_1514 (O_1514,N_19683,N_19630);
and UO_1515 (O_1515,N_19307,N_19251);
and UO_1516 (O_1516,N_19846,N_19516);
nor UO_1517 (O_1517,N_19403,N_19617);
and UO_1518 (O_1518,N_19489,N_19403);
or UO_1519 (O_1519,N_19923,N_19543);
or UO_1520 (O_1520,N_19280,N_19868);
nor UO_1521 (O_1521,N_19431,N_19440);
nand UO_1522 (O_1522,N_19991,N_19729);
nand UO_1523 (O_1523,N_19346,N_19453);
xor UO_1524 (O_1524,N_19343,N_19962);
nor UO_1525 (O_1525,N_19459,N_19364);
nand UO_1526 (O_1526,N_19479,N_19402);
nand UO_1527 (O_1527,N_19275,N_19797);
and UO_1528 (O_1528,N_19819,N_19773);
nand UO_1529 (O_1529,N_19521,N_19543);
xnor UO_1530 (O_1530,N_19485,N_19403);
nor UO_1531 (O_1531,N_19816,N_19701);
or UO_1532 (O_1532,N_19278,N_19825);
and UO_1533 (O_1533,N_19548,N_19989);
nand UO_1534 (O_1534,N_19677,N_19784);
and UO_1535 (O_1535,N_19619,N_19960);
nand UO_1536 (O_1536,N_19604,N_19641);
and UO_1537 (O_1537,N_19671,N_19828);
nand UO_1538 (O_1538,N_19878,N_19372);
nor UO_1539 (O_1539,N_19661,N_19533);
or UO_1540 (O_1540,N_19724,N_19744);
xnor UO_1541 (O_1541,N_19916,N_19424);
xor UO_1542 (O_1542,N_19201,N_19930);
xor UO_1543 (O_1543,N_19531,N_19397);
nor UO_1544 (O_1544,N_19957,N_19487);
and UO_1545 (O_1545,N_19374,N_19426);
nand UO_1546 (O_1546,N_19834,N_19934);
or UO_1547 (O_1547,N_19914,N_19865);
nand UO_1548 (O_1548,N_19710,N_19452);
or UO_1549 (O_1549,N_19623,N_19941);
xor UO_1550 (O_1550,N_19618,N_19795);
and UO_1551 (O_1551,N_19794,N_19313);
nor UO_1552 (O_1552,N_19717,N_19902);
and UO_1553 (O_1553,N_19467,N_19258);
nor UO_1554 (O_1554,N_19303,N_19920);
nand UO_1555 (O_1555,N_19614,N_19874);
xnor UO_1556 (O_1556,N_19441,N_19893);
and UO_1557 (O_1557,N_19222,N_19340);
nor UO_1558 (O_1558,N_19939,N_19959);
or UO_1559 (O_1559,N_19452,N_19658);
xnor UO_1560 (O_1560,N_19807,N_19885);
nand UO_1561 (O_1561,N_19518,N_19551);
or UO_1562 (O_1562,N_19439,N_19450);
nor UO_1563 (O_1563,N_19225,N_19461);
or UO_1564 (O_1564,N_19755,N_19515);
nor UO_1565 (O_1565,N_19776,N_19267);
nor UO_1566 (O_1566,N_19354,N_19267);
or UO_1567 (O_1567,N_19963,N_19719);
xnor UO_1568 (O_1568,N_19269,N_19707);
xnor UO_1569 (O_1569,N_19825,N_19652);
nor UO_1570 (O_1570,N_19697,N_19916);
or UO_1571 (O_1571,N_19711,N_19980);
or UO_1572 (O_1572,N_19375,N_19502);
or UO_1573 (O_1573,N_19694,N_19330);
nand UO_1574 (O_1574,N_19898,N_19925);
nand UO_1575 (O_1575,N_19573,N_19365);
or UO_1576 (O_1576,N_19351,N_19326);
and UO_1577 (O_1577,N_19365,N_19883);
nand UO_1578 (O_1578,N_19618,N_19672);
xnor UO_1579 (O_1579,N_19806,N_19310);
nor UO_1580 (O_1580,N_19433,N_19284);
nand UO_1581 (O_1581,N_19794,N_19887);
nor UO_1582 (O_1582,N_19758,N_19274);
or UO_1583 (O_1583,N_19906,N_19477);
nand UO_1584 (O_1584,N_19281,N_19671);
or UO_1585 (O_1585,N_19752,N_19438);
and UO_1586 (O_1586,N_19875,N_19304);
nor UO_1587 (O_1587,N_19398,N_19662);
or UO_1588 (O_1588,N_19311,N_19352);
nor UO_1589 (O_1589,N_19992,N_19945);
nor UO_1590 (O_1590,N_19923,N_19893);
xor UO_1591 (O_1591,N_19741,N_19779);
and UO_1592 (O_1592,N_19884,N_19539);
or UO_1593 (O_1593,N_19900,N_19454);
nor UO_1594 (O_1594,N_19800,N_19483);
nor UO_1595 (O_1595,N_19741,N_19342);
nand UO_1596 (O_1596,N_19524,N_19283);
nor UO_1597 (O_1597,N_19992,N_19696);
xor UO_1598 (O_1598,N_19904,N_19815);
nor UO_1599 (O_1599,N_19330,N_19201);
nor UO_1600 (O_1600,N_19487,N_19264);
nand UO_1601 (O_1601,N_19739,N_19515);
nand UO_1602 (O_1602,N_19628,N_19406);
nor UO_1603 (O_1603,N_19268,N_19218);
xnor UO_1604 (O_1604,N_19356,N_19328);
nand UO_1605 (O_1605,N_19232,N_19253);
xor UO_1606 (O_1606,N_19661,N_19435);
or UO_1607 (O_1607,N_19229,N_19280);
and UO_1608 (O_1608,N_19336,N_19708);
xor UO_1609 (O_1609,N_19439,N_19872);
or UO_1610 (O_1610,N_19516,N_19541);
and UO_1611 (O_1611,N_19700,N_19843);
xnor UO_1612 (O_1612,N_19482,N_19942);
xnor UO_1613 (O_1613,N_19695,N_19513);
nand UO_1614 (O_1614,N_19274,N_19655);
and UO_1615 (O_1615,N_19797,N_19351);
nand UO_1616 (O_1616,N_19800,N_19439);
and UO_1617 (O_1617,N_19353,N_19294);
xor UO_1618 (O_1618,N_19278,N_19518);
nor UO_1619 (O_1619,N_19899,N_19508);
nor UO_1620 (O_1620,N_19756,N_19789);
and UO_1621 (O_1621,N_19259,N_19992);
or UO_1622 (O_1622,N_19601,N_19705);
and UO_1623 (O_1623,N_19986,N_19695);
xnor UO_1624 (O_1624,N_19934,N_19993);
xor UO_1625 (O_1625,N_19368,N_19768);
and UO_1626 (O_1626,N_19469,N_19895);
xor UO_1627 (O_1627,N_19782,N_19973);
nor UO_1628 (O_1628,N_19470,N_19500);
and UO_1629 (O_1629,N_19627,N_19411);
and UO_1630 (O_1630,N_19314,N_19566);
and UO_1631 (O_1631,N_19382,N_19832);
nand UO_1632 (O_1632,N_19707,N_19921);
nor UO_1633 (O_1633,N_19335,N_19420);
xnor UO_1634 (O_1634,N_19409,N_19526);
nor UO_1635 (O_1635,N_19904,N_19932);
nand UO_1636 (O_1636,N_19663,N_19209);
or UO_1637 (O_1637,N_19499,N_19702);
xor UO_1638 (O_1638,N_19317,N_19306);
or UO_1639 (O_1639,N_19599,N_19256);
xor UO_1640 (O_1640,N_19730,N_19822);
or UO_1641 (O_1641,N_19556,N_19807);
xor UO_1642 (O_1642,N_19766,N_19845);
xnor UO_1643 (O_1643,N_19218,N_19489);
and UO_1644 (O_1644,N_19973,N_19430);
nand UO_1645 (O_1645,N_19378,N_19451);
nor UO_1646 (O_1646,N_19791,N_19955);
or UO_1647 (O_1647,N_19413,N_19588);
nand UO_1648 (O_1648,N_19920,N_19906);
nor UO_1649 (O_1649,N_19635,N_19925);
nand UO_1650 (O_1650,N_19987,N_19295);
and UO_1651 (O_1651,N_19264,N_19426);
nand UO_1652 (O_1652,N_19781,N_19943);
xor UO_1653 (O_1653,N_19633,N_19391);
and UO_1654 (O_1654,N_19209,N_19660);
xnor UO_1655 (O_1655,N_19782,N_19548);
nand UO_1656 (O_1656,N_19590,N_19692);
nor UO_1657 (O_1657,N_19421,N_19735);
nor UO_1658 (O_1658,N_19712,N_19215);
nor UO_1659 (O_1659,N_19806,N_19339);
nand UO_1660 (O_1660,N_19762,N_19421);
or UO_1661 (O_1661,N_19336,N_19211);
nand UO_1662 (O_1662,N_19888,N_19432);
and UO_1663 (O_1663,N_19662,N_19582);
xor UO_1664 (O_1664,N_19741,N_19236);
nand UO_1665 (O_1665,N_19760,N_19729);
nor UO_1666 (O_1666,N_19697,N_19385);
nand UO_1667 (O_1667,N_19510,N_19972);
xnor UO_1668 (O_1668,N_19445,N_19809);
nand UO_1669 (O_1669,N_19226,N_19516);
nand UO_1670 (O_1670,N_19689,N_19614);
nor UO_1671 (O_1671,N_19270,N_19630);
or UO_1672 (O_1672,N_19981,N_19252);
nand UO_1673 (O_1673,N_19977,N_19508);
and UO_1674 (O_1674,N_19600,N_19808);
nand UO_1675 (O_1675,N_19959,N_19370);
xor UO_1676 (O_1676,N_19950,N_19597);
and UO_1677 (O_1677,N_19956,N_19764);
nand UO_1678 (O_1678,N_19939,N_19440);
and UO_1679 (O_1679,N_19770,N_19488);
nor UO_1680 (O_1680,N_19887,N_19548);
xnor UO_1681 (O_1681,N_19556,N_19285);
nand UO_1682 (O_1682,N_19254,N_19565);
or UO_1683 (O_1683,N_19259,N_19456);
nor UO_1684 (O_1684,N_19688,N_19856);
or UO_1685 (O_1685,N_19692,N_19598);
xnor UO_1686 (O_1686,N_19905,N_19843);
or UO_1687 (O_1687,N_19313,N_19470);
or UO_1688 (O_1688,N_19487,N_19508);
nand UO_1689 (O_1689,N_19981,N_19705);
nand UO_1690 (O_1690,N_19415,N_19826);
and UO_1691 (O_1691,N_19800,N_19520);
xor UO_1692 (O_1692,N_19488,N_19711);
nor UO_1693 (O_1693,N_19573,N_19823);
nor UO_1694 (O_1694,N_19786,N_19643);
or UO_1695 (O_1695,N_19834,N_19291);
nor UO_1696 (O_1696,N_19518,N_19950);
nand UO_1697 (O_1697,N_19970,N_19502);
xor UO_1698 (O_1698,N_19687,N_19709);
xnor UO_1699 (O_1699,N_19204,N_19525);
nand UO_1700 (O_1700,N_19948,N_19232);
nand UO_1701 (O_1701,N_19471,N_19207);
or UO_1702 (O_1702,N_19633,N_19474);
nor UO_1703 (O_1703,N_19853,N_19576);
or UO_1704 (O_1704,N_19828,N_19887);
nor UO_1705 (O_1705,N_19971,N_19305);
nand UO_1706 (O_1706,N_19825,N_19333);
or UO_1707 (O_1707,N_19713,N_19683);
nand UO_1708 (O_1708,N_19572,N_19787);
nor UO_1709 (O_1709,N_19643,N_19626);
nand UO_1710 (O_1710,N_19385,N_19226);
nand UO_1711 (O_1711,N_19515,N_19700);
nor UO_1712 (O_1712,N_19425,N_19515);
or UO_1713 (O_1713,N_19271,N_19754);
nor UO_1714 (O_1714,N_19882,N_19613);
xnor UO_1715 (O_1715,N_19586,N_19563);
or UO_1716 (O_1716,N_19734,N_19917);
nand UO_1717 (O_1717,N_19998,N_19805);
xor UO_1718 (O_1718,N_19703,N_19455);
nor UO_1719 (O_1719,N_19817,N_19769);
nand UO_1720 (O_1720,N_19327,N_19677);
and UO_1721 (O_1721,N_19746,N_19482);
nor UO_1722 (O_1722,N_19931,N_19309);
nand UO_1723 (O_1723,N_19571,N_19746);
nand UO_1724 (O_1724,N_19542,N_19282);
xnor UO_1725 (O_1725,N_19534,N_19852);
nand UO_1726 (O_1726,N_19287,N_19472);
nand UO_1727 (O_1727,N_19641,N_19246);
nor UO_1728 (O_1728,N_19201,N_19305);
nor UO_1729 (O_1729,N_19331,N_19851);
or UO_1730 (O_1730,N_19303,N_19457);
and UO_1731 (O_1731,N_19650,N_19207);
xnor UO_1732 (O_1732,N_19494,N_19395);
xnor UO_1733 (O_1733,N_19306,N_19985);
xor UO_1734 (O_1734,N_19569,N_19473);
or UO_1735 (O_1735,N_19212,N_19741);
nor UO_1736 (O_1736,N_19955,N_19906);
and UO_1737 (O_1737,N_19482,N_19628);
or UO_1738 (O_1738,N_19252,N_19514);
or UO_1739 (O_1739,N_19802,N_19208);
xor UO_1740 (O_1740,N_19368,N_19965);
or UO_1741 (O_1741,N_19758,N_19930);
xnor UO_1742 (O_1742,N_19492,N_19202);
or UO_1743 (O_1743,N_19576,N_19911);
and UO_1744 (O_1744,N_19597,N_19457);
or UO_1745 (O_1745,N_19429,N_19620);
nand UO_1746 (O_1746,N_19569,N_19796);
xnor UO_1747 (O_1747,N_19425,N_19802);
and UO_1748 (O_1748,N_19714,N_19809);
nand UO_1749 (O_1749,N_19209,N_19415);
or UO_1750 (O_1750,N_19484,N_19888);
or UO_1751 (O_1751,N_19979,N_19500);
xnor UO_1752 (O_1752,N_19240,N_19359);
nand UO_1753 (O_1753,N_19297,N_19292);
xor UO_1754 (O_1754,N_19647,N_19732);
nor UO_1755 (O_1755,N_19850,N_19959);
and UO_1756 (O_1756,N_19829,N_19646);
nand UO_1757 (O_1757,N_19226,N_19589);
xor UO_1758 (O_1758,N_19440,N_19963);
and UO_1759 (O_1759,N_19776,N_19341);
nor UO_1760 (O_1760,N_19826,N_19908);
or UO_1761 (O_1761,N_19518,N_19352);
nand UO_1762 (O_1762,N_19418,N_19411);
and UO_1763 (O_1763,N_19993,N_19933);
nand UO_1764 (O_1764,N_19471,N_19811);
and UO_1765 (O_1765,N_19683,N_19633);
nor UO_1766 (O_1766,N_19404,N_19924);
or UO_1767 (O_1767,N_19992,N_19332);
and UO_1768 (O_1768,N_19256,N_19821);
xor UO_1769 (O_1769,N_19447,N_19570);
nand UO_1770 (O_1770,N_19264,N_19235);
and UO_1771 (O_1771,N_19806,N_19477);
and UO_1772 (O_1772,N_19675,N_19312);
and UO_1773 (O_1773,N_19885,N_19816);
and UO_1774 (O_1774,N_19539,N_19208);
nor UO_1775 (O_1775,N_19890,N_19658);
nand UO_1776 (O_1776,N_19942,N_19398);
and UO_1777 (O_1777,N_19252,N_19742);
nand UO_1778 (O_1778,N_19247,N_19666);
nor UO_1779 (O_1779,N_19852,N_19920);
nand UO_1780 (O_1780,N_19201,N_19711);
or UO_1781 (O_1781,N_19665,N_19351);
or UO_1782 (O_1782,N_19966,N_19426);
nand UO_1783 (O_1783,N_19411,N_19377);
nand UO_1784 (O_1784,N_19322,N_19712);
or UO_1785 (O_1785,N_19917,N_19314);
nand UO_1786 (O_1786,N_19696,N_19409);
xor UO_1787 (O_1787,N_19803,N_19751);
and UO_1788 (O_1788,N_19454,N_19735);
and UO_1789 (O_1789,N_19455,N_19545);
or UO_1790 (O_1790,N_19346,N_19848);
or UO_1791 (O_1791,N_19738,N_19872);
nor UO_1792 (O_1792,N_19696,N_19293);
and UO_1793 (O_1793,N_19683,N_19688);
nor UO_1794 (O_1794,N_19670,N_19675);
xor UO_1795 (O_1795,N_19540,N_19508);
xor UO_1796 (O_1796,N_19586,N_19255);
xnor UO_1797 (O_1797,N_19218,N_19982);
nor UO_1798 (O_1798,N_19680,N_19330);
nor UO_1799 (O_1799,N_19508,N_19802);
nor UO_1800 (O_1800,N_19930,N_19486);
and UO_1801 (O_1801,N_19579,N_19416);
nor UO_1802 (O_1802,N_19579,N_19381);
nor UO_1803 (O_1803,N_19660,N_19262);
nand UO_1804 (O_1804,N_19745,N_19889);
or UO_1805 (O_1805,N_19916,N_19827);
nand UO_1806 (O_1806,N_19581,N_19444);
nor UO_1807 (O_1807,N_19577,N_19681);
nor UO_1808 (O_1808,N_19266,N_19633);
nor UO_1809 (O_1809,N_19929,N_19533);
nand UO_1810 (O_1810,N_19734,N_19462);
xor UO_1811 (O_1811,N_19839,N_19572);
and UO_1812 (O_1812,N_19839,N_19219);
or UO_1813 (O_1813,N_19268,N_19802);
or UO_1814 (O_1814,N_19313,N_19271);
or UO_1815 (O_1815,N_19581,N_19830);
or UO_1816 (O_1816,N_19754,N_19496);
and UO_1817 (O_1817,N_19387,N_19284);
or UO_1818 (O_1818,N_19974,N_19443);
nor UO_1819 (O_1819,N_19271,N_19863);
nand UO_1820 (O_1820,N_19490,N_19494);
or UO_1821 (O_1821,N_19876,N_19859);
nand UO_1822 (O_1822,N_19292,N_19461);
xnor UO_1823 (O_1823,N_19637,N_19504);
and UO_1824 (O_1824,N_19734,N_19340);
xor UO_1825 (O_1825,N_19440,N_19457);
nor UO_1826 (O_1826,N_19393,N_19297);
and UO_1827 (O_1827,N_19880,N_19860);
and UO_1828 (O_1828,N_19581,N_19293);
nand UO_1829 (O_1829,N_19884,N_19716);
nor UO_1830 (O_1830,N_19898,N_19248);
nor UO_1831 (O_1831,N_19880,N_19974);
and UO_1832 (O_1832,N_19920,N_19366);
nand UO_1833 (O_1833,N_19855,N_19774);
nor UO_1834 (O_1834,N_19309,N_19850);
and UO_1835 (O_1835,N_19880,N_19273);
nand UO_1836 (O_1836,N_19813,N_19900);
xor UO_1837 (O_1837,N_19252,N_19933);
nand UO_1838 (O_1838,N_19277,N_19233);
xor UO_1839 (O_1839,N_19201,N_19359);
nor UO_1840 (O_1840,N_19425,N_19748);
or UO_1841 (O_1841,N_19773,N_19647);
and UO_1842 (O_1842,N_19326,N_19647);
xnor UO_1843 (O_1843,N_19948,N_19383);
nand UO_1844 (O_1844,N_19397,N_19662);
nor UO_1845 (O_1845,N_19623,N_19467);
nand UO_1846 (O_1846,N_19450,N_19509);
and UO_1847 (O_1847,N_19587,N_19873);
nor UO_1848 (O_1848,N_19342,N_19920);
and UO_1849 (O_1849,N_19269,N_19209);
nor UO_1850 (O_1850,N_19296,N_19961);
nand UO_1851 (O_1851,N_19538,N_19518);
or UO_1852 (O_1852,N_19716,N_19561);
nor UO_1853 (O_1853,N_19493,N_19484);
nand UO_1854 (O_1854,N_19836,N_19235);
xnor UO_1855 (O_1855,N_19581,N_19677);
nor UO_1856 (O_1856,N_19710,N_19580);
or UO_1857 (O_1857,N_19759,N_19571);
and UO_1858 (O_1858,N_19438,N_19765);
nand UO_1859 (O_1859,N_19940,N_19233);
nand UO_1860 (O_1860,N_19611,N_19570);
xor UO_1861 (O_1861,N_19370,N_19973);
xor UO_1862 (O_1862,N_19720,N_19624);
or UO_1863 (O_1863,N_19359,N_19402);
and UO_1864 (O_1864,N_19993,N_19657);
xnor UO_1865 (O_1865,N_19647,N_19718);
or UO_1866 (O_1866,N_19240,N_19502);
nor UO_1867 (O_1867,N_19726,N_19824);
xnor UO_1868 (O_1868,N_19325,N_19204);
and UO_1869 (O_1869,N_19758,N_19736);
and UO_1870 (O_1870,N_19992,N_19338);
xnor UO_1871 (O_1871,N_19708,N_19957);
xnor UO_1872 (O_1872,N_19674,N_19926);
xnor UO_1873 (O_1873,N_19542,N_19857);
nand UO_1874 (O_1874,N_19590,N_19308);
nand UO_1875 (O_1875,N_19602,N_19350);
nand UO_1876 (O_1876,N_19427,N_19888);
and UO_1877 (O_1877,N_19814,N_19912);
or UO_1878 (O_1878,N_19945,N_19368);
nand UO_1879 (O_1879,N_19966,N_19342);
or UO_1880 (O_1880,N_19956,N_19997);
xnor UO_1881 (O_1881,N_19732,N_19407);
and UO_1882 (O_1882,N_19674,N_19975);
xnor UO_1883 (O_1883,N_19788,N_19448);
nor UO_1884 (O_1884,N_19703,N_19324);
and UO_1885 (O_1885,N_19629,N_19472);
or UO_1886 (O_1886,N_19634,N_19976);
and UO_1887 (O_1887,N_19490,N_19325);
and UO_1888 (O_1888,N_19321,N_19202);
nand UO_1889 (O_1889,N_19232,N_19620);
or UO_1890 (O_1890,N_19658,N_19674);
or UO_1891 (O_1891,N_19899,N_19649);
and UO_1892 (O_1892,N_19369,N_19768);
nand UO_1893 (O_1893,N_19885,N_19248);
or UO_1894 (O_1894,N_19959,N_19575);
or UO_1895 (O_1895,N_19816,N_19699);
nor UO_1896 (O_1896,N_19443,N_19898);
and UO_1897 (O_1897,N_19292,N_19870);
nor UO_1898 (O_1898,N_19317,N_19346);
or UO_1899 (O_1899,N_19479,N_19637);
or UO_1900 (O_1900,N_19583,N_19358);
xor UO_1901 (O_1901,N_19608,N_19879);
nor UO_1902 (O_1902,N_19510,N_19764);
nand UO_1903 (O_1903,N_19852,N_19362);
and UO_1904 (O_1904,N_19934,N_19303);
or UO_1905 (O_1905,N_19267,N_19250);
or UO_1906 (O_1906,N_19957,N_19790);
nor UO_1907 (O_1907,N_19373,N_19765);
nor UO_1908 (O_1908,N_19793,N_19710);
xnor UO_1909 (O_1909,N_19699,N_19489);
nand UO_1910 (O_1910,N_19818,N_19775);
or UO_1911 (O_1911,N_19630,N_19723);
nor UO_1912 (O_1912,N_19903,N_19521);
nor UO_1913 (O_1913,N_19575,N_19230);
and UO_1914 (O_1914,N_19826,N_19718);
and UO_1915 (O_1915,N_19581,N_19401);
xor UO_1916 (O_1916,N_19950,N_19542);
nor UO_1917 (O_1917,N_19489,N_19631);
nand UO_1918 (O_1918,N_19634,N_19360);
xor UO_1919 (O_1919,N_19703,N_19953);
and UO_1920 (O_1920,N_19409,N_19791);
nand UO_1921 (O_1921,N_19324,N_19448);
nand UO_1922 (O_1922,N_19461,N_19203);
or UO_1923 (O_1923,N_19712,N_19329);
and UO_1924 (O_1924,N_19217,N_19972);
xnor UO_1925 (O_1925,N_19555,N_19685);
or UO_1926 (O_1926,N_19450,N_19917);
nor UO_1927 (O_1927,N_19248,N_19764);
or UO_1928 (O_1928,N_19618,N_19620);
or UO_1929 (O_1929,N_19908,N_19346);
xor UO_1930 (O_1930,N_19919,N_19338);
or UO_1931 (O_1931,N_19534,N_19606);
or UO_1932 (O_1932,N_19265,N_19343);
nand UO_1933 (O_1933,N_19711,N_19588);
nand UO_1934 (O_1934,N_19357,N_19673);
and UO_1935 (O_1935,N_19659,N_19718);
nand UO_1936 (O_1936,N_19228,N_19513);
or UO_1937 (O_1937,N_19574,N_19738);
nand UO_1938 (O_1938,N_19270,N_19420);
or UO_1939 (O_1939,N_19950,N_19255);
xor UO_1940 (O_1940,N_19603,N_19963);
nand UO_1941 (O_1941,N_19427,N_19664);
nand UO_1942 (O_1942,N_19349,N_19323);
and UO_1943 (O_1943,N_19849,N_19742);
nor UO_1944 (O_1944,N_19758,N_19874);
nor UO_1945 (O_1945,N_19341,N_19826);
or UO_1946 (O_1946,N_19944,N_19877);
and UO_1947 (O_1947,N_19869,N_19940);
nor UO_1948 (O_1948,N_19646,N_19246);
and UO_1949 (O_1949,N_19323,N_19777);
and UO_1950 (O_1950,N_19907,N_19368);
or UO_1951 (O_1951,N_19259,N_19321);
nor UO_1952 (O_1952,N_19600,N_19700);
xnor UO_1953 (O_1953,N_19567,N_19383);
xnor UO_1954 (O_1954,N_19513,N_19929);
or UO_1955 (O_1955,N_19660,N_19688);
and UO_1956 (O_1956,N_19685,N_19407);
xor UO_1957 (O_1957,N_19640,N_19268);
xor UO_1958 (O_1958,N_19601,N_19663);
xnor UO_1959 (O_1959,N_19645,N_19317);
and UO_1960 (O_1960,N_19372,N_19376);
and UO_1961 (O_1961,N_19460,N_19774);
nor UO_1962 (O_1962,N_19690,N_19413);
nand UO_1963 (O_1963,N_19654,N_19215);
or UO_1964 (O_1964,N_19711,N_19619);
or UO_1965 (O_1965,N_19350,N_19905);
and UO_1966 (O_1966,N_19890,N_19598);
nor UO_1967 (O_1967,N_19346,N_19435);
nand UO_1968 (O_1968,N_19602,N_19271);
nand UO_1969 (O_1969,N_19537,N_19962);
xnor UO_1970 (O_1970,N_19779,N_19852);
and UO_1971 (O_1971,N_19420,N_19607);
and UO_1972 (O_1972,N_19865,N_19686);
or UO_1973 (O_1973,N_19790,N_19912);
xnor UO_1974 (O_1974,N_19303,N_19719);
xor UO_1975 (O_1975,N_19468,N_19921);
and UO_1976 (O_1976,N_19594,N_19452);
nand UO_1977 (O_1977,N_19488,N_19272);
xnor UO_1978 (O_1978,N_19260,N_19571);
nor UO_1979 (O_1979,N_19840,N_19876);
nand UO_1980 (O_1980,N_19700,N_19891);
and UO_1981 (O_1981,N_19912,N_19624);
xor UO_1982 (O_1982,N_19503,N_19867);
or UO_1983 (O_1983,N_19369,N_19763);
or UO_1984 (O_1984,N_19331,N_19840);
or UO_1985 (O_1985,N_19972,N_19777);
xnor UO_1986 (O_1986,N_19867,N_19972);
nor UO_1987 (O_1987,N_19559,N_19680);
or UO_1988 (O_1988,N_19647,N_19305);
nand UO_1989 (O_1989,N_19580,N_19470);
and UO_1990 (O_1990,N_19543,N_19935);
and UO_1991 (O_1991,N_19342,N_19505);
nor UO_1992 (O_1992,N_19484,N_19693);
and UO_1993 (O_1993,N_19206,N_19811);
xor UO_1994 (O_1994,N_19332,N_19249);
nand UO_1995 (O_1995,N_19928,N_19211);
or UO_1996 (O_1996,N_19971,N_19586);
or UO_1997 (O_1997,N_19957,N_19723);
xnor UO_1998 (O_1998,N_19361,N_19200);
and UO_1999 (O_1999,N_19833,N_19665);
nand UO_2000 (O_2000,N_19920,N_19961);
nand UO_2001 (O_2001,N_19343,N_19640);
or UO_2002 (O_2002,N_19514,N_19611);
nor UO_2003 (O_2003,N_19727,N_19605);
and UO_2004 (O_2004,N_19294,N_19560);
nand UO_2005 (O_2005,N_19769,N_19251);
nor UO_2006 (O_2006,N_19711,N_19777);
or UO_2007 (O_2007,N_19699,N_19344);
nor UO_2008 (O_2008,N_19673,N_19782);
nand UO_2009 (O_2009,N_19748,N_19501);
or UO_2010 (O_2010,N_19278,N_19621);
nand UO_2011 (O_2011,N_19998,N_19944);
xor UO_2012 (O_2012,N_19416,N_19293);
and UO_2013 (O_2013,N_19236,N_19835);
nand UO_2014 (O_2014,N_19969,N_19504);
nor UO_2015 (O_2015,N_19489,N_19374);
nor UO_2016 (O_2016,N_19713,N_19699);
and UO_2017 (O_2017,N_19914,N_19288);
xor UO_2018 (O_2018,N_19582,N_19401);
or UO_2019 (O_2019,N_19695,N_19982);
or UO_2020 (O_2020,N_19782,N_19275);
nor UO_2021 (O_2021,N_19979,N_19266);
nand UO_2022 (O_2022,N_19490,N_19554);
and UO_2023 (O_2023,N_19211,N_19597);
and UO_2024 (O_2024,N_19869,N_19245);
nor UO_2025 (O_2025,N_19891,N_19571);
and UO_2026 (O_2026,N_19217,N_19304);
nand UO_2027 (O_2027,N_19337,N_19364);
xor UO_2028 (O_2028,N_19968,N_19507);
nor UO_2029 (O_2029,N_19498,N_19920);
or UO_2030 (O_2030,N_19596,N_19245);
and UO_2031 (O_2031,N_19442,N_19259);
xor UO_2032 (O_2032,N_19859,N_19852);
nand UO_2033 (O_2033,N_19221,N_19487);
or UO_2034 (O_2034,N_19404,N_19418);
or UO_2035 (O_2035,N_19616,N_19431);
nand UO_2036 (O_2036,N_19930,N_19464);
nor UO_2037 (O_2037,N_19893,N_19547);
nand UO_2038 (O_2038,N_19427,N_19436);
and UO_2039 (O_2039,N_19915,N_19791);
or UO_2040 (O_2040,N_19333,N_19907);
nor UO_2041 (O_2041,N_19357,N_19979);
nor UO_2042 (O_2042,N_19522,N_19508);
and UO_2043 (O_2043,N_19608,N_19417);
or UO_2044 (O_2044,N_19746,N_19329);
and UO_2045 (O_2045,N_19886,N_19511);
or UO_2046 (O_2046,N_19588,N_19766);
xnor UO_2047 (O_2047,N_19847,N_19288);
or UO_2048 (O_2048,N_19481,N_19949);
nor UO_2049 (O_2049,N_19285,N_19808);
and UO_2050 (O_2050,N_19972,N_19220);
and UO_2051 (O_2051,N_19831,N_19925);
or UO_2052 (O_2052,N_19356,N_19600);
nand UO_2053 (O_2053,N_19547,N_19465);
or UO_2054 (O_2054,N_19594,N_19738);
or UO_2055 (O_2055,N_19553,N_19552);
nor UO_2056 (O_2056,N_19826,N_19726);
nand UO_2057 (O_2057,N_19411,N_19796);
and UO_2058 (O_2058,N_19820,N_19362);
nor UO_2059 (O_2059,N_19541,N_19494);
nor UO_2060 (O_2060,N_19486,N_19418);
and UO_2061 (O_2061,N_19233,N_19534);
or UO_2062 (O_2062,N_19663,N_19367);
xor UO_2063 (O_2063,N_19504,N_19280);
nand UO_2064 (O_2064,N_19338,N_19504);
nor UO_2065 (O_2065,N_19474,N_19207);
or UO_2066 (O_2066,N_19626,N_19229);
nand UO_2067 (O_2067,N_19955,N_19619);
or UO_2068 (O_2068,N_19211,N_19835);
or UO_2069 (O_2069,N_19862,N_19329);
nor UO_2070 (O_2070,N_19531,N_19555);
and UO_2071 (O_2071,N_19949,N_19365);
or UO_2072 (O_2072,N_19855,N_19575);
xnor UO_2073 (O_2073,N_19278,N_19692);
or UO_2074 (O_2074,N_19561,N_19269);
and UO_2075 (O_2075,N_19749,N_19392);
or UO_2076 (O_2076,N_19513,N_19714);
nor UO_2077 (O_2077,N_19412,N_19513);
or UO_2078 (O_2078,N_19497,N_19323);
nand UO_2079 (O_2079,N_19626,N_19293);
nor UO_2080 (O_2080,N_19510,N_19945);
nand UO_2081 (O_2081,N_19258,N_19982);
nor UO_2082 (O_2082,N_19610,N_19304);
nand UO_2083 (O_2083,N_19550,N_19241);
or UO_2084 (O_2084,N_19429,N_19231);
nor UO_2085 (O_2085,N_19583,N_19702);
xor UO_2086 (O_2086,N_19510,N_19738);
nand UO_2087 (O_2087,N_19217,N_19332);
nor UO_2088 (O_2088,N_19667,N_19749);
xnor UO_2089 (O_2089,N_19619,N_19292);
and UO_2090 (O_2090,N_19376,N_19405);
nand UO_2091 (O_2091,N_19841,N_19787);
nand UO_2092 (O_2092,N_19374,N_19537);
xor UO_2093 (O_2093,N_19769,N_19942);
nand UO_2094 (O_2094,N_19309,N_19845);
nand UO_2095 (O_2095,N_19759,N_19615);
xor UO_2096 (O_2096,N_19462,N_19301);
xor UO_2097 (O_2097,N_19662,N_19994);
xnor UO_2098 (O_2098,N_19848,N_19699);
or UO_2099 (O_2099,N_19698,N_19935);
xor UO_2100 (O_2100,N_19959,N_19978);
and UO_2101 (O_2101,N_19688,N_19627);
nand UO_2102 (O_2102,N_19279,N_19496);
or UO_2103 (O_2103,N_19601,N_19379);
nor UO_2104 (O_2104,N_19532,N_19724);
or UO_2105 (O_2105,N_19888,N_19998);
xor UO_2106 (O_2106,N_19413,N_19444);
nor UO_2107 (O_2107,N_19253,N_19401);
or UO_2108 (O_2108,N_19379,N_19306);
or UO_2109 (O_2109,N_19262,N_19668);
and UO_2110 (O_2110,N_19786,N_19820);
nand UO_2111 (O_2111,N_19799,N_19764);
and UO_2112 (O_2112,N_19245,N_19693);
nor UO_2113 (O_2113,N_19382,N_19801);
nand UO_2114 (O_2114,N_19536,N_19396);
nor UO_2115 (O_2115,N_19822,N_19646);
or UO_2116 (O_2116,N_19812,N_19720);
xor UO_2117 (O_2117,N_19959,N_19658);
and UO_2118 (O_2118,N_19802,N_19947);
xor UO_2119 (O_2119,N_19973,N_19495);
nor UO_2120 (O_2120,N_19437,N_19624);
nand UO_2121 (O_2121,N_19311,N_19503);
and UO_2122 (O_2122,N_19826,N_19967);
or UO_2123 (O_2123,N_19826,N_19663);
nand UO_2124 (O_2124,N_19784,N_19912);
nand UO_2125 (O_2125,N_19301,N_19516);
nand UO_2126 (O_2126,N_19690,N_19628);
nor UO_2127 (O_2127,N_19663,N_19526);
nor UO_2128 (O_2128,N_19412,N_19887);
nor UO_2129 (O_2129,N_19868,N_19434);
xnor UO_2130 (O_2130,N_19524,N_19757);
nor UO_2131 (O_2131,N_19674,N_19638);
xor UO_2132 (O_2132,N_19661,N_19715);
or UO_2133 (O_2133,N_19556,N_19248);
or UO_2134 (O_2134,N_19381,N_19311);
or UO_2135 (O_2135,N_19211,N_19491);
xor UO_2136 (O_2136,N_19908,N_19261);
nor UO_2137 (O_2137,N_19892,N_19342);
xnor UO_2138 (O_2138,N_19794,N_19445);
and UO_2139 (O_2139,N_19267,N_19670);
nand UO_2140 (O_2140,N_19606,N_19271);
nor UO_2141 (O_2141,N_19491,N_19315);
or UO_2142 (O_2142,N_19884,N_19261);
or UO_2143 (O_2143,N_19728,N_19989);
and UO_2144 (O_2144,N_19314,N_19887);
xnor UO_2145 (O_2145,N_19850,N_19357);
xnor UO_2146 (O_2146,N_19503,N_19223);
or UO_2147 (O_2147,N_19876,N_19861);
xor UO_2148 (O_2148,N_19460,N_19988);
and UO_2149 (O_2149,N_19400,N_19646);
nor UO_2150 (O_2150,N_19584,N_19467);
and UO_2151 (O_2151,N_19855,N_19666);
or UO_2152 (O_2152,N_19685,N_19354);
xnor UO_2153 (O_2153,N_19627,N_19577);
and UO_2154 (O_2154,N_19972,N_19734);
or UO_2155 (O_2155,N_19287,N_19667);
xor UO_2156 (O_2156,N_19698,N_19617);
nor UO_2157 (O_2157,N_19220,N_19501);
nand UO_2158 (O_2158,N_19906,N_19764);
nor UO_2159 (O_2159,N_19298,N_19746);
or UO_2160 (O_2160,N_19438,N_19216);
nor UO_2161 (O_2161,N_19541,N_19275);
nor UO_2162 (O_2162,N_19278,N_19292);
xnor UO_2163 (O_2163,N_19620,N_19962);
nand UO_2164 (O_2164,N_19279,N_19390);
nor UO_2165 (O_2165,N_19497,N_19464);
xnor UO_2166 (O_2166,N_19778,N_19663);
and UO_2167 (O_2167,N_19950,N_19265);
nor UO_2168 (O_2168,N_19326,N_19606);
or UO_2169 (O_2169,N_19697,N_19226);
nor UO_2170 (O_2170,N_19499,N_19801);
and UO_2171 (O_2171,N_19351,N_19691);
xor UO_2172 (O_2172,N_19274,N_19478);
and UO_2173 (O_2173,N_19491,N_19265);
and UO_2174 (O_2174,N_19646,N_19514);
nand UO_2175 (O_2175,N_19417,N_19548);
nand UO_2176 (O_2176,N_19528,N_19676);
and UO_2177 (O_2177,N_19487,N_19795);
nor UO_2178 (O_2178,N_19468,N_19673);
nor UO_2179 (O_2179,N_19499,N_19954);
and UO_2180 (O_2180,N_19527,N_19297);
nor UO_2181 (O_2181,N_19795,N_19855);
or UO_2182 (O_2182,N_19398,N_19725);
and UO_2183 (O_2183,N_19606,N_19907);
or UO_2184 (O_2184,N_19756,N_19933);
or UO_2185 (O_2185,N_19359,N_19477);
or UO_2186 (O_2186,N_19937,N_19529);
or UO_2187 (O_2187,N_19350,N_19479);
nand UO_2188 (O_2188,N_19242,N_19628);
and UO_2189 (O_2189,N_19465,N_19347);
and UO_2190 (O_2190,N_19278,N_19434);
or UO_2191 (O_2191,N_19643,N_19510);
or UO_2192 (O_2192,N_19877,N_19895);
or UO_2193 (O_2193,N_19594,N_19961);
nor UO_2194 (O_2194,N_19271,N_19220);
or UO_2195 (O_2195,N_19814,N_19445);
nor UO_2196 (O_2196,N_19988,N_19924);
nor UO_2197 (O_2197,N_19681,N_19226);
and UO_2198 (O_2198,N_19281,N_19711);
xor UO_2199 (O_2199,N_19995,N_19492);
or UO_2200 (O_2200,N_19702,N_19860);
or UO_2201 (O_2201,N_19858,N_19552);
xnor UO_2202 (O_2202,N_19257,N_19319);
or UO_2203 (O_2203,N_19404,N_19744);
or UO_2204 (O_2204,N_19767,N_19785);
nor UO_2205 (O_2205,N_19592,N_19401);
xnor UO_2206 (O_2206,N_19999,N_19827);
or UO_2207 (O_2207,N_19459,N_19711);
and UO_2208 (O_2208,N_19456,N_19403);
nor UO_2209 (O_2209,N_19778,N_19405);
and UO_2210 (O_2210,N_19244,N_19482);
nor UO_2211 (O_2211,N_19695,N_19797);
nand UO_2212 (O_2212,N_19355,N_19937);
nor UO_2213 (O_2213,N_19702,N_19537);
xnor UO_2214 (O_2214,N_19257,N_19393);
nand UO_2215 (O_2215,N_19730,N_19729);
nand UO_2216 (O_2216,N_19539,N_19436);
or UO_2217 (O_2217,N_19524,N_19800);
nand UO_2218 (O_2218,N_19550,N_19376);
nor UO_2219 (O_2219,N_19636,N_19682);
xor UO_2220 (O_2220,N_19505,N_19563);
or UO_2221 (O_2221,N_19448,N_19377);
nand UO_2222 (O_2222,N_19598,N_19238);
xnor UO_2223 (O_2223,N_19227,N_19500);
xor UO_2224 (O_2224,N_19692,N_19779);
or UO_2225 (O_2225,N_19800,N_19791);
and UO_2226 (O_2226,N_19861,N_19710);
and UO_2227 (O_2227,N_19382,N_19917);
and UO_2228 (O_2228,N_19541,N_19567);
and UO_2229 (O_2229,N_19629,N_19851);
and UO_2230 (O_2230,N_19606,N_19369);
xor UO_2231 (O_2231,N_19885,N_19957);
or UO_2232 (O_2232,N_19221,N_19734);
nor UO_2233 (O_2233,N_19838,N_19870);
xnor UO_2234 (O_2234,N_19388,N_19201);
nand UO_2235 (O_2235,N_19676,N_19916);
nand UO_2236 (O_2236,N_19713,N_19992);
nor UO_2237 (O_2237,N_19907,N_19647);
or UO_2238 (O_2238,N_19570,N_19425);
nand UO_2239 (O_2239,N_19951,N_19585);
or UO_2240 (O_2240,N_19360,N_19644);
or UO_2241 (O_2241,N_19509,N_19527);
or UO_2242 (O_2242,N_19508,N_19945);
nand UO_2243 (O_2243,N_19937,N_19656);
nor UO_2244 (O_2244,N_19341,N_19357);
nor UO_2245 (O_2245,N_19650,N_19713);
or UO_2246 (O_2246,N_19838,N_19825);
nor UO_2247 (O_2247,N_19958,N_19758);
and UO_2248 (O_2248,N_19234,N_19933);
nor UO_2249 (O_2249,N_19605,N_19312);
or UO_2250 (O_2250,N_19334,N_19718);
and UO_2251 (O_2251,N_19468,N_19476);
or UO_2252 (O_2252,N_19724,N_19785);
and UO_2253 (O_2253,N_19369,N_19676);
nand UO_2254 (O_2254,N_19547,N_19455);
nand UO_2255 (O_2255,N_19313,N_19734);
nand UO_2256 (O_2256,N_19274,N_19215);
or UO_2257 (O_2257,N_19882,N_19805);
nor UO_2258 (O_2258,N_19523,N_19936);
and UO_2259 (O_2259,N_19498,N_19746);
xor UO_2260 (O_2260,N_19733,N_19444);
and UO_2261 (O_2261,N_19345,N_19737);
nand UO_2262 (O_2262,N_19234,N_19964);
or UO_2263 (O_2263,N_19922,N_19678);
nand UO_2264 (O_2264,N_19986,N_19470);
nand UO_2265 (O_2265,N_19318,N_19576);
nand UO_2266 (O_2266,N_19642,N_19516);
or UO_2267 (O_2267,N_19594,N_19960);
nand UO_2268 (O_2268,N_19223,N_19750);
nand UO_2269 (O_2269,N_19990,N_19527);
nor UO_2270 (O_2270,N_19867,N_19326);
xor UO_2271 (O_2271,N_19325,N_19342);
xor UO_2272 (O_2272,N_19909,N_19381);
or UO_2273 (O_2273,N_19970,N_19744);
nor UO_2274 (O_2274,N_19702,N_19579);
or UO_2275 (O_2275,N_19625,N_19394);
nand UO_2276 (O_2276,N_19201,N_19849);
nand UO_2277 (O_2277,N_19936,N_19670);
xnor UO_2278 (O_2278,N_19273,N_19530);
nor UO_2279 (O_2279,N_19326,N_19438);
and UO_2280 (O_2280,N_19668,N_19637);
nand UO_2281 (O_2281,N_19483,N_19297);
xor UO_2282 (O_2282,N_19870,N_19321);
xor UO_2283 (O_2283,N_19208,N_19844);
nand UO_2284 (O_2284,N_19408,N_19203);
nand UO_2285 (O_2285,N_19347,N_19565);
xnor UO_2286 (O_2286,N_19381,N_19941);
or UO_2287 (O_2287,N_19859,N_19623);
nand UO_2288 (O_2288,N_19809,N_19566);
and UO_2289 (O_2289,N_19480,N_19211);
and UO_2290 (O_2290,N_19329,N_19948);
or UO_2291 (O_2291,N_19956,N_19527);
nand UO_2292 (O_2292,N_19307,N_19436);
nor UO_2293 (O_2293,N_19898,N_19267);
nor UO_2294 (O_2294,N_19422,N_19893);
nor UO_2295 (O_2295,N_19913,N_19691);
and UO_2296 (O_2296,N_19432,N_19883);
nor UO_2297 (O_2297,N_19239,N_19410);
or UO_2298 (O_2298,N_19573,N_19267);
nor UO_2299 (O_2299,N_19246,N_19712);
or UO_2300 (O_2300,N_19400,N_19460);
nand UO_2301 (O_2301,N_19306,N_19305);
and UO_2302 (O_2302,N_19606,N_19812);
or UO_2303 (O_2303,N_19667,N_19216);
or UO_2304 (O_2304,N_19867,N_19396);
nand UO_2305 (O_2305,N_19204,N_19839);
and UO_2306 (O_2306,N_19395,N_19769);
or UO_2307 (O_2307,N_19595,N_19737);
nand UO_2308 (O_2308,N_19645,N_19958);
and UO_2309 (O_2309,N_19413,N_19692);
and UO_2310 (O_2310,N_19925,N_19245);
and UO_2311 (O_2311,N_19363,N_19765);
nand UO_2312 (O_2312,N_19672,N_19995);
nand UO_2313 (O_2313,N_19910,N_19271);
nand UO_2314 (O_2314,N_19382,N_19262);
or UO_2315 (O_2315,N_19424,N_19586);
nand UO_2316 (O_2316,N_19341,N_19394);
nand UO_2317 (O_2317,N_19235,N_19354);
nand UO_2318 (O_2318,N_19723,N_19933);
xnor UO_2319 (O_2319,N_19229,N_19597);
or UO_2320 (O_2320,N_19333,N_19348);
nor UO_2321 (O_2321,N_19838,N_19552);
nor UO_2322 (O_2322,N_19421,N_19560);
xnor UO_2323 (O_2323,N_19934,N_19730);
nand UO_2324 (O_2324,N_19427,N_19831);
nand UO_2325 (O_2325,N_19888,N_19289);
nand UO_2326 (O_2326,N_19614,N_19629);
nor UO_2327 (O_2327,N_19515,N_19394);
xor UO_2328 (O_2328,N_19632,N_19494);
nor UO_2329 (O_2329,N_19590,N_19246);
and UO_2330 (O_2330,N_19652,N_19860);
nand UO_2331 (O_2331,N_19608,N_19895);
nor UO_2332 (O_2332,N_19864,N_19522);
and UO_2333 (O_2333,N_19651,N_19835);
or UO_2334 (O_2334,N_19341,N_19223);
nor UO_2335 (O_2335,N_19732,N_19936);
nand UO_2336 (O_2336,N_19806,N_19605);
or UO_2337 (O_2337,N_19777,N_19330);
and UO_2338 (O_2338,N_19735,N_19791);
nand UO_2339 (O_2339,N_19822,N_19281);
xor UO_2340 (O_2340,N_19731,N_19941);
xor UO_2341 (O_2341,N_19797,N_19254);
xor UO_2342 (O_2342,N_19763,N_19643);
and UO_2343 (O_2343,N_19317,N_19542);
nand UO_2344 (O_2344,N_19963,N_19327);
nor UO_2345 (O_2345,N_19399,N_19246);
and UO_2346 (O_2346,N_19228,N_19866);
xor UO_2347 (O_2347,N_19257,N_19337);
or UO_2348 (O_2348,N_19483,N_19828);
and UO_2349 (O_2349,N_19311,N_19473);
nor UO_2350 (O_2350,N_19671,N_19290);
nor UO_2351 (O_2351,N_19497,N_19306);
nor UO_2352 (O_2352,N_19898,N_19457);
xor UO_2353 (O_2353,N_19413,N_19299);
and UO_2354 (O_2354,N_19551,N_19607);
or UO_2355 (O_2355,N_19557,N_19956);
or UO_2356 (O_2356,N_19301,N_19305);
and UO_2357 (O_2357,N_19203,N_19226);
nand UO_2358 (O_2358,N_19748,N_19728);
nand UO_2359 (O_2359,N_19808,N_19731);
nand UO_2360 (O_2360,N_19411,N_19529);
and UO_2361 (O_2361,N_19235,N_19997);
nand UO_2362 (O_2362,N_19634,N_19896);
or UO_2363 (O_2363,N_19368,N_19802);
or UO_2364 (O_2364,N_19596,N_19386);
or UO_2365 (O_2365,N_19506,N_19526);
and UO_2366 (O_2366,N_19450,N_19353);
nand UO_2367 (O_2367,N_19285,N_19613);
and UO_2368 (O_2368,N_19640,N_19638);
and UO_2369 (O_2369,N_19678,N_19875);
xor UO_2370 (O_2370,N_19370,N_19514);
nand UO_2371 (O_2371,N_19333,N_19338);
or UO_2372 (O_2372,N_19783,N_19208);
nand UO_2373 (O_2373,N_19469,N_19703);
nand UO_2374 (O_2374,N_19403,N_19745);
xnor UO_2375 (O_2375,N_19275,N_19842);
xor UO_2376 (O_2376,N_19780,N_19506);
xor UO_2377 (O_2377,N_19835,N_19262);
or UO_2378 (O_2378,N_19602,N_19985);
nand UO_2379 (O_2379,N_19382,N_19980);
xor UO_2380 (O_2380,N_19220,N_19779);
nor UO_2381 (O_2381,N_19933,N_19902);
xnor UO_2382 (O_2382,N_19693,N_19287);
or UO_2383 (O_2383,N_19259,N_19355);
xnor UO_2384 (O_2384,N_19547,N_19889);
nand UO_2385 (O_2385,N_19908,N_19310);
xor UO_2386 (O_2386,N_19823,N_19634);
and UO_2387 (O_2387,N_19794,N_19689);
or UO_2388 (O_2388,N_19379,N_19799);
nand UO_2389 (O_2389,N_19577,N_19346);
nand UO_2390 (O_2390,N_19606,N_19871);
and UO_2391 (O_2391,N_19498,N_19893);
nor UO_2392 (O_2392,N_19958,N_19613);
or UO_2393 (O_2393,N_19267,N_19293);
or UO_2394 (O_2394,N_19499,N_19701);
nor UO_2395 (O_2395,N_19833,N_19805);
nor UO_2396 (O_2396,N_19728,N_19674);
and UO_2397 (O_2397,N_19849,N_19624);
nand UO_2398 (O_2398,N_19786,N_19546);
nand UO_2399 (O_2399,N_19947,N_19474);
or UO_2400 (O_2400,N_19697,N_19374);
or UO_2401 (O_2401,N_19532,N_19682);
nand UO_2402 (O_2402,N_19951,N_19413);
nand UO_2403 (O_2403,N_19676,N_19393);
xnor UO_2404 (O_2404,N_19543,N_19390);
nand UO_2405 (O_2405,N_19463,N_19232);
xnor UO_2406 (O_2406,N_19504,N_19683);
xnor UO_2407 (O_2407,N_19433,N_19807);
or UO_2408 (O_2408,N_19916,N_19734);
xnor UO_2409 (O_2409,N_19526,N_19319);
or UO_2410 (O_2410,N_19840,N_19858);
or UO_2411 (O_2411,N_19721,N_19808);
xor UO_2412 (O_2412,N_19969,N_19652);
xnor UO_2413 (O_2413,N_19754,N_19214);
and UO_2414 (O_2414,N_19363,N_19224);
or UO_2415 (O_2415,N_19383,N_19258);
nor UO_2416 (O_2416,N_19398,N_19540);
or UO_2417 (O_2417,N_19676,N_19919);
xnor UO_2418 (O_2418,N_19942,N_19224);
nand UO_2419 (O_2419,N_19631,N_19237);
and UO_2420 (O_2420,N_19879,N_19881);
or UO_2421 (O_2421,N_19962,N_19636);
or UO_2422 (O_2422,N_19303,N_19669);
nand UO_2423 (O_2423,N_19298,N_19602);
and UO_2424 (O_2424,N_19998,N_19417);
nand UO_2425 (O_2425,N_19229,N_19763);
or UO_2426 (O_2426,N_19800,N_19654);
nand UO_2427 (O_2427,N_19295,N_19851);
nor UO_2428 (O_2428,N_19260,N_19966);
and UO_2429 (O_2429,N_19710,N_19342);
or UO_2430 (O_2430,N_19333,N_19422);
or UO_2431 (O_2431,N_19889,N_19721);
nand UO_2432 (O_2432,N_19221,N_19760);
nor UO_2433 (O_2433,N_19407,N_19774);
xor UO_2434 (O_2434,N_19302,N_19941);
xnor UO_2435 (O_2435,N_19394,N_19666);
nor UO_2436 (O_2436,N_19509,N_19698);
nand UO_2437 (O_2437,N_19385,N_19887);
nor UO_2438 (O_2438,N_19861,N_19488);
or UO_2439 (O_2439,N_19397,N_19834);
xnor UO_2440 (O_2440,N_19244,N_19288);
nor UO_2441 (O_2441,N_19633,N_19305);
and UO_2442 (O_2442,N_19782,N_19404);
xor UO_2443 (O_2443,N_19315,N_19695);
nand UO_2444 (O_2444,N_19972,N_19552);
and UO_2445 (O_2445,N_19850,N_19984);
or UO_2446 (O_2446,N_19246,N_19427);
xnor UO_2447 (O_2447,N_19247,N_19478);
xor UO_2448 (O_2448,N_19478,N_19702);
nand UO_2449 (O_2449,N_19926,N_19609);
or UO_2450 (O_2450,N_19689,N_19946);
and UO_2451 (O_2451,N_19591,N_19668);
nand UO_2452 (O_2452,N_19679,N_19730);
or UO_2453 (O_2453,N_19311,N_19414);
nand UO_2454 (O_2454,N_19255,N_19631);
nand UO_2455 (O_2455,N_19925,N_19731);
nor UO_2456 (O_2456,N_19923,N_19410);
nor UO_2457 (O_2457,N_19246,N_19487);
xor UO_2458 (O_2458,N_19345,N_19843);
nor UO_2459 (O_2459,N_19228,N_19230);
xnor UO_2460 (O_2460,N_19771,N_19574);
and UO_2461 (O_2461,N_19894,N_19460);
nor UO_2462 (O_2462,N_19432,N_19610);
xor UO_2463 (O_2463,N_19351,N_19735);
and UO_2464 (O_2464,N_19275,N_19633);
or UO_2465 (O_2465,N_19561,N_19906);
nor UO_2466 (O_2466,N_19274,N_19716);
or UO_2467 (O_2467,N_19474,N_19869);
and UO_2468 (O_2468,N_19412,N_19567);
nand UO_2469 (O_2469,N_19451,N_19429);
nand UO_2470 (O_2470,N_19634,N_19726);
and UO_2471 (O_2471,N_19548,N_19741);
and UO_2472 (O_2472,N_19822,N_19395);
or UO_2473 (O_2473,N_19698,N_19592);
nand UO_2474 (O_2474,N_19781,N_19879);
nor UO_2475 (O_2475,N_19838,N_19874);
nand UO_2476 (O_2476,N_19691,N_19888);
nand UO_2477 (O_2477,N_19268,N_19417);
xnor UO_2478 (O_2478,N_19345,N_19366);
nor UO_2479 (O_2479,N_19295,N_19262);
or UO_2480 (O_2480,N_19350,N_19731);
or UO_2481 (O_2481,N_19231,N_19711);
and UO_2482 (O_2482,N_19310,N_19730);
nor UO_2483 (O_2483,N_19689,N_19848);
or UO_2484 (O_2484,N_19931,N_19780);
xnor UO_2485 (O_2485,N_19870,N_19564);
or UO_2486 (O_2486,N_19782,N_19549);
xor UO_2487 (O_2487,N_19745,N_19530);
nor UO_2488 (O_2488,N_19516,N_19634);
or UO_2489 (O_2489,N_19362,N_19434);
xor UO_2490 (O_2490,N_19972,N_19524);
nor UO_2491 (O_2491,N_19655,N_19626);
nor UO_2492 (O_2492,N_19723,N_19784);
nand UO_2493 (O_2493,N_19285,N_19914);
and UO_2494 (O_2494,N_19362,N_19715);
or UO_2495 (O_2495,N_19287,N_19789);
nand UO_2496 (O_2496,N_19363,N_19981);
nor UO_2497 (O_2497,N_19610,N_19462);
nand UO_2498 (O_2498,N_19729,N_19697);
nor UO_2499 (O_2499,N_19721,N_19454);
endmodule