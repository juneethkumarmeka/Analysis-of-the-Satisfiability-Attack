module basic_500_3000_500_30_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_289,In_315);
nor U1 (N_1,In_425,In_367);
and U2 (N_2,In_160,In_346);
or U3 (N_3,In_209,In_230);
or U4 (N_4,In_228,In_11);
or U5 (N_5,In_214,In_396);
or U6 (N_6,In_181,In_254);
nand U7 (N_7,In_222,In_47);
nor U8 (N_8,In_395,In_393);
or U9 (N_9,In_342,In_296);
nand U10 (N_10,In_18,In_251);
and U11 (N_11,In_198,In_167);
nand U12 (N_12,In_320,In_57);
and U13 (N_13,In_2,In_80);
nand U14 (N_14,In_485,In_443);
nor U15 (N_15,In_187,In_460);
nand U16 (N_16,In_362,In_189);
and U17 (N_17,In_233,In_34);
or U18 (N_18,In_406,In_133);
and U19 (N_19,In_441,In_308);
or U20 (N_20,In_39,In_434);
and U21 (N_21,In_426,In_468);
or U22 (N_22,In_427,In_288);
and U23 (N_23,In_445,In_72);
nand U24 (N_24,In_210,In_50);
nand U25 (N_25,In_405,In_201);
and U26 (N_26,In_202,In_299);
nand U27 (N_27,In_484,In_217);
nor U28 (N_28,In_136,In_118);
and U29 (N_29,In_370,In_5);
and U30 (N_30,In_90,In_175);
nand U31 (N_31,In_389,In_9);
or U32 (N_32,In_52,In_205);
nand U33 (N_33,In_411,In_446);
or U34 (N_34,In_237,In_125);
nor U35 (N_35,In_221,In_65);
nor U36 (N_36,In_302,In_323);
and U37 (N_37,In_357,In_195);
or U38 (N_38,In_190,In_131);
nand U39 (N_39,In_374,In_25);
or U40 (N_40,In_339,In_74);
and U41 (N_41,In_345,In_83);
nand U42 (N_42,In_23,In_36);
or U43 (N_43,In_191,In_193);
nand U44 (N_44,In_338,In_212);
nand U45 (N_45,In_303,In_22);
or U46 (N_46,In_277,In_482);
nand U47 (N_47,In_317,In_192);
nor U48 (N_48,In_135,In_358);
or U49 (N_49,In_111,In_140);
nand U50 (N_50,In_282,In_264);
nand U51 (N_51,In_248,In_69);
and U52 (N_52,In_499,In_404);
and U53 (N_53,In_120,In_351);
nor U54 (N_54,In_142,In_32);
and U55 (N_55,In_223,In_84);
nand U56 (N_56,In_108,In_143);
nor U57 (N_57,In_3,In_477);
and U58 (N_58,In_487,In_206);
or U59 (N_59,In_44,In_494);
nand U60 (N_60,In_4,In_10);
nor U61 (N_61,In_227,In_493);
and U62 (N_62,In_162,In_98);
nor U63 (N_63,In_438,In_124);
xnor U64 (N_64,In_461,In_319);
nand U65 (N_65,In_163,In_376);
nor U66 (N_66,In_380,In_82);
or U67 (N_67,In_188,In_349);
and U68 (N_68,In_259,In_271);
nand U69 (N_69,In_153,In_306);
or U70 (N_70,In_15,In_348);
nor U71 (N_71,In_197,In_244);
nand U72 (N_72,In_99,In_149);
nand U73 (N_73,In_56,In_86);
and U74 (N_74,In_75,In_126);
nand U75 (N_75,In_311,In_401);
nor U76 (N_76,In_437,In_343);
nand U77 (N_77,In_378,In_298);
nor U78 (N_78,In_260,In_177);
or U79 (N_79,In_454,In_114);
and U80 (N_80,In_43,In_421);
xor U81 (N_81,In_322,In_449);
nand U82 (N_82,In_440,In_46);
and U83 (N_83,In_372,In_49);
nor U84 (N_84,In_356,In_444);
or U85 (N_85,In_20,In_176);
nand U86 (N_86,In_469,In_432);
nand U87 (N_87,In_331,In_375);
nor U88 (N_88,In_88,In_159);
nand U89 (N_89,In_157,In_414);
and U90 (N_90,In_337,In_392);
and U91 (N_91,In_60,In_495);
and U92 (N_92,In_285,In_424);
or U93 (N_93,In_16,In_387);
and U94 (N_94,In_294,In_341);
or U95 (N_95,In_247,In_253);
nand U96 (N_96,In_292,In_168);
and U97 (N_97,In_498,In_194);
or U98 (N_98,In_450,In_249);
nor U99 (N_99,In_101,In_266);
nand U100 (N_100,In_369,In_78);
nor U101 (N_101,In_272,In_310);
nand U102 (N_102,In_408,In_107);
and U103 (N_103,In_238,In_184);
and U104 (N_104,N_71,In_474);
or U105 (N_105,In_382,In_324);
or U106 (N_106,N_0,In_430);
or U107 (N_107,In_256,In_458);
or U108 (N_108,N_40,In_179);
and U109 (N_109,In_95,In_200);
nand U110 (N_110,In_312,In_154);
or U111 (N_111,N_98,In_383);
and U112 (N_112,N_70,N_44);
or U113 (N_113,In_258,In_123);
nand U114 (N_114,N_39,In_27);
and U115 (N_115,In_475,In_470);
and U116 (N_116,In_270,N_51);
nand U117 (N_117,In_229,N_91);
or U118 (N_118,In_412,N_14);
or U119 (N_119,N_37,In_19);
and U120 (N_120,In_486,In_496);
nand U121 (N_121,In_129,In_483);
xor U122 (N_122,In_66,In_488);
nand U123 (N_123,N_10,In_59);
and U124 (N_124,In_436,In_145);
nor U125 (N_125,In_330,In_419);
or U126 (N_126,In_472,In_284);
nor U127 (N_127,In_431,In_459);
nor U128 (N_128,In_365,N_8);
nand U129 (N_129,In_155,N_62);
nand U130 (N_130,In_17,N_42);
nor U131 (N_131,In_232,N_66);
or U132 (N_132,In_373,N_52);
nand U133 (N_133,In_0,In_106);
nor U134 (N_134,In_327,In_185);
and U135 (N_135,In_26,In_161);
nor U136 (N_136,N_13,In_381);
nor U137 (N_137,In_473,N_65);
nor U138 (N_138,N_58,In_301);
or U139 (N_139,In_169,In_335);
nand U140 (N_140,N_77,In_418);
and U141 (N_141,In_433,In_61);
and U142 (N_142,In_55,N_83);
or U143 (N_143,In_79,In_64);
and U144 (N_144,In_203,In_326);
nor U145 (N_145,N_86,N_96);
and U146 (N_146,In_278,In_141);
nor U147 (N_147,In_417,N_34);
nor U148 (N_148,In_220,In_307);
and U149 (N_149,In_213,N_68);
and U150 (N_150,In_252,N_28);
and U151 (N_151,In_150,In_313);
nand U152 (N_152,In_239,In_448);
nor U153 (N_153,In_267,N_49);
or U154 (N_154,In_216,In_37);
nor U155 (N_155,N_1,In_235);
and U156 (N_156,In_489,N_76);
nor U157 (N_157,In_388,N_97);
or U158 (N_158,N_59,In_127);
and U159 (N_159,N_79,N_78);
nand U160 (N_160,In_132,In_96);
or U161 (N_161,N_85,In_110);
and U162 (N_162,N_11,In_407);
nor U163 (N_163,N_82,In_68);
or U164 (N_164,In_172,N_12);
or U165 (N_165,In_347,In_109);
nand U166 (N_166,In_415,N_29);
or U167 (N_167,N_5,In_451);
nand U168 (N_168,In_263,In_447);
nor U169 (N_169,In_314,In_226);
and U170 (N_170,In_462,In_104);
nor U171 (N_171,N_99,In_280);
nand U172 (N_172,In_379,N_74);
or U173 (N_173,In_148,In_164);
nand U174 (N_174,In_384,In_97);
nand U175 (N_175,In_138,In_340);
and U176 (N_176,In_453,In_279);
nor U177 (N_177,In_71,In_144);
or U178 (N_178,In_147,In_245);
or U179 (N_179,N_19,In_14);
nor U180 (N_180,In_146,N_87);
and U181 (N_181,In_268,In_265);
nor U182 (N_182,N_7,N_41);
and U183 (N_183,In_410,N_38);
nand U184 (N_184,In_40,In_361);
nand U185 (N_185,In_478,In_309);
or U186 (N_186,In_178,In_492);
or U187 (N_187,In_35,N_30);
or U188 (N_188,In_87,N_61);
xor U189 (N_189,In_416,In_183);
and U190 (N_190,In_385,In_219);
or U191 (N_191,In_397,In_275);
or U192 (N_192,In_171,In_355);
nand U193 (N_193,N_17,N_43);
and U194 (N_194,N_64,In_42);
nand U195 (N_195,In_180,In_479);
nand U196 (N_196,In_152,In_121);
or U197 (N_197,In_439,N_56);
and U198 (N_198,In_48,In_332);
or U199 (N_199,N_4,N_18);
or U200 (N_200,In_300,In_134);
or U201 (N_201,N_105,In_352);
or U202 (N_202,In_41,In_413);
or U203 (N_203,In_452,In_409);
and U204 (N_204,N_138,In_466);
and U205 (N_205,In_103,N_157);
nor U206 (N_206,N_69,In_390);
nor U207 (N_207,N_131,In_386);
or U208 (N_208,In_6,N_125);
or U209 (N_209,In_208,In_63);
and U210 (N_210,N_80,N_2);
nor U211 (N_211,In_45,N_166);
nand U212 (N_212,In_242,N_147);
or U213 (N_213,In_112,In_476);
or U214 (N_214,N_93,In_286);
nor U215 (N_215,N_104,In_257);
or U216 (N_216,N_159,N_45);
or U217 (N_217,N_109,In_28);
nor U218 (N_218,N_150,In_255);
and U219 (N_219,In_81,In_243);
and U220 (N_220,In_305,In_480);
or U221 (N_221,In_38,In_139);
nor U222 (N_222,N_46,N_170);
nor U223 (N_223,In_295,N_15);
or U224 (N_224,In_359,In_102);
and U225 (N_225,In_224,N_180);
nand U226 (N_226,N_156,In_457);
or U227 (N_227,N_55,In_70);
and U228 (N_228,N_22,N_186);
and U229 (N_229,N_95,In_353);
or U230 (N_230,In_465,N_57);
nand U231 (N_231,N_126,N_176);
nand U232 (N_232,In_354,In_471);
nand U233 (N_233,In_119,N_161);
nand U234 (N_234,N_172,N_142);
nor U235 (N_235,N_169,In_368);
and U236 (N_236,N_165,In_261);
and U237 (N_237,N_31,N_73);
nand U238 (N_238,In_497,In_360);
nor U239 (N_239,In_394,In_321);
nand U240 (N_240,In_105,In_423);
or U241 (N_241,N_9,N_146);
nand U242 (N_242,In_186,N_128);
or U243 (N_243,N_196,N_132);
nand U244 (N_244,N_48,In_122);
nand U245 (N_245,N_181,N_179);
or U246 (N_246,In_269,N_103);
or U247 (N_247,N_152,N_120);
nor U248 (N_248,N_116,N_107);
nor U249 (N_249,In_377,In_73);
and U250 (N_250,N_88,N_158);
nand U251 (N_251,In_92,In_246);
and U252 (N_252,In_350,In_91);
nor U253 (N_253,In_117,In_218);
nor U254 (N_254,In_293,N_193);
nand U255 (N_255,In_51,N_119);
nor U256 (N_256,N_81,In_371);
or U257 (N_257,N_189,N_27);
or U258 (N_258,N_185,N_24);
and U259 (N_259,N_53,N_101);
nand U260 (N_260,N_127,N_25);
and U261 (N_261,N_26,In_344);
or U262 (N_262,In_199,In_165);
or U263 (N_263,N_198,In_403);
and U264 (N_264,N_195,N_182);
or U265 (N_265,N_188,In_54);
or U266 (N_266,N_151,In_273);
and U267 (N_267,In_170,In_29);
or U268 (N_268,N_113,In_336);
or U269 (N_269,N_144,N_133);
nor U270 (N_270,N_187,In_116);
or U271 (N_271,N_102,N_177);
and U272 (N_272,In_234,N_197);
nor U273 (N_273,In_420,In_467);
nor U274 (N_274,In_128,N_106);
or U275 (N_275,N_178,In_33);
or U276 (N_276,In_196,In_363);
nor U277 (N_277,N_145,N_111);
nand U278 (N_278,In_283,N_121);
nand U279 (N_279,In_262,N_23);
nand U280 (N_280,In_62,In_429);
nand U281 (N_281,N_89,In_281);
nand U282 (N_282,In_481,In_402);
and U283 (N_283,N_153,In_156);
or U284 (N_284,In_366,In_290);
and U285 (N_285,In_93,N_160);
or U286 (N_286,N_194,N_190);
and U287 (N_287,In_276,In_100);
and U288 (N_288,In_334,N_140);
or U289 (N_289,In_204,N_16);
and U290 (N_290,In_364,In_8);
or U291 (N_291,N_50,N_141);
nand U292 (N_292,In_58,In_236);
nand U293 (N_293,In_463,N_191);
nor U294 (N_294,N_199,N_33);
and U295 (N_295,N_94,N_32);
nand U296 (N_296,In_391,In_85);
or U297 (N_297,N_174,N_92);
nor U298 (N_298,In_287,N_175);
nand U299 (N_299,N_154,In_115);
and U300 (N_300,In_215,N_21);
nor U301 (N_301,N_275,In_12);
or U302 (N_302,N_235,In_398);
or U303 (N_303,N_279,N_136);
or U304 (N_304,N_84,N_212);
or U305 (N_305,N_122,In_94);
nand U306 (N_306,In_7,N_243);
nor U307 (N_307,N_238,N_232);
and U308 (N_308,N_293,N_265);
nand U309 (N_309,N_6,In_13);
nand U310 (N_310,N_90,N_255);
or U311 (N_311,N_236,N_163);
nand U312 (N_312,N_134,N_281);
nand U313 (N_313,N_272,N_219);
or U314 (N_314,N_224,N_202);
and U315 (N_315,N_268,N_237);
or U316 (N_316,N_227,In_464);
nand U317 (N_317,In_399,N_183);
nand U318 (N_318,In_1,N_210);
and U319 (N_319,In_325,N_143);
xor U320 (N_320,In_422,N_278);
nor U321 (N_321,In_31,In_318);
nand U322 (N_322,In_428,In_89);
nand U323 (N_323,N_3,In_76);
nor U324 (N_324,In_211,N_296);
or U325 (N_325,In_240,In_231);
nand U326 (N_326,N_283,In_442);
or U327 (N_327,N_256,N_110);
and U328 (N_328,In_113,N_297);
nor U329 (N_329,N_290,N_205);
nand U330 (N_330,N_241,N_253);
and U331 (N_331,In_491,In_456);
nand U332 (N_332,N_245,N_167);
nand U333 (N_333,N_288,N_207);
nor U334 (N_334,N_47,N_260);
nor U335 (N_335,N_287,N_206);
nand U336 (N_336,N_266,N_229);
or U337 (N_337,N_289,In_158);
nand U338 (N_338,N_75,In_53);
nor U339 (N_339,In_304,N_223);
nand U340 (N_340,N_271,N_130);
and U341 (N_341,In_182,N_100);
nand U342 (N_342,N_252,N_221);
nand U343 (N_343,N_216,N_123);
nand U344 (N_344,In_21,N_226);
nor U345 (N_345,N_251,In_291);
and U346 (N_346,N_214,N_67);
and U347 (N_347,N_263,N_264);
nand U348 (N_348,N_164,In_250);
and U349 (N_349,In_151,N_108);
and U350 (N_350,N_276,N_269);
and U351 (N_351,N_171,N_112);
or U352 (N_352,In_207,N_209);
or U353 (N_353,N_204,N_135);
and U354 (N_354,N_148,N_213);
and U355 (N_355,N_250,N_220);
nand U356 (N_356,N_270,N_162);
and U357 (N_357,N_114,In_328);
nand U358 (N_358,N_184,In_316);
nand U359 (N_359,N_201,N_240);
nor U360 (N_360,N_203,In_455);
nor U361 (N_361,N_248,N_242);
nand U362 (N_362,In_435,In_490);
and U363 (N_363,N_234,N_254);
or U364 (N_364,N_60,In_174);
nor U365 (N_365,N_139,In_225);
nor U366 (N_366,N_282,In_30);
or U367 (N_367,In_241,N_292);
nand U368 (N_368,N_267,N_222);
nand U369 (N_369,N_230,In_333);
nor U370 (N_370,N_208,N_280);
or U371 (N_371,N_259,N_217);
and U372 (N_372,N_218,N_261);
nor U373 (N_373,N_291,N_249);
nor U374 (N_374,N_35,N_118);
or U375 (N_375,N_129,N_117);
or U376 (N_376,In_329,N_137);
nor U377 (N_377,In_24,In_137);
nor U378 (N_378,In_274,N_273);
and U379 (N_379,N_244,N_36);
or U380 (N_380,N_200,In_166);
or U381 (N_381,N_63,N_115);
nand U382 (N_382,N_211,In_297);
or U383 (N_383,N_277,In_173);
and U384 (N_384,N_168,N_298);
and U385 (N_385,N_247,N_149);
nor U386 (N_386,N_155,N_231);
nor U387 (N_387,N_257,N_294);
nor U388 (N_388,N_228,N_72);
and U389 (N_389,N_173,N_215);
nand U390 (N_390,N_20,N_262);
and U391 (N_391,In_77,N_124);
nor U392 (N_392,N_286,In_67);
and U393 (N_393,N_192,N_239);
nand U394 (N_394,N_233,N_246);
nor U395 (N_395,N_258,N_284);
nand U396 (N_396,N_299,N_274);
and U397 (N_397,In_400,N_295);
and U398 (N_398,In_130,N_285);
and U399 (N_399,N_225,N_54);
and U400 (N_400,N_316,N_348);
nor U401 (N_401,N_373,N_353);
nand U402 (N_402,N_309,N_378);
or U403 (N_403,N_356,N_349);
or U404 (N_404,N_352,N_385);
nand U405 (N_405,N_359,N_389);
or U406 (N_406,N_360,N_321);
nor U407 (N_407,N_336,N_350);
and U408 (N_408,N_342,N_397);
nand U409 (N_409,N_323,N_375);
or U410 (N_410,N_333,N_383);
xnor U411 (N_411,N_366,N_335);
and U412 (N_412,N_364,N_395);
nor U413 (N_413,N_393,N_345);
nor U414 (N_414,N_367,N_399);
or U415 (N_415,N_315,N_310);
nand U416 (N_416,N_390,N_392);
and U417 (N_417,N_384,N_379);
and U418 (N_418,N_330,N_371);
nor U419 (N_419,N_329,N_320);
nand U420 (N_420,N_362,N_365);
nor U421 (N_421,N_388,N_340);
nor U422 (N_422,N_341,N_377);
and U423 (N_423,N_338,N_368);
and U424 (N_424,N_347,N_318);
or U425 (N_425,N_358,N_387);
and U426 (N_426,N_357,N_331);
or U427 (N_427,N_381,N_391);
nand U428 (N_428,N_325,N_317);
nor U429 (N_429,N_306,N_369);
and U430 (N_430,N_319,N_361);
nor U431 (N_431,N_355,N_372);
nand U432 (N_432,N_370,N_334);
or U433 (N_433,N_302,N_314);
and U434 (N_434,N_346,N_396);
or U435 (N_435,N_398,N_324);
and U436 (N_436,N_351,N_363);
and U437 (N_437,N_328,N_326);
and U438 (N_438,N_374,N_305);
or U439 (N_439,N_300,N_303);
and U440 (N_440,N_386,N_307);
or U441 (N_441,N_337,N_354);
nand U442 (N_442,N_327,N_382);
and U443 (N_443,N_376,N_311);
nand U444 (N_444,N_344,N_313);
nor U445 (N_445,N_312,N_380);
and U446 (N_446,N_304,N_339);
nand U447 (N_447,N_332,N_343);
nor U448 (N_448,N_322,N_394);
or U449 (N_449,N_301,N_308);
nand U450 (N_450,N_399,N_392);
or U451 (N_451,N_340,N_333);
or U452 (N_452,N_384,N_339);
nor U453 (N_453,N_366,N_399);
and U454 (N_454,N_340,N_391);
nand U455 (N_455,N_308,N_303);
or U456 (N_456,N_395,N_308);
nand U457 (N_457,N_377,N_384);
nand U458 (N_458,N_322,N_377);
or U459 (N_459,N_398,N_389);
nor U460 (N_460,N_360,N_362);
and U461 (N_461,N_384,N_320);
xor U462 (N_462,N_350,N_332);
and U463 (N_463,N_371,N_352);
or U464 (N_464,N_389,N_336);
nor U465 (N_465,N_399,N_328);
and U466 (N_466,N_347,N_353);
and U467 (N_467,N_360,N_378);
and U468 (N_468,N_349,N_327);
or U469 (N_469,N_390,N_361);
nor U470 (N_470,N_393,N_339);
and U471 (N_471,N_340,N_387);
or U472 (N_472,N_345,N_396);
or U473 (N_473,N_303,N_389);
and U474 (N_474,N_309,N_383);
xor U475 (N_475,N_346,N_312);
nand U476 (N_476,N_345,N_349);
and U477 (N_477,N_366,N_393);
or U478 (N_478,N_358,N_397);
nand U479 (N_479,N_354,N_380);
and U480 (N_480,N_358,N_344);
or U481 (N_481,N_339,N_320);
nand U482 (N_482,N_379,N_335);
nand U483 (N_483,N_378,N_346);
or U484 (N_484,N_375,N_394);
or U485 (N_485,N_396,N_334);
nor U486 (N_486,N_340,N_347);
or U487 (N_487,N_385,N_391);
and U488 (N_488,N_347,N_386);
nor U489 (N_489,N_394,N_317);
nand U490 (N_490,N_357,N_324);
or U491 (N_491,N_375,N_333);
and U492 (N_492,N_339,N_335);
nand U493 (N_493,N_391,N_326);
nand U494 (N_494,N_311,N_324);
nand U495 (N_495,N_318,N_369);
nor U496 (N_496,N_337,N_318);
nand U497 (N_497,N_372,N_398);
nor U498 (N_498,N_367,N_343);
nand U499 (N_499,N_325,N_359);
and U500 (N_500,N_473,N_417);
nor U501 (N_501,N_481,N_411);
nor U502 (N_502,N_459,N_490);
xnor U503 (N_503,N_453,N_458);
xor U504 (N_504,N_404,N_493);
and U505 (N_505,N_487,N_491);
or U506 (N_506,N_433,N_418);
and U507 (N_507,N_401,N_451);
and U508 (N_508,N_450,N_470);
nand U509 (N_509,N_494,N_436);
nand U510 (N_510,N_438,N_441);
or U511 (N_511,N_456,N_443);
and U512 (N_512,N_403,N_449);
or U513 (N_513,N_448,N_416);
nor U514 (N_514,N_496,N_474);
nor U515 (N_515,N_483,N_402);
and U516 (N_516,N_432,N_471);
and U517 (N_517,N_414,N_425);
nand U518 (N_518,N_424,N_455);
nor U519 (N_519,N_465,N_434);
nor U520 (N_520,N_407,N_460);
nand U521 (N_521,N_408,N_454);
and U522 (N_522,N_498,N_480);
nand U523 (N_523,N_400,N_415);
and U524 (N_524,N_423,N_440);
nor U525 (N_525,N_413,N_477);
xor U526 (N_526,N_463,N_478);
or U527 (N_527,N_497,N_447);
nor U528 (N_528,N_462,N_428);
and U529 (N_529,N_469,N_461);
nand U530 (N_530,N_482,N_486);
nand U531 (N_531,N_452,N_442);
and U532 (N_532,N_475,N_405);
and U533 (N_533,N_410,N_406);
nand U534 (N_534,N_489,N_437);
nor U535 (N_535,N_430,N_468);
and U536 (N_536,N_495,N_431);
nor U537 (N_537,N_467,N_464);
nand U538 (N_538,N_445,N_485);
or U539 (N_539,N_476,N_492);
nand U540 (N_540,N_422,N_499);
nand U541 (N_541,N_446,N_419);
nand U542 (N_542,N_427,N_479);
and U543 (N_543,N_412,N_421);
and U544 (N_544,N_488,N_426);
or U545 (N_545,N_435,N_409);
and U546 (N_546,N_439,N_466);
nor U547 (N_547,N_429,N_484);
or U548 (N_548,N_472,N_457);
nand U549 (N_549,N_444,N_420);
nor U550 (N_550,N_410,N_411);
nor U551 (N_551,N_425,N_434);
and U552 (N_552,N_480,N_472);
and U553 (N_553,N_422,N_400);
nand U554 (N_554,N_479,N_461);
and U555 (N_555,N_426,N_410);
xor U556 (N_556,N_413,N_456);
nand U557 (N_557,N_454,N_433);
nor U558 (N_558,N_491,N_495);
nor U559 (N_559,N_444,N_419);
and U560 (N_560,N_421,N_495);
and U561 (N_561,N_452,N_468);
and U562 (N_562,N_438,N_496);
or U563 (N_563,N_499,N_444);
nand U564 (N_564,N_420,N_411);
or U565 (N_565,N_483,N_446);
and U566 (N_566,N_460,N_492);
and U567 (N_567,N_493,N_497);
nor U568 (N_568,N_480,N_495);
or U569 (N_569,N_410,N_448);
nand U570 (N_570,N_480,N_487);
and U571 (N_571,N_405,N_480);
nand U572 (N_572,N_468,N_417);
nor U573 (N_573,N_451,N_417);
and U574 (N_574,N_491,N_410);
or U575 (N_575,N_492,N_481);
or U576 (N_576,N_483,N_468);
nor U577 (N_577,N_407,N_483);
nand U578 (N_578,N_402,N_481);
nor U579 (N_579,N_410,N_465);
and U580 (N_580,N_480,N_400);
or U581 (N_581,N_437,N_431);
or U582 (N_582,N_427,N_404);
and U583 (N_583,N_433,N_402);
and U584 (N_584,N_486,N_468);
and U585 (N_585,N_475,N_433);
nor U586 (N_586,N_461,N_439);
and U587 (N_587,N_491,N_494);
and U588 (N_588,N_427,N_499);
nand U589 (N_589,N_473,N_452);
and U590 (N_590,N_410,N_422);
nor U591 (N_591,N_437,N_469);
and U592 (N_592,N_456,N_455);
and U593 (N_593,N_498,N_471);
nand U594 (N_594,N_464,N_422);
nor U595 (N_595,N_449,N_408);
and U596 (N_596,N_440,N_434);
nand U597 (N_597,N_451,N_408);
nor U598 (N_598,N_477,N_469);
and U599 (N_599,N_490,N_454);
and U600 (N_600,N_517,N_558);
or U601 (N_601,N_544,N_542);
or U602 (N_602,N_557,N_548);
nor U603 (N_603,N_589,N_578);
and U604 (N_604,N_599,N_556);
and U605 (N_605,N_511,N_519);
or U606 (N_606,N_592,N_567);
nor U607 (N_607,N_560,N_561);
or U608 (N_608,N_528,N_510);
or U609 (N_609,N_541,N_587);
or U610 (N_610,N_506,N_573);
and U611 (N_611,N_520,N_574);
or U612 (N_612,N_543,N_547);
nor U613 (N_613,N_593,N_572);
nand U614 (N_614,N_531,N_563);
and U615 (N_615,N_545,N_550);
nor U616 (N_616,N_504,N_529);
and U617 (N_617,N_562,N_507);
nand U618 (N_618,N_530,N_516);
nor U619 (N_619,N_584,N_554);
nor U620 (N_620,N_539,N_534);
nand U621 (N_621,N_570,N_582);
nor U622 (N_622,N_586,N_590);
nor U623 (N_623,N_526,N_597);
nand U624 (N_624,N_552,N_555);
nor U625 (N_625,N_591,N_537);
and U626 (N_626,N_564,N_515);
nand U627 (N_627,N_525,N_522);
and U628 (N_628,N_596,N_553);
and U629 (N_629,N_551,N_514);
and U630 (N_630,N_518,N_508);
or U631 (N_631,N_594,N_533);
or U632 (N_632,N_568,N_540);
or U633 (N_633,N_538,N_503);
and U634 (N_634,N_581,N_559);
nand U635 (N_635,N_583,N_512);
nand U636 (N_636,N_588,N_509);
and U637 (N_637,N_569,N_576);
nor U638 (N_638,N_598,N_500);
nor U639 (N_639,N_549,N_513);
nand U640 (N_640,N_501,N_523);
nand U641 (N_641,N_524,N_535);
and U642 (N_642,N_580,N_546);
and U643 (N_643,N_585,N_566);
or U644 (N_644,N_536,N_565);
and U645 (N_645,N_521,N_527);
or U646 (N_646,N_577,N_532);
or U647 (N_647,N_575,N_595);
nor U648 (N_648,N_571,N_505);
and U649 (N_649,N_579,N_502);
and U650 (N_650,N_571,N_565);
or U651 (N_651,N_506,N_551);
nor U652 (N_652,N_595,N_527);
nor U653 (N_653,N_598,N_543);
and U654 (N_654,N_520,N_549);
nand U655 (N_655,N_538,N_532);
or U656 (N_656,N_575,N_512);
and U657 (N_657,N_570,N_572);
and U658 (N_658,N_539,N_531);
or U659 (N_659,N_557,N_567);
and U660 (N_660,N_534,N_504);
and U661 (N_661,N_503,N_554);
nand U662 (N_662,N_520,N_578);
nor U663 (N_663,N_510,N_511);
nor U664 (N_664,N_580,N_562);
nand U665 (N_665,N_521,N_506);
and U666 (N_666,N_570,N_566);
nand U667 (N_667,N_547,N_519);
nand U668 (N_668,N_557,N_581);
nand U669 (N_669,N_546,N_500);
nand U670 (N_670,N_562,N_547);
and U671 (N_671,N_585,N_598);
nor U672 (N_672,N_538,N_505);
or U673 (N_673,N_591,N_516);
nand U674 (N_674,N_596,N_577);
xnor U675 (N_675,N_514,N_537);
or U676 (N_676,N_574,N_579);
nor U677 (N_677,N_516,N_528);
nor U678 (N_678,N_596,N_551);
xor U679 (N_679,N_513,N_514);
or U680 (N_680,N_599,N_530);
and U681 (N_681,N_580,N_592);
nor U682 (N_682,N_530,N_569);
nor U683 (N_683,N_571,N_541);
xnor U684 (N_684,N_566,N_525);
nor U685 (N_685,N_554,N_578);
nor U686 (N_686,N_521,N_505);
nand U687 (N_687,N_550,N_592);
or U688 (N_688,N_513,N_563);
or U689 (N_689,N_530,N_584);
or U690 (N_690,N_557,N_518);
nand U691 (N_691,N_596,N_534);
nand U692 (N_692,N_595,N_505);
and U693 (N_693,N_553,N_537);
nand U694 (N_694,N_559,N_507);
nand U695 (N_695,N_503,N_546);
or U696 (N_696,N_576,N_591);
or U697 (N_697,N_548,N_572);
nand U698 (N_698,N_545,N_561);
nand U699 (N_699,N_577,N_598);
and U700 (N_700,N_683,N_692);
or U701 (N_701,N_670,N_629);
nand U702 (N_702,N_614,N_665);
or U703 (N_703,N_676,N_600);
nor U704 (N_704,N_611,N_619);
or U705 (N_705,N_609,N_626);
and U706 (N_706,N_673,N_691);
nand U707 (N_707,N_654,N_605);
or U708 (N_708,N_641,N_632);
nor U709 (N_709,N_690,N_608);
and U710 (N_710,N_660,N_689);
nand U711 (N_711,N_645,N_694);
and U712 (N_712,N_618,N_613);
nor U713 (N_713,N_688,N_638);
and U714 (N_714,N_634,N_628);
or U715 (N_715,N_653,N_644);
nor U716 (N_716,N_674,N_677);
nand U717 (N_717,N_686,N_684);
and U718 (N_718,N_639,N_695);
or U719 (N_719,N_621,N_687);
and U720 (N_720,N_698,N_606);
nor U721 (N_721,N_651,N_612);
nand U722 (N_722,N_648,N_679);
or U723 (N_723,N_640,N_603);
nor U724 (N_724,N_655,N_617);
or U725 (N_725,N_623,N_699);
nand U726 (N_726,N_615,N_668);
and U727 (N_727,N_616,N_633);
nor U728 (N_728,N_678,N_607);
or U729 (N_729,N_646,N_625);
nand U730 (N_730,N_637,N_622);
nor U731 (N_731,N_680,N_627);
or U732 (N_732,N_631,N_604);
nor U733 (N_733,N_601,N_696);
and U734 (N_734,N_666,N_697);
nor U735 (N_735,N_656,N_620);
and U736 (N_736,N_649,N_647);
and U737 (N_737,N_685,N_659);
nand U738 (N_738,N_650,N_682);
nand U739 (N_739,N_672,N_663);
nor U740 (N_740,N_671,N_643);
nand U741 (N_741,N_635,N_658);
nand U742 (N_742,N_675,N_630);
nor U743 (N_743,N_667,N_610);
or U744 (N_744,N_652,N_624);
and U745 (N_745,N_642,N_693);
nor U746 (N_746,N_661,N_657);
nand U747 (N_747,N_602,N_664);
or U748 (N_748,N_669,N_636);
or U749 (N_749,N_662,N_681);
or U750 (N_750,N_619,N_625);
or U751 (N_751,N_642,N_694);
and U752 (N_752,N_696,N_645);
and U753 (N_753,N_600,N_678);
or U754 (N_754,N_619,N_665);
nor U755 (N_755,N_673,N_611);
or U756 (N_756,N_601,N_662);
nor U757 (N_757,N_680,N_696);
nand U758 (N_758,N_676,N_693);
nor U759 (N_759,N_637,N_682);
and U760 (N_760,N_678,N_681);
and U761 (N_761,N_643,N_699);
nand U762 (N_762,N_681,N_645);
and U763 (N_763,N_648,N_623);
or U764 (N_764,N_662,N_630);
nand U765 (N_765,N_632,N_611);
nor U766 (N_766,N_669,N_600);
and U767 (N_767,N_624,N_699);
nand U768 (N_768,N_608,N_698);
and U769 (N_769,N_626,N_673);
or U770 (N_770,N_691,N_699);
nand U771 (N_771,N_632,N_618);
nand U772 (N_772,N_662,N_628);
and U773 (N_773,N_674,N_631);
and U774 (N_774,N_618,N_652);
nand U775 (N_775,N_667,N_628);
or U776 (N_776,N_602,N_692);
nand U777 (N_777,N_672,N_661);
nand U778 (N_778,N_648,N_661);
or U779 (N_779,N_610,N_648);
nand U780 (N_780,N_686,N_672);
and U781 (N_781,N_648,N_665);
and U782 (N_782,N_696,N_623);
or U783 (N_783,N_695,N_613);
nand U784 (N_784,N_696,N_686);
nand U785 (N_785,N_693,N_666);
or U786 (N_786,N_631,N_679);
nand U787 (N_787,N_615,N_646);
or U788 (N_788,N_607,N_638);
and U789 (N_789,N_619,N_681);
and U790 (N_790,N_691,N_618);
and U791 (N_791,N_667,N_699);
or U792 (N_792,N_644,N_602);
nand U793 (N_793,N_660,N_648);
and U794 (N_794,N_612,N_648);
and U795 (N_795,N_660,N_655);
nor U796 (N_796,N_646,N_633);
nand U797 (N_797,N_651,N_676);
or U798 (N_798,N_612,N_665);
nor U799 (N_799,N_612,N_622);
or U800 (N_800,N_706,N_774);
nor U801 (N_801,N_799,N_790);
nand U802 (N_802,N_761,N_767);
nand U803 (N_803,N_762,N_729);
or U804 (N_804,N_741,N_777);
and U805 (N_805,N_758,N_719);
nor U806 (N_806,N_736,N_794);
nand U807 (N_807,N_735,N_721);
nor U808 (N_808,N_763,N_730);
nand U809 (N_809,N_705,N_704);
nand U810 (N_810,N_737,N_771);
or U811 (N_811,N_717,N_709);
and U812 (N_812,N_795,N_779);
nand U813 (N_813,N_703,N_742);
or U814 (N_814,N_712,N_796);
nand U815 (N_815,N_778,N_788);
nor U816 (N_816,N_747,N_759);
or U817 (N_817,N_789,N_720);
nand U818 (N_818,N_723,N_797);
or U819 (N_819,N_772,N_727);
and U820 (N_820,N_754,N_728);
nand U821 (N_821,N_773,N_775);
or U822 (N_822,N_748,N_766);
nor U823 (N_823,N_722,N_770);
and U824 (N_824,N_731,N_738);
nand U825 (N_825,N_750,N_769);
nand U826 (N_826,N_700,N_715);
and U827 (N_827,N_702,N_787);
or U828 (N_828,N_725,N_782);
or U829 (N_829,N_707,N_793);
nor U830 (N_830,N_739,N_708);
nand U831 (N_831,N_716,N_791);
and U832 (N_832,N_744,N_765);
nor U833 (N_833,N_781,N_751);
nand U834 (N_834,N_755,N_746);
and U835 (N_835,N_784,N_732);
nor U836 (N_836,N_733,N_710);
nand U837 (N_837,N_757,N_740);
or U838 (N_838,N_713,N_711);
nor U839 (N_839,N_798,N_714);
or U840 (N_840,N_783,N_776);
nor U841 (N_841,N_764,N_726);
and U842 (N_842,N_753,N_718);
nand U843 (N_843,N_743,N_701);
nand U844 (N_844,N_724,N_780);
nor U845 (N_845,N_792,N_734);
or U846 (N_846,N_768,N_760);
nor U847 (N_847,N_749,N_786);
or U848 (N_848,N_756,N_752);
and U849 (N_849,N_785,N_745);
and U850 (N_850,N_799,N_758);
and U851 (N_851,N_768,N_796);
nand U852 (N_852,N_748,N_705);
or U853 (N_853,N_783,N_720);
and U854 (N_854,N_789,N_744);
nand U855 (N_855,N_746,N_779);
or U856 (N_856,N_762,N_784);
or U857 (N_857,N_730,N_760);
nand U858 (N_858,N_703,N_711);
and U859 (N_859,N_777,N_732);
and U860 (N_860,N_731,N_709);
or U861 (N_861,N_701,N_726);
nor U862 (N_862,N_782,N_766);
nand U863 (N_863,N_747,N_776);
nor U864 (N_864,N_724,N_736);
nand U865 (N_865,N_755,N_730);
and U866 (N_866,N_790,N_776);
or U867 (N_867,N_734,N_773);
nor U868 (N_868,N_782,N_789);
or U869 (N_869,N_753,N_746);
and U870 (N_870,N_787,N_795);
nand U871 (N_871,N_768,N_700);
or U872 (N_872,N_798,N_742);
or U873 (N_873,N_705,N_749);
or U874 (N_874,N_730,N_707);
or U875 (N_875,N_738,N_777);
nand U876 (N_876,N_767,N_705);
or U877 (N_877,N_747,N_791);
or U878 (N_878,N_776,N_792);
and U879 (N_879,N_790,N_739);
and U880 (N_880,N_738,N_711);
xor U881 (N_881,N_711,N_794);
xnor U882 (N_882,N_739,N_706);
nor U883 (N_883,N_748,N_735);
nor U884 (N_884,N_794,N_726);
nand U885 (N_885,N_764,N_742);
or U886 (N_886,N_738,N_798);
and U887 (N_887,N_756,N_722);
nand U888 (N_888,N_799,N_723);
nand U889 (N_889,N_716,N_746);
nand U890 (N_890,N_788,N_702);
nor U891 (N_891,N_791,N_728);
xnor U892 (N_892,N_781,N_752);
nor U893 (N_893,N_708,N_793);
or U894 (N_894,N_742,N_792);
and U895 (N_895,N_788,N_720);
and U896 (N_896,N_715,N_730);
and U897 (N_897,N_716,N_710);
nor U898 (N_898,N_731,N_762);
or U899 (N_899,N_744,N_723);
nor U900 (N_900,N_828,N_826);
and U901 (N_901,N_807,N_849);
and U902 (N_902,N_824,N_883);
nand U903 (N_903,N_858,N_866);
and U904 (N_904,N_879,N_832);
nor U905 (N_905,N_861,N_888);
nand U906 (N_906,N_851,N_802);
and U907 (N_907,N_816,N_865);
and U908 (N_908,N_846,N_872);
nor U909 (N_909,N_889,N_871);
nor U910 (N_910,N_899,N_848);
or U911 (N_911,N_819,N_868);
nand U912 (N_912,N_880,N_839);
or U913 (N_913,N_894,N_829);
nand U914 (N_914,N_821,N_811);
and U915 (N_915,N_838,N_814);
nor U916 (N_916,N_809,N_867);
and U917 (N_917,N_827,N_820);
or U918 (N_918,N_898,N_804);
and U919 (N_919,N_891,N_840);
or U920 (N_920,N_853,N_886);
or U921 (N_921,N_857,N_887);
nand U922 (N_922,N_837,N_864);
nor U923 (N_923,N_801,N_847);
or U924 (N_924,N_815,N_800);
nor U925 (N_925,N_810,N_878);
nand U926 (N_926,N_859,N_825);
nor U927 (N_927,N_890,N_817);
or U928 (N_928,N_812,N_836);
and U929 (N_929,N_835,N_823);
nor U930 (N_930,N_841,N_895);
xor U931 (N_931,N_844,N_881);
nor U932 (N_932,N_822,N_854);
or U933 (N_933,N_805,N_875);
nor U934 (N_934,N_863,N_896);
or U935 (N_935,N_808,N_855);
nand U936 (N_936,N_856,N_842);
or U937 (N_937,N_818,N_870);
nand U938 (N_938,N_843,N_897);
or U939 (N_939,N_874,N_873);
nand U940 (N_940,N_877,N_852);
or U941 (N_941,N_834,N_813);
nand U942 (N_942,N_860,N_830);
nor U943 (N_943,N_831,N_893);
or U944 (N_944,N_884,N_806);
nand U945 (N_945,N_850,N_869);
nand U946 (N_946,N_876,N_803);
nor U947 (N_947,N_845,N_833);
and U948 (N_948,N_862,N_885);
or U949 (N_949,N_882,N_892);
nand U950 (N_950,N_895,N_856);
nand U951 (N_951,N_820,N_891);
xnor U952 (N_952,N_844,N_896);
and U953 (N_953,N_867,N_804);
and U954 (N_954,N_896,N_866);
and U955 (N_955,N_852,N_802);
nand U956 (N_956,N_878,N_893);
and U957 (N_957,N_896,N_867);
nand U958 (N_958,N_865,N_850);
and U959 (N_959,N_815,N_818);
and U960 (N_960,N_890,N_803);
nand U961 (N_961,N_868,N_855);
nor U962 (N_962,N_820,N_881);
or U963 (N_963,N_821,N_864);
nor U964 (N_964,N_876,N_877);
nor U965 (N_965,N_892,N_819);
nor U966 (N_966,N_829,N_800);
and U967 (N_967,N_873,N_802);
or U968 (N_968,N_882,N_873);
and U969 (N_969,N_844,N_880);
nor U970 (N_970,N_885,N_833);
nor U971 (N_971,N_863,N_885);
nand U972 (N_972,N_851,N_840);
or U973 (N_973,N_880,N_819);
or U974 (N_974,N_863,N_801);
nor U975 (N_975,N_844,N_897);
or U976 (N_976,N_890,N_826);
nor U977 (N_977,N_816,N_868);
or U978 (N_978,N_875,N_840);
and U979 (N_979,N_865,N_833);
and U980 (N_980,N_831,N_878);
or U981 (N_981,N_810,N_887);
or U982 (N_982,N_886,N_826);
and U983 (N_983,N_832,N_878);
or U984 (N_984,N_800,N_859);
and U985 (N_985,N_876,N_843);
or U986 (N_986,N_877,N_861);
nand U987 (N_987,N_813,N_888);
and U988 (N_988,N_869,N_866);
nand U989 (N_989,N_811,N_883);
or U990 (N_990,N_871,N_895);
and U991 (N_991,N_842,N_803);
nand U992 (N_992,N_873,N_885);
nor U993 (N_993,N_843,N_801);
or U994 (N_994,N_818,N_800);
or U995 (N_995,N_814,N_888);
and U996 (N_996,N_800,N_871);
and U997 (N_997,N_891,N_895);
nand U998 (N_998,N_875,N_855);
and U999 (N_999,N_813,N_876);
nand U1000 (N_1000,N_906,N_956);
nand U1001 (N_1001,N_943,N_974);
and U1002 (N_1002,N_977,N_948);
nor U1003 (N_1003,N_904,N_909);
or U1004 (N_1004,N_951,N_903);
and U1005 (N_1005,N_912,N_946);
and U1006 (N_1006,N_957,N_964);
nand U1007 (N_1007,N_966,N_952);
nor U1008 (N_1008,N_921,N_901);
and U1009 (N_1009,N_944,N_938);
nor U1010 (N_1010,N_962,N_985);
or U1011 (N_1011,N_900,N_907);
and U1012 (N_1012,N_945,N_959);
nor U1013 (N_1013,N_917,N_931);
nor U1014 (N_1014,N_984,N_999);
nor U1015 (N_1015,N_950,N_969);
or U1016 (N_1016,N_940,N_982);
nor U1017 (N_1017,N_942,N_914);
or U1018 (N_1018,N_955,N_923);
or U1019 (N_1019,N_934,N_973);
nand U1020 (N_1020,N_920,N_902);
nor U1021 (N_1021,N_961,N_989);
nand U1022 (N_1022,N_963,N_993);
xnor U1023 (N_1023,N_992,N_929);
or U1024 (N_1024,N_926,N_939);
nand U1025 (N_1025,N_972,N_918);
and U1026 (N_1026,N_910,N_997);
nand U1027 (N_1027,N_990,N_937);
nand U1028 (N_1028,N_970,N_935);
nor U1029 (N_1029,N_922,N_981);
nand U1030 (N_1030,N_928,N_932);
or U1031 (N_1031,N_915,N_953);
and U1032 (N_1032,N_933,N_908);
xor U1033 (N_1033,N_930,N_924);
or U1034 (N_1034,N_991,N_960);
xor U1035 (N_1035,N_996,N_987);
nand U1036 (N_1036,N_958,N_968);
nand U1037 (N_1037,N_954,N_998);
or U1038 (N_1038,N_905,N_986);
or U1039 (N_1039,N_965,N_983);
or U1040 (N_1040,N_927,N_913);
nand U1041 (N_1041,N_995,N_947);
nand U1042 (N_1042,N_925,N_949);
or U1043 (N_1043,N_971,N_988);
nand U1044 (N_1044,N_936,N_976);
nor U1045 (N_1045,N_941,N_911);
nand U1046 (N_1046,N_979,N_980);
and U1047 (N_1047,N_967,N_916);
nor U1048 (N_1048,N_978,N_994);
and U1049 (N_1049,N_975,N_919);
and U1050 (N_1050,N_921,N_939);
and U1051 (N_1051,N_934,N_965);
nand U1052 (N_1052,N_904,N_929);
nor U1053 (N_1053,N_945,N_919);
nand U1054 (N_1054,N_908,N_922);
and U1055 (N_1055,N_903,N_921);
nand U1056 (N_1056,N_998,N_905);
or U1057 (N_1057,N_958,N_992);
nand U1058 (N_1058,N_940,N_962);
and U1059 (N_1059,N_958,N_902);
and U1060 (N_1060,N_973,N_902);
nor U1061 (N_1061,N_947,N_991);
or U1062 (N_1062,N_910,N_955);
or U1063 (N_1063,N_961,N_972);
nor U1064 (N_1064,N_925,N_943);
and U1065 (N_1065,N_922,N_932);
or U1066 (N_1066,N_934,N_995);
nor U1067 (N_1067,N_900,N_983);
nor U1068 (N_1068,N_997,N_986);
nand U1069 (N_1069,N_937,N_945);
and U1070 (N_1070,N_914,N_948);
nor U1071 (N_1071,N_967,N_980);
nand U1072 (N_1072,N_924,N_957);
nor U1073 (N_1073,N_997,N_933);
nand U1074 (N_1074,N_993,N_962);
nor U1075 (N_1075,N_939,N_984);
nand U1076 (N_1076,N_974,N_996);
nand U1077 (N_1077,N_914,N_972);
and U1078 (N_1078,N_995,N_904);
or U1079 (N_1079,N_907,N_980);
and U1080 (N_1080,N_917,N_918);
nand U1081 (N_1081,N_991,N_953);
nand U1082 (N_1082,N_914,N_970);
and U1083 (N_1083,N_932,N_906);
nand U1084 (N_1084,N_939,N_950);
or U1085 (N_1085,N_946,N_969);
and U1086 (N_1086,N_964,N_924);
nand U1087 (N_1087,N_960,N_966);
nand U1088 (N_1088,N_983,N_960);
and U1089 (N_1089,N_952,N_987);
nand U1090 (N_1090,N_992,N_966);
or U1091 (N_1091,N_962,N_915);
and U1092 (N_1092,N_908,N_946);
or U1093 (N_1093,N_908,N_973);
nand U1094 (N_1094,N_962,N_957);
and U1095 (N_1095,N_911,N_985);
nor U1096 (N_1096,N_917,N_998);
or U1097 (N_1097,N_994,N_904);
nor U1098 (N_1098,N_981,N_900);
and U1099 (N_1099,N_917,N_905);
nor U1100 (N_1100,N_1043,N_1073);
and U1101 (N_1101,N_1093,N_1037);
or U1102 (N_1102,N_1034,N_1033);
nand U1103 (N_1103,N_1044,N_1057);
nand U1104 (N_1104,N_1065,N_1015);
nand U1105 (N_1105,N_1014,N_1042);
and U1106 (N_1106,N_1025,N_1078);
or U1107 (N_1107,N_1009,N_1017);
or U1108 (N_1108,N_1061,N_1022);
or U1109 (N_1109,N_1007,N_1028);
nor U1110 (N_1110,N_1000,N_1011);
and U1111 (N_1111,N_1077,N_1050);
nor U1112 (N_1112,N_1038,N_1096);
nand U1113 (N_1113,N_1045,N_1085);
and U1114 (N_1114,N_1010,N_1074);
nor U1115 (N_1115,N_1071,N_1002);
and U1116 (N_1116,N_1001,N_1026);
nor U1117 (N_1117,N_1004,N_1008);
nand U1118 (N_1118,N_1099,N_1082);
nor U1119 (N_1119,N_1092,N_1060);
nor U1120 (N_1120,N_1047,N_1070);
or U1121 (N_1121,N_1066,N_1097);
nor U1122 (N_1122,N_1013,N_1087);
nand U1123 (N_1123,N_1049,N_1086);
xor U1124 (N_1124,N_1051,N_1005);
and U1125 (N_1125,N_1076,N_1055);
or U1126 (N_1126,N_1053,N_1023);
nand U1127 (N_1127,N_1083,N_1068);
and U1128 (N_1128,N_1084,N_1021);
or U1129 (N_1129,N_1052,N_1035);
nor U1130 (N_1130,N_1046,N_1098);
and U1131 (N_1131,N_1088,N_1030);
and U1132 (N_1132,N_1036,N_1059);
or U1133 (N_1133,N_1029,N_1039);
nand U1134 (N_1134,N_1019,N_1024);
and U1135 (N_1135,N_1016,N_1056);
and U1136 (N_1136,N_1040,N_1072);
or U1137 (N_1137,N_1091,N_1075);
nand U1138 (N_1138,N_1054,N_1041);
or U1139 (N_1139,N_1006,N_1067);
or U1140 (N_1140,N_1032,N_1003);
and U1141 (N_1141,N_1048,N_1090);
and U1142 (N_1142,N_1058,N_1089);
or U1143 (N_1143,N_1069,N_1094);
and U1144 (N_1144,N_1080,N_1027);
nand U1145 (N_1145,N_1031,N_1081);
nand U1146 (N_1146,N_1018,N_1020);
nand U1147 (N_1147,N_1095,N_1062);
nand U1148 (N_1148,N_1079,N_1064);
nor U1149 (N_1149,N_1012,N_1063);
nor U1150 (N_1150,N_1007,N_1047);
nor U1151 (N_1151,N_1005,N_1024);
nand U1152 (N_1152,N_1053,N_1046);
nor U1153 (N_1153,N_1042,N_1090);
nor U1154 (N_1154,N_1091,N_1054);
or U1155 (N_1155,N_1041,N_1092);
or U1156 (N_1156,N_1047,N_1042);
nand U1157 (N_1157,N_1023,N_1011);
nor U1158 (N_1158,N_1091,N_1035);
and U1159 (N_1159,N_1016,N_1025);
nor U1160 (N_1160,N_1021,N_1027);
and U1161 (N_1161,N_1078,N_1006);
or U1162 (N_1162,N_1012,N_1067);
nand U1163 (N_1163,N_1062,N_1029);
nor U1164 (N_1164,N_1019,N_1086);
or U1165 (N_1165,N_1066,N_1061);
nor U1166 (N_1166,N_1020,N_1044);
nand U1167 (N_1167,N_1074,N_1018);
nand U1168 (N_1168,N_1017,N_1089);
or U1169 (N_1169,N_1049,N_1000);
and U1170 (N_1170,N_1094,N_1044);
nor U1171 (N_1171,N_1079,N_1035);
nand U1172 (N_1172,N_1066,N_1035);
nand U1173 (N_1173,N_1021,N_1034);
or U1174 (N_1174,N_1096,N_1006);
nand U1175 (N_1175,N_1081,N_1045);
nand U1176 (N_1176,N_1081,N_1033);
nor U1177 (N_1177,N_1079,N_1083);
and U1178 (N_1178,N_1037,N_1061);
nor U1179 (N_1179,N_1031,N_1086);
nor U1180 (N_1180,N_1094,N_1018);
or U1181 (N_1181,N_1024,N_1012);
nand U1182 (N_1182,N_1005,N_1071);
or U1183 (N_1183,N_1023,N_1061);
nor U1184 (N_1184,N_1026,N_1073);
nand U1185 (N_1185,N_1083,N_1060);
nor U1186 (N_1186,N_1082,N_1047);
or U1187 (N_1187,N_1050,N_1073);
nand U1188 (N_1188,N_1050,N_1005);
nand U1189 (N_1189,N_1056,N_1017);
and U1190 (N_1190,N_1063,N_1033);
or U1191 (N_1191,N_1077,N_1045);
and U1192 (N_1192,N_1066,N_1031);
or U1193 (N_1193,N_1030,N_1063);
and U1194 (N_1194,N_1078,N_1087);
and U1195 (N_1195,N_1041,N_1049);
nor U1196 (N_1196,N_1035,N_1009);
nor U1197 (N_1197,N_1051,N_1004);
and U1198 (N_1198,N_1009,N_1038);
nor U1199 (N_1199,N_1010,N_1036);
nand U1200 (N_1200,N_1190,N_1129);
nand U1201 (N_1201,N_1184,N_1171);
nor U1202 (N_1202,N_1166,N_1112);
nor U1203 (N_1203,N_1142,N_1198);
or U1204 (N_1204,N_1177,N_1138);
or U1205 (N_1205,N_1106,N_1187);
nor U1206 (N_1206,N_1183,N_1186);
or U1207 (N_1207,N_1102,N_1149);
and U1208 (N_1208,N_1117,N_1147);
and U1209 (N_1209,N_1157,N_1169);
or U1210 (N_1210,N_1113,N_1188);
and U1211 (N_1211,N_1123,N_1170);
or U1212 (N_1212,N_1132,N_1193);
or U1213 (N_1213,N_1192,N_1124);
nor U1214 (N_1214,N_1194,N_1182);
and U1215 (N_1215,N_1118,N_1144);
and U1216 (N_1216,N_1125,N_1191);
nor U1217 (N_1217,N_1148,N_1164);
or U1218 (N_1218,N_1101,N_1167);
nand U1219 (N_1219,N_1120,N_1126);
or U1220 (N_1220,N_1160,N_1179);
nor U1221 (N_1221,N_1131,N_1158);
and U1222 (N_1222,N_1181,N_1108);
nand U1223 (N_1223,N_1121,N_1172);
or U1224 (N_1224,N_1135,N_1146);
or U1225 (N_1225,N_1161,N_1134);
or U1226 (N_1226,N_1145,N_1168);
nand U1227 (N_1227,N_1154,N_1156);
and U1228 (N_1228,N_1185,N_1196);
nor U1229 (N_1229,N_1127,N_1128);
nand U1230 (N_1230,N_1155,N_1159);
nand U1231 (N_1231,N_1178,N_1133);
and U1232 (N_1232,N_1175,N_1165);
nor U1233 (N_1233,N_1119,N_1162);
nor U1234 (N_1234,N_1116,N_1153);
nor U1235 (N_1235,N_1173,N_1109);
nand U1236 (N_1236,N_1199,N_1104);
nand U1237 (N_1237,N_1180,N_1174);
and U1238 (N_1238,N_1107,N_1141);
nand U1239 (N_1239,N_1163,N_1110);
nor U1240 (N_1240,N_1105,N_1137);
nor U1241 (N_1241,N_1114,N_1103);
or U1242 (N_1242,N_1197,N_1189);
and U1243 (N_1243,N_1111,N_1122);
nand U1244 (N_1244,N_1139,N_1143);
nand U1245 (N_1245,N_1150,N_1176);
nand U1246 (N_1246,N_1130,N_1195);
nor U1247 (N_1247,N_1136,N_1115);
nand U1248 (N_1248,N_1152,N_1140);
nand U1249 (N_1249,N_1100,N_1151);
nor U1250 (N_1250,N_1156,N_1193);
and U1251 (N_1251,N_1151,N_1149);
or U1252 (N_1252,N_1136,N_1108);
or U1253 (N_1253,N_1181,N_1168);
or U1254 (N_1254,N_1194,N_1172);
nand U1255 (N_1255,N_1142,N_1129);
and U1256 (N_1256,N_1109,N_1152);
nand U1257 (N_1257,N_1169,N_1168);
nor U1258 (N_1258,N_1159,N_1194);
nor U1259 (N_1259,N_1183,N_1122);
nor U1260 (N_1260,N_1138,N_1148);
and U1261 (N_1261,N_1158,N_1171);
nand U1262 (N_1262,N_1181,N_1177);
or U1263 (N_1263,N_1123,N_1195);
or U1264 (N_1264,N_1142,N_1182);
nand U1265 (N_1265,N_1145,N_1178);
nand U1266 (N_1266,N_1156,N_1176);
and U1267 (N_1267,N_1177,N_1194);
nand U1268 (N_1268,N_1189,N_1147);
or U1269 (N_1269,N_1103,N_1109);
and U1270 (N_1270,N_1177,N_1161);
nor U1271 (N_1271,N_1177,N_1195);
and U1272 (N_1272,N_1108,N_1144);
or U1273 (N_1273,N_1129,N_1172);
and U1274 (N_1274,N_1146,N_1122);
or U1275 (N_1275,N_1194,N_1100);
and U1276 (N_1276,N_1134,N_1150);
or U1277 (N_1277,N_1170,N_1142);
or U1278 (N_1278,N_1181,N_1101);
and U1279 (N_1279,N_1111,N_1182);
nor U1280 (N_1280,N_1107,N_1108);
or U1281 (N_1281,N_1103,N_1189);
or U1282 (N_1282,N_1199,N_1128);
and U1283 (N_1283,N_1183,N_1125);
and U1284 (N_1284,N_1121,N_1111);
and U1285 (N_1285,N_1182,N_1121);
or U1286 (N_1286,N_1162,N_1122);
and U1287 (N_1287,N_1115,N_1149);
and U1288 (N_1288,N_1128,N_1124);
nor U1289 (N_1289,N_1178,N_1148);
or U1290 (N_1290,N_1167,N_1115);
or U1291 (N_1291,N_1111,N_1118);
nor U1292 (N_1292,N_1162,N_1156);
nand U1293 (N_1293,N_1136,N_1195);
nor U1294 (N_1294,N_1173,N_1199);
or U1295 (N_1295,N_1118,N_1180);
nor U1296 (N_1296,N_1150,N_1131);
nand U1297 (N_1297,N_1199,N_1108);
nor U1298 (N_1298,N_1176,N_1197);
and U1299 (N_1299,N_1145,N_1160);
or U1300 (N_1300,N_1253,N_1274);
and U1301 (N_1301,N_1297,N_1259);
nand U1302 (N_1302,N_1258,N_1265);
nor U1303 (N_1303,N_1213,N_1220);
and U1304 (N_1304,N_1207,N_1233);
and U1305 (N_1305,N_1249,N_1268);
nor U1306 (N_1306,N_1209,N_1251);
nor U1307 (N_1307,N_1202,N_1206);
nor U1308 (N_1308,N_1252,N_1267);
or U1309 (N_1309,N_1289,N_1266);
nor U1310 (N_1310,N_1255,N_1230);
nor U1311 (N_1311,N_1227,N_1235);
nand U1312 (N_1312,N_1234,N_1244);
and U1313 (N_1313,N_1270,N_1285);
nand U1314 (N_1314,N_1247,N_1257);
and U1315 (N_1315,N_1239,N_1210);
nor U1316 (N_1316,N_1275,N_1224);
or U1317 (N_1317,N_1283,N_1222);
nor U1318 (N_1318,N_1221,N_1250);
or U1319 (N_1319,N_1205,N_1236);
nor U1320 (N_1320,N_1272,N_1292);
nor U1321 (N_1321,N_1276,N_1240);
or U1322 (N_1322,N_1286,N_1228);
and U1323 (N_1323,N_1200,N_1204);
nand U1324 (N_1324,N_1260,N_1242);
nor U1325 (N_1325,N_1298,N_1291);
nand U1326 (N_1326,N_1225,N_1296);
and U1327 (N_1327,N_1269,N_1278);
and U1328 (N_1328,N_1263,N_1288);
nand U1329 (N_1329,N_1279,N_1254);
or U1330 (N_1330,N_1203,N_1246);
or U1331 (N_1331,N_1223,N_1261);
and U1332 (N_1332,N_1284,N_1219);
or U1333 (N_1333,N_1226,N_1243);
nor U1334 (N_1334,N_1280,N_1290);
nand U1335 (N_1335,N_1256,N_1248);
nand U1336 (N_1336,N_1216,N_1215);
nor U1337 (N_1337,N_1245,N_1277);
or U1338 (N_1338,N_1201,N_1264);
nor U1339 (N_1339,N_1229,N_1294);
nor U1340 (N_1340,N_1212,N_1217);
and U1341 (N_1341,N_1211,N_1262);
or U1342 (N_1342,N_1271,N_1282);
and U1343 (N_1343,N_1281,N_1218);
or U1344 (N_1344,N_1299,N_1231);
and U1345 (N_1345,N_1214,N_1295);
nand U1346 (N_1346,N_1237,N_1273);
nor U1347 (N_1347,N_1287,N_1238);
and U1348 (N_1348,N_1208,N_1293);
nor U1349 (N_1349,N_1241,N_1232);
nor U1350 (N_1350,N_1230,N_1241);
nand U1351 (N_1351,N_1293,N_1264);
nor U1352 (N_1352,N_1288,N_1285);
or U1353 (N_1353,N_1236,N_1253);
nor U1354 (N_1354,N_1256,N_1241);
nor U1355 (N_1355,N_1276,N_1225);
or U1356 (N_1356,N_1270,N_1206);
or U1357 (N_1357,N_1287,N_1286);
nor U1358 (N_1358,N_1217,N_1288);
nor U1359 (N_1359,N_1289,N_1246);
and U1360 (N_1360,N_1218,N_1262);
and U1361 (N_1361,N_1239,N_1245);
nor U1362 (N_1362,N_1295,N_1227);
or U1363 (N_1363,N_1220,N_1240);
and U1364 (N_1364,N_1267,N_1257);
nor U1365 (N_1365,N_1200,N_1234);
nor U1366 (N_1366,N_1244,N_1260);
or U1367 (N_1367,N_1213,N_1256);
nor U1368 (N_1368,N_1275,N_1289);
and U1369 (N_1369,N_1227,N_1276);
and U1370 (N_1370,N_1207,N_1229);
or U1371 (N_1371,N_1240,N_1264);
nand U1372 (N_1372,N_1291,N_1285);
and U1373 (N_1373,N_1226,N_1237);
and U1374 (N_1374,N_1229,N_1293);
nand U1375 (N_1375,N_1244,N_1241);
nor U1376 (N_1376,N_1226,N_1266);
nand U1377 (N_1377,N_1267,N_1223);
or U1378 (N_1378,N_1243,N_1256);
and U1379 (N_1379,N_1299,N_1285);
and U1380 (N_1380,N_1255,N_1251);
nand U1381 (N_1381,N_1246,N_1284);
nor U1382 (N_1382,N_1274,N_1279);
nor U1383 (N_1383,N_1215,N_1202);
and U1384 (N_1384,N_1251,N_1284);
nor U1385 (N_1385,N_1244,N_1223);
nand U1386 (N_1386,N_1237,N_1220);
nor U1387 (N_1387,N_1298,N_1239);
nor U1388 (N_1388,N_1265,N_1219);
or U1389 (N_1389,N_1285,N_1260);
nand U1390 (N_1390,N_1226,N_1227);
or U1391 (N_1391,N_1249,N_1260);
and U1392 (N_1392,N_1285,N_1258);
nand U1393 (N_1393,N_1279,N_1207);
nand U1394 (N_1394,N_1293,N_1223);
or U1395 (N_1395,N_1215,N_1297);
and U1396 (N_1396,N_1214,N_1230);
nand U1397 (N_1397,N_1212,N_1221);
and U1398 (N_1398,N_1205,N_1289);
nor U1399 (N_1399,N_1286,N_1275);
nor U1400 (N_1400,N_1385,N_1309);
nor U1401 (N_1401,N_1382,N_1306);
nand U1402 (N_1402,N_1376,N_1327);
and U1403 (N_1403,N_1392,N_1334);
nor U1404 (N_1404,N_1355,N_1318);
and U1405 (N_1405,N_1378,N_1329);
or U1406 (N_1406,N_1348,N_1386);
nor U1407 (N_1407,N_1379,N_1328);
nand U1408 (N_1408,N_1313,N_1350);
or U1409 (N_1409,N_1333,N_1361);
or U1410 (N_1410,N_1396,N_1398);
nand U1411 (N_1411,N_1391,N_1384);
and U1412 (N_1412,N_1305,N_1387);
and U1413 (N_1413,N_1357,N_1349);
nor U1414 (N_1414,N_1300,N_1336);
and U1415 (N_1415,N_1352,N_1359);
nor U1416 (N_1416,N_1372,N_1341);
nand U1417 (N_1417,N_1368,N_1314);
and U1418 (N_1418,N_1343,N_1363);
and U1419 (N_1419,N_1301,N_1337);
or U1420 (N_1420,N_1307,N_1340);
or U1421 (N_1421,N_1308,N_1390);
and U1422 (N_1422,N_1338,N_1393);
or U1423 (N_1423,N_1344,N_1389);
or U1424 (N_1424,N_1304,N_1369);
nor U1425 (N_1425,N_1325,N_1324);
nor U1426 (N_1426,N_1377,N_1310);
nand U1427 (N_1427,N_1321,N_1383);
nand U1428 (N_1428,N_1322,N_1358);
xor U1429 (N_1429,N_1375,N_1326);
and U1430 (N_1430,N_1356,N_1362);
nor U1431 (N_1431,N_1347,N_1335);
nand U1432 (N_1432,N_1332,N_1354);
and U1433 (N_1433,N_1345,N_1365);
nand U1434 (N_1434,N_1353,N_1388);
nand U1435 (N_1435,N_1302,N_1395);
and U1436 (N_1436,N_1371,N_1381);
nor U1437 (N_1437,N_1380,N_1346);
and U1438 (N_1438,N_1394,N_1316);
and U1439 (N_1439,N_1370,N_1360);
nor U1440 (N_1440,N_1303,N_1374);
nor U1441 (N_1441,N_1315,N_1339);
nand U1442 (N_1442,N_1366,N_1312);
nor U1443 (N_1443,N_1367,N_1399);
nand U1444 (N_1444,N_1397,N_1330);
nand U1445 (N_1445,N_1323,N_1342);
nand U1446 (N_1446,N_1373,N_1351);
nand U1447 (N_1447,N_1320,N_1311);
nor U1448 (N_1448,N_1364,N_1317);
or U1449 (N_1449,N_1319,N_1331);
or U1450 (N_1450,N_1303,N_1301);
or U1451 (N_1451,N_1330,N_1367);
or U1452 (N_1452,N_1346,N_1317);
nor U1453 (N_1453,N_1358,N_1382);
nor U1454 (N_1454,N_1336,N_1350);
and U1455 (N_1455,N_1308,N_1386);
nor U1456 (N_1456,N_1316,N_1324);
or U1457 (N_1457,N_1336,N_1313);
nor U1458 (N_1458,N_1302,N_1323);
nor U1459 (N_1459,N_1313,N_1311);
or U1460 (N_1460,N_1310,N_1399);
and U1461 (N_1461,N_1310,N_1387);
nand U1462 (N_1462,N_1326,N_1358);
nand U1463 (N_1463,N_1304,N_1368);
or U1464 (N_1464,N_1393,N_1333);
nor U1465 (N_1465,N_1348,N_1365);
or U1466 (N_1466,N_1300,N_1341);
or U1467 (N_1467,N_1359,N_1325);
and U1468 (N_1468,N_1357,N_1368);
nor U1469 (N_1469,N_1391,N_1334);
or U1470 (N_1470,N_1306,N_1367);
nand U1471 (N_1471,N_1302,N_1398);
or U1472 (N_1472,N_1399,N_1372);
or U1473 (N_1473,N_1335,N_1369);
or U1474 (N_1474,N_1350,N_1337);
nor U1475 (N_1475,N_1339,N_1389);
nor U1476 (N_1476,N_1360,N_1343);
and U1477 (N_1477,N_1376,N_1364);
nand U1478 (N_1478,N_1378,N_1343);
and U1479 (N_1479,N_1369,N_1365);
nor U1480 (N_1480,N_1339,N_1376);
or U1481 (N_1481,N_1328,N_1351);
nand U1482 (N_1482,N_1355,N_1352);
nor U1483 (N_1483,N_1382,N_1388);
and U1484 (N_1484,N_1339,N_1391);
nor U1485 (N_1485,N_1363,N_1383);
or U1486 (N_1486,N_1361,N_1334);
or U1487 (N_1487,N_1361,N_1353);
nor U1488 (N_1488,N_1388,N_1352);
and U1489 (N_1489,N_1310,N_1348);
and U1490 (N_1490,N_1398,N_1331);
and U1491 (N_1491,N_1319,N_1392);
nand U1492 (N_1492,N_1336,N_1332);
nor U1493 (N_1493,N_1324,N_1326);
nor U1494 (N_1494,N_1392,N_1397);
nand U1495 (N_1495,N_1318,N_1302);
nand U1496 (N_1496,N_1385,N_1306);
nor U1497 (N_1497,N_1320,N_1344);
nand U1498 (N_1498,N_1337,N_1335);
nor U1499 (N_1499,N_1350,N_1335);
or U1500 (N_1500,N_1459,N_1490);
or U1501 (N_1501,N_1415,N_1446);
or U1502 (N_1502,N_1435,N_1409);
nand U1503 (N_1503,N_1462,N_1466);
nand U1504 (N_1504,N_1456,N_1472);
and U1505 (N_1505,N_1455,N_1471);
and U1506 (N_1506,N_1478,N_1488);
nor U1507 (N_1507,N_1404,N_1485);
and U1508 (N_1508,N_1417,N_1448);
and U1509 (N_1509,N_1452,N_1438);
nand U1510 (N_1510,N_1439,N_1483);
or U1511 (N_1511,N_1467,N_1473);
xor U1512 (N_1512,N_1414,N_1422);
nand U1513 (N_1513,N_1420,N_1492);
or U1514 (N_1514,N_1425,N_1498);
and U1515 (N_1515,N_1461,N_1454);
and U1516 (N_1516,N_1480,N_1401);
nor U1517 (N_1517,N_1476,N_1423);
nor U1518 (N_1518,N_1445,N_1431);
and U1519 (N_1519,N_1405,N_1416);
xor U1520 (N_1520,N_1487,N_1436);
nor U1521 (N_1521,N_1486,N_1493);
nand U1522 (N_1522,N_1497,N_1407);
and U1523 (N_1523,N_1434,N_1491);
and U1524 (N_1524,N_1496,N_1457);
xnor U1525 (N_1525,N_1465,N_1463);
and U1526 (N_1526,N_1433,N_1470);
or U1527 (N_1527,N_1411,N_1477);
nand U1528 (N_1528,N_1447,N_1479);
nor U1529 (N_1529,N_1442,N_1408);
or U1530 (N_1530,N_1427,N_1410);
nor U1531 (N_1531,N_1421,N_1458);
nor U1532 (N_1532,N_1453,N_1451);
nand U1533 (N_1533,N_1494,N_1418);
and U1534 (N_1534,N_1428,N_1424);
and U1535 (N_1535,N_1402,N_1413);
nor U1536 (N_1536,N_1444,N_1460);
and U1537 (N_1537,N_1489,N_1495);
nor U1538 (N_1538,N_1400,N_1482);
or U1539 (N_1539,N_1403,N_1468);
nor U1540 (N_1540,N_1432,N_1481);
and U1541 (N_1541,N_1499,N_1475);
nand U1542 (N_1542,N_1440,N_1437);
nor U1543 (N_1543,N_1429,N_1412);
and U1544 (N_1544,N_1484,N_1419);
nor U1545 (N_1545,N_1430,N_1449);
or U1546 (N_1546,N_1469,N_1426);
nor U1547 (N_1547,N_1406,N_1474);
and U1548 (N_1548,N_1450,N_1443);
nor U1549 (N_1549,N_1464,N_1441);
or U1550 (N_1550,N_1491,N_1452);
and U1551 (N_1551,N_1457,N_1420);
and U1552 (N_1552,N_1432,N_1457);
nand U1553 (N_1553,N_1417,N_1434);
nand U1554 (N_1554,N_1416,N_1409);
nand U1555 (N_1555,N_1434,N_1418);
or U1556 (N_1556,N_1458,N_1454);
and U1557 (N_1557,N_1498,N_1424);
nand U1558 (N_1558,N_1492,N_1482);
nor U1559 (N_1559,N_1407,N_1485);
nor U1560 (N_1560,N_1465,N_1448);
or U1561 (N_1561,N_1422,N_1474);
or U1562 (N_1562,N_1478,N_1416);
and U1563 (N_1563,N_1447,N_1490);
nand U1564 (N_1564,N_1493,N_1435);
nor U1565 (N_1565,N_1430,N_1437);
nand U1566 (N_1566,N_1443,N_1435);
nand U1567 (N_1567,N_1405,N_1448);
nor U1568 (N_1568,N_1484,N_1486);
xnor U1569 (N_1569,N_1417,N_1487);
nand U1570 (N_1570,N_1434,N_1454);
nor U1571 (N_1571,N_1422,N_1436);
nand U1572 (N_1572,N_1486,N_1403);
nand U1573 (N_1573,N_1419,N_1470);
nor U1574 (N_1574,N_1413,N_1437);
nand U1575 (N_1575,N_1493,N_1465);
and U1576 (N_1576,N_1452,N_1401);
and U1577 (N_1577,N_1424,N_1429);
nor U1578 (N_1578,N_1451,N_1486);
and U1579 (N_1579,N_1444,N_1479);
or U1580 (N_1580,N_1490,N_1426);
and U1581 (N_1581,N_1466,N_1468);
or U1582 (N_1582,N_1462,N_1410);
nor U1583 (N_1583,N_1476,N_1449);
or U1584 (N_1584,N_1461,N_1426);
xnor U1585 (N_1585,N_1400,N_1479);
nor U1586 (N_1586,N_1439,N_1493);
nor U1587 (N_1587,N_1496,N_1486);
or U1588 (N_1588,N_1400,N_1406);
nand U1589 (N_1589,N_1488,N_1422);
nand U1590 (N_1590,N_1454,N_1448);
and U1591 (N_1591,N_1443,N_1409);
or U1592 (N_1592,N_1490,N_1446);
and U1593 (N_1593,N_1412,N_1489);
and U1594 (N_1594,N_1414,N_1433);
nand U1595 (N_1595,N_1496,N_1436);
and U1596 (N_1596,N_1422,N_1499);
nor U1597 (N_1597,N_1446,N_1421);
nor U1598 (N_1598,N_1414,N_1439);
nand U1599 (N_1599,N_1443,N_1411);
nand U1600 (N_1600,N_1562,N_1564);
or U1601 (N_1601,N_1516,N_1596);
nor U1602 (N_1602,N_1584,N_1583);
nor U1603 (N_1603,N_1511,N_1557);
or U1604 (N_1604,N_1598,N_1542);
and U1605 (N_1605,N_1568,N_1512);
nand U1606 (N_1606,N_1515,N_1591);
nor U1607 (N_1607,N_1588,N_1540);
or U1608 (N_1608,N_1525,N_1541);
nor U1609 (N_1609,N_1523,N_1529);
or U1610 (N_1610,N_1587,N_1551);
or U1611 (N_1611,N_1522,N_1517);
or U1612 (N_1612,N_1574,N_1509);
and U1613 (N_1613,N_1545,N_1592);
nor U1614 (N_1614,N_1501,N_1552);
nand U1615 (N_1615,N_1543,N_1559);
and U1616 (N_1616,N_1570,N_1510);
nor U1617 (N_1617,N_1544,N_1535);
or U1618 (N_1618,N_1573,N_1579);
xor U1619 (N_1619,N_1549,N_1558);
or U1620 (N_1620,N_1520,N_1585);
and U1621 (N_1621,N_1589,N_1528);
nor U1622 (N_1622,N_1597,N_1586);
or U1623 (N_1623,N_1537,N_1565);
and U1624 (N_1624,N_1554,N_1504);
and U1625 (N_1625,N_1563,N_1503);
and U1626 (N_1626,N_1576,N_1578);
nor U1627 (N_1627,N_1593,N_1531);
and U1628 (N_1628,N_1526,N_1536);
nor U1629 (N_1629,N_1566,N_1580);
and U1630 (N_1630,N_1594,N_1539);
nor U1631 (N_1631,N_1581,N_1507);
and U1632 (N_1632,N_1595,N_1508);
nand U1633 (N_1633,N_1590,N_1518);
nor U1634 (N_1634,N_1532,N_1505);
or U1635 (N_1635,N_1577,N_1547);
and U1636 (N_1636,N_1533,N_1514);
nor U1637 (N_1637,N_1569,N_1506);
and U1638 (N_1638,N_1502,N_1571);
nand U1639 (N_1639,N_1556,N_1524);
or U1640 (N_1640,N_1534,N_1575);
nor U1641 (N_1641,N_1530,N_1567);
nand U1642 (N_1642,N_1513,N_1500);
and U1643 (N_1643,N_1555,N_1553);
or U1644 (N_1644,N_1527,N_1519);
nand U1645 (N_1645,N_1548,N_1582);
nor U1646 (N_1646,N_1599,N_1572);
nand U1647 (N_1647,N_1561,N_1550);
nand U1648 (N_1648,N_1538,N_1521);
nor U1649 (N_1649,N_1560,N_1546);
and U1650 (N_1650,N_1563,N_1546);
or U1651 (N_1651,N_1559,N_1512);
nor U1652 (N_1652,N_1535,N_1571);
or U1653 (N_1653,N_1586,N_1595);
or U1654 (N_1654,N_1579,N_1552);
or U1655 (N_1655,N_1566,N_1534);
nor U1656 (N_1656,N_1534,N_1519);
nor U1657 (N_1657,N_1529,N_1595);
nand U1658 (N_1658,N_1557,N_1530);
xnor U1659 (N_1659,N_1590,N_1568);
nand U1660 (N_1660,N_1593,N_1595);
and U1661 (N_1661,N_1544,N_1550);
or U1662 (N_1662,N_1529,N_1519);
nand U1663 (N_1663,N_1562,N_1535);
nor U1664 (N_1664,N_1552,N_1591);
nor U1665 (N_1665,N_1542,N_1500);
nand U1666 (N_1666,N_1535,N_1507);
nand U1667 (N_1667,N_1564,N_1531);
or U1668 (N_1668,N_1539,N_1504);
and U1669 (N_1669,N_1506,N_1578);
or U1670 (N_1670,N_1584,N_1524);
nor U1671 (N_1671,N_1568,N_1587);
nand U1672 (N_1672,N_1589,N_1563);
nor U1673 (N_1673,N_1588,N_1551);
and U1674 (N_1674,N_1536,N_1568);
nand U1675 (N_1675,N_1516,N_1556);
or U1676 (N_1676,N_1578,N_1510);
nor U1677 (N_1677,N_1523,N_1540);
nand U1678 (N_1678,N_1518,N_1564);
or U1679 (N_1679,N_1527,N_1575);
and U1680 (N_1680,N_1598,N_1507);
nor U1681 (N_1681,N_1565,N_1589);
nor U1682 (N_1682,N_1568,N_1559);
and U1683 (N_1683,N_1541,N_1517);
nor U1684 (N_1684,N_1544,N_1537);
nand U1685 (N_1685,N_1594,N_1511);
nand U1686 (N_1686,N_1539,N_1560);
nand U1687 (N_1687,N_1505,N_1580);
and U1688 (N_1688,N_1510,N_1528);
nor U1689 (N_1689,N_1589,N_1574);
nand U1690 (N_1690,N_1540,N_1504);
nor U1691 (N_1691,N_1582,N_1506);
or U1692 (N_1692,N_1563,N_1534);
nor U1693 (N_1693,N_1500,N_1597);
nor U1694 (N_1694,N_1583,N_1533);
and U1695 (N_1695,N_1579,N_1578);
and U1696 (N_1696,N_1560,N_1503);
or U1697 (N_1697,N_1573,N_1532);
nor U1698 (N_1698,N_1506,N_1554);
nor U1699 (N_1699,N_1500,N_1564);
or U1700 (N_1700,N_1629,N_1651);
or U1701 (N_1701,N_1654,N_1670);
nand U1702 (N_1702,N_1611,N_1622);
or U1703 (N_1703,N_1658,N_1603);
nor U1704 (N_1704,N_1668,N_1614);
and U1705 (N_1705,N_1641,N_1683);
and U1706 (N_1706,N_1632,N_1619);
nand U1707 (N_1707,N_1694,N_1672);
nor U1708 (N_1708,N_1636,N_1631);
nor U1709 (N_1709,N_1613,N_1689);
or U1710 (N_1710,N_1627,N_1690);
nand U1711 (N_1711,N_1692,N_1676);
nor U1712 (N_1712,N_1663,N_1648);
nand U1713 (N_1713,N_1698,N_1643);
and U1714 (N_1714,N_1644,N_1695);
or U1715 (N_1715,N_1645,N_1688);
nor U1716 (N_1716,N_1665,N_1621);
or U1717 (N_1717,N_1691,N_1617);
nor U1718 (N_1718,N_1693,N_1661);
or U1719 (N_1719,N_1681,N_1673);
nand U1720 (N_1720,N_1615,N_1649);
and U1721 (N_1721,N_1675,N_1669);
and U1722 (N_1722,N_1600,N_1640);
nand U1723 (N_1723,N_1653,N_1623);
or U1724 (N_1724,N_1697,N_1642);
nor U1725 (N_1725,N_1671,N_1606);
or U1726 (N_1726,N_1626,N_1667);
and U1727 (N_1727,N_1680,N_1609);
nand U1728 (N_1728,N_1635,N_1628);
nand U1729 (N_1729,N_1679,N_1655);
or U1730 (N_1730,N_1678,N_1620);
and U1731 (N_1731,N_1659,N_1616);
nand U1732 (N_1732,N_1624,N_1684);
and U1733 (N_1733,N_1607,N_1638);
nor U1734 (N_1734,N_1656,N_1639);
and U1735 (N_1735,N_1662,N_1686);
or U1736 (N_1736,N_1610,N_1682);
nor U1737 (N_1737,N_1652,N_1647);
and U1738 (N_1738,N_1602,N_1612);
nor U1739 (N_1739,N_1608,N_1604);
and U1740 (N_1740,N_1699,N_1601);
nor U1741 (N_1741,N_1685,N_1618);
nand U1742 (N_1742,N_1650,N_1696);
or U1743 (N_1743,N_1657,N_1605);
nor U1744 (N_1744,N_1687,N_1664);
and U1745 (N_1745,N_1674,N_1634);
or U1746 (N_1746,N_1677,N_1646);
or U1747 (N_1747,N_1630,N_1637);
nor U1748 (N_1748,N_1666,N_1633);
nor U1749 (N_1749,N_1625,N_1660);
and U1750 (N_1750,N_1632,N_1604);
or U1751 (N_1751,N_1654,N_1601);
nor U1752 (N_1752,N_1686,N_1650);
nand U1753 (N_1753,N_1652,N_1606);
nand U1754 (N_1754,N_1686,N_1645);
and U1755 (N_1755,N_1691,N_1620);
nand U1756 (N_1756,N_1680,N_1626);
nor U1757 (N_1757,N_1687,N_1674);
or U1758 (N_1758,N_1643,N_1617);
or U1759 (N_1759,N_1605,N_1625);
nor U1760 (N_1760,N_1618,N_1698);
and U1761 (N_1761,N_1644,N_1632);
and U1762 (N_1762,N_1691,N_1631);
nor U1763 (N_1763,N_1613,N_1621);
nor U1764 (N_1764,N_1659,N_1674);
nor U1765 (N_1765,N_1641,N_1661);
nand U1766 (N_1766,N_1658,N_1686);
and U1767 (N_1767,N_1686,N_1633);
xnor U1768 (N_1768,N_1656,N_1635);
nor U1769 (N_1769,N_1628,N_1632);
nand U1770 (N_1770,N_1678,N_1627);
or U1771 (N_1771,N_1688,N_1670);
nor U1772 (N_1772,N_1672,N_1654);
nand U1773 (N_1773,N_1695,N_1679);
nor U1774 (N_1774,N_1688,N_1660);
or U1775 (N_1775,N_1649,N_1646);
nor U1776 (N_1776,N_1646,N_1666);
nor U1777 (N_1777,N_1678,N_1653);
nor U1778 (N_1778,N_1623,N_1618);
and U1779 (N_1779,N_1609,N_1608);
or U1780 (N_1780,N_1699,N_1604);
or U1781 (N_1781,N_1622,N_1669);
nand U1782 (N_1782,N_1628,N_1681);
or U1783 (N_1783,N_1651,N_1642);
nand U1784 (N_1784,N_1614,N_1674);
nor U1785 (N_1785,N_1654,N_1614);
or U1786 (N_1786,N_1681,N_1621);
nor U1787 (N_1787,N_1651,N_1694);
nand U1788 (N_1788,N_1666,N_1655);
and U1789 (N_1789,N_1678,N_1641);
nand U1790 (N_1790,N_1621,N_1626);
and U1791 (N_1791,N_1677,N_1691);
nand U1792 (N_1792,N_1684,N_1667);
and U1793 (N_1793,N_1663,N_1686);
nor U1794 (N_1794,N_1651,N_1679);
and U1795 (N_1795,N_1606,N_1620);
or U1796 (N_1796,N_1695,N_1655);
nand U1797 (N_1797,N_1689,N_1675);
and U1798 (N_1798,N_1664,N_1686);
or U1799 (N_1799,N_1626,N_1652);
and U1800 (N_1800,N_1785,N_1743);
nor U1801 (N_1801,N_1786,N_1729);
and U1802 (N_1802,N_1755,N_1713);
or U1803 (N_1803,N_1773,N_1775);
nor U1804 (N_1804,N_1744,N_1715);
nand U1805 (N_1805,N_1769,N_1737);
and U1806 (N_1806,N_1712,N_1719);
and U1807 (N_1807,N_1752,N_1738);
or U1808 (N_1808,N_1794,N_1795);
nand U1809 (N_1809,N_1761,N_1706);
nor U1810 (N_1810,N_1768,N_1747);
xor U1811 (N_1811,N_1776,N_1745);
and U1812 (N_1812,N_1700,N_1753);
and U1813 (N_1813,N_1790,N_1726);
and U1814 (N_1814,N_1704,N_1718);
or U1815 (N_1815,N_1716,N_1748);
nor U1816 (N_1816,N_1791,N_1739);
and U1817 (N_1817,N_1778,N_1732);
nand U1818 (N_1818,N_1721,N_1707);
nand U1819 (N_1819,N_1777,N_1764);
nand U1820 (N_1820,N_1735,N_1724);
or U1821 (N_1821,N_1772,N_1740);
and U1822 (N_1822,N_1703,N_1770);
nor U1823 (N_1823,N_1774,N_1731);
nand U1824 (N_1824,N_1758,N_1787);
nor U1825 (N_1825,N_1711,N_1798);
nand U1826 (N_1826,N_1710,N_1754);
nand U1827 (N_1827,N_1742,N_1727);
nor U1828 (N_1828,N_1750,N_1788);
nor U1829 (N_1829,N_1779,N_1723);
or U1830 (N_1830,N_1781,N_1783);
and U1831 (N_1831,N_1771,N_1725);
or U1832 (N_1832,N_1762,N_1701);
nand U1833 (N_1833,N_1717,N_1741);
and U1834 (N_1834,N_1765,N_1766);
and U1835 (N_1835,N_1789,N_1782);
and U1836 (N_1836,N_1702,N_1714);
or U1837 (N_1837,N_1708,N_1746);
and U1838 (N_1838,N_1733,N_1767);
and U1839 (N_1839,N_1736,N_1705);
and U1840 (N_1840,N_1756,N_1760);
nor U1841 (N_1841,N_1734,N_1763);
or U1842 (N_1842,N_1792,N_1749);
or U1843 (N_1843,N_1780,N_1730);
nand U1844 (N_1844,N_1793,N_1722);
nor U1845 (N_1845,N_1759,N_1751);
and U1846 (N_1846,N_1799,N_1796);
or U1847 (N_1847,N_1728,N_1757);
or U1848 (N_1848,N_1720,N_1784);
or U1849 (N_1849,N_1709,N_1797);
or U1850 (N_1850,N_1707,N_1771);
nor U1851 (N_1851,N_1746,N_1705);
nand U1852 (N_1852,N_1741,N_1783);
nor U1853 (N_1853,N_1745,N_1704);
or U1854 (N_1854,N_1787,N_1795);
or U1855 (N_1855,N_1770,N_1794);
nor U1856 (N_1856,N_1729,N_1753);
or U1857 (N_1857,N_1703,N_1793);
nand U1858 (N_1858,N_1788,N_1789);
or U1859 (N_1859,N_1711,N_1756);
and U1860 (N_1860,N_1793,N_1782);
or U1861 (N_1861,N_1748,N_1738);
nand U1862 (N_1862,N_1723,N_1769);
or U1863 (N_1863,N_1776,N_1725);
nor U1864 (N_1864,N_1752,N_1737);
or U1865 (N_1865,N_1759,N_1712);
or U1866 (N_1866,N_1754,N_1748);
nor U1867 (N_1867,N_1768,N_1758);
nor U1868 (N_1868,N_1792,N_1739);
nand U1869 (N_1869,N_1797,N_1756);
nor U1870 (N_1870,N_1707,N_1755);
nand U1871 (N_1871,N_1792,N_1736);
nor U1872 (N_1872,N_1764,N_1751);
or U1873 (N_1873,N_1793,N_1715);
or U1874 (N_1874,N_1745,N_1790);
nand U1875 (N_1875,N_1779,N_1706);
and U1876 (N_1876,N_1738,N_1792);
nor U1877 (N_1877,N_1772,N_1753);
nand U1878 (N_1878,N_1705,N_1795);
nor U1879 (N_1879,N_1793,N_1754);
and U1880 (N_1880,N_1757,N_1706);
or U1881 (N_1881,N_1773,N_1799);
or U1882 (N_1882,N_1700,N_1738);
or U1883 (N_1883,N_1783,N_1798);
or U1884 (N_1884,N_1760,N_1795);
and U1885 (N_1885,N_1734,N_1705);
nand U1886 (N_1886,N_1710,N_1782);
nor U1887 (N_1887,N_1704,N_1741);
and U1888 (N_1888,N_1789,N_1768);
and U1889 (N_1889,N_1721,N_1731);
or U1890 (N_1890,N_1773,N_1748);
nor U1891 (N_1891,N_1798,N_1733);
and U1892 (N_1892,N_1783,N_1787);
nand U1893 (N_1893,N_1741,N_1773);
nand U1894 (N_1894,N_1779,N_1784);
nor U1895 (N_1895,N_1791,N_1730);
nand U1896 (N_1896,N_1745,N_1713);
nor U1897 (N_1897,N_1733,N_1740);
and U1898 (N_1898,N_1799,N_1757);
and U1899 (N_1899,N_1785,N_1742);
or U1900 (N_1900,N_1878,N_1807);
and U1901 (N_1901,N_1830,N_1825);
and U1902 (N_1902,N_1895,N_1885);
and U1903 (N_1903,N_1868,N_1853);
or U1904 (N_1904,N_1823,N_1871);
and U1905 (N_1905,N_1877,N_1816);
or U1906 (N_1906,N_1874,N_1862);
xnor U1907 (N_1907,N_1858,N_1847);
or U1908 (N_1908,N_1812,N_1886);
or U1909 (N_1909,N_1839,N_1811);
nor U1910 (N_1910,N_1815,N_1840);
nor U1911 (N_1911,N_1863,N_1873);
or U1912 (N_1912,N_1827,N_1883);
nor U1913 (N_1913,N_1801,N_1891);
nand U1914 (N_1914,N_1829,N_1844);
nand U1915 (N_1915,N_1896,N_1899);
or U1916 (N_1916,N_1897,N_1884);
nand U1917 (N_1917,N_1864,N_1842);
nand U1918 (N_1918,N_1861,N_1805);
and U1919 (N_1919,N_1870,N_1892);
and U1920 (N_1920,N_1894,N_1845);
or U1921 (N_1921,N_1820,N_1869);
nand U1922 (N_1922,N_1887,N_1826);
or U1923 (N_1923,N_1851,N_1879);
and U1924 (N_1924,N_1833,N_1843);
nor U1925 (N_1925,N_1867,N_1808);
nor U1926 (N_1926,N_1837,N_1865);
nor U1927 (N_1927,N_1836,N_1814);
and U1928 (N_1928,N_1809,N_1898);
and U1929 (N_1929,N_1866,N_1880);
nand U1930 (N_1930,N_1838,N_1893);
and U1931 (N_1931,N_1806,N_1855);
or U1932 (N_1932,N_1859,N_1835);
and U1933 (N_1933,N_1856,N_1803);
and U1934 (N_1934,N_1860,N_1817);
nand U1935 (N_1935,N_1875,N_1821);
and U1936 (N_1936,N_1881,N_1890);
nor U1937 (N_1937,N_1876,N_1841);
nor U1938 (N_1938,N_1834,N_1819);
and U1939 (N_1939,N_1848,N_1822);
nor U1940 (N_1940,N_1810,N_1888);
nor U1941 (N_1941,N_1804,N_1813);
and U1942 (N_1942,N_1828,N_1831);
nor U1943 (N_1943,N_1854,N_1882);
and U1944 (N_1944,N_1889,N_1802);
nor U1945 (N_1945,N_1832,N_1852);
xor U1946 (N_1946,N_1872,N_1857);
nor U1947 (N_1947,N_1850,N_1800);
nand U1948 (N_1948,N_1824,N_1846);
or U1949 (N_1949,N_1818,N_1849);
and U1950 (N_1950,N_1889,N_1873);
nor U1951 (N_1951,N_1869,N_1891);
or U1952 (N_1952,N_1858,N_1835);
nand U1953 (N_1953,N_1865,N_1879);
and U1954 (N_1954,N_1852,N_1859);
nand U1955 (N_1955,N_1887,N_1812);
or U1956 (N_1956,N_1816,N_1817);
or U1957 (N_1957,N_1829,N_1823);
or U1958 (N_1958,N_1889,N_1844);
and U1959 (N_1959,N_1898,N_1887);
and U1960 (N_1960,N_1897,N_1853);
and U1961 (N_1961,N_1836,N_1878);
or U1962 (N_1962,N_1862,N_1851);
nand U1963 (N_1963,N_1828,N_1846);
nor U1964 (N_1964,N_1818,N_1897);
or U1965 (N_1965,N_1800,N_1844);
nor U1966 (N_1966,N_1895,N_1833);
nor U1967 (N_1967,N_1817,N_1849);
nor U1968 (N_1968,N_1873,N_1856);
nand U1969 (N_1969,N_1810,N_1801);
nand U1970 (N_1970,N_1884,N_1837);
nand U1971 (N_1971,N_1813,N_1866);
and U1972 (N_1972,N_1827,N_1843);
or U1973 (N_1973,N_1886,N_1882);
or U1974 (N_1974,N_1865,N_1871);
nand U1975 (N_1975,N_1879,N_1874);
nor U1976 (N_1976,N_1869,N_1859);
or U1977 (N_1977,N_1890,N_1815);
or U1978 (N_1978,N_1886,N_1888);
nand U1979 (N_1979,N_1871,N_1864);
and U1980 (N_1980,N_1850,N_1806);
and U1981 (N_1981,N_1898,N_1866);
and U1982 (N_1982,N_1828,N_1812);
nand U1983 (N_1983,N_1868,N_1875);
and U1984 (N_1984,N_1804,N_1850);
and U1985 (N_1985,N_1835,N_1846);
and U1986 (N_1986,N_1825,N_1851);
nand U1987 (N_1987,N_1827,N_1835);
nand U1988 (N_1988,N_1863,N_1802);
or U1989 (N_1989,N_1828,N_1837);
nand U1990 (N_1990,N_1864,N_1868);
nor U1991 (N_1991,N_1867,N_1829);
nand U1992 (N_1992,N_1884,N_1829);
nand U1993 (N_1993,N_1868,N_1897);
and U1994 (N_1994,N_1838,N_1858);
or U1995 (N_1995,N_1849,N_1847);
nand U1996 (N_1996,N_1881,N_1869);
nor U1997 (N_1997,N_1831,N_1817);
nand U1998 (N_1998,N_1823,N_1821);
nor U1999 (N_1999,N_1896,N_1830);
nor U2000 (N_2000,N_1947,N_1967);
nor U2001 (N_2001,N_1981,N_1954);
or U2002 (N_2002,N_1908,N_1999);
nand U2003 (N_2003,N_1905,N_1909);
nor U2004 (N_2004,N_1902,N_1972);
nand U2005 (N_2005,N_1918,N_1946);
nand U2006 (N_2006,N_1955,N_1929);
and U2007 (N_2007,N_1921,N_1997);
and U2008 (N_2008,N_1951,N_1978);
nor U2009 (N_2009,N_1957,N_1958);
nand U2010 (N_2010,N_1991,N_1937);
nor U2011 (N_2011,N_1989,N_1906);
or U2012 (N_2012,N_1984,N_1959);
nor U2013 (N_2013,N_1971,N_1940);
nor U2014 (N_2014,N_1930,N_1965);
and U2015 (N_2015,N_1962,N_1924);
nor U2016 (N_2016,N_1996,N_1952);
or U2017 (N_2017,N_1915,N_1956);
nor U2018 (N_2018,N_1976,N_1975);
nor U2019 (N_2019,N_1919,N_1966);
and U2020 (N_2020,N_1953,N_1987);
xnor U2021 (N_2021,N_1903,N_1993);
nor U2022 (N_2022,N_1963,N_1970);
and U2023 (N_2023,N_1934,N_1920);
nor U2024 (N_2024,N_1995,N_1904);
nand U2025 (N_2025,N_1948,N_1925);
nand U2026 (N_2026,N_1922,N_1979);
nand U2027 (N_2027,N_1938,N_1933);
nand U2028 (N_2028,N_1973,N_1914);
nor U2029 (N_2029,N_1986,N_1910);
nand U2030 (N_2030,N_1950,N_1968);
or U2031 (N_2031,N_1943,N_1932);
and U2032 (N_2032,N_1911,N_1985);
or U2033 (N_2033,N_1969,N_1917);
and U2034 (N_2034,N_1942,N_1982);
and U2035 (N_2035,N_1927,N_1974);
nand U2036 (N_2036,N_1907,N_1912);
and U2037 (N_2037,N_1900,N_1928);
and U2038 (N_2038,N_1961,N_1988);
and U2039 (N_2039,N_1926,N_1994);
and U2040 (N_2040,N_1944,N_1941);
nand U2041 (N_2041,N_1936,N_1945);
nor U2042 (N_2042,N_1949,N_1913);
or U2043 (N_2043,N_1977,N_1916);
or U2044 (N_2044,N_1983,N_1990);
and U2045 (N_2045,N_1931,N_1992);
nand U2046 (N_2046,N_1923,N_1964);
and U2047 (N_2047,N_1960,N_1998);
and U2048 (N_2048,N_1901,N_1939);
or U2049 (N_2049,N_1980,N_1935);
or U2050 (N_2050,N_1944,N_1909);
nand U2051 (N_2051,N_1987,N_1997);
and U2052 (N_2052,N_1936,N_1923);
nor U2053 (N_2053,N_1951,N_1907);
nand U2054 (N_2054,N_1966,N_1999);
and U2055 (N_2055,N_1911,N_1980);
nand U2056 (N_2056,N_1970,N_1964);
and U2057 (N_2057,N_1981,N_1955);
and U2058 (N_2058,N_1928,N_1927);
and U2059 (N_2059,N_1987,N_1940);
or U2060 (N_2060,N_1945,N_1913);
and U2061 (N_2061,N_1933,N_1960);
nor U2062 (N_2062,N_1923,N_1949);
nand U2063 (N_2063,N_1936,N_1908);
nor U2064 (N_2064,N_1904,N_1974);
nor U2065 (N_2065,N_1963,N_1926);
nor U2066 (N_2066,N_1910,N_1987);
nor U2067 (N_2067,N_1914,N_1951);
or U2068 (N_2068,N_1951,N_1995);
nor U2069 (N_2069,N_1962,N_1974);
or U2070 (N_2070,N_1938,N_1993);
nand U2071 (N_2071,N_1958,N_1929);
nor U2072 (N_2072,N_1914,N_1964);
nand U2073 (N_2073,N_1984,N_1945);
and U2074 (N_2074,N_1924,N_1947);
nor U2075 (N_2075,N_1999,N_1949);
nand U2076 (N_2076,N_1913,N_1936);
nor U2077 (N_2077,N_1979,N_1942);
nand U2078 (N_2078,N_1981,N_1984);
nor U2079 (N_2079,N_1954,N_1935);
nand U2080 (N_2080,N_1954,N_1996);
and U2081 (N_2081,N_1927,N_1945);
nand U2082 (N_2082,N_1974,N_1938);
nor U2083 (N_2083,N_1980,N_1992);
nand U2084 (N_2084,N_1936,N_1939);
nand U2085 (N_2085,N_1961,N_1939);
and U2086 (N_2086,N_1911,N_1981);
nand U2087 (N_2087,N_1959,N_1972);
nor U2088 (N_2088,N_1981,N_1992);
nand U2089 (N_2089,N_1932,N_1916);
nor U2090 (N_2090,N_1930,N_1931);
nor U2091 (N_2091,N_1918,N_1965);
or U2092 (N_2092,N_1900,N_1985);
nor U2093 (N_2093,N_1965,N_1962);
xor U2094 (N_2094,N_1974,N_1963);
or U2095 (N_2095,N_1903,N_1913);
nor U2096 (N_2096,N_1904,N_1989);
and U2097 (N_2097,N_1948,N_1967);
nor U2098 (N_2098,N_1969,N_1912);
nor U2099 (N_2099,N_1983,N_1948);
nor U2100 (N_2100,N_2077,N_2063);
and U2101 (N_2101,N_2031,N_2083);
and U2102 (N_2102,N_2015,N_2017);
nand U2103 (N_2103,N_2042,N_2024);
nand U2104 (N_2104,N_2068,N_2036);
nand U2105 (N_2105,N_2090,N_2050);
nand U2106 (N_2106,N_2074,N_2045);
nand U2107 (N_2107,N_2080,N_2094);
nand U2108 (N_2108,N_2071,N_2041);
or U2109 (N_2109,N_2034,N_2095);
nand U2110 (N_2110,N_2049,N_2084);
nor U2111 (N_2111,N_2005,N_2073);
nand U2112 (N_2112,N_2099,N_2023);
nor U2113 (N_2113,N_2048,N_2053);
nand U2114 (N_2114,N_2059,N_2032);
nand U2115 (N_2115,N_2087,N_2093);
or U2116 (N_2116,N_2027,N_2029);
and U2117 (N_2117,N_2019,N_2052);
nand U2118 (N_2118,N_2044,N_2020);
or U2119 (N_2119,N_2009,N_2057);
nor U2120 (N_2120,N_2067,N_2086);
and U2121 (N_2121,N_2060,N_2081);
nor U2122 (N_2122,N_2003,N_2066);
and U2123 (N_2123,N_2091,N_2070);
nor U2124 (N_2124,N_2078,N_2000);
nor U2125 (N_2125,N_2006,N_2039);
xor U2126 (N_2126,N_2011,N_2037);
nor U2127 (N_2127,N_2061,N_2016);
and U2128 (N_2128,N_2012,N_2054);
nor U2129 (N_2129,N_2075,N_2013);
nand U2130 (N_2130,N_2001,N_2082);
nor U2131 (N_2131,N_2025,N_2043);
xnor U2132 (N_2132,N_2018,N_2097);
nand U2133 (N_2133,N_2007,N_2069);
or U2134 (N_2134,N_2072,N_2079);
and U2135 (N_2135,N_2056,N_2008);
nand U2136 (N_2136,N_2096,N_2092);
nor U2137 (N_2137,N_2028,N_2047);
nor U2138 (N_2138,N_2051,N_2010);
or U2139 (N_2139,N_2062,N_2022);
nor U2140 (N_2140,N_2002,N_2046);
nand U2141 (N_2141,N_2064,N_2065);
xor U2142 (N_2142,N_2040,N_2085);
nor U2143 (N_2143,N_2088,N_2076);
nand U2144 (N_2144,N_2055,N_2030);
nand U2145 (N_2145,N_2058,N_2026);
nand U2146 (N_2146,N_2038,N_2098);
and U2147 (N_2147,N_2004,N_2035);
or U2148 (N_2148,N_2033,N_2089);
or U2149 (N_2149,N_2021,N_2014);
xnor U2150 (N_2150,N_2062,N_2080);
nor U2151 (N_2151,N_2034,N_2038);
nand U2152 (N_2152,N_2062,N_2026);
nand U2153 (N_2153,N_2063,N_2051);
nand U2154 (N_2154,N_2004,N_2006);
nor U2155 (N_2155,N_2066,N_2056);
and U2156 (N_2156,N_2010,N_2092);
nor U2157 (N_2157,N_2004,N_2058);
nor U2158 (N_2158,N_2030,N_2088);
nand U2159 (N_2159,N_2073,N_2030);
nor U2160 (N_2160,N_2035,N_2076);
and U2161 (N_2161,N_2099,N_2071);
nand U2162 (N_2162,N_2042,N_2056);
and U2163 (N_2163,N_2034,N_2093);
nor U2164 (N_2164,N_2095,N_2067);
nand U2165 (N_2165,N_2030,N_2038);
nand U2166 (N_2166,N_2040,N_2051);
nor U2167 (N_2167,N_2047,N_2016);
nor U2168 (N_2168,N_2038,N_2025);
and U2169 (N_2169,N_2030,N_2074);
and U2170 (N_2170,N_2061,N_2098);
nand U2171 (N_2171,N_2073,N_2070);
nor U2172 (N_2172,N_2011,N_2067);
or U2173 (N_2173,N_2002,N_2061);
nand U2174 (N_2174,N_2066,N_2015);
and U2175 (N_2175,N_2091,N_2046);
nand U2176 (N_2176,N_2000,N_2007);
nand U2177 (N_2177,N_2008,N_2088);
or U2178 (N_2178,N_2026,N_2081);
and U2179 (N_2179,N_2028,N_2048);
nor U2180 (N_2180,N_2006,N_2028);
nand U2181 (N_2181,N_2056,N_2061);
or U2182 (N_2182,N_2098,N_2064);
nor U2183 (N_2183,N_2061,N_2029);
nand U2184 (N_2184,N_2021,N_2078);
nand U2185 (N_2185,N_2025,N_2092);
nor U2186 (N_2186,N_2094,N_2057);
nor U2187 (N_2187,N_2013,N_2078);
nor U2188 (N_2188,N_2064,N_2030);
nor U2189 (N_2189,N_2068,N_2093);
nor U2190 (N_2190,N_2024,N_2027);
nand U2191 (N_2191,N_2086,N_2097);
nor U2192 (N_2192,N_2035,N_2059);
nor U2193 (N_2193,N_2056,N_2010);
and U2194 (N_2194,N_2021,N_2093);
nor U2195 (N_2195,N_2072,N_2085);
nand U2196 (N_2196,N_2035,N_2013);
or U2197 (N_2197,N_2035,N_2090);
or U2198 (N_2198,N_2036,N_2017);
nor U2199 (N_2199,N_2072,N_2038);
and U2200 (N_2200,N_2182,N_2176);
nand U2201 (N_2201,N_2168,N_2186);
and U2202 (N_2202,N_2181,N_2194);
nand U2203 (N_2203,N_2135,N_2132);
nand U2204 (N_2204,N_2122,N_2196);
and U2205 (N_2205,N_2187,N_2198);
or U2206 (N_2206,N_2179,N_2153);
and U2207 (N_2207,N_2162,N_2121);
or U2208 (N_2208,N_2103,N_2171);
nor U2209 (N_2209,N_2114,N_2126);
nand U2210 (N_2210,N_2124,N_2192);
or U2211 (N_2211,N_2151,N_2195);
and U2212 (N_2212,N_2111,N_2115);
or U2213 (N_2213,N_2112,N_2180);
nand U2214 (N_2214,N_2127,N_2144);
or U2215 (N_2215,N_2190,N_2150);
or U2216 (N_2216,N_2119,N_2154);
and U2217 (N_2217,N_2141,N_2128);
nand U2218 (N_2218,N_2133,N_2152);
and U2219 (N_2219,N_2110,N_2143);
nor U2220 (N_2220,N_2185,N_2172);
nor U2221 (N_2221,N_2167,N_2164);
and U2222 (N_2222,N_2170,N_2100);
or U2223 (N_2223,N_2120,N_2129);
nand U2224 (N_2224,N_2197,N_2136);
nor U2225 (N_2225,N_2130,N_2188);
and U2226 (N_2226,N_2161,N_2125);
and U2227 (N_2227,N_2173,N_2199);
nor U2228 (N_2228,N_2107,N_2157);
nor U2229 (N_2229,N_2166,N_2113);
nor U2230 (N_2230,N_2193,N_2175);
or U2231 (N_2231,N_2155,N_2137);
nand U2232 (N_2232,N_2108,N_2183);
nand U2233 (N_2233,N_2163,N_2148);
or U2234 (N_2234,N_2165,N_2131);
nand U2235 (N_2235,N_2177,N_2104);
nand U2236 (N_2236,N_2142,N_2191);
nand U2237 (N_2237,N_2147,N_2139);
nand U2238 (N_2238,N_2140,N_2189);
nor U2239 (N_2239,N_2146,N_2102);
nor U2240 (N_2240,N_2116,N_2174);
or U2241 (N_2241,N_2117,N_2106);
or U2242 (N_2242,N_2160,N_2149);
or U2243 (N_2243,N_2105,N_2101);
and U2244 (N_2244,N_2156,N_2138);
or U2245 (N_2245,N_2178,N_2158);
nor U2246 (N_2246,N_2123,N_2134);
nand U2247 (N_2247,N_2145,N_2159);
nor U2248 (N_2248,N_2169,N_2109);
nand U2249 (N_2249,N_2118,N_2184);
and U2250 (N_2250,N_2117,N_2134);
or U2251 (N_2251,N_2179,N_2122);
and U2252 (N_2252,N_2125,N_2182);
nand U2253 (N_2253,N_2184,N_2181);
nor U2254 (N_2254,N_2195,N_2191);
or U2255 (N_2255,N_2173,N_2198);
nand U2256 (N_2256,N_2188,N_2113);
nor U2257 (N_2257,N_2172,N_2141);
and U2258 (N_2258,N_2193,N_2173);
nand U2259 (N_2259,N_2152,N_2154);
nor U2260 (N_2260,N_2155,N_2199);
or U2261 (N_2261,N_2120,N_2100);
and U2262 (N_2262,N_2146,N_2167);
or U2263 (N_2263,N_2194,N_2127);
xor U2264 (N_2264,N_2167,N_2179);
or U2265 (N_2265,N_2102,N_2172);
or U2266 (N_2266,N_2196,N_2147);
nor U2267 (N_2267,N_2189,N_2172);
nand U2268 (N_2268,N_2161,N_2145);
nand U2269 (N_2269,N_2155,N_2102);
and U2270 (N_2270,N_2179,N_2196);
nor U2271 (N_2271,N_2111,N_2141);
nor U2272 (N_2272,N_2160,N_2161);
nor U2273 (N_2273,N_2138,N_2196);
nor U2274 (N_2274,N_2138,N_2166);
nor U2275 (N_2275,N_2139,N_2152);
nor U2276 (N_2276,N_2144,N_2148);
and U2277 (N_2277,N_2191,N_2104);
and U2278 (N_2278,N_2118,N_2178);
nand U2279 (N_2279,N_2163,N_2123);
nor U2280 (N_2280,N_2181,N_2139);
or U2281 (N_2281,N_2106,N_2103);
and U2282 (N_2282,N_2195,N_2170);
nand U2283 (N_2283,N_2172,N_2198);
or U2284 (N_2284,N_2112,N_2125);
nor U2285 (N_2285,N_2124,N_2162);
nand U2286 (N_2286,N_2156,N_2176);
nor U2287 (N_2287,N_2140,N_2119);
nor U2288 (N_2288,N_2158,N_2113);
nor U2289 (N_2289,N_2170,N_2145);
nor U2290 (N_2290,N_2161,N_2105);
nand U2291 (N_2291,N_2161,N_2169);
and U2292 (N_2292,N_2183,N_2181);
nor U2293 (N_2293,N_2121,N_2187);
or U2294 (N_2294,N_2129,N_2170);
nor U2295 (N_2295,N_2123,N_2169);
nand U2296 (N_2296,N_2138,N_2153);
and U2297 (N_2297,N_2157,N_2103);
or U2298 (N_2298,N_2118,N_2168);
nor U2299 (N_2299,N_2170,N_2176);
and U2300 (N_2300,N_2208,N_2282);
nand U2301 (N_2301,N_2224,N_2237);
or U2302 (N_2302,N_2291,N_2201);
nand U2303 (N_2303,N_2250,N_2242);
and U2304 (N_2304,N_2216,N_2219);
nand U2305 (N_2305,N_2234,N_2265);
and U2306 (N_2306,N_2248,N_2294);
and U2307 (N_2307,N_2232,N_2231);
nand U2308 (N_2308,N_2252,N_2200);
nor U2309 (N_2309,N_2257,N_2293);
and U2310 (N_2310,N_2285,N_2246);
and U2311 (N_2311,N_2278,N_2238);
nand U2312 (N_2312,N_2251,N_2255);
nor U2313 (N_2313,N_2207,N_2260);
and U2314 (N_2314,N_2262,N_2220);
nand U2315 (N_2315,N_2283,N_2245);
and U2316 (N_2316,N_2267,N_2281);
nor U2317 (N_2317,N_2206,N_2299);
nor U2318 (N_2318,N_2229,N_2214);
nor U2319 (N_2319,N_2249,N_2254);
nor U2320 (N_2320,N_2226,N_2259);
xnor U2321 (N_2321,N_2202,N_2211);
nand U2322 (N_2322,N_2236,N_2289);
nand U2323 (N_2323,N_2221,N_2290);
nand U2324 (N_2324,N_2209,N_2243);
nor U2325 (N_2325,N_2292,N_2258);
nand U2326 (N_2326,N_2217,N_2223);
or U2327 (N_2327,N_2205,N_2225);
or U2328 (N_2328,N_2230,N_2268);
or U2329 (N_2329,N_2222,N_2215);
nand U2330 (N_2330,N_2276,N_2244);
and U2331 (N_2331,N_2256,N_2263);
and U2332 (N_2332,N_2233,N_2261);
and U2333 (N_2333,N_2271,N_2213);
and U2334 (N_2334,N_2203,N_2235);
or U2335 (N_2335,N_2297,N_2296);
nor U2336 (N_2336,N_2228,N_2247);
or U2337 (N_2337,N_2295,N_2227);
nand U2338 (N_2338,N_2274,N_2269);
nand U2339 (N_2339,N_2204,N_2273);
or U2340 (N_2340,N_2298,N_2272);
or U2341 (N_2341,N_2253,N_2279);
and U2342 (N_2342,N_2264,N_2266);
or U2343 (N_2343,N_2277,N_2240);
or U2344 (N_2344,N_2210,N_2270);
nand U2345 (N_2345,N_2288,N_2284);
nor U2346 (N_2346,N_2275,N_2239);
and U2347 (N_2347,N_2241,N_2287);
or U2348 (N_2348,N_2218,N_2212);
and U2349 (N_2349,N_2280,N_2286);
xor U2350 (N_2350,N_2277,N_2282);
nand U2351 (N_2351,N_2209,N_2281);
or U2352 (N_2352,N_2205,N_2203);
and U2353 (N_2353,N_2281,N_2218);
xor U2354 (N_2354,N_2201,N_2228);
nand U2355 (N_2355,N_2263,N_2258);
or U2356 (N_2356,N_2291,N_2208);
or U2357 (N_2357,N_2289,N_2229);
or U2358 (N_2358,N_2254,N_2206);
and U2359 (N_2359,N_2258,N_2267);
nand U2360 (N_2360,N_2279,N_2248);
or U2361 (N_2361,N_2215,N_2216);
and U2362 (N_2362,N_2270,N_2266);
or U2363 (N_2363,N_2238,N_2297);
or U2364 (N_2364,N_2292,N_2273);
nand U2365 (N_2365,N_2233,N_2279);
or U2366 (N_2366,N_2255,N_2237);
or U2367 (N_2367,N_2237,N_2223);
nand U2368 (N_2368,N_2219,N_2218);
nor U2369 (N_2369,N_2217,N_2296);
nor U2370 (N_2370,N_2238,N_2262);
and U2371 (N_2371,N_2282,N_2274);
nor U2372 (N_2372,N_2242,N_2254);
nand U2373 (N_2373,N_2294,N_2273);
nor U2374 (N_2374,N_2221,N_2229);
nand U2375 (N_2375,N_2218,N_2277);
and U2376 (N_2376,N_2263,N_2212);
nand U2377 (N_2377,N_2204,N_2232);
and U2378 (N_2378,N_2296,N_2289);
and U2379 (N_2379,N_2220,N_2278);
and U2380 (N_2380,N_2287,N_2203);
and U2381 (N_2381,N_2257,N_2295);
nand U2382 (N_2382,N_2261,N_2248);
and U2383 (N_2383,N_2233,N_2259);
nand U2384 (N_2384,N_2271,N_2203);
nand U2385 (N_2385,N_2262,N_2259);
or U2386 (N_2386,N_2239,N_2244);
nand U2387 (N_2387,N_2208,N_2210);
nor U2388 (N_2388,N_2226,N_2289);
nor U2389 (N_2389,N_2256,N_2251);
or U2390 (N_2390,N_2246,N_2293);
or U2391 (N_2391,N_2243,N_2248);
nor U2392 (N_2392,N_2283,N_2296);
nor U2393 (N_2393,N_2208,N_2222);
and U2394 (N_2394,N_2253,N_2252);
nor U2395 (N_2395,N_2280,N_2229);
nand U2396 (N_2396,N_2245,N_2296);
nand U2397 (N_2397,N_2216,N_2232);
xnor U2398 (N_2398,N_2203,N_2247);
nand U2399 (N_2399,N_2243,N_2213);
nor U2400 (N_2400,N_2357,N_2316);
nand U2401 (N_2401,N_2376,N_2332);
or U2402 (N_2402,N_2382,N_2328);
or U2403 (N_2403,N_2396,N_2300);
or U2404 (N_2404,N_2341,N_2363);
nor U2405 (N_2405,N_2365,N_2393);
and U2406 (N_2406,N_2339,N_2317);
or U2407 (N_2407,N_2353,N_2348);
nand U2408 (N_2408,N_2346,N_2347);
nor U2409 (N_2409,N_2337,N_2399);
xnor U2410 (N_2410,N_2319,N_2338);
nand U2411 (N_2411,N_2358,N_2342);
nand U2412 (N_2412,N_2318,N_2307);
or U2413 (N_2413,N_2374,N_2373);
nor U2414 (N_2414,N_2364,N_2370);
nand U2415 (N_2415,N_2372,N_2359);
and U2416 (N_2416,N_2313,N_2312);
or U2417 (N_2417,N_2394,N_2384);
or U2418 (N_2418,N_2375,N_2361);
or U2419 (N_2419,N_2360,N_2344);
nor U2420 (N_2420,N_2336,N_2349);
and U2421 (N_2421,N_2322,N_2371);
nand U2422 (N_2422,N_2321,N_2330);
nor U2423 (N_2423,N_2326,N_2323);
and U2424 (N_2424,N_2308,N_2383);
and U2425 (N_2425,N_2380,N_2356);
and U2426 (N_2426,N_2389,N_2355);
nand U2427 (N_2427,N_2390,N_2302);
or U2428 (N_2428,N_2367,N_2352);
and U2429 (N_2429,N_2320,N_2331);
or U2430 (N_2430,N_2304,N_2362);
nand U2431 (N_2431,N_2381,N_2354);
nor U2432 (N_2432,N_2377,N_2350);
nor U2433 (N_2433,N_2369,N_2315);
nor U2434 (N_2434,N_2309,N_2386);
or U2435 (N_2435,N_2305,N_2340);
and U2436 (N_2436,N_2397,N_2345);
or U2437 (N_2437,N_2391,N_2311);
and U2438 (N_2438,N_2324,N_2392);
nand U2439 (N_2439,N_2314,N_2327);
nor U2440 (N_2440,N_2303,N_2378);
or U2441 (N_2441,N_2351,N_2366);
and U2442 (N_2442,N_2368,N_2387);
nor U2443 (N_2443,N_2398,N_2388);
and U2444 (N_2444,N_2306,N_2335);
or U2445 (N_2445,N_2395,N_2325);
and U2446 (N_2446,N_2301,N_2334);
or U2447 (N_2447,N_2343,N_2385);
and U2448 (N_2448,N_2333,N_2329);
or U2449 (N_2449,N_2379,N_2310);
nand U2450 (N_2450,N_2341,N_2374);
and U2451 (N_2451,N_2352,N_2364);
and U2452 (N_2452,N_2324,N_2303);
or U2453 (N_2453,N_2335,N_2364);
or U2454 (N_2454,N_2363,N_2305);
and U2455 (N_2455,N_2310,N_2315);
or U2456 (N_2456,N_2394,N_2340);
and U2457 (N_2457,N_2332,N_2384);
and U2458 (N_2458,N_2387,N_2356);
xnor U2459 (N_2459,N_2385,N_2314);
or U2460 (N_2460,N_2310,N_2396);
nand U2461 (N_2461,N_2399,N_2307);
nand U2462 (N_2462,N_2306,N_2328);
and U2463 (N_2463,N_2346,N_2360);
or U2464 (N_2464,N_2304,N_2335);
or U2465 (N_2465,N_2318,N_2385);
and U2466 (N_2466,N_2341,N_2308);
nand U2467 (N_2467,N_2358,N_2313);
nand U2468 (N_2468,N_2348,N_2305);
and U2469 (N_2469,N_2349,N_2367);
and U2470 (N_2470,N_2351,N_2321);
nor U2471 (N_2471,N_2399,N_2379);
nor U2472 (N_2472,N_2346,N_2323);
nand U2473 (N_2473,N_2374,N_2394);
nand U2474 (N_2474,N_2374,N_2347);
and U2475 (N_2475,N_2338,N_2343);
and U2476 (N_2476,N_2323,N_2338);
nor U2477 (N_2477,N_2334,N_2327);
or U2478 (N_2478,N_2351,N_2395);
nor U2479 (N_2479,N_2362,N_2356);
or U2480 (N_2480,N_2395,N_2312);
and U2481 (N_2481,N_2388,N_2393);
nand U2482 (N_2482,N_2392,N_2374);
nor U2483 (N_2483,N_2325,N_2391);
or U2484 (N_2484,N_2357,N_2387);
nand U2485 (N_2485,N_2348,N_2374);
nor U2486 (N_2486,N_2321,N_2304);
nor U2487 (N_2487,N_2393,N_2367);
nand U2488 (N_2488,N_2332,N_2300);
nor U2489 (N_2489,N_2320,N_2347);
nand U2490 (N_2490,N_2379,N_2331);
or U2491 (N_2491,N_2361,N_2353);
nand U2492 (N_2492,N_2387,N_2317);
or U2493 (N_2493,N_2361,N_2329);
nand U2494 (N_2494,N_2341,N_2362);
nor U2495 (N_2495,N_2396,N_2344);
nand U2496 (N_2496,N_2385,N_2350);
nor U2497 (N_2497,N_2372,N_2349);
nand U2498 (N_2498,N_2310,N_2359);
or U2499 (N_2499,N_2311,N_2370);
or U2500 (N_2500,N_2413,N_2403);
and U2501 (N_2501,N_2459,N_2499);
nand U2502 (N_2502,N_2409,N_2492);
and U2503 (N_2503,N_2461,N_2429);
and U2504 (N_2504,N_2471,N_2469);
or U2505 (N_2505,N_2462,N_2473);
or U2506 (N_2506,N_2416,N_2440);
nand U2507 (N_2507,N_2453,N_2447);
nor U2508 (N_2508,N_2478,N_2423);
and U2509 (N_2509,N_2466,N_2442);
or U2510 (N_2510,N_2415,N_2483);
nand U2511 (N_2511,N_2475,N_2428);
or U2512 (N_2512,N_2407,N_2420);
or U2513 (N_2513,N_2401,N_2460);
or U2514 (N_2514,N_2439,N_2422);
nand U2515 (N_2515,N_2463,N_2402);
nor U2516 (N_2516,N_2497,N_2456);
nand U2517 (N_2517,N_2465,N_2406);
nand U2518 (N_2518,N_2446,N_2437);
nand U2519 (N_2519,N_2432,N_2411);
and U2520 (N_2520,N_2477,N_2484);
or U2521 (N_2521,N_2457,N_2464);
nand U2522 (N_2522,N_2436,N_2489);
or U2523 (N_2523,N_2410,N_2425);
nor U2524 (N_2524,N_2458,N_2467);
nor U2525 (N_2525,N_2498,N_2400);
xor U2526 (N_2526,N_2449,N_2485);
and U2527 (N_2527,N_2490,N_2433);
nand U2528 (N_2528,N_2496,N_2414);
or U2529 (N_2529,N_2444,N_2408);
nand U2530 (N_2530,N_2405,N_2486);
nor U2531 (N_2531,N_2452,N_2482);
nand U2532 (N_2532,N_2427,N_2443);
or U2533 (N_2533,N_2424,N_2404);
nor U2534 (N_2534,N_2417,N_2448);
or U2535 (N_2535,N_2430,N_2450);
and U2536 (N_2536,N_2434,N_2470);
nand U2537 (N_2537,N_2476,N_2472);
or U2538 (N_2538,N_2445,N_2474);
and U2539 (N_2539,N_2493,N_2480);
or U2540 (N_2540,N_2481,N_2441);
and U2541 (N_2541,N_2426,N_2438);
nor U2542 (N_2542,N_2495,N_2468);
nor U2543 (N_2543,N_2491,N_2435);
nand U2544 (N_2544,N_2454,N_2412);
and U2545 (N_2545,N_2419,N_2431);
and U2546 (N_2546,N_2488,N_2421);
nand U2547 (N_2547,N_2455,N_2418);
nand U2548 (N_2548,N_2479,N_2494);
nor U2549 (N_2549,N_2451,N_2487);
or U2550 (N_2550,N_2454,N_2409);
nor U2551 (N_2551,N_2464,N_2407);
nor U2552 (N_2552,N_2403,N_2441);
and U2553 (N_2553,N_2448,N_2406);
and U2554 (N_2554,N_2434,N_2492);
nand U2555 (N_2555,N_2453,N_2498);
nor U2556 (N_2556,N_2452,N_2421);
or U2557 (N_2557,N_2482,N_2445);
nand U2558 (N_2558,N_2444,N_2488);
nor U2559 (N_2559,N_2499,N_2424);
or U2560 (N_2560,N_2487,N_2475);
nand U2561 (N_2561,N_2447,N_2422);
nor U2562 (N_2562,N_2434,N_2450);
nand U2563 (N_2563,N_2407,N_2440);
or U2564 (N_2564,N_2458,N_2486);
nor U2565 (N_2565,N_2463,N_2459);
or U2566 (N_2566,N_2418,N_2493);
or U2567 (N_2567,N_2482,N_2462);
nand U2568 (N_2568,N_2493,N_2464);
nor U2569 (N_2569,N_2438,N_2472);
nor U2570 (N_2570,N_2473,N_2492);
and U2571 (N_2571,N_2475,N_2423);
nor U2572 (N_2572,N_2452,N_2426);
and U2573 (N_2573,N_2459,N_2489);
nor U2574 (N_2574,N_2476,N_2466);
nand U2575 (N_2575,N_2463,N_2410);
or U2576 (N_2576,N_2407,N_2488);
nor U2577 (N_2577,N_2489,N_2446);
nand U2578 (N_2578,N_2439,N_2499);
nand U2579 (N_2579,N_2480,N_2403);
nor U2580 (N_2580,N_2439,N_2452);
and U2581 (N_2581,N_2482,N_2402);
or U2582 (N_2582,N_2449,N_2457);
xnor U2583 (N_2583,N_2405,N_2432);
nand U2584 (N_2584,N_2475,N_2439);
nor U2585 (N_2585,N_2461,N_2477);
and U2586 (N_2586,N_2469,N_2419);
nand U2587 (N_2587,N_2458,N_2412);
and U2588 (N_2588,N_2451,N_2448);
nand U2589 (N_2589,N_2400,N_2453);
nor U2590 (N_2590,N_2437,N_2489);
or U2591 (N_2591,N_2473,N_2450);
nand U2592 (N_2592,N_2408,N_2474);
nand U2593 (N_2593,N_2410,N_2497);
xor U2594 (N_2594,N_2432,N_2495);
or U2595 (N_2595,N_2460,N_2442);
nor U2596 (N_2596,N_2479,N_2400);
and U2597 (N_2597,N_2492,N_2441);
nor U2598 (N_2598,N_2423,N_2487);
nand U2599 (N_2599,N_2469,N_2472);
nor U2600 (N_2600,N_2508,N_2524);
or U2601 (N_2601,N_2587,N_2591);
nand U2602 (N_2602,N_2529,N_2550);
nand U2603 (N_2603,N_2528,N_2553);
nand U2604 (N_2604,N_2581,N_2560);
nor U2605 (N_2605,N_2584,N_2505);
nor U2606 (N_2606,N_2547,N_2596);
nor U2607 (N_2607,N_2548,N_2551);
and U2608 (N_2608,N_2506,N_2582);
nand U2609 (N_2609,N_2503,N_2579);
and U2610 (N_2610,N_2535,N_2507);
nand U2611 (N_2611,N_2564,N_2549);
nor U2612 (N_2612,N_2565,N_2588);
nand U2613 (N_2613,N_2570,N_2557);
nand U2614 (N_2614,N_2578,N_2554);
or U2615 (N_2615,N_2522,N_2538);
or U2616 (N_2616,N_2527,N_2531);
nand U2617 (N_2617,N_2530,N_2519);
and U2618 (N_2618,N_2501,N_2574);
nand U2619 (N_2619,N_2563,N_2572);
or U2620 (N_2620,N_2543,N_2515);
or U2621 (N_2621,N_2556,N_2580);
nand U2622 (N_2622,N_2562,N_2592);
nand U2623 (N_2623,N_2567,N_2537);
or U2624 (N_2624,N_2552,N_2504);
nor U2625 (N_2625,N_2517,N_2534);
or U2626 (N_2626,N_2594,N_2571);
or U2627 (N_2627,N_2509,N_2546);
or U2628 (N_2628,N_2595,N_2577);
or U2629 (N_2629,N_2502,N_2576);
and U2630 (N_2630,N_2518,N_2541);
or U2631 (N_2631,N_2512,N_2569);
nor U2632 (N_2632,N_2510,N_2568);
nand U2633 (N_2633,N_2589,N_2516);
nand U2634 (N_2634,N_2521,N_2544);
nor U2635 (N_2635,N_2500,N_2599);
nor U2636 (N_2636,N_2511,N_2542);
nand U2637 (N_2637,N_2520,N_2539);
nand U2638 (N_2638,N_2575,N_2558);
and U2639 (N_2639,N_2583,N_2590);
nor U2640 (N_2640,N_2598,N_2525);
nor U2641 (N_2641,N_2533,N_2593);
and U2642 (N_2642,N_2559,N_2597);
and U2643 (N_2643,N_2523,N_2573);
and U2644 (N_2644,N_2540,N_2514);
nor U2645 (N_2645,N_2561,N_2555);
and U2646 (N_2646,N_2585,N_2513);
nor U2647 (N_2647,N_2586,N_2566);
and U2648 (N_2648,N_2526,N_2532);
and U2649 (N_2649,N_2545,N_2536);
nor U2650 (N_2650,N_2508,N_2561);
and U2651 (N_2651,N_2529,N_2589);
nor U2652 (N_2652,N_2540,N_2549);
nand U2653 (N_2653,N_2504,N_2555);
nand U2654 (N_2654,N_2527,N_2505);
nor U2655 (N_2655,N_2517,N_2562);
or U2656 (N_2656,N_2541,N_2531);
nand U2657 (N_2657,N_2587,N_2539);
xnor U2658 (N_2658,N_2587,N_2548);
and U2659 (N_2659,N_2511,N_2594);
nand U2660 (N_2660,N_2537,N_2535);
or U2661 (N_2661,N_2573,N_2594);
and U2662 (N_2662,N_2579,N_2593);
and U2663 (N_2663,N_2518,N_2528);
nor U2664 (N_2664,N_2540,N_2542);
or U2665 (N_2665,N_2538,N_2586);
or U2666 (N_2666,N_2565,N_2544);
nand U2667 (N_2667,N_2566,N_2503);
and U2668 (N_2668,N_2584,N_2533);
nor U2669 (N_2669,N_2575,N_2525);
or U2670 (N_2670,N_2535,N_2545);
and U2671 (N_2671,N_2593,N_2598);
nand U2672 (N_2672,N_2599,N_2531);
and U2673 (N_2673,N_2541,N_2573);
nand U2674 (N_2674,N_2546,N_2541);
or U2675 (N_2675,N_2589,N_2519);
or U2676 (N_2676,N_2545,N_2565);
and U2677 (N_2677,N_2553,N_2531);
or U2678 (N_2678,N_2583,N_2544);
nor U2679 (N_2679,N_2540,N_2548);
or U2680 (N_2680,N_2552,N_2540);
or U2681 (N_2681,N_2507,N_2583);
nor U2682 (N_2682,N_2529,N_2502);
and U2683 (N_2683,N_2593,N_2524);
nor U2684 (N_2684,N_2524,N_2521);
or U2685 (N_2685,N_2514,N_2535);
and U2686 (N_2686,N_2564,N_2570);
nor U2687 (N_2687,N_2598,N_2510);
or U2688 (N_2688,N_2591,N_2507);
nand U2689 (N_2689,N_2552,N_2546);
and U2690 (N_2690,N_2596,N_2550);
nand U2691 (N_2691,N_2534,N_2587);
and U2692 (N_2692,N_2540,N_2583);
nand U2693 (N_2693,N_2506,N_2597);
or U2694 (N_2694,N_2521,N_2530);
nor U2695 (N_2695,N_2549,N_2505);
nor U2696 (N_2696,N_2582,N_2519);
or U2697 (N_2697,N_2583,N_2586);
nor U2698 (N_2698,N_2586,N_2547);
nor U2699 (N_2699,N_2526,N_2597);
or U2700 (N_2700,N_2636,N_2686);
nor U2701 (N_2701,N_2655,N_2677);
nand U2702 (N_2702,N_2666,N_2600);
nor U2703 (N_2703,N_2695,N_2626);
or U2704 (N_2704,N_2649,N_2633);
and U2705 (N_2705,N_2652,N_2604);
or U2706 (N_2706,N_2643,N_2673);
nand U2707 (N_2707,N_2699,N_2618);
or U2708 (N_2708,N_2610,N_2692);
and U2709 (N_2709,N_2653,N_2627);
and U2710 (N_2710,N_2608,N_2651);
and U2711 (N_2711,N_2609,N_2620);
or U2712 (N_2712,N_2662,N_2638);
nor U2713 (N_2713,N_2697,N_2661);
nand U2714 (N_2714,N_2683,N_2664);
and U2715 (N_2715,N_2696,N_2650);
or U2716 (N_2716,N_2622,N_2623);
and U2717 (N_2717,N_2682,N_2624);
and U2718 (N_2718,N_2690,N_2634);
nand U2719 (N_2719,N_2637,N_2679);
and U2720 (N_2720,N_2607,N_2644);
nand U2721 (N_2721,N_2648,N_2681);
or U2722 (N_2722,N_2641,N_2605);
nand U2723 (N_2723,N_2630,N_2606);
or U2724 (N_2724,N_2680,N_2611);
nand U2725 (N_2725,N_2656,N_2640);
nor U2726 (N_2726,N_2629,N_2659);
and U2727 (N_2727,N_2635,N_2668);
or U2728 (N_2728,N_2689,N_2621);
or U2729 (N_2729,N_2672,N_2687);
nand U2730 (N_2730,N_2675,N_2601);
xor U2731 (N_2731,N_2658,N_2645);
nor U2732 (N_2732,N_2613,N_2614);
and U2733 (N_2733,N_2669,N_2693);
nand U2734 (N_2734,N_2676,N_2617);
nor U2735 (N_2735,N_2642,N_2674);
or U2736 (N_2736,N_2628,N_2678);
nand U2737 (N_2737,N_2663,N_2685);
nor U2738 (N_2738,N_2667,N_2602);
nand U2739 (N_2739,N_2625,N_2670);
nand U2740 (N_2740,N_2660,N_2688);
nor U2741 (N_2741,N_2694,N_2616);
and U2742 (N_2742,N_2691,N_2671);
nor U2743 (N_2743,N_2684,N_2615);
or U2744 (N_2744,N_2646,N_2657);
or U2745 (N_2745,N_2632,N_2647);
or U2746 (N_2746,N_2639,N_2603);
nand U2747 (N_2747,N_2619,N_2698);
or U2748 (N_2748,N_2612,N_2631);
nor U2749 (N_2749,N_2654,N_2665);
nand U2750 (N_2750,N_2684,N_2699);
nor U2751 (N_2751,N_2656,N_2625);
nand U2752 (N_2752,N_2653,N_2615);
nand U2753 (N_2753,N_2600,N_2623);
nor U2754 (N_2754,N_2621,N_2690);
nand U2755 (N_2755,N_2617,N_2651);
nand U2756 (N_2756,N_2667,N_2614);
and U2757 (N_2757,N_2635,N_2684);
nand U2758 (N_2758,N_2657,N_2661);
or U2759 (N_2759,N_2684,N_2664);
or U2760 (N_2760,N_2632,N_2611);
and U2761 (N_2761,N_2668,N_2699);
and U2762 (N_2762,N_2651,N_2669);
or U2763 (N_2763,N_2661,N_2651);
nor U2764 (N_2764,N_2673,N_2630);
or U2765 (N_2765,N_2686,N_2613);
or U2766 (N_2766,N_2638,N_2631);
nor U2767 (N_2767,N_2665,N_2632);
or U2768 (N_2768,N_2606,N_2649);
nor U2769 (N_2769,N_2650,N_2618);
or U2770 (N_2770,N_2695,N_2623);
nand U2771 (N_2771,N_2665,N_2662);
nand U2772 (N_2772,N_2621,N_2662);
nand U2773 (N_2773,N_2618,N_2691);
nor U2774 (N_2774,N_2681,N_2612);
xnor U2775 (N_2775,N_2611,N_2688);
and U2776 (N_2776,N_2619,N_2674);
or U2777 (N_2777,N_2607,N_2624);
or U2778 (N_2778,N_2671,N_2690);
nand U2779 (N_2779,N_2633,N_2642);
nand U2780 (N_2780,N_2696,N_2631);
or U2781 (N_2781,N_2685,N_2697);
nor U2782 (N_2782,N_2602,N_2625);
and U2783 (N_2783,N_2683,N_2620);
or U2784 (N_2784,N_2699,N_2608);
or U2785 (N_2785,N_2685,N_2617);
and U2786 (N_2786,N_2611,N_2657);
or U2787 (N_2787,N_2652,N_2682);
nand U2788 (N_2788,N_2672,N_2682);
or U2789 (N_2789,N_2641,N_2603);
and U2790 (N_2790,N_2601,N_2605);
or U2791 (N_2791,N_2646,N_2649);
and U2792 (N_2792,N_2621,N_2687);
nor U2793 (N_2793,N_2630,N_2678);
and U2794 (N_2794,N_2651,N_2690);
or U2795 (N_2795,N_2617,N_2672);
and U2796 (N_2796,N_2668,N_2652);
nor U2797 (N_2797,N_2617,N_2606);
and U2798 (N_2798,N_2639,N_2646);
nor U2799 (N_2799,N_2694,N_2666);
and U2800 (N_2800,N_2735,N_2750);
or U2801 (N_2801,N_2749,N_2725);
nor U2802 (N_2802,N_2779,N_2763);
and U2803 (N_2803,N_2777,N_2790);
nor U2804 (N_2804,N_2738,N_2797);
nor U2805 (N_2805,N_2716,N_2767);
nor U2806 (N_2806,N_2791,N_2719);
nor U2807 (N_2807,N_2727,N_2713);
and U2808 (N_2808,N_2705,N_2785);
and U2809 (N_2809,N_2778,N_2742);
nor U2810 (N_2810,N_2703,N_2771);
nor U2811 (N_2811,N_2783,N_2766);
nor U2812 (N_2812,N_2711,N_2709);
and U2813 (N_2813,N_2700,N_2724);
and U2814 (N_2814,N_2758,N_2752);
nand U2815 (N_2815,N_2747,N_2755);
nand U2816 (N_2816,N_2780,N_2781);
or U2817 (N_2817,N_2708,N_2710);
or U2818 (N_2818,N_2794,N_2726);
nand U2819 (N_2819,N_2731,N_2718);
nor U2820 (N_2820,N_2744,N_2789);
nor U2821 (N_2821,N_2796,N_2740);
or U2822 (N_2822,N_2756,N_2760);
nor U2823 (N_2823,N_2736,N_2764);
and U2824 (N_2824,N_2774,N_2714);
or U2825 (N_2825,N_2765,N_2745);
nor U2826 (N_2826,N_2720,N_2776);
and U2827 (N_2827,N_2773,N_2786);
nand U2828 (N_2828,N_2704,N_2723);
or U2829 (N_2829,N_2772,N_2702);
and U2830 (N_2830,N_2782,N_2754);
nand U2831 (N_2831,N_2739,N_2769);
nand U2832 (N_2832,N_2715,N_2712);
nor U2833 (N_2833,N_2721,N_2741);
or U2834 (N_2834,N_2706,N_2730);
nand U2835 (N_2835,N_2746,N_2761);
or U2836 (N_2836,N_2748,N_2751);
and U2837 (N_2837,N_2734,N_2737);
xor U2838 (N_2838,N_2707,N_2775);
nor U2839 (N_2839,N_2753,N_2722);
or U2840 (N_2840,N_2762,N_2733);
or U2841 (N_2841,N_2732,N_2792);
or U2842 (N_2842,N_2768,N_2757);
nor U2843 (N_2843,N_2798,N_2787);
or U2844 (N_2844,N_2728,N_2701);
nor U2845 (N_2845,N_2759,N_2793);
or U2846 (N_2846,N_2743,N_2799);
nor U2847 (N_2847,N_2770,N_2795);
nand U2848 (N_2848,N_2729,N_2717);
nand U2849 (N_2849,N_2784,N_2788);
and U2850 (N_2850,N_2727,N_2756);
and U2851 (N_2851,N_2768,N_2764);
and U2852 (N_2852,N_2728,N_2772);
or U2853 (N_2853,N_2746,N_2792);
and U2854 (N_2854,N_2735,N_2783);
nand U2855 (N_2855,N_2742,N_2724);
nand U2856 (N_2856,N_2760,N_2731);
and U2857 (N_2857,N_2729,N_2771);
and U2858 (N_2858,N_2730,N_2788);
or U2859 (N_2859,N_2772,N_2776);
nand U2860 (N_2860,N_2726,N_2769);
or U2861 (N_2861,N_2770,N_2769);
or U2862 (N_2862,N_2708,N_2702);
or U2863 (N_2863,N_2744,N_2787);
or U2864 (N_2864,N_2786,N_2776);
and U2865 (N_2865,N_2704,N_2795);
or U2866 (N_2866,N_2724,N_2711);
nand U2867 (N_2867,N_2724,N_2765);
and U2868 (N_2868,N_2758,N_2777);
and U2869 (N_2869,N_2782,N_2746);
and U2870 (N_2870,N_2723,N_2738);
nor U2871 (N_2871,N_2778,N_2737);
nand U2872 (N_2872,N_2703,N_2700);
and U2873 (N_2873,N_2774,N_2770);
and U2874 (N_2874,N_2734,N_2768);
and U2875 (N_2875,N_2704,N_2789);
nor U2876 (N_2876,N_2793,N_2774);
and U2877 (N_2877,N_2793,N_2755);
and U2878 (N_2878,N_2773,N_2751);
nor U2879 (N_2879,N_2740,N_2719);
or U2880 (N_2880,N_2708,N_2798);
or U2881 (N_2881,N_2786,N_2734);
and U2882 (N_2882,N_2746,N_2726);
nor U2883 (N_2883,N_2726,N_2783);
and U2884 (N_2884,N_2767,N_2770);
nor U2885 (N_2885,N_2728,N_2731);
or U2886 (N_2886,N_2767,N_2798);
nand U2887 (N_2887,N_2784,N_2785);
or U2888 (N_2888,N_2766,N_2782);
and U2889 (N_2889,N_2769,N_2719);
and U2890 (N_2890,N_2727,N_2795);
and U2891 (N_2891,N_2744,N_2763);
or U2892 (N_2892,N_2758,N_2782);
nor U2893 (N_2893,N_2749,N_2770);
and U2894 (N_2894,N_2703,N_2794);
or U2895 (N_2895,N_2794,N_2775);
nand U2896 (N_2896,N_2766,N_2770);
nand U2897 (N_2897,N_2711,N_2712);
nand U2898 (N_2898,N_2703,N_2746);
nand U2899 (N_2899,N_2734,N_2749);
nand U2900 (N_2900,N_2805,N_2826);
nor U2901 (N_2901,N_2854,N_2845);
or U2902 (N_2902,N_2884,N_2861);
nor U2903 (N_2903,N_2887,N_2892);
and U2904 (N_2904,N_2831,N_2853);
nand U2905 (N_2905,N_2875,N_2891);
or U2906 (N_2906,N_2877,N_2852);
xnor U2907 (N_2907,N_2881,N_2866);
or U2908 (N_2908,N_2888,N_2872);
and U2909 (N_2909,N_2862,N_2815);
and U2910 (N_2910,N_2812,N_2844);
nand U2911 (N_2911,N_2898,N_2878);
and U2912 (N_2912,N_2802,N_2827);
or U2913 (N_2913,N_2829,N_2803);
nor U2914 (N_2914,N_2868,N_2897);
and U2915 (N_2915,N_2836,N_2810);
nor U2916 (N_2916,N_2804,N_2816);
nand U2917 (N_2917,N_2842,N_2830);
and U2918 (N_2918,N_2806,N_2859);
nor U2919 (N_2919,N_2819,N_2896);
and U2920 (N_2920,N_2869,N_2801);
or U2921 (N_2921,N_2835,N_2874);
nand U2922 (N_2922,N_2886,N_2864);
nand U2923 (N_2923,N_2840,N_2857);
and U2924 (N_2924,N_2825,N_2846);
nor U2925 (N_2925,N_2848,N_2837);
or U2926 (N_2926,N_2843,N_2832);
and U2927 (N_2927,N_2871,N_2885);
nand U2928 (N_2928,N_2820,N_2899);
and U2929 (N_2929,N_2809,N_2823);
nand U2930 (N_2930,N_2876,N_2847);
and U2931 (N_2931,N_2851,N_2849);
nand U2932 (N_2932,N_2824,N_2860);
and U2933 (N_2933,N_2822,N_2811);
nor U2934 (N_2934,N_2856,N_2870);
or U2935 (N_2935,N_2818,N_2873);
or U2936 (N_2936,N_2850,N_2807);
and U2937 (N_2937,N_2863,N_2889);
and U2938 (N_2938,N_2858,N_2883);
or U2939 (N_2939,N_2880,N_2814);
and U2940 (N_2940,N_2839,N_2841);
nand U2941 (N_2941,N_2838,N_2855);
nor U2942 (N_2942,N_2894,N_2834);
nand U2943 (N_2943,N_2821,N_2882);
nand U2944 (N_2944,N_2813,N_2808);
nor U2945 (N_2945,N_2865,N_2833);
and U2946 (N_2946,N_2895,N_2800);
nor U2947 (N_2947,N_2879,N_2893);
nand U2948 (N_2948,N_2828,N_2890);
nand U2949 (N_2949,N_2867,N_2817);
or U2950 (N_2950,N_2899,N_2841);
nor U2951 (N_2951,N_2805,N_2809);
or U2952 (N_2952,N_2868,N_2812);
or U2953 (N_2953,N_2860,N_2813);
nor U2954 (N_2954,N_2872,N_2855);
or U2955 (N_2955,N_2856,N_2877);
or U2956 (N_2956,N_2869,N_2831);
nor U2957 (N_2957,N_2877,N_2883);
nand U2958 (N_2958,N_2835,N_2859);
nand U2959 (N_2959,N_2884,N_2859);
nand U2960 (N_2960,N_2868,N_2875);
nand U2961 (N_2961,N_2812,N_2898);
or U2962 (N_2962,N_2848,N_2814);
nor U2963 (N_2963,N_2882,N_2852);
and U2964 (N_2964,N_2800,N_2841);
nand U2965 (N_2965,N_2817,N_2888);
nand U2966 (N_2966,N_2833,N_2800);
and U2967 (N_2967,N_2867,N_2805);
or U2968 (N_2968,N_2887,N_2816);
and U2969 (N_2969,N_2879,N_2841);
and U2970 (N_2970,N_2886,N_2812);
or U2971 (N_2971,N_2853,N_2898);
and U2972 (N_2972,N_2815,N_2857);
or U2973 (N_2973,N_2801,N_2885);
or U2974 (N_2974,N_2840,N_2802);
and U2975 (N_2975,N_2894,N_2814);
or U2976 (N_2976,N_2813,N_2877);
and U2977 (N_2977,N_2817,N_2851);
and U2978 (N_2978,N_2835,N_2800);
and U2979 (N_2979,N_2894,N_2846);
and U2980 (N_2980,N_2802,N_2890);
or U2981 (N_2981,N_2889,N_2871);
nor U2982 (N_2982,N_2804,N_2872);
nand U2983 (N_2983,N_2814,N_2841);
nor U2984 (N_2984,N_2825,N_2829);
nand U2985 (N_2985,N_2843,N_2824);
and U2986 (N_2986,N_2806,N_2888);
or U2987 (N_2987,N_2898,N_2806);
nor U2988 (N_2988,N_2815,N_2848);
nand U2989 (N_2989,N_2805,N_2894);
and U2990 (N_2990,N_2818,N_2809);
and U2991 (N_2991,N_2880,N_2816);
or U2992 (N_2992,N_2892,N_2846);
nor U2993 (N_2993,N_2887,N_2831);
nand U2994 (N_2994,N_2856,N_2866);
or U2995 (N_2995,N_2869,N_2837);
or U2996 (N_2996,N_2892,N_2865);
or U2997 (N_2997,N_2821,N_2806);
nand U2998 (N_2998,N_2884,N_2837);
or U2999 (N_2999,N_2802,N_2888);
nand UO_0 (O_0,N_2968,N_2907);
nand UO_1 (O_1,N_2964,N_2962);
and UO_2 (O_2,N_2915,N_2965);
nand UO_3 (O_3,N_2989,N_2997);
or UO_4 (O_4,N_2992,N_2945);
nand UO_5 (O_5,N_2970,N_2912);
or UO_6 (O_6,N_2981,N_2908);
and UO_7 (O_7,N_2969,N_2914);
or UO_8 (O_8,N_2988,N_2937);
nand UO_9 (O_9,N_2961,N_2949);
and UO_10 (O_10,N_2947,N_2923);
and UO_11 (O_11,N_2932,N_2938);
nand UO_12 (O_12,N_2951,N_2903);
nand UO_13 (O_13,N_2979,N_2921);
nand UO_14 (O_14,N_2924,N_2943);
or UO_15 (O_15,N_2955,N_2925);
nor UO_16 (O_16,N_2948,N_2952);
nor UO_17 (O_17,N_2919,N_2976);
nor UO_18 (O_18,N_2933,N_2995);
and UO_19 (O_19,N_2930,N_2927);
nand UO_20 (O_20,N_2985,N_2906);
nand UO_21 (O_21,N_2958,N_2905);
nand UO_22 (O_22,N_2986,N_2918);
or UO_23 (O_23,N_2956,N_2998);
and UO_24 (O_24,N_2913,N_2996);
nand UO_25 (O_25,N_2939,N_2994);
and UO_26 (O_26,N_2922,N_2910);
nand UO_27 (O_27,N_2987,N_2917);
or UO_28 (O_28,N_2901,N_2935);
nand UO_29 (O_29,N_2936,N_2960);
nand UO_30 (O_30,N_2946,N_2954);
nand UO_31 (O_31,N_2920,N_2928);
xnor UO_32 (O_32,N_2977,N_2900);
nand UO_33 (O_33,N_2916,N_2902);
nor UO_34 (O_34,N_2993,N_2972);
nand UO_35 (O_35,N_2904,N_2975);
and UO_36 (O_36,N_2911,N_2967);
or UO_37 (O_37,N_2990,N_2957);
and UO_38 (O_38,N_2973,N_2929);
or UO_39 (O_39,N_2984,N_2966);
nor UO_40 (O_40,N_2909,N_2974);
nand UO_41 (O_41,N_2991,N_2983);
or UO_42 (O_42,N_2941,N_2940);
and UO_43 (O_43,N_2978,N_2971);
nand UO_44 (O_44,N_2999,N_2934);
or UO_45 (O_45,N_2944,N_2953);
nand UO_46 (O_46,N_2980,N_2926);
nor UO_47 (O_47,N_2982,N_2942);
or UO_48 (O_48,N_2963,N_2950);
xor UO_49 (O_49,N_2959,N_2931);
and UO_50 (O_50,N_2914,N_2933);
nor UO_51 (O_51,N_2901,N_2967);
nand UO_52 (O_52,N_2920,N_2998);
or UO_53 (O_53,N_2921,N_2947);
or UO_54 (O_54,N_2967,N_2964);
or UO_55 (O_55,N_2945,N_2967);
nor UO_56 (O_56,N_2980,N_2986);
and UO_57 (O_57,N_2964,N_2970);
and UO_58 (O_58,N_2952,N_2921);
nor UO_59 (O_59,N_2991,N_2978);
xnor UO_60 (O_60,N_2914,N_2984);
nor UO_61 (O_61,N_2901,N_2999);
nor UO_62 (O_62,N_2905,N_2931);
nor UO_63 (O_63,N_2905,N_2998);
or UO_64 (O_64,N_2907,N_2997);
nand UO_65 (O_65,N_2913,N_2953);
and UO_66 (O_66,N_2927,N_2996);
nor UO_67 (O_67,N_2903,N_2964);
nor UO_68 (O_68,N_2961,N_2902);
and UO_69 (O_69,N_2910,N_2960);
and UO_70 (O_70,N_2905,N_2925);
nand UO_71 (O_71,N_2981,N_2903);
nand UO_72 (O_72,N_2923,N_2975);
and UO_73 (O_73,N_2948,N_2960);
or UO_74 (O_74,N_2976,N_2959);
nand UO_75 (O_75,N_2917,N_2958);
nor UO_76 (O_76,N_2935,N_2979);
and UO_77 (O_77,N_2936,N_2946);
or UO_78 (O_78,N_2940,N_2967);
or UO_79 (O_79,N_2925,N_2970);
and UO_80 (O_80,N_2934,N_2948);
and UO_81 (O_81,N_2989,N_2942);
and UO_82 (O_82,N_2997,N_2978);
nand UO_83 (O_83,N_2916,N_2982);
nand UO_84 (O_84,N_2960,N_2969);
nand UO_85 (O_85,N_2995,N_2999);
nand UO_86 (O_86,N_2993,N_2922);
nor UO_87 (O_87,N_2916,N_2961);
nand UO_88 (O_88,N_2997,N_2911);
and UO_89 (O_89,N_2920,N_2974);
nor UO_90 (O_90,N_2964,N_2984);
xor UO_91 (O_91,N_2906,N_2988);
nand UO_92 (O_92,N_2926,N_2908);
nand UO_93 (O_93,N_2944,N_2950);
nand UO_94 (O_94,N_2900,N_2985);
or UO_95 (O_95,N_2930,N_2907);
nand UO_96 (O_96,N_2992,N_2958);
and UO_97 (O_97,N_2970,N_2995);
or UO_98 (O_98,N_2915,N_2946);
or UO_99 (O_99,N_2977,N_2948);
and UO_100 (O_100,N_2926,N_2915);
or UO_101 (O_101,N_2942,N_2931);
nor UO_102 (O_102,N_2994,N_2906);
nor UO_103 (O_103,N_2929,N_2976);
or UO_104 (O_104,N_2902,N_2970);
or UO_105 (O_105,N_2934,N_2959);
xnor UO_106 (O_106,N_2903,N_2998);
nor UO_107 (O_107,N_2948,N_2987);
or UO_108 (O_108,N_2998,N_2945);
or UO_109 (O_109,N_2997,N_2930);
and UO_110 (O_110,N_2960,N_2968);
nor UO_111 (O_111,N_2995,N_2921);
nand UO_112 (O_112,N_2969,N_2925);
nor UO_113 (O_113,N_2986,N_2911);
and UO_114 (O_114,N_2900,N_2979);
nand UO_115 (O_115,N_2984,N_2926);
nand UO_116 (O_116,N_2913,N_2959);
nand UO_117 (O_117,N_2987,N_2902);
and UO_118 (O_118,N_2919,N_2916);
and UO_119 (O_119,N_2913,N_2973);
nand UO_120 (O_120,N_2941,N_2999);
and UO_121 (O_121,N_2949,N_2950);
nand UO_122 (O_122,N_2901,N_2920);
and UO_123 (O_123,N_2947,N_2951);
nand UO_124 (O_124,N_2948,N_2963);
and UO_125 (O_125,N_2959,N_2980);
nand UO_126 (O_126,N_2983,N_2917);
nand UO_127 (O_127,N_2903,N_2906);
nand UO_128 (O_128,N_2911,N_2971);
nor UO_129 (O_129,N_2985,N_2967);
and UO_130 (O_130,N_2996,N_2924);
or UO_131 (O_131,N_2959,N_2941);
nor UO_132 (O_132,N_2910,N_2966);
nand UO_133 (O_133,N_2946,N_2938);
or UO_134 (O_134,N_2908,N_2959);
nor UO_135 (O_135,N_2903,N_2988);
or UO_136 (O_136,N_2987,N_2937);
and UO_137 (O_137,N_2930,N_2941);
nand UO_138 (O_138,N_2950,N_2945);
nor UO_139 (O_139,N_2944,N_2988);
nand UO_140 (O_140,N_2983,N_2980);
nand UO_141 (O_141,N_2986,N_2943);
or UO_142 (O_142,N_2964,N_2908);
and UO_143 (O_143,N_2995,N_2975);
or UO_144 (O_144,N_2973,N_2900);
and UO_145 (O_145,N_2958,N_2929);
and UO_146 (O_146,N_2932,N_2953);
nand UO_147 (O_147,N_2950,N_2965);
nor UO_148 (O_148,N_2930,N_2933);
xor UO_149 (O_149,N_2924,N_2936);
nand UO_150 (O_150,N_2911,N_2903);
and UO_151 (O_151,N_2946,N_2948);
nand UO_152 (O_152,N_2994,N_2913);
nor UO_153 (O_153,N_2955,N_2919);
or UO_154 (O_154,N_2972,N_2987);
and UO_155 (O_155,N_2926,N_2931);
nor UO_156 (O_156,N_2950,N_2980);
and UO_157 (O_157,N_2941,N_2950);
nor UO_158 (O_158,N_2981,N_2936);
nand UO_159 (O_159,N_2993,N_2983);
and UO_160 (O_160,N_2944,N_2993);
nand UO_161 (O_161,N_2932,N_2923);
and UO_162 (O_162,N_2919,N_2901);
and UO_163 (O_163,N_2952,N_2922);
nor UO_164 (O_164,N_2929,N_2940);
or UO_165 (O_165,N_2909,N_2910);
or UO_166 (O_166,N_2977,N_2932);
nor UO_167 (O_167,N_2960,N_2926);
nand UO_168 (O_168,N_2982,N_2911);
nand UO_169 (O_169,N_2992,N_2916);
or UO_170 (O_170,N_2946,N_2967);
nor UO_171 (O_171,N_2994,N_2907);
nor UO_172 (O_172,N_2918,N_2939);
nor UO_173 (O_173,N_2966,N_2969);
and UO_174 (O_174,N_2903,N_2960);
or UO_175 (O_175,N_2957,N_2950);
nor UO_176 (O_176,N_2984,N_2974);
nand UO_177 (O_177,N_2923,N_2920);
and UO_178 (O_178,N_2921,N_2974);
nand UO_179 (O_179,N_2987,N_2900);
or UO_180 (O_180,N_2967,N_2974);
and UO_181 (O_181,N_2956,N_2970);
nor UO_182 (O_182,N_2956,N_2917);
and UO_183 (O_183,N_2961,N_2913);
and UO_184 (O_184,N_2911,N_2972);
or UO_185 (O_185,N_2906,N_2975);
nor UO_186 (O_186,N_2916,N_2920);
or UO_187 (O_187,N_2908,N_2994);
and UO_188 (O_188,N_2979,N_2937);
nand UO_189 (O_189,N_2996,N_2908);
nor UO_190 (O_190,N_2908,N_2944);
nand UO_191 (O_191,N_2919,N_2969);
and UO_192 (O_192,N_2989,N_2902);
nand UO_193 (O_193,N_2962,N_2904);
nand UO_194 (O_194,N_2913,N_2923);
nor UO_195 (O_195,N_2955,N_2939);
nand UO_196 (O_196,N_2999,N_2985);
xnor UO_197 (O_197,N_2926,N_2909);
nand UO_198 (O_198,N_2921,N_2924);
or UO_199 (O_199,N_2969,N_2996);
and UO_200 (O_200,N_2980,N_2998);
nand UO_201 (O_201,N_2950,N_2975);
and UO_202 (O_202,N_2997,N_2995);
and UO_203 (O_203,N_2998,N_2927);
nor UO_204 (O_204,N_2914,N_2921);
or UO_205 (O_205,N_2971,N_2951);
and UO_206 (O_206,N_2963,N_2949);
xor UO_207 (O_207,N_2984,N_2980);
and UO_208 (O_208,N_2957,N_2916);
nand UO_209 (O_209,N_2970,N_2946);
nand UO_210 (O_210,N_2965,N_2969);
or UO_211 (O_211,N_2994,N_2990);
xnor UO_212 (O_212,N_2933,N_2903);
nand UO_213 (O_213,N_2984,N_2999);
or UO_214 (O_214,N_2926,N_2957);
nand UO_215 (O_215,N_2915,N_2921);
or UO_216 (O_216,N_2969,N_2999);
nand UO_217 (O_217,N_2939,N_2954);
or UO_218 (O_218,N_2959,N_2960);
or UO_219 (O_219,N_2967,N_2959);
nor UO_220 (O_220,N_2930,N_2987);
and UO_221 (O_221,N_2978,N_2922);
nor UO_222 (O_222,N_2907,N_2970);
nand UO_223 (O_223,N_2987,N_2984);
or UO_224 (O_224,N_2972,N_2957);
and UO_225 (O_225,N_2932,N_2997);
nor UO_226 (O_226,N_2946,N_2926);
or UO_227 (O_227,N_2995,N_2981);
nand UO_228 (O_228,N_2975,N_2961);
nand UO_229 (O_229,N_2982,N_2975);
nand UO_230 (O_230,N_2973,N_2917);
nand UO_231 (O_231,N_2982,N_2959);
nor UO_232 (O_232,N_2959,N_2965);
and UO_233 (O_233,N_2970,N_2973);
nor UO_234 (O_234,N_2972,N_2906);
nand UO_235 (O_235,N_2906,N_2948);
or UO_236 (O_236,N_2970,N_2915);
nand UO_237 (O_237,N_2939,N_2984);
and UO_238 (O_238,N_2956,N_2964);
nor UO_239 (O_239,N_2984,N_2916);
or UO_240 (O_240,N_2917,N_2921);
nand UO_241 (O_241,N_2958,N_2934);
and UO_242 (O_242,N_2942,N_2963);
xor UO_243 (O_243,N_2996,N_2916);
or UO_244 (O_244,N_2945,N_2957);
or UO_245 (O_245,N_2904,N_2993);
nand UO_246 (O_246,N_2944,N_2935);
or UO_247 (O_247,N_2966,N_2943);
or UO_248 (O_248,N_2999,N_2964);
and UO_249 (O_249,N_2912,N_2915);
nor UO_250 (O_250,N_2941,N_2978);
nor UO_251 (O_251,N_2980,N_2933);
nor UO_252 (O_252,N_2937,N_2991);
nor UO_253 (O_253,N_2975,N_2902);
nand UO_254 (O_254,N_2949,N_2980);
nor UO_255 (O_255,N_2936,N_2977);
nand UO_256 (O_256,N_2935,N_2954);
nor UO_257 (O_257,N_2944,N_2996);
and UO_258 (O_258,N_2994,N_2903);
nor UO_259 (O_259,N_2931,N_2961);
nand UO_260 (O_260,N_2988,N_2969);
nor UO_261 (O_261,N_2955,N_2927);
and UO_262 (O_262,N_2979,N_2965);
nand UO_263 (O_263,N_2982,N_2990);
and UO_264 (O_264,N_2945,N_2960);
nor UO_265 (O_265,N_2977,N_2947);
or UO_266 (O_266,N_2961,N_2917);
nor UO_267 (O_267,N_2989,N_2929);
and UO_268 (O_268,N_2914,N_2909);
or UO_269 (O_269,N_2955,N_2978);
nand UO_270 (O_270,N_2990,N_2981);
or UO_271 (O_271,N_2937,N_2914);
and UO_272 (O_272,N_2990,N_2971);
or UO_273 (O_273,N_2916,N_2967);
and UO_274 (O_274,N_2952,N_2994);
and UO_275 (O_275,N_2931,N_2952);
nor UO_276 (O_276,N_2900,N_2995);
nor UO_277 (O_277,N_2911,N_2974);
and UO_278 (O_278,N_2960,N_2944);
and UO_279 (O_279,N_2967,N_2932);
nor UO_280 (O_280,N_2996,N_2952);
nor UO_281 (O_281,N_2986,N_2950);
nor UO_282 (O_282,N_2962,N_2976);
nand UO_283 (O_283,N_2989,N_2988);
nand UO_284 (O_284,N_2917,N_2970);
nor UO_285 (O_285,N_2929,N_2938);
nor UO_286 (O_286,N_2902,N_2925);
nor UO_287 (O_287,N_2981,N_2933);
or UO_288 (O_288,N_2928,N_2930);
or UO_289 (O_289,N_2936,N_2940);
or UO_290 (O_290,N_2999,N_2973);
and UO_291 (O_291,N_2961,N_2947);
and UO_292 (O_292,N_2923,N_2922);
nor UO_293 (O_293,N_2981,N_2921);
nand UO_294 (O_294,N_2953,N_2940);
nor UO_295 (O_295,N_2942,N_2970);
nand UO_296 (O_296,N_2915,N_2900);
and UO_297 (O_297,N_2960,N_2931);
nor UO_298 (O_298,N_2956,N_2985);
and UO_299 (O_299,N_2942,N_2905);
and UO_300 (O_300,N_2978,N_2934);
or UO_301 (O_301,N_2901,N_2970);
nor UO_302 (O_302,N_2970,N_2908);
nand UO_303 (O_303,N_2920,N_2994);
or UO_304 (O_304,N_2917,N_2960);
or UO_305 (O_305,N_2954,N_2904);
and UO_306 (O_306,N_2949,N_2928);
nand UO_307 (O_307,N_2998,N_2907);
or UO_308 (O_308,N_2981,N_2909);
nand UO_309 (O_309,N_2982,N_2937);
nand UO_310 (O_310,N_2923,N_2997);
and UO_311 (O_311,N_2954,N_2975);
nand UO_312 (O_312,N_2923,N_2962);
or UO_313 (O_313,N_2979,N_2933);
nand UO_314 (O_314,N_2956,N_2902);
nor UO_315 (O_315,N_2920,N_2946);
nand UO_316 (O_316,N_2939,N_2995);
or UO_317 (O_317,N_2948,N_2932);
nor UO_318 (O_318,N_2927,N_2993);
nor UO_319 (O_319,N_2983,N_2947);
nor UO_320 (O_320,N_2942,N_2913);
and UO_321 (O_321,N_2946,N_2971);
and UO_322 (O_322,N_2921,N_2993);
nor UO_323 (O_323,N_2988,N_2918);
nor UO_324 (O_324,N_2962,N_2902);
or UO_325 (O_325,N_2992,N_2962);
nor UO_326 (O_326,N_2926,N_2993);
or UO_327 (O_327,N_2977,N_2906);
and UO_328 (O_328,N_2942,N_2971);
or UO_329 (O_329,N_2974,N_2959);
nor UO_330 (O_330,N_2941,N_2965);
or UO_331 (O_331,N_2981,N_2997);
and UO_332 (O_332,N_2914,N_2967);
nand UO_333 (O_333,N_2925,N_2908);
nand UO_334 (O_334,N_2972,N_2950);
nor UO_335 (O_335,N_2935,N_2929);
and UO_336 (O_336,N_2904,N_2935);
nand UO_337 (O_337,N_2965,N_2996);
and UO_338 (O_338,N_2998,N_2944);
and UO_339 (O_339,N_2917,N_2962);
and UO_340 (O_340,N_2995,N_2923);
nand UO_341 (O_341,N_2989,N_2982);
or UO_342 (O_342,N_2987,N_2955);
nor UO_343 (O_343,N_2932,N_2905);
and UO_344 (O_344,N_2949,N_2964);
nand UO_345 (O_345,N_2901,N_2985);
or UO_346 (O_346,N_2903,N_2977);
nand UO_347 (O_347,N_2958,N_2984);
nand UO_348 (O_348,N_2986,N_2928);
nor UO_349 (O_349,N_2981,N_2950);
nand UO_350 (O_350,N_2928,N_2937);
or UO_351 (O_351,N_2965,N_2966);
and UO_352 (O_352,N_2993,N_2903);
and UO_353 (O_353,N_2914,N_2901);
and UO_354 (O_354,N_2957,N_2952);
or UO_355 (O_355,N_2910,N_2946);
nor UO_356 (O_356,N_2952,N_2904);
nand UO_357 (O_357,N_2925,N_2956);
and UO_358 (O_358,N_2983,N_2905);
nor UO_359 (O_359,N_2973,N_2934);
nand UO_360 (O_360,N_2947,N_2974);
or UO_361 (O_361,N_2925,N_2998);
nand UO_362 (O_362,N_2951,N_2909);
and UO_363 (O_363,N_2949,N_2916);
and UO_364 (O_364,N_2940,N_2934);
or UO_365 (O_365,N_2981,N_2922);
and UO_366 (O_366,N_2996,N_2905);
and UO_367 (O_367,N_2973,N_2990);
and UO_368 (O_368,N_2998,N_2955);
nor UO_369 (O_369,N_2985,N_2976);
or UO_370 (O_370,N_2999,N_2914);
and UO_371 (O_371,N_2980,N_2942);
nor UO_372 (O_372,N_2968,N_2981);
and UO_373 (O_373,N_2917,N_2903);
or UO_374 (O_374,N_2920,N_2922);
or UO_375 (O_375,N_2937,N_2939);
xnor UO_376 (O_376,N_2935,N_2988);
or UO_377 (O_377,N_2903,N_2943);
and UO_378 (O_378,N_2934,N_2986);
nand UO_379 (O_379,N_2949,N_2989);
nand UO_380 (O_380,N_2968,N_2943);
nand UO_381 (O_381,N_2911,N_2926);
nor UO_382 (O_382,N_2992,N_2909);
nand UO_383 (O_383,N_2925,N_2948);
and UO_384 (O_384,N_2978,N_2949);
nor UO_385 (O_385,N_2923,N_2941);
or UO_386 (O_386,N_2942,N_2924);
nor UO_387 (O_387,N_2962,N_2953);
and UO_388 (O_388,N_2940,N_2962);
and UO_389 (O_389,N_2906,N_2984);
nor UO_390 (O_390,N_2963,N_2919);
nor UO_391 (O_391,N_2908,N_2995);
or UO_392 (O_392,N_2902,N_2992);
nor UO_393 (O_393,N_2981,N_2924);
and UO_394 (O_394,N_2913,N_2924);
nor UO_395 (O_395,N_2939,N_2935);
or UO_396 (O_396,N_2918,N_2949);
or UO_397 (O_397,N_2964,N_2996);
nand UO_398 (O_398,N_2930,N_2977);
nor UO_399 (O_399,N_2999,N_2921);
nor UO_400 (O_400,N_2918,N_2963);
and UO_401 (O_401,N_2983,N_2928);
nand UO_402 (O_402,N_2967,N_2986);
and UO_403 (O_403,N_2957,N_2964);
or UO_404 (O_404,N_2927,N_2925);
and UO_405 (O_405,N_2980,N_2981);
and UO_406 (O_406,N_2957,N_2983);
and UO_407 (O_407,N_2945,N_2988);
or UO_408 (O_408,N_2983,N_2995);
nor UO_409 (O_409,N_2998,N_2910);
nand UO_410 (O_410,N_2979,N_2922);
and UO_411 (O_411,N_2980,N_2916);
and UO_412 (O_412,N_2935,N_2991);
nand UO_413 (O_413,N_2980,N_2900);
or UO_414 (O_414,N_2912,N_2944);
nor UO_415 (O_415,N_2927,N_2933);
and UO_416 (O_416,N_2948,N_2996);
nand UO_417 (O_417,N_2914,N_2987);
and UO_418 (O_418,N_2905,N_2907);
or UO_419 (O_419,N_2985,N_2913);
nand UO_420 (O_420,N_2955,N_2930);
nor UO_421 (O_421,N_2999,N_2966);
or UO_422 (O_422,N_2960,N_2921);
nor UO_423 (O_423,N_2919,N_2960);
or UO_424 (O_424,N_2963,N_2926);
xor UO_425 (O_425,N_2993,N_2999);
nand UO_426 (O_426,N_2979,N_2908);
nor UO_427 (O_427,N_2935,N_2982);
and UO_428 (O_428,N_2904,N_2996);
and UO_429 (O_429,N_2962,N_2947);
or UO_430 (O_430,N_2923,N_2937);
nor UO_431 (O_431,N_2919,N_2999);
or UO_432 (O_432,N_2908,N_2900);
nor UO_433 (O_433,N_2913,N_2982);
and UO_434 (O_434,N_2954,N_2928);
nor UO_435 (O_435,N_2929,N_2916);
and UO_436 (O_436,N_2907,N_2990);
nor UO_437 (O_437,N_2965,N_2929);
nor UO_438 (O_438,N_2984,N_2978);
and UO_439 (O_439,N_2937,N_2972);
and UO_440 (O_440,N_2927,N_2961);
nor UO_441 (O_441,N_2939,N_2916);
nand UO_442 (O_442,N_2910,N_2920);
or UO_443 (O_443,N_2968,N_2940);
and UO_444 (O_444,N_2949,N_2981);
and UO_445 (O_445,N_2900,N_2914);
nor UO_446 (O_446,N_2983,N_2941);
xor UO_447 (O_447,N_2992,N_2934);
or UO_448 (O_448,N_2917,N_2967);
nor UO_449 (O_449,N_2920,N_2919);
nand UO_450 (O_450,N_2903,N_2904);
and UO_451 (O_451,N_2947,N_2914);
nor UO_452 (O_452,N_2946,N_2968);
nor UO_453 (O_453,N_2912,N_2918);
and UO_454 (O_454,N_2921,N_2937);
and UO_455 (O_455,N_2979,N_2918);
xor UO_456 (O_456,N_2911,N_2975);
nor UO_457 (O_457,N_2931,N_2954);
or UO_458 (O_458,N_2998,N_2993);
nand UO_459 (O_459,N_2939,N_2985);
or UO_460 (O_460,N_2909,N_2929);
nor UO_461 (O_461,N_2979,N_2945);
nor UO_462 (O_462,N_2912,N_2968);
or UO_463 (O_463,N_2968,N_2962);
nor UO_464 (O_464,N_2927,N_2910);
nor UO_465 (O_465,N_2973,N_2959);
nand UO_466 (O_466,N_2963,N_2971);
and UO_467 (O_467,N_2912,N_2989);
nor UO_468 (O_468,N_2968,N_2967);
nor UO_469 (O_469,N_2913,N_2926);
nor UO_470 (O_470,N_2923,N_2948);
and UO_471 (O_471,N_2933,N_2972);
nor UO_472 (O_472,N_2960,N_2914);
and UO_473 (O_473,N_2915,N_2995);
or UO_474 (O_474,N_2972,N_2981);
and UO_475 (O_475,N_2994,N_2925);
and UO_476 (O_476,N_2922,N_2998);
nand UO_477 (O_477,N_2985,N_2959);
nor UO_478 (O_478,N_2908,N_2918);
nor UO_479 (O_479,N_2935,N_2909);
or UO_480 (O_480,N_2994,N_2993);
nand UO_481 (O_481,N_2971,N_2970);
nand UO_482 (O_482,N_2988,N_2986);
nand UO_483 (O_483,N_2997,N_2993);
nand UO_484 (O_484,N_2989,N_2996);
and UO_485 (O_485,N_2929,N_2978);
nand UO_486 (O_486,N_2991,N_2913);
or UO_487 (O_487,N_2999,N_2975);
nand UO_488 (O_488,N_2969,N_2956);
or UO_489 (O_489,N_2954,N_2993);
or UO_490 (O_490,N_2902,N_2947);
nand UO_491 (O_491,N_2950,N_2928);
and UO_492 (O_492,N_2959,N_2999);
and UO_493 (O_493,N_2986,N_2969);
nor UO_494 (O_494,N_2960,N_2970);
nor UO_495 (O_495,N_2974,N_2990);
or UO_496 (O_496,N_2948,N_2942);
or UO_497 (O_497,N_2940,N_2921);
or UO_498 (O_498,N_2909,N_2916);
nand UO_499 (O_499,N_2975,N_2900);
endmodule