module basic_500_3000_500_40_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_219,In_463);
nand U1 (N_1,In_354,In_175);
or U2 (N_2,In_404,In_308);
nand U3 (N_3,In_149,In_464);
nand U4 (N_4,In_227,In_208);
and U5 (N_5,In_465,In_148);
nor U6 (N_6,In_255,In_339);
or U7 (N_7,In_21,In_203);
or U8 (N_8,In_406,In_191);
nor U9 (N_9,In_84,In_104);
nand U10 (N_10,In_487,In_40);
nand U11 (N_11,In_498,In_475);
nand U12 (N_12,In_454,In_410);
nand U13 (N_13,In_393,In_216);
and U14 (N_14,In_81,In_172);
nand U15 (N_15,In_446,In_474);
nand U16 (N_16,In_164,In_229);
or U17 (N_17,In_397,In_422);
and U18 (N_18,In_118,In_232);
nor U19 (N_19,In_234,In_39);
or U20 (N_20,In_356,In_87);
and U21 (N_21,In_161,In_253);
or U22 (N_22,In_94,In_467);
or U23 (N_23,In_184,In_176);
nand U24 (N_24,In_379,In_257);
nand U25 (N_25,In_270,In_8);
and U26 (N_26,In_294,In_70);
nand U27 (N_27,In_77,In_156);
nand U28 (N_28,In_144,In_380);
nor U29 (N_29,In_471,In_490);
or U30 (N_30,In_10,In_412);
or U31 (N_31,In_86,In_388);
or U32 (N_32,In_246,In_181);
nand U33 (N_33,In_190,In_486);
nand U34 (N_34,In_480,In_185);
nand U35 (N_35,In_137,In_83);
and U36 (N_36,In_368,In_66);
and U37 (N_37,In_193,In_38);
and U38 (N_38,In_192,In_302);
and U39 (N_39,In_428,In_279);
nor U40 (N_40,In_129,In_252);
nand U41 (N_41,In_331,In_24);
or U42 (N_42,In_153,In_79);
or U43 (N_43,In_430,In_115);
nor U44 (N_44,In_455,In_108);
nand U45 (N_45,In_305,In_365);
nor U46 (N_46,In_78,In_14);
and U47 (N_47,In_346,In_29);
and U48 (N_48,In_326,In_65);
or U49 (N_49,In_320,In_28);
and U50 (N_50,In_462,In_220);
and U51 (N_51,In_132,In_371);
nand U52 (N_52,In_385,In_286);
or U53 (N_53,In_19,In_399);
or U54 (N_54,In_291,In_324);
nand U55 (N_55,In_206,In_240);
nor U56 (N_56,In_3,In_413);
xor U57 (N_57,In_167,In_401);
nand U58 (N_58,In_12,In_95);
and U59 (N_59,In_9,In_180);
and U60 (N_60,In_492,In_235);
nor U61 (N_61,In_424,In_47);
nand U62 (N_62,In_169,In_30);
or U63 (N_63,In_389,In_280);
and U64 (N_64,In_398,In_458);
nand U65 (N_65,In_131,In_1);
nand U66 (N_66,In_374,In_445);
nor U67 (N_67,In_186,In_448);
nand U68 (N_68,In_441,In_233);
nor U69 (N_69,In_112,In_447);
and U70 (N_70,In_459,In_143);
and U71 (N_71,In_466,In_214);
nand U72 (N_72,In_369,In_157);
and U73 (N_73,In_418,In_5);
or U74 (N_74,In_323,In_198);
and U75 (N_75,In_306,In_439);
nand U76 (N_76,In_272,In_489);
nand U77 (N_77,In_293,In_62);
xnor U78 (N_78,In_20,N_16);
nor U79 (N_79,In_163,In_444);
or U80 (N_80,In_244,N_61);
and U81 (N_81,In_48,In_373);
or U82 (N_82,In_242,In_134);
or U83 (N_83,In_284,N_50);
nand U84 (N_84,N_48,N_19);
or U85 (N_85,In_386,In_338);
or U86 (N_86,In_15,In_375);
nor U87 (N_87,In_178,In_25);
or U88 (N_88,In_37,In_217);
nand U89 (N_89,In_179,In_419);
or U90 (N_90,In_289,N_15);
nand U91 (N_91,N_60,N_7);
and U92 (N_92,In_150,In_63);
nor U93 (N_93,In_400,N_28);
and U94 (N_94,In_92,In_493);
and U95 (N_95,N_73,In_296);
or U96 (N_96,In_189,In_42);
or U97 (N_97,In_473,In_348);
and U98 (N_98,N_51,In_360);
or U99 (N_99,In_350,In_353);
and U100 (N_100,In_23,N_59);
and U101 (N_101,In_391,In_195);
and U102 (N_102,In_225,N_38);
or U103 (N_103,In_482,In_295);
or U104 (N_104,In_89,In_243);
nor U105 (N_105,In_145,In_45);
nand U106 (N_106,In_432,In_314);
nand U107 (N_107,In_138,In_333);
nand U108 (N_108,In_165,In_59);
nand U109 (N_109,In_33,In_322);
and U110 (N_110,In_98,In_120);
nor U111 (N_111,In_174,In_276);
or U112 (N_112,In_200,In_440);
nand U113 (N_113,In_58,In_469);
and U114 (N_114,N_53,In_34);
nand U115 (N_115,N_6,In_249);
and U116 (N_116,In_114,In_13);
and U117 (N_117,In_96,In_158);
or U118 (N_118,N_65,In_248);
or U119 (N_119,In_22,In_151);
or U120 (N_120,In_122,In_409);
nand U121 (N_121,In_290,In_27);
and U122 (N_122,In_362,In_457);
and U123 (N_123,In_263,In_57);
or U124 (N_124,In_188,In_32);
nor U125 (N_125,In_76,In_160);
nand U126 (N_126,In_139,In_256);
nor U127 (N_127,In_100,In_130);
or U128 (N_128,In_69,In_135);
nor U129 (N_129,In_285,In_2);
and U130 (N_130,N_72,In_266);
or U131 (N_131,In_159,N_41);
nand U132 (N_132,In_258,In_381);
and U133 (N_133,N_11,In_402);
nor U134 (N_134,In_363,In_251);
and U135 (N_135,In_202,In_0);
or U136 (N_136,In_116,In_152);
nand U137 (N_137,In_105,In_337);
xnor U138 (N_138,In_301,In_72);
nor U139 (N_139,In_357,In_335);
nor U140 (N_140,In_264,In_405);
nor U141 (N_141,In_147,In_275);
and U142 (N_142,In_491,In_124);
nor U143 (N_143,In_154,In_103);
and U144 (N_144,In_330,In_146);
nand U145 (N_145,In_73,In_75);
nand U146 (N_146,In_64,In_456);
nand U147 (N_147,In_341,In_499);
nor U148 (N_148,N_55,N_27);
or U149 (N_149,In_481,N_35);
nand U150 (N_150,In_355,In_327);
nor U151 (N_151,In_230,N_32);
nor U152 (N_152,In_378,In_476);
and U153 (N_153,N_75,N_0);
nor U154 (N_154,In_318,In_166);
nor U155 (N_155,In_278,In_417);
and U156 (N_156,N_83,In_194);
and U157 (N_157,In_102,N_99);
nor U158 (N_158,N_132,In_171);
or U159 (N_159,In_56,In_182);
nand U160 (N_160,In_82,In_488);
or U161 (N_161,In_361,In_347);
nand U162 (N_162,In_241,In_17);
nor U163 (N_163,N_18,In_218);
or U164 (N_164,In_90,N_80);
nand U165 (N_165,In_427,In_387);
nor U166 (N_166,In_207,N_10);
and U167 (N_167,N_1,In_237);
or U168 (N_168,In_383,In_372);
and U169 (N_169,N_91,In_16);
nand U170 (N_170,N_89,N_40);
nor U171 (N_171,N_70,In_317);
nand U172 (N_172,In_53,In_49);
nand U173 (N_173,In_74,In_483);
and U174 (N_174,N_103,N_37);
nand U175 (N_175,N_114,N_9);
and U176 (N_176,In_414,In_162);
or U177 (N_177,In_31,N_140);
nor U178 (N_178,N_87,N_113);
nor U179 (N_179,N_62,In_50);
or U180 (N_180,In_36,N_131);
or U181 (N_181,In_6,N_49);
or U182 (N_182,In_97,In_312);
or U183 (N_183,In_221,In_61);
or U184 (N_184,In_425,In_332);
nand U185 (N_185,In_484,In_325);
nor U186 (N_186,In_421,In_247);
and U187 (N_187,In_367,N_13);
and U188 (N_188,In_433,In_41);
or U189 (N_189,In_71,In_415);
and U190 (N_190,In_460,In_396);
nand U191 (N_191,In_187,In_311);
nand U192 (N_192,In_315,In_298);
nor U193 (N_193,N_86,N_136);
or U194 (N_194,In_91,In_210);
nand U195 (N_195,In_170,N_66);
or U196 (N_196,In_222,N_110);
or U197 (N_197,N_138,N_39);
nor U198 (N_198,In_283,In_168);
or U199 (N_199,In_259,In_68);
and U200 (N_200,N_88,N_94);
nand U201 (N_201,N_77,N_82);
or U202 (N_202,In_128,In_408);
or U203 (N_203,In_111,In_452);
nor U204 (N_204,In_67,In_420);
nor U205 (N_205,In_7,N_3);
nand U206 (N_206,In_261,In_44);
or U207 (N_207,N_109,In_351);
and U208 (N_208,In_213,N_64);
nand U209 (N_209,In_468,In_359);
nand U210 (N_210,In_403,In_262);
nand U211 (N_211,In_236,N_47);
and U212 (N_212,In_140,N_31);
nand U213 (N_213,N_102,In_110);
nor U214 (N_214,In_277,In_224);
and U215 (N_215,N_76,N_98);
xor U216 (N_216,In_342,In_99);
and U217 (N_217,In_438,N_68);
and U218 (N_218,In_431,N_56);
nor U219 (N_219,In_245,N_63);
nor U220 (N_220,N_2,N_58);
or U221 (N_221,N_122,In_345);
nor U222 (N_222,N_118,In_382);
nand U223 (N_223,In_250,In_470);
nand U224 (N_224,In_377,N_90);
nor U225 (N_225,N_85,N_127);
nand U226 (N_226,N_4,In_334);
nand U227 (N_227,N_23,In_392);
or U228 (N_228,N_218,In_376);
and U229 (N_229,In_260,N_96);
nor U230 (N_230,In_358,N_160);
or U231 (N_231,N_172,N_104);
or U232 (N_232,In_267,N_142);
or U233 (N_233,In_485,In_46);
or U234 (N_234,N_79,In_155);
and U235 (N_235,N_100,In_328);
nor U236 (N_236,N_215,In_478);
or U237 (N_237,N_188,N_166);
or U238 (N_238,N_180,N_25);
nor U239 (N_239,In_226,In_197);
and U240 (N_240,N_134,N_165);
nand U241 (N_241,N_153,N_185);
or U242 (N_242,N_183,N_181);
or U243 (N_243,N_42,In_435);
or U244 (N_244,In_273,N_24);
and U245 (N_245,In_416,In_126);
nor U246 (N_246,N_202,In_395);
nor U247 (N_247,In_142,In_479);
nand U248 (N_248,N_187,N_179);
or U249 (N_249,In_352,N_173);
or U250 (N_250,N_108,In_196);
or U251 (N_251,N_149,In_390);
nand U252 (N_252,N_157,In_177);
nand U253 (N_253,N_164,N_176);
nor U254 (N_254,In_349,In_52);
nor U255 (N_255,In_394,N_57);
and U256 (N_256,In_450,N_152);
and U257 (N_257,N_111,In_321);
nor U258 (N_258,In_60,N_105);
and U259 (N_259,In_442,N_84);
nand U260 (N_260,In_223,N_162);
or U261 (N_261,N_175,In_310);
and U262 (N_262,N_154,In_437);
nand U263 (N_263,In_271,N_81);
and U264 (N_264,N_26,N_159);
nand U265 (N_265,In_496,N_174);
nand U266 (N_266,In_303,N_135);
or U267 (N_267,In_127,In_201);
nand U268 (N_268,In_461,N_222);
nor U269 (N_269,N_147,N_123);
or U270 (N_270,N_192,In_117);
xnor U271 (N_271,In_495,In_35);
and U272 (N_272,N_190,In_11);
nand U273 (N_273,In_313,N_212);
or U274 (N_274,N_119,In_136);
or U275 (N_275,N_139,In_423);
nor U276 (N_276,N_211,N_12);
nand U277 (N_277,In_297,In_370);
nor U278 (N_278,In_101,In_113);
or U279 (N_279,In_212,N_30);
nor U280 (N_280,In_497,N_167);
and U281 (N_281,In_434,N_204);
nor U282 (N_282,N_146,N_143);
nor U283 (N_283,In_411,In_4);
nand U284 (N_284,N_43,In_384);
nand U285 (N_285,In_426,N_46);
xor U286 (N_286,In_449,In_443);
nand U287 (N_287,N_128,In_18);
nor U288 (N_288,In_51,N_155);
nor U289 (N_289,In_477,N_182);
nor U290 (N_290,N_213,N_210);
nand U291 (N_291,N_106,N_201);
nor U292 (N_292,In_133,N_200);
nand U293 (N_293,In_209,In_123);
nand U294 (N_294,In_239,In_319);
or U295 (N_295,N_33,N_178);
nor U296 (N_296,N_145,N_44);
nor U297 (N_297,N_195,In_429);
and U298 (N_298,N_171,N_29);
and U299 (N_299,N_129,N_126);
or U300 (N_300,In_211,In_281);
and U301 (N_301,N_240,N_112);
nand U302 (N_302,N_45,In_307);
nor U303 (N_303,N_245,N_193);
nor U304 (N_304,In_121,N_276);
nor U305 (N_305,N_232,N_69);
and U306 (N_306,N_293,N_246);
and U307 (N_307,N_272,N_241);
nand U308 (N_308,N_283,In_304);
nand U309 (N_309,N_219,N_78);
and U310 (N_310,N_107,N_34);
nand U311 (N_311,In_336,N_170);
nor U312 (N_312,N_228,N_17);
nand U313 (N_313,N_298,N_299);
nor U314 (N_314,N_217,In_107);
and U315 (N_315,N_256,In_343);
and U316 (N_316,N_254,In_282);
and U317 (N_317,N_287,N_238);
nor U318 (N_318,In_316,In_287);
nand U319 (N_319,N_156,N_230);
nand U320 (N_320,N_8,N_92);
nor U321 (N_321,N_169,In_309);
or U322 (N_322,N_295,N_225);
or U323 (N_323,N_93,N_294);
nor U324 (N_324,In_407,In_265);
nor U325 (N_325,N_284,N_253);
and U326 (N_326,In_254,N_168);
or U327 (N_327,N_289,In_106);
and U328 (N_328,N_291,N_67);
and U329 (N_329,N_280,N_71);
nor U330 (N_330,In_199,N_271);
or U331 (N_331,N_275,N_262);
nor U332 (N_332,N_235,N_197);
and U333 (N_333,In_85,N_141);
nand U334 (N_334,In_43,N_116);
or U335 (N_335,N_285,N_36);
and U336 (N_336,In_183,In_494);
nand U337 (N_337,N_121,In_299);
nor U338 (N_338,N_52,N_163);
nor U339 (N_339,In_436,N_124);
nor U340 (N_340,In_88,N_22);
nor U341 (N_341,In_366,N_279);
nand U342 (N_342,In_238,N_101);
and U343 (N_343,N_273,In_288);
or U344 (N_344,N_198,N_277);
or U345 (N_345,N_243,N_74);
nand U346 (N_346,N_158,N_194);
and U347 (N_347,In_269,N_269);
nor U348 (N_348,N_144,N_297);
or U349 (N_349,N_278,N_130);
or U350 (N_350,N_137,In_340);
nor U351 (N_351,N_281,In_215);
and U352 (N_352,N_296,N_191);
nor U353 (N_353,N_227,N_233);
nor U354 (N_354,N_261,N_117);
and U355 (N_355,In_109,N_220);
nand U356 (N_356,N_224,N_292);
nor U357 (N_357,N_186,N_189);
and U358 (N_358,N_226,In_119);
or U359 (N_359,N_290,N_115);
nor U360 (N_360,N_97,In_125);
nand U361 (N_361,N_268,N_95);
nor U362 (N_362,N_184,N_266);
nand U363 (N_363,N_255,N_21);
or U364 (N_364,In_228,N_263);
nor U365 (N_365,N_209,In_451);
or U366 (N_366,In_141,In_292);
or U367 (N_367,N_161,N_203);
nor U368 (N_368,N_231,N_274);
and U369 (N_369,N_148,N_257);
or U370 (N_370,In_364,N_54);
and U371 (N_371,In_274,N_207);
nor U372 (N_372,N_248,N_288);
nand U373 (N_373,In_231,N_221);
or U374 (N_374,In_329,In_54);
nor U375 (N_375,N_358,N_322);
nor U376 (N_376,N_270,N_20);
and U377 (N_377,N_310,N_150);
or U378 (N_378,N_330,N_319);
nand U379 (N_379,N_199,N_332);
or U380 (N_380,N_214,N_326);
nor U381 (N_381,N_252,N_300);
and U382 (N_382,N_353,N_320);
and U383 (N_383,N_229,N_350);
nor U384 (N_384,N_368,In_268);
and U385 (N_385,N_205,N_267);
nor U386 (N_386,N_301,N_206);
nor U387 (N_387,N_335,N_325);
and U388 (N_388,N_333,N_304);
nor U389 (N_389,N_302,N_329);
nor U390 (N_390,N_234,N_344);
or U391 (N_391,N_151,N_264);
nor U392 (N_392,N_259,In_93);
nand U393 (N_393,N_258,In_80);
nand U394 (N_394,N_236,N_286);
nor U395 (N_395,N_120,N_342);
nor U396 (N_396,N_340,N_321);
nand U397 (N_397,N_360,N_314);
nand U398 (N_398,N_363,N_208);
and U399 (N_399,N_336,N_351);
or U400 (N_400,N_338,In_344);
and U401 (N_401,N_323,N_216);
nor U402 (N_402,N_316,N_369);
or U403 (N_403,N_352,N_327);
or U404 (N_404,N_328,N_318);
or U405 (N_405,N_346,N_354);
nand U406 (N_406,In_173,N_349);
and U407 (N_407,N_362,N_356);
and U408 (N_408,N_306,N_247);
nand U409 (N_409,In_55,In_26);
or U410 (N_410,N_337,N_324);
nor U411 (N_411,N_355,N_312);
nand U412 (N_412,N_315,N_311);
and U413 (N_413,N_308,N_371);
nand U414 (N_414,N_366,N_250);
or U415 (N_415,N_237,N_305);
and U416 (N_416,N_359,In_205);
or U417 (N_417,N_307,N_244);
and U418 (N_418,N_341,N_309);
or U419 (N_419,N_334,N_364);
and U420 (N_420,In_300,N_348);
or U421 (N_421,N_125,N_242);
or U422 (N_422,N_361,N_249);
or U423 (N_423,N_14,N_177);
and U424 (N_424,N_239,In_453);
nor U425 (N_425,N_196,N_372);
and U426 (N_426,N_347,N_339);
or U427 (N_427,N_282,N_317);
and U428 (N_428,N_5,N_223);
nor U429 (N_429,N_370,N_265);
or U430 (N_430,N_365,N_260);
or U431 (N_431,N_133,N_303);
and U432 (N_432,N_251,N_343);
nor U433 (N_433,In_472,N_331);
nor U434 (N_434,In_204,N_367);
and U435 (N_435,N_313,N_374);
nor U436 (N_436,N_345,N_357);
or U437 (N_437,N_373,In_300);
and U438 (N_438,N_366,N_264);
nand U439 (N_439,N_352,In_80);
nor U440 (N_440,N_264,N_373);
nand U441 (N_441,N_199,N_367);
and U442 (N_442,N_373,N_249);
nand U443 (N_443,N_223,N_306);
and U444 (N_444,N_326,N_252);
nor U445 (N_445,N_352,N_234);
and U446 (N_446,N_244,N_303);
or U447 (N_447,N_336,N_309);
nor U448 (N_448,N_331,N_372);
nand U449 (N_449,N_133,N_196);
or U450 (N_450,N_446,N_444);
nor U451 (N_451,N_397,N_411);
nor U452 (N_452,N_420,N_422);
and U453 (N_453,N_384,N_394);
or U454 (N_454,N_445,N_423);
or U455 (N_455,N_408,N_386);
nand U456 (N_456,N_441,N_432);
nor U457 (N_457,N_410,N_389);
nor U458 (N_458,N_424,N_396);
or U459 (N_459,N_431,N_398);
nand U460 (N_460,N_388,N_442);
and U461 (N_461,N_399,N_376);
and U462 (N_462,N_390,N_434);
nor U463 (N_463,N_402,N_425);
and U464 (N_464,N_375,N_439);
or U465 (N_465,N_403,N_438);
and U466 (N_466,N_392,N_379);
nor U467 (N_467,N_443,N_409);
nor U468 (N_468,N_412,N_415);
nor U469 (N_469,N_393,N_401);
nand U470 (N_470,N_430,N_405);
nand U471 (N_471,N_378,N_381);
nand U472 (N_472,N_427,N_413);
nor U473 (N_473,N_391,N_400);
and U474 (N_474,N_416,N_437);
nand U475 (N_475,N_433,N_395);
or U476 (N_476,N_421,N_435);
or U477 (N_477,N_448,N_426);
and U478 (N_478,N_383,N_406);
and U479 (N_479,N_407,N_385);
and U480 (N_480,N_417,N_414);
and U481 (N_481,N_382,N_429);
nand U482 (N_482,N_380,N_377);
or U483 (N_483,N_449,N_419);
nor U484 (N_484,N_428,N_440);
nor U485 (N_485,N_387,N_436);
nand U486 (N_486,N_447,N_404);
and U487 (N_487,N_418,N_426);
nor U488 (N_488,N_402,N_432);
and U489 (N_489,N_426,N_399);
and U490 (N_490,N_401,N_436);
and U491 (N_491,N_393,N_380);
nand U492 (N_492,N_400,N_398);
nand U493 (N_493,N_415,N_396);
nand U494 (N_494,N_427,N_441);
nand U495 (N_495,N_431,N_395);
nand U496 (N_496,N_421,N_397);
and U497 (N_497,N_416,N_428);
and U498 (N_498,N_415,N_400);
or U499 (N_499,N_375,N_420);
and U500 (N_500,N_439,N_403);
nand U501 (N_501,N_386,N_390);
or U502 (N_502,N_449,N_389);
and U503 (N_503,N_382,N_438);
nand U504 (N_504,N_397,N_446);
and U505 (N_505,N_419,N_423);
or U506 (N_506,N_421,N_404);
nand U507 (N_507,N_442,N_400);
or U508 (N_508,N_445,N_394);
nand U509 (N_509,N_379,N_449);
nor U510 (N_510,N_441,N_442);
or U511 (N_511,N_415,N_407);
nor U512 (N_512,N_409,N_416);
nand U513 (N_513,N_405,N_423);
and U514 (N_514,N_375,N_418);
or U515 (N_515,N_401,N_408);
nand U516 (N_516,N_406,N_376);
nor U517 (N_517,N_440,N_402);
nand U518 (N_518,N_417,N_387);
nor U519 (N_519,N_419,N_385);
or U520 (N_520,N_418,N_383);
nor U521 (N_521,N_431,N_418);
nand U522 (N_522,N_378,N_404);
and U523 (N_523,N_448,N_435);
and U524 (N_524,N_399,N_388);
nor U525 (N_525,N_466,N_512);
and U526 (N_526,N_460,N_515);
nand U527 (N_527,N_471,N_517);
or U528 (N_528,N_457,N_478);
and U529 (N_529,N_509,N_482);
and U530 (N_530,N_487,N_463);
nand U531 (N_531,N_514,N_510);
nand U532 (N_532,N_494,N_522);
nand U533 (N_533,N_453,N_505);
or U534 (N_534,N_518,N_481);
or U535 (N_535,N_454,N_516);
or U536 (N_536,N_480,N_484);
nand U537 (N_537,N_459,N_524);
and U538 (N_538,N_488,N_479);
nand U539 (N_539,N_461,N_492);
and U540 (N_540,N_468,N_469);
xnor U541 (N_541,N_477,N_503);
nor U542 (N_542,N_483,N_473);
and U543 (N_543,N_493,N_456);
or U544 (N_544,N_499,N_523);
nor U545 (N_545,N_451,N_501);
nand U546 (N_546,N_465,N_520);
and U547 (N_547,N_486,N_472);
nand U548 (N_548,N_467,N_455);
nand U549 (N_549,N_474,N_462);
nor U550 (N_550,N_495,N_508);
or U551 (N_551,N_458,N_491);
nor U552 (N_552,N_507,N_485);
nand U553 (N_553,N_506,N_504);
or U554 (N_554,N_476,N_452);
or U555 (N_555,N_470,N_496);
and U556 (N_556,N_450,N_502);
nor U557 (N_557,N_497,N_521);
or U558 (N_558,N_511,N_500);
nor U559 (N_559,N_513,N_464);
and U560 (N_560,N_519,N_489);
and U561 (N_561,N_490,N_498);
nand U562 (N_562,N_475,N_474);
or U563 (N_563,N_481,N_482);
nand U564 (N_564,N_453,N_490);
nor U565 (N_565,N_487,N_456);
nor U566 (N_566,N_473,N_501);
nor U567 (N_567,N_494,N_523);
nor U568 (N_568,N_479,N_503);
or U569 (N_569,N_452,N_451);
or U570 (N_570,N_500,N_495);
nand U571 (N_571,N_474,N_524);
nor U572 (N_572,N_505,N_465);
or U573 (N_573,N_509,N_466);
nor U574 (N_574,N_474,N_471);
nor U575 (N_575,N_478,N_492);
or U576 (N_576,N_456,N_491);
nor U577 (N_577,N_501,N_517);
nor U578 (N_578,N_518,N_464);
nor U579 (N_579,N_467,N_499);
nand U580 (N_580,N_459,N_480);
nor U581 (N_581,N_480,N_478);
and U582 (N_582,N_450,N_451);
and U583 (N_583,N_478,N_499);
and U584 (N_584,N_504,N_468);
nand U585 (N_585,N_497,N_464);
or U586 (N_586,N_450,N_477);
or U587 (N_587,N_506,N_498);
nand U588 (N_588,N_475,N_480);
nor U589 (N_589,N_454,N_501);
nor U590 (N_590,N_468,N_524);
nand U591 (N_591,N_517,N_489);
nand U592 (N_592,N_484,N_523);
and U593 (N_593,N_516,N_497);
nor U594 (N_594,N_478,N_513);
and U595 (N_595,N_479,N_513);
nand U596 (N_596,N_464,N_458);
xnor U597 (N_597,N_487,N_506);
nor U598 (N_598,N_452,N_454);
nand U599 (N_599,N_518,N_477);
nand U600 (N_600,N_534,N_599);
and U601 (N_601,N_527,N_554);
nor U602 (N_602,N_595,N_571);
nor U603 (N_603,N_579,N_564);
and U604 (N_604,N_591,N_573);
or U605 (N_605,N_560,N_544);
nand U606 (N_606,N_533,N_598);
nand U607 (N_607,N_578,N_535);
and U608 (N_608,N_528,N_584);
nor U609 (N_609,N_588,N_559);
or U610 (N_610,N_563,N_572);
nand U611 (N_611,N_550,N_581);
or U612 (N_612,N_575,N_548);
nand U613 (N_613,N_594,N_580);
or U614 (N_614,N_526,N_585);
and U615 (N_615,N_547,N_592);
and U616 (N_616,N_593,N_541);
nand U617 (N_617,N_558,N_566);
and U618 (N_618,N_537,N_538);
nor U619 (N_619,N_567,N_590);
nor U620 (N_620,N_568,N_551);
nor U621 (N_621,N_582,N_586);
nor U622 (N_622,N_553,N_540);
and U623 (N_623,N_577,N_539);
or U624 (N_624,N_596,N_536);
nor U625 (N_625,N_530,N_574);
nand U626 (N_626,N_561,N_525);
and U627 (N_627,N_531,N_565);
nand U628 (N_628,N_552,N_562);
or U629 (N_629,N_542,N_597);
or U630 (N_630,N_583,N_546);
nor U631 (N_631,N_529,N_557);
nor U632 (N_632,N_569,N_545);
or U633 (N_633,N_549,N_576);
and U634 (N_634,N_532,N_556);
nand U635 (N_635,N_555,N_543);
and U636 (N_636,N_587,N_589);
and U637 (N_637,N_570,N_587);
and U638 (N_638,N_554,N_565);
and U639 (N_639,N_566,N_553);
or U640 (N_640,N_560,N_537);
or U641 (N_641,N_559,N_568);
nand U642 (N_642,N_569,N_543);
nor U643 (N_643,N_530,N_593);
nand U644 (N_644,N_568,N_579);
and U645 (N_645,N_540,N_542);
or U646 (N_646,N_525,N_589);
or U647 (N_647,N_594,N_571);
or U648 (N_648,N_576,N_527);
and U649 (N_649,N_533,N_530);
and U650 (N_650,N_571,N_597);
nor U651 (N_651,N_583,N_579);
and U652 (N_652,N_525,N_590);
and U653 (N_653,N_579,N_588);
or U654 (N_654,N_563,N_574);
nand U655 (N_655,N_544,N_561);
nand U656 (N_656,N_596,N_581);
or U657 (N_657,N_586,N_580);
or U658 (N_658,N_562,N_553);
nand U659 (N_659,N_583,N_584);
and U660 (N_660,N_583,N_532);
or U661 (N_661,N_566,N_556);
or U662 (N_662,N_599,N_550);
nand U663 (N_663,N_575,N_530);
nor U664 (N_664,N_533,N_537);
or U665 (N_665,N_530,N_526);
nor U666 (N_666,N_590,N_587);
nand U667 (N_667,N_534,N_541);
or U668 (N_668,N_545,N_580);
nand U669 (N_669,N_548,N_554);
and U670 (N_670,N_533,N_574);
or U671 (N_671,N_526,N_591);
or U672 (N_672,N_562,N_566);
and U673 (N_673,N_538,N_572);
nor U674 (N_674,N_578,N_557);
and U675 (N_675,N_632,N_619);
or U676 (N_676,N_670,N_665);
or U677 (N_677,N_629,N_654);
nor U678 (N_678,N_655,N_646);
or U679 (N_679,N_674,N_627);
and U680 (N_680,N_666,N_633);
and U681 (N_681,N_603,N_650);
nand U682 (N_682,N_615,N_620);
and U683 (N_683,N_611,N_631);
or U684 (N_684,N_637,N_667);
nor U685 (N_685,N_652,N_641);
or U686 (N_686,N_653,N_656);
nor U687 (N_687,N_638,N_659);
and U688 (N_688,N_609,N_601);
and U689 (N_689,N_606,N_673);
and U690 (N_690,N_643,N_616);
or U691 (N_691,N_602,N_648);
or U692 (N_692,N_625,N_604);
or U693 (N_693,N_617,N_628);
nor U694 (N_694,N_608,N_644);
nor U695 (N_695,N_651,N_649);
or U696 (N_696,N_664,N_607);
and U697 (N_697,N_613,N_647);
nor U698 (N_698,N_614,N_658);
or U699 (N_699,N_621,N_639);
nand U700 (N_700,N_640,N_671);
nor U701 (N_701,N_645,N_623);
nor U702 (N_702,N_624,N_622);
nand U703 (N_703,N_672,N_661);
nor U704 (N_704,N_636,N_626);
or U705 (N_705,N_663,N_660);
nand U706 (N_706,N_642,N_610);
or U707 (N_707,N_600,N_630);
or U708 (N_708,N_634,N_657);
or U709 (N_709,N_669,N_618);
nand U710 (N_710,N_662,N_605);
or U711 (N_711,N_612,N_668);
nand U712 (N_712,N_635,N_651);
nand U713 (N_713,N_664,N_629);
and U714 (N_714,N_615,N_626);
and U715 (N_715,N_647,N_644);
or U716 (N_716,N_632,N_606);
and U717 (N_717,N_635,N_618);
and U718 (N_718,N_671,N_644);
nand U719 (N_719,N_652,N_672);
nand U720 (N_720,N_624,N_667);
and U721 (N_721,N_638,N_662);
or U722 (N_722,N_669,N_631);
and U723 (N_723,N_651,N_642);
nand U724 (N_724,N_631,N_625);
nand U725 (N_725,N_627,N_609);
nor U726 (N_726,N_619,N_611);
nand U727 (N_727,N_645,N_616);
nand U728 (N_728,N_605,N_628);
or U729 (N_729,N_601,N_623);
or U730 (N_730,N_648,N_616);
nor U731 (N_731,N_631,N_628);
and U732 (N_732,N_617,N_646);
nor U733 (N_733,N_655,N_612);
or U734 (N_734,N_654,N_631);
or U735 (N_735,N_622,N_659);
xnor U736 (N_736,N_632,N_649);
and U737 (N_737,N_645,N_611);
or U738 (N_738,N_642,N_659);
nand U739 (N_739,N_648,N_650);
nor U740 (N_740,N_605,N_668);
or U741 (N_741,N_665,N_651);
and U742 (N_742,N_625,N_663);
or U743 (N_743,N_642,N_636);
and U744 (N_744,N_609,N_665);
nor U745 (N_745,N_626,N_653);
xnor U746 (N_746,N_667,N_615);
nand U747 (N_747,N_644,N_626);
nand U748 (N_748,N_606,N_651);
and U749 (N_749,N_657,N_652);
and U750 (N_750,N_731,N_687);
or U751 (N_751,N_702,N_683);
or U752 (N_752,N_700,N_706);
nand U753 (N_753,N_730,N_686);
nand U754 (N_754,N_717,N_684);
or U755 (N_755,N_718,N_693);
nand U756 (N_756,N_749,N_746);
nor U757 (N_757,N_695,N_698);
or U758 (N_758,N_716,N_747);
or U759 (N_759,N_710,N_734);
or U760 (N_760,N_676,N_694);
nand U761 (N_761,N_707,N_745);
or U762 (N_762,N_678,N_725);
or U763 (N_763,N_689,N_735);
and U764 (N_764,N_711,N_696);
or U765 (N_765,N_715,N_722);
xnor U766 (N_766,N_708,N_692);
and U767 (N_767,N_737,N_729);
and U768 (N_768,N_677,N_739);
or U769 (N_769,N_748,N_713);
nor U770 (N_770,N_701,N_680);
or U771 (N_771,N_744,N_728);
nor U772 (N_772,N_726,N_727);
nand U773 (N_773,N_675,N_719);
and U774 (N_774,N_682,N_703);
or U775 (N_775,N_681,N_738);
nand U776 (N_776,N_723,N_688);
nand U777 (N_777,N_709,N_690);
nand U778 (N_778,N_714,N_736);
or U779 (N_779,N_721,N_704);
nor U780 (N_780,N_742,N_733);
nor U781 (N_781,N_732,N_720);
and U782 (N_782,N_685,N_705);
and U783 (N_783,N_712,N_740);
nor U784 (N_784,N_691,N_697);
nand U785 (N_785,N_679,N_741);
nand U786 (N_786,N_699,N_724);
nor U787 (N_787,N_743,N_690);
nor U788 (N_788,N_711,N_702);
nor U789 (N_789,N_738,N_722);
and U790 (N_790,N_709,N_701);
nand U791 (N_791,N_676,N_744);
and U792 (N_792,N_736,N_720);
nand U793 (N_793,N_681,N_737);
nand U794 (N_794,N_682,N_685);
nand U795 (N_795,N_691,N_685);
nor U796 (N_796,N_737,N_705);
nor U797 (N_797,N_677,N_707);
nor U798 (N_798,N_739,N_703);
or U799 (N_799,N_746,N_739);
or U800 (N_800,N_694,N_687);
or U801 (N_801,N_677,N_729);
nor U802 (N_802,N_709,N_689);
or U803 (N_803,N_713,N_683);
nand U804 (N_804,N_685,N_696);
or U805 (N_805,N_725,N_685);
nor U806 (N_806,N_705,N_746);
and U807 (N_807,N_676,N_675);
and U808 (N_808,N_740,N_727);
nand U809 (N_809,N_707,N_695);
and U810 (N_810,N_710,N_704);
and U811 (N_811,N_698,N_745);
nand U812 (N_812,N_742,N_708);
nor U813 (N_813,N_710,N_700);
nor U814 (N_814,N_708,N_741);
nand U815 (N_815,N_712,N_685);
or U816 (N_816,N_708,N_733);
nor U817 (N_817,N_705,N_720);
or U818 (N_818,N_737,N_732);
and U819 (N_819,N_731,N_683);
or U820 (N_820,N_741,N_740);
nand U821 (N_821,N_702,N_723);
or U822 (N_822,N_713,N_702);
nor U823 (N_823,N_708,N_718);
xor U824 (N_824,N_721,N_679);
and U825 (N_825,N_804,N_802);
nand U826 (N_826,N_784,N_797);
nand U827 (N_827,N_777,N_791);
and U828 (N_828,N_796,N_789);
nand U829 (N_829,N_755,N_790);
or U830 (N_830,N_793,N_787);
nor U831 (N_831,N_823,N_763);
and U832 (N_832,N_758,N_779);
and U833 (N_833,N_753,N_770);
or U834 (N_834,N_785,N_809);
and U835 (N_835,N_817,N_807);
and U836 (N_836,N_773,N_757);
nor U837 (N_837,N_803,N_780);
and U838 (N_838,N_794,N_762);
and U839 (N_839,N_810,N_805);
or U840 (N_840,N_768,N_750);
or U841 (N_841,N_767,N_759);
nor U842 (N_842,N_756,N_815);
nand U843 (N_843,N_778,N_806);
or U844 (N_844,N_800,N_820);
or U845 (N_845,N_801,N_818);
nor U846 (N_846,N_798,N_782);
or U847 (N_847,N_824,N_822);
nand U848 (N_848,N_783,N_786);
nor U849 (N_849,N_799,N_808);
and U850 (N_850,N_764,N_819);
and U851 (N_851,N_752,N_771);
nor U852 (N_852,N_795,N_821);
and U853 (N_853,N_814,N_769);
or U854 (N_854,N_792,N_775);
nand U855 (N_855,N_751,N_776);
nor U856 (N_856,N_760,N_811);
or U857 (N_857,N_816,N_774);
nor U858 (N_858,N_812,N_761);
nor U859 (N_859,N_766,N_754);
nor U860 (N_860,N_765,N_781);
nor U861 (N_861,N_772,N_788);
nand U862 (N_862,N_813,N_764);
and U863 (N_863,N_792,N_761);
nor U864 (N_864,N_781,N_815);
nand U865 (N_865,N_772,N_767);
or U866 (N_866,N_805,N_803);
nand U867 (N_867,N_792,N_802);
nor U868 (N_868,N_824,N_784);
or U869 (N_869,N_815,N_779);
or U870 (N_870,N_771,N_802);
xor U871 (N_871,N_751,N_788);
and U872 (N_872,N_823,N_795);
nand U873 (N_873,N_791,N_757);
and U874 (N_874,N_778,N_767);
nor U875 (N_875,N_760,N_765);
nor U876 (N_876,N_815,N_813);
and U877 (N_877,N_815,N_757);
and U878 (N_878,N_812,N_820);
and U879 (N_879,N_764,N_783);
or U880 (N_880,N_777,N_812);
or U881 (N_881,N_750,N_779);
or U882 (N_882,N_801,N_808);
nor U883 (N_883,N_822,N_807);
nor U884 (N_884,N_823,N_772);
nand U885 (N_885,N_796,N_807);
and U886 (N_886,N_816,N_777);
nand U887 (N_887,N_816,N_778);
nor U888 (N_888,N_756,N_783);
or U889 (N_889,N_769,N_813);
nand U890 (N_890,N_791,N_781);
nor U891 (N_891,N_784,N_800);
or U892 (N_892,N_764,N_770);
and U893 (N_893,N_796,N_791);
and U894 (N_894,N_757,N_784);
nor U895 (N_895,N_770,N_790);
or U896 (N_896,N_772,N_765);
nor U897 (N_897,N_809,N_754);
nand U898 (N_898,N_777,N_770);
and U899 (N_899,N_775,N_759);
nand U900 (N_900,N_864,N_843);
and U901 (N_901,N_854,N_886);
and U902 (N_902,N_841,N_859);
nand U903 (N_903,N_870,N_894);
nor U904 (N_904,N_869,N_828);
nor U905 (N_905,N_831,N_899);
and U906 (N_906,N_849,N_892);
nor U907 (N_907,N_840,N_871);
nor U908 (N_908,N_856,N_826);
and U909 (N_909,N_891,N_834);
and U910 (N_910,N_874,N_845);
nand U911 (N_911,N_827,N_830);
nand U912 (N_912,N_868,N_885);
nor U913 (N_913,N_895,N_897);
nor U914 (N_914,N_873,N_860);
nor U915 (N_915,N_887,N_836);
nand U916 (N_916,N_855,N_842);
and U917 (N_917,N_884,N_880);
or U918 (N_918,N_846,N_829);
nand U919 (N_919,N_853,N_852);
nor U920 (N_920,N_857,N_882);
or U921 (N_921,N_893,N_862);
nand U922 (N_922,N_865,N_839);
nand U923 (N_923,N_825,N_861);
nand U924 (N_924,N_876,N_890);
nor U925 (N_925,N_838,N_867);
nand U926 (N_926,N_847,N_863);
nor U927 (N_927,N_844,N_879);
nand U928 (N_928,N_898,N_833);
and U929 (N_929,N_837,N_878);
nor U930 (N_930,N_875,N_896);
nand U931 (N_931,N_832,N_877);
nor U932 (N_932,N_851,N_835);
nor U933 (N_933,N_889,N_848);
and U934 (N_934,N_850,N_858);
nor U935 (N_935,N_881,N_888);
nand U936 (N_936,N_883,N_866);
or U937 (N_937,N_872,N_868);
or U938 (N_938,N_885,N_827);
nand U939 (N_939,N_847,N_868);
or U940 (N_940,N_863,N_876);
and U941 (N_941,N_851,N_878);
and U942 (N_942,N_869,N_866);
and U943 (N_943,N_831,N_898);
nor U944 (N_944,N_844,N_866);
nor U945 (N_945,N_858,N_867);
or U946 (N_946,N_843,N_887);
and U947 (N_947,N_869,N_832);
nor U948 (N_948,N_838,N_895);
nor U949 (N_949,N_855,N_888);
nand U950 (N_950,N_849,N_867);
nor U951 (N_951,N_852,N_890);
nor U952 (N_952,N_847,N_862);
nor U953 (N_953,N_826,N_896);
and U954 (N_954,N_899,N_837);
or U955 (N_955,N_840,N_857);
nand U956 (N_956,N_874,N_842);
or U957 (N_957,N_861,N_863);
nand U958 (N_958,N_880,N_841);
or U959 (N_959,N_871,N_843);
nor U960 (N_960,N_825,N_831);
nand U961 (N_961,N_875,N_886);
or U962 (N_962,N_849,N_851);
nand U963 (N_963,N_868,N_846);
nor U964 (N_964,N_867,N_888);
nor U965 (N_965,N_891,N_844);
nor U966 (N_966,N_861,N_850);
nor U967 (N_967,N_826,N_895);
and U968 (N_968,N_875,N_889);
or U969 (N_969,N_872,N_838);
and U970 (N_970,N_848,N_845);
nand U971 (N_971,N_856,N_883);
nand U972 (N_972,N_846,N_832);
nand U973 (N_973,N_851,N_841);
and U974 (N_974,N_899,N_858);
nor U975 (N_975,N_934,N_935);
nor U976 (N_976,N_943,N_960);
nor U977 (N_977,N_967,N_928);
and U978 (N_978,N_955,N_945);
or U979 (N_979,N_954,N_925);
nand U980 (N_980,N_913,N_917);
nor U981 (N_981,N_900,N_939);
nand U982 (N_982,N_937,N_911);
and U983 (N_983,N_970,N_966);
and U984 (N_984,N_974,N_958);
nand U985 (N_985,N_963,N_959);
or U986 (N_986,N_918,N_949);
nor U987 (N_987,N_936,N_901);
nand U988 (N_988,N_968,N_903);
and U989 (N_989,N_919,N_971);
or U990 (N_990,N_946,N_910);
or U991 (N_991,N_957,N_941);
nand U992 (N_992,N_938,N_953);
or U993 (N_993,N_929,N_920);
or U994 (N_994,N_961,N_950);
xor U995 (N_995,N_940,N_914);
or U996 (N_996,N_922,N_973);
or U997 (N_997,N_942,N_965);
nor U998 (N_998,N_909,N_923);
and U999 (N_999,N_932,N_972);
nand U1000 (N_1000,N_962,N_912);
or U1001 (N_1001,N_921,N_931);
or U1002 (N_1002,N_904,N_969);
and U1003 (N_1003,N_951,N_927);
and U1004 (N_1004,N_947,N_930);
or U1005 (N_1005,N_905,N_956);
or U1006 (N_1006,N_944,N_924);
and U1007 (N_1007,N_952,N_948);
or U1008 (N_1008,N_906,N_964);
nor U1009 (N_1009,N_902,N_933);
nor U1010 (N_1010,N_915,N_926);
nor U1011 (N_1011,N_907,N_916);
nand U1012 (N_1012,N_908,N_919);
and U1013 (N_1013,N_958,N_912);
nor U1014 (N_1014,N_922,N_963);
or U1015 (N_1015,N_968,N_947);
and U1016 (N_1016,N_902,N_963);
and U1017 (N_1017,N_913,N_944);
or U1018 (N_1018,N_957,N_945);
nor U1019 (N_1019,N_954,N_932);
and U1020 (N_1020,N_956,N_911);
nand U1021 (N_1021,N_926,N_959);
and U1022 (N_1022,N_963,N_950);
nor U1023 (N_1023,N_916,N_906);
or U1024 (N_1024,N_918,N_906);
and U1025 (N_1025,N_951,N_919);
nor U1026 (N_1026,N_911,N_912);
or U1027 (N_1027,N_912,N_901);
nand U1028 (N_1028,N_916,N_908);
or U1029 (N_1029,N_909,N_973);
or U1030 (N_1030,N_935,N_908);
or U1031 (N_1031,N_956,N_925);
and U1032 (N_1032,N_936,N_932);
and U1033 (N_1033,N_956,N_914);
nand U1034 (N_1034,N_907,N_905);
and U1035 (N_1035,N_944,N_961);
and U1036 (N_1036,N_908,N_948);
and U1037 (N_1037,N_922,N_943);
and U1038 (N_1038,N_937,N_957);
and U1039 (N_1039,N_906,N_948);
nand U1040 (N_1040,N_938,N_925);
or U1041 (N_1041,N_945,N_924);
nand U1042 (N_1042,N_903,N_951);
xnor U1043 (N_1043,N_919,N_928);
xnor U1044 (N_1044,N_973,N_929);
nor U1045 (N_1045,N_925,N_936);
or U1046 (N_1046,N_965,N_961);
and U1047 (N_1047,N_921,N_901);
and U1048 (N_1048,N_911,N_961);
and U1049 (N_1049,N_913,N_953);
nor U1050 (N_1050,N_981,N_1014);
and U1051 (N_1051,N_1003,N_1011);
nor U1052 (N_1052,N_1023,N_1041);
and U1053 (N_1053,N_1026,N_1036);
and U1054 (N_1054,N_1017,N_1001);
or U1055 (N_1055,N_1000,N_984);
and U1056 (N_1056,N_975,N_989);
or U1057 (N_1057,N_1016,N_979);
and U1058 (N_1058,N_1047,N_1018);
nor U1059 (N_1059,N_993,N_1024);
and U1060 (N_1060,N_1021,N_997);
and U1061 (N_1061,N_990,N_988);
nand U1062 (N_1062,N_1012,N_980);
and U1063 (N_1063,N_1022,N_1048);
and U1064 (N_1064,N_1015,N_1045);
nor U1065 (N_1065,N_998,N_1040);
or U1066 (N_1066,N_1044,N_1007);
nor U1067 (N_1067,N_1025,N_1020);
or U1068 (N_1068,N_1010,N_1009);
nor U1069 (N_1069,N_1043,N_1039);
nor U1070 (N_1070,N_1034,N_982);
and U1071 (N_1071,N_1049,N_978);
nor U1072 (N_1072,N_1033,N_976);
and U1073 (N_1073,N_1038,N_1037);
nor U1074 (N_1074,N_1032,N_991);
nor U1075 (N_1075,N_1006,N_985);
and U1076 (N_1076,N_987,N_1029);
nor U1077 (N_1077,N_1004,N_977);
nor U1078 (N_1078,N_992,N_1042);
nand U1079 (N_1079,N_996,N_1046);
and U1080 (N_1080,N_1028,N_1013);
or U1081 (N_1081,N_1035,N_999);
nor U1082 (N_1082,N_994,N_1005);
nand U1083 (N_1083,N_983,N_1030);
nand U1084 (N_1084,N_986,N_1027);
nand U1085 (N_1085,N_1031,N_1002);
and U1086 (N_1086,N_1019,N_995);
and U1087 (N_1087,N_1008,N_995);
nand U1088 (N_1088,N_1026,N_1003);
nor U1089 (N_1089,N_1002,N_1005);
or U1090 (N_1090,N_999,N_1018);
nor U1091 (N_1091,N_1006,N_994);
nor U1092 (N_1092,N_995,N_1015);
nor U1093 (N_1093,N_1008,N_987);
or U1094 (N_1094,N_991,N_1008);
or U1095 (N_1095,N_980,N_1002);
or U1096 (N_1096,N_1027,N_981);
and U1097 (N_1097,N_1028,N_1033);
or U1098 (N_1098,N_1019,N_1039);
nand U1099 (N_1099,N_979,N_1040);
or U1100 (N_1100,N_1023,N_1003);
or U1101 (N_1101,N_1028,N_995);
nand U1102 (N_1102,N_1032,N_978);
and U1103 (N_1103,N_1027,N_1048);
nor U1104 (N_1104,N_1021,N_1025);
or U1105 (N_1105,N_1002,N_991);
and U1106 (N_1106,N_991,N_1035);
and U1107 (N_1107,N_1012,N_1025);
nor U1108 (N_1108,N_983,N_1001);
nand U1109 (N_1109,N_1012,N_1031);
and U1110 (N_1110,N_994,N_1003);
or U1111 (N_1111,N_1034,N_978);
and U1112 (N_1112,N_988,N_1036);
nor U1113 (N_1113,N_978,N_1000);
nand U1114 (N_1114,N_1002,N_1039);
nand U1115 (N_1115,N_1037,N_996);
and U1116 (N_1116,N_1014,N_975);
nand U1117 (N_1117,N_1008,N_1034);
nor U1118 (N_1118,N_1033,N_1022);
and U1119 (N_1119,N_990,N_981);
nor U1120 (N_1120,N_975,N_1038);
and U1121 (N_1121,N_1032,N_992);
and U1122 (N_1122,N_1004,N_1042);
nand U1123 (N_1123,N_1020,N_987);
and U1124 (N_1124,N_984,N_1043);
nor U1125 (N_1125,N_1064,N_1051);
or U1126 (N_1126,N_1083,N_1118);
nand U1127 (N_1127,N_1111,N_1088);
nor U1128 (N_1128,N_1065,N_1109);
and U1129 (N_1129,N_1057,N_1097);
nand U1130 (N_1130,N_1085,N_1089);
nand U1131 (N_1131,N_1073,N_1055);
nor U1132 (N_1132,N_1120,N_1062);
or U1133 (N_1133,N_1092,N_1071);
and U1134 (N_1134,N_1114,N_1074);
nand U1135 (N_1135,N_1122,N_1061);
nand U1136 (N_1136,N_1087,N_1081);
or U1137 (N_1137,N_1121,N_1091);
nand U1138 (N_1138,N_1116,N_1124);
nand U1139 (N_1139,N_1054,N_1094);
and U1140 (N_1140,N_1093,N_1108);
nor U1141 (N_1141,N_1105,N_1076);
nor U1142 (N_1142,N_1086,N_1075);
and U1143 (N_1143,N_1101,N_1079);
nand U1144 (N_1144,N_1100,N_1107);
nor U1145 (N_1145,N_1069,N_1082);
nor U1146 (N_1146,N_1059,N_1050);
nand U1147 (N_1147,N_1103,N_1058);
or U1148 (N_1148,N_1123,N_1106);
nand U1149 (N_1149,N_1056,N_1096);
nor U1150 (N_1150,N_1070,N_1066);
nand U1151 (N_1151,N_1060,N_1104);
nand U1152 (N_1152,N_1067,N_1068);
nor U1153 (N_1153,N_1099,N_1078);
and U1154 (N_1154,N_1053,N_1110);
or U1155 (N_1155,N_1077,N_1119);
or U1156 (N_1156,N_1102,N_1112);
and U1157 (N_1157,N_1090,N_1084);
nand U1158 (N_1158,N_1098,N_1063);
nor U1159 (N_1159,N_1052,N_1095);
or U1160 (N_1160,N_1072,N_1113);
nand U1161 (N_1161,N_1117,N_1080);
nand U1162 (N_1162,N_1115,N_1064);
or U1163 (N_1163,N_1068,N_1057);
nand U1164 (N_1164,N_1118,N_1063);
and U1165 (N_1165,N_1088,N_1052);
or U1166 (N_1166,N_1092,N_1079);
or U1167 (N_1167,N_1051,N_1057);
nor U1168 (N_1168,N_1096,N_1074);
and U1169 (N_1169,N_1070,N_1114);
nor U1170 (N_1170,N_1079,N_1124);
or U1171 (N_1171,N_1061,N_1060);
nand U1172 (N_1172,N_1087,N_1096);
nor U1173 (N_1173,N_1120,N_1081);
nand U1174 (N_1174,N_1089,N_1058);
and U1175 (N_1175,N_1114,N_1101);
and U1176 (N_1176,N_1108,N_1111);
nand U1177 (N_1177,N_1105,N_1089);
or U1178 (N_1178,N_1053,N_1063);
or U1179 (N_1179,N_1093,N_1110);
or U1180 (N_1180,N_1084,N_1070);
nand U1181 (N_1181,N_1082,N_1090);
or U1182 (N_1182,N_1107,N_1089);
or U1183 (N_1183,N_1050,N_1060);
nor U1184 (N_1184,N_1095,N_1088);
and U1185 (N_1185,N_1072,N_1075);
nor U1186 (N_1186,N_1065,N_1105);
and U1187 (N_1187,N_1089,N_1108);
or U1188 (N_1188,N_1071,N_1076);
or U1189 (N_1189,N_1100,N_1063);
or U1190 (N_1190,N_1097,N_1112);
and U1191 (N_1191,N_1060,N_1083);
or U1192 (N_1192,N_1107,N_1070);
or U1193 (N_1193,N_1081,N_1118);
nor U1194 (N_1194,N_1078,N_1061);
or U1195 (N_1195,N_1068,N_1073);
and U1196 (N_1196,N_1120,N_1085);
nor U1197 (N_1197,N_1051,N_1053);
nor U1198 (N_1198,N_1117,N_1085);
or U1199 (N_1199,N_1089,N_1116);
nand U1200 (N_1200,N_1127,N_1163);
or U1201 (N_1201,N_1140,N_1125);
and U1202 (N_1202,N_1192,N_1194);
and U1203 (N_1203,N_1141,N_1135);
nand U1204 (N_1204,N_1158,N_1197);
nor U1205 (N_1205,N_1130,N_1153);
nand U1206 (N_1206,N_1162,N_1169);
and U1207 (N_1207,N_1170,N_1182);
nand U1208 (N_1208,N_1176,N_1160);
nor U1209 (N_1209,N_1172,N_1188);
xor U1210 (N_1210,N_1173,N_1132);
nand U1211 (N_1211,N_1144,N_1198);
and U1212 (N_1212,N_1161,N_1164);
and U1213 (N_1213,N_1168,N_1171);
nor U1214 (N_1214,N_1143,N_1181);
and U1215 (N_1215,N_1138,N_1147);
nor U1216 (N_1216,N_1155,N_1145);
nand U1217 (N_1217,N_1159,N_1193);
or U1218 (N_1218,N_1167,N_1189);
and U1219 (N_1219,N_1131,N_1184);
or U1220 (N_1220,N_1134,N_1152);
nand U1221 (N_1221,N_1154,N_1136);
nand U1222 (N_1222,N_1137,N_1175);
and U1223 (N_1223,N_1190,N_1151);
and U1224 (N_1224,N_1191,N_1165);
or U1225 (N_1225,N_1150,N_1195);
nand U1226 (N_1226,N_1129,N_1177);
and U1227 (N_1227,N_1183,N_1149);
and U1228 (N_1228,N_1185,N_1179);
nand U1229 (N_1229,N_1156,N_1187);
nand U1230 (N_1230,N_1166,N_1196);
nand U1231 (N_1231,N_1146,N_1126);
or U1232 (N_1232,N_1133,N_1186);
or U1233 (N_1233,N_1157,N_1178);
and U1234 (N_1234,N_1128,N_1180);
nor U1235 (N_1235,N_1148,N_1199);
nor U1236 (N_1236,N_1139,N_1174);
or U1237 (N_1237,N_1142,N_1196);
or U1238 (N_1238,N_1185,N_1176);
or U1239 (N_1239,N_1186,N_1181);
nand U1240 (N_1240,N_1134,N_1174);
xor U1241 (N_1241,N_1159,N_1162);
or U1242 (N_1242,N_1135,N_1144);
nor U1243 (N_1243,N_1152,N_1151);
or U1244 (N_1244,N_1152,N_1169);
or U1245 (N_1245,N_1193,N_1154);
or U1246 (N_1246,N_1149,N_1194);
nand U1247 (N_1247,N_1188,N_1134);
and U1248 (N_1248,N_1134,N_1182);
nand U1249 (N_1249,N_1167,N_1160);
or U1250 (N_1250,N_1145,N_1181);
and U1251 (N_1251,N_1172,N_1152);
nor U1252 (N_1252,N_1170,N_1135);
and U1253 (N_1253,N_1147,N_1150);
or U1254 (N_1254,N_1195,N_1129);
and U1255 (N_1255,N_1153,N_1174);
nand U1256 (N_1256,N_1140,N_1164);
and U1257 (N_1257,N_1192,N_1161);
and U1258 (N_1258,N_1172,N_1171);
nand U1259 (N_1259,N_1192,N_1157);
and U1260 (N_1260,N_1197,N_1178);
or U1261 (N_1261,N_1180,N_1193);
nand U1262 (N_1262,N_1184,N_1169);
or U1263 (N_1263,N_1146,N_1133);
nand U1264 (N_1264,N_1149,N_1166);
or U1265 (N_1265,N_1137,N_1193);
nor U1266 (N_1266,N_1182,N_1175);
nor U1267 (N_1267,N_1144,N_1136);
xnor U1268 (N_1268,N_1130,N_1143);
xnor U1269 (N_1269,N_1139,N_1195);
or U1270 (N_1270,N_1137,N_1156);
nor U1271 (N_1271,N_1177,N_1176);
or U1272 (N_1272,N_1179,N_1144);
nor U1273 (N_1273,N_1132,N_1126);
or U1274 (N_1274,N_1127,N_1169);
nor U1275 (N_1275,N_1264,N_1236);
and U1276 (N_1276,N_1240,N_1223);
or U1277 (N_1277,N_1226,N_1224);
and U1278 (N_1278,N_1234,N_1247);
nand U1279 (N_1279,N_1266,N_1273);
nor U1280 (N_1280,N_1213,N_1246);
nand U1281 (N_1281,N_1255,N_1259);
or U1282 (N_1282,N_1248,N_1204);
nor U1283 (N_1283,N_1258,N_1239);
nand U1284 (N_1284,N_1260,N_1257);
and U1285 (N_1285,N_1211,N_1237);
nand U1286 (N_1286,N_1262,N_1227);
nand U1287 (N_1287,N_1235,N_1209);
nor U1288 (N_1288,N_1201,N_1212);
or U1289 (N_1289,N_1202,N_1261);
or U1290 (N_1290,N_1215,N_1205);
nand U1291 (N_1291,N_1217,N_1263);
nand U1292 (N_1292,N_1216,N_1203);
nor U1293 (N_1293,N_1252,N_1231);
and U1294 (N_1294,N_1265,N_1268);
nand U1295 (N_1295,N_1210,N_1256);
or U1296 (N_1296,N_1230,N_1222);
nor U1297 (N_1297,N_1274,N_1270);
or U1298 (N_1298,N_1267,N_1244);
and U1299 (N_1299,N_1272,N_1269);
and U1300 (N_1300,N_1229,N_1238);
or U1301 (N_1301,N_1242,N_1220);
nand U1302 (N_1302,N_1207,N_1271);
nand U1303 (N_1303,N_1250,N_1200);
and U1304 (N_1304,N_1232,N_1243);
or U1305 (N_1305,N_1221,N_1254);
nand U1306 (N_1306,N_1206,N_1233);
or U1307 (N_1307,N_1253,N_1218);
nor U1308 (N_1308,N_1225,N_1241);
nand U1309 (N_1309,N_1219,N_1249);
or U1310 (N_1310,N_1228,N_1245);
nand U1311 (N_1311,N_1251,N_1214);
nand U1312 (N_1312,N_1208,N_1218);
or U1313 (N_1313,N_1211,N_1264);
or U1314 (N_1314,N_1260,N_1221);
or U1315 (N_1315,N_1207,N_1223);
nor U1316 (N_1316,N_1237,N_1256);
or U1317 (N_1317,N_1268,N_1233);
and U1318 (N_1318,N_1206,N_1250);
and U1319 (N_1319,N_1250,N_1218);
and U1320 (N_1320,N_1251,N_1259);
and U1321 (N_1321,N_1252,N_1256);
or U1322 (N_1322,N_1210,N_1242);
and U1323 (N_1323,N_1218,N_1266);
or U1324 (N_1324,N_1244,N_1228);
nor U1325 (N_1325,N_1222,N_1224);
nand U1326 (N_1326,N_1270,N_1221);
nor U1327 (N_1327,N_1274,N_1235);
nor U1328 (N_1328,N_1207,N_1244);
nand U1329 (N_1329,N_1204,N_1263);
and U1330 (N_1330,N_1223,N_1248);
or U1331 (N_1331,N_1250,N_1202);
xnor U1332 (N_1332,N_1232,N_1203);
or U1333 (N_1333,N_1265,N_1207);
nand U1334 (N_1334,N_1246,N_1240);
and U1335 (N_1335,N_1242,N_1246);
nand U1336 (N_1336,N_1214,N_1204);
and U1337 (N_1337,N_1212,N_1214);
nor U1338 (N_1338,N_1222,N_1212);
and U1339 (N_1339,N_1255,N_1228);
and U1340 (N_1340,N_1222,N_1221);
and U1341 (N_1341,N_1254,N_1207);
nor U1342 (N_1342,N_1255,N_1252);
nor U1343 (N_1343,N_1211,N_1265);
or U1344 (N_1344,N_1204,N_1231);
and U1345 (N_1345,N_1209,N_1231);
nor U1346 (N_1346,N_1234,N_1229);
and U1347 (N_1347,N_1231,N_1242);
nor U1348 (N_1348,N_1248,N_1249);
nand U1349 (N_1349,N_1262,N_1263);
nor U1350 (N_1350,N_1302,N_1295);
nand U1351 (N_1351,N_1299,N_1325);
and U1352 (N_1352,N_1337,N_1339);
nor U1353 (N_1353,N_1324,N_1290);
xor U1354 (N_1354,N_1326,N_1284);
or U1355 (N_1355,N_1298,N_1346);
and U1356 (N_1356,N_1309,N_1280);
or U1357 (N_1357,N_1320,N_1303);
and U1358 (N_1358,N_1322,N_1317);
nor U1359 (N_1359,N_1286,N_1316);
nor U1360 (N_1360,N_1301,N_1341);
and U1361 (N_1361,N_1310,N_1342);
or U1362 (N_1362,N_1311,N_1327);
and U1363 (N_1363,N_1313,N_1277);
and U1364 (N_1364,N_1335,N_1276);
nor U1365 (N_1365,N_1312,N_1292);
nor U1366 (N_1366,N_1336,N_1278);
nand U1367 (N_1367,N_1300,N_1330);
nand U1368 (N_1368,N_1285,N_1305);
nand U1369 (N_1369,N_1291,N_1340);
nor U1370 (N_1370,N_1347,N_1314);
nand U1371 (N_1371,N_1321,N_1283);
and U1372 (N_1372,N_1323,N_1293);
or U1373 (N_1373,N_1279,N_1304);
nand U1374 (N_1374,N_1328,N_1315);
nand U1375 (N_1375,N_1334,N_1348);
xor U1376 (N_1376,N_1289,N_1288);
or U1377 (N_1377,N_1294,N_1344);
nand U1378 (N_1378,N_1332,N_1297);
and U1379 (N_1379,N_1345,N_1319);
nor U1380 (N_1380,N_1275,N_1329);
and U1381 (N_1381,N_1296,N_1343);
or U1382 (N_1382,N_1349,N_1307);
or U1383 (N_1383,N_1282,N_1287);
or U1384 (N_1384,N_1308,N_1333);
or U1385 (N_1385,N_1338,N_1318);
nor U1386 (N_1386,N_1281,N_1306);
nand U1387 (N_1387,N_1331,N_1288);
or U1388 (N_1388,N_1325,N_1307);
and U1389 (N_1389,N_1307,N_1336);
or U1390 (N_1390,N_1308,N_1305);
or U1391 (N_1391,N_1284,N_1340);
nand U1392 (N_1392,N_1330,N_1319);
and U1393 (N_1393,N_1295,N_1303);
or U1394 (N_1394,N_1287,N_1275);
and U1395 (N_1395,N_1295,N_1346);
nand U1396 (N_1396,N_1315,N_1344);
or U1397 (N_1397,N_1340,N_1282);
nand U1398 (N_1398,N_1295,N_1277);
and U1399 (N_1399,N_1319,N_1328);
or U1400 (N_1400,N_1333,N_1295);
nor U1401 (N_1401,N_1337,N_1307);
and U1402 (N_1402,N_1290,N_1327);
and U1403 (N_1403,N_1295,N_1345);
nand U1404 (N_1404,N_1320,N_1302);
nand U1405 (N_1405,N_1278,N_1342);
nor U1406 (N_1406,N_1277,N_1345);
and U1407 (N_1407,N_1308,N_1346);
nor U1408 (N_1408,N_1347,N_1342);
and U1409 (N_1409,N_1309,N_1324);
and U1410 (N_1410,N_1327,N_1299);
and U1411 (N_1411,N_1344,N_1317);
and U1412 (N_1412,N_1335,N_1278);
nand U1413 (N_1413,N_1311,N_1313);
nand U1414 (N_1414,N_1335,N_1347);
nand U1415 (N_1415,N_1324,N_1305);
nand U1416 (N_1416,N_1283,N_1304);
or U1417 (N_1417,N_1334,N_1284);
or U1418 (N_1418,N_1342,N_1345);
and U1419 (N_1419,N_1281,N_1280);
nand U1420 (N_1420,N_1300,N_1341);
nor U1421 (N_1421,N_1308,N_1349);
and U1422 (N_1422,N_1305,N_1304);
nor U1423 (N_1423,N_1339,N_1296);
nor U1424 (N_1424,N_1310,N_1296);
xnor U1425 (N_1425,N_1414,N_1407);
nor U1426 (N_1426,N_1365,N_1409);
or U1427 (N_1427,N_1405,N_1396);
nand U1428 (N_1428,N_1372,N_1421);
nor U1429 (N_1429,N_1406,N_1415);
or U1430 (N_1430,N_1410,N_1361);
xnor U1431 (N_1431,N_1364,N_1419);
nor U1432 (N_1432,N_1418,N_1355);
and U1433 (N_1433,N_1362,N_1350);
or U1434 (N_1434,N_1371,N_1402);
nor U1435 (N_1435,N_1351,N_1399);
and U1436 (N_1436,N_1375,N_1369);
and U1437 (N_1437,N_1356,N_1408);
and U1438 (N_1438,N_1383,N_1404);
and U1439 (N_1439,N_1380,N_1368);
nor U1440 (N_1440,N_1403,N_1422);
or U1441 (N_1441,N_1416,N_1395);
nor U1442 (N_1442,N_1378,N_1393);
or U1443 (N_1443,N_1420,N_1417);
and U1444 (N_1444,N_1413,N_1357);
nand U1445 (N_1445,N_1423,N_1359);
or U1446 (N_1446,N_1382,N_1424);
nor U1447 (N_1447,N_1389,N_1386);
nand U1448 (N_1448,N_1377,N_1398);
or U1449 (N_1449,N_1374,N_1366);
nor U1450 (N_1450,N_1367,N_1388);
and U1451 (N_1451,N_1392,N_1354);
nor U1452 (N_1452,N_1363,N_1353);
nand U1453 (N_1453,N_1390,N_1360);
and U1454 (N_1454,N_1376,N_1352);
nand U1455 (N_1455,N_1381,N_1412);
or U1456 (N_1456,N_1400,N_1411);
nor U1457 (N_1457,N_1373,N_1401);
and U1458 (N_1458,N_1397,N_1358);
and U1459 (N_1459,N_1370,N_1385);
nand U1460 (N_1460,N_1394,N_1384);
or U1461 (N_1461,N_1387,N_1391);
nor U1462 (N_1462,N_1379,N_1382);
or U1463 (N_1463,N_1375,N_1365);
nand U1464 (N_1464,N_1414,N_1406);
and U1465 (N_1465,N_1422,N_1388);
and U1466 (N_1466,N_1419,N_1418);
nand U1467 (N_1467,N_1394,N_1385);
nor U1468 (N_1468,N_1380,N_1420);
and U1469 (N_1469,N_1422,N_1411);
xnor U1470 (N_1470,N_1408,N_1372);
and U1471 (N_1471,N_1355,N_1352);
xnor U1472 (N_1472,N_1382,N_1414);
and U1473 (N_1473,N_1350,N_1366);
nand U1474 (N_1474,N_1416,N_1393);
nand U1475 (N_1475,N_1417,N_1375);
xnor U1476 (N_1476,N_1374,N_1388);
and U1477 (N_1477,N_1422,N_1417);
and U1478 (N_1478,N_1394,N_1395);
and U1479 (N_1479,N_1421,N_1382);
nor U1480 (N_1480,N_1424,N_1404);
or U1481 (N_1481,N_1357,N_1359);
or U1482 (N_1482,N_1362,N_1422);
nor U1483 (N_1483,N_1387,N_1381);
nor U1484 (N_1484,N_1361,N_1365);
nor U1485 (N_1485,N_1396,N_1364);
or U1486 (N_1486,N_1397,N_1392);
nand U1487 (N_1487,N_1365,N_1395);
or U1488 (N_1488,N_1358,N_1375);
and U1489 (N_1489,N_1356,N_1378);
or U1490 (N_1490,N_1409,N_1355);
nor U1491 (N_1491,N_1398,N_1373);
or U1492 (N_1492,N_1355,N_1405);
or U1493 (N_1493,N_1416,N_1355);
nand U1494 (N_1494,N_1370,N_1371);
xor U1495 (N_1495,N_1353,N_1406);
nand U1496 (N_1496,N_1380,N_1361);
and U1497 (N_1497,N_1399,N_1392);
nand U1498 (N_1498,N_1376,N_1390);
or U1499 (N_1499,N_1378,N_1411);
nor U1500 (N_1500,N_1483,N_1461);
and U1501 (N_1501,N_1469,N_1465);
or U1502 (N_1502,N_1439,N_1467);
nand U1503 (N_1503,N_1444,N_1449);
and U1504 (N_1504,N_1491,N_1470);
nor U1505 (N_1505,N_1446,N_1497);
nand U1506 (N_1506,N_1478,N_1482);
or U1507 (N_1507,N_1442,N_1476);
and U1508 (N_1508,N_1448,N_1487);
nor U1509 (N_1509,N_1447,N_1485);
or U1510 (N_1510,N_1489,N_1450);
or U1511 (N_1511,N_1432,N_1425);
nor U1512 (N_1512,N_1434,N_1438);
nand U1513 (N_1513,N_1486,N_1427);
nor U1514 (N_1514,N_1480,N_1431);
and U1515 (N_1515,N_1436,N_1435);
nor U1516 (N_1516,N_1456,N_1466);
or U1517 (N_1517,N_1428,N_1490);
nor U1518 (N_1518,N_1468,N_1426);
nand U1519 (N_1519,N_1493,N_1437);
nor U1520 (N_1520,N_1445,N_1484);
and U1521 (N_1521,N_1481,N_1488);
and U1522 (N_1522,N_1477,N_1451);
nand U1523 (N_1523,N_1440,N_1457);
nand U1524 (N_1524,N_1475,N_1454);
nor U1525 (N_1525,N_1462,N_1499);
or U1526 (N_1526,N_1459,N_1460);
and U1527 (N_1527,N_1452,N_1433);
nand U1528 (N_1528,N_1472,N_1463);
nor U1529 (N_1529,N_1496,N_1443);
and U1530 (N_1530,N_1473,N_1492);
nand U1531 (N_1531,N_1455,N_1453);
nor U1532 (N_1532,N_1494,N_1458);
nor U1533 (N_1533,N_1471,N_1479);
and U1534 (N_1534,N_1441,N_1495);
nand U1535 (N_1535,N_1430,N_1429);
nor U1536 (N_1536,N_1474,N_1498);
nand U1537 (N_1537,N_1464,N_1445);
and U1538 (N_1538,N_1433,N_1459);
and U1539 (N_1539,N_1467,N_1469);
nand U1540 (N_1540,N_1455,N_1463);
nor U1541 (N_1541,N_1440,N_1479);
nand U1542 (N_1542,N_1471,N_1436);
nor U1543 (N_1543,N_1477,N_1470);
and U1544 (N_1544,N_1480,N_1466);
nor U1545 (N_1545,N_1441,N_1463);
nor U1546 (N_1546,N_1492,N_1430);
nand U1547 (N_1547,N_1465,N_1483);
nand U1548 (N_1548,N_1454,N_1456);
nand U1549 (N_1549,N_1436,N_1437);
nand U1550 (N_1550,N_1474,N_1453);
nand U1551 (N_1551,N_1450,N_1452);
or U1552 (N_1552,N_1427,N_1470);
nor U1553 (N_1553,N_1460,N_1495);
and U1554 (N_1554,N_1425,N_1492);
nor U1555 (N_1555,N_1481,N_1433);
or U1556 (N_1556,N_1472,N_1431);
and U1557 (N_1557,N_1440,N_1456);
nand U1558 (N_1558,N_1483,N_1474);
and U1559 (N_1559,N_1480,N_1470);
nand U1560 (N_1560,N_1437,N_1449);
xor U1561 (N_1561,N_1429,N_1426);
nand U1562 (N_1562,N_1499,N_1433);
and U1563 (N_1563,N_1456,N_1483);
nor U1564 (N_1564,N_1452,N_1427);
nor U1565 (N_1565,N_1486,N_1491);
or U1566 (N_1566,N_1496,N_1463);
and U1567 (N_1567,N_1463,N_1436);
nand U1568 (N_1568,N_1473,N_1476);
and U1569 (N_1569,N_1441,N_1446);
nor U1570 (N_1570,N_1443,N_1482);
nor U1571 (N_1571,N_1498,N_1482);
nand U1572 (N_1572,N_1491,N_1427);
nor U1573 (N_1573,N_1429,N_1482);
nor U1574 (N_1574,N_1444,N_1438);
nor U1575 (N_1575,N_1564,N_1507);
and U1576 (N_1576,N_1573,N_1541);
nand U1577 (N_1577,N_1550,N_1508);
or U1578 (N_1578,N_1533,N_1520);
nand U1579 (N_1579,N_1537,N_1523);
nor U1580 (N_1580,N_1558,N_1571);
or U1581 (N_1581,N_1549,N_1538);
or U1582 (N_1582,N_1511,N_1551);
or U1583 (N_1583,N_1522,N_1529);
nand U1584 (N_1584,N_1552,N_1524);
nor U1585 (N_1585,N_1502,N_1559);
or U1586 (N_1586,N_1509,N_1544);
or U1587 (N_1587,N_1547,N_1556);
nand U1588 (N_1588,N_1553,N_1535);
nor U1589 (N_1589,N_1501,N_1521);
nand U1590 (N_1590,N_1527,N_1512);
nor U1591 (N_1591,N_1572,N_1560);
nor U1592 (N_1592,N_1510,N_1534);
nor U1593 (N_1593,N_1528,N_1543);
and U1594 (N_1594,N_1531,N_1506);
or U1595 (N_1595,N_1503,N_1526);
and U1596 (N_1596,N_1536,N_1532);
nor U1597 (N_1597,N_1540,N_1518);
and U1598 (N_1598,N_1563,N_1557);
nand U1599 (N_1599,N_1562,N_1505);
and U1600 (N_1600,N_1567,N_1546);
or U1601 (N_1601,N_1555,N_1568);
nor U1602 (N_1602,N_1570,N_1504);
nor U1603 (N_1603,N_1519,N_1514);
or U1604 (N_1604,N_1561,N_1517);
nor U1605 (N_1605,N_1569,N_1530);
or U1606 (N_1606,N_1516,N_1545);
nor U1607 (N_1607,N_1513,N_1574);
or U1608 (N_1608,N_1566,N_1542);
or U1609 (N_1609,N_1548,N_1515);
and U1610 (N_1610,N_1565,N_1539);
nor U1611 (N_1611,N_1554,N_1525);
nor U1612 (N_1612,N_1500,N_1505);
nor U1613 (N_1613,N_1502,N_1501);
and U1614 (N_1614,N_1517,N_1507);
nor U1615 (N_1615,N_1570,N_1574);
and U1616 (N_1616,N_1529,N_1525);
or U1617 (N_1617,N_1523,N_1530);
nor U1618 (N_1618,N_1531,N_1507);
or U1619 (N_1619,N_1526,N_1564);
or U1620 (N_1620,N_1560,N_1506);
and U1621 (N_1621,N_1540,N_1557);
nand U1622 (N_1622,N_1516,N_1544);
nand U1623 (N_1623,N_1550,N_1558);
nor U1624 (N_1624,N_1539,N_1517);
xor U1625 (N_1625,N_1516,N_1558);
nor U1626 (N_1626,N_1560,N_1538);
nand U1627 (N_1627,N_1552,N_1572);
nor U1628 (N_1628,N_1559,N_1508);
or U1629 (N_1629,N_1571,N_1534);
nand U1630 (N_1630,N_1551,N_1540);
or U1631 (N_1631,N_1546,N_1516);
xor U1632 (N_1632,N_1505,N_1536);
nand U1633 (N_1633,N_1550,N_1570);
and U1634 (N_1634,N_1538,N_1564);
xor U1635 (N_1635,N_1524,N_1523);
or U1636 (N_1636,N_1572,N_1551);
nand U1637 (N_1637,N_1513,N_1558);
and U1638 (N_1638,N_1524,N_1512);
or U1639 (N_1639,N_1520,N_1529);
and U1640 (N_1640,N_1509,N_1557);
and U1641 (N_1641,N_1546,N_1518);
nand U1642 (N_1642,N_1574,N_1544);
or U1643 (N_1643,N_1535,N_1557);
nand U1644 (N_1644,N_1573,N_1522);
and U1645 (N_1645,N_1562,N_1552);
nor U1646 (N_1646,N_1541,N_1572);
and U1647 (N_1647,N_1530,N_1568);
nor U1648 (N_1648,N_1544,N_1520);
and U1649 (N_1649,N_1548,N_1538);
nand U1650 (N_1650,N_1590,N_1625);
nand U1651 (N_1651,N_1613,N_1614);
nand U1652 (N_1652,N_1637,N_1638);
and U1653 (N_1653,N_1575,N_1623);
nand U1654 (N_1654,N_1648,N_1577);
or U1655 (N_1655,N_1597,N_1644);
nand U1656 (N_1656,N_1634,N_1585);
nand U1657 (N_1657,N_1620,N_1626);
nand U1658 (N_1658,N_1583,N_1604);
nand U1659 (N_1659,N_1611,N_1600);
and U1660 (N_1660,N_1593,N_1606);
nand U1661 (N_1661,N_1586,N_1615);
nand U1662 (N_1662,N_1612,N_1622);
or U1663 (N_1663,N_1595,N_1581);
or U1664 (N_1664,N_1587,N_1643);
and U1665 (N_1665,N_1588,N_1602);
or U1666 (N_1666,N_1639,N_1618);
and U1667 (N_1667,N_1645,N_1582);
and U1668 (N_1668,N_1589,N_1632);
nor U1669 (N_1669,N_1627,N_1619);
or U1670 (N_1670,N_1605,N_1621);
nand U1671 (N_1671,N_1579,N_1630);
or U1672 (N_1672,N_1598,N_1649);
nand U1673 (N_1673,N_1601,N_1610);
or U1674 (N_1674,N_1631,N_1647);
nor U1675 (N_1675,N_1576,N_1642);
or U1676 (N_1676,N_1635,N_1592);
or U1677 (N_1677,N_1584,N_1608);
nor U1678 (N_1678,N_1640,N_1628);
nand U1679 (N_1679,N_1591,N_1629);
xnor U1680 (N_1680,N_1646,N_1594);
nor U1681 (N_1681,N_1636,N_1603);
and U1682 (N_1682,N_1633,N_1616);
or U1683 (N_1683,N_1607,N_1596);
and U1684 (N_1684,N_1609,N_1580);
and U1685 (N_1685,N_1641,N_1617);
nand U1686 (N_1686,N_1624,N_1578);
nor U1687 (N_1687,N_1599,N_1618);
and U1688 (N_1688,N_1622,N_1627);
nand U1689 (N_1689,N_1586,N_1640);
nor U1690 (N_1690,N_1579,N_1605);
nor U1691 (N_1691,N_1609,N_1592);
nand U1692 (N_1692,N_1593,N_1600);
or U1693 (N_1693,N_1638,N_1640);
or U1694 (N_1694,N_1605,N_1580);
xnor U1695 (N_1695,N_1619,N_1644);
or U1696 (N_1696,N_1586,N_1631);
and U1697 (N_1697,N_1623,N_1597);
nor U1698 (N_1698,N_1646,N_1609);
or U1699 (N_1699,N_1631,N_1620);
or U1700 (N_1700,N_1628,N_1587);
and U1701 (N_1701,N_1635,N_1576);
xor U1702 (N_1702,N_1632,N_1622);
nor U1703 (N_1703,N_1609,N_1611);
nor U1704 (N_1704,N_1647,N_1615);
nand U1705 (N_1705,N_1627,N_1584);
or U1706 (N_1706,N_1622,N_1587);
nor U1707 (N_1707,N_1623,N_1579);
and U1708 (N_1708,N_1633,N_1580);
nor U1709 (N_1709,N_1610,N_1646);
or U1710 (N_1710,N_1618,N_1582);
nor U1711 (N_1711,N_1582,N_1634);
or U1712 (N_1712,N_1583,N_1627);
or U1713 (N_1713,N_1600,N_1642);
or U1714 (N_1714,N_1604,N_1646);
and U1715 (N_1715,N_1592,N_1576);
and U1716 (N_1716,N_1581,N_1643);
and U1717 (N_1717,N_1581,N_1632);
and U1718 (N_1718,N_1612,N_1636);
nand U1719 (N_1719,N_1629,N_1623);
and U1720 (N_1720,N_1593,N_1641);
nor U1721 (N_1721,N_1631,N_1628);
nand U1722 (N_1722,N_1582,N_1621);
nor U1723 (N_1723,N_1579,N_1595);
nand U1724 (N_1724,N_1642,N_1635);
and U1725 (N_1725,N_1682,N_1661);
nand U1726 (N_1726,N_1698,N_1702);
nand U1727 (N_1727,N_1674,N_1724);
and U1728 (N_1728,N_1656,N_1669);
and U1729 (N_1729,N_1719,N_1650);
or U1730 (N_1730,N_1670,N_1672);
and U1731 (N_1731,N_1680,N_1685);
nand U1732 (N_1732,N_1666,N_1710);
or U1733 (N_1733,N_1658,N_1665);
nand U1734 (N_1734,N_1668,N_1691);
nand U1735 (N_1735,N_1690,N_1700);
nand U1736 (N_1736,N_1652,N_1718);
and U1737 (N_1737,N_1696,N_1717);
and U1738 (N_1738,N_1660,N_1716);
nand U1739 (N_1739,N_1655,N_1706);
and U1740 (N_1740,N_1707,N_1720);
nand U1741 (N_1741,N_1677,N_1703);
nor U1742 (N_1742,N_1697,N_1688);
nor U1743 (N_1743,N_1711,N_1701);
xor U1744 (N_1744,N_1705,N_1659);
nor U1745 (N_1745,N_1671,N_1714);
and U1746 (N_1746,N_1675,N_1676);
and U1747 (N_1747,N_1662,N_1713);
or U1748 (N_1748,N_1723,N_1699);
nor U1749 (N_1749,N_1715,N_1692);
or U1750 (N_1750,N_1651,N_1653);
or U1751 (N_1751,N_1709,N_1722);
and U1752 (N_1752,N_1693,N_1654);
xnor U1753 (N_1753,N_1678,N_1679);
nand U1754 (N_1754,N_1681,N_1687);
nand U1755 (N_1755,N_1712,N_1683);
or U1756 (N_1756,N_1721,N_1664);
or U1757 (N_1757,N_1704,N_1694);
and U1758 (N_1758,N_1657,N_1708);
or U1759 (N_1759,N_1695,N_1667);
and U1760 (N_1760,N_1673,N_1684);
nand U1761 (N_1761,N_1663,N_1686);
and U1762 (N_1762,N_1689,N_1712);
or U1763 (N_1763,N_1718,N_1669);
xor U1764 (N_1764,N_1666,N_1711);
and U1765 (N_1765,N_1693,N_1711);
nor U1766 (N_1766,N_1697,N_1718);
and U1767 (N_1767,N_1673,N_1686);
or U1768 (N_1768,N_1697,N_1676);
nand U1769 (N_1769,N_1674,N_1675);
nand U1770 (N_1770,N_1673,N_1669);
nand U1771 (N_1771,N_1654,N_1679);
nand U1772 (N_1772,N_1694,N_1706);
or U1773 (N_1773,N_1664,N_1703);
nor U1774 (N_1774,N_1695,N_1687);
and U1775 (N_1775,N_1686,N_1709);
nand U1776 (N_1776,N_1661,N_1658);
or U1777 (N_1777,N_1668,N_1664);
nor U1778 (N_1778,N_1685,N_1675);
and U1779 (N_1779,N_1679,N_1677);
and U1780 (N_1780,N_1670,N_1714);
and U1781 (N_1781,N_1683,N_1694);
and U1782 (N_1782,N_1667,N_1693);
and U1783 (N_1783,N_1664,N_1679);
nand U1784 (N_1784,N_1699,N_1696);
and U1785 (N_1785,N_1695,N_1679);
and U1786 (N_1786,N_1657,N_1707);
and U1787 (N_1787,N_1707,N_1710);
nor U1788 (N_1788,N_1656,N_1666);
nand U1789 (N_1789,N_1687,N_1659);
or U1790 (N_1790,N_1665,N_1708);
or U1791 (N_1791,N_1693,N_1690);
or U1792 (N_1792,N_1710,N_1679);
and U1793 (N_1793,N_1652,N_1693);
nor U1794 (N_1794,N_1662,N_1692);
and U1795 (N_1795,N_1689,N_1723);
nand U1796 (N_1796,N_1670,N_1689);
nand U1797 (N_1797,N_1679,N_1704);
nor U1798 (N_1798,N_1676,N_1715);
nor U1799 (N_1799,N_1664,N_1672);
nand U1800 (N_1800,N_1759,N_1749);
nand U1801 (N_1801,N_1773,N_1738);
nand U1802 (N_1802,N_1797,N_1792);
nor U1803 (N_1803,N_1727,N_1763);
nand U1804 (N_1804,N_1740,N_1754);
and U1805 (N_1805,N_1772,N_1739);
xnor U1806 (N_1806,N_1781,N_1768);
nor U1807 (N_1807,N_1752,N_1761);
or U1808 (N_1808,N_1753,N_1765);
nor U1809 (N_1809,N_1737,N_1793);
xor U1810 (N_1810,N_1757,N_1775);
nor U1811 (N_1811,N_1780,N_1748);
or U1812 (N_1812,N_1743,N_1750);
nor U1813 (N_1813,N_1788,N_1760);
or U1814 (N_1814,N_1769,N_1730);
or U1815 (N_1815,N_1787,N_1796);
nor U1816 (N_1816,N_1756,N_1770);
or U1817 (N_1817,N_1747,N_1762);
nor U1818 (N_1818,N_1771,N_1786);
and U1819 (N_1819,N_1778,N_1767);
and U1820 (N_1820,N_1776,N_1736);
and U1821 (N_1821,N_1791,N_1744);
and U1822 (N_1822,N_1766,N_1790);
nor U1823 (N_1823,N_1774,N_1732);
xor U1824 (N_1824,N_1777,N_1799);
or U1825 (N_1825,N_1783,N_1726);
nand U1826 (N_1826,N_1729,N_1784);
nor U1827 (N_1827,N_1728,N_1734);
xnor U1828 (N_1828,N_1758,N_1751);
nor U1829 (N_1829,N_1794,N_1795);
and U1830 (N_1830,N_1782,N_1735);
nand U1831 (N_1831,N_1733,N_1746);
or U1832 (N_1832,N_1742,N_1725);
and U1833 (N_1833,N_1745,N_1741);
and U1834 (N_1834,N_1764,N_1785);
and U1835 (N_1835,N_1755,N_1789);
and U1836 (N_1836,N_1798,N_1779);
or U1837 (N_1837,N_1731,N_1727);
nor U1838 (N_1838,N_1775,N_1755);
nor U1839 (N_1839,N_1791,N_1798);
nor U1840 (N_1840,N_1764,N_1787);
or U1841 (N_1841,N_1795,N_1765);
or U1842 (N_1842,N_1727,N_1768);
and U1843 (N_1843,N_1766,N_1767);
and U1844 (N_1844,N_1781,N_1785);
and U1845 (N_1845,N_1725,N_1797);
or U1846 (N_1846,N_1732,N_1725);
or U1847 (N_1847,N_1725,N_1756);
nor U1848 (N_1848,N_1778,N_1745);
or U1849 (N_1849,N_1772,N_1731);
nand U1850 (N_1850,N_1730,N_1768);
nand U1851 (N_1851,N_1762,N_1736);
and U1852 (N_1852,N_1756,N_1729);
nor U1853 (N_1853,N_1789,N_1774);
xor U1854 (N_1854,N_1799,N_1773);
nor U1855 (N_1855,N_1779,N_1731);
or U1856 (N_1856,N_1779,N_1787);
or U1857 (N_1857,N_1777,N_1758);
nor U1858 (N_1858,N_1781,N_1749);
or U1859 (N_1859,N_1740,N_1728);
nor U1860 (N_1860,N_1741,N_1764);
and U1861 (N_1861,N_1789,N_1785);
and U1862 (N_1862,N_1728,N_1762);
nand U1863 (N_1863,N_1740,N_1791);
and U1864 (N_1864,N_1753,N_1776);
nor U1865 (N_1865,N_1777,N_1769);
nand U1866 (N_1866,N_1733,N_1792);
nand U1867 (N_1867,N_1765,N_1793);
nor U1868 (N_1868,N_1773,N_1781);
nand U1869 (N_1869,N_1794,N_1799);
nand U1870 (N_1870,N_1741,N_1756);
and U1871 (N_1871,N_1776,N_1790);
or U1872 (N_1872,N_1737,N_1738);
nor U1873 (N_1873,N_1733,N_1782);
nor U1874 (N_1874,N_1735,N_1758);
and U1875 (N_1875,N_1819,N_1809);
and U1876 (N_1876,N_1833,N_1806);
and U1877 (N_1877,N_1822,N_1869);
or U1878 (N_1878,N_1864,N_1850);
nor U1879 (N_1879,N_1871,N_1847);
and U1880 (N_1880,N_1835,N_1813);
or U1881 (N_1881,N_1844,N_1839);
nor U1882 (N_1882,N_1865,N_1862);
nand U1883 (N_1883,N_1816,N_1827);
or U1884 (N_1884,N_1866,N_1863);
nand U1885 (N_1885,N_1825,N_1817);
nor U1886 (N_1886,N_1802,N_1846);
nor U1887 (N_1887,N_1841,N_1826);
nand U1888 (N_1888,N_1855,N_1872);
and U1889 (N_1889,N_1868,N_1859);
or U1890 (N_1890,N_1848,N_1845);
nand U1891 (N_1891,N_1838,N_1830);
and U1892 (N_1892,N_1832,N_1852);
nor U1893 (N_1893,N_1870,N_1812);
and U1894 (N_1894,N_1861,N_1840);
nand U1895 (N_1895,N_1849,N_1814);
or U1896 (N_1896,N_1823,N_1867);
nand U1897 (N_1897,N_1842,N_1834);
nand U1898 (N_1898,N_1800,N_1856);
or U1899 (N_1899,N_1805,N_1810);
or U1900 (N_1900,N_1873,N_1836);
nand U1901 (N_1901,N_1828,N_1815);
nand U1902 (N_1902,N_1874,N_1851);
xnor U1903 (N_1903,N_1811,N_1854);
or U1904 (N_1904,N_1804,N_1831);
or U1905 (N_1905,N_1818,N_1837);
nand U1906 (N_1906,N_1829,N_1801);
nor U1907 (N_1907,N_1843,N_1821);
and U1908 (N_1908,N_1857,N_1860);
and U1909 (N_1909,N_1820,N_1803);
nand U1910 (N_1910,N_1807,N_1824);
nor U1911 (N_1911,N_1858,N_1808);
or U1912 (N_1912,N_1853,N_1822);
nand U1913 (N_1913,N_1815,N_1858);
and U1914 (N_1914,N_1838,N_1855);
or U1915 (N_1915,N_1866,N_1816);
or U1916 (N_1916,N_1812,N_1845);
nand U1917 (N_1917,N_1812,N_1831);
or U1918 (N_1918,N_1831,N_1823);
or U1919 (N_1919,N_1803,N_1872);
nor U1920 (N_1920,N_1864,N_1874);
or U1921 (N_1921,N_1834,N_1830);
xnor U1922 (N_1922,N_1832,N_1806);
and U1923 (N_1923,N_1815,N_1840);
nor U1924 (N_1924,N_1860,N_1830);
nand U1925 (N_1925,N_1863,N_1804);
nand U1926 (N_1926,N_1835,N_1812);
nor U1927 (N_1927,N_1834,N_1852);
or U1928 (N_1928,N_1864,N_1839);
and U1929 (N_1929,N_1827,N_1870);
nor U1930 (N_1930,N_1869,N_1861);
nand U1931 (N_1931,N_1840,N_1864);
and U1932 (N_1932,N_1805,N_1830);
nand U1933 (N_1933,N_1820,N_1869);
nor U1934 (N_1934,N_1819,N_1837);
nor U1935 (N_1935,N_1843,N_1849);
and U1936 (N_1936,N_1824,N_1872);
and U1937 (N_1937,N_1819,N_1803);
nand U1938 (N_1938,N_1814,N_1865);
nand U1939 (N_1939,N_1818,N_1860);
or U1940 (N_1940,N_1841,N_1800);
nor U1941 (N_1941,N_1834,N_1846);
and U1942 (N_1942,N_1837,N_1850);
nor U1943 (N_1943,N_1836,N_1809);
or U1944 (N_1944,N_1868,N_1843);
and U1945 (N_1945,N_1850,N_1819);
nor U1946 (N_1946,N_1818,N_1868);
nor U1947 (N_1947,N_1807,N_1820);
and U1948 (N_1948,N_1825,N_1849);
and U1949 (N_1949,N_1846,N_1870);
xnor U1950 (N_1950,N_1916,N_1939);
nand U1951 (N_1951,N_1910,N_1890);
and U1952 (N_1952,N_1921,N_1946);
xor U1953 (N_1953,N_1928,N_1906);
xor U1954 (N_1954,N_1933,N_1913);
nand U1955 (N_1955,N_1927,N_1878);
and U1956 (N_1956,N_1932,N_1908);
or U1957 (N_1957,N_1889,N_1886);
nand U1958 (N_1958,N_1875,N_1912);
nor U1959 (N_1959,N_1943,N_1899);
nand U1960 (N_1960,N_1876,N_1941);
or U1961 (N_1961,N_1909,N_1877);
and U1962 (N_1962,N_1905,N_1942);
nor U1963 (N_1963,N_1919,N_1888);
or U1964 (N_1964,N_1922,N_1938);
or U1965 (N_1965,N_1882,N_1923);
and U1966 (N_1966,N_1948,N_1936);
nor U1967 (N_1967,N_1937,N_1885);
nand U1968 (N_1968,N_1915,N_1902);
and U1969 (N_1969,N_1935,N_1891);
nand U1970 (N_1970,N_1920,N_1893);
or U1971 (N_1971,N_1907,N_1879);
or U1972 (N_1972,N_1934,N_1925);
or U1973 (N_1973,N_1901,N_1924);
or U1974 (N_1974,N_1929,N_1926);
nand U1975 (N_1975,N_1947,N_1900);
or U1976 (N_1976,N_1898,N_1945);
and U1977 (N_1977,N_1903,N_1892);
and U1978 (N_1978,N_1884,N_1880);
nor U1979 (N_1979,N_1940,N_1914);
nand U1980 (N_1980,N_1881,N_1949);
nand U1981 (N_1981,N_1931,N_1897);
or U1982 (N_1982,N_1894,N_1917);
and U1983 (N_1983,N_1918,N_1930);
or U1984 (N_1984,N_1895,N_1896);
nand U1985 (N_1985,N_1883,N_1944);
and U1986 (N_1986,N_1904,N_1887);
nand U1987 (N_1987,N_1911,N_1888);
nor U1988 (N_1988,N_1901,N_1936);
and U1989 (N_1989,N_1898,N_1919);
or U1990 (N_1990,N_1917,N_1934);
nor U1991 (N_1991,N_1925,N_1897);
and U1992 (N_1992,N_1938,N_1894);
or U1993 (N_1993,N_1936,N_1909);
nand U1994 (N_1994,N_1935,N_1881);
and U1995 (N_1995,N_1889,N_1913);
nor U1996 (N_1996,N_1910,N_1918);
and U1997 (N_1997,N_1899,N_1885);
or U1998 (N_1998,N_1918,N_1936);
or U1999 (N_1999,N_1901,N_1933);
or U2000 (N_2000,N_1896,N_1947);
nand U2001 (N_2001,N_1884,N_1913);
nor U2002 (N_2002,N_1900,N_1877);
and U2003 (N_2003,N_1915,N_1935);
and U2004 (N_2004,N_1893,N_1911);
nor U2005 (N_2005,N_1934,N_1901);
nand U2006 (N_2006,N_1927,N_1924);
nor U2007 (N_2007,N_1923,N_1890);
or U2008 (N_2008,N_1883,N_1905);
nor U2009 (N_2009,N_1884,N_1888);
and U2010 (N_2010,N_1939,N_1898);
and U2011 (N_2011,N_1875,N_1898);
nand U2012 (N_2012,N_1923,N_1901);
and U2013 (N_2013,N_1882,N_1878);
nand U2014 (N_2014,N_1891,N_1909);
nand U2015 (N_2015,N_1945,N_1912);
nor U2016 (N_2016,N_1929,N_1928);
nand U2017 (N_2017,N_1921,N_1896);
and U2018 (N_2018,N_1937,N_1932);
and U2019 (N_2019,N_1898,N_1889);
or U2020 (N_2020,N_1915,N_1908);
or U2021 (N_2021,N_1883,N_1932);
and U2022 (N_2022,N_1937,N_1912);
nand U2023 (N_2023,N_1924,N_1896);
or U2024 (N_2024,N_1885,N_1916);
or U2025 (N_2025,N_2008,N_2023);
or U2026 (N_2026,N_1997,N_1955);
nor U2027 (N_2027,N_1967,N_1951);
nand U2028 (N_2028,N_1988,N_2002);
or U2029 (N_2029,N_1972,N_2001);
nand U2030 (N_2030,N_1960,N_2012);
or U2031 (N_2031,N_1992,N_1999);
nor U2032 (N_2032,N_1975,N_2006);
or U2033 (N_2033,N_1989,N_1981);
nor U2034 (N_2034,N_1983,N_1966);
or U2035 (N_2035,N_1979,N_2000);
nor U2036 (N_2036,N_2013,N_2022);
and U2037 (N_2037,N_1973,N_1970);
or U2038 (N_2038,N_2024,N_1956);
nand U2039 (N_2039,N_1968,N_2010);
nor U2040 (N_2040,N_1986,N_2005);
and U2041 (N_2041,N_1991,N_2019);
nand U2042 (N_2042,N_2009,N_2018);
nand U2043 (N_2043,N_1971,N_1953);
nand U2044 (N_2044,N_1987,N_2014);
and U2045 (N_2045,N_1978,N_1985);
or U2046 (N_2046,N_1982,N_1993);
or U2047 (N_2047,N_1994,N_2003);
or U2048 (N_2048,N_1974,N_1952);
nor U2049 (N_2049,N_2007,N_1995);
and U2050 (N_2050,N_2004,N_2011);
nand U2051 (N_2051,N_2017,N_2020);
and U2052 (N_2052,N_1963,N_2021);
nor U2053 (N_2053,N_1984,N_1977);
nand U2054 (N_2054,N_1990,N_2015);
or U2055 (N_2055,N_1959,N_1964);
nor U2056 (N_2056,N_1961,N_1962);
nor U2057 (N_2057,N_1980,N_1957);
nor U2058 (N_2058,N_1958,N_2016);
or U2059 (N_2059,N_1969,N_1954);
or U2060 (N_2060,N_1965,N_1976);
nor U2061 (N_2061,N_1998,N_1996);
or U2062 (N_2062,N_1950,N_2018);
nor U2063 (N_2063,N_1950,N_1951);
or U2064 (N_2064,N_1983,N_1995);
and U2065 (N_2065,N_1996,N_2018);
and U2066 (N_2066,N_2016,N_2020);
nand U2067 (N_2067,N_1974,N_1979);
nor U2068 (N_2068,N_2011,N_2001);
nor U2069 (N_2069,N_2016,N_1955);
or U2070 (N_2070,N_2002,N_1973);
or U2071 (N_2071,N_1992,N_1960);
nand U2072 (N_2072,N_1968,N_1997);
or U2073 (N_2073,N_1967,N_2014);
nand U2074 (N_2074,N_1984,N_1950);
or U2075 (N_2075,N_1978,N_1992);
nand U2076 (N_2076,N_1966,N_1972);
nand U2077 (N_2077,N_1990,N_1951);
nor U2078 (N_2078,N_1951,N_1999);
nand U2079 (N_2079,N_2011,N_1976);
nand U2080 (N_2080,N_1974,N_2023);
nor U2081 (N_2081,N_2000,N_2007);
nor U2082 (N_2082,N_1995,N_1981);
and U2083 (N_2083,N_2002,N_1990);
or U2084 (N_2084,N_1989,N_2003);
or U2085 (N_2085,N_1971,N_1986);
or U2086 (N_2086,N_1973,N_1955);
nor U2087 (N_2087,N_2012,N_2022);
nand U2088 (N_2088,N_1997,N_1984);
nand U2089 (N_2089,N_1961,N_1982);
and U2090 (N_2090,N_1965,N_2000);
or U2091 (N_2091,N_1976,N_1995);
nor U2092 (N_2092,N_1992,N_1981);
nand U2093 (N_2093,N_1950,N_1995);
nand U2094 (N_2094,N_1959,N_1991);
or U2095 (N_2095,N_1957,N_1983);
and U2096 (N_2096,N_1963,N_1989);
nand U2097 (N_2097,N_2017,N_1965);
and U2098 (N_2098,N_1998,N_1977);
and U2099 (N_2099,N_1968,N_1969);
or U2100 (N_2100,N_2093,N_2045);
or U2101 (N_2101,N_2099,N_2031);
xor U2102 (N_2102,N_2048,N_2087);
xor U2103 (N_2103,N_2049,N_2090);
and U2104 (N_2104,N_2091,N_2041);
nor U2105 (N_2105,N_2034,N_2080);
and U2106 (N_2106,N_2066,N_2078);
nand U2107 (N_2107,N_2053,N_2089);
and U2108 (N_2108,N_2088,N_2030);
and U2109 (N_2109,N_2073,N_2070);
nor U2110 (N_2110,N_2067,N_2092);
nor U2111 (N_2111,N_2046,N_2064);
and U2112 (N_2112,N_2036,N_2029);
or U2113 (N_2113,N_2038,N_2052);
nor U2114 (N_2114,N_2047,N_2068);
and U2115 (N_2115,N_2082,N_2026);
or U2116 (N_2116,N_2097,N_2061);
nand U2117 (N_2117,N_2081,N_2060);
nor U2118 (N_2118,N_2079,N_2063);
or U2119 (N_2119,N_2039,N_2065);
nor U2120 (N_2120,N_2056,N_2083);
and U2121 (N_2121,N_2040,N_2084);
nor U2122 (N_2122,N_2096,N_2069);
and U2123 (N_2123,N_2033,N_2077);
or U2124 (N_2124,N_2044,N_2072);
and U2125 (N_2125,N_2085,N_2025);
and U2126 (N_2126,N_2054,N_2055);
nor U2127 (N_2127,N_2076,N_2050);
and U2128 (N_2128,N_2059,N_2094);
and U2129 (N_2129,N_2037,N_2075);
and U2130 (N_2130,N_2095,N_2032);
or U2131 (N_2131,N_2098,N_2028);
or U2132 (N_2132,N_2058,N_2043);
and U2133 (N_2133,N_2086,N_2042);
nand U2134 (N_2134,N_2027,N_2051);
nor U2135 (N_2135,N_2035,N_2074);
and U2136 (N_2136,N_2071,N_2057);
nor U2137 (N_2137,N_2062,N_2084);
nand U2138 (N_2138,N_2060,N_2048);
nor U2139 (N_2139,N_2071,N_2065);
nor U2140 (N_2140,N_2057,N_2042);
or U2141 (N_2141,N_2060,N_2046);
nor U2142 (N_2142,N_2089,N_2099);
nand U2143 (N_2143,N_2084,N_2027);
nor U2144 (N_2144,N_2094,N_2046);
or U2145 (N_2145,N_2053,N_2092);
and U2146 (N_2146,N_2034,N_2026);
nand U2147 (N_2147,N_2087,N_2040);
or U2148 (N_2148,N_2091,N_2089);
and U2149 (N_2149,N_2029,N_2072);
and U2150 (N_2150,N_2073,N_2067);
nor U2151 (N_2151,N_2076,N_2090);
nor U2152 (N_2152,N_2050,N_2040);
nor U2153 (N_2153,N_2082,N_2070);
nor U2154 (N_2154,N_2082,N_2058);
and U2155 (N_2155,N_2091,N_2099);
nor U2156 (N_2156,N_2037,N_2034);
nor U2157 (N_2157,N_2093,N_2050);
nand U2158 (N_2158,N_2066,N_2051);
or U2159 (N_2159,N_2076,N_2064);
nor U2160 (N_2160,N_2051,N_2067);
and U2161 (N_2161,N_2050,N_2031);
nor U2162 (N_2162,N_2038,N_2064);
nand U2163 (N_2163,N_2071,N_2053);
or U2164 (N_2164,N_2039,N_2026);
and U2165 (N_2165,N_2070,N_2053);
nor U2166 (N_2166,N_2036,N_2057);
or U2167 (N_2167,N_2029,N_2099);
or U2168 (N_2168,N_2035,N_2091);
nor U2169 (N_2169,N_2034,N_2072);
xor U2170 (N_2170,N_2061,N_2082);
nor U2171 (N_2171,N_2048,N_2042);
and U2172 (N_2172,N_2081,N_2026);
or U2173 (N_2173,N_2078,N_2059);
nor U2174 (N_2174,N_2099,N_2094);
xor U2175 (N_2175,N_2111,N_2105);
and U2176 (N_2176,N_2108,N_2119);
or U2177 (N_2177,N_2121,N_2142);
or U2178 (N_2178,N_2165,N_2153);
nand U2179 (N_2179,N_2169,N_2173);
nor U2180 (N_2180,N_2161,N_2174);
xor U2181 (N_2181,N_2124,N_2113);
or U2182 (N_2182,N_2141,N_2138);
nand U2183 (N_2183,N_2150,N_2156);
nor U2184 (N_2184,N_2149,N_2168);
or U2185 (N_2185,N_2160,N_2152);
and U2186 (N_2186,N_2145,N_2131);
xnor U2187 (N_2187,N_2107,N_2157);
or U2188 (N_2188,N_2159,N_2170);
nor U2189 (N_2189,N_2106,N_2135);
nand U2190 (N_2190,N_2118,N_2102);
nor U2191 (N_2191,N_2146,N_2101);
and U2192 (N_2192,N_2116,N_2123);
and U2193 (N_2193,N_2122,N_2163);
nor U2194 (N_2194,N_2147,N_2130);
or U2195 (N_2195,N_2104,N_2172);
or U2196 (N_2196,N_2166,N_2154);
or U2197 (N_2197,N_2109,N_2120);
nor U2198 (N_2198,N_2139,N_2144);
nor U2199 (N_2199,N_2127,N_2148);
nand U2200 (N_2200,N_2115,N_2136);
and U2201 (N_2201,N_2167,N_2140);
and U2202 (N_2202,N_2112,N_2110);
or U2203 (N_2203,N_2129,N_2133);
nand U2204 (N_2204,N_2143,N_2100);
nor U2205 (N_2205,N_2103,N_2126);
and U2206 (N_2206,N_2125,N_2137);
nor U2207 (N_2207,N_2117,N_2164);
nor U2208 (N_2208,N_2134,N_2171);
nand U2209 (N_2209,N_2162,N_2151);
and U2210 (N_2210,N_2114,N_2132);
or U2211 (N_2211,N_2158,N_2128);
and U2212 (N_2212,N_2155,N_2120);
and U2213 (N_2213,N_2161,N_2116);
nor U2214 (N_2214,N_2135,N_2137);
nand U2215 (N_2215,N_2132,N_2121);
nor U2216 (N_2216,N_2137,N_2112);
and U2217 (N_2217,N_2163,N_2112);
nand U2218 (N_2218,N_2132,N_2128);
nand U2219 (N_2219,N_2108,N_2163);
and U2220 (N_2220,N_2120,N_2104);
nor U2221 (N_2221,N_2146,N_2100);
nand U2222 (N_2222,N_2124,N_2150);
nor U2223 (N_2223,N_2137,N_2168);
nor U2224 (N_2224,N_2126,N_2108);
and U2225 (N_2225,N_2149,N_2133);
and U2226 (N_2226,N_2103,N_2127);
nor U2227 (N_2227,N_2153,N_2129);
nor U2228 (N_2228,N_2116,N_2169);
and U2229 (N_2229,N_2141,N_2102);
and U2230 (N_2230,N_2140,N_2130);
or U2231 (N_2231,N_2101,N_2134);
or U2232 (N_2232,N_2108,N_2153);
nor U2233 (N_2233,N_2117,N_2120);
and U2234 (N_2234,N_2151,N_2113);
or U2235 (N_2235,N_2112,N_2173);
nor U2236 (N_2236,N_2107,N_2126);
or U2237 (N_2237,N_2123,N_2105);
xor U2238 (N_2238,N_2168,N_2140);
or U2239 (N_2239,N_2131,N_2168);
nor U2240 (N_2240,N_2115,N_2167);
nand U2241 (N_2241,N_2145,N_2170);
and U2242 (N_2242,N_2167,N_2160);
and U2243 (N_2243,N_2119,N_2167);
or U2244 (N_2244,N_2141,N_2157);
or U2245 (N_2245,N_2118,N_2148);
xor U2246 (N_2246,N_2146,N_2135);
or U2247 (N_2247,N_2152,N_2150);
nand U2248 (N_2248,N_2139,N_2134);
nor U2249 (N_2249,N_2105,N_2127);
or U2250 (N_2250,N_2178,N_2238);
and U2251 (N_2251,N_2244,N_2197);
nand U2252 (N_2252,N_2211,N_2232);
nand U2253 (N_2253,N_2214,N_2210);
and U2254 (N_2254,N_2202,N_2239);
or U2255 (N_2255,N_2184,N_2209);
xnor U2256 (N_2256,N_2228,N_2205);
or U2257 (N_2257,N_2246,N_2237);
nand U2258 (N_2258,N_2188,N_2181);
nor U2259 (N_2259,N_2221,N_2216);
or U2260 (N_2260,N_2229,N_2193);
nor U2261 (N_2261,N_2231,N_2186);
or U2262 (N_2262,N_2218,N_2190);
and U2263 (N_2263,N_2176,N_2199);
or U2264 (N_2264,N_2224,N_2243);
nand U2265 (N_2265,N_2213,N_2207);
or U2266 (N_2266,N_2227,N_2212);
and U2267 (N_2267,N_2182,N_2194);
or U2268 (N_2268,N_2247,N_2175);
nand U2269 (N_2269,N_2235,N_2234);
and U2270 (N_2270,N_2191,N_2185);
and U2271 (N_2271,N_2215,N_2198);
nand U2272 (N_2272,N_2230,N_2192);
and U2273 (N_2273,N_2249,N_2180);
or U2274 (N_2274,N_2240,N_2219);
or U2275 (N_2275,N_2241,N_2204);
nor U2276 (N_2276,N_2200,N_2242);
and U2277 (N_2277,N_2245,N_2206);
nand U2278 (N_2278,N_2183,N_2203);
nand U2279 (N_2279,N_2233,N_2177);
nor U2280 (N_2280,N_2226,N_2222);
nor U2281 (N_2281,N_2189,N_2195);
and U2282 (N_2282,N_2236,N_2201);
and U2283 (N_2283,N_2208,N_2217);
nand U2284 (N_2284,N_2220,N_2225);
and U2285 (N_2285,N_2187,N_2248);
nor U2286 (N_2286,N_2223,N_2179);
and U2287 (N_2287,N_2196,N_2191);
or U2288 (N_2288,N_2244,N_2181);
nand U2289 (N_2289,N_2234,N_2231);
and U2290 (N_2290,N_2234,N_2217);
or U2291 (N_2291,N_2245,N_2210);
nor U2292 (N_2292,N_2209,N_2203);
or U2293 (N_2293,N_2196,N_2247);
and U2294 (N_2294,N_2204,N_2187);
and U2295 (N_2295,N_2201,N_2227);
or U2296 (N_2296,N_2226,N_2175);
and U2297 (N_2297,N_2185,N_2214);
nand U2298 (N_2298,N_2242,N_2217);
or U2299 (N_2299,N_2222,N_2210);
nor U2300 (N_2300,N_2218,N_2191);
and U2301 (N_2301,N_2233,N_2212);
and U2302 (N_2302,N_2224,N_2223);
and U2303 (N_2303,N_2213,N_2219);
or U2304 (N_2304,N_2184,N_2238);
nor U2305 (N_2305,N_2248,N_2190);
nand U2306 (N_2306,N_2205,N_2187);
or U2307 (N_2307,N_2211,N_2204);
or U2308 (N_2308,N_2188,N_2193);
nand U2309 (N_2309,N_2216,N_2201);
and U2310 (N_2310,N_2229,N_2217);
and U2311 (N_2311,N_2216,N_2215);
nand U2312 (N_2312,N_2187,N_2242);
nand U2313 (N_2313,N_2247,N_2245);
or U2314 (N_2314,N_2245,N_2234);
or U2315 (N_2315,N_2249,N_2207);
nand U2316 (N_2316,N_2248,N_2225);
or U2317 (N_2317,N_2223,N_2209);
nand U2318 (N_2318,N_2197,N_2222);
nor U2319 (N_2319,N_2247,N_2227);
or U2320 (N_2320,N_2179,N_2185);
nor U2321 (N_2321,N_2228,N_2240);
and U2322 (N_2322,N_2246,N_2179);
and U2323 (N_2323,N_2186,N_2226);
nor U2324 (N_2324,N_2184,N_2221);
and U2325 (N_2325,N_2261,N_2252);
xnor U2326 (N_2326,N_2282,N_2257);
nor U2327 (N_2327,N_2253,N_2307);
or U2328 (N_2328,N_2317,N_2310);
and U2329 (N_2329,N_2308,N_2322);
or U2330 (N_2330,N_2303,N_2275);
and U2331 (N_2331,N_2289,N_2280);
or U2332 (N_2332,N_2288,N_2268);
and U2333 (N_2333,N_2254,N_2294);
nand U2334 (N_2334,N_2255,N_2301);
xor U2335 (N_2335,N_2296,N_2285);
and U2336 (N_2336,N_2274,N_2306);
or U2337 (N_2337,N_2319,N_2292);
nand U2338 (N_2338,N_2321,N_2324);
or U2339 (N_2339,N_2258,N_2315);
or U2340 (N_2340,N_2304,N_2286);
nor U2341 (N_2341,N_2312,N_2269);
nand U2342 (N_2342,N_2323,N_2314);
or U2343 (N_2343,N_2284,N_2276);
nand U2344 (N_2344,N_2271,N_2302);
and U2345 (N_2345,N_2299,N_2281);
nand U2346 (N_2346,N_2309,N_2278);
nand U2347 (N_2347,N_2318,N_2290);
and U2348 (N_2348,N_2297,N_2279);
and U2349 (N_2349,N_2300,N_2283);
and U2350 (N_2350,N_2259,N_2270);
nand U2351 (N_2351,N_2316,N_2272);
nand U2352 (N_2352,N_2262,N_2293);
or U2353 (N_2353,N_2320,N_2260);
nand U2354 (N_2354,N_2266,N_2305);
or U2355 (N_2355,N_2273,N_2263);
or U2356 (N_2356,N_2287,N_2267);
nor U2357 (N_2357,N_2250,N_2256);
xnor U2358 (N_2358,N_2311,N_2298);
nand U2359 (N_2359,N_2277,N_2291);
xnor U2360 (N_2360,N_2295,N_2251);
nand U2361 (N_2361,N_2265,N_2264);
or U2362 (N_2362,N_2313,N_2316);
and U2363 (N_2363,N_2289,N_2287);
nor U2364 (N_2364,N_2287,N_2297);
nand U2365 (N_2365,N_2253,N_2291);
and U2366 (N_2366,N_2273,N_2306);
and U2367 (N_2367,N_2276,N_2324);
nor U2368 (N_2368,N_2263,N_2257);
nand U2369 (N_2369,N_2271,N_2303);
nor U2370 (N_2370,N_2270,N_2296);
nor U2371 (N_2371,N_2250,N_2301);
and U2372 (N_2372,N_2287,N_2253);
and U2373 (N_2373,N_2274,N_2302);
and U2374 (N_2374,N_2260,N_2259);
nor U2375 (N_2375,N_2270,N_2303);
nor U2376 (N_2376,N_2295,N_2267);
nand U2377 (N_2377,N_2260,N_2251);
nor U2378 (N_2378,N_2323,N_2286);
and U2379 (N_2379,N_2267,N_2290);
or U2380 (N_2380,N_2323,N_2279);
nor U2381 (N_2381,N_2316,N_2271);
nand U2382 (N_2382,N_2265,N_2309);
nor U2383 (N_2383,N_2276,N_2278);
and U2384 (N_2384,N_2302,N_2268);
nor U2385 (N_2385,N_2318,N_2296);
and U2386 (N_2386,N_2312,N_2303);
nor U2387 (N_2387,N_2261,N_2309);
or U2388 (N_2388,N_2286,N_2315);
nor U2389 (N_2389,N_2256,N_2287);
nand U2390 (N_2390,N_2252,N_2297);
nand U2391 (N_2391,N_2317,N_2262);
xor U2392 (N_2392,N_2270,N_2318);
nor U2393 (N_2393,N_2270,N_2278);
nand U2394 (N_2394,N_2281,N_2289);
nand U2395 (N_2395,N_2311,N_2281);
nand U2396 (N_2396,N_2320,N_2274);
or U2397 (N_2397,N_2289,N_2272);
nor U2398 (N_2398,N_2276,N_2250);
or U2399 (N_2399,N_2279,N_2304);
nand U2400 (N_2400,N_2371,N_2376);
nand U2401 (N_2401,N_2330,N_2366);
nand U2402 (N_2402,N_2374,N_2395);
or U2403 (N_2403,N_2340,N_2389);
and U2404 (N_2404,N_2362,N_2399);
nor U2405 (N_2405,N_2360,N_2326);
and U2406 (N_2406,N_2367,N_2329);
nand U2407 (N_2407,N_2336,N_2357);
and U2408 (N_2408,N_2347,N_2358);
nor U2409 (N_2409,N_2349,N_2373);
or U2410 (N_2410,N_2333,N_2355);
nor U2411 (N_2411,N_2387,N_2351);
nand U2412 (N_2412,N_2375,N_2398);
xnor U2413 (N_2413,N_2334,N_2331);
nor U2414 (N_2414,N_2341,N_2332);
or U2415 (N_2415,N_2345,N_2350);
and U2416 (N_2416,N_2378,N_2352);
xor U2417 (N_2417,N_2386,N_2348);
nand U2418 (N_2418,N_2327,N_2377);
nand U2419 (N_2419,N_2382,N_2380);
nand U2420 (N_2420,N_2394,N_2392);
or U2421 (N_2421,N_2381,N_2354);
or U2422 (N_2422,N_2363,N_2343);
nand U2423 (N_2423,N_2328,N_2356);
nand U2424 (N_2424,N_2361,N_2342);
and U2425 (N_2425,N_2364,N_2379);
or U2426 (N_2426,N_2346,N_2393);
nor U2427 (N_2427,N_2397,N_2369);
nand U2428 (N_2428,N_2325,N_2391);
and U2429 (N_2429,N_2337,N_2388);
and U2430 (N_2430,N_2390,N_2359);
and U2431 (N_2431,N_2339,N_2368);
or U2432 (N_2432,N_2344,N_2353);
or U2433 (N_2433,N_2365,N_2396);
and U2434 (N_2434,N_2383,N_2335);
nor U2435 (N_2435,N_2384,N_2372);
or U2436 (N_2436,N_2338,N_2370);
nor U2437 (N_2437,N_2385,N_2376);
nor U2438 (N_2438,N_2335,N_2355);
and U2439 (N_2439,N_2349,N_2387);
or U2440 (N_2440,N_2342,N_2383);
nand U2441 (N_2441,N_2390,N_2367);
nor U2442 (N_2442,N_2372,N_2338);
nor U2443 (N_2443,N_2340,N_2385);
nand U2444 (N_2444,N_2370,N_2372);
nor U2445 (N_2445,N_2334,N_2381);
or U2446 (N_2446,N_2374,N_2353);
and U2447 (N_2447,N_2353,N_2387);
or U2448 (N_2448,N_2397,N_2390);
or U2449 (N_2449,N_2363,N_2382);
nor U2450 (N_2450,N_2350,N_2372);
nor U2451 (N_2451,N_2335,N_2389);
or U2452 (N_2452,N_2352,N_2337);
and U2453 (N_2453,N_2396,N_2374);
nor U2454 (N_2454,N_2330,N_2371);
nor U2455 (N_2455,N_2356,N_2368);
and U2456 (N_2456,N_2325,N_2351);
nand U2457 (N_2457,N_2359,N_2367);
nand U2458 (N_2458,N_2360,N_2389);
nand U2459 (N_2459,N_2360,N_2348);
nand U2460 (N_2460,N_2359,N_2396);
or U2461 (N_2461,N_2348,N_2345);
nor U2462 (N_2462,N_2363,N_2331);
and U2463 (N_2463,N_2330,N_2333);
nor U2464 (N_2464,N_2359,N_2380);
nor U2465 (N_2465,N_2352,N_2342);
nor U2466 (N_2466,N_2393,N_2366);
nor U2467 (N_2467,N_2331,N_2359);
and U2468 (N_2468,N_2348,N_2374);
nand U2469 (N_2469,N_2332,N_2349);
nor U2470 (N_2470,N_2351,N_2374);
nor U2471 (N_2471,N_2383,N_2378);
nor U2472 (N_2472,N_2360,N_2338);
or U2473 (N_2473,N_2361,N_2354);
nand U2474 (N_2474,N_2372,N_2352);
nor U2475 (N_2475,N_2461,N_2426);
or U2476 (N_2476,N_2468,N_2427);
nor U2477 (N_2477,N_2451,N_2438);
nand U2478 (N_2478,N_2439,N_2459);
nand U2479 (N_2479,N_2428,N_2454);
xnor U2480 (N_2480,N_2416,N_2402);
nand U2481 (N_2481,N_2448,N_2456);
or U2482 (N_2482,N_2462,N_2410);
nand U2483 (N_2483,N_2474,N_2409);
nand U2484 (N_2484,N_2430,N_2440);
nor U2485 (N_2485,N_2437,N_2404);
nand U2486 (N_2486,N_2465,N_2435);
nor U2487 (N_2487,N_2467,N_2469);
or U2488 (N_2488,N_2434,N_2403);
or U2489 (N_2489,N_2418,N_2466);
or U2490 (N_2490,N_2457,N_2460);
or U2491 (N_2491,N_2425,N_2422);
or U2492 (N_2492,N_2412,N_2453);
nand U2493 (N_2493,N_2446,N_2441);
nand U2494 (N_2494,N_2413,N_2444);
and U2495 (N_2495,N_2405,N_2442);
nand U2496 (N_2496,N_2447,N_2415);
nor U2497 (N_2497,N_2452,N_2429);
and U2498 (N_2498,N_2400,N_2420);
nor U2499 (N_2499,N_2406,N_2423);
and U2500 (N_2500,N_2421,N_2431);
or U2501 (N_2501,N_2414,N_2470);
nand U2502 (N_2502,N_2432,N_2408);
nor U2503 (N_2503,N_2417,N_2424);
and U2504 (N_2504,N_2450,N_2458);
or U2505 (N_2505,N_2411,N_2401);
and U2506 (N_2506,N_2463,N_2449);
nor U2507 (N_2507,N_2407,N_2419);
or U2508 (N_2508,N_2436,N_2445);
nand U2509 (N_2509,N_2473,N_2471);
and U2510 (N_2510,N_2472,N_2464);
nor U2511 (N_2511,N_2455,N_2443);
nand U2512 (N_2512,N_2433,N_2468);
or U2513 (N_2513,N_2421,N_2424);
nand U2514 (N_2514,N_2461,N_2471);
nor U2515 (N_2515,N_2431,N_2464);
nand U2516 (N_2516,N_2429,N_2405);
or U2517 (N_2517,N_2407,N_2429);
and U2518 (N_2518,N_2400,N_2431);
nand U2519 (N_2519,N_2416,N_2470);
nor U2520 (N_2520,N_2433,N_2473);
nor U2521 (N_2521,N_2438,N_2424);
or U2522 (N_2522,N_2429,N_2433);
nand U2523 (N_2523,N_2425,N_2418);
and U2524 (N_2524,N_2442,N_2435);
or U2525 (N_2525,N_2432,N_2422);
or U2526 (N_2526,N_2404,N_2454);
nand U2527 (N_2527,N_2425,N_2466);
nor U2528 (N_2528,N_2459,N_2438);
nor U2529 (N_2529,N_2424,N_2435);
nor U2530 (N_2530,N_2472,N_2400);
or U2531 (N_2531,N_2404,N_2411);
or U2532 (N_2532,N_2426,N_2405);
nand U2533 (N_2533,N_2443,N_2437);
nand U2534 (N_2534,N_2431,N_2419);
nor U2535 (N_2535,N_2419,N_2469);
and U2536 (N_2536,N_2471,N_2434);
nand U2537 (N_2537,N_2446,N_2427);
or U2538 (N_2538,N_2461,N_2442);
nor U2539 (N_2539,N_2457,N_2426);
or U2540 (N_2540,N_2430,N_2416);
nor U2541 (N_2541,N_2400,N_2449);
nand U2542 (N_2542,N_2461,N_2459);
nand U2543 (N_2543,N_2432,N_2429);
and U2544 (N_2544,N_2442,N_2423);
or U2545 (N_2545,N_2428,N_2471);
nand U2546 (N_2546,N_2422,N_2447);
and U2547 (N_2547,N_2458,N_2470);
and U2548 (N_2548,N_2460,N_2418);
nor U2549 (N_2549,N_2457,N_2449);
or U2550 (N_2550,N_2477,N_2505);
or U2551 (N_2551,N_2500,N_2518);
or U2552 (N_2552,N_2498,N_2487);
and U2553 (N_2553,N_2517,N_2479);
nor U2554 (N_2554,N_2501,N_2544);
nor U2555 (N_2555,N_2536,N_2481);
nand U2556 (N_2556,N_2491,N_2483);
and U2557 (N_2557,N_2548,N_2537);
nor U2558 (N_2558,N_2546,N_2516);
nor U2559 (N_2559,N_2475,N_2535);
or U2560 (N_2560,N_2485,N_2490);
or U2561 (N_2561,N_2496,N_2520);
and U2562 (N_2562,N_2542,N_2524);
nand U2563 (N_2563,N_2506,N_2476);
and U2564 (N_2564,N_2531,N_2545);
or U2565 (N_2565,N_2527,N_2549);
nor U2566 (N_2566,N_2521,N_2511);
nand U2567 (N_2567,N_2522,N_2528);
nand U2568 (N_2568,N_2519,N_2502);
nand U2569 (N_2569,N_2529,N_2507);
or U2570 (N_2570,N_2533,N_2499);
nor U2571 (N_2571,N_2486,N_2508);
nand U2572 (N_2572,N_2525,N_2492);
nand U2573 (N_2573,N_2489,N_2482);
or U2574 (N_2574,N_2540,N_2538);
nor U2575 (N_2575,N_2523,N_2493);
nor U2576 (N_2576,N_2478,N_2513);
and U2577 (N_2577,N_2484,N_2480);
or U2578 (N_2578,N_2509,N_2512);
or U2579 (N_2579,N_2532,N_2543);
or U2580 (N_2580,N_2497,N_2494);
and U2581 (N_2581,N_2515,N_2495);
or U2582 (N_2582,N_2514,N_2526);
nand U2583 (N_2583,N_2539,N_2488);
or U2584 (N_2584,N_2504,N_2534);
nand U2585 (N_2585,N_2541,N_2510);
and U2586 (N_2586,N_2503,N_2547);
and U2587 (N_2587,N_2530,N_2490);
nand U2588 (N_2588,N_2506,N_2539);
and U2589 (N_2589,N_2538,N_2516);
or U2590 (N_2590,N_2477,N_2488);
or U2591 (N_2591,N_2541,N_2506);
nand U2592 (N_2592,N_2483,N_2528);
and U2593 (N_2593,N_2524,N_2518);
or U2594 (N_2594,N_2512,N_2479);
or U2595 (N_2595,N_2532,N_2540);
or U2596 (N_2596,N_2538,N_2498);
and U2597 (N_2597,N_2482,N_2490);
or U2598 (N_2598,N_2479,N_2477);
or U2599 (N_2599,N_2535,N_2498);
or U2600 (N_2600,N_2526,N_2541);
or U2601 (N_2601,N_2514,N_2497);
nand U2602 (N_2602,N_2546,N_2534);
or U2603 (N_2603,N_2498,N_2533);
nor U2604 (N_2604,N_2530,N_2495);
nor U2605 (N_2605,N_2494,N_2488);
or U2606 (N_2606,N_2493,N_2541);
and U2607 (N_2607,N_2502,N_2534);
or U2608 (N_2608,N_2543,N_2516);
nor U2609 (N_2609,N_2549,N_2500);
nand U2610 (N_2610,N_2504,N_2543);
and U2611 (N_2611,N_2504,N_2523);
and U2612 (N_2612,N_2527,N_2532);
and U2613 (N_2613,N_2488,N_2495);
and U2614 (N_2614,N_2516,N_2544);
and U2615 (N_2615,N_2545,N_2530);
nor U2616 (N_2616,N_2485,N_2475);
nor U2617 (N_2617,N_2485,N_2497);
nor U2618 (N_2618,N_2521,N_2490);
nor U2619 (N_2619,N_2481,N_2516);
nor U2620 (N_2620,N_2506,N_2524);
xor U2621 (N_2621,N_2537,N_2517);
nor U2622 (N_2622,N_2479,N_2524);
and U2623 (N_2623,N_2484,N_2540);
or U2624 (N_2624,N_2528,N_2541);
nand U2625 (N_2625,N_2585,N_2618);
nor U2626 (N_2626,N_2610,N_2622);
and U2627 (N_2627,N_2567,N_2577);
and U2628 (N_2628,N_2602,N_2554);
nor U2629 (N_2629,N_2561,N_2596);
nor U2630 (N_2630,N_2582,N_2614);
and U2631 (N_2631,N_2593,N_2624);
nand U2632 (N_2632,N_2592,N_2575);
or U2633 (N_2633,N_2551,N_2599);
and U2634 (N_2634,N_2581,N_2583);
or U2635 (N_2635,N_2615,N_2595);
nand U2636 (N_2636,N_2556,N_2550);
nand U2637 (N_2637,N_2576,N_2584);
nor U2638 (N_2638,N_2617,N_2570);
nor U2639 (N_2639,N_2574,N_2563);
nor U2640 (N_2640,N_2589,N_2601);
xor U2641 (N_2641,N_2569,N_2564);
nor U2642 (N_2642,N_2560,N_2580);
nor U2643 (N_2643,N_2587,N_2557);
nand U2644 (N_2644,N_2571,N_2619);
nor U2645 (N_2645,N_2568,N_2604);
and U2646 (N_2646,N_2608,N_2590);
nor U2647 (N_2647,N_2597,N_2579);
and U2648 (N_2648,N_2600,N_2578);
nand U2649 (N_2649,N_2606,N_2552);
or U2650 (N_2650,N_2616,N_2573);
nand U2651 (N_2651,N_2605,N_2603);
or U2652 (N_2652,N_2559,N_2555);
nor U2653 (N_2653,N_2558,N_2553);
and U2654 (N_2654,N_2613,N_2566);
nand U2655 (N_2655,N_2565,N_2621);
nor U2656 (N_2656,N_2623,N_2598);
nor U2657 (N_2657,N_2620,N_2611);
nand U2658 (N_2658,N_2562,N_2609);
nor U2659 (N_2659,N_2612,N_2607);
nor U2660 (N_2660,N_2572,N_2586);
and U2661 (N_2661,N_2588,N_2594);
and U2662 (N_2662,N_2591,N_2587);
and U2663 (N_2663,N_2604,N_2563);
nor U2664 (N_2664,N_2610,N_2582);
nor U2665 (N_2665,N_2597,N_2619);
nand U2666 (N_2666,N_2611,N_2565);
and U2667 (N_2667,N_2550,N_2566);
nor U2668 (N_2668,N_2551,N_2556);
nor U2669 (N_2669,N_2604,N_2607);
nor U2670 (N_2670,N_2585,N_2582);
and U2671 (N_2671,N_2567,N_2580);
and U2672 (N_2672,N_2587,N_2624);
nand U2673 (N_2673,N_2596,N_2564);
and U2674 (N_2674,N_2559,N_2551);
nor U2675 (N_2675,N_2593,N_2586);
nand U2676 (N_2676,N_2583,N_2563);
nand U2677 (N_2677,N_2621,N_2579);
or U2678 (N_2678,N_2607,N_2611);
nand U2679 (N_2679,N_2590,N_2602);
or U2680 (N_2680,N_2606,N_2586);
nand U2681 (N_2681,N_2554,N_2590);
nand U2682 (N_2682,N_2557,N_2575);
nand U2683 (N_2683,N_2621,N_2577);
nand U2684 (N_2684,N_2618,N_2581);
and U2685 (N_2685,N_2574,N_2562);
xor U2686 (N_2686,N_2587,N_2582);
nor U2687 (N_2687,N_2596,N_2600);
and U2688 (N_2688,N_2589,N_2624);
and U2689 (N_2689,N_2554,N_2555);
nor U2690 (N_2690,N_2553,N_2605);
or U2691 (N_2691,N_2571,N_2604);
nand U2692 (N_2692,N_2619,N_2566);
nand U2693 (N_2693,N_2590,N_2607);
nand U2694 (N_2694,N_2612,N_2575);
nor U2695 (N_2695,N_2585,N_2580);
and U2696 (N_2696,N_2586,N_2573);
nor U2697 (N_2697,N_2556,N_2559);
nor U2698 (N_2698,N_2553,N_2620);
nor U2699 (N_2699,N_2569,N_2582);
and U2700 (N_2700,N_2693,N_2658);
and U2701 (N_2701,N_2652,N_2669);
nor U2702 (N_2702,N_2643,N_2640);
nand U2703 (N_2703,N_2689,N_2667);
and U2704 (N_2704,N_2692,N_2639);
or U2705 (N_2705,N_2690,N_2694);
and U2706 (N_2706,N_2696,N_2680);
nor U2707 (N_2707,N_2674,N_2671);
nor U2708 (N_2708,N_2633,N_2698);
and U2709 (N_2709,N_2697,N_2654);
nand U2710 (N_2710,N_2648,N_2655);
nor U2711 (N_2711,N_2675,N_2656);
and U2712 (N_2712,N_2657,N_2672);
nand U2713 (N_2713,N_2676,N_2683);
or U2714 (N_2714,N_2645,N_2646);
and U2715 (N_2715,N_2631,N_2681);
nand U2716 (N_2716,N_2673,N_2630);
and U2717 (N_2717,N_2695,N_2660);
nor U2718 (N_2718,N_2641,N_2628);
nand U2719 (N_2719,N_2663,N_2626);
nor U2720 (N_2720,N_2666,N_2635);
or U2721 (N_2721,N_2627,N_2691);
nand U2722 (N_2722,N_2634,N_2638);
xnor U2723 (N_2723,N_2662,N_2688);
nand U2724 (N_2724,N_2647,N_2625);
nor U2725 (N_2725,N_2632,N_2642);
or U2726 (N_2726,N_2653,N_2685);
nor U2727 (N_2727,N_2649,N_2651);
nand U2728 (N_2728,N_2687,N_2659);
nor U2729 (N_2729,N_2661,N_2678);
nand U2730 (N_2730,N_2668,N_2636);
nor U2731 (N_2731,N_2684,N_2664);
or U2732 (N_2732,N_2629,N_2679);
nor U2733 (N_2733,N_2677,N_2682);
or U2734 (N_2734,N_2699,N_2650);
and U2735 (N_2735,N_2686,N_2670);
and U2736 (N_2736,N_2637,N_2644);
nand U2737 (N_2737,N_2665,N_2690);
or U2738 (N_2738,N_2661,N_2654);
nand U2739 (N_2739,N_2699,N_2654);
nor U2740 (N_2740,N_2693,N_2645);
and U2741 (N_2741,N_2635,N_2643);
nand U2742 (N_2742,N_2625,N_2652);
and U2743 (N_2743,N_2695,N_2676);
and U2744 (N_2744,N_2648,N_2687);
nand U2745 (N_2745,N_2661,N_2692);
and U2746 (N_2746,N_2653,N_2657);
or U2747 (N_2747,N_2639,N_2688);
nor U2748 (N_2748,N_2677,N_2691);
and U2749 (N_2749,N_2693,N_2643);
nor U2750 (N_2750,N_2697,N_2680);
or U2751 (N_2751,N_2684,N_2627);
nand U2752 (N_2752,N_2644,N_2680);
or U2753 (N_2753,N_2656,N_2653);
nand U2754 (N_2754,N_2695,N_2690);
or U2755 (N_2755,N_2658,N_2646);
nand U2756 (N_2756,N_2643,N_2689);
nor U2757 (N_2757,N_2647,N_2684);
xnor U2758 (N_2758,N_2690,N_2663);
or U2759 (N_2759,N_2657,N_2691);
nand U2760 (N_2760,N_2633,N_2699);
xor U2761 (N_2761,N_2684,N_2678);
and U2762 (N_2762,N_2641,N_2666);
nor U2763 (N_2763,N_2659,N_2650);
or U2764 (N_2764,N_2671,N_2644);
or U2765 (N_2765,N_2687,N_2696);
and U2766 (N_2766,N_2681,N_2698);
and U2767 (N_2767,N_2666,N_2683);
or U2768 (N_2768,N_2687,N_2634);
nand U2769 (N_2769,N_2652,N_2695);
nor U2770 (N_2770,N_2677,N_2685);
nor U2771 (N_2771,N_2646,N_2662);
nand U2772 (N_2772,N_2673,N_2653);
nor U2773 (N_2773,N_2677,N_2697);
and U2774 (N_2774,N_2659,N_2686);
nand U2775 (N_2775,N_2717,N_2706);
nand U2776 (N_2776,N_2728,N_2748);
nor U2777 (N_2777,N_2703,N_2749);
nand U2778 (N_2778,N_2729,N_2708);
and U2779 (N_2779,N_2762,N_2715);
nand U2780 (N_2780,N_2746,N_2716);
xor U2781 (N_2781,N_2734,N_2711);
nand U2782 (N_2782,N_2764,N_2763);
nand U2783 (N_2783,N_2705,N_2740);
and U2784 (N_2784,N_2719,N_2738);
and U2785 (N_2785,N_2720,N_2713);
nor U2786 (N_2786,N_2743,N_2723);
and U2787 (N_2787,N_2773,N_2701);
or U2788 (N_2788,N_2759,N_2768);
nand U2789 (N_2789,N_2767,N_2712);
or U2790 (N_2790,N_2752,N_2747);
nor U2791 (N_2791,N_2700,N_2718);
nor U2792 (N_2792,N_2761,N_2757);
or U2793 (N_2793,N_2731,N_2758);
nand U2794 (N_2794,N_2769,N_2735);
xor U2795 (N_2795,N_2755,N_2766);
nor U2796 (N_2796,N_2704,N_2760);
and U2797 (N_2797,N_2737,N_2709);
or U2798 (N_2798,N_2765,N_2742);
nand U2799 (N_2799,N_2736,N_2721);
and U2800 (N_2800,N_2739,N_2741);
nand U2801 (N_2801,N_2772,N_2732);
or U2802 (N_2802,N_2756,N_2745);
and U2803 (N_2803,N_2770,N_2751);
nand U2804 (N_2804,N_2730,N_2722);
nor U2805 (N_2805,N_2714,N_2733);
and U2806 (N_2806,N_2771,N_2744);
and U2807 (N_2807,N_2710,N_2702);
and U2808 (N_2808,N_2707,N_2753);
nand U2809 (N_2809,N_2724,N_2727);
or U2810 (N_2810,N_2725,N_2774);
nand U2811 (N_2811,N_2726,N_2754);
nand U2812 (N_2812,N_2750,N_2747);
and U2813 (N_2813,N_2748,N_2743);
and U2814 (N_2814,N_2720,N_2773);
or U2815 (N_2815,N_2742,N_2764);
nor U2816 (N_2816,N_2763,N_2727);
nand U2817 (N_2817,N_2738,N_2740);
nor U2818 (N_2818,N_2700,N_2729);
and U2819 (N_2819,N_2742,N_2703);
nor U2820 (N_2820,N_2704,N_2751);
or U2821 (N_2821,N_2753,N_2770);
nand U2822 (N_2822,N_2732,N_2770);
nand U2823 (N_2823,N_2719,N_2747);
nand U2824 (N_2824,N_2719,N_2702);
nand U2825 (N_2825,N_2758,N_2710);
nand U2826 (N_2826,N_2758,N_2726);
nand U2827 (N_2827,N_2727,N_2768);
nand U2828 (N_2828,N_2748,N_2716);
and U2829 (N_2829,N_2700,N_2704);
nand U2830 (N_2830,N_2739,N_2703);
or U2831 (N_2831,N_2734,N_2722);
or U2832 (N_2832,N_2743,N_2722);
or U2833 (N_2833,N_2743,N_2720);
nor U2834 (N_2834,N_2701,N_2732);
nor U2835 (N_2835,N_2712,N_2713);
and U2836 (N_2836,N_2766,N_2714);
nand U2837 (N_2837,N_2701,N_2708);
and U2838 (N_2838,N_2712,N_2720);
nor U2839 (N_2839,N_2755,N_2708);
nor U2840 (N_2840,N_2712,N_2748);
and U2841 (N_2841,N_2741,N_2744);
and U2842 (N_2842,N_2747,N_2717);
nand U2843 (N_2843,N_2765,N_2750);
or U2844 (N_2844,N_2766,N_2712);
or U2845 (N_2845,N_2735,N_2702);
and U2846 (N_2846,N_2705,N_2743);
nand U2847 (N_2847,N_2716,N_2745);
and U2848 (N_2848,N_2774,N_2712);
and U2849 (N_2849,N_2751,N_2724);
and U2850 (N_2850,N_2780,N_2819);
nand U2851 (N_2851,N_2818,N_2795);
nor U2852 (N_2852,N_2804,N_2805);
and U2853 (N_2853,N_2844,N_2789);
nand U2854 (N_2854,N_2782,N_2794);
or U2855 (N_2855,N_2812,N_2811);
nand U2856 (N_2856,N_2828,N_2824);
and U2857 (N_2857,N_2842,N_2796);
or U2858 (N_2858,N_2832,N_2843);
and U2859 (N_2859,N_2830,N_2841);
nor U2860 (N_2860,N_2839,N_2799);
or U2861 (N_2861,N_2810,N_2836);
nor U2862 (N_2862,N_2803,N_2833);
nor U2863 (N_2863,N_2845,N_2790);
nand U2864 (N_2864,N_2835,N_2847);
nor U2865 (N_2865,N_2776,N_2813);
or U2866 (N_2866,N_2787,N_2781);
or U2867 (N_2867,N_2829,N_2808);
and U2868 (N_2868,N_2816,N_2792);
nand U2869 (N_2869,N_2801,N_2807);
nor U2870 (N_2870,N_2783,N_2834);
nor U2871 (N_2871,N_2814,N_2797);
nand U2872 (N_2872,N_2815,N_2775);
nand U2873 (N_2873,N_2846,N_2802);
nand U2874 (N_2874,N_2798,N_2822);
or U2875 (N_2875,N_2784,N_2838);
or U2876 (N_2876,N_2820,N_2777);
nor U2877 (N_2877,N_2806,N_2788);
nor U2878 (N_2878,N_2821,N_2848);
nor U2879 (N_2879,N_2817,N_2793);
nor U2880 (N_2880,N_2831,N_2823);
nor U2881 (N_2881,N_2825,N_2786);
nor U2882 (N_2882,N_2840,N_2849);
and U2883 (N_2883,N_2809,N_2800);
nand U2884 (N_2884,N_2779,N_2778);
xor U2885 (N_2885,N_2785,N_2827);
and U2886 (N_2886,N_2826,N_2837);
and U2887 (N_2887,N_2791,N_2813);
nor U2888 (N_2888,N_2802,N_2830);
and U2889 (N_2889,N_2845,N_2824);
or U2890 (N_2890,N_2838,N_2816);
nor U2891 (N_2891,N_2833,N_2831);
and U2892 (N_2892,N_2776,N_2810);
and U2893 (N_2893,N_2808,N_2846);
and U2894 (N_2894,N_2820,N_2800);
or U2895 (N_2895,N_2806,N_2843);
nand U2896 (N_2896,N_2819,N_2798);
and U2897 (N_2897,N_2848,N_2790);
and U2898 (N_2898,N_2821,N_2833);
and U2899 (N_2899,N_2820,N_2806);
and U2900 (N_2900,N_2783,N_2832);
nor U2901 (N_2901,N_2794,N_2777);
and U2902 (N_2902,N_2839,N_2806);
or U2903 (N_2903,N_2832,N_2849);
nand U2904 (N_2904,N_2841,N_2790);
nor U2905 (N_2905,N_2795,N_2779);
xor U2906 (N_2906,N_2797,N_2816);
xnor U2907 (N_2907,N_2797,N_2821);
nand U2908 (N_2908,N_2844,N_2826);
and U2909 (N_2909,N_2846,N_2814);
nand U2910 (N_2910,N_2817,N_2820);
and U2911 (N_2911,N_2830,N_2823);
or U2912 (N_2912,N_2799,N_2846);
nand U2913 (N_2913,N_2836,N_2782);
nor U2914 (N_2914,N_2835,N_2788);
nand U2915 (N_2915,N_2828,N_2812);
or U2916 (N_2916,N_2802,N_2825);
and U2917 (N_2917,N_2778,N_2844);
nand U2918 (N_2918,N_2778,N_2838);
nor U2919 (N_2919,N_2829,N_2798);
nor U2920 (N_2920,N_2840,N_2809);
nor U2921 (N_2921,N_2794,N_2849);
and U2922 (N_2922,N_2820,N_2848);
nor U2923 (N_2923,N_2781,N_2823);
nand U2924 (N_2924,N_2841,N_2807);
nor U2925 (N_2925,N_2900,N_2919);
nor U2926 (N_2926,N_2889,N_2920);
nand U2927 (N_2927,N_2863,N_2911);
nand U2928 (N_2928,N_2906,N_2883);
nand U2929 (N_2929,N_2875,N_2890);
and U2930 (N_2930,N_2877,N_2871);
and U2931 (N_2931,N_2893,N_2864);
nand U2932 (N_2932,N_2891,N_2905);
and U2933 (N_2933,N_2880,N_2850);
or U2934 (N_2934,N_2859,N_2868);
nor U2935 (N_2935,N_2885,N_2903);
nor U2936 (N_2936,N_2853,N_2898);
nand U2937 (N_2937,N_2901,N_2886);
nor U2938 (N_2938,N_2854,N_2897);
nor U2939 (N_2939,N_2922,N_2851);
or U2940 (N_2940,N_2908,N_2895);
and U2941 (N_2941,N_2862,N_2872);
or U2942 (N_2942,N_2865,N_2907);
nand U2943 (N_2943,N_2887,N_2896);
nor U2944 (N_2944,N_2857,N_2852);
or U2945 (N_2945,N_2855,N_2866);
and U2946 (N_2946,N_2910,N_2916);
or U2947 (N_2947,N_2902,N_2904);
and U2948 (N_2948,N_2892,N_2917);
and U2949 (N_2949,N_2869,N_2921);
nand U2950 (N_2950,N_2888,N_2894);
xor U2951 (N_2951,N_2915,N_2867);
nor U2952 (N_2952,N_2879,N_2861);
nand U2953 (N_2953,N_2881,N_2874);
and U2954 (N_2954,N_2856,N_2899);
or U2955 (N_2955,N_2882,N_2924);
nor U2956 (N_2956,N_2912,N_2873);
and U2957 (N_2957,N_2914,N_2860);
and U2958 (N_2958,N_2913,N_2909);
or U2959 (N_2959,N_2878,N_2876);
or U2960 (N_2960,N_2918,N_2858);
nand U2961 (N_2961,N_2870,N_2884);
or U2962 (N_2962,N_2923,N_2912);
nand U2963 (N_2963,N_2911,N_2910);
nor U2964 (N_2964,N_2865,N_2895);
nor U2965 (N_2965,N_2906,N_2859);
nor U2966 (N_2966,N_2875,N_2886);
or U2967 (N_2967,N_2915,N_2873);
nor U2968 (N_2968,N_2884,N_2921);
nor U2969 (N_2969,N_2890,N_2863);
nand U2970 (N_2970,N_2877,N_2879);
or U2971 (N_2971,N_2920,N_2899);
nand U2972 (N_2972,N_2906,N_2899);
or U2973 (N_2973,N_2880,N_2870);
and U2974 (N_2974,N_2923,N_2901);
and U2975 (N_2975,N_2919,N_2902);
and U2976 (N_2976,N_2887,N_2914);
nand U2977 (N_2977,N_2909,N_2868);
nor U2978 (N_2978,N_2876,N_2858);
or U2979 (N_2979,N_2861,N_2895);
nor U2980 (N_2980,N_2853,N_2892);
nand U2981 (N_2981,N_2905,N_2887);
nor U2982 (N_2982,N_2890,N_2893);
or U2983 (N_2983,N_2853,N_2885);
and U2984 (N_2984,N_2913,N_2869);
or U2985 (N_2985,N_2858,N_2901);
nand U2986 (N_2986,N_2875,N_2918);
nand U2987 (N_2987,N_2856,N_2887);
nand U2988 (N_2988,N_2876,N_2880);
and U2989 (N_2989,N_2881,N_2879);
and U2990 (N_2990,N_2911,N_2868);
nor U2991 (N_2991,N_2912,N_2870);
nand U2992 (N_2992,N_2891,N_2883);
nand U2993 (N_2993,N_2865,N_2915);
or U2994 (N_2994,N_2868,N_2906);
and U2995 (N_2995,N_2889,N_2862);
or U2996 (N_2996,N_2909,N_2910);
or U2997 (N_2997,N_2866,N_2896);
nor U2998 (N_2998,N_2858,N_2881);
nand U2999 (N_2999,N_2880,N_2889);
or UO_0 (O_0,N_2950,N_2977);
nand UO_1 (O_1,N_2971,N_2994);
or UO_2 (O_2,N_2926,N_2949);
nor UO_3 (O_3,N_2939,N_2993);
or UO_4 (O_4,N_2938,N_2969);
and UO_5 (O_5,N_2927,N_2944);
or UO_6 (O_6,N_2995,N_2946);
or UO_7 (O_7,N_2933,N_2992);
and UO_8 (O_8,N_2988,N_2956);
and UO_9 (O_9,N_2940,N_2998);
nand UO_10 (O_10,N_2935,N_2964);
nand UO_11 (O_11,N_2955,N_2930);
nand UO_12 (O_12,N_2962,N_2960);
nand UO_13 (O_13,N_2970,N_2997);
nand UO_14 (O_14,N_2932,N_2973);
and UO_15 (O_15,N_2979,N_2996);
and UO_16 (O_16,N_2929,N_2931);
nor UO_17 (O_17,N_2957,N_2976);
nor UO_18 (O_18,N_2958,N_2983);
nand UO_19 (O_19,N_2981,N_2954);
nor UO_20 (O_20,N_2959,N_2942);
or UO_21 (O_21,N_2963,N_2934);
nand UO_22 (O_22,N_2941,N_2943);
nand UO_23 (O_23,N_2987,N_2952);
or UO_24 (O_24,N_2986,N_2989);
or UO_25 (O_25,N_2936,N_2948);
nand UO_26 (O_26,N_2982,N_2972);
and UO_27 (O_27,N_2975,N_2978);
nor UO_28 (O_28,N_2980,N_2974);
nand UO_29 (O_29,N_2999,N_2945);
nor UO_30 (O_30,N_2953,N_2925);
xor UO_31 (O_31,N_2951,N_2991);
nor UO_32 (O_32,N_2928,N_2937);
and UO_33 (O_33,N_2966,N_2990);
nand UO_34 (O_34,N_2967,N_2947);
nor UO_35 (O_35,N_2965,N_2968);
nor UO_36 (O_36,N_2961,N_2984);
nor UO_37 (O_37,N_2985,N_2992);
nand UO_38 (O_38,N_2950,N_2976);
nor UO_39 (O_39,N_2983,N_2984);
or UO_40 (O_40,N_2949,N_2993);
or UO_41 (O_41,N_2959,N_2928);
or UO_42 (O_42,N_2983,N_2928);
or UO_43 (O_43,N_2933,N_2980);
nor UO_44 (O_44,N_2986,N_2979);
nor UO_45 (O_45,N_2945,N_2994);
and UO_46 (O_46,N_2925,N_2989);
nand UO_47 (O_47,N_2963,N_2979);
and UO_48 (O_48,N_2989,N_2946);
nor UO_49 (O_49,N_2947,N_2971);
and UO_50 (O_50,N_2983,N_2969);
nand UO_51 (O_51,N_2948,N_2930);
nor UO_52 (O_52,N_2962,N_2978);
nand UO_53 (O_53,N_2958,N_2995);
and UO_54 (O_54,N_2942,N_2973);
nand UO_55 (O_55,N_2993,N_2936);
or UO_56 (O_56,N_2933,N_2956);
and UO_57 (O_57,N_2934,N_2993);
nand UO_58 (O_58,N_2958,N_2950);
nor UO_59 (O_59,N_2976,N_2987);
nor UO_60 (O_60,N_2983,N_2935);
nand UO_61 (O_61,N_2969,N_2982);
or UO_62 (O_62,N_2967,N_2973);
or UO_63 (O_63,N_2970,N_2961);
nand UO_64 (O_64,N_2970,N_2940);
and UO_65 (O_65,N_2984,N_2949);
and UO_66 (O_66,N_2981,N_2961);
nor UO_67 (O_67,N_2940,N_2939);
nor UO_68 (O_68,N_2938,N_2987);
nor UO_69 (O_69,N_2935,N_2942);
nor UO_70 (O_70,N_2964,N_2999);
nor UO_71 (O_71,N_2971,N_2972);
or UO_72 (O_72,N_2990,N_2971);
or UO_73 (O_73,N_2994,N_2960);
nand UO_74 (O_74,N_2931,N_2978);
nor UO_75 (O_75,N_2943,N_2947);
or UO_76 (O_76,N_2973,N_2976);
nand UO_77 (O_77,N_2979,N_2947);
or UO_78 (O_78,N_2933,N_2987);
nand UO_79 (O_79,N_2951,N_2952);
or UO_80 (O_80,N_2946,N_2973);
nand UO_81 (O_81,N_2939,N_2979);
nand UO_82 (O_82,N_2925,N_2941);
nor UO_83 (O_83,N_2997,N_2934);
nor UO_84 (O_84,N_2947,N_2996);
nand UO_85 (O_85,N_2996,N_2933);
nor UO_86 (O_86,N_2927,N_2977);
or UO_87 (O_87,N_2949,N_2966);
nand UO_88 (O_88,N_2979,N_2985);
nand UO_89 (O_89,N_2966,N_2974);
nand UO_90 (O_90,N_2926,N_2943);
and UO_91 (O_91,N_2943,N_2988);
and UO_92 (O_92,N_2961,N_2956);
and UO_93 (O_93,N_2984,N_2939);
or UO_94 (O_94,N_2934,N_2961);
nand UO_95 (O_95,N_2937,N_2930);
and UO_96 (O_96,N_2942,N_2950);
nor UO_97 (O_97,N_2987,N_2948);
nor UO_98 (O_98,N_2949,N_2980);
and UO_99 (O_99,N_2978,N_2940);
or UO_100 (O_100,N_2957,N_2967);
and UO_101 (O_101,N_2936,N_2995);
nand UO_102 (O_102,N_2993,N_2945);
or UO_103 (O_103,N_2951,N_2994);
nor UO_104 (O_104,N_2953,N_2974);
nor UO_105 (O_105,N_2947,N_2998);
nor UO_106 (O_106,N_2929,N_2943);
and UO_107 (O_107,N_2977,N_2953);
nor UO_108 (O_108,N_2985,N_2976);
and UO_109 (O_109,N_2978,N_2988);
and UO_110 (O_110,N_2956,N_2991);
or UO_111 (O_111,N_2977,N_2968);
or UO_112 (O_112,N_2936,N_2943);
or UO_113 (O_113,N_2955,N_2976);
or UO_114 (O_114,N_2960,N_2944);
nor UO_115 (O_115,N_2946,N_2926);
and UO_116 (O_116,N_2949,N_2982);
and UO_117 (O_117,N_2996,N_2991);
and UO_118 (O_118,N_2946,N_2949);
or UO_119 (O_119,N_2951,N_2959);
or UO_120 (O_120,N_2957,N_2958);
and UO_121 (O_121,N_2985,N_2947);
and UO_122 (O_122,N_2995,N_2973);
or UO_123 (O_123,N_2991,N_2985);
nor UO_124 (O_124,N_2940,N_2985);
nand UO_125 (O_125,N_2957,N_2960);
nand UO_126 (O_126,N_2952,N_2961);
or UO_127 (O_127,N_2929,N_2982);
or UO_128 (O_128,N_2944,N_2970);
nor UO_129 (O_129,N_2974,N_2936);
nor UO_130 (O_130,N_2959,N_2965);
nand UO_131 (O_131,N_2936,N_2954);
nand UO_132 (O_132,N_2968,N_2942);
nand UO_133 (O_133,N_2964,N_2981);
nor UO_134 (O_134,N_2977,N_2928);
or UO_135 (O_135,N_2998,N_2945);
and UO_136 (O_136,N_2996,N_2969);
nor UO_137 (O_137,N_2980,N_2971);
and UO_138 (O_138,N_2997,N_2982);
nor UO_139 (O_139,N_2969,N_2945);
or UO_140 (O_140,N_2933,N_2947);
nand UO_141 (O_141,N_2948,N_2966);
nand UO_142 (O_142,N_2978,N_2976);
nand UO_143 (O_143,N_2975,N_2959);
or UO_144 (O_144,N_2951,N_2990);
nor UO_145 (O_145,N_2937,N_2940);
or UO_146 (O_146,N_2968,N_2943);
or UO_147 (O_147,N_2965,N_2998);
or UO_148 (O_148,N_2961,N_2951);
nand UO_149 (O_149,N_2933,N_2937);
nor UO_150 (O_150,N_2955,N_2941);
nor UO_151 (O_151,N_2965,N_2995);
nor UO_152 (O_152,N_2996,N_2962);
nand UO_153 (O_153,N_2986,N_2991);
nand UO_154 (O_154,N_2926,N_2967);
nand UO_155 (O_155,N_2935,N_2991);
and UO_156 (O_156,N_2977,N_2984);
or UO_157 (O_157,N_2990,N_2977);
and UO_158 (O_158,N_2955,N_2927);
and UO_159 (O_159,N_2993,N_2959);
or UO_160 (O_160,N_2948,N_2979);
or UO_161 (O_161,N_2962,N_2930);
nand UO_162 (O_162,N_2960,N_2930);
nand UO_163 (O_163,N_2955,N_2942);
and UO_164 (O_164,N_2927,N_2930);
nor UO_165 (O_165,N_2952,N_2972);
nor UO_166 (O_166,N_2993,N_2958);
or UO_167 (O_167,N_2993,N_2981);
nor UO_168 (O_168,N_2959,N_2937);
or UO_169 (O_169,N_2963,N_2981);
nor UO_170 (O_170,N_2962,N_2949);
nor UO_171 (O_171,N_2971,N_2957);
and UO_172 (O_172,N_2934,N_2931);
nor UO_173 (O_173,N_2992,N_2988);
or UO_174 (O_174,N_2926,N_2966);
nor UO_175 (O_175,N_2948,N_2943);
and UO_176 (O_176,N_2986,N_2976);
nand UO_177 (O_177,N_2990,N_2961);
nand UO_178 (O_178,N_2966,N_2975);
and UO_179 (O_179,N_2978,N_2952);
and UO_180 (O_180,N_2951,N_2980);
or UO_181 (O_181,N_2932,N_2937);
and UO_182 (O_182,N_2959,N_2933);
and UO_183 (O_183,N_2949,N_2932);
and UO_184 (O_184,N_2944,N_2998);
nand UO_185 (O_185,N_2968,N_2952);
or UO_186 (O_186,N_2971,N_2974);
and UO_187 (O_187,N_2936,N_2933);
nand UO_188 (O_188,N_2956,N_2984);
nand UO_189 (O_189,N_2968,N_2971);
nor UO_190 (O_190,N_2948,N_2945);
or UO_191 (O_191,N_2926,N_2941);
nand UO_192 (O_192,N_2978,N_2947);
and UO_193 (O_193,N_2938,N_2991);
nand UO_194 (O_194,N_2970,N_2935);
and UO_195 (O_195,N_2964,N_2957);
nand UO_196 (O_196,N_2988,N_2939);
nand UO_197 (O_197,N_2982,N_2928);
and UO_198 (O_198,N_2940,N_2954);
and UO_199 (O_199,N_2944,N_2925);
or UO_200 (O_200,N_2944,N_2964);
nor UO_201 (O_201,N_2979,N_2936);
nand UO_202 (O_202,N_2968,N_2990);
or UO_203 (O_203,N_2942,N_2963);
nand UO_204 (O_204,N_2983,N_2955);
and UO_205 (O_205,N_2931,N_2990);
or UO_206 (O_206,N_2958,N_2969);
or UO_207 (O_207,N_2953,N_2966);
or UO_208 (O_208,N_2992,N_2945);
nor UO_209 (O_209,N_2974,N_2988);
nand UO_210 (O_210,N_2937,N_2952);
nand UO_211 (O_211,N_2994,N_2983);
and UO_212 (O_212,N_2954,N_2999);
or UO_213 (O_213,N_2936,N_2997);
or UO_214 (O_214,N_2929,N_2997);
or UO_215 (O_215,N_2943,N_2945);
nand UO_216 (O_216,N_2962,N_2950);
nor UO_217 (O_217,N_2971,N_2959);
and UO_218 (O_218,N_2981,N_2956);
and UO_219 (O_219,N_2938,N_2973);
and UO_220 (O_220,N_2978,N_2996);
nor UO_221 (O_221,N_2998,N_2978);
nor UO_222 (O_222,N_2959,N_2983);
or UO_223 (O_223,N_2926,N_2954);
nor UO_224 (O_224,N_2931,N_2995);
nand UO_225 (O_225,N_2961,N_2989);
nand UO_226 (O_226,N_2940,N_2929);
nand UO_227 (O_227,N_2929,N_2995);
nor UO_228 (O_228,N_2995,N_2989);
and UO_229 (O_229,N_2985,N_2997);
or UO_230 (O_230,N_2941,N_2937);
nor UO_231 (O_231,N_2952,N_2982);
or UO_232 (O_232,N_2992,N_2981);
and UO_233 (O_233,N_2959,N_2968);
or UO_234 (O_234,N_2959,N_2943);
and UO_235 (O_235,N_2972,N_2978);
xor UO_236 (O_236,N_2937,N_2950);
or UO_237 (O_237,N_2956,N_2944);
nand UO_238 (O_238,N_2942,N_2969);
or UO_239 (O_239,N_2947,N_2987);
nor UO_240 (O_240,N_2968,N_2949);
nand UO_241 (O_241,N_2978,N_2970);
or UO_242 (O_242,N_2960,N_2932);
and UO_243 (O_243,N_2967,N_2975);
nor UO_244 (O_244,N_2931,N_2959);
nand UO_245 (O_245,N_2944,N_2980);
and UO_246 (O_246,N_2982,N_2938);
and UO_247 (O_247,N_2929,N_2984);
nand UO_248 (O_248,N_2947,N_2997);
and UO_249 (O_249,N_2956,N_2997);
and UO_250 (O_250,N_2994,N_2936);
nand UO_251 (O_251,N_2980,N_2954);
nand UO_252 (O_252,N_2989,N_2930);
nor UO_253 (O_253,N_2969,N_2929);
or UO_254 (O_254,N_2950,N_2951);
nand UO_255 (O_255,N_2942,N_2992);
nor UO_256 (O_256,N_2967,N_2959);
and UO_257 (O_257,N_2944,N_2974);
nor UO_258 (O_258,N_2988,N_2959);
or UO_259 (O_259,N_2990,N_2942);
or UO_260 (O_260,N_2928,N_2931);
or UO_261 (O_261,N_2946,N_2933);
nand UO_262 (O_262,N_2942,N_2930);
or UO_263 (O_263,N_2982,N_2943);
nand UO_264 (O_264,N_2928,N_2979);
and UO_265 (O_265,N_2970,N_2956);
nand UO_266 (O_266,N_2965,N_2985);
and UO_267 (O_267,N_2945,N_2944);
or UO_268 (O_268,N_2991,N_2957);
xnor UO_269 (O_269,N_2929,N_2976);
nand UO_270 (O_270,N_2993,N_2976);
or UO_271 (O_271,N_2969,N_2946);
nor UO_272 (O_272,N_2960,N_2934);
or UO_273 (O_273,N_2981,N_2937);
nor UO_274 (O_274,N_2998,N_2929);
and UO_275 (O_275,N_2932,N_2945);
nand UO_276 (O_276,N_2932,N_2996);
and UO_277 (O_277,N_2964,N_2939);
xor UO_278 (O_278,N_2962,N_2989);
nand UO_279 (O_279,N_2979,N_2927);
or UO_280 (O_280,N_2935,N_2936);
or UO_281 (O_281,N_2998,N_2966);
and UO_282 (O_282,N_2975,N_2945);
nor UO_283 (O_283,N_2946,N_2963);
nand UO_284 (O_284,N_2996,N_2990);
and UO_285 (O_285,N_2959,N_2976);
nor UO_286 (O_286,N_2949,N_2929);
nand UO_287 (O_287,N_2999,N_2973);
nand UO_288 (O_288,N_2938,N_2981);
or UO_289 (O_289,N_2953,N_2979);
or UO_290 (O_290,N_2946,N_2948);
nor UO_291 (O_291,N_2982,N_2953);
nor UO_292 (O_292,N_2996,N_2989);
or UO_293 (O_293,N_2940,N_2963);
and UO_294 (O_294,N_2964,N_2936);
or UO_295 (O_295,N_2963,N_2996);
and UO_296 (O_296,N_2989,N_2983);
or UO_297 (O_297,N_2931,N_2932);
or UO_298 (O_298,N_2997,N_2938);
nor UO_299 (O_299,N_2997,N_2981);
nor UO_300 (O_300,N_2967,N_2951);
nand UO_301 (O_301,N_2951,N_2964);
or UO_302 (O_302,N_2947,N_2934);
and UO_303 (O_303,N_2961,N_2982);
nand UO_304 (O_304,N_2984,N_2970);
nand UO_305 (O_305,N_2952,N_2995);
or UO_306 (O_306,N_2989,N_2981);
nand UO_307 (O_307,N_2957,N_2953);
nand UO_308 (O_308,N_2991,N_2978);
and UO_309 (O_309,N_2987,N_2989);
or UO_310 (O_310,N_2982,N_2926);
nand UO_311 (O_311,N_2947,N_2993);
and UO_312 (O_312,N_2971,N_2996);
nor UO_313 (O_313,N_2957,N_2926);
nand UO_314 (O_314,N_2983,N_2952);
nand UO_315 (O_315,N_2987,N_2932);
or UO_316 (O_316,N_2977,N_2933);
nor UO_317 (O_317,N_2952,N_2934);
or UO_318 (O_318,N_2982,N_2965);
nand UO_319 (O_319,N_2953,N_2976);
or UO_320 (O_320,N_2978,N_2957);
nand UO_321 (O_321,N_2954,N_2929);
nor UO_322 (O_322,N_2975,N_2937);
nor UO_323 (O_323,N_2975,N_2977);
or UO_324 (O_324,N_2983,N_2999);
and UO_325 (O_325,N_2958,N_2944);
nand UO_326 (O_326,N_2970,N_2941);
or UO_327 (O_327,N_2993,N_2954);
and UO_328 (O_328,N_2977,N_2930);
nand UO_329 (O_329,N_2960,N_2926);
nor UO_330 (O_330,N_2994,N_2996);
nor UO_331 (O_331,N_2932,N_2947);
and UO_332 (O_332,N_2980,N_2937);
nor UO_333 (O_333,N_2962,N_2936);
or UO_334 (O_334,N_2994,N_2953);
and UO_335 (O_335,N_2984,N_2959);
nor UO_336 (O_336,N_2946,N_2958);
and UO_337 (O_337,N_2998,N_2936);
nand UO_338 (O_338,N_2990,N_2956);
nand UO_339 (O_339,N_2983,N_2974);
nor UO_340 (O_340,N_2991,N_2994);
nand UO_341 (O_341,N_2951,N_2983);
and UO_342 (O_342,N_2944,N_2950);
and UO_343 (O_343,N_2973,N_2954);
or UO_344 (O_344,N_2977,N_2996);
nand UO_345 (O_345,N_2997,N_2954);
and UO_346 (O_346,N_2976,N_2961);
or UO_347 (O_347,N_2971,N_2995);
or UO_348 (O_348,N_2995,N_2969);
and UO_349 (O_349,N_2991,N_2967);
or UO_350 (O_350,N_2956,N_2996);
and UO_351 (O_351,N_2937,N_2973);
nand UO_352 (O_352,N_2988,N_2996);
and UO_353 (O_353,N_2931,N_2940);
nor UO_354 (O_354,N_2978,N_2942);
and UO_355 (O_355,N_2935,N_2978);
and UO_356 (O_356,N_2970,N_2925);
nor UO_357 (O_357,N_2972,N_2946);
nand UO_358 (O_358,N_2990,N_2949);
and UO_359 (O_359,N_2961,N_2930);
and UO_360 (O_360,N_2953,N_2967);
nand UO_361 (O_361,N_2998,N_2994);
or UO_362 (O_362,N_2965,N_2956);
nand UO_363 (O_363,N_2982,N_2978);
or UO_364 (O_364,N_2928,N_2978);
nor UO_365 (O_365,N_2929,N_2974);
or UO_366 (O_366,N_2959,N_2949);
and UO_367 (O_367,N_2989,N_2973);
or UO_368 (O_368,N_2934,N_2933);
and UO_369 (O_369,N_2987,N_2991);
nand UO_370 (O_370,N_2985,N_2969);
or UO_371 (O_371,N_2964,N_2980);
nand UO_372 (O_372,N_2935,N_2959);
nand UO_373 (O_373,N_2988,N_2967);
or UO_374 (O_374,N_2931,N_2933);
nor UO_375 (O_375,N_2951,N_2982);
and UO_376 (O_376,N_2997,N_2948);
or UO_377 (O_377,N_2940,N_2955);
and UO_378 (O_378,N_2959,N_2952);
nor UO_379 (O_379,N_2957,N_2962);
nand UO_380 (O_380,N_2996,N_2967);
or UO_381 (O_381,N_2957,N_2943);
nor UO_382 (O_382,N_2952,N_2962);
nor UO_383 (O_383,N_2933,N_2993);
nand UO_384 (O_384,N_2947,N_2946);
nand UO_385 (O_385,N_2984,N_2990);
or UO_386 (O_386,N_2989,N_2999);
or UO_387 (O_387,N_2931,N_2980);
or UO_388 (O_388,N_2949,N_2927);
or UO_389 (O_389,N_2967,N_2993);
and UO_390 (O_390,N_2932,N_2941);
xnor UO_391 (O_391,N_2952,N_2945);
and UO_392 (O_392,N_2966,N_2995);
nor UO_393 (O_393,N_2931,N_2997);
nor UO_394 (O_394,N_2999,N_2968);
and UO_395 (O_395,N_2957,N_2984);
or UO_396 (O_396,N_2942,N_2944);
or UO_397 (O_397,N_2986,N_2960);
xnor UO_398 (O_398,N_2937,N_2929);
nand UO_399 (O_399,N_2995,N_2959);
xnor UO_400 (O_400,N_2957,N_2987);
nor UO_401 (O_401,N_2993,N_2998);
or UO_402 (O_402,N_2933,N_2929);
or UO_403 (O_403,N_2927,N_2995);
nor UO_404 (O_404,N_2959,N_2936);
nor UO_405 (O_405,N_2955,N_2937);
or UO_406 (O_406,N_2969,N_2939);
nand UO_407 (O_407,N_2956,N_2978);
nand UO_408 (O_408,N_2956,N_2947);
or UO_409 (O_409,N_2925,N_2980);
xor UO_410 (O_410,N_2951,N_2978);
or UO_411 (O_411,N_2951,N_2995);
xnor UO_412 (O_412,N_2996,N_2928);
and UO_413 (O_413,N_2977,N_2926);
nand UO_414 (O_414,N_2960,N_2927);
nor UO_415 (O_415,N_2984,N_2946);
or UO_416 (O_416,N_2944,N_2962);
or UO_417 (O_417,N_2982,N_2936);
nor UO_418 (O_418,N_2951,N_2956);
nand UO_419 (O_419,N_2966,N_2973);
or UO_420 (O_420,N_2994,N_2973);
nand UO_421 (O_421,N_2992,N_2984);
nand UO_422 (O_422,N_2957,N_2950);
and UO_423 (O_423,N_2955,N_2971);
nor UO_424 (O_424,N_2968,N_2955);
and UO_425 (O_425,N_2928,N_2935);
nand UO_426 (O_426,N_2988,N_2985);
nor UO_427 (O_427,N_2959,N_2926);
and UO_428 (O_428,N_2932,N_2990);
nor UO_429 (O_429,N_2953,N_2930);
and UO_430 (O_430,N_2999,N_2946);
or UO_431 (O_431,N_2968,N_2939);
nand UO_432 (O_432,N_2987,N_2995);
and UO_433 (O_433,N_2982,N_2992);
and UO_434 (O_434,N_2949,N_2958);
and UO_435 (O_435,N_2963,N_2978);
or UO_436 (O_436,N_2994,N_2972);
or UO_437 (O_437,N_2945,N_2936);
nor UO_438 (O_438,N_2955,N_2992);
or UO_439 (O_439,N_2971,N_2937);
nand UO_440 (O_440,N_2946,N_2967);
nor UO_441 (O_441,N_2941,N_2974);
and UO_442 (O_442,N_2940,N_2994);
or UO_443 (O_443,N_2948,N_2992);
nand UO_444 (O_444,N_2957,N_2956);
or UO_445 (O_445,N_2960,N_2970);
or UO_446 (O_446,N_2945,N_2997);
and UO_447 (O_447,N_2985,N_2935);
nor UO_448 (O_448,N_2980,N_2927);
or UO_449 (O_449,N_2997,N_2993);
and UO_450 (O_450,N_2969,N_2986);
nand UO_451 (O_451,N_2931,N_2935);
and UO_452 (O_452,N_2995,N_2949);
and UO_453 (O_453,N_2957,N_2990);
nor UO_454 (O_454,N_2957,N_2996);
and UO_455 (O_455,N_2939,N_2955);
or UO_456 (O_456,N_2932,N_2927);
nand UO_457 (O_457,N_2947,N_2964);
or UO_458 (O_458,N_2969,N_2960);
nand UO_459 (O_459,N_2981,N_2945);
nand UO_460 (O_460,N_2972,N_2968);
nor UO_461 (O_461,N_2932,N_2936);
or UO_462 (O_462,N_2980,N_2957);
nand UO_463 (O_463,N_2995,N_2963);
nand UO_464 (O_464,N_2925,N_2940);
nand UO_465 (O_465,N_2930,N_2988);
and UO_466 (O_466,N_2960,N_2973);
nor UO_467 (O_467,N_2958,N_2933);
and UO_468 (O_468,N_2966,N_2955);
or UO_469 (O_469,N_2961,N_2960);
or UO_470 (O_470,N_2934,N_2955);
nor UO_471 (O_471,N_2960,N_2965);
nand UO_472 (O_472,N_2995,N_2996);
and UO_473 (O_473,N_2971,N_2964);
nand UO_474 (O_474,N_2975,N_2958);
and UO_475 (O_475,N_2963,N_2999);
nor UO_476 (O_476,N_2985,N_2983);
nor UO_477 (O_477,N_2987,N_2925);
and UO_478 (O_478,N_2950,N_2953);
or UO_479 (O_479,N_2939,N_2999);
nand UO_480 (O_480,N_2961,N_2974);
nor UO_481 (O_481,N_2957,N_2949);
or UO_482 (O_482,N_2937,N_2984);
nor UO_483 (O_483,N_2988,N_2997);
nand UO_484 (O_484,N_2976,N_2979);
nand UO_485 (O_485,N_2996,N_2974);
nor UO_486 (O_486,N_2994,N_2962);
nor UO_487 (O_487,N_2977,N_2991);
nor UO_488 (O_488,N_2940,N_2986);
nand UO_489 (O_489,N_2925,N_2946);
xor UO_490 (O_490,N_2962,N_2995);
or UO_491 (O_491,N_2971,N_2935);
nand UO_492 (O_492,N_2926,N_2979);
nand UO_493 (O_493,N_2967,N_2955);
nor UO_494 (O_494,N_2980,N_2959);
and UO_495 (O_495,N_2994,N_2930);
nor UO_496 (O_496,N_2935,N_2982);
nor UO_497 (O_497,N_2947,N_2948);
nand UO_498 (O_498,N_2941,N_2972);
or UO_499 (O_499,N_2955,N_2947);
endmodule