module basic_500_3000_500_60_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_484,In_410);
and U1 (N_1,In_321,In_13);
nand U2 (N_2,In_173,In_190);
nor U3 (N_3,In_59,In_87);
nand U4 (N_4,In_332,In_337);
or U5 (N_5,In_349,In_10);
and U6 (N_6,In_462,In_358);
nand U7 (N_7,In_88,In_17);
or U8 (N_8,In_4,In_89);
or U9 (N_9,In_48,In_133);
nand U10 (N_10,In_193,In_413);
nor U11 (N_11,In_288,In_379);
nor U12 (N_12,In_207,In_401);
nand U13 (N_13,In_493,In_257);
or U14 (N_14,In_440,In_252);
and U15 (N_15,In_483,In_294);
and U16 (N_16,In_452,In_97);
or U17 (N_17,In_128,In_340);
or U18 (N_18,In_351,In_138);
nor U19 (N_19,In_277,In_402);
or U20 (N_20,In_446,In_261);
nand U21 (N_21,In_110,In_375);
nand U22 (N_22,In_223,In_82);
nand U23 (N_23,In_296,In_362);
nand U24 (N_24,In_453,In_369);
or U25 (N_25,In_79,In_469);
or U26 (N_26,In_158,In_271);
and U27 (N_27,In_45,In_155);
nor U28 (N_28,In_329,In_90);
or U29 (N_29,In_154,In_5);
or U30 (N_30,In_255,In_202);
and U31 (N_31,In_253,In_224);
nand U32 (N_32,In_25,In_393);
or U33 (N_33,In_258,In_227);
nor U34 (N_34,In_474,In_436);
and U35 (N_35,In_44,In_392);
and U36 (N_36,In_194,In_54);
or U37 (N_37,In_342,In_73);
or U38 (N_38,In_335,In_274);
or U39 (N_39,In_231,In_353);
and U40 (N_40,In_419,In_459);
and U41 (N_41,In_177,In_273);
and U42 (N_42,In_414,In_303);
xnor U43 (N_43,In_400,In_75);
or U44 (N_44,In_421,In_8);
and U45 (N_45,In_112,In_473);
nor U46 (N_46,In_430,In_256);
nand U47 (N_47,In_368,In_22);
nor U48 (N_48,In_433,In_210);
nand U49 (N_49,In_361,In_39);
or U50 (N_50,In_407,N_36);
and U51 (N_51,N_48,In_55);
nor U52 (N_52,In_383,In_309);
nand U53 (N_53,In_448,In_30);
nand U54 (N_54,N_37,In_397);
and U55 (N_55,In_298,In_31);
nor U56 (N_56,In_53,In_374);
or U57 (N_57,In_416,In_239);
nand U58 (N_58,In_324,In_427);
and U59 (N_59,In_153,In_479);
and U60 (N_60,In_186,In_322);
and U61 (N_61,In_29,In_346);
nor U62 (N_62,In_310,In_144);
and U63 (N_63,In_219,In_27);
and U64 (N_64,In_56,N_28);
and U65 (N_65,In_94,N_4);
or U66 (N_66,In_142,In_12);
or U67 (N_67,In_319,In_225);
and U68 (N_68,In_377,In_381);
nor U69 (N_69,In_476,In_454);
and U70 (N_70,In_355,N_44);
nor U71 (N_71,In_344,N_16);
nor U72 (N_72,In_103,In_40);
nor U73 (N_73,In_447,In_143);
nand U74 (N_74,In_395,N_38);
or U75 (N_75,In_92,In_263);
nor U76 (N_76,In_130,N_25);
nand U77 (N_77,In_157,In_260);
nor U78 (N_78,In_187,In_9);
nor U79 (N_79,In_406,In_471);
nor U80 (N_80,In_347,In_359);
nor U81 (N_81,In_266,In_450);
and U82 (N_82,In_485,In_162);
xor U83 (N_83,In_185,In_60);
or U84 (N_84,In_293,In_443);
nor U85 (N_85,In_241,In_404);
or U86 (N_86,In_146,In_1);
nor U87 (N_87,In_119,N_5);
or U88 (N_88,In_465,In_482);
and U89 (N_89,In_478,In_64);
or U90 (N_90,In_233,In_281);
and U91 (N_91,In_279,In_308);
nand U92 (N_92,N_12,In_171);
or U93 (N_93,In_318,In_242);
and U94 (N_94,In_323,In_434);
or U95 (N_95,In_71,N_29);
or U96 (N_96,N_45,In_246);
nand U97 (N_97,N_30,In_93);
or U98 (N_98,In_262,N_43);
nor U99 (N_99,In_69,In_264);
nand U100 (N_100,In_269,In_161);
or U101 (N_101,In_78,In_109);
or U102 (N_102,N_26,In_472);
nand U103 (N_103,N_18,In_405);
nor U104 (N_104,In_115,In_411);
nand U105 (N_105,In_200,In_123);
and U106 (N_106,N_35,In_57);
nor U107 (N_107,In_166,In_84);
or U108 (N_108,In_18,In_339);
nor U109 (N_109,N_83,In_265);
nand U110 (N_110,In_350,In_438);
or U111 (N_111,N_19,In_26);
nand U112 (N_112,N_0,N_2);
nand U113 (N_113,N_57,In_126);
and U114 (N_114,In_189,In_248);
nand U115 (N_115,In_174,In_285);
nor U116 (N_116,In_304,In_147);
or U117 (N_117,In_480,In_106);
and U118 (N_118,In_498,In_209);
or U119 (N_119,In_389,In_267);
nand U120 (N_120,N_14,In_150);
nor U121 (N_121,In_399,In_311);
or U122 (N_122,In_387,N_88);
or U123 (N_123,In_102,In_65);
nand U124 (N_124,In_403,N_59);
nor U125 (N_125,In_165,In_365);
or U126 (N_126,In_116,In_328);
and U127 (N_127,In_140,In_212);
nor U128 (N_128,In_356,In_461);
or U129 (N_129,N_76,In_481);
nand U130 (N_130,In_366,N_20);
nor U131 (N_131,In_240,In_2);
or U132 (N_132,In_390,N_97);
or U133 (N_133,In_470,In_391);
nand U134 (N_134,In_348,In_238);
or U135 (N_135,N_52,In_114);
or U136 (N_136,In_178,In_47);
and U137 (N_137,In_228,N_78);
or U138 (N_138,In_292,In_297);
nand U139 (N_139,In_326,In_33);
or U140 (N_140,In_35,In_120);
nand U141 (N_141,N_3,In_132);
and U142 (N_142,In_156,In_254);
nand U143 (N_143,In_188,In_108);
nor U144 (N_144,N_56,In_287);
and U145 (N_145,N_58,In_81);
nor U146 (N_146,In_259,In_409);
and U147 (N_147,In_15,N_86);
and U148 (N_148,In_66,N_96);
nand U149 (N_149,In_497,In_289);
nand U150 (N_150,N_22,In_336);
xnor U151 (N_151,In_74,In_139);
nor U152 (N_152,In_317,In_76);
and U153 (N_153,N_103,N_99);
nor U154 (N_154,In_169,In_98);
nor U155 (N_155,In_492,N_66);
nor U156 (N_156,In_195,In_284);
xor U157 (N_157,N_74,In_159);
and U158 (N_158,In_70,In_32);
or U159 (N_159,In_0,N_89);
nor U160 (N_160,In_488,N_115);
and U161 (N_161,In_86,N_63);
nand U162 (N_162,In_251,In_179);
nand U163 (N_163,In_220,N_85);
and U164 (N_164,In_437,In_145);
nor U165 (N_165,In_117,N_116);
or U166 (N_166,In_275,In_468);
nor U167 (N_167,In_232,In_198);
and U168 (N_168,In_245,In_7);
and U169 (N_169,In_286,In_184);
or U170 (N_170,N_147,In_272);
nand U171 (N_171,In_163,N_82);
or U172 (N_172,N_133,In_475);
or U173 (N_173,In_343,N_75);
nor U174 (N_174,In_201,N_91);
nor U175 (N_175,In_301,In_49);
and U176 (N_176,In_352,In_101);
or U177 (N_177,In_172,N_92);
nor U178 (N_178,In_477,In_218);
nand U179 (N_179,N_11,In_168);
nand U180 (N_180,N_1,N_79);
or U181 (N_181,In_208,In_363);
or U182 (N_182,N_67,N_93);
nor U183 (N_183,N_132,In_37);
nand U184 (N_184,In_249,In_214);
nor U185 (N_185,In_445,N_98);
nand U186 (N_186,In_222,In_23);
or U187 (N_187,In_16,In_464);
or U188 (N_188,N_6,N_24);
or U189 (N_189,In_458,N_90);
nand U190 (N_190,N_69,N_134);
and U191 (N_191,In_62,In_398);
and U192 (N_192,In_136,In_376);
and U193 (N_193,In_134,In_432);
nor U194 (N_194,In_426,In_372);
or U195 (N_195,N_123,N_13);
nor U196 (N_196,N_15,In_302);
or U197 (N_197,In_425,In_85);
nand U198 (N_198,N_68,In_72);
or U199 (N_199,In_370,In_334);
or U200 (N_200,N_107,N_53);
and U201 (N_201,In_180,In_268);
or U202 (N_202,In_206,In_243);
nor U203 (N_203,N_102,In_282);
nand U204 (N_204,In_38,N_138);
and U205 (N_205,In_113,N_172);
or U206 (N_206,N_151,N_163);
or U207 (N_207,In_290,In_19);
nand U208 (N_208,In_467,In_11);
and U209 (N_209,N_42,N_178);
nor U210 (N_210,In_176,N_55);
or U211 (N_211,In_96,In_305);
and U212 (N_212,In_211,In_280);
or U213 (N_213,N_170,N_32);
and U214 (N_214,In_95,In_489);
nand U215 (N_215,N_144,In_320);
nand U216 (N_216,N_9,In_325);
nand U217 (N_217,In_466,N_183);
and U218 (N_218,N_49,N_140);
or U219 (N_219,In_456,N_70);
or U220 (N_220,In_135,In_276);
or U221 (N_221,In_291,In_373);
nand U222 (N_222,N_148,N_72);
or U223 (N_223,In_192,In_423);
nor U224 (N_224,In_83,In_28);
nor U225 (N_225,In_151,In_216);
nand U226 (N_226,In_111,In_34);
nor U227 (N_227,N_136,N_10);
nand U228 (N_228,N_194,N_109);
and U229 (N_229,In_384,N_162);
nand U230 (N_230,N_113,N_62);
nor U231 (N_231,N_149,In_441);
or U232 (N_232,In_236,In_230);
and U233 (N_233,In_364,In_61);
nand U234 (N_234,In_80,N_186);
nand U235 (N_235,In_50,N_73);
or U236 (N_236,N_94,N_100);
nand U237 (N_237,In_333,N_166);
nor U238 (N_238,N_120,In_215);
or U239 (N_239,N_158,In_141);
nand U240 (N_240,In_43,In_444);
or U241 (N_241,In_14,In_314);
nor U242 (N_242,In_229,In_24);
or U243 (N_243,N_108,In_182);
or U244 (N_244,In_394,N_80);
or U245 (N_245,N_154,N_21);
nor U246 (N_246,In_46,In_307);
nor U247 (N_247,N_41,N_153);
and U248 (N_248,In_235,In_420);
or U249 (N_249,N_185,In_496);
nand U250 (N_250,N_33,N_236);
nor U251 (N_251,N_249,N_169);
nor U252 (N_252,N_177,N_54);
or U253 (N_253,N_234,In_367);
nor U254 (N_254,In_435,N_137);
nand U255 (N_255,N_143,N_106);
nand U256 (N_256,N_214,N_181);
nand U257 (N_257,N_159,In_203);
and U258 (N_258,In_152,N_146);
or U259 (N_259,In_129,N_65);
or U260 (N_260,N_77,In_122);
and U261 (N_261,In_204,N_165);
or U262 (N_262,In_91,N_224);
nand U263 (N_263,In_455,N_173);
nand U264 (N_264,N_200,N_226);
nor U265 (N_265,In_52,N_211);
nor U266 (N_266,In_160,N_205);
nand U267 (N_267,N_152,N_213);
or U268 (N_268,In_58,In_3);
or U269 (N_269,In_418,In_457);
nor U270 (N_270,N_201,N_8);
and U271 (N_271,In_199,N_118);
nand U272 (N_272,In_244,N_161);
or U273 (N_273,N_232,N_212);
and U274 (N_274,In_181,N_245);
nor U275 (N_275,N_167,N_190);
and U276 (N_276,N_124,In_99);
and U277 (N_277,In_137,In_164);
nor U278 (N_278,In_283,N_216);
or U279 (N_279,In_191,In_345);
nand U280 (N_280,N_182,N_51);
nand U281 (N_281,In_131,In_205);
and U282 (N_282,In_388,N_179);
nand U283 (N_283,N_225,N_203);
and U284 (N_284,N_175,N_191);
nor U285 (N_285,In_494,N_126);
and U286 (N_286,N_61,In_170);
nor U287 (N_287,N_202,N_204);
nand U288 (N_288,In_396,In_67);
nor U289 (N_289,In_415,N_114);
or U290 (N_290,In_51,In_442);
nand U291 (N_291,N_87,N_243);
or U292 (N_292,N_128,In_149);
or U293 (N_293,N_129,N_50);
nor U294 (N_294,N_231,In_118);
nor U295 (N_295,In_183,N_240);
or U296 (N_296,N_141,In_491);
or U297 (N_297,In_382,In_270);
and U298 (N_298,In_463,In_175);
nand U299 (N_299,In_21,In_422);
nor U300 (N_300,N_81,N_7);
or U301 (N_301,N_288,N_40);
nand U302 (N_302,In_495,N_168);
nor U303 (N_303,N_244,N_279);
or U304 (N_304,N_222,N_289);
or U305 (N_305,In_42,In_20);
or U306 (N_306,In_385,N_254);
and U307 (N_307,N_135,N_117);
and U308 (N_308,N_285,In_100);
nor U309 (N_309,N_267,In_428);
xnor U310 (N_310,In_424,N_258);
nor U311 (N_311,In_499,In_371);
and U312 (N_312,In_338,In_380);
nor U313 (N_313,In_121,N_276);
nor U314 (N_314,N_252,N_253);
and U315 (N_315,N_230,N_187);
xor U316 (N_316,N_291,In_250);
and U317 (N_317,In_6,In_124);
nor U318 (N_318,In_148,N_233);
nor U319 (N_319,In_300,N_237);
nand U320 (N_320,In_460,N_270);
or U321 (N_321,N_274,In_63);
and U322 (N_322,N_150,In_354);
and U323 (N_323,N_101,N_250);
nand U324 (N_324,N_268,In_36);
or U325 (N_325,N_156,N_155);
or U326 (N_326,N_235,In_412);
nor U327 (N_327,N_171,In_357);
nand U328 (N_328,N_228,In_234);
and U329 (N_329,N_121,N_260);
nor U330 (N_330,N_206,N_248);
nand U331 (N_331,In_125,N_119);
nand U332 (N_332,In_127,In_408);
or U333 (N_333,N_157,N_189);
nor U334 (N_334,N_256,N_130);
nor U335 (N_335,N_284,N_125);
or U336 (N_336,N_131,In_439);
and U337 (N_337,N_105,In_107);
nand U338 (N_338,In_213,N_265);
nor U339 (N_339,N_95,In_313);
nand U340 (N_340,N_197,N_227);
nand U341 (N_341,In_316,In_105);
nor U342 (N_342,N_239,N_275);
and U343 (N_343,N_198,N_273);
and U344 (N_344,In_221,In_417);
or U345 (N_345,In_315,N_111);
and U346 (N_346,N_195,N_84);
nor U347 (N_347,N_262,N_261);
and U348 (N_348,In_278,N_295);
nor U349 (N_349,In_68,In_341);
nand U350 (N_350,In_306,N_317);
or U351 (N_351,In_167,N_139);
and U352 (N_352,In_299,N_313);
and U353 (N_353,N_251,N_337);
nor U354 (N_354,N_266,N_286);
nand U355 (N_355,N_302,N_320);
nand U356 (N_356,N_34,In_429);
nand U357 (N_357,N_188,N_283);
and U358 (N_358,In_331,N_344);
nand U359 (N_359,N_349,N_184);
nor U360 (N_360,N_247,N_269);
or U361 (N_361,N_272,N_281);
nand U362 (N_362,N_255,N_348);
and U363 (N_363,N_304,In_451);
nor U364 (N_364,N_263,N_278);
nand U365 (N_365,N_343,N_328);
nor U366 (N_366,In_196,N_221);
or U367 (N_367,N_314,N_287);
and U368 (N_368,N_296,N_309);
and U369 (N_369,N_329,N_27);
or U370 (N_370,N_180,N_331);
nor U371 (N_371,N_104,In_431);
and U372 (N_372,N_23,N_297);
nor U373 (N_373,N_305,N_322);
and U374 (N_374,N_325,N_218);
and U375 (N_375,In_487,N_259);
or U376 (N_376,N_46,N_215);
nand U377 (N_377,N_312,N_246);
nor U378 (N_378,N_280,N_319);
and U379 (N_379,N_321,N_299);
or U380 (N_380,N_47,N_324);
nand U381 (N_381,N_271,N_292);
or U382 (N_382,N_199,N_64);
or U383 (N_383,N_229,In_360);
or U384 (N_384,N_310,In_312);
or U385 (N_385,N_315,N_127);
or U386 (N_386,N_311,N_160);
nand U387 (N_387,N_257,N_145);
nand U388 (N_388,In_378,N_238);
or U389 (N_389,N_210,N_341);
and U390 (N_390,In_330,N_192);
nor U391 (N_391,In_486,N_110);
and U392 (N_392,N_122,N_323);
xnor U393 (N_393,In_237,N_290);
and U394 (N_394,In_104,In_449);
or U395 (N_395,N_298,N_332);
and U396 (N_396,N_220,In_247);
nor U397 (N_397,In_490,N_264);
and U398 (N_398,N_316,N_342);
nand U399 (N_399,N_219,N_293);
or U400 (N_400,N_318,N_336);
nand U401 (N_401,N_300,N_294);
or U402 (N_402,N_372,N_366);
and U403 (N_403,N_380,N_303);
or U404 (N_404,N_17,N_398);
or U405 (N_405,N_346,N_306);
or U406 (N_406,N_207,N_381);
nor U407 (N_407,N_396,N_383);
nand U408 (N_408,N_371,N_385);
nand U409 (N_409,N_338,In_386);
nand U410 (N_410,N_142,N_378);
nor U411 (N_411,N_379,N_347);
nand U412 (N_412,N_388,N_356);
nand U413 (N_413,N_364,N_394);
nand U414 (N_414,N_363,N_196);
and U415 (N_415,N_368,N_375);
or U416 (N_416,N_365,N_241);
nor U417 (N_417,N_392,N_393);
nand U418 (N_418,N_60,N_355);
nor U419 (N_419,N_395,N_373);
nand U420 (N_420,N_208,N_370);
or U421 (N_421,N_301,In_197);
nand U422 (N_422,N_358,N_39);
nor U423 (N_423,In_295,N_326);
nand U424 (N_424,In_41,N_352);
or U425 (N_425,N_390,N_382);
nor U426 (N_426,N_242,In_327);
and U427 (N_427,N_330,N_327);
nor U428 (N_428,N_282,N_339);
or U429 (N_429,N_377,N_357);
nor U430 (N_430,N_308,N_354);
nand U431 (N_431,N_397,In_77);
nor U432 (N_432,N_193,N_335);
nor U433 (N_433,N_359,N_353);
or U434 (N_434,N_164,N_334);
and U435 (N_435,N_391,N_174);
or U436 (N_436,N_376,N_277);
or U437 (N_437,N_369,N_387);
or U438 (N_438,N_386,N_384);
nand U439 (N_439,N_389,N_399);
or U440 (N_440,N_345,N_367);
or U441 (N_441,N_340,N_223);
nor U442 (N_442,N_333,N_112);
and U443 (N_443,N_71,In_226);
nand U444 (N_444,N_374,N_351);
nand U445 (N_445,N_176,In_217);
or U446 (N_446,N_362,N_217);
nand U447 (N_447,N_361,N_350);
nand U448 (N_448,N_209,N_31);
or U449 (N_449,N_307,N_360);
and U450 (N_450,N_415,N_433);
nor U451 (N_451,N_404,N_423);
nand U452 (N_452,N_428,N_447);
nand U453 (N_453,N_444,N_448);
and U454 (N_454,N_430,N_412);
nand U455 (N_455,N_420,N_449);
nand U456 (N_456,N_413,N_418);
or U457 (N_457,N_419,N_407);
and U458 (N_458,N_431,N_446);
nor U459 (N_459,N_406,N_442);
and U460 (N_460,N_409,N_426);
and U461 (N_461,N_432,N_417);
or U462 (N_462,N_440,N_429);
or U463 (N_463,N_402,N_405);
or U464 (N_464,N_435,N_422);
nand U465 (N_465,N_403,N_414);
nor U466 (N_466,N_438,N_441);
xnor U467 (N_467,N_439,N_436);
nor U468 (N_468,N_424,N_434);
nand U469 (N_469,N_445,N_427);
and U470 (N_470,N_400,N_437);
nand U471 (N_471,N_411,N_408);
nand U472 (N_472,N_416,N_410);
or U473 (N_473,N_401,N_425);
nor U474 (N_474,N_443,N_421);
xnor U475 (N_475,N_430,N_432);
nor U476 (N_476,N_449,N_426);
or U477 (N_477,N_438,N_418);
xnor U478 (N_478,N_416,N_418);
nand U479 (N_479,N_411,N_404);
or U480 (N_480,N_404,N_426);
nand U481 (N_481,N_425,N_429);
nor U482 (N_482,N_406,N_413);
nor U483 (N_483,N_434,N_440);
nand U484 (N_484,N_445,N_410);
and U485 (N_485,N_449,N_416);
nand U486 (N_486,N_416,N_439);
nor U487 (N_487,N_420,N_442);
nor U488 (N_488,N_414,N_413);
or U489 (N_489,N_425,N_431);
nor U490 (N_490,N_420,N_417);
nand U491 (N_491,N_400,N_449);
or U492 (N_492,N_446,N_405);
and U493 (N_493,N_416,N_446);
nor U494 (N_494,N_447,N_430);
nor U495 (N_495,N_436,N_419);
nor U496 (N_496,N_419,N_426);
nor U497 (N_497,N_410,N_443);
or U498 (N_498,N_424,N_421);
or U499 (N_499,N_411,N_429);
or U500 (N_500,N_456,N_450);
or U501 (N_501,N_466,N_498);
xnor U502 (N_502,N_487,N_478);
nor U503 (N_503,N_464,N_495);
and U504 (N_504,N_472,N_480);
nand U505 (N_505,N_455,N_485);
and U506 (N_506,N_467,N_493);
nand U507 (N_507,N_463,N_490);
nor U508 (N_508,N_489,N_494);
nor U509 (N_509,N_470,N_479);
and U510 (N_510,N_454,N_452);
nand U511 (N_511,N_484,N_462);
or U512 (N_512,N_457,N_492);
or U513 (N_513,N_499,N_453);
and U514 (N_514,N_461,N_491);
nand U515 (N_515,N_486,N_483);
nand U516 (N_516,N_476,N_488);
nor U517 (N_517,N_473,N_451);
or U518 (N_518,N_458,N_477);
and U519 (N_519,N_497,N_469);
or U520 (N_520,N_496,N_465);
nand U521 (N_521,N_459,N_481);
nor U522 (N_522,N_474,N_460);
or U523 (N_523,N_468,N_475);
xnor U524 (N_524,N_482,N_471);
nor U525 (N_525,N_470,N_474);
nor U526 (N_526,N_463,N_465);
or U527 (N_527,N_459,N_480);
nand U528 (N_528,N_499,N_451);
or U529 (N_529,N_496,N_468);
or U530 (N_530,N_495,N_493);
or U531 (N_531,N_467,N_466);
or U532 (N_532,N_459,N_488);
nor U533 (N_533,N_492,N_498);
nand U534 (N_534,N_452,N_473);
nand U535 (N_535,N_497,N_462);
nor U536 (N_536,N_459,N_471);
nand U537 (N_537,N_491,N_492);
and U538 (N_538,N_482,N_472);
nand U539 (N_539,N_479,N_485);
or U540 (N_540,N_451,N_456);
xnor U541 (N_541,N_468,N_493);
nor U542 (N_542,N_474,N_479);
nand U543 (N_543,N_465,N_486);
and U544 (N_544,N_490,N_497);
nand U545 (N_545,N_491,N_453);
and U546 (N_546,N_486,N_478);
and U547 (N_547,N_469,N_493);
nor U548 (N_548,N_451,N_491);
nand U549 (N_549,N_463,N_487);
nor U550 (N_550,N_514,N_506);
nor U551 (N_551,N_510,N_521);
or U552 (N_552,N_526,N_525);
and U553 (N_553,N_511,N_516);
nor U554 (N_554,N_528,N_549);
or U555 (N_555,N_503,N_501);
nand U556 (N_556,N_515,N_534);
and U557 (N_557,N_542,N_513);
and U558 (N_558,N_547,N_519);
nor U559 (N_559,N_504,N_500);
and U560 (N_560,N_530,N_502);
nor U561 (N_561,N_533,N_527);
nand U562 (N_562,N_531,N_548);
or U563 (N_563,N_537,N_520);
nand U564 (N_564,N_517,N_512);
and U565 (N_565,N_536,N_529);
nand U566 (N_566,N_532,N_543);
or U567 (N_567,N_522,N_507);
nand U568 (N_568,N_540,N_524);
or U569 (N_569,N_539,N_523);
and U570 (N_570,N_538,N_546);
xnor U571 (N_571,N_518,N_509);
nor U572 (N_572,N_541,N_544);
and U573 (N_573,N_535,N_505);
or U574 (N_574,N_508,N_545);
and U575 (N_575,N_521,N_517);
nand U576 (N_576,N_500,N_532);
nand U577 (N_577,N_524,N_545);
or U578 (N_578,N_516,N_521);
nor U579 (N_579,N_548,N_515);
nor U580 (N_580,N_545,N_519);
or U581 (N_581,N_542,N_539);
and U582 (N_582,N_544,N_508);
or U583 (N_583,N_521,N_523);
and U584 (N_584,N_533,N_510);
nand U585 (N_585,N_540,N_506);
nand U586 (N_586,N_549,N_534);
or U587 (N_587,N_528,N_504);
or U588 (N_588,N_505,N_524);
nand U589 (N_589,N_538,N_511);
nor U590 (N_590,N_544,N_519);
nand U591 (N_591,N_520,N_529);
or U592 (N_592,N_522,N_535);
and U593 (N_593,N_539,N_533);
nand U594 (N_594,N_517,N_502);
or U595 (N_595,N_504,N_523);
and U596 (N_596,N_542,N_526);
nand U597 (N_597,N_516,N_515);
nor U598 (N_598,N_523,N_529);
nand U599 (N_599,N_546,N_525);
or U600 (N_600,N_559,N_595);
or U601 (N_601,N_556,N_578);
nand U602 (N_602,N_561,N_572);
nor U603 (N_603,N_558,N_593);
nand U604 (N_604,N_568,N_550);
or U605 (N_605,N_557,N_562);
or U606 (N_606,N_570,N_554);
nor U607 (N_607,N_571,N_589);
and U608 (N_608,N_591,N_575);
nand U609 (N_609,N_574,N_553);
and U610 (N_610,N_599,N_567);
nor U611 (N_611,N_566,N_586);
or U612 (N_612,N_563,N_598);
or U613 (N_613,N_577,N_597);
and U614 (N_614,N_596,N_594);
or U615 (N_615,N_592,N_581);
xnor U616 (N_616,N_560,N_580);
or U617 (N_617,N_584,N_555);
or U618 (N_618,N_576,N_573);
nand U619 (N_619,N_551,N_588);
nor U620 (N_620,N_552,N_579);
or U621 (N_621,N_565,N_582);
or U622 (N_622,N_583,N_587);
or U623 (N_623,N_569,N_590);
or U624 (N_624,N_564,N_585);
or U625 (N_625,N_555,N_575);
nor U626 (N_626,N_583,N_593);
and U627 (N_627,N_569,N_595);
or U628 (N_628,N_573,N_593);
nor U629 (N_629,N_591,N_574);
or U630 (N_630,N_560,N_554);
nor U631 (N_631,N_566,N_579);
nor U632 (N_632,N_579,N_597);
nor U633 (N_633,N_569,N_560);
or U634 (N_634,N_596,N_554);
nor U635 (N_635,N_591,N_585);
nand U636 (N_636,N_559,N_570);
xnor U637 (N_637,N_597,N_559);
nor U638 (N_638,N_556,N_553);
or U639 (N_639,N_582,N_561);
and U640 (N_640,N_565,N_568);
nand U641 (N_641,N_594,N_595);
or U642 (N_642,N_563,N_552);
nand U643 (N_643,N_590,N_578);
nand U644 (N_644,N_599,N_565);
nor U645 (N_645,N_568,N_596);
and U646 (N_646,N_576,N_581);
and U647 (N_647,N_597,N_565);
or U648 (N_648,N_583,N_577);
or U649 (N_649,N_557,N_553);
nor U650 (N_650,N_636,N_621);
or U651 (N_651,N_633,N_629);
nor U652 (N_652,N_622,N_641);
and U653 (N_653,N_604,N_628);
or U654 (N_654,N_634,N_600);
and U655 (N_655,N_625,N_619);
nor U656 (N_656,N_608,N_623);
and U657 (N_657,N_602,N_632);
nand U658 (N_658,N_644,N_649);
nor U659 (N_659,N_630,N_635);
or U660 (N_660,N_614,N_612);
nand U661 (N_661,N_603,N_631);
and U662 (N_662,N_638,N_643);
or U663 (N_663,N_646,N_637);
nand U664 (N_664,N_607,N_647);
nand U665 (N_665,N_626,N_606);
and U666 (N_666,N_645,N_617);
xnor U667 (N_667,N_609,N_642);
nor U668 (N_668,N_648,N_610);
nand U669 (N_669,N_601,N_640);
and U670 (N_670,N_620,N_639);
and U671 (N_671,N_616,N_627);
nand U672 (N_672,N_613,N_624);
and U673 (N_673,N_605,N_615);
nand U674 (N_674,N_611,N_618);
nor U675 (N_675,N_625,N_646);
and U676 (N_676,N_623,N_648);
nor U677 (N_677,N_642,N_634);
nor U678 (N_678,N_623,N_626);
nand U679 (N_679,N_601,N_638);
and U680 (N_680,N_614,N_608);
nor U681 (N_681,N_643,N_603);
and U682 (N_682,N_647,N_626);
nor U683 (N_683,N_605,N_611);
and U684 (N_684,N_631,N_643);
nor U685 (N_685,N_604,N_646);
nand U686 (N_686,N_645,N_625);
or U687 (N_687,N_633,N_607);
or U688 (N_688,N_604,N_619);
nor U689 (N_689,N_643,N_621);
and U690 (N_690,N_601,N_602);
nor U691 (N_691,N_616,N_604);
nand U692 (N_692,N_605,N_603);
nor U693 (N_693,N_630,N_610);
and U694 (N_694,N_642,N_616);
nand U695 (N_695,N_601,N_643);
or U696 (N_696,N_611,N_610);
nor U697 (N_697,N_600,N_648);
and U698 (N_698,N_630,N_608);
nand U699 (N_699,N_647,N_643);
nor U700 (N_700,N_697,N_650);
and U701 (N_701,N_680,N_665);
nor U702 (N_702,N_684,N_692);
or U703 (N_703,N_690,N_667);
nand U704 (N_704,N_666,N_661);
or U705 (N_705,N_672,N_674);
nor U706 (N_706,N_691,N_657);
or U707 (N_707,N_696,N_699);
or U708 (N_708,N_695,N_686);
nand U709 (N_709,N_659,N_651);
and U710 (N_710,N_658,N_656);
nand U711 (N_711,N_678,N_687);
nand U712 (N_712,N_675,N_670);
nand U713 (N_713,N_698,N_683);
and U714 (N_714,N_669,N_654);
nor U715 (N_715,N_671,N_685);
and U716 (N_716,N_660,N_682);
nand U717 (N_717,N_652,N_676);
nand U718 (N_718,N_662,N_688);
or U719 (N_719,N_689,N_653);
and U720 (N_720,N_663,N_664);
and U721 (N_721,N_668,N_694);
and U722 (N_722,N_679,N_693);
or U723 (N_723,N_677,N_673);
nand U724 (N_724,N_655,N_681);
nand U725 (N_725,N_691,N_698);
or U726 (N_726,N_675,N_681);
nand U727 (N_727,N_675,N_662);
nor U728 (N_728,N_683,N_690);
nor U729 (N_729,N_659,N_690);
nor U730 (N_730,N_679,N_658);
and U731 (N_731,N_685,N_662);
nor U732 (N_732,N_685,N_683);
and U733 (N_733,N_660,N_695);
nand U734 (N_734,N_690,N_658);
nand U735 (N_735,N_699,N_662);
nor U736 (N_736,N_672,N_664);
nor U737 (N_737,N_669,N_665);
and U738 (N_738,N_677,N_665);
or U739 (N_739,N_677,N_693);
or U740 (N_740,N_681,N_653);
or U741 (N_741,N_687,N_691);
and U742 (N_742,N_680,N_658);
and U743 (N_743,N_673,N_657);
or U744 (N_744,N_681,N_661);
or U745 (N_745,N_670,N_674);
nor U746 (N_746,N_666,N_692);
nor U747 (N_747,N_692,N_690);
nor U748 (N_748,N_683,N_676);
xor U749 (N_749,N_655,N_660);
and U750 (N_750,N_718,N_741);
nor U751 (N_751,N_740,N_749);
or U752 (N_752,N_711,N_728);
and U753 (N_753,N_737,N_705);
and U754 (N_754,N_742,N_730);
nor U755 (N_755,N_726,N_729);
nand U756 (N_756,N_747,N_745);
nor U757 (N_757,N_738,N_707);
and U758 (N_758,N_704,N_724);
and U759 (N_759,N_735,N_709);
nor U760 (N_760,N_708,N_715);
and U761 (N_761,N_720,N_702);
and U762 (N_762,N_744,N_731);
or U763 (N_763,N_714,N_721);
nor U764 (N_764,N_748,N_716);
and U765 (N_765,N_706,N_712);
or U766 (N_766,N_746,N_736);
and U767 (N_767,N_701,N_710);
nor U768 (N_768,N_717,N_722);
nor U769 (N_769,N_743,N_732);
nand U770 (N_770,N_739,N_725);
or U771 (N_771,N_719,N_727);
nand U772 (N_772,N_700,N_733);
and U773 (N_773,N_713,N_703);
nor U774 (N_774,N_734,N_723);
nor U775 (N_775,N_705,N_704);
and U776 (N_776,N_743,N_706);
or U777 (N_777,N_747,N_705);
and U778 (N_778,N_720,N_709);
or U779 (N_779,N_721,N_748);
or U780 (N_780,N_731,N_748);
or U781 (N_781,N_736,N_730);
and U782 (N_782,N_745,N_727);
nand U783 (N_783,N_702,N_708);
nand U784 (N_784,N_742,N_706);
or U785 (N_785,N_719,N_748);
or U786 (N_786,N_727,N_734);
or U787 (N_787,N_708,N_733);
nor U788 (N_788,N_724,N_707);
nor U789 (N_789,N_740,N_743);
and U790 (N_790,N_727,N_723);
or U791 (N_791,N_707,N_722);
nor U792 (N_792,N_726,N_744);
or U793 (N_793,N_730,N_743);
nand U794 (N_794,N_702,N_725);
and U795 (N_795,N_735,N_706);
or U796 (N_796,N_718,N_706);
nor U797 (N_797,N_747,N_720);
nor U798 (N_798,N_711,N_735);
nor U799 (N_799,N_714,N_716);
nand U800 (N_800,N_763,N_785);
and U801 (N_801,N_787,N_754);
and U802 (N_802,N_768,N_798);
and U803 (N_803,N_799,N_751);
and U804 (N_804,N_784,N_794);
or U805 (N_805,N_792,N_790);
or U806 (N_806,N_752,N_791);
and U807 (N_807,N_789,N_786);
nor U808 (N_808,N_776,N_758);
or U809 (N_809,N_760,N_773);
or U810 (N_810,N_780,N_782);
nor U811 (N_811,N_769,N_777);
and U812 (N_812,N_774,N_750);
or U813 (N_813,N_764,N_771);
and U814 (N_814,N_788,N_781);
or U815 (N_815,N_761,N_767);
nand U816 (N_816,N_783,N_759);
nand U817 (N_817,N_775,N_779);
nor U818 (N_818,N_765,N_756);
and U819 (N_819,N_793,N_797);
nor U820 (N_820,N_778,N_770);
nor U821 (N_821,N_753,N_755);
and U822 (N_822,N_757,N_796);
nand U823 (N_823,N_772,N_762);
nor U824 (N_824,N_766,N_795);
nor U825 (N_825,N_785,N_776);
nand U826 (N_826,N_774,N_778);
nor U827 (N_827,N_781,N_785);
and U828 (N_828,N_759,N_795);
nand U829 (N_829,N_787,N_777);
and U830 (N_830,N_787,N_752);
or U831 (N_831,N_752,N_766);
and U832 (N_832,N_761,N_756);
nor U833 (N_833,N_767,N_799);
or U834 (N_834,N_794,N_771);
nand U835 (N_835,N_767,N_768);
nand U836 (N_836,N_757,N_783);
or U837 (N_837,N_752,N_761);
and U838 (N_838,N_770,N_774);
nor U839 (N_839,N_783,N_772);
and U840 (N_840,N_768,N_775);
nand U841 (N_841,N_761,N_782);
nand U842 (N_842,N_782,N_756);
nor U843 (N_843,N_760,N_774);
and U844 (N_844,N_799,N_769);
and U845 (N_845,N_756,N_785);
nand U846 (N_846,N_765,N_758);
nand U847 (N_847,N_761,N_798);
or U848 (N_848,N_786,N_750);
or U849 (N_849,N_785,N_798);
nand U850 (N_850,N_819,N_834);
nor U851 (N_851,N_806,N_838);
nor U852 (N_852,N_811,N_845);
nand U853 (N_853,N_825,N_849);
nor U854 (N_854,N_821,N_808);
nand U855 (N_855,N_813,N_815);
and U856 (N_856,N_812,N_805);
or U857 (N_857,N_810,N_827);
and U858 (N_858,N_848,N_828);
nor U859 (N_859,N_842,N_823);
and U860 (N_860,N_822,N_837);
nor U861 (N_861,N_820,N_809);
or U862 (N_862,N_831,N_818);
nand U863 (N_863,N_817,N_802);
xor U864 (N_864,N_800,N_844);
or U865 (N_865,N_839,N_841);
and U866 (N_866,N_830,N_835);
nand U867 (N_867,N_801,N_833);
nand U868 (N_868,N_824,N_843);
nand U869 (N_869,N_804,N_847);
nand U870 (N_870,N_807,N_816);
nand U871 (N_871,N_814,N_826);
nor U872 (N_872,N_832,N_840);
nand U873 (N_873,N_803,N_846);
nor U874 (N_874,N_836,N_829);
nor U875 (N_875,N_815,N_806);
or U876 (N_876,N_833,N_824);
or U877 (N_877,N_845,N_821);
nand U878 (N_878,N_801,N_826);
nand U879 (N_879,N_846,N_844);
nand U880 (N_880,N_819,N_811);
and U881 (N_881,N_829,N_818);
or U882 (N_882,N_811,N_805);
nand U883 (N_883,N_821,N_830);
nor U884 (N_884,N_836,N_841);
xnor U885 (N_885,N_809,N_825);
xnor U886 (N_886,N_828,N_835);
and U887 (N_887,N_832,N_844);
nor U888 (N_888,N_829,N_803);
and U889 (N_889,N_813,N_843);
or U890 (N_890,N_846,N_845);
and U891 (N_891,N_840,N_810);
nor U892 (N_892,N_839,N_800);
or U893 (N_893,N_818,N_819);
nor U894 (N_894,N_835,N_818);
or U895 (N_895,N_825,N_814);
nor U896 (N_896,N_800,N_835);
nand U897 (N_897,N_844,N_843);
and U898 (N_898,N_812,N_825);
nand U899 (N_899,N_848,N_809);
and U900 (N_900,N_866,N_886);
nor U901 (N_901,N_898,N_862);
and U902 (N_902,N_859,N_881);
and U903 (N_903,N_863,N_858);
nand U904 (N_904,N_891,N_880);
nand U905 (N_905,N_875,N_874);
and U906 (N_906,N_860,N_851);
and U907 (N_907,N_854,N_868);
and U908 (N_908,N_895,N_883);
nor U909 (N_909,N_873,N_857);
nand U910 (N_910,N_894,N_877);
nor U911 (N_911,N_872,N_871);
xnor U912 (N_912,N_888,N_852);
or U913 (N_913,N_896,N_887);
or U914 (N_914,N_869,N_889);
and U915 (N_915,N_884,N_897);
and U916 (N_916,N_882,N_899);
and U917 (N_917,N_892,N_855);
xnor U918 (N_918,N_878,N_870);
and U919 (N_919,N_879,N_867);
and U920 (N_920,N_850,N_853);
and U921 (N_921,N_893,N_861);
nand U922 (N_922,N_876,N_865);
nand U923 (N_923,N_890,N_856);
or U924 (N_924,N_864,N_885);
or U925 (N_925,N_881,N_868);
nor U926 (N_926,N_852,N_866);
and U927 (N_927,N_871,N_887);
or U928 (N_928,N_881,N_861);
nand U929 (N_929,N_878,N_886);
nor U930 (N_930,N_897,N_853);
or U931 (N_931,N_866,N_875);
and U932 (N_932,N_897,N_888);
and U933 (N_933,N_878,N_877);
nand U934 (N_934,N_881,N_856);
nor U935 (N_935,N_855,N_862);
nor U936 (N_936,N_890,N_867);
nand U937 (N_937,N_892,N_885);
nor U938 (N_938,N_882,N_870);
and U939 (N_939,N_893,N_863);
and U940 (N_940,N_878,N_894);
nor U941 (N_941,N_854,N_885);
and U942 (N_942,N_856,N_886);
nand U943 (N_943,N_874,N_861);
and U944 (N_944,N_862,N_887);
or U945 (N_945,N_894,N_898);
xor U946 (N_946,N_891,N_889);
nor U947 (N_947,N_896,N_893);
nand U948 (N_948,N_891,N_859);
nor U949 (N_949,N_870,N_883);
or U950 (N_950,N_935,N_929);
or U951 (N_951,N_949,N_936);
nand U952 (N_952,N_919,N_925);
or U953 (N_953,N_933,N_903);
nand U954 (N_954,N_900,N_911);
nor U955 (N_955,N_934,N_904);
nand U956 (N_956,N_923,N_901);
nor U957 (N_957,N_913,N_939);
nand U958 (N_958,N_942,N_947);
and U959 (N_959,N_905,N_938);
nor U960 (N_960,N_926,N_948);
and U961 (N_961,N_924,N_937);
or U962 (N_962,N_920,N_902);
and U963 (N_963,N_917,N_943);
or U964 (N_964,N_912,N_910);
and U965 (N_965,N_914,N_916);
or U966 (N_966,N_907,N_918);
or U967 (N_967,N_908,N_944);
nor U968 (N_968,N_932,N_909);
and U969 (N_969,N_921,N_906);
or U970 (N_970,N_931,N_915);
nand U971 (N_971,N_946,N_930);
and U972 (N_972,N_940,N_927);
nor U973 (N_973,N_928,N_945);
nor U974 (N_974,N_922,N_941);
and U975 (N_975,N_934,N_903);
or U976 (N_976,N_945,N_902);
or U977 (N_977,N_915,N_923);
and U978 (N_978,N_937,N_901);
or U979 (N_979,N_904,N_940);
and U980 (N_980,N_933,N_946);
and U981 (N_981,N_902,N_934);
or U982 (N_982,N_935,N_947);
or U983 (N_983,N_944,N_914);
or U984 (N_984,N_919,N_922);
or U985 (N_985,N_941,N_910);
nand U986 (N_986,N_943,N_927);
nand U987 (N_987,N_926,N_912);
nand U988 (N_988,N_924,N_932);
nand U989 (N_989,N_935,N_911);
or U990 (N_990,N_924,N_914);
and U991 (N_991,N_908,N_936);
xnor U992 (N_992,N_914,N_908);
and U993 (N_993,N_914,N_923);
nor U994 (N_994,N_935,N_902);
or U995 (N_995,N_936,N_922);
nor U996 (N_996,N_942,N_933);
or U997 (N_997,N_929,N_902);
and U998 (N_998,N_940,N_912);
and U999 (N_999,N_909,N_906);
nand U1000 (N_1000,N_976,N_974);
nand U1001 (N_1001,N_952,N_961);
and U1002 (N_1002,N_950,N_989);
or U1003 (N_1003,N_981,N_957);
nand U1004 (N_1004,N_954,N_984);
and U1005 (N_1005,N_994,N_958);
and U1006 (N_1006,N_959,N_970);
nand U1007 (N_1007,N_960,N_973);
nand U1008 (N_1008,N_953,N_993);
nand U1009 (N_1009,N_999,N_986);
nand U1010 (N_1010,N_971,N_998);
nand U1011 (N_1011,N_985,N_968);
and U1012 (N_1012,N_996,N_990);
nor U1013 (N_1013,N_967,N_982);
and U1014 (N_1014,N_956,N_997);
or U1015 (N_1015,N_980,N_978);
nor U1016 (N_1016,N_951,N_995);
and U1017 (N_1017,N_992,N_979);
or U1018 (N_1018,N_955,N_988);
and U1019 (N_1019,N_983,N_987);
nand U1020 (N_1020,N_972,N_962);
nand U1021 (N_1021,N_969,N_965);
xnor U1022 (N_1022,N_977,N_966);
or U1023 (N_1023,N_991,N_975);
xor U1024 (N_1024,N_963,N_964);
or U1025 (N_1025,N_971,N_997);
or U1026 (N_1026,N_982,N_996);
or U1027 (N_1027,N_963,N_957);
xnor U1028 (N_1028,N_995,N_964);
nor U1029 (N_1029,N_961,N_990);
or U1030 (N_1030,N_981,N_960);
nor U1031 (N_1031,N_951,N_983);
and U1032 (N_1032,N_999,N_968);
nand U1033 (N_1033,N_984,N_972);
nand U1034 (N_1034,N_957,N_951);
nor U1035 (N_1035,N_990,N_954);
and U1036 (N_1036,N_986,N_976);
nand U1037 (N_1037,N_951,N_986);
or U1038 (N_1038,N_966,N_983);
nor U1039 (N_1039,N_973,N_987);
and U1040 (N_1040,N_950,N_952);
nand U1041 (N_1041,N_995,N_991);
nor U1042 (N_1042,N_958,N_999);
and U1043 (N_1043,N_986,N_997);
nand U1044 (N_1044,N_962,N_991);
and U1045 (N_1045,N_997,N_989);
nor U1046 (N_1046,N_965,N_994);
nand U1047 (N_1047,N_971,N_992);
or U1048 (N_1048,N_970,N_993);
nand U1049 (N_1049,N_955,N_963);
nand U1050 (N_1050,N_1047,N_1039);
nand U1051 (N_1051,N_1020,N_1033);
nor U1052 (N_1052,N_1018,N_1011);
or U1053 (N_1053,N_1005,N_1001);
nand U1054 (N_1054,N_1028,N_1035);
nor U1055 (N_1055,N_1037,N_1013);
nor U1056 (N_1056,N_1032,N_1036);
and U1057 (N_1057,N_1010,N_1030);
or U1058 (N_1058,N_1038,N_1041);
nand U1059 (N_1059,N_1017,N_1024);
nor U1060 (N_1060,N_1019,N_1016);
nor U1061 (N_1061,N_1023,N_1003);
nand U1062 (N_1062,N_1021,N_1007);
nor U1063 (N_1063,N_1009,N_1025);
nor U1064 (N_1064,N_1014,N_1004);
or U1065 (N_1065,N_1049,N_1048);
nand U1066 (N_1066,N_1043,N_1027);
nor U1067 (N_1067,N_1008,N_1042);
and U1068 (N_1068,N_1000,N_1040);
and U1069 (N_1069,N_1026,N_1046);
and U1070 (N_1070,N_1045,N_1002);
and U1071 (N_1071,N_1015,N_1012);
or U1072 (N_1072,N_1031,N_1044);
nand U1073 (N_1073,N_1006,N_1022);
or U1074 (N_1074,N_1034,N_1029);
or U1075 (N_1075,N_1016,N_1018);
or U1076 (N_1076,N_1030,N_1000);
nor U1077 (N_1077,N_1017,N_1032);
nor U1078 (N_1078,N_1033,N_1035);
and U1079 (N_1079,N_1022,N_1037);
or U1080 (N_1080,N_1027,N_1007);
nand U1081 (N_1081,N_1033,N_1041);
and U1082 (N_1082,N_1004,N_1047);
or U1083 (N_1083,N_1048,N_1006);
or U1084 (N_1084,N_1043,N_1012);
or U1085 (N_1085,N_1031,N_1008);
nor U1086 (N_1086,N_1041,N_1046);
nor U1087 (N_1087,N_1046,N_1018);
nor U1088 (N_1088,N_1040,N_1034);
and U1089 (N_1089,N_1037,N_1010);
nand U1090 (N_1090,N_1034,N_1030);
nor U1091 (N_1091,N_1043,N_1009);
nor U1092 (N_1092,N_1037,N_1034);
nor U1093 (N_1093,N_1008,N_1017);
and U1094 (N_1094,N_1004,N_1028);
and U1095 (N_1095,N_1023,N_1042);
and U1096 (N_1096,N_1034,N_1023);
or U1097 (N_1097,N_1005,N_1048);
nand U1098 (N_1098,N_1034,N_1036);
nand U1099 (N_1099,N_1012,N_1007);
or U1100 (N_1100,N_1068,N_1078);
nor U1101 (N_1101,N_1054,N_1095);
nand U1102 (N_1102,N_1088,N_1092);
and U1103 (N_1103,N_1062,N_1067);
nand U1104 (N_1104,N_1069,N_1063);
and U1105 (N_1105,N_1072,N_1082);
or U1106 (N_1106,N_1096,N_1065);
or U1107 (N_1107,N_1080,N_1098);
or U1108 (N_1108,N_1089,N_1050);
nor U1109 (N_1109,N_1077,N_1053);
xnor U1110 (N_1110,N_1057,N_1093);
or U1111 (N_1111,N_1060,N_1079);
or U1112 (N_1112,N_1055,N_1076);
nand U1113 (N_1113,N_1097,N_1083);
nor U1114 (N_1114,N_1051,N_1073);
and U1115 (N_1115,N_1084,N_1059);
or U1116 (N_1116,N_1061,N_1074);
or U1117 (N_1117,N_1075,N_1070);
and U1118 (N_1118,N_1087,N_1085);
and U1119 (N_1119,N_1090,N_1086);
or U1120 (N_1120,N_1064,N_1091);
or U1121 (N_1121,N_1081,N_1094);
or U1122 (N_1122,N_1056,N_1099);
or U1123 (N_1123,N_1052,N_1071);
nand U1124 (N_1124,N_1058,N_1066);
nand U1125 (N_1125,N_1056,N_1074);
or U1126 (N_1126,N_1071,N_1055);
nor U1127 (N_1127,N_1069,N_1074);
or U1128 (N_1128,N_1075,N_1067);
and U1129 (N_1129,N_1072,N_1050);
nor U1130 (N_1130,N_1058,N_1090);
nor U1131 (N_1131,N_1078,N_1058);
nand U1132 (N_1132,N_1082,N_1056);
and U1133 (N_1133,N_1066,N_1087);
or U1134 (N_1134,N_1090,N_1056);
and U1135 (N_1135,N_1077,N_1078);
nand U1136 (N_1136,N_1081,N_1098);
nor U1137 (N_1137,N_1089,N_1059);
nand U1138 (N_1138,N_1052,N_1067);
and U1139 (N_1139,N_1088,N_1079);
nand U1140 (N_1140,N_1077,N_1076);
nand U1141 (N_1141,N_1087,N_1056);
or U1142 (N_1142,N_1092,N_1065);
and U1143 (N_1143,N_1054,N_1052);
or U1144 (N_1144,N_1099,N_1074);
nor U1145 (N_1145,N_1086,N_1053);
nor U1146 (N_1146,N_1097,N_1089);
or U1147 (N_1147,N_1057,N_1069);
and U1148 (N_1148,N_1056,N_1067);
or U1149 (N_1149,N_1065,N_1061);
nor U1150 (N_1150,N_1137,N_1104);
nand U1151 (N_1151,N_1116,N_1107);
nor U1152 (N_1152,N_1112,N_1133);
and U1153 (N_1153,N_1127,N_1139);
nand U1154 (N_1154,N_1134,N_1145);
and U1155 (N_1155,N_1126,N_1132);
and U1156 (N_1156,N_1108,N_1122);
nand U1157 (N_1157,N_1109,N_1100);
xor U1158 (N_1158,N_1118,N_1114);
nor U1159 (N_1159,N_1119,N_1136);
nor U1160 (N_1160,N_1140,N_1121);
and U1161 (N_1161,N_1141,N_1124);
nor U1162 (N_1162,N_1117,N_1147);
and U1163 (N_1163,N_1105,N_1125);
and U1164 (N_1164,N_1143,N_1130);
nand U1165 (N_1165,N_1128,N_1120);
nor U1166 (N_1166,N_1106,N_1149);
nor U1167 (N_1167,N_1148,N_1144);
nand U1168 (N_1168,N_1129,N_1135);
or U1169 (N_1169,N_1142,N_1146);
or U1170 (N_1170,N_1113,N_1103);
and U1171 (N_1171,N_1101,N_1131);
or U1172 (N_1172,N_1102,N_1111);
or U1173 (N_1173,N_1123,N_1110);
or U1174 (N_1174,N_1115,N_1138);
or U1175 (N_1175,N_1128,N_1112);
or U1176 (N_1176,N_1106,N_1131);
or U1177 (N_1177,N_1124,N_1132);
and U1178 (N_1178,N_1100,N_1128);
nand U1179 (N_1179,N_1147,N_1136);
nand U1180 (N_1180,N_1107,N_1130);
nor U1181 (N_1181,N_1106,N_1113);
nor U1182 (N_1182,N_1109,N_1123);
and U1183 (N_1183,N_1103,N_1143);
nand U1184 (N_1184,N_1114,N_1117);
nor U1185 (N_1185,N_1105,N_1127);
and U1186 (N_1186,N_1139,N_1144);
or U1187 (N_1187,N_1138,N_1123);
nor U1188 (N_1188,N_1147,N_1134);
xor U1189 (N_1189,N_1118,N_1135);
nor U1190 (N_1190,N_1120,N_1122);
nand U1191 (N_1191,N_1135,N_1115);
or U1192 (N_1192,N_1121,N_1105);
nand U1193 (N_1193,N_1106,N_1123);
nor U1194 (N_1194,N_1123,N_1139);
xor U1195 (N_1195,N_1129,N_1123);
and U1196 (N_1196,N_1140,N_1106);
xor U1197 (N_1197,N_1120,N_1123);
and U1198 (N_1198,N_1107,N_1105);
xor U1199 (N_1199,N_1124,N_1108);
nor U1200 (N_1200,N_1158,N_1150);
and U1201 (N_1201,N_1198,N_1160);
or U1202 (N_1202,N_1166,N_1168);
and U1203 (N_1203,N_1182,N_1188);
or U1204 (N_1204,N_1162,N_1192);
and U1205 (N_1205,N_1153,N_1187);
and U1206 (N_1206,N_1181,N_1199);
nand U1207 (N_1207,N_1156,N_1195);
or U1208 (N_1208,N_1193,N_1157);
and U1209 (N_1209,N_1167,N_1183);
and U1210 (N_1210,N_1155,N_1184);
and U1211 (N_1211,N_1177,N_1175);
nor U1212 (N_1212,N_1194,N_1185);
or U1213 (N_1213,N_1159,N_1176);
nor U1214 (N_1214,N_1171,N_1196);
or U1215 (N_1215,N_1178,N_1172);
nand U1216 (N_1216,N_1152,N_1191);
nand U1217 (N_1217,N_1151,N_1169);
or U1218 (N_1218,N_1161,N_1164);
nand U1219 (N_1219,N_1190,N_1189);
and U1220 (N_1220,N_1154,N_1186);
nor U1221 (N_1221,N_1173,N_1180);
nor U1222 (N_1222,N_1163,N_1170);
nor U1223 (N_1223,N_1174,N_1165);
nand U1224 (N_1224,N_1179,N_1197);
nor U1225 (N_1225,N_1175,N_1161);
nand U1226 (N_1226,N_1167,N_1171);
or U1227 (N_1227,N_1190,N_1181);
nand U1228 (N_1228,N_1190,N_1162);
nand U1229 (N_1229,N_1168,N_1178);
or U1230 (N_1230,N_1170,N_1174);
nor U1231 (N_1231,N_1162,N_1163);
or U1232 (N_1232,N_1198,N_1168);
nand U1233 (N_1233,N_1195,N_1184);
nand U1234 (N_1234,N_1151,N_1161);
and U1235 (N_1235,N_1193,N_1195);
and U1236 (N_1236,N_1177,N_1176);
xor U1237 (N_1237,N_1166,N_1197);
or U1238 (N_1238,N_1151,N_1177);
nand U1239 (N_1239,N_1151,N_1173);
and U1240 (N_1240,N_1150,N_1195);
nor U1241 (N_1241,N_1156,N_1175);
nor U1242 (N_1242,N_1192,N_1169);
and U1243 (N_1243,N_1185,N_1186);
xor U1244 (N_1244,N_1158,N_1171);
nand U1245 (N_1245,N_1178,N_1182);
and U1246 (N_1246,N_1170,N_1150);
nor U1247 (N_1247,N_1195,N_1177);
nor U1248 (N_1248,N_1187,N_1188);
nand U1249 (N_1249,N_1187,N_1164);
and U1250 (N_1250,N_1210,N_1222);
and U1251 (N_1251,N_1204,N_1206);
nand U1252 (N_1252,N_1240,N_1203);
nor U1253 (N_1253,N_1223,N_1216);
or U1254 (N_1254,N_1246,N_1230);
nand U1255 (N_1255,N_1237,N_1202);
and U1256 (N_1256,N_1239,N_1233);
or U1257 (N_1257,N_1211,N_1235);
xnor U1258 (N_1258,N_1220,N_1245);
nor U1259 (N_1259,N_1248,N_1215);
or U1260 (N_1260,N_1242,N_1208);
and U1261 (N_1261,N_1227,N_1228);
or U1262 (N_1262,N_1221,N_1229);
nor U1263 (N_1263,N_1232,N_1201);
and U1264 (N_1264,N_1249,N_1236);
or U1265 (N_1265,N_1225,N_1200);
or U1266 (N_1266,N_1209,N_1224);
nor U1267 (N_1267,N_1219,N_1205);
and U1268 (N_1268,N_1241,N_1234);
or U1269 (N_1269,N_1238,N_1218);
and U1270 (N_1270,N_1243,N_1214);
and U1271 (N_1271,N_1212,N_1247);
nand U1272 (N_1272,N_1244,N_1207);
nor U1273 (N_1273,N_1217,N_1231);
and U1274 (N_1274,N_1226,N_1213);
nand U1275 (N_1275,N_1206,N_1237);
or U1276 (N_1276,N_1247,N_1201);
nand U1277 (N_1277,N_1223,N_1245);
nand U1278 (N_1278,N_1247,N_1200);
nor U1279 (N_1279,N_1225,N_1213);
nor U1280 (N_1280,N_1223,N_1247);
nor U1281 (N_1281,N_1216,N_1217);
or U1282 (N_1282,N_1225,N_1240);
or U1283 (N_1283,N_1223,N_1220);
and U1284 (N_1284,N_1232,N_1221);
and U1285 (N_1285,N_1216,N_1209);
nor U1286 (N_1286,N_1213,N_1240);
nor U1287 (N_1287,N_1220,N_1240);
or U1288 (N_1288,N_1230,N_1206);
nand U1289 (N_1289,N_1228,N_1218);
or U1290 (N_1290,N_1214,N_1224);
xnor U1291 (N_1291,N_1240,N_1238);
nor U1292 (N_1292,N_1223,N_1237);
nand U1293 (N_1293,N_1209,N_1235);
or U1294 (N_1294,N_1220,N_1214);
and U1295 (N_1295,N_1229,N_1203);
nand U1296 (N_1296,N_1241,N_1224);
or U1297 (N_1297,N_1203,N_1219);
nand U1298 (N_1298,N_1249,N_1219);
nor U1299 (N_1299,N_1239,N_1215);
and U1300 (N_1300,N_1277,N_1270);
or U1301 (N_1301,N_1263,N_1285);
or U1302 (N_1302,N_1297,N_1294);
and U1303 (N_1303,N_1256,N_1250);
and U1304 (N_1304,N_1278,N_1287);
and U1305 (N_1305,N_1266,N_1279);
or U1306 (N_1306,N_1299,N_1255);
nand U1307 (N_1307,N_1293,N_1253);
nand U1308 (N_1308,N_1288,N_1292);
nand U1309 (N_1309,N_1296,N_1254);
or U1310 (N_1310,N_1291,N_1290);
nand U1311 (N_1311,N_1257,N_1283);
or U1312 (N_1312,N_1289,N_1268);
nand U1313 (N_1313,N_1259,N_1261);
nand U1314 (N_1314,N_1258,N_1264);
and U1315 (N_1315,N_1282,N_1262);
nand U1316 (N_1316,N_1272,N_1271);
and U1317 (N_1317,N_1286,N_1267);
or U1318 (N_1318,N_1281,N_1252);
and U1319 (N_1319,N_1280,N_1274);
nand U1320 (N_1320,N_1265,N_1276);
nand U1321 (N_1321,N_1298,N_1284);
or U1322 (N_1322,N_1269,N_1251);
or U1323 (N_1323,N_1275,N_1295);
and U1324 (N_1324,N_1273,N_1260);
nor U1325 (N_1325,N_1278,N_1286);
or U1326 (N_1326,N_1267,N_1273);
nor U1327 (N_1327,N_1252,N_1279);
nand U1328 (N_1328,N_1297,N_1255);
nand U1329 (N_1329,N_1277,N_1266);
and U1330 (N_1330,N_1267,N_1259);
nor U1331 (N_1331,N_1277,N_1274);
nand U1332 (N_1332,N_1285,N_1295);
nand U1333 (N_1333,N_1262,N_1287);
and U1334 (N_1334,N_1264,N_1270);
and U1335 (N_1335,N_1290,N_1285);
nand U1336 (N_1336,N_1256,N_1283);
nor U1337 (N_1337,N_1299,N_1271);
or U1338 (N_1338,N_1264,N_1295);
nor U1339 (N_1339,N_1271,N_1269);
nor U1340 (N_1340,N_1288,N_1280);
and U1341 (N_1341,N_1280,N_1268);
or U1342 (N_1342,N_1266,N_1281);
and U1343 (N_1343,N_1290,N_1296);
or U1344 (N_1344,N_1294,N_1262);
or U1345 (N_1345,N_1297,N_1266);
and U1346 (N_1346,N_1276,N_1278);
nor U1347 (N_1347,N_1289,N_1269);
or U1348 (N_1348,N_1295,N_1271);
or U1349 (N_1349,N_1280,N_1251);
and U1350 (N_1350,N_1348,N_1323);
and U1351 (N_1351,N_1306,N_1300);
or U1352 (N_1352,N_1344,N_1328);
nor U1353 (N_1353,N_1308,N_1339);
nand U1354 (N_1354,N_1309,N_1321);
nand U1355 (N_1355,N_1337,N_1303);
or U1356 (N_1356,N_1301,N_1318);
nor U1357 (N_1357,N_1331,N_1326);
nand U1358 (N_1358,N_1342,N_1305);
or U1359 (N_1359,N_1349,N_1335);
nand U1360 (N_1360,N_1319,N_1315);
nand U1361 (N_1361,N_1311,N_1307);
or U1362 (N_1362,N_1312,N_1343);
and U1363 (N_1363,N_1338,N_1310);
nor U1364 (N_1364,N_1314,N_1334);
nand U1365 (N_1365,N_1341,N_1330);
nand U1366 (N_1366,N_1316,N_1313);
and U1367 (N_1367,N_1327,N_1332);
nand U1368 (N_1368,N_1322,N_1320);
nand U1369 (N_1369,N_1302,N_1317);
nor U1370 (N_1370,N_1325,N_1329);
nor U1371 (N_1371,N_1345,N_1340);
nand U1372 (N_1372,N_1304,N_1333);
nor U1373 (N_1373,N_1347,N_1336);
or U1374 (N_1374,N_1346,N_1324);
or U1375 (N_1375,N_1340,N_1315);
or U1376 (N_1376,N_1326,N_1340);
or U1377 (N_1377,N_1306,N_1308);
or U1378 (N_1378,N_1336,N_1346);
nor U1379 (N_1379,N_1325,N_1310);
or U1380 (N_1380,N_1301,N_1329);
or U1381 (N_1381,N_1311,N_1333);
nand U1382 (N_1382,N_1323,N_1339);
nor U1383 (N_1383,N_1304,N_1323);
and U1384 (N_1384,N_1303,N_1324);
or U1385 (N_1385,N_1349,N_1317);
and U1386 (N_1386,N_1326,N_1337);
and U1387 (N_1387,N_1349,N_1344);
and U1388 (N_1388,N_1324,N_1330);
nand U1389 (N_1389,N_1326,N_1318);
nor U1390 (N_1390,N_1324,N_1302);
and U1391 (N_1391,N_1342,N_1304);
nand U1392 (N_1392,N_1307,N_1328);
nor U1393 (N_1393,N_1301,N_1342);
nand U1394 (N_1394,N_1328,N_1303);
or U1395 (N_1395,N_1315,N_1345);
or U1396 (N_1396,N_1311,N_1336);
and U1397 (N_1397,N_1305,N_1300);
or U1398 (N_1398,N_1330,N_1319);
or U1399 (N_1399,N_1319,N_1332);
and U1400 (N_1400,N_1360,N_1367);
nand U1401 (N_1401,N_1384,N_1355);
or U1402 (N_1402,N_1375,N_1356);
and U1403 (N_1403,N_1388,N_1376);
or U1404 (N_1404,N_1383,N_1370);
or U1405 (N_1405,N_1369,N_1366);
and U1406 (N_1406,N_1393,N_1396);
or U1407 (N_1407,N_1365,N_1350);
or U1408 (N_1408,N_1379,N_1387);
or U1409 (N_1409,N_1372,N_1353);
and U1410 (N_1410,N_1395,N_1354);
and U1411 (N_1411,N_1363,N_1380);
and U1412 (N_1412,N_1378,N_1352);
or U1413 (N_1413,N_1374,N_1389);
nand U1414 (N_1414,N_1358,N_1361);
nand U1415 (N_1415,N_1391,N_1357);
or U1416 (N_1416,N_1382,N_1390);
and U1417 (N_1417,N_1368,N_1394);
or U1418 (N_1418,N_1385,N_1381);
or U1419 (N_1419,N_1397,N_1373);
nand U1420 (N_1420,N_1386,N_1399);
and U1421 (N_1421,N_1362,N_1398);
or U1422 (N_1422,N_1371,N_1351);
nor U1423 (N_1423,N_1364,N_1359);
or U1424 (N_1424,N_1392,N_1377);
nor U1425 (N_1425,N_1374,N_1359);
or U1426 (N_1426,N_1385,N_1380);
and U1427 (N_1427,N_1379,N_1353);
nand U1428 (N_1428,N_1357,N_1359);
and U1429 (N_1429,N_1384,N_1363);
nor U1430 (N_1430,N_1395,N_1365);
or U1431 (N_1431,N_1379,N_1378);
and U1432 (N_1432,N_1392,N_1399);
or U1433 (N_1433,N_1380,N_1389);
or U1434 (N_1434,N_1365,N_1379);
or U1435 (N_1435,N_1376,N_1385);
nor U1436 (N_1436,N_1384,N_1389);
or U1437 (N_1437,N_1364,N_1399);
nand U1438 (N_1438,N_1353,N_1373);
or U1439 (N_1439,N_1396,N_1376);
nand U1440 (N_1440,N_1390,N_1371);
nor U1441 (N_1441,N_1354,N_1388);
nor U1442 (N_1442,N_1374,N_1397);
and U1443 (N_1443,N_1393,N_1390);
and U1444 (N_1444,N_1390,N_1377);
xor U1445 (N_1445,N_1373,N_1357);
nand U1446 (N_1446,N_1394,N_1385);
or U1447 (N_1447,N_1387,N_1360);
or U1448 (N_1448,N_1399,N_1375);
or U1449 (N_1449,N_1374,N_1371);
nand U1450 (N_1450,N_1406,N_1413);
nand U1451 (N_1451,N_1425,N_1442);
and U1452 (N_1452,N_1436,N_1449);
or U1453 (N_1453,N_1434,N_1441);
nand U1454 (N_1454,N_1411,N_1445);
and U1455 (N_1455,N_1408,N_1447);
nor U1456 (N_1456,N_1437,N_1429);
and U1457 (N_1457,N_1421,N_1409);
nor U1458 (N_1458,N_1443,N_1431);
or U1459 (N_1459,N_1402,N_1404);
nand U1460 (N_1460,N_1424,N_1414);
or U1461 (N_1461,N_1415,N_1401);
nand U1462 (N_1462,N_1419,N_1416);
or U1463 (N_1463,N_1422,N_1400);
nor U1464 (N_1464,N_1417,N_1428);
or U1465 (N_1465,N_1438,N_1427);
nand U1466 (N_1466,N_1432,N_1430);
nor U1467 (N_1467,N_1407,N_1444);
and U1468 (N_1468,N_1405,N_1448);
nor U1469 (N_1469,N_1435,N_1439);
nand U1470 (N_1470,N_1423,N_1410);
and U1471 (N_1471,N_1433,N_1446);
nand U1472 (N_1472,N_1403,N_1420);
or U1473 (N_1473,N_1440,N_1426);
and U1474 (N_1474,N_1418,N_1412);
nand U1475 (N_1475,N_1442,N_1428);
nand U1476 (N_1476,N_1419,N_1437);
and U1477 (N_1477,N_1411,N_1402);
nor U1478 (N_1478,N_1444,N_1410);
or U1479 (N_1479,N_1440,N_1412);
or U1480 (N_1480,N_1419,N_1435);
nor U1481 (N_1481,N_1434,N_1440);
xor U1482 (N_1482,N_1429,N_1400);
or U1483 (N_1483,N_1446,N_1445);
nand U1484 (N_1484,N_1416,N_1425);
and U1485 (N_1485,N_1407,N_1422);
or U1486 (N_1486,N_1426,N_1439);
and U1487 (N_1487,N_1408,N_1439);
nand U1488 (N_1488,N_1430,N_1436);
or U1489 (N_1489,N_1420,N_1433);
or U1490 (N_1490,N_1440,N_1415);
and U1491 (N_1491,N_1409,N_1403);
nor U1492 (N_1492,N_1435,N_1406);
nor U1493 (N_1493,N_1441,N_1444);
nor U1494 (N_1494,N_1432,N_1415);
nor U1495 (N_1495,N_1422,N_1410);
or U1496 (N_1496,N_1429,N_1427);
nor U1497 (N_1497,N_1400,N_1405);
xor U1498 (N_1498,N_1422,N_1447);
nand U1499 (N_1499,N_1445,N_1438);
nor U1500 (N_1500,N_1457,N_1472);
or U1501 (N_1501,N_1462,N_1497);
nor U1502 (N_1502,N_1488,N_1461);
nand U1503 (N_1503,N_1474,N_1465);
nand U1504 (N_1504,N_1475,N_1491);
nor U1505 (N_1505,N_1489,N_1470);
nand U1506 (N_1506,N_1478,N_1494);
and U1507 (N_1507,N_1499,N_1493);
nand U1508 (N_1508,N_1498,N_1496);
or U1509 (N_1509,N_1463,N_1484);
or U1510 (N_1510,N_1490,N_1452);
or U1511 (N_1511,N_1466,N_1492);
nor U1512 (N_1512,N_1486,N_1469);
or U1513 (N_1513,N_1480,N_1468);
or U1514 (N_1514,N_1459,N_1453);
nor U1515 (N_1515,N_1464,N_1485);
and U1516 (N_1516,N_1450,N_1456);
nor U1517 (N_1517,N_1451,N_1482);
nand U1518 (N_1518,N_1476,N_1471);
or U1519 (N_1519,N_1477,N_1460);
nand U1520 (N_1520,N_1479,N_1455);
nand U1521 (N_1521,N_1481,N_1495);
nor U1522 (N_1522,N_1473,N_1454);
or U1523 (N_1523,N_1483,N_1458);
nand U1524 (N_1524,N_1487,N_1467);
or U1525 (N_1525,N_1476,N_1492);
or U1526 (N_1526,N_1482,N_1464);
and U1527 (N_1527,N_1459,N_1491);
and U1528 (N_1528,N_1472,N_1496);
nand U1529 (N_1529,N_1490,N_1472);
nor U1530 (N_1530,N_1482,N_1476);
nor U1531 (N_1531,N_1488,N_1478);
and U1532 (N_1532,N_1481,N_1496);
nor U1533 (N_1533,N_1480,N_1492);
or U1534 (N_1534,N_1459,N_1456);
nand U1535 (N_1535,N_1456,N_1458);
nor U1536 (N_1536,N_1481,N_1469);
or U1537 (N_1537,N_1469,N_1474);
nor U1538 (N_1538,N_1488,N_1497);
nand U1539 (N_1539,N_1474,N_1490);
or U1540 (N_1540,N_1459,N_1498);
nor U1541 (N_1541,N_1469,N_1487);
nor U1542 (N_1542,N_1472,N_1480);
nand U1543 (N_1543,N_1458,N_1496);
nor U1544 (N_1544,N_1466,N_1481);
and U1545 (N_1545,N_1486,N_1487);
or U1546 (N_1546,N_1475,N_1460);
or U1547 (N_1547,N_1481,N_1465);
nor U1548 (N_1548,N_1469,N_1453);
and U1549 (N_1549,N_1495,N_1450);
xor U1550 (N_1550,N_1522,N_1532);
or U1551 (N_1551,N_1545,N_1517);
and U1552 (N_1552,N_1546,N_1521);
nand U1553 (N_1553,N_1541,N_1519);
nor U1554 (N_1554,N_1505,N_1531);
nor U1555 (N_1555,N_1533,N_1549);
or U1556 (N_1556,N_1527,N_1530);
and U1557 (N_1557,N_1515,N_1539);
nand U1558 (N_1558,N_1503,N_1524);
nand U1559 (N_1559,N_1544,N_1511);
nand U1560 (N_1560,N_1500,N_1529);
nor U1561 (N_1561,N_1537,N_1523);
nor U1562 (N_1562,N_1502,N_1518);
or U1563 (N_1563,N_1514,N_1513);
nor U1564 (N_1564,N_1526,N_1536);
nand U1565 (N_1565,N_1508,N_1504);
nand U1566 (N_1566,N_1512,N_1516);
nor U1567 (N_1567,N_1525,N_1510);
xnor U1568 (N_1568,N_1507,N_1538);
and U1569 (N_1569,N_1534,N_1528);
and U1570 (N_1570,N_1540,N_1506);
nand U1571 (N_1571,N_1547,N_1548);
and U1572 (N_1572,N_1543,N_1535);
nor U1573 (N_1573,N_1501,N_1509);
and U1574 (N_1574,N_1520,N_1542);
nor U1575 (N_1575,N_1533,N_1510);
nor U1576 (N_1576,N_1533,N_1531);
nand U1577 (N_1577,N_1533,N_1502);
nand U1578 (N_1578,N_1545,N_1507);
and U1579 (N_1579,N_1517,N_1527);
nor U1580 (N_1580,N_1504,N_1529);
nand U1581 (N_1581,N_1533,N_1538);
nand U1582 (N_1582,N_1512,N_1519);
or U1583 (N_1583,N_1526,N_1549);
and U1584 (N_1584,N_1527,N_1545);
or U1585 (N_1585,N_1536,N_1512);
or U1586 (N_1586,N_1520,N_1521);
or U1587 (N_1587,N_1520,N_1530);
nand U1588 (N_1588,N_1545,N_1502);
or U1589 (N_1589,N_1514,N_1512);
or U1590 (N_1590,N_1536,N_1548);
or U1591 (N_1591,N_1500,N_1518);
nor U1592 (N_1592,N_1511,N_1532);
nor U1593 (N_1593,N_1538,N_1511);
and U1594 (N_1594,N_1516,N_1545);
nand U1595 (N_1595,N_1513,N_1549);
nand U1596 (N_1596,N_1511,N_1540);
or U1597 (N_1597,N_1519,N_1528);
and U1598 (N_1598,N_1549,N_1531);
nand U1599 (N_1599,N_1529,N_1535);
nor U1600 (N_1600,N_1597,N_1595);
nand U1601 (N_1601,N_1573,N_1574);
nand U1602 (N_1602,N_1551,N_1568);
or U1603 (N_1603,N_1594,N_1586);
and U1604 (N_1604,N_1581,N_1567);
or U1605 (N_1605,N_1564,N_1552);
and U1606 (N_1606,N_1578,N_1592);
and U1607 (N_1607,N_1579,N_1560);
or U1608 (N_1608,N_1575,N_1591);
xnor U1609 (N_1609,N_1582,N_1550);
nor U1610 (N_1610,N_1565,N_1598);
and U1611 (N_1611,N_1557,N_1593);
and U1612 (N_1612,N_1596,N_1584);
nand U1613 (N_1613,N_1566,N_1553);
nand U1614 (N_1614,N_1555,N_1590);
and U1615 (N_1615,N_1572,N_1570);
and U1616 (N_1616,N_1558,N_1576);
or U1617 (N_1617,N_1562,N_1571);
nor U1618 (N_1618,N_1569,N_1585);
or U1619 (N_1619,N_1587,N_1559);
nand U1620 (N_1620,N_1554,N_1583);
and U1621 (N_1621,N_1561,N_1599);
and U1622 (N_1622,N_1577,N_1580);
nand U1623 (N_1623,N_1563,N_1556);
nand U1624 (N_1624,N_1589,N_1588);
and U1625 (N_1625,N_1593,N_1582);
nor U1626 (N_1626,N_1582,N_1590);
nor U1627 (N_1627,N_1584,N_1597);
or U1628 (N_1628,N_1572,N_1554);
nand U1629 (N_1629,N_1581,N_1575);
nand U1630 (N_1630,N_1577,N_1596);
nor U1631 (N_1631,N_1555,N_1569);
nor U1632 (N_1632,N_1575,N_1598);
nand U1633 (N_1633,N_1552,N_1569);
nor U1634 (N_1634,N_1591,N_1553);
nand U1635 (N_1635,N_1597,N_1576);
or U1636 (N_1636,N_1584,N_1593);
nor U1637 (N_1637,N_1594,N_1575);
nor U1638 (N_1638,N_1593,N_1581);
nor U1639 (N_1639,N_1572,N_1573);
nor U1640 (N_1640,N_1596,N_1564);
or U1641 (N_1641,N_1599,N_1557);
nand U1642 (N_1642,N_1567,N_1583);
or U1643 (N_1643,N_1571,N_1572);
nand U1644 (N_1644,N_1563,N_1576);
and U1645 (N_1645,N_1584,N_1566);
nand U1646 (N_1646,N_1577,N_1552);
nand U1647 (N_1647,N_1585,N_1577);
nand U1648 (N_1648,N_1569,N_1579);
nand U1649 (N_1649,N_1579,N_1580);
nand U1650 (N_1650,N_1646,N_1600);
nand U1651 (N_1651,N_1622,N_1611);
nand U1652 (N_1652,N_1627,N_1639);
and U1653 (N_1653,N_1619,N_1647);
and U1654 (N_1654,N_1624,N_1610);
and U1655 (N_1655,N_1601,N_1603);
and U1656 (N_1656,N_1604,N_1607);
or U1657 (N_1657,N_1625,N_1628);
nand U1658 (N_1658,N_1616,N_1636);
nand U1659 (N_1659,N_1641,N_1615);
nor U1660 (N_1660,N_1618,N_1634);
or U1661 (N_1661,N_1637,N_1612);
or U1662 (N_1662,N_1609,N_1631);
nand U1663 (N_1663,N_1648,N_1614);
and U1664 (N_1664,N_1630,N_1608);
nand U1665 (N_1665,N_1605,N_1620);
nand U1666 (N_1666,N_1617,N_1644);
nor U1667 (N_1667,N_1640,N_1643);
nand U1668 (N_1668,N_1638,N_1621);
and U1669 (N_1669,N_1602,N_1629);
or U1670 (N_1670,N_1626,N_1632);
or U1671 (N_1671,N_1623,N_1613);
and U1672 (N_1672,N_1645,N_1606);
nand U1673 (N_1673,N_1649,N_1642);
and U1674 (N_1674,N_1635,N_1633);
or U1675 (N_1675,N_1629,N_1623);
and U1676 (N_1676,N_1645,N_1610);
nand U1677 (N_1677,N_1641,N_1629);
or U1678 (N_1678,N_1632,N_1637);
and U1679 (N_1679,N_1601,N_1620);
and U1680 (N_1680,N_1644,N_1620);
nor U1681 (N_1681,N_1637,N_1620);
nand U1682 (N_1682,N_1646,N_1638);
or U1683 (N_1683,N_1644,N_1634);
nor U1684 (N_1684,N_1611,N_1616);
nor U1685 (N_1685,N_1637,N_1608);
or U1686 (N_1686,N_1645,N_1644);
or U1687 (N_1687,N_1635,N_1631);
nand U1688 (N_1688,N_1649,N_1619);
or U1689 (N_1689,N_1649,N_1608);
and U1690 (N_1690,N_1615,N_1631);
nor U1691 (N_1691,N_1645,N_1613);
and U1692 (N_1692,N_1614,N_1621);
or U1693 (N_1693,N_1633,N_1639);
nor U1694 (N_1694,N_1608,N_1612);
nor U1695 (N_1695,N_1642,N_1645);
nor U1696 (N_1696,N_1631,N_1606);
and U1697 (N_1697,N_1604,N_1628);
and U1698 (N_1698,N_1625,N_1631);
nor U1699 (N_1699,N_1601,N_1624);
or U1700 (N_1700,N_1677,N_1680);
nand U1701 (N_1701,N_1668,N_1676);
nor U1702 (N_1702,N_1682,N_1652);
and U1703 (N_1703,N_1685,N_1690);
nor U1704 (N_1704,N_1695,N_1671);
or U1705 (N_1705,N_1692,N_1679);
nor U1706 (N_1706,N_1689,N_1670);
or U1707 (N_1707,N_1678,N_1675);
nor U1708 (N_1708,N_1686,N_1659);
nand U1709 (N_1709,N_1672,N_1693);
and U1710 (N_1710,N_1655,N_1674);
nor U1711 (N_1711,N_1650,N_1669);
or U1712 (N_1712,N_1664,N_1696);
nand U1713 (N_1713,N_1663,N_1698);
and U1714 (N_1714,N_1651,N_1681);
or U1715 (N_1715,N_1691,N_1657);
nand U1716 (N_1716,N_1673,N_1684);
nor U1717 (N_1717,N_1654,N_1666);
nor U1718 (N_1718,N_1656,N_1665);
nand U1719 (N_1719,N_1667,N_1658);
or U1720 (N_1720,N_1662,N_1697);
nand U1721 (N_1721,N_1660,N_1699);
xnor U1722 (N_1722,N_1653,N_1661);
and U1723 (N_1723,N_1683,N_1688);
and U1724 (N_1724,N_1687,N_1694);
nor U1725 (N_1725,N_1671,N_1682);
or U1726 (N_1726,N_1690,N_1695);
and U1727 (N_1727,N_1688,N_1687);
and U1728 (N_1728,N_1664,N_1677);
nand U1729 (N_1729,N_1686,N_1664);
or U1730 (N_1730,N_1669,N_1698);
and U1731 (N_1731,N_1666,N_1690);
or U1732 (N_1732,N_1694,N_1695);
nor U1733 (N_1733,N_1689,N_1662);
nor U1734 (N_1734,N_1665,N_1674);
nand U1735 (N_1735,N_1651,N_1683);
or U1736 (N_1736,N_1690,N_1664);
nor U1737 (N_1737,N_1692,N_1695);
nor U1738 (N_1738,N_1665,N_1676);
or U1739 (N_1739,N_1651,N_1685);
nor U1740 (N_1740,N_1674,N_1690);
nand U1741 (N_1741,N_1669,N_1686);
or U1742 (N_1742,N_1696,N_1672);
and U1743 (N_1743,N_1663,N_1689);
and U1744 (N_1744,N_1666,N_1676);
and U1745 (N_1745,N_1653,N_1657);
or U1746 (N_1746,N_1687,N_1689);
nand U1747 (N_1747,N_1666,N_1658);
or U1748 (N_1748,N_1683,N_1660);
and U1749 (N_1749,N_1694,N_1676);
or U1750 (N_1750,N_1705,N_1720);
nand U1751 (N_1751,N_1736,N_1746);
and U1752 (N_1752,N_1725,N_1748);
and U1753 (N_1753,N_1712,N_1733);
or U1754 (N_1754,N_1729,N_1741);
or U1755 (N_1755,N_1737,N_1745);
nor U1756 (N_1756,N_1727,N_1703);
and U1757 (N_1757,N_1708,N_1719);
or U1758 (N_1758,N_1742,N_1743);
or U1759 (N_1759,N_1730,N_1714);
or U1760 (N_1760,N_1735,N_1739);
and U1761 (N_1761,N_1716,N_1749);
nor U1762 (N_1762,N_1724,N_1713);
and U1763 (N_1763,N_1706,N_1709);
nor U1764 (N_1764,N_1717,N_1715);
nand U1765 (N_1765,N_1744,N_1738);
nor U1766 (N_1766,N_1711,N_1740);
nor U1767 (N_1767,N_1701,N_1731);
or U1768 (N_1768,N_1702,N_1707);
nand U1769 (N_1769,N_1718,N_1728);
nand U1770 (N_1770,N_1726,N_1732);
nand U1771 (N_1771,N_1723,N_1721);
or U1772 (N_1772,N_1710,N_1704);
nand U1773 (N_1773,N_1722,N_1734);
nor U1774 (N_1774,N_1747,N_1700);
and U1775 (N_1775,N_1724,N_1700);
nand U1776 (N_1776,N_1716,N_1738);
nand U1777 (N_1777,N_1722,N_1724);
nor U1778 (N_1778,N_1724,N_1723);
nand U1779 (N_1779,N_1734,N_1725);
and U1780 (N_1780,N_1733,N_1725);
nand U1781 (N_1781,N_1714,N_1708);
nand U1782 (N_1782,N_1730,N_1705);
nor U1783 (N_1783,N_1726,N_1704);
nand U1784 (N_1784,N_1733,N_1736);
nand U1785 (N_1785,N_1733,N_1739);
nor U1786 (N_1786,N_1715,N_1742);
nor U1787 (N_1787,N_1725,N_1706);
or U1788 (N_1788,N_1734,N_1702);
nand U1789 (N_1789,N_1711,N_1743);
nand U1790 (N_1790,N_1703,N_1729);
nand U1791 (N_1791,N_1743,N_1740);
or U1792 (N_1792,N_1712,N_1749);
nor U1793 (N_1793,N_1726,N_1749);
or U1794 (N_1794,N_1729,N_1706);
and U1795 (N_1795,N_1744,N_1739);
or U1796 (N_1796,N_1707,N_1722);
or U1797 (N_1797,N_1739,N_1713);
and U1798 (N_1798,N_1727,N_1729);
nand U1799 (N_1799,N_1739,N_1709);
or U1800 (N_1800,N_1799,N_1765);
or U1801 (N_1801,N_1761,N_1785);
or U1802 (N_1802,N_1778,N_1796);
and U1803 (N_1803,N_1771,N_1784);
nand U1804 (N_1804,N_1763,N_1781);
and U1805 (N_1805,N_1782,N_1754);
or U1806 (N_1806,N_1792,N_1774);
or U1807 (N_1807,N_1770,N_1794);
nand U1808 (N_1808,N_1764,N_1777);
or U1809 (N_1809,N_1769,N_1772);
and U1810 (N_1810,N_1768,N_1773);
or U1811 (N_1811,N_1776,N_1760);
or U1812 (N_1812,N_1793,N_1753);
and U1813 (N_1813,N_1758,N_1788);
or U1814 (N_1814,N_1797,N_1787);
or U1815 (N_1815,N_1756,N_1752);
nand U1816 (N_1816,N_1779,N_1751);
or U1817 (N_1817,N_1750,N_1786);
or U1818 (N_1818,N_1795,N_1780);
or U1819 (N_1819,N_1798,N_1791);
nor U1820 (N_1820,N_1762,N_1783);
nand U1821 (N_1821,N_1775,N_1790);
nor U1822 (N_1822,N_1789,N_1766);
and U1823 (N_1823,N_1759,N_1755);
nand U1824 (N_1824,N_1767,N_1757);
nor U1825 (N_1825,N_1777,N_1793);
nand U1826 (N_1826,N_1767,N_1778);
nor U1827 (N_1827,N_1780,N_1779);
nand U1828 (N_1828,N_1755,N_1779);
or U1829 (N_1829,N_1794,N_1790);
nor U1830 (N_1830,N_1756,N_1767);
nand U1831 (N_1831,N_1790,N_1797);
nand U1832 (N_1832,N_1796,N_1785);
nor U1833 (N_1833,N_1785,N_1798);
and U1834 (N_1834,N_1789,N_1773);
or U1835 (N_1835,N_1782,N_1795);
nor U1836 (N_1836,N_1785,N_1792);
or U1837 (N_1837,N_1783,N_1788);
and U1838 (N_1838,N_1767,N_1766);
nand U1839 (N_1839,N_1797,N_1778);
nor U1840 (N_1840,N_1760,N_1799);
nand U1841 (N_1841,N_1790,N_1762);
nor U1842 (N_1842,N_1794,N_1754);
nor U1843 (N_1843,N_1788,N_1782);
nor U1844 (N_1844,N_1798,N_1779);
or U1845 (N_1845,N_1795,N_1784);
nand U1846 (N_1846,N_1786,N_1796);
or U1847 (N_1847,N_1797,N_1781);
or U1848 (N_1848,N_1799,N_1774);
or U1849 (N_1849,N_1758,N_1791);
or U1850 (N_1850,N_1847,N_1843);
and U1851 (N_1851,N_1817,N_1834);
nor U1852 (N_1852,N_1837,N_1819);
nor U1853 (N_1853,N_1829,N_1836);
and U1854 (N_1854,N_1818,N_1845);
nor U1855 (N_1855,N_1844,N_1806);
nand U1856 (N_1856,N_1813,N_1800);
nand U1857 (N_1857,N_1825,N_1808);
and U1858 (N_1858,N_1846,N_1841);
nand U1859 (N_1859,N_1805,N_1826);
or U1860 (N_1860,N_1810,N_1814);
or U1861 (N_1861,N_1821,N_1801);
and U1862 (N_1862,N_1838,N_1820);
nand U1863 (N_1863,N_1822,N_1809);
or U1864 (N_1864,N_1830,N_1849);
nor U1865 (N_1865,N_1811,N_1842);
nand U1866 (N_1866,N_1833,N_1804);
nand U1867 (N_1867,N_1840,N_1835);
nand U1868 (N_1868,N_1807,N_1802);
nand U1869 (N_1869,N_1848,N_1812);
nor U1870 (N_1870,N_1828,N_1824);
or U1871 (N_1871,N_1815,N_1839);
and U1872 (N_1872,N_1832,N_1803);
and U1873 (N_1873,N_1823,N_1831);
nor U1874 (N_1874,N_1816,N_1827);
and U1875 (N_1875,N_1800,N_1834);
nor U1876 (N_1876,N_1838,N_1845);
nor U1877 (N_1877,N_1803,N_1823);
nor U1878 (N_1878,N_1817,N_1830);
nor U1879 (N_1879,N_1832,N_1821);
nand U1880 (N_1880,N_1824,N_1811);
and U1881 (N_1881,N_1814,N_1800);
nand U1882 (N_1882,N_1832,N_1836);
nand U1883 (N_1883,N_1824,N_1822);
nor U1884 (N_1884,N_1835,N_1849);
and U1885 (N_1885,N_1807,N_1836);
and U1886 (N_1886,N_1831,N_1832);
nor U1887 (N_1887,N_1800,N_1803);
or U1888 (N_1888,N_1814,N_1828);
nor U1889 (N_1889,N_1800,N_1807);
and U1890 (N_1890,N_1810,N_1820);
xnor U1891 (N_1891,N_1800,N_1846);
and U1892 (N_1892,N_1820,N_1807);
nor U1893 (N_1893,N_1811,N_1825);
nor U1894 (N_1894,N_1827,N_1821);
and U1895 (N_1895,N_1836,N_1839);
and U1896 (N_1896,N_1812,N_1818);
nor U1897 (N_1897,N_1803,N_1834);
nand U1898 (N_1898,N_1846,N_1837);
nor U1899 (N_1899,N_1810,N_1804);
and U1900 (N_1900,N_1881,N_1898);
and U1901 (N_1901,N_1888,N_1851);
and U1902 (N_1902,N_1882,N_1871);
nor U1903 (N_1903,N_1879,N_1854);
nand U1904 (N_1904,N_1890,N_1857);
and U1905 (N_1905,N_1877,N_1886);
nor U1906 (N_1906,N_1884,N_1897);
nor U1907 (N_1907,N_1872,N_1889);
and U1908 (N_1908,N_1875,N_1891);
or U1909 (N_1909,N_1883,N_1870);
nand U1910 (N_1910,N_1899,N_1887);
and U1911 (N_1911,N_1873,N_1855);
nor U1912 (N_1912,N_1880,N_1853);
nor U1913 (N_1913,N_1864,N_1856);
or U1914 (N_1914,N_1861,N_1892);
nor U1915 (N_1915,N_1895,N_1852);
xnor U1916 (N_1916,N_1878,N_1866);
nand U1917 (N_1917,N_1868,N_1893);
nand U1918 (N_1918,N_1876,N_1894);
nor U1919 (N_1919,N_1869,N_1858);
or U1920 (N_1920,N_1867,N_1865);
and U1921 (N_1921,N_1874,N_1860);
nor U1922 (N_1922,N_1863,N_1896);
and U1923 (N_1923,N_1862,N_1859);
and U1924 (N_1924,N_1850,N_1885);
or U1925 (N_1925,N_1896,N_1862);
nand U1926 (N_1926,N_1856,N_1877);
nor U1927 (N_1927,N_1865,N_1877);
or U1928 (N_1928,N_1872,N_1875);
nor U1929 (N_1929,N_1893,N_1898);
or U1930 (N_1930,N_1875,N_1860);
and U1931 (N_1931,N_1863,N_1867);
nor U1932 (N_1932,N_1889,N_1859);
nor U1933 (N_1933,N_1889,N_1866);
and U1934 (N_1934,N_1881,N_1851);
nor U1935 (N_1935,N_1872,N_1863);
nand U1936 (N_1936,N_1875,N_1857);
and U1937 (N_1937,N_1858,N_1891);
nand U1938 (N_1938,N_1884,N_1869);
and U1939 (N_1939,N_1887,N_1879);
nor U1940 (N_1940,N_1897,N_1885);
nand U1941 (N_1941,N_1869,N_1897);
nor U1942 (N_1942,N_1879,N_1875);
nand U1943 (N_1943,N_1862,N_1855);
nor U1944 (N_1944,N_1878,N_1893);
and U1945 (N_1945,N_1898,N_1888);
nor U1946 (N_1946,N_1896,N_1870);
nand U1947 (N_1947,N_1859,N_1867);
and U1948 (N_1948,N_1876,N_1870);
or U1949 (N_1949,N_1882,N_1892);
nand U1950 (N_1950,N_1918,N_1948);
and U1951 (N_1951,N_1919,N_1931);
and U1952 (N_1952,N_1923,N_1922);
nand U1953 (N_1953,N_1930,N_1940);
nor U1954 (N_1954,N_1926,N_1939);
nor U1955 (N_1955,N_1938,N_1934);
nand U1956 (N_1956,N_1902,N_1907);
nand U1957 (N_1957,N_1906,N_1947);
nor U1958 (N_1958,N_1927,N_1903);
or U1959 (N_1959,N_1932,N_1921);
and U1960 (N_1960,N_1929,N_1904);
or U1961 (N_1961,N_1915,N_1925);
nor U1962 (N_1962,N_1949,N_1901);
nor U1963 (N_1963,N_1913,N_1912);
nor U1964 (N_1964,N_1936,N_1909);
or U1965 (N_1965,N_1928,N_1941);
nand U1966 (N_1966,N_1933,N_1924);
nor U1967 (N_1967,N_1944,N_1900);
nor U1968 (N_1968,N_1916,N_1946);
nor U1969 (N_1969,N_1908,N_1911);
nor U1970 (N_1970,N_1905,N_1917);
nand U1971 (N_1971,N_1914,N_1935);
nor U1972 (N_1972,N_1920,N_1942);
nor U1973 (N_1973,N_1943,N_1937);
nor U1974 (N_1974,N_1945,N_1910);
and U1975 (N_1975,N_1902,N_1920);
or U1976 (N_1976,N_1915,N_1918);
or U1977 (N_1977,N_1941,N_1932);
and U1978 (N_1978,N_1910,N_1912);
nor U1979 (N_1979,N_1909,N_1918);
nand U1980 (N_1980,N_1921,N_1949);
or U1981 (N_1981,N_1920,N_1923);
nor U1982 (N_1982,N_1924,N_1930);
xnor U1983 (N_1983,N_1937,N_1944);
and U1984 (N_1984,N_1948,N_1921);
or U1985 (N_1985,N_1915,N_1938);
and U1986 (N_1986,N_1901,N_1933);
nor U1987 (N_1987,N_1923,N_1929);
and U1988 (N_1988,N_1911,N_1910);
nor U1989 (N_1989,N_1917,N_1931);
nand U1990 (N_1990,N_1936,N_1942);
and U1991 (N_1991,N_1949,N_1937);
nand U1992 (N_1992,N_1912,N_1923);
or U1993 (N_1993,N_1949,N_1945);
nand U1994 (N_1994,N_1939,N_1933);
nand U1995 (N_1995,N_1939,N_1936);
and U1996 (N_1996,N_1902,N_1946);
and U1997 (N_1997,N_1940,N_1914);
nor U1998 (N_1998,N_1928,N_1914);
or U1999 (N_1999,N_1905,N_1911);
or U2000 (N_2000,N_1995,N_1997);
or U2001 (N_2001,N_1975,N_1988);
or U2002 (N_2002,N_1979,N_1963);
or U2003 (N_2003,N_1953,N_1980);
nand U2004 (N_2004,N_1985,N_1982);
nand U2005 (N_2005,N_1977,N_1957);
or U2006 (N_2006,N_1960,N_1973);
or U2007 (N_2007,N_1994,N_1971);
nor U2008 (N_2008,N_1969,N_1966);
and U2009 (N_2009,N_1952,N_1967);
and U2010 (N_2010,N_1987,N_1968);
and U2011 (N_2011,N_1996,N_1998);
and U2012 (N_2012,N_1981,N_1964);
and U2013 (N_2013,N_1974,N_1958);
or U2014 (N_2014,N_1959,N_1993);
and U2015 (N_2015,N_1954,N_1950);
and U2016 (N_2016,N_1983,N_1991);
or U2017 (N_2017,N_1992,N_1976);
nand U2018 (N_2018,N_1961,N_1972);
nand U2019 (N_2019,N_1989,N_1970);
nand U2020 (N_2020,N_1999,N_1986);
nor U2021 (N_2021,N_1956,N_1984);
and U2022 (N_2022,N_1955,N_1965);
and U2023 (N_2023,N_1990,N_1978);
nor U2024 (N_2024,N_1962,N_1951);
nand U2025 (N_2025,N_1988,N_1958);
nor U2026 (N_2026,N_1980,N_1956);
nor U2027 (N_2027,N_1969,N_1987);
and U2028 (N_2028,N_1981,N_1959);
nor U2029 (N_2029,N_1981,N_1995);
nor U2030 (N_2030,N_1960,N_1961);
or U2031 (N_2031,N_1990,N_1967);
nor U2032 (N_2032,N_1975,N_1982);
nand U2033 (N_2033,N_1961,N_1957);
or U2034 (N_2034,N_1958,N_1956);
nand U2035 (N_2035,N_1950,N_1976);
nor U2036 (N_2036,N_1967,N_1954);
and U2037 (N_2037,N_1985,N_1979);
and U2038 (N_2038,N_1980,N_1969);
or U2039 (N_2039,N_1984,N_1976);
nor U2040 (N_2040,N_1984,N_1988);
nand U2041 (N_2041,N_1987,N_1999);
nor U2042 (N_2042,N_1994,N_1979);
nor U2043 (N_2043,N_1995,N_1958);
or U2044 (N_2044,N_1992,N_1977);
nor U2045 (N_2045,N_1992,N_1979);
or U2046 (N_2046,N_1995,N_1957);
nor U2047 (N_2047,N_1986,N_1953);
and U2048 (N_2048,N_1961,N_1990);
nor U2049 (N_2049,N_1961,N_1973);
and U2050 (N_2050,N_2033,N_2012);
or U2051 (N_2051,N_2026,N_2038);
nand U2052 (N_2052,N_2025,N_2035);
nand U2053 (N_2053,N_2010,N_2004);
nor U2054 (N_2054,N_2023,N_2008);
nand U2055 (N_2055,N_2022,N_2016);
or U2056 (N_2056,N_2049,N_2034);
and U2057 (N_2057,N_2029,N_2011);
and U2058 (N_2058,N_2037,N_2036);
nor U2059 (N_2059,N_2047,N_2046);
or U2060 (N_2060,N_2021,N_2000);
nand U2061 (N_2061,N_2039,N_2028);
nand U2062 (N_2062,N_2040,N_2043);
nor U2063 (N_2063,N_2041,N_2001);
and U2064 (N_2064,N_2032,N_2044);
and U2065 (N_2065,N_2020,N_2005);
xor U2066 (N_2066,N_2002,N_2024);
xnor U2067 (N_2067,N_2030,N_2031);
or U2068 (N_2068,N_2006,N_2019);
and U2069 (N_2069,N_2027,N_2014);
or U2070 (N_2070,N_2045,N_2048);
nor U2071 (N_2071,N_2007,N_2017);
and U2072 (N_2072,N_2042,N_2009);
nand U2073 (N_2073,N_2018,N_2015);
nor U2074 (N_2074,N_2003,N_2013);
and U2075 (N_2075,N_2039,N_2011);
nand U2076 (N_2076,N_2049,N_2048);
or U2077 (N_2077,N_2028,N_2041);
or U2078 (N_2078,N_2028,N_2033);
and U2079 (N_2079,N_2005,N_2041);
nor U2080 (N_2080,N_2042,N_2045);
and U2081 (N_2081,N_2003,N_2008);
and U2082 (N_2082,N_2041,N_2035);
or U2083 (N_2083,N_2026,N_2045);
nor U2084 (N_2084,N_2031,N_2000);
or U2085 (N_2085,N_2038,N_2041);
and U2086 (N_2086,N_2024,N_2037);
or U2087 (N_2087,N_2041,N_2012);
nor U2088 (N_2088,N_2001,N_2032);
nand U2089 (N_2089,N_2011,N_2048);
nor U2090 (N_2090,N_2033,N_2049);
nor U2091 (N_2091,N_2009,N_2000);
nor U2092 (N_2092,N_2035,N_2006);
and U2093 (N_2093,N_2047,N_2041);
nand U2094 (N_2094,N_2040,N_2032);
nand U2095 (N_2095,N_2021,N_2048);
nor U2096 (N_2096,N_2011,N_2002);
xor U2097 (N_2097,N_2004,N_2023);
and U2098 (N_2098,N_2040,N_2002);
nand U2099 (N_2099,N_2029,N_2047);
nor U2100 (N_2100,N_2086,N_2051);
or U2101 (N_2101,N_2074,N_2055);
or U2102 (N_2102,N_2089,N_2090);
or U2103 (N_2103,N_2066,N_2080);
nand U2104 (N_2104,N_2076,N_2072);
or U2105 (N_2105,N_2053,N_2096);
nand U2106 (N_2106,N_2094,N_2092);
or U2107 (N_2107,N_2088,N_2052);
and U2108 (N_2108,N_2079,N_2070);
and U2109 (N_2109,N_2064,N_2099);
nand U2110 (N_2110,N_2050,N_2068);
or U2111 (N_2111,N_2077,N_2069);
and U2112 (N_2112,N_2085,N_2095);
and U2113 (N_2113,N_2065,N_2084);
nand U2114 (N_2114,N_2073,N_2081);
and U2115 (N_2115,N_2067,N_2097);
nor U2116 (N_2116,N_2054,N_2061);
nand U2117 (N_2117,N_2082,N_2093);
nor U2118 (N_2118,N_2058,N_2083);
nor U2119 (N_2119,N_2060,N_2059);
nor U2120 (N_2120,N_2078,N_2057);
and U2121 (N_2121,N_2098,N_2063);
nor U2122 (N_2122,N_2087,N_2075);
and U2123 (N_2123,N_2056,N_2062);
or U2124 (N_2124,N_2071,N_2091);
nand U2125 (N_2125,N_2074,N_2052);
or U2126 (N_2126,N_2074,N_2093);
or U2127 (N_2127,N_2054,N_2072);
nor U2128 (N_2128,N_2096,N_2050);
and U2129 (N_2129,N_2072,N_2097);
and U2130 (N_2130,N_2057,N_2091);
nand U2131 (N_2131,N_2099,N_2094);
nand U2132 (N_2132,N_2072,N_2084);
and U2133 (N_2133,N_2051,N_2092);
or U2134 (N_2134,N_2056,N_2088);
nor U2135 (N_2135,N_2069,N_2051);
or U2136 (N_2136,N_2053,N_2078);
nor U2137 (N_2137,N_2083,N_2068);
or U2138 (N_2138,N_2058,N_2053);
nand U2139 (N_2139,N_2098,N_2070);
or U2140 (N_2140,N_2069,N_2092);
nor U2141 (N_2141,N_2086,N_2056);
nor U2142 (N_2142,N_2075,N_2058);
or U2143 (N_2143,N_2065,N_2064);
xor U2144 (N_2144,N_2073,N_2068);
nand U2145 (N_2145,N_2060,N_2098);
xor U2146 (N_2146,N_2078,N_2062);
and U2147 (N_2147,N_2093,N_2096);
or U2148 (N_2148,N_2070,N_2071);
nand U2149 (N_2149,N_2087,N_2062);
or U2150 (N_2150,N_2121,N_2115);
and U2151 (N_2151,N_2103,N_2135);
nand U2152 (N_2152,N_2148,N_2130);
nand U2153 (N_2153,N_2147,N_2128);
or U2154 (N_2154,N_2114,N_2112);
nor U2155 (N_2155,N_2119,N_2117);
nor U2156 (N_2156,N_2108,N_2145);
nand U2157 (N_2157,N_2101,N_2134);
nand U2158 (N_2158,N_2137,N_2143);
nand U2159 (N_2159,N_2125,N_2110);
and U2160 (N_2160,N_2118,N_2133);
and U2161 (N_2161,N_2100,N_2142);
or U2162 (N_2162,N_2126,N_2123);
and U2163 (N_2163,N_2132,N_2120);
nor U2164 (N_2164,N_2113,N_2124);
nor U2165 (N_2165,N_2146,N_2107);
nor U2166 (N_2166,N_2129,N_2122);
and U2167 (N_2167,N_2149,N_2144);
and U2168 (N_2168,N_2136,N_2105);
and U2169 (N_2169,N_2111,N_2102);
nand U2170 (N_2170,N_2109,N_2127);
or U2171 (N_2171,N_2131,N_2116);
and U2172 (N_2172,N_2139,N_2141);
nand U2173 (N_2173,N_2104,N_2106);
nor U2174 (N_2174,N_2140,N_2138);
nand U2175 (N_2175,N_2143,N_2130);
nand U2176 (N_2176,N_2141,N_2117);
nor U2177 (N_2177,N_2137,N_2121);
nand U2178 (N_2178,N_2103,N_2110);
nor U2179 (N_2179,N_2117,N_2122);
nor U2180 (N_2180,N_2141,N_2105);
nand U2181 (N_2181,N_2147,N_2146);
nor U2182 (N_2182,N_2113,N_2138);
nor U2183 (N_2183,N_2117,N_2113);
or U2184 (N_2184,N_2136,N_2143);
or U2185 (N_2185,N_2105,N_2147);
nand U2186 (N_2186,N_2116,N_2148);
nand U2187 (N_2187,N_2141,N_2137);
or U2188 (N_2188,N_2133,N_2127);
nand U2189 (N_2189,N_2149,N_2101);
nand U2190 (N_2190,N_2106,N_2130);
nor U2191 (N_2191,N_2118,N_2107);
nor U2192 (N_2192,N_2126,N_2122);
and U2193 (N_2193,N_2135,N_2115);
and U2194 (N_2194,N_2149,N_2121);
and U2195 (N_2195,N_2120,N_2105);
and U2196 (N_2196,N_2145,N_2135);
or U2197 (N_2197,N_2133,N_2124);
or U2198 (N_2198,N_2103,N_2149);
and U2199 (N_2199,N_2137,N_2109);
or U2200 (N_2200,N_2191,N_2174);
nor U2201 (N_2201,N_2193,N_2185);
and U2202 (N_2202,N_2176,N_2150);
nor U2203 (N_2203,N_2186,N_2167);
and U2204 (N_2204,N_2161,N_2195);
or U2205 (N_2205,N_2152,N_2164);
nor U2206 (N_2206,N_2170,N_2181);
and U2207 (N_2207,N_2151,N_2154);
or U2208 (N_2208,N_2178,N_2160);
or U2209 (N_2209,N_2155,N_2197);
nand U2210 (N_2210,N_2180,N_2168);
nor U2211 (N_2211,N_2190,N_2165);
nand U2212 (N_2212,N_2188,N_2184);
or U2213 (N_2213,N_2173,N_2199);
xnor U2214 (N_2214,N_2192,N_2153);
or U2215 (N_2215,N_2156,N_2196);
nand U2216 (N_2216,N_2189,N_2175);
or U2217 (N_2217,N_2163,N_2183);
nand U2218 (N_2218,N_2159,N_2171);
nor U2219 (N_2219,N_2179,N_2157);
and U2220 (N_2220,N_2162,N_2169);
and U2221 (N_2221,N_2172,N_2198);
or U2222 (N_2222,N_2158,N_2194);
nand U2223 (N_2223,N_2166,N_2187);
or U2224 (N_2224,N_2177,N_2182);
nor U2225 (N_2225,N_2192,N_2179);
xnor U2226 (N_2226,N_2183,N_2187);
and U2227 (N_2227,N_2158,N_2152);
and U2228 (N_2228,N_2160,N_2150);
or U2229 (N_2229,N_2186,N_2164);
nor U2230 (N_2230,N_2169,N_2178);
or U2231 (N_2231,N_2154,N_2159);
nor U2232 (N_2232,N_2188,N_2172);
or U2233 (N_2233,N_2166,N_2190);
nor U2234 (N_2234,N_2164,N_2177);
nor U2235 (N_2235,N_2156,N_2183);
or U2236 (N_2236,N_2195,N_2156);
nand U2237 (N_2237,N_2153,N_2197);
or U2238 (N_2238,N_2175,N_2193);
nor U2239 (N_2239,N_2194,N_2184);
or U2240 (N_2240,N_2152,N_2172);
nand U2241 (N_2241,N_2167,N_2162);
or U2242 (N_2242,N_2173,N_2159);
or U2243 (N_2243,N_2181,N_2178);
nand U2244 (N_2244,N_2162,N_2179);
nor U2245 (N_2245,N_2174,N_2155);
or U2246 (N_2246,N_2150,N_2195);
and U2247 (N_2247,N_2187,N_2167);
nor U2248 (N_2248,N_2157,N_2184);
and U2249 (N_2249,N_2152,N_2159);
and U2250 (N_2250,N_2206,N_2222);
or U2251 (N_2251,N_2229,N_2249);
nand U2252 (N_2252,N_2213,N_2227);
nand U2253 (N_2253,N_2240,N_2245);
or U2254 (N_2254,N_2216,N_2204);
or U2255 (N_2255,N_2223,N_2248);
nand U2256 (N_2256,N_2235,N_2203);
and U2257 (N_2257,N_2211,N_2232);
and U2258 (N_2258,N_2210,N_2231);
or U2259 (N_2259,N_2246,N_2215);
nor U2260 (N_2260,N_2221,N_2236);
nor U2261 (N_2261,N_2214,N_2207);
or U2262 (N_2262,N_2243,N_2201);
and U2263 (N_2263,N_2205,N_2219);
nor U2264 (N_2264,N_2233,N_2226);
nor U2265 (N_2265,N_2244,N_2224);
nor U2266 (N_2266,N_2230,N_2239);
nand U2267 (N_2267,N_2241,N_2200);
or U2268 (N_2268,N_2202,N_2220);
nand U2269 (N_2269,N_2242,N_2217);
and U2270 (N_2270,N_2225,N_2237);
or U2271 (N_2271,N_2209,N_2238);
nor U2272 (N_2272,N_2228,N_2218);
nand U2273 (N_2273,N_2247,N_2212);
and U2274 (N_2274,N_2234,N_2208);
and U2275 (N_2275,N_2229,N_2241);
nand U2276 (N_2276,N_2232,N_2235);
nor U2277 (N_2277,N_2212,N_2224);
or U2278 (N_2278,N_2209,N_2243);
nor U2279 (N_2279,N_2226,N_2240);
nand U2280 (N_2280,N_2226,N_2206);
nor U2281 (N_2281,N_2206,N_2246);
nor U2282 (N_2282,N_2228,N_2216);
nor U2283 (N_2283,N_2242,N_2248);
or U2284 (N_2284,N_2222,N_2228);
nor U2285 (N_2285,N_2207,N_2225);
nor U2286 (N_2286,N_2217,N_2216);
or U2287 (N_2287,N_2201,N_2228);
nor U2288 (N_2288,N_2224,N_2210);
nand U2289 (N_2289,N_2200,N_2202);
nand U2290 (N_2290,N_2218,N_2234);
or U2291 (N_2291,N_2220,N_2212);
and U2292 (N_2292,N_2205,N_2237);
and U2293 (N_2293,N_2216,N_2248);
nor U2294 (N_2294,N_2214,N_2225);
nand U2295 (N_2295,N_2249,N_2226);
nand U2296 (N_2296,N_2219,N_2241);
and U2297 (N_2297,N_2217,N_2232);
and U2298 (N_2298,N_2242,N_2201);
and U2299 (N_2299,N_2233,N_2200);
nor U2300 (N_2300,N_2269,N_2281);
nand U2301 (N_2301,N_2296,N_2294);
or U2302 (N_2302,N_2278,N_2289);
nor U2303 (N_2303,N_2274,N_2267);
nor U2304 (N_2304,N_2284,N_2250);
nand U2305 (N_2305,N_2259,N_2280);
nor U2306 (N_2306,N_2253,N_2263);
nor U2307 (N_2307,N_2283,N_2255);
nand U2308 (N_2308,N_2279,N_2260);
nand U2309 (N_2309,N_2295,N_2270);
nor U2310 (N_2310,N_2286,N_2276);
or U2311 (N_2311,N_2298,N_2291);
nor U2312 (N_2312,N_2277,N_2288);
or U2313 (N_2313,N_2266,N_2252);
nor U2314 (N_2314,N_2258,N_2256);
nor U2315 (N_2315,N_2275,N_2254);
and U2316 (N_2316,N_2297,N_2285);
or U2317 (N_2317,N_2272,N_2262);
and U2318 (N_2318,N_2292,N_2273);
nand U2319 (N_2319,N_2271,N_2251);
or U2320 (N_2320,N_2261,N_2293);
or U2321 (N_2321,N_2282,N_2257);
nand U2322 (N_2322,N_2299,N_2265);
nand U2323 (N_2323,N_2268,N_2264);
and U2324 (N_2324,N_2287,N_2290);
and U2325 (N_2325,N_2289,N_2283);
nand U2326 (N_2326,N_2273,N_2259);
or U2327 (N_2327,N_2274,N_2266);
or U2328 (N_2328,N_2290,N_2264);
nand U2329 (N_2329,N_2298,N_2256);
nor U2330 (N_2330,N_2270,N_2251);
and U2331 (N_2331,N_2277,N_2266);
nor U2332 (N_2332,N_2273,N_2271);
or U2333 (N_2333,N_2266,N_2281);
or U2334 (N_2334,N_2288,N_2289);
and U2335 (N_2335,N_2297,N_2298);
or U2336 (N_2336,N_2299,N_2268);
nand U2337 (N_2337,N_2264,N_2258);
or U2338 (N_2338,N_2253,N_2276);
nand U2339 (N_2339,N_2289,N_2276);
nand U2340 (N_2340,N_2285,N_2263);
nand U2341 (N_2341,N_2253,N_2265);
and U2342 (N_2342,N_2278,N_2251);
or U2343 (N_2343,N_2263,N_2273);
and U2344 (N_2344,N_2273,N_2267);
nand U2345 (N_2345,N_2288,N_2270);
or U2346 (N_2346,N_2263,N_2286);
nor U2347 (N_2347,N_2281,N_2267);
nor U2348 (N_2348,N_2284,N_2297);
nand U2349 (N_2349,N_2299,N_2295);
and U2350 (N_2350,N_2308,N_2322);
or U2351 (N_2351,N_2309,N_2310);
or U2352 (N_2352,N_2301,N_2307);
or U2353 (N_2353,N_2331,N_2304);
or U2354 (N_2354,N_2303,N_2341);
nor U2355 (N_2355,N_2324,N_2343);
nor U2356 (N_2356,N_2349,N_2345);
or U2357 (N_2357,N_2348,N_2317);
nand U2358 (N_2358,N_2344,N_2325);
nand U2359 (N_2359,N_2334,N_2330);
nor U2360 (N_2360,N_2339,N_2329);
nor U2361 (N_2361,N_2327,N_2333);
and U2362 (N_2362,N_2312,N_2337);
and U2363 (N_2363,N_2313,N_2326);
or U2364 (N_2364,N_2335,N_2336);
nor U2365 (N_2365,N_2340,N_2318);
and U2366 (N_2366,N_2328,N_2342);
nor U2367 (N_2367,N_2315,N_2321);
or U2368 (N_2368,N_2319,N_2338);
or U2369 (N_2369,N_2311,N_2323);
nor U2370 (N_2370,N_2314,N_2316);
nor U2371 (N_2371,N_2302,N_2347);
nor U2372 (N_2372,N_2300,N_2332);
nor U2373 (N_2373,N_2346,N_2320);
nand U2374 (N_2374,N_2306,N_2305);
nor U2375 (N_2375,N_2318,N_2342);
and U2376 (N_2376,N_2319,N_2339);
and U2377 (N_2377,N_2323,N_2343);
nor U2378 (N_2378,N_2338,N_2307);
nand U2379 (N_2379,N_2333,N_2303);
nor U2380 (N_2380,N_2327,N_2329);
or U2381 (N_2381,N_2323,N_2302);
nor U2382 (N_2382,N_2339,N_2343);
or U2383 (N_2383,N_2334,N_2310);
nand U2384 (N_2384,N_2327,N_2346);
nand U2385 (N_2385,N_2329,N_2345);
nor U2386 (N_2386,N_2328,N_2340);
nand U2387 (N_2387,N_2324,N_2338);
nor U2388 (N_2388,N_2340,N_2317);
nor U2389 (N_2389,N_2317,N_2320);
and U2390 (N_2390,N_2346,N_2344);
nand U2391 (N_2391,N_2329,N_2338);
and U2392 (N_2392,N_2319,N_2334);
and U2393 (N_2393,N_2324,N_2331);
nor U2394 (N_2394,N_2314,N_2346);
nand U2395 (N_2395,N_2320,N_2319);
nor U2396 (N_2396,N_2311,N_2331);
and U2397 (N_2397,N_2321,N_2318);
nand U2398 (N_2398,N_2311,N_2335);
and U2399 (N_2399,N_2325,N_2336);
or U2400 (N_2400,N_2393,N_2386);
nand U2401 (N_2401,N_2390,N_2371);
nand U2402 (N_2402,N_2377,N_2366);
nor U2403 (N_2403,N_2368,N_2396);
and U2404 (N_2404,N_2376,N_2387);
or U2405 (N_2405,N_2355,N_2399);
nor U2406 (N_2406,N_2357,N_2395);
nor U2407 (N_2407,N_2354,N_2391);
or U2408 (N_2408,N_2359,N_2381);
or U2409 (N_2409,N_2375,N_2392);
nand U2410 (N_2410,N_2385,N_2380);
nand U2411 (N_2411,N_2384,N_2373);
nor U2412 (N_2412,N_2382,N_2362);
nor U2413 (N_2413,N_2356,N_2363);
or U2414 (N_2414,N_2379,N_2398);
and U2415 (N_2415,N_2383,N_2394);
nand U2416 (N_2416,N_2370,N_2367);
nor U2417 (N_2417,N_2397,N_2365);
nor U2418 (N_2418,N_2353,N_2378);
nand U2419 (N_2419,N_2389,N_2361);
and U2420 (N_2420,N_2352,N_2350);
nor U2421 (N_2421,N_2351,N_2369);
and U2422 (N_2422,N_2358,N_2372);
nand U2423 (N_2423,N_2360,N_2388);
or U2424 (N_2424,N_2364,N_2374);
or U2425 (N_2425,N_2370,N_2392);
and U2426 (N_2426,N_2353,N_2398);
or U2427 (N_2427,N_2361,N_2375);
or U2428 (N_2428,N_2354,N_2363);
nand U2429 (N_2429,N_2384,N_2389);
nor U2430 (N_2430,N_2388,N_2385);
nor U2431 (N_2431,N_2383,N_2386);
nor U2432 (N_2432,N_2368,N_2382);
nand U2433 (N_2433,N_2389,N_2374);
nand U2434 (N_2434,N_2388,N_2356);
and U2435 (N_2435,N_2388,N_2397);
or U2436 (N_2436,N_2371,N_2392);
or U2437 (N_2437,N_2352,N_2391);
and U2438 (N_2438,N_2366,N_2375);
xnor U2439 (N_2439,N_2387,N_2369);
or U2440 (N_2440,N_2372,N_2363);
nor U2441 (N_2441,N_2394,N_2396);
nand U2442 (N_2442,N_2389,N_2355);
nor U2443 (N_2443,N_2388,N_2382);
or U2444 (N_2444,N_2367,N_2393);
nor U2445 (N_2445,N_2353,N_2375);
nor U2446 (N_2446,N_2383,N_2376);
nor U2447 (N_2447,N_2355,N_2383);
and U2448 (N_2448,N_2373,N_2356);
or U2449 (N_2449,N_2387,N_2386);
or U2450 (N_2450,N_2412,N_2427);
nor U2451 (N_2451,N_2413,N_2428);
nand U2452 (N_2452,N_2417,N_2434);
nor U2453 (N_2453,N_2438,N_2445);
and U2454 (N_2454,N_2431,N_2421);
or U2455 (N_2455,N_2419,N_2448);
nand U2456 (N_2456,N_2426,N_2414);
xor U2457 (N_2457,N_2401,N_2447);
nor U2458 (N_2458,N_2436,N_2449);
and U2459 (N_2459,N_2422,N_2415);
nand U2460 (N_2460,N_2424,N_2443);
and U2461 (N_2461,N_2402,N_2437);
nand U2462 (N_2462,N_2430,N_2441);
and U2463 (N_2463,N_2404,N_2410);
or U2464 (N_2464,N_2429,N_2432);
and U2465 (N_2465,N_2403,N_2406);
xnor U2466 (N_2466,N_2408,N_2411);
nor U2467 (N_2467,N_2423,N_2444);
and U2468 (N_2468,N_2442,N_2405);
or U2469 (N_2469,N_2420,N_2418);
xor U2470 (N_2470,N_2440,N_2435);
or U2471 (N_2471,N_2446,N_2409);
nand U2472 (N_2472,N_2407,N_2439);
nand U2473 (N_2473,N_2433,N_2416);
nor U2474 (N_2474,N_2400,N_2425);
nand U2475 (N_2475,N_2404,N_2441);
nor U2476 (N_2476,N_2448,N_2434);
nand U2477 (N_2477,N_2409,N_2406);
xnor U2478 (N_2478,N_2412,N_2413);
or U2479 (N_2479,N_2411,N_2449);
nor U2480 (N_2480,N_2424,N_2446);
and U2481 (N_2481,N_2420,N_2417);
and U2482 (N_2482,N_2424,N_2404);
or U2483 (N_2483,N_2424,N_2435);
xor U2484 (N_2484,N_2443,N_2431);
or U2485 (N_2485,N_2441,N_2443);
and U2486 (N_2486,N_2421,N_2448);
or U2487 (N_2487,N_2426,N_2436);
and U2488 (N_2488,N_2408,N_2432);
or U2489 (N_2489,N_2445,N_2448);
or U2490 (N_2490,N_2406,N_2434);
nor U2491 (N_2491,N_2424,N_2437);
and U2492 (N_2492,N_2435,N_2400);
nand U2493 (N_2493,N_2419,N_2404);
and U2494 (N_2494,N_2438,N_2401);
or U2495 (N_2495,N_2407,N_2444);
nand U2496 (N_2496,N_2439,N_2416);
or U2497 (N_2497,N_2410,N_2441);
and U2498 (N_2498,N_2401,N_2427);
or U2499 (N_2499,N_2400,N_2406);
nor U2500 (N_2500,N_2465,N_2490);
nand U2501 (N_2501,N_2487,N_2454);
nor U2502 (N_2502,N_2450,N_2471);
nand U2503 (N_2503,N_2452,N_2489);
and U2504 (N_2504,N_2478,N_2498);
and U2505 (N_2505,N_2468,N_2493);
or U2506 (N_2506,N_2467,N_2463);
and U2507 (N_2507,N_2474,N_2484);
nand U2508 (N_2508,N_2458,N_2470);
or U2509 (N_2509,N_2494,N_2455);
and U2510 (N_2510,N_2482,N_2473);
or U2511 (N_2511,N_2462,N_2492);
and U2512 (N_2512,N_2481,N_2466);
nand U2513 (N_2513,N_2495,N_2499);
nor U2514 (N_2514,N_2475,N_2460);
and U2515 (N_2515,N_2477,N_2472);
and U2516 (N_2516,N_2480,N_2451);
and U2517 (N_2517,N_2496,N_2476);
and U2518 (N_2518,N_2459,N_2464);
and U2519 (N_2519,N_2491,N_2456);
nand U2520 (N_2520,N_2488,N_2461);
and U2521 (N_2521,N_2483,N_2485);
or U2522 (N_2522,N_2469,N_2453);
and U2523 (N_2523,N_2457,N_2486);
nand U2524 (N_2524,N_2497,N_2479);
nor U2525 (N_2525,N_2483,N_2481);
and U2526 (N_2526,N_2467,N_2464);
or U2527 (N_2527,N_2486,N_2478);
nand U2528 (N_2528,N_2487,N_2460);
and U2529 (N_2529,N_2474,N_2452);
and U2530 (N_2530,N_2492,N_2484);
nor U2531 (N_2531,N_2463,N_2495);
nand U2532 (N_2532,N_2456,N_2473);
and U2533 (N_2533,N_2450,N_2477);
or U2534 (N_2534,N_2456,N_2471);
and U2535 (N_2535,N_2454,N_2451);
nor U2536 (N_2536,N_2498,N_2492);
nand U2537 (N_2537,N_2465,N_2475);
nor U2538 (N_2538,N_2495,N_2450);
nand U2539 (N_2539,N_2456,N_2487);
or U2540 (N_2540,N_2482,N_2490);
and U2541 (N_2541,N_2472,N_2494);
nor U2542 (N_2542,N_2463,N_2453);
or U2543 (N_2543,N_2471,N_2475);
nor U2544 (N_2544,N_2470,N_2499);
nor U2545 (N_2545,N_2485,N_2454);
nor U2546 (N_2546,N_2479,N_2461);
and U2547 (N_2547,N_2462,N_2459);
or U2548 (N_2548,N_2490,N_2476);
nor U2549 (N_2549,N_2453,N_2476);
nand U2550 (N_2550,N_2541,N_2536);
and U2551 (N_2551,N_2545,N_2512);
nand U2552 (N_2552,N_2535,N_2533);
nor U2553 (N_2553,N_2548,N_2534);
nor U2554 (N_2554,N_2505,N_2513);
or U2555 (N_2555,N_2524,N_2546);
or U2556 (N_2556,N_2540,N_2538);
nor U2557 (N_2557,N_2543,N_2503);
and U2558 (N_2558,N_2510,N_2547);
nand U2559 (N_2559,N_2526,N_2529);
or U2560 (N_2560,N_2542,N_2521);
and U2561 (N_2561,N_2504,N_2549);
or U2562 (N_2562,N_2530,N_2528);
nand U2563 (N_2563,N_2508,N_2516);
or U2564 (N_2564,N_2537,N_2507);
and U2565 (N_2565,N_2523,N_2527);
or U2566 (N_2566,N_2506,N_2517);
and U2567 (N_2567,N_2531,N_2544);
or U2568 (N_2568,N_2525,N_2539);
and U2569 (N_2569,N_2501,N_2522);
and U2570 (N_2570,N_2509,N_2500);
or U2571 (N_2571,N_2532,N_2518);
xnor U2572 (N_2572,N_2502,N_2514);
and U2573 (N_2573,N_2519,N_2515);
or U2574 (N_2574,N_2520,N_2511);
xor U2575 (N_2575,N_2538,N_2532);
and U2576 (N_2576,N_2512,N_2529);
nor U2577 (N_2577,N_2532,N_2524);
nand U2578 (N_2578,N_2546,N_2541);
and U2579 (N_2579,N_2540,N_2507);
nor U2580 (N_2580,N_2518,N_2535);
or U2581 (N_2581,N_2523,N_2545);
xnor U2582 (N_2582,N_2521,N_2531);
or U2583 (N_2583,N_2503,N_2531);
nand U2584 (N_2584,N_2506,N_2539);
nor U2585 (N_2585,N_2517,N_2527);
or U2586 (N_2586,N_2504,N_2543);
and U2587 (N_2587,N_2546,N_2539);
and U2588 (N_2588,N_2511,N_2513);
nand U2589 (N_2589,N_2514,N_2533);
nor U2590 (N_2590,N_2538,N_2502);
nand U2591 (N_2591,N_2513,N_2508);
and U2592 (N_2592,N_2526,N_2538);
nand U2593 (N_2593,N_2540,N_2508);
nor U2594 (N_2594,N_2513,N_2537);
nand U2595 (N_2595,N_2501,N_2517);
or U2596 (N_2596,N_2509,N_2527);
and U2597 (N_2597,N_2532,N_2517);
nor U2598 (N_2598,N_2546,N_2518);
nor U2599 (N_2599,N_2536,N_2548);
nor U2600 (N_2600,N_2596,N_2576);
or U2601 (N_2601,N_2556,N_2569);
and U2602 (N_2602,N_2554,N_2587);
or U2603 (N_2603,N_2599,N_2571);
or U2604 (N_2604,N_2593,N_2577);
and U2605 (N_2605,N_2586,N_2573);
and U2606 (N_2606,N_2575,N_2581);
nor U2607 (N_2607,N_2568,N_2572);
nand U2608 (N_2608,N_2550,N_2558);
nor U2609 (N_2609,N_2559,N_2592);
and U2610 (N_2610,N_2580,N_2564);
nand U2611 (N_2611,N_2552,N_2561);
nand U2612 (N_2612,N_2562,N_2565);
nor U2613 (N_2613,N_2560,N_2583);
and U2614 (N_2614,N_2551,N_2563);
nor U2615 (N_2615,N_2557,N_2597);
or U2616 (N_2616,N_2591,N_2570);
or U2617 (N_2617,N_2579,N_2594);
and U2618 (N_2618,N_2566,N_2595);
and U2619 (N_2619,N_2553,N_2584);
and U2620 (N_2620,N_2585,N_2589);
and U2621 (N_2621,N_2574,N_2555);
nor U2622 (N_2622,N_2582,N_2578);
or U2623 (N_2623,N_2598,N_2590);
or U2624 (N_2624,N_2567,N_2588);
nor U2625 (N_2625,N_2586,N_2556);
and U2626 (N_2626,N_2561,N_2556);
and U2627 (N_2627,N_2561,N_2567);
and U2628 (N_2628,N_2567,N_2598);
and U2629 (N_2629,N_2553,N_2597);
or U2630 (N_2630,N_2553,N_2593);
or U2631 (N_2631,N_2557,N_2572);
nor U2632 (N_2632,N_2587,N_2557);
or U2633 (N_2633,N_2597,N_2558);
nor U2634 (N_2634,N_2592,N_2568);
or U2635 (N_2635,N_2568,N_2590);
nand U2636 (N_2636,N_2556,N_2592);
nand U2637 (N_2637,N_2569,N_2573);
or U2638 (N_2638,N_2587,N_2563);
and U2639 (N_2639,N_2583,N_2580);
nand U2640 (N_2640,N_2551,N_2559);
nor U2641 (N_2641,N_2575,N_2582);
nor U2642 (N_2642,N_2555,N_2557);
or U2643 (N_2643,N_2573,N_2579);
nand U2644 (N_2644,N_2596,N_2555);
or U2645 (N_2645,N_2560,N_2585);
nor U2646 (N_2646,N_2591,N_2574);
and U2647 (N_2647,N_2559,N_2552);
or U2648 (N_2648,N_2567,N_2596);
and U2649 (N_2649,N_2590,N_2571);
nor U2650 (N_2650,N_2619,N_2629);
and U2651 (N_2651,N_2637,N_2636);
nor U2652 (N_2652,N_2607,N_2632);
nand U2653 (N_2653,N_2606,N_2649);
nand U2654 (N_2654,N_2645,N_2627);
and U2655 (N_2655,N_2610,N_2626);
and U2656 (N_2656,N_2638,N_2623);
nand U2657 (N_2657,N_2630,N_2646);
or U2658 (N_2658,N_2631,N_2605);
nor U2659 (N_2659,N_2621,N_2643);
or U2660 (N_2660,N_2603,N_2642);
nor U2661 (N_2661,N_2618,N_2616);
and U2662 (N_2662,N_2625,N_2602);
nand U2663 (N_2663,N_2611,N_2641);
nand U2664 (N_2664,N_2634,N_2628);
nor U2665 (N_2665,N_2635,N_2644);
or U2666 (N_2666,N_2600,N_2612);
and U2667 (N_2667,N_2613,N_2608);
or U2668 (N_2668,N_2639,N_2633);
or U2669 (N_2669,N_2624,N_2615);
nor U2670 (N_2670,N_2620,N_2622);
and U2671 (N_2671,N_2601,N_2604);
or U2672 (N_2672,N_2648,N_2614);
or U2673 (N_2673,N_2640,N_2609);
nand U2674 (N_2674,N_2647,N_2617);
nand U2675 (N_2675,N_2609,N_2621);
nor U2676 (N_2676,N_2604,N_2611);
nor U2677 (N_2677,N_2642,N_2640);
and U2678 (N_2678,N_2619,N_2647);
nand U2679 (N_2679,N_2614,N_2621);
nor U2680 (N_2680,N_2623,N_2604);
and U2681 (N_2681,N_2612,N_2614);
nand U2682 (N_2682,N_2603,N_2631);
nor U2683 (N_2683,N_2632,N_2605);
nand U2684 (N_2684,N_2609,N_2626);
and U2685 (N_2685,N_2623,N_2620);
or U2686 (N_2686,N_2616,N_2624);
nand U2687 (N_2687,N_2648,N_2605);
and U2688 (N_2688,N_2620,N_2630);
xnor U2689 (N_2689,N_2624,N_2621);
and U2690 (N_2690,N_2620,N_2637);
nor U2691 (N_2691,N_2631,N_2630);
and U2692 (N_2692,N_2633,N_2606);
nand U2693 (N_2693,N_2619,N_2602);
nor U2694 (N_2694,N_2611,N_2644);
or U2695 (N_2695,N_2637,N_2610);
or U2696 (N_2696,N_2619,N_2612);
or U2697 (N_2697,N_2600,N_2626);
and U2698 (N_2698,N_2601,N_2642);
xor U2699 (N_2699,N_2618,N_2638);
and U2700 (N_2700,N_2688,N_2651);
nand U2701 (N_2701,N_2662,N_2659);
xnor U2702 (N_2702,N_2673,N_2697);
or U2703 (N_2703,N_2685,N_2661);
nand U2704 (N_2704,N_2658,N_2660);
nand U2705 (N_2705,N_2667,N_2653);
or U2706 (N_2706,N_2678,N_2682);
nand U2707 (N_2707,N_2652,N_2671);
or U2708 (N_2708,N_2656,N_2664);
nor U2709 (N_2709,N_2699,N_2686);
and U2710 (N_2710,N_2670,N_2689);
or U2711 (N_2711,N_2695,N_2663);
nor U2712 (N_2712,N_2668,N_2654);
nand U2713 (N_2713,N_2692,N_2694);
and U2714 (N_2714,N_2680,N_2674);
or U2715 (N_2715,N_2675,N_2698);
or U2716 (N_2716,N_2691,N_2655);
and U2717 (N_2717,N_2690,N_2684);
nand U2718 (N_2718,N_2665,N_2677);
nor U2719 (N_2719,N_2693,N_2650);
and U2720 (N_2720,N_2672,N_2681);
nor U2721 (N_2721,N_2683,N_2657);
nor U2722 (N_2722,N_2687,N_2696);
nor U2723 (N_2723,N_2679,N_2666);
nand U2724 (N_2724,N_2669,N_2676);
or U2725 (N_2725,N_2699,N_2683);
nor U2726 (N_2726,N_2676,N_2692);
nand U2727 (N_2727,N_2688,N_2695);
and U2728 (N_2728,N_2650,N_2668);
nor U2729 (N_2729,N_2675,N_2679);
nand U2730 (N_2730,N_2674,N_2671);
and U2731 (N_2731,N_2659,N_2656);
and U2732 (N_2732,N_2650,N_2674);
and U2733 (N_2733,N_2663,N_2653);
nand U2734 (N_2734,N_2689,N_2652);
nand U2735 (N_2735,N_2652,N_2656);
xor U2736 (N_2736,N_2687,N_2692);
nand U2737 (N_2737,N_2694,N_2652);
or U2738 (N_2738,N_2693,N_2694);
and U2739 (N_2739,N_2673,N_2699);
xnor U2740 (N_2740,N_2683,N_2679);
nor U2741 (N_2741,N_2686,N_2697);
nor U2742 (N_2742,N_2696,N_2678);
nand U2743 (N_2743,N_2698,N_2659);
or U2744 (N_2744,N_2668,N_2672);
and U2745 (N_2745,N_2678,N_2671);
or U2746 (N_2746,N_2676,N_2673);
nor U2747 (N_2747,N_2674,N_2682);
and U2748 (N_2748,N_2699,N_2691);
nor U2749 (N_2749,N_2680,N_2667);
or U2750 (N_2750,N_2722,N_2748);
or U2751 (N_2751,N_2735,N_2704);
nor U2752 (N_2752,N_2729,N_2739);
nand U2753 (N_2753,N_2700,N_2721);
and U2754 (N_2754,N_2733,N_2723);
and U2755 (N_2755,N_2737,N_2726);
nand U2756 (N_2756,N_2731,N_2728);
and U2757 (N_2757,N_2742,N_2716);
and U2758 (N_2758,N_2705,N_2715);
and U2759 (N_2759,N_2709,N_2725);
or U2760 (N_2760,N_2727,N_2734);
or U2761 (N_2761,N_2701,N_2707);
nor U2762 (N_2762,N_2749,N_2724);
nand U2763 (N_2763,N_2718,N_2741);
nor U2764 (N_2764,N_2703,N_2712);
and U2765 (N_2765,N_2710,N_2732);
and U2766 (N_2766,N_2713,N_2740);
and U2767 (N_2767,N_2747,N_2746);
or U2768 (N_2768,N_2736,N_2708);
or U2769 (N_2769,N_2706,N_2702);
nand U2770 (N_2770,N_2738,N_2720);
or U2771 (N_2771,N_2730,N_2719);
nand U2772 (N_2772,N_2717,N_2711);
and U2773 (N_2773,N_2743,N_2714);
nand U2774 (N_2774,N_2745,N_2744);
and U2775 (N_2775,N_2709,N_2707);
or U2776 (N_2776,N_2742,N_2735);
or U2777 (N_2777,N_2736,N_2703);
or U2778 (N_2778,N_2726,N_2746);
and U2779 (N_2779,N_2712,N_2738);
and U2780 (N_2780,N_2716,N_2743);
nor U2781 (N_2781,N_2733,N_2740);
nor U2782 (N_2782,N_2747,N_2743);
nor U2783 (N_2783,N_2716,N_2711);
nand U2784 (N_2784,N_2700,N_2705);
nand U2785 (N_2785,N_2733,N_2729);
and U2786 (N_2786,N_2734,N_2747);
xnor U2787 (N_2787,N_2737,N_2728);
or U2788 (N_2788,N_2709,N_2722);
or U2789 (N_2789,N_2734,N_2730);
and U2790 (N_2790,N_2716,N_2730);
nor U2791 (N_2791,N_2714,N_2702);
or U2792 (N_2792,N_2705,N_2748);
or U2793 (N_2793,N_2701,N_2749);
nor U2794 (N_2794,N_2746,N_2713);
xor U2795 (N_2795,N_2714,N_2737);
nor U2796 (N_2796,N_2726,N_2700);
and U2797 (N_2797,N_2737,N_2721);
nand U2798 (N_2798,N_2733,N_2749);
and U2799 (N_2799,N_2725,N_2711);
or U2800 (N_2800,N_2777,N_2761);
or U2801 (N_2801,N_2753,N_2760);
or U2802 (N_2802,N_2785,N_2757);
or U2803 (N_2803,N_2787,N_2796);
nand U2804 (N_2804,N_2766,N_2773);
nand U2805 (N_2805,N_2771,N_2791);
nand U2806 (N_2806,N_2783,N_2776);
or U2807 (N_2807,N_2762,N_2790);
or U2808 (N_2808,N_2786,N_2792);
and U2809 (N_2809,N_2751,N_2794);
or U2810 (N_2810,N_2793,N_2770);
xor U2811 (N_2811,N_2795,N_2781);
and U2812 (N_2812,N_2754,N_2788);
nor U2813 (N_2813,N_2756,N_2772);
nand U2814 (N_2814,N_2782,N_2768);
nor U2815 (N_2815,N_2784,N_2789);
nand U2816 (N_2816,N_2755,N_2759);
or U2817 (N_2817,N_2752,N_2798);
nor U2818 (N_2818,N_2775,N_2758);
or U2819 (N_2819,N_2750,N_2767);
nor U2820 (N_2820,N_2764,N_2778);
nand U2821 (N_2821,N_2799,N_2765);
and U2822 (N_2822,N_2797,N_2763);
and U2823 (N_2823,N_2780,N_2769);
nand U2824 (N_2824,N_2774,N_2779);
and U2825 (N_2825,N_2780,N_2752);
and U2826 (N_2826,N_2794,N_2755);
nand U2827 (N_2827,N_2750,N_2799);
nor U2828 (N_2828,N_2787,N_2795);
and U2829 (N_2829,N_2781,N_2761);
and U2830 (N_2830,N_2781,N_2766);
nand U2831 (N_2831,N_2752,N_2794);
nand U2832 (N_2832,N_2774,N_2786);
or U2833 (N_2833,N_2787,N_2789);
nor U2834 (N_2834,N_2783,N_2773);
nand U2835 (N_2835,N_2761,N_2766);
and U2836 (N_2836,N_2772,N_2786);
nor U2837 (N_2837,N_2771,N_2778);
nor U2838 (N_2838,N_2782,N_2750);
nand U2839 (N_2839,N_2766,N_2795);
nor U2840 (N_2840,N_2772,N_2773);
or U2841 (N_2841,N_2779,N_2787);
and U2842 (N_2842,N_2764,N_2788);
or U2843 (N_2843,N_2763,N_2795);
nor U2844 (N_2844,N_2767,N_2751);
or U2845 (N_2845,N_2757,N_2778);
nand U2846 (N_2846,N_2757,N_2765);
or U2847 (N_2847,N_2766,N_2779);
nor U2848 (N_2848,N_2770,N_2767);
nor U2849 (N_2849,N_2757,N_2777);
or U2850 (N_2850,N_2827,N_2802);
nor U2851 (N_2851,N_2818,N_2842);
and U2852 (N_2852,N_2807,N_2822);
nor U2853 (N_2853,N_2812,N_2817);
nand U2854 (N_2854,N_2823,N_2820);
or U2855 (N_2855,N_2832,N_2849);
nor U2856 (N_2856,N_2813,N_2819);
or U2857 (N_2857,N_2829,N_2843);
or U2858 (N_2858,N_2806,N_2833);
nor U2859 (N_2859,N_2830,N_2805);
or U2860 (N_2860,N_2841,N_2815);
nor U2861 (N_2861,N_2831,N_2837);
nand U2862 (N_2862,N_2834,N_2824);
nor U2863 (N_2863,N_2839,N_2816);
nand U2864 (N_2864,N_2804,N_2826);
nand U2865 (N_2865,N_2840,N_2835);
nand U2866 (N_2866,N_2809,N_2800);
and U2867 (N_2867,N_2801,N_2847);
nand U2868 (N_2868,N_2846,N_2844);
nor U2869 (N_2869,N_2838,N_2808);
or U2870 (N_2870,N_2814,N_2821);
and U2871 (N_2871,N_2828,N_2803);
nor U2872 (N_2872,N_2811,N_2848);
and U2873 (N_2873,N_2845,N_2810);
nor U2874 (N_2874,N_2836,N_2825);
nor U2875 (N_2875,N_2841,N_2803);
and U2876 (N_2876,N_2836,N_2837);
and U2877 (N_2877,N_2801,N_2831);
nor U2878 (N_2878,N_2815,N_2811);
and U2879 (N_2879,N_2833,N_2809);
nand U2880 (N_2880,N_2815,N_2821);
and U2881 (N_2881,N_2824,N_2833);
or U2882 (N_2882,N_2811,N_2823);
nand U2883 (N_2883,N_2826,N_2843);
nor U2884 (N_2884,N_2848,N_2825);
nor U2885 (N_2885,N_2839,N_2806);
and U2886 (N_2886,N_2814,N_2804);
or U2887 (N_2887,N_2812,N_2840);
nor U2888 (N_2888,N_2825,N_2811);
nand U2889 (N_2889,N_2823,N_2834);
nand U2890 (N_2890,N_2808,N_2805);
and U2891 (N_2891,N_2823,N_2812);
and U2892 (N_2892,N_2848,N_2845);
or U2893 (N_2893,N_2848,N_2817);
and U2894 (N_2894,N_2810,N_2800);
nor U2895 (N_2895,N_2837,N_2827);
and U2896 (N_2896,N_2817,N_2820);
or U2897 (N_2897,N_2829,N_2831);
and U2898 (N_2898,N_2809,N_2825);
nor U2899 (N_2899,N_2838,N_2814);
and U2900 (N_2900,N_2859,N_2899);
nor U2901 (N_2901,N_2894,N_2896);
and U2902 (N_2902,N_2893,N_2889);
and U2903 (N_2903,N_2881,N_2862);
or U2904 (N_2904,N_2851,N_2883);
or U2905 (N_2905,N_2877,N_2898);
nand U2906 (N_2906,N_2880,N_2860);
and U2907 (N_2907,N_2886,N_2897);
and U2908 (N_2908,N_2875,N_2861);
or U2909 (N_2909,N_2867,N_2890);
or U2910 (N_2910,N_2857,N_2884);
or U2911 (N_2911,N_2870,N_2866);
nor U2912 (N_2912,N_2872,N_2885);
or U2913 (N_2913,N_2856,N_2854);
and U2914 (N_2914,N_2874,N_2852);
nor U2915 (N_2915,N_2882,N_2864);
nand U2916 (N_2916,N_2869,N_2871);
nor U2917 (N_2917,N_2887,N_2863);
and U2918 (N_2918,N_2855,N_2888);
and U2919 (N_2919,N_2868,N_2850);
nor U2920 (N_2920,N_2876,N_2865);
and U2921 (N_2921,N_2858,N_2895);
and U2922 (N_2922,N_2892,N_2878);
nor U2923 (N_2923,N_2873,N_2891);
nand U2924 (N_2924,N_2879,N_2853);
nor U2925 (N_2925,N_2876,N_2889);
and U2926 (N_2926,N_2856,N_2890);
or U2927 (N_2927,N_2892,N_2866);
nand U2928 (N_2928,N_2850,N_2895);
nor U2929 (N_2929,N_2884,N_2896);
and U2930 (N_2930,N_2863,N_2885);
and U2931 (N_2931,N_2886,N_2891);
nand U2932 (N_2932,N_2874,N_2857);
and U2933 (N_2933,N_2897,N_2899);
or U2934 (N_2934,N_2884,N_2851);
or U2935 (N_2935,N_2868,N_2878);
or U2936 (N_2936,N_2883,N_2884);
or U2937 (N_2937,N_2893,N_2864);
or U2938 (N_2938,N_2857,N_2872);
or U2939 (N_2939,N_2866,N_2868);
and U2940 (N_2940,N_2879,N_2861);
or U2941 (N_2941,N_2856,N_2885);
nor U2942 (N_2942,N_2899,N_2863);
or U2943 (N_2943,N_2854,N_2891);
or U2944 (N_2944,N_2893,N_2874);
nor U2945 (N_2945,N_2878,N_2897);
nand U2946 (N_2946,N_2861,N_2890);
nand U2947 (N_2947,N_2850,N_2878);
and U2948 (N_2948,N_2852,N_2867);
nand U2949 (N_2949,N_2893,N_2892);
nor U2950 (N_2950,N_2928,N_2929);
and U2951 (N_2951,N_2901,N_2941);
or U2952 (N_2952,N_2943,N_2914);
or U2953 (N_2953,N_2934,N_2917);
or U2954 (N_2954,N_2942,N_2937);
nand U2955 (N_2955,N_2911,N_2912);
nor U2956 (N_2956,N_2908,N_2906);
and U2957 (N_2957,N_2931,N_2925);
and U2958 (N_2958,N_2945,N_2900);
nand U2959 (N_2959,N_2946,N_2902);
or U2960 (N_2960,N_2936,N_2935);
or U2961 (N_2961,N_2938,N_2926);
or U2962 (N_2962,N_2920,N_2907);
and U2963 (N_2963,N_2913,N_2944);
or U2964 (N_2964,N_2924,N_2922);
nand U2965 (N_2965,N_2904,N_2939);
or U2966 (N_2966,N_2948,N_2915);
or U2967 (N_2967,N_2947,N_2918);
nor U2968 (N_2968,N_2903,N_2921);
and U2969 (N_2969,N_2927,N_2940);
nand U2970 (N_2970,N_2932,N_2909);
nand U2971 (N_2971,N_2933,N_2910);
nand U2972 (N_2972,N_2930,N_2916);
or U2973 (N_2973,N_2919,N_2949);
and U2974 (N_2974,N_2905,N_2923);
or U2975 (N_2975,N_2921,N_2901);
and U2976 (N_2976,N_2919,N_2903);
nor U2977 (N_2977,N_2911,N_2941);
or U2978 (N_2978,N_2906,N_2949);
and U2979 (N_2979,N_2933,N_2918);
and U2980 (N_2980,N_2933,N_2906);
and U2981 (N_2981,N_2903,N_2929);
nor U2982 (N_2982,N_2947,N_2933);
or U2983 (N_2983,N_2934,N_2904);
nor U2984 (N_2984,N_2948,N_2921);
nor U2985 (N_2985,N_2917,N_2933);
or U2986 (N_2986,N_2939,N_2918);
nand U2987 (N_2987,N_2947,N_2939);
and U2988 (N_2988,N_2921,N_2932);
or U2989 (N_2989,N_2903,N_2902);
and U2990 (N_2990,N_2930,N_2920);
and U2991 (N_2991,N_2943,N_2905);
or U2992 (N_2992,N_2906,N_2911);
nor U2993 (N_2993,N_2943,N_2942);
nor U2994 (N_2994,N_2945,N_2934);
or U2995 (N_2995,N_2901,N_2908);
nor U2996 (N_2996,N_2924,N_2908);
nor U2997 (N_2997,N_2920,N_2940);
or U2998 (N_2998,N_2926,N_2924);
xnor U2999 (N_2999,N_2949,N_2942);
nor UO_0 (O_0,N_2969,N_2988);
nand UO_1 (O_1,N_2960,N_2970);
nand UO_2 (O_2,N_2995,N_2984);
nand UO_3 (O_3,N_2950,N_2992);
and UO_4 (O_4,N_2952,N_2990);
and UO_5 (O_5,N_2953,N_2963);
and UO_6 (O_6,N_2987,N_2978);
and UO_7 (O_7,N_2954,N_2957);
or UO_8 (O_8,N_2982,N_2986);
and UO_9 (O_9,N_2951,N_2991);
and UO_10 (O_10,N_2959,N_2999);
nand UO_11 (O_11,N_2968,N_2983);
or UO_12 (O_12,N_2967,N_2971);
or UO_13 (O_13,N_2993,N_2976);
or UO_14 (O_14,N_2972,N_2985);
nand UO_15 (O_15,N_2965,N_2955);
nor UO_16 (O_16,N_2977,N_2964);
nor UO_17 (O_17,N_2997,N_2962);
or UO_18 (O_18,N_2996,N_2956);
or UO_19 (O_19,N_2973,N_2989);
nand UO_20 (O_20,N_2979,N_2975);
nand UO_21 (O_21,N_2958,N_2961);
nor UO_22 (O_22,N_2980,N_2974);
nor UO_23 (O_23,N_2998,N_2966);
nor UO_24 (O_24,N_2994,N_2981);
nand UO_25 (O_25,N_2953,N_2983);
or UO_26 (O_26,N_2982,N_2994);
or UO_27 (O_27,N_2961,N_2968);
nor UO_28 (O_28,N_2956,N_2950);
and UO_29 (O_29,N_2956,N_2981);
and UO_30 (O_30,N_2954,N_2983);
nor UO_31 (O_31,N_2984,N_2990);
or UO_32 (O_32,N_2986,N_2992);
nand UO_33 (O_33,N_2987,N_2955);
nand UO_34 (O_34,N_2967,N_2975);
xnor UO_35 (O_35,N_2963,N_2970);
and UO_36 (O_36,N_2989,N_2982);
and UO_37 (O_37,N_2963,N_2960);
nand UO_38 (O_38,N_2964,N_2951);
nand UO_39 (O_39,N_2974,N_2968);
nand UO_40 (O_40,N_2979,N_2998);
or UO_41 (O_41,N_2973,N_2964);
and UO_42 (O_42,N_2962,N_2985);
nand UO_43 (O_43,N_2997,N_2998);
nor UO_44 (O_44,N_2991,N_2954);
and UO_45 (O_45,N_2994,N_2990);
nand UO_46 (O_46,N_2978,N_2952);
nand UO_47 (O_47,N_2951,N_2956);
nor UO_48 (O_48,N_2970,N_2976);
and UO_49 (O_49,N_2950,N_2981);
nor UO_50 (O_50,N_2953,N_2967);
nand UO_51 (O_51,N_2955,N_2992);
or UO_52 (O_52,N_2989,N_2959);
nand UO_53 (O_53,N_2997,N_2968);
or UO_54 (O_54,N_2966,N_2983);
and UO_55 (O_55,N_2975,N_2970);
and UO_56 (O_56,N_2984,N_2991);
and UO_57 (O_57,N_2959,N_2985);
nor UO_58 (O_58,N_2981,N_2974);
nand UO_59 (O_59,N_2970,N_2953);
or UO_60 (O_60,N_2986,N_2978);
or UO_61 (O_61,N_2966,N_2953);
nor UO_62 (O_62,N_2961,N_2971);
nor UO_63 (O_63,N_2954,N_2966);
nor UO_64 (O_64,N_2959,N_2975);
and UO_65 (O_65,N_2993,N_2955);
nand UO_66 (O_66,N_2950,N_2979);
and UO_67 (O_67,N_2986,N_2950);
nand UO_68 (O_68,N_2991,N_2987);
and UO_69 (O_69,N_2983,N_2992);
or UO_70 (O_70,N_2977,N_2962);
nor UO_71 (O_71,N_2984,N_2965);
nor UO_72 (O_72,N_2989,N_2977);
nand UO_73 (O_73,N_2969,N_2982);
and UO_74 (O_74,N_2971,N_2989);
nor UO_75 (O_75,N_2988,N_2978);
and UO_76 (O_76,N_2984,N_2983);
nand UO_77 (O_77,N_2976,N_2977);
xor UO_78 (O_78,N_2959,N_2968);
nor UO_79 (O_79,N_2999,N_2993);
or UO_80 (O_80,N_2997,N_2990);
nand UO_81 (O_81,N_2968,N_2979);
nor UO_82 (O_82,N_2998,N_2955);
nand UO_83 (O_83,N_2968,N_2964);
and UO_84 (O_84,N_2974,N_2972);
and UO_85 (O_85,N_2968,N_2988);
or UO_86 (O_86,N_2993,N_2985);
nand UO_87 (O_87,N_2998,N_2958);
nor UO_88 (O_88,N_2991,N_2994);
nand UO_89 (O_89,N_2979,N_2987);
or UO_90 (O_90,N_2993,N_2996);
and UO_91 (O_91,N_2956,N_2982);
nand UO_92 (O_92,N_2988,N_2999);
nand UO_93 (O_93,N_2974,N_2997);
and UO_94 (O_94,N_2951,N_2996);
nand UO_95 (O_95,N_2997,N_2984);
nor UO_96 (O_96,N_2964,N_2970);
nor UO_97 (O_97,N_2972,N_2963);
or UO_98 (O_98,N_2950,N_2964);
or UO_99 (O_99,N_2973,N_2984);
and UO_100 (O_100,N_2977,N_2961);
nor UO_101 (O_101,N_2975,N_2989);
nand UO_102 (O_102,N_2984,N_2968);
nor UO_103 (O_103,N_2991,N_2966);
nand UO_104 (O_104,N_2989,N_2984);
nand UO_105 (O_105,N_2969,N_2958);
or UO_106 (O_106,N_2970,N_2998);
or UO_107 (O_107,N_2965,N_2990);
nand UO_108 (O_108,N_2988,N_2972);
nor UO_109 (O_109,N_2959,N_2957);
nand UO_110 (O_110,N_2987,N_2953);
or UO_111 (O_111,N_2995,N_2987);
and UO_112 (O_112,N_2956,N_2964);
nand UO_113 (O_113,N_2952,N_2977);
or UO_114 (O_114,N_2974,N_2975);
and UO_115 (O_115,N_2969,N_2968);
nor UO_116 (O_116,N_2976,N_2996);
or UO_117 (O_117,N_2985,N_2955);
nor UO_118 (O_118,N_2997,N_2956);
nand UO_119 (O_119,N_2991,N_2985);
nand UO_120 (O_120,N_2964,N_2981);
nand UO_121 (O_121,N_2972,N_2997);
or UO_122 (O_122,N_2953,N_2951);
or UO_123 (O_123,N_2996,N_2963);
nor UO_124 (O_124,N_2971,N_2998);
and UO_125 (O_125,N_2985,N_2967);
nand UO_126 (O_126,N_2966,N_2959);
and UO_127 (O_127,N_2980,N_2972);
nand UO_128 (O_128,N_2983,N_2957);
nor UO_129 (O_129,N_2978,N_2969);
nor UO_130 (O_130,N_2950,N_2970);
nor UO_131 (O_131,N_2966,N_2974);
nor UO_132 (O_132,N_2983,N_2988);
nand UO_133 (O_133,N_2985,N_2986);
or UO_134 (O_134,N_2970,N_2958);
nand UO_135 (O_135,N_2968,N_2973);
or UO_136 (O_136,N_2978,N_2990);
or UO_137 (O_137,N_2982,N_2993);
and UO_138 (O_138,N_2973,N_2976);
nor UO_139 (O_139,N_2956,N_2993);
nand UO_140 (O_140,N_2955,N_2976);
nand UO_141 (O_141,N_2959,N_2972);
and UO_142 (O_142,N_2996,N_2953);
or UO_143 (O_143,N_2992,N_2961);
nor UO_144 (O_144,N_2957,N_2951);
or UO_145 (O_145,N_2993,N_2969);
or UO_146 (O_146,N_2965,N_2952);
and UO_147 (O_147,N_2967,N_2950);
nand UO_148 (O_148,N_2955,N_2961);
nor UO_149 (O_149,N_2960,N_2988);
and UO_150 (O_150,N_2978,N_2957);
nor UO_151 (O_151,N_2973,N_2959);
or UO_152 (O_152,N_2967,N_2965);
nand UO_153 (O_153,N_2956,N_2971);
and UO_154 (O_154,N_2990,N_2987);
and UO_155 (O_155,N_2987,N_2950);
nor UO_156 (O_156,N_2963,N_2983);
and UO_157 (O_157,N_2969,N_2996);
or UO_158 (O_158,N_2971,N_2981);
or UO_159 (O_159,N_2961,N_2960);
nand UO_160 (O_160,N_2969,N_2999);
nand UO_161 (O_161,N_2975,N_2987);
nand UO_162 (O_162,N_2974,N_2988);
and UO_163 (O_163,N_2969,N_2966);
nor UO_164 (O_164,N_2966,N_2972);
and UO_165 (O_165,N_2950,N_2968);
or UO_166 (O_166,N_2952,N_2958);
or UO_167 (O_167,N_2968,N_2986);
nand UO_168 (O_168,N_2959,N_2956);
or UO_169 (O_169,N_2969,N_2984);
and UO_170 (O_170,N_2961,N_2998);
nand UO_171 (O_171,N_2987,N_2963);
nand UO_172 (O_172,N_2974,N_2956);
and UO_173 (O_173,N_2956,N_2965);
nand UO_174 (O_174,N_2980,N_2957);
and UO_175 (O_175,N_2987,N_2974);
nor UO_176 (O_176,N_2982,N_2968);
nand UO_177 (O_177,N_2995,N_2954);
xnor UO_178 (O_178,N_2980,N_2992);
and UO_179 (O_179,N_2953,N_2973);
nand UO_180 (O_180,N_2965,N_2968);
or UO_181 (O_181,N_2998,N_2999);
and UO_182 (O_182,N_2961,N_2978);
or UO_183 (O_183,N_2987,N_2983);
nor UO_184 (O_184,N_2954,N_2987);
nand UO_185 (O_185,N_2963,N_2977);
or UO_186 (O_186,N_2954,N_2982);
nand UO_187 (O_187,N_2987,N_2973);
or UO_188 (O_188,N_2997,N_2967);
or UO_189 (O_189,N_2991,N_2997);
nor UO_190 (O_190,N_2996,N_2973);
and UO_191 (O_191,N_2989,N_2974);
nor UO_192 (O_192,N_2972,N_2953);
nand UO_193 (O_193,N_2950,N_2954);
nor UO_194 (O_194,N_2990,N_2998);
nand UO_195 (O_195,N_2955,N_2954);
nor UO_196 (O_196,N_2954,N_2984);
nand UO_197 (O_197,N_2957,N_2968);
nand UO_198 (O_198,N_2998,N_2993);
nand UO_199 (O_199,N_2990,N_2955);
nor UO_200 (O_200,N_2986,N_2977);
nor UO_201 (O_201,N_2979,N_2993);
nand UO_202 (O_202,N_2983,N_2979);
and UO_203 (O_203,N_2967,N_2991);
and UO_204 (O_204,N_2956,N_2973);
or UO_205 (O_205,N_2962,N_2954);
or UO_206 (O_206,N_2997,N_2992);
nand UO_207 (O_207,N_2999,N_2989);
nand UO_208 (O_208,N_2988,N_2985);
nand UO_209 (O_209,N_2979,N_2966);
or UO_210 (O_210,N_2956,N_2963);
and UO_211 (O_211,N_2990,N_2996);
nand UO_212 (O_212,N_2958,N_2957);
nor UO_213 (O_213,N_2970,N_2973);
or UO_214 (O_214,N_2985,N_2956);
or UO_215 (O_215,N_2978,N_2979);
xor UO_216 (O_216,N_2960,N_2964);
and UO_217 (O_217,N_2966,N_2985);
or UO_218 (O_218,N_2979,N_2969);
and UO_219 (O_219,N_2961,N_2950);
nand UO_220 (O_220,N_2987,N_2998);
nand UO_221 (O_221,N_2988,N_2976);
and UO_222 (O_222,N_2973,N_2997);
or UO_223 (O_223,N_2972,N_2976);
and UO_224 (O_224,N_2993,N_2980);
or UO_225 (O_225,N_2988,N_2957);
and UO_226 (O_226,N_2977,N_2983);
and UO_227 (O_227,N_2958,N_2976);
or UO_228 (O_228,N_2997,N_2978);
or UO_229 (O_229,N_2976,N_2989);
nor UO_230 (O_230,N_2958,N_2972);
nand UO_231 (O_231,N_2970,N_2978);
nand UO_232 (O_232,N_2997,N_2980);
nor UO_233 (O_233,N_2988,N_2959);
nor UO_234 (O_234,N_2994,N_2989);
and UO_235 (O_235,N_2957,N_2960);
nand UO_236 (O_236,N_2986,N_2971);
nand UO_237 (O_237,N_2959,N_2974);
nand UO_238 (O_238,N_2984,N_2962);
and UO_239 (O_239,N_2959,N_2983);
or UO_240 (O_240,N_2979,N_2972);
nor UO_241 (O_241,N_2969,N_2998);
or UO_242 (O_242,N_2982,N_2950);
nor UO_243 (O_243,N_2989,N_2970);
nand UO_244 (O_244,N_2976,N_2954);
or UO_245 (O_245,N_2974,N_2985);
and UO_246 (O_246,N_2988,N_2967);
nand UO_247 (O_247,N_2968,N_2976);
or UO_248 (O_248,N_2955,N_2986);
or UO_249 (O_249,N_2992,N_2969);
nor UO_250 (O_250,N_2963,N_2961);
nor UO_251 (O_251,N_2950,N_2985);
nor UO_252 (O_252,N_2995,N_2997);
or UO_253 (O_253,N_2996,N_2981);
and UO_254 (O_254,N_2986,N_2952);
or UO_255 (O_255,N_2953,N_2979);
nor UO_256 (O_256,N_2966,N_2971);
nor UO_257 (O_257,N_2983,N_2964);
nor UO_258 (O_258,N_2952,N_2988);
and UO_259 (O_259,N_2981,N_2969);
and UO_260 (O_260,N_2965,N_2970);
or UO_261 (O_261,N_2990,N_2986);
or UO_262 (O_262,N_2950,N_2988);
nor UO_263 (O_263,N_2996,N_2989);
nor UO_264 (O_264,N_2965,N_2991);
and UO_265 (O_265,N_2968,N_2955);
and UO_266 (O_266,N_2998,N_2963);
nor UO_267 (O_267,N_2972,N_2951);
nand UO_268 (O_268,N_2991,N_2979);
and UO_269 (O_269,N_2966,N_2990);
and UO_270 (O_270,N_2967,N_2958);
and UO_271 (O_271,N_2954,N_2967);
or UO_272 (O_272,N_2979,N_2980);
nor UO_273 (O_273,N_2973,N_2999);
or UO_274 (O_274,N_2981,N_2988);
nor UO_275 (O_275,N_2984,N_2976);
and UO_276 (O_276,N_2962,N_2976);
or UO_277 (O_277,N_2980,N_2985);
and UO_278 (O_278,N_2982,N_2977);
and UO_279 (O_279,N_2959,N_2994);
nor UO_280 (O_280,N_2980,N_2991);
nand UO_281 (O_281,N_2953,N_2957);
or UO_282 (O_282,N_2976,N_2957);
nor UO_283 (O_283,N_2973,N_2986);
nor UO_284 (O_284,N_2971,N_2984);
nand UO_285 (O_285,N_2952,N_2964);
nor UO_286 (O_286,N_2954,N_2998);
or UO_287 (O_287,N_2993,N_2997);
nand UO_288 (O_288,N_2953,N_2994);
nand UO_289 (O_289,N_2959,N_2950);
and UO_290 (O_290,N_2993,N_2978);
and UO_291 (O_291,N_2975,N_2977);
nor UO_292 (O_292,N_2965,N_2964);
nor UO_293 (O_293,N_2988,N_2987);
nand UO_294 (O_294,N_2983,N_2970);
or UO_295 (O_295,N_2997,N_2950);
or UO_296 (O_296,N_2981,N_2995);
and UO_297 (O_297,N_2964,N_2957);
nor UO_298 (O_298,N_2975,N_2952);
or UO_299 (O_299,N_2994,N_2975);
nand UO_300 (O_300,N_2955,N_2966);
nor UO_301 (O_301,N_2993,N_2971);
nand UO_302 (O_302,N_2996,N_2959);
or UO_303 (O_303,N_2974,N_2967);
and UO_304 (O_304,N_2995,N_2969);
nand UO_305 (O_305,N_2955,N_2974);
or UO_306 (O_306,N_2967,N_2993);
nand UO_307 (O_307,N_2996,N_2992);
xnor UO_308 (O_308,N_2956,N_2980);
nor UO_309 (O_309,N_2996,N_2970);
nor UO_310 (O_310,N_2962,N_2980);
nand UO_311 (O_311,N_2999,N_2956);
or UO_312 (O_312,N_2964,N_2993);
or UO_313 (O_313,N_2987,N_2952);
or UO_314 (O_314,N_2953,N_2978);
or UO_315 (O_315,N_2985,N_2984);
and UO_316 (O_316,N_2972,N_2969);
nor UO_317 (O_317,N_2954,N_2972);
nor UO_318 (O_318,N_2992,N_2959);
nand UO_319 (O_319,N_2965,N_2998);
nand UO_320 (O_320,N_2989,N_2972);
and UO_321 (O_321,N_2956,N_2970);
and UO_322 (O_322,N_2965,N_2988);
nor UO_323 (O_323,N_2992,N_2981);
or UO_324 (O_324,N_2950,N_2958);
nand UO_325 (O_325,N_2992,N_2971);
or UO_326 (O_326,N_2987,N_2977);
and UO_327 (O_327,N_2998,N_2983);
nor UO_328 (O_328,N_2957,N_2991);
nand UO_329 (O_329,N_2951,N_2995);
or UO_330 (O_330,N_2960,N_2976);
nand UO_331 (O_331,N_2995,N_2994);
and UO_332 (O_332,N_2992,N_2952);
nand UO_333 (O_333,N_2982,N_2980);
nand UO_334 (O_334,N_2972,N_2999);
xor UO_335 (O_335,N_2992,N_2988);
or UO_336 (O_336,N_2983,N_2974);
or UO_337 (O_337,N_2958,N_2986);
nor UO_338 (O_338,N_2951,N_2962);
or UO_339 (O_339,N_2991,N_2995);
nand UO_340 (O_340,N_2994,N_2963);
nor UO_341 (O_341,N_2980,N_2968);
or UO_342 (O_342,N_2981,N_2993);
nand UO_343 (O_343,N_2999,N_2987);
nor UO_344 (O_344,N_2998,N_2985);
nand UO_345 (O_345,N_2998,N_2959);
and UO_346 (O_346,N_2974,N_2952);
nor UO_347 (O_347,N_2996,N_2955);
nor UO_348 (O_348,N_2970,N_2987);
or UO_349 (O_349,N_2975,N_2984);
nor UO_350 (O_350,N_2959,N_2955);
and UO_351 (O_351,N_2953,N_2952);
and UO_352 (O_352,N_2988,N_2984);
and UO_353 (O_353,N_2976,N_2975);
or UO_354 (O_354,N_2962,N_2973);
and UO_355 (O_355,N_2958,N_2999);
nand UO_356 (O_356,N_2951,N_2974);
nand UO_357 (O_357,N_2992,N_2964);
nor UO_358 (O_358,N_2957,N_2982);
nand UO_359 (O_359,N_2954,N_2994);
nand UO_360 (O_360,N_2989,N_2995);
nor UO_361 (O_361,N_2952,N_2956);
and UO_362 (O_362,N_2986,N_2969);
and UO_363 (O_363,N_2985,N_2976);
or UO_364 (O_364,N_2999,N_2971);
or UO_365 (O_365,N_2952,N_2981);
and UO_366 (O_366,N_2973,N_2977);
or UO_367 (O_367,N_2978,N_2956);
or UO_368 (O_368,N_2965,N_2958);
and UO_369 (O_369,N_2998,N_2992);
nor UO_370 (O_370,N_2958,N_2981);
nand UO_371 (O_371,N_2979,N_2951);
nand UO_372 (O_372,N_2984,N_2986);
nand UO_373 (O_373,N_2956,N_2954);
nand UO_374 (O_374,N_2981,N_2962);
xor UO_375 (O_375,N_2959,N_2997);
and UO_376 (O_376,N_2981,N_2984);
nand UO_377 (O_377,N_2952,N_2951);
and UO_378 (O_378,N_2967,N_2990);
nor UO_379 (O_379,N_2990,N_2956);
or UO_380 (O_380,N_2993,N_2992);
nor UO_381 (O_381,N_2998,N_2996);
nand UO_382 (O_382,N_2985,N_2989);
and UO_383 (O_383,N_2960,N_2958);
nand UO_384 (O_384,N_2982,N_2988);
or UO_385 (O_385,N_2963,N_2997);
and UO_386 (O_386,N_2993,N_2973);
and UO_387 (O_387,N_2967,N_2972);
nand UO_388 (O_388,N_2969,N_2961);
and UO_389 (O_389,N_2976,N_2971);
nand UO_390 (O_390,N_2951,N_2980);
nor UO_391 (O_391,N_2981,N_2954);
and UO_392 (O_392,N_2977,N_2992);
and UO_393 (O_393,N_2993,N_2970);
nand UO_394 (O_394,N_2977,N_2950);
and UO_395 (O_395,N_2990,N_2979);
nand UO_396 (O_396,N_2956,N_2998);
or UO_397 (O_397,N_2964,N_2954);
nor UO_398 (O_398,N_2953,N_2977);
nand UO_399 (O_399,N_2987,N_2956);
or UO_400 (O_400,N_2971,N_2987);
nor UO_401 (O_401,N_2950,N_2999);
and UO_402 (O_402,N_2955,N_2970);
and UO_403 (O_403,N_2986,N_2997);
nor UO_404 (O_404,N_2966,N_2962);
and UO_405 (O_405,N_2997,N_2985);
and UO_406 (O_406,N_2993,N_2975);
nor UO_407 (O_407,N_2975,N_2955);
nor UO_408 (O_408,N_2951,N_2971);
nor UO_409 (O_409,N_2994,N_2978);
or UO_410 (O_410,N_2963,N_2999);
nand UO_411 (O_411,N_2960,N_2999);
and UO_412 (O_412,N_2991,N_2990);
nor UO_413 (O_413,N_2957,N_2963);
and UO_414 (O_414,N_2976,N_2974);
or UO_415 (O_415,N_2969,N_2991);
and UO_416 (O_416,N_2995,N_2971);
nor UO_417 (O_417,N_2958,N_2990);
or UO_418 (O_418,N_2964,N_2976);
nand UO_419 (O_419,N_2961,N_2985);
nor UO_420 (O_420,N_2972,N_2993);
nand UO_421 (O_421,N_2997,N_2953);
and UO_422 (O_422,N_2956,N_2995);
or UO_423 (O_423,N_2965,N_2969);
and UO_424 (O_424,N_2966,N_2950);
or UO_425 (O_425,N_2992,N_2966);
nand UO_426 (O_426,N_2972,N_2991);
nand UO_427 (O_427,N_2956,N_2983);
or UO_428 (O_428,N_2967,N_2966);
and UO_429 (O_429,N_2958,N_2964);
xor UO_430 (O_430,N_2959,N_2995);
nor UO_431 (O_431,N_2985,N_2992);
and UO_432 (O_432,N_2989,N_2952);
and UO_433 (O_433,N_2970,N_2968);
and UO_434 (O_434,N_2979,N_2989);
and UO_435 (O_435,N_2951,N_2987);
and UO_436 (O_436,N_2992,N_2958);
and UO_437 (O_437,N_2992,N_2962);
or UO_438 (O_438,N_2973,N_2992);
nor UO_439 (O_439,N_2960,N_2987);
or UO_440 (O_440,N_2995,N_2950);
nor UO_441 (O_441,N_2969,N_2954);
or UO_442 (O_442,N_2955,N_2964);
nor UO_443 (O_443,N_2953,N_2981);
or UO_444 (O_444,N_2967,N_2961);
nand UO_445 (O_445,N_2987,N_2964);
or UO_446 (O_446,N_2978,N_2977);
nand UO_447 (O_447,N_2993,N_2965);
nor UO_448 (O_448,N_2970,N_2974);
or UO_449 (O_449,N_2950,N_2973);
xor UO_450 (O_450,N_2998,N_2981);
nand UO_451 (O_451,N_2987,N_2989);
nand UO_452 (O_452,N_2995,N_2973);
or UO_453 (O_453,N_2993,N_2962);
or UO_454 (O_454,N_2971,N_2980);
or UO_455 (O_455,N_2959,N_2967);
and UO_456 (O_456,N_2990,N_2970);
nor UO_457 (O_457,N_2971,N_2970);
and UO_458 (O_458,N_2988,N_2970);
and UO_459 (O_459,N_2950,N_2984);
nor UO_460 (O_460,N_2999,N_2994);
nand UO_461 (O_461,N_2953,N_2991);
nor UO_462 (O_462,N_2978,N_2996);
nand UO_463 (O_463,N_2975,N_2968);
and UO_464 (O_464,N_2990,N_2968);
or UO_465 (O_465,N_2990,N_2993);
nand UO_466 (O_466,N_2978,N_2975);
nor UO_467 (O_467,N_2984,N_2992);
nor UO_468 (O_468,N_2999,N_2955);
nor UO_469 (O_469,N_2976,N_2992);
or UO_470 (O_470,N_2953,N_2985);
nand UO_471 (O_471,N_2970,N_2962);
nor UO_472 (O_472,N_2953,N_2968);
or UO_473 (O_473,N_2985,N_2951);
nand UO_474 (O_474,N_2991,N_2968);
nor UO_475 (O_475,N_2969,N_2951);
nor UO_476 (O_476,N_2996,N_2965);
nor UO_477 (O_477,N_2999,N_2967);
nand UO_478 (O_478,N_2977,N_2955);
or UO_479 (O_479,N_2955,N_2950);
nor UO_480 (O_480,N_2975,N_2972);
and UO_481 (O_481,N_2958,N_2979);
nand UO_482 (O_482,N_2962,N_2965);
nor UO_483 (O_483,N_2967,N_2998);
nor UO_484 (O_484,N_2959,N_2981);
nand UO_485 (O_485,N_2990,N_2972);
or UO_486 (O_486,N_2981,N_2985);
nor UO_487 (O_487,N_2998,N_2980);
or UO_488 (O_488,N_2967,N_2983);
and UO_489 (O_489,N_2988,N_2973);
nand UO_490 (O_490,N_2965,N_2978);
and UO_491 (O_491,N_2992,N_2968);
nor UO_492 (O_492,N_2976,N_2994);
nand UO_493 (O_493,N_2992,N_2970);
and UO_494 (O_494,N_2999,N_2979);
nor UO_495 (O_495,N_2951,N_2975);
nor UO_496 (O_496,N_2999,N_2966);
nor UO_497 (O_497,N_2991,N_2955);
nor UO_498 (O_498,N_2957,N_2962);
nor UO_499 (O_499,N_2965,N_2987);
endmodule