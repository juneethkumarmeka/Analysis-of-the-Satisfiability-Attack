module basic_500_3000_500_15_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_111,In_57);
or U1 (N_1,In_375,In_62);
and U2 (N_2,In_225,In_130);
and U3 (N_3,In_455,In_96);
nand U4 (N_4,In_429,In_388);
xor U5 (N_5,In_401,In_14);
nand U6 (N_6,In_410,In_485);
or U7 (N_7,In_12,In_55);
and U8 (N_8,In_241,In_149);
nand U9 (N_9,In_293,In_174);
nand U10 (N_10,In_324,In_93);
and U11 (N_11,In_143,In_328);
nor U12 (N_12,In_80,In_396);
or U13 (N_13,In_307,In_76);
or U14 (N_14,In_342,In_22);
xnor U15 (N_15,In_56,In_374);
nand U16 (N_16,In_382,In_197);
nand U17 (N_17,In_425,In_196);
or U18 (N_18,In_448,In_7);
and U19 (N_19,In_191,In_32);
or U20 (N_20,In_424,In_415);
nand U21 (N_21,In_418,In_101);
and U22 (N_22,In_217,In_372);
and U23 (N_23,In_239,In_150);
or U24 (N_24,In_236,In_271);
nand U25 (N_25,In_257,In_341);
nor U26 (N_26,In_330,In_118);
nor U27 (N_27,In_145,In_497);
and U28 (N_28,In_19,In_454);
and U29 (N_29,In_490,In_30);
or U30 (N_30,In_253,In_313);
and U31 (N_31,In_232,In_492);
or U32 (N_32,In_365,In_302);
and U33 (N_33,In_488,In_254);
nor U34 (N_34,In_376,In_121);
and U35 (N_35,In_384,In_157);
and U36 (N_36,In_228,In_499);
nor U37 (N_37,In_269,In_61);
nor U38 (N_38,In_114,In_468);
and U39 (N_39,In_29,In_144);
or U40 (N_40,In_479,In_434);
nand U41 (N_41,In_360,In_91);
nand U42 (N_42,In_36,In_49);
nor U43 (N_43,In_39,In_286);
nor U44 (N_44,In_176,In_266);
nor U45 (N_45,In_216,In_465);
and U46 (N_46,In_427,In_387);
nand U47 (N_47,In_426,In_474);
and U48 (N_48,In_24,In_278);
or U49 (N_49,In_208,In_167);
nand U50 (N_50,In_87,In_346);
and U51 (N_51,In_211,In_132);
nand U52 (N_52,In_243,In_270);
and U53 (N_53,In_475,In_206);
and U54 (N_54,In_212,In_326);
nor U55 (N_55,In_136,In_102);
nand U56 (N_56,In_173,In_398);
nand U57 (N_57,In_294,In_332);
and U58 (N_58,In_100,In_158);
and U59 (N_59,In_430,In_357);
nor U60 (N_60,In_73,In_127);
nand U61 (N_61,In_117,In_83);
nand U62 (N_62,In_33,In_95);
or U63 (N_63,In_94,In_9);
nand U64 (N_64,In_390,In_188);
nand U65 (N_65,In_477,In_155);
and U66 (N_66,In_171,In_120);
or U67 (N_67,In_399,In_289);
nand U68 (N_68,In_116,In_381);
nand U69 (N_69,In_353,In_43);
and U70 (N_70,In_284,In_123);
nor U71 (N_71,In_316,In_133);
nor U72 (N_72,In_135,In_414);
and U73 (N_73,In_77,In_223);
or U74 (N_74,In_476,In_105);
nor U75 (N_75,In_323,In_125);
or U76 (N_76,In_69,In_457);
nor U77 (N_77,In_162,In_305);
xor U78 (N_78,In_233,In_129);
or U79 (N_79,In_273,In_74);
or U80 (N_80,In_296,In_459);
and U81 (N_81,In_4,In_470);
nand U82 (N_82,In_442,In_297);
or U83 (N_83,In_291,In_147);
nor U84 (N_84,In_168,In_53);
nor U85 (N_85,In_276,In_338);
nand U86 (N_86,In_215,In_438);
nor U87 (N_87,In_137,In_109);
or U88 (N_88,In_199,In_303);
nand U89 (N_89,In_301,In_25);
nand U90 (N_90,In_447,In_169);
and U91 (N_91,In_140,In_52);
nor U92 (N_92,In_200,In_90);
nand U93 (N_93,In_264,In_50);
nor U94 (N_94,In_213,In_54);
nor U95 (N_95,In_412,In_146);
or U96 (N_96,In_138,In_484);
or U97 (N_97,In_195,In_107);
and U98 (N_98,In_15,In_234);
nor U99 (N_99,In_428,In_26);
and U100 (N_100,In_325,In_126);
nand U101 (N_101,In_115,In_249);
nand U102 (N_102,In_343,In_192);
and U103 (N_103,In_178,In_10);
nand U104 (N_104,In_203,In_153);
and U105 (N_105,In_344,In_462);
nor U106 (N_106,In_395,In_481);
and U107 (N_107,In_432,In_31);
nor U108 (N_108,In_373,In_42);
and U109 (N_109,In_315,In_131);
and U110 (N_110,In_445,In_306);
and U111 (N_111,In_159,In_184);
nor U112 (N_112,In_435,In_416);
or U113 (N_113,In_16,In_44);
or U114 (N_114,In_423,In_108);
nand U115 (N_115,In_461,In_163);
and U116 (N_116,In_279,In_71);
nor U117 (N_117,In_437,In_106);
nand U118 (N_118,In_245,In_321);
and U119 (N_119,In_274,In_392);
or U120 (N_120,In_230,In_210);
nand U121 (N_121,In_84,In_371);
nor U122 (N_122,In_48,In_128);
nand U123 (N_123,In_487,In_363);
and U124 (N_124,In_281,In_359);
nand U125 (N_125,In_397,In_65);
nand U126 (N_126,In_6,In_17);
nand U127 (N_127,In_472,In_112);
and U128 (N_128,In_367,In_406);
nand U129 (N_129,In_496,In_408);
or U130 (N_130,In_483,In_463);
or U131 (N_131,In_443,In_41);
nand U132 (N_132,In_165,In_175);
nand U133 (N_133,In_142,In_421);
or U134 (N_134,In_322,In_259);
nor U135 (N_135,In_329,In_187);
or U136 (N_136,In_304,In_263);
or U137 (N_137,In_104,In_214);
nand U138 (N_138,In_11,In_393);
and U139 (N_139,In_5,In_8);
nand U140 (N_140,In_119,In_161);
nand U141 (N_141,In_280,In_309);
nand U142 (N_142,In_402,In_282);
nand U143 (N_143,In_453,In_334);
nor U144 (N_144,In_170,In_231);
nand U145 (N_145,In_413,In_179);
nand U146 (N_146,In_275,In_478);
nand U147 (N_147,In_335,In_495);
nand U148 (N_148,In_154,In_333);
and U149 (N_149,In_164,In_141);
nand U150 (N_150,In_72,In_452);
nor U151 (N_151,In_378,In_417);
nand U152 (N_152,In_407,In_183);
nand U153 (N_153,In_201,In_82);
or U154 (N_154,In_21,In_347);
nand U155 (N_155,In_218,In_222);
and U156 (N_156,In_238,In_489);
and U157 (N_157,In_419,In_411);
nor U158 (N_158,In_229,In_148);
or U159 (N_159,In_400,In_268);
nor U160 (N_160,In_366,In_277);
nand U161 (N_161,In_193,In_156);
nand U162 (N_162,In_308,In_172);
or U163 (N_163,In_103,In_262);
and U164 (N_164,In_242,In_422);
nand U165 (N_165,In_207,In_63);
and U166 (N_166,In_471,In_311);
nand U167 (N_167,In_13,In_272);
and U168 (N_168,In_202,In_295);
nand U169 (N_169,In_290,In_35);
nand U170 (N_170,In_405,In_458);
or U171 (N_171,In_85,In_247);
nor U172 (N_172,In_113,In_404);
nand U173 (N_173,In_38,In_166);
and U174 (N_174,In_244,In_337);
nand U175 (N_175,In_23,In_385);
nor U176 (N_176,In_354,In_75);
nor U177 (N_177,In_473,In_2);
nand U178 (N_178,In_287,In_377);
or U179 (N_179,In_285,In_292);
nand U180 (N_180,In_358,In_441);
or U181 (N_181,In_185,In_312);
nor U182 (N_182,In_433,In_391);
nor U183 (N_183,In_498,In_383);
or U184 (N_184,In_99,In_181);
nand U185 (N_185,In_480,In_491);
nand U186 (N_186,In_124,In_18);
nor U187 (N_187,In_482,In_98);
nor U188 (N_188,In_320,In_389);
and U189 (N_189,In_70,In_160);
or U190 (N_190,In_37,In_251);
or U191 (N_191,In_352,In_370);
and U192 (N_192,In_318,In_194);
nand U193 (N_193,In_394,In_51);
nor U194 (N_194,In_369,In_331);
and U195 (N_195,In_189,In_226);
and U196 (N_196,In_227,In_224);
nand U197 (N_197,In_351,In_340);
nand U198 (N_198,In_209,In_420);
nand U199 (N_199,In_299,In_205);
or U200 (N_200,N_4,N_186);
or U201 (N_201,N_94,N_90);
nand U202 (N_202,In_314,N_191);
nand U203 (N_203,N_26,N_55);
nand U204 (N_204,N_59,In_466);
and U205 (N_205,In_339,In_350);
nand U206 (N_206,In_3,N_167);
nand U207 (N_207,N_79,In_221);
nor U208 (N_208,In_349,N_169);
and U209 (N_209,N_115,N_76);
nand U210 (N_210,N_80,N_149);
or U211 (N_211,In_258,In_252);
or U212 (N_212,N_97,N_91);
nor U213 (N_213,N_96,N_144);
and U214 (N_214,In_494,N_38);
nor U215 (N_215,N_151,In_368);
nor U216 (N_216,In_190,N_28);
nand U217 (N_217,In_380,N_163);
nor U218 (N_218,In_486,In_67);
or U219 (N_219,N_110,N_177);
nor U220 (N_220,N_48,N_143);
nand U221 (N_221,N_39,N_146);
and U222 (N_222,In_28,N_182);
xor U223 (N_223,N_20,N_180);
nand U224 (N_224,N_187,N_137);
and U225 (N_225,N_195,N_74);
nor U226 (N_226,N_10,N_71);
nor U227 (N_227,N_17,In_78);
nor U228 (N_228,N_21,In_220);
nand U229 (N_229,N_173,N_68);
nand U230 (N_230,In_255,In_310);
and U231 (N_231,In_355,N_166);
xnor U232 (N_232,N_148,In_451);
or U233 (N_233,N_155,In_182);
nand U234 (N_234,N_120,N_78);
or U235 (N_235,In_110,N_69);
and U236 (N_236,N_86,N_136);
nand U237 (N_237,N_46,N_14);
and U238 (N_238,In_450,In_345);
or U239 (N_239,N_70,N_108);
nand U240 (N_240,N_112,N_124);
or U241 (N_241,In_469,N_84);
nand U242 (N_242,N_154,In_386);
and U243 (N_243,N_13,In_265);
nor U244 (N_244,N_7,N_25);
or U245 (N_245,In_409,In_464);
nor U246 (N_246,N_123,N_36);
and U247 (N_247,N_42,In_81);
nand U248 (N_248,In_40,N_85);
nor U249 (N_249,N_122,In_139);
and U250 (N_250,N_98,In_319);
nand U251 (N_251,In_267,N_116);
nor U252 (N_252,In_336,N_160);
and U253 (N_253,In_79,N_88);
or U254 (N_254,N_50,N_53);
or U255 (N_255,In_59,N_118);
and U256 (N_256,N_31,In_248);
or U257 (N_257,N_60,N_52);
and U258 (N_258,In_356,N_142);
or U259 (N_259,N_117,N_125);
nor U260 (N_260,In_219,N_95);
nor U261 (N_261,N_72,N_157);
or U262 (N_262,In_237,N_127);
nand U263 (N_263,N_192,N_105);
nor U264 (N_264,N_6,In_86);
or U265 (N_265,In_403,N_67);
nand U266 (N_266,N_147,N_24);
nand U267 (N_267,In_449,N_18);
nor U268 (N_268,N_193,N_41);
and U269 (N_269,In_177,N_83);
and U270 (N_270,N_73,N_128);
or U271 (N_271,N_61,N_129);
nand U272 (N_272,N_23,N_45);
nand U273 (N_273,N_171,In_68);
and U274 (N_274,In_327,N_111);
nor U275 (N_275,N_27,N_102);
nand U276 (N_276,N_176,In_446);
and U277 (N_277,N_178,In_246);
or U278 (N_278,In_436,N_133);
and U279 (N_279,N_16,N_196);
or U280 (N_280,N_141,In_235);
nor U281 (N_281,N_185,N_77);
nand U282 (N_282,In_456,In_467);
and U283 (N_283,N_175,N_121);
nand U284 (N_284,In_261,N_37);
or U285 (N_285,N_64,N_92);
or U286 (N_286,In_64,N_198);
nand U287 (N_287,N_170,N_51);
nor U288 (N_288,N_140,N_19);
nor U289 (N_289,N_58,N_183);
or U290 (N_290,In_444,In_122);
nor U291 (N_291,N_103,In_283);
nand U292 (N_292,In_66,N_32);
nor U293 (N_293,N_75,N_150);
and U294 (N_294,N_189,N_82);
nor U295 (N_295,N_33,In_20);
nor U296 (N_296,In_348,N_43);
nor U297 (N_297,In_89,N_22);
or U298 (N_298,N_47,In_431);
nand U299 (N_299,N_152,N_107);
nand U300 (N_300,In_151,N_165);
nor U301 (N_301,N_126,N_30);
nand U302 (N_302,N_139,N_159);
nor U303 (N_303,N_138,N_145);
or U304 (N_304,In_45,N_3);
nor U305 (N_305,In_493,N_172);
nor U306 (N_306,In_379,In_298);
and U307 (N_307,N_62,In_186);
and U308 (N_308,In_364,N_100);
or U309 (N_309,N_131,In_60);
and U310 (N_310,N_106,N_56);
nor U311 (N_311,N_99,N_164);
and U312 (N_312,In_0,N_190);
xor U313 (N_313,In_361,In_460);
or U314 (N_314,N_66,N_153);
and U315 (N_315,N_65,N_63);
nand U316 (N_316,N_134,N_54);
nand U317 (N_317,N_132,In_97);
and U318 (N_318,In_47,N_135);
nand U319 (N_319,In_300,In_440);
or U320 (N_320,N_109,In_362);
nand U321 (N_321,In_260,N_194);
and U322 (N_322,In_288,N_130);
nand U323 (N_323,N_161,N_188);
nand U324 (N_324,N_11,N_113);
and U325 (N_325,N_162,N_168);
nor U326 (N_326,In_88,N_104);
nand U327 (N_327,In_152,In_92);
nor U328 (N_328,In_134,In_250);
and U329 (N_329,N_35,N_184);
or U330 (N_330,N_49,N_87);
nand U331 (N_331,In_198,In_180);
nand U332 (N_332,N_9,In_256);
nor U333 (N_333,N_174,In_34);
nor U334 (N_334,N_158,N_57);
or U335 (N_335,N_114,In_240);
nor U336 (N_336,In_204,N_40);
nor U337 (N_337,In_317,N_93);
nor U338 (N_338,N_8,N_81);
nor U339 (N_339,In_58,In_27);
nand U340 (N_340,In_46,N_101);
and U341 (N_341,N_34,N_2);
and U342 (N_342,N_0,N_44);
or U343 (N_343,In_439,N_156);
and U344 (N_344,N_181,N_89);
and U345 (N_345,N_15,N_12);
nor U346 (N_346,N_119,N_29);
nand U347 (N_347,N_1,N_199);
nand U348 (N_348,In_1,N_197);
or U349 (N_349,N_179,N_5);
or U350 (N_350,N_183,N_48);
nand U351 (N_351,N_144,In_464);
nand U352 (N_352,N_140,N_125);
or U353 (N_353,N_25,N_67);
nand U354 (N_354,N_112,N_192);
or U355 (N_355,N_16,N_199);
or U356 (N_356,N_115,In_456);
and U357 (N_357,N_96,N_164);
and U358 (N_358,In_58,N_135);
nand U359 (N_359,N_144,In_237);
nand U360 (N_360,N_192,N_4);
nand U361 (N_361,N_21,N_74);
nor U362 (N_362,N_107,N_110);
or U363 (N_363,In_0,N_146);
or U364 (N_364,In_60,N_144);
nor U365 (N_365,In_3,N_164);
or U366 (N_366,In_456,N_42);
and U367 (N_367,N_22,N_35);
nand U368 (N_368,N_102,In_88);
or U369 (N_369,N_96,N_0);
nor U370 (N_370,In_27,N_144);
and U371 (N_371,In_288,N_2);
or U372 (N_372,N_190,N_113);
or U373 (N_373,In_450,N_185);
and U374 (N_374,N_42,In_78);
nand U375 (N_375,N_21,In_68);
and U376 (N_376,N_72,N_175);
and U377 (N_377,In_467,N_122);
and U378 (N_378,In_260,In_248);
nand U379 (N_379,In_345,N_41);
or U380 (N_380,N_130,N_148);
or U381 (N_381,In_446,N_85);
and U382 (N_382,N_168,N_14);
or U383 (N_383,N_148,N_34);
or U384 (N_384,In_368,N_172);
and U385 (N_385,In_380,N_89);
nand U386 (N_386,In_134,N_62);
or U387 (N_387,In_317,N_100);
and U388 (N_388,N_158,N_194);
and U389 (N_389,N_90,N_74);
nand U390 (N_390,N_10,In_248);
or U391 (N_391,In_327,In_88);
nor U392 (N_392,N_31,N_25);
or U393 (N_393,N_105,N_117);
and U394 (N_394,N_32,N_118);
or U395 (N_395,N_162,N_58);
or U396 (N_396,In_469,In_494);
and U397 (N_397,N_3,In_409);
or U398 (N_398,In_3,N_162);
nand U399 (N_399,In_348,N_119);
or U400 (N_400,N_240,N_251);
and U401 (N_401,N_282,N_245);
or U402 (N_402,N_369,N_288);
nor U403 (N_403,N_330,N_265);
nor U404 (N_404,N_278,N_225);
nor U405 (N_405,N_283,N_319);
nand U406 (N_406,N_348,N_289);
or U407 (N_407,N_274,N_394);
and U408 (N_408,N_391,N_386);
nand U409 (N_409,N_370,N_211);
and U410 (N_410,N_349,N_350);
and U411 (N_411,N_229,N_228);
nor U412 (N_412,N_208,N_373);
and U413 (N_413,N_300,N_247);
or U414 (N_414,N_261,N_295);
nor U415 (N_415,N_390,N_396);
nand U416 (N_416,N_382,N_316);
nand U417 (N_417,N_205,N_259);
xnor U418 (N_418,N_346,N_226);
nor U419 (N_419,N_356,N_358);
and U420 (N_420,N_341,N_262);
nand U421 (N_421,N_311,N_351);
nand U422 (N_422,N_270,N_306);
nor U423 (N_423,N_204,N_287);
nand U424 (N_424,N_244,N_257);
nand U425 (N_425,N_273,N_359);
nor U426 (N_426,N_281,N_398);
or U427 (N_427,N_277,N_243);
or U428 (N_428,N_347,N_333);
nor U429 (N_429,N_286,N_294);
nand U430 (N_430,N_342,N_309);
nand U431 (N_431,N_354,N_301);
nor U432 (N_432,N_332,N_293);
nand U433 (N_433,N_307,N_399);
and U434 (N_434,N_305,N_378);
and U435 (N_435,N_355,N_233);
and U436 (N_436,N_320,N_336);
and U437 (N_437,N_365,N_387);
nor U438 (N_438,N_222,N_337);
or U439 (N_439,N_328,N_318);
and U440 (N_440,N_214,N_321);
nor U441 (N_441,N_324,N_224);
nor U442 (N_442,N_368,N_326);
nand U443 (N_443,N_323,N_264);
nand U444 (N_444,N_327,N_302);
and U445 (N_445,N_375,N_303);
or U446 (N_446,N_280,N_260);
or U447 (N_447,N_297,N_212);
nand U448 (N_448,N_380,N_381);
nand U449 (N_449,N_232,N_344);
nand U450 (N_450,N_213,N_361);
nor U451 (N_451,N_299,N_235);
nor U452 (N_452,N_236,N_360);
and U453 (N_453,N_338,N_219);
nand U454 (N_454,N_221,N_241);
and U455 (N_455,N_252,N_268);
or U456 (N_456,N_366,N_317);
or U457 (N_457,N_395,N_230);
nor U458 (N_458,N_335,N_239);
nand U459 (N_459,N_308,N_379);
or U460 (N_460,N_352,N_314);
nor U461 (N_461,N_371,N_315);
nand U462 (N_462,N_209,N_364);
nor U463 (N_463,N_322,N_267);
nor U464 (N_464,N_384,N_217);
or U465 (N_465,N_279,N_246);
and U466 (N_466,N_210,N_292);
and U467 (N_467,N_377,N_250);
nand U468 (N_468,N_353,N_340);
or U469 (N_469,N_263,N_266);
and U470 (N_470,N_272,N_220);
nand U471 (N_471,N_313,N_256);
and U472 (N_472,N_372,N_201);
nor U473 (N_473,N_255,N_276);
and U474 (N_474,N_339,N_290);
or U475 (N_475,N_393,N_234);
and U476 (N_476,N_218,N_357);
or U477 (N_477,N_334,N_345);
or U478 (N_478,N_227,N_362);
nor U479 (N_479,N_253,N_258);
nor U480 (N_480,N_296,N_254);
nand U481 (N_481,N_376,N_248);
and U482 (N_482,N_374,N_388);
nor U483 (N_483,N_223,N_310);
or U484 (N_484,N_284,N_237);
nor U485 (N_485,N_206,N_200);
nor U486 (N_486,N_249,N_304);
and U487 (N_487,N_363,N_271);
and U488 (N_488,N_275,N_397);
or U489 (N_489,N_203,N_343);
and U490 (N_490,N_216,N_285);
and U491 (N_491,N_291,N_238);
nand U492 (N_492,N_325,N_392);
nand U493 (N_493,N_298,N_207);
nor U494 (N_494,N_385,N_367);
or U495 (N_495,N_331,N_202);
and U496 (N_496,N_383,N_329);
or U497 (N_497,N_269,N_312);
nand U498 (N_498,N_389,N_215);
or U499 (N_499,N_242,N_231);
and U500 (N_500,N_274,N_337);
and U501 (N_501,N_398,N_308);
nor U502 (N_502,N_321,N_336);
and U503 (N_503,N_295,N_342);
nand U504 (N_504,N_263,N_244);
and U505 (N_505,N_378,N_233);
nand U506 (N_506,N_245,N_263);
or U507 (N_507,N_203,N_337);
nor U508 (N_508,N_263,N_226);
nand U509 (N_509,N_366,N_364);
or U510 (N_510,N_367,N_231);
nor U511 (N_511,N_307,N_250);
and U512 (N_512,N_324,N_281);
nand U513 (N_513,N_236,N_314);
and U514 (N_514,N_218,N_368);
nand U515 (N_515,N_268,N_397);
nor U516 (N_516,N_269,N_355);
nor U517 (N_517,N_334,N_201);
or U518 (N_518,N_216,N_246);
or U519 (N_519,N_254,N_311);
and U520 (N_520,N_311,N_346);
and U521 (N_521,N_247,N_254);
nand U522 (N_522,N_354,N_306);
and U523 (N_523,N_285,N_247);
nand U524 (N_524,N_206,N_246);
nand U525 (N_525,N_355,N_286);
xor U526 (N_526,N_271,N_352);
or U527 (N_527,N_288,N_323);
and U528 (N_528,N_309,N_313);
or U529 (N_529,N_258,N_392);
or U530 (N_530,N_255,N_295);
nand U531 (N_531,N_292,N_296);
and U532 (N_532,N_229,N_299);
and U533 (N_533,N_346,N_200);
and U534 (N_534,N_368,N_329);
nor U535 (N_535,N_365,N_273);
and U536 (N_536,N_212,N_332);
and U537 (N_537,N_217,N_243);
or U538 (N_538,N_321,N_257);
or U539 (N_539,N_247,N_346);
or U540 (N_540,N_200,N_271);
nand U541 (N_541,N_222,N_366);
and U542 (N_542,N_303,N_267);
nand U543 (N_543,N_333,N_368);
and U544 (N_544,N_201,N_271);
nand U545 (N_545,N_303,N_357);
or U546 (N_546,N_283,N_368);
nor U547 (N_547,N_386,N_263);
nor U548 (N_548,N_318,N_267);
nand U549 (N_549,N_207,N_381);
nor U550 (N_550,N_276,N_308);
nor U551 (N_551,N_386,N_332);
and U552 (N_552,N_310,N_342);
nor U553 (N_553,N_289,N_270);
xnor U554 (N_554,N_321,N_352);
or U555 (N_555,N_287,N_295);
nor U556 (N_556,N_235,N_262);
nand U557 (N_557,N_398,N_220);
nand U558 (N_558,N_205,N_395);
and U559 (N_559,N_303,N_392);
or U560 (N_560,N_223,N_358);
nor U561 (N_561,N_234,N_297);
and U562 (N_562,N_212,N_260);
nand U563 (N_563,N_388,N_342);
nor U564 (N_564,N_293,N_322);
or U565 (N_565,N_200,N_337);
nand U566 (N_566,N_222,N_350);
and U567 (N_567,N_201,N_294);
and U568 (N_568,N_292,N_354);
nor U569 (N_569,N_303,N_322);
or U570 (N_570,N_249,N_297);
nor U571 (N_571,N_316,N_277);
nand U572 (N_572,N_224,N_307);
and U573 (N_573,N_277,N_343);
nor U574 (N_574,N_340,N_364);
or U575 (N_575,N_293,N_295);
or U576 (N_576,N_296,N_206);
and U577 (N_577,N_309,N_238);
nor U578 (N_578,N_215,N_262);
and U579 (N_579,N_389,N_347);
or U580 (N_580,N_211,N_235);
nand U581 (N_581,N_346,N_336);
or U582 (N_582,N_332,N_263);
nand U583 (N_583,N_363,N_366);
nand U584 (N_584,N_201,N_303);
nor U585 (N_585,N_392,N_270);
and U586 (N_586,N_258,N_296);
or U587 (N_587,N_345,N_224);
nor U588 (N_588,N_394,N_206);
and U589 (N_589,N_300,N_396);
nand U590 (N_590,N_273,N_232);
nor U591 (N_591,N_374,N_324);
nor U592 (N_592,N_305,N_357);
nand U593 (N_593,N_221,N_303);
nand U594 (N_594,N_224,N_213);
nand U595 (N_595,N_378,N_224);
and U596 (N_596,N_361,N_383);
or U597 (N_597,N_384,N_275);
nand U598 (N_598,N_293,N_221);
and U599 (N_599,N_374,N_358);
or U600 (N_600,N_591,N_428);
or U601 (N_601,N_485,N_549);
or U602 (N_602,N_460,N_580);
or U603 (N_603,N_444,N_496);
or U604 (N_604,N_478,N_400);
and U605 (N_605,N_585,N_482);
or U606 (N_606,N_524,N_554);
nor U607 (N_607,N_424,N_583);
nand U608 (N_608,N_414,N_555);
nor U609 (N_609,N_582,N_465);
nand U610 (N_610,N_566,N_476);
and U611 (N_611,N_479,N_432);
or U612 (N_612,N_522,N_550);
or U613 (N_613,N_408,N_407);
and U614 (N_614,N_520,N_447);
and U615 (N_615,N_545,N_598);
nand U616 (N_616,N_527,N_574);
or U617 (N_617,N_501,N_544);
or U618 (N_618,N_551,N_421);
or U619 (N_619,N_588,N_516);
nand U620 (N_620,N_471,N_584);
nand U621 (N_621,N_451,N_487);
nor U622 (N_622,N_434,N_406);
nand U623 (N_623,N_529,N_419);
and U624 (N_624,N_436,N_514);
and U625 (N_625,N_570,N_491);
and U626 (N_626,N_538,N_474);
or U627 (N_627,N_472,N_578);
or U628 (N_628,N_416,N_542);
nor U629 (N_629,N_457,N_442);
nor U630 (N_630,N_531,N_521);
nand U631 (N_631,N_528,N_559);
and U632 (N_632,N_553,N_563);
and U633 (N_633,N_448,N_467);
nand U634 (N_634,N_470,N_540);
nor U635 (N_635,N_493,N_483);
or U636 (N_636,N_430,N_511);
nand U637 (N_637,N_537,N_552);
and U638 (N_638,N_415,N_426);
or U639 (N_639,N_423,N_492);
and U640 (N_640,N_513,N_490);
and U641 (N_641,N_469,N_562);
and U642 (N_642,N_402,N_463);
and U643 (N_643,N_569,N_548);
and U644 (N_644,N_568,N_523);
nand U645 (N_645,N_572,N_567);
and U646 (N_646,N_449,N_495);
or U647 (N_647,N_507,N_401);
or U648 (N_648,N_577,N_592);
or U649 (N_649,N_500,N_453);
and U650 (N_650,N_440,N_435);
and U651 (N_651,N_508,N_509);
nor U652 (N_652,N_445,N_475);
nor U653 (N_653,N_404,N_573);
nand U654 (N_654,N_437,N_502);
nor U655 (N_655,N_536,N_427);
or U656 (N_656,N_473,N_441);
nor U657 (N_657,N_481,N_593);
and U658 (N_658,N_547,N_539);
and U659 (N_659,N_543,N_599);
and U660 (N_660,N_546,N_576);
nand U661 (N_661,N_497,N_403);
nor U662 (N_662,N_561,N_462);
nor U663 (N_663,N_597,N_564);
and U664 (N_664,N_412,N_594);
nor U665 (N_665,N_534,N_459);
nor U666 (N_666,N_420,N_504);
nand U667 (N_667,N_590,N_480);
and U668 (N_668,N_499,N_418);
nor U669 (N_669,N_443,N_595);
and U670 (N_670,N_517,N_422);
and U671 (N_671,N_503,N_532);
nand U672 (N_672,N_586,N_596);
nor U673 (N_673,N_587,N_439);
nand U674 (N_674,N_454,N_530);
and U675 (N_675,N_510,N_425);
nand U676 (N_676,N_515,N_575);
or U677 (N_677,N_484,N_494);
and U678 (N_678,N_505,N_488);
nand U679 (N_679,N_533,N_535);
and U680 (N_680,N_519,N_405);
nand U681 (N_681,N_431,N_579);
nor U682 (N_682,N_571,N_433);
nand U683 (N_683,N_461,N_446);
nand U684 (N_684,N_411,N_455);
nand U685 (N_685,N_506,N_438);
nor U686 (N_686,N_489,N_468);
and U687 (N_687,N_486,N_409);
or U688 (N_688,N_429,N_498);
nand U689 (N_689,N_556,N_477);
nor U690 (N_690,N_413,N_417);
and U691 (N_691,N_466,N_557);
and U692 (N_692,N_518,N_456);
and U693 (N_693,N_558,N_565);
nor U694 (N_694,N_410,N_581);
and U695 (N_695,N_525,N_512);
nor U696 (N_696,N_452,N_464);
and U697 (N_697,N_450,N_458);
or U698 (N_698,N_541,N_589);
nor U699 (N_699,N_526,N_560);
and U700 (N_700,N_429,N_477);
nor U701 (N_701,N_553,N_518);
nand U702 (N_702,N_590,N_533);
nor U703 (N_703,N_408,N_518);
nor U704 (N_704,N_428,N_413);
and U705 (N_705,N_536,N_470);
or U706 (N_706,N_477,N_410);
and U707 (N_707,N_558,N_562);
or U708 (N_708,N_563,N_570);
nand U709 (N_709,N_582,N_587);
nor U710 (N_710,N_545,N_584);
and U711 (N_711,N_499,N_474);
or U712 (N_712,N_487,N_446);
nor U713 (N_713,N_447,N_537);
nor U714 (N_714,N_464,N_590);
nor U715 (N_715,N_542,N_471);
nor U716 (N_716,N_541,N_511);
or U717 (N_717,N_581,N_528);
nor U718 (N_718,N_589,N_566);
or U719 (N_719,N_556,N_517);
nand U720 (N_720,N_539,N_577);
nor U721 (N_721,N_434,N_568);
nand U722 (N_722,N_422,N_414);
nand U723 (N_723,N_576,N_431);
or U724 (N_724,N_461,N_529);
nor U725 (N_725,N_437,N_489);
nor U726 (N_726,N_598,N_451);
and U727 (N_727,N_405,N_457);
or U728 (N_728,N_521,N_458);
and U729 (N_729,N_552,N_551);
and U730 (N_730,N_534,N_512);
or U731 (N_731,N_552,N_533);
and U732 (N_732,N_455,N_536);
nand U733 (N_733,N_441,N_514);
or U734 (N_734,N_478,N_450);
or U735 (N_735,N_495,N_584);
nand U736 (N_736,N_482,N_449);
nor U737 (N_737,N_406,N_521);
or U738 (N_738,N_422,N_586);
nor U739 (N_739,N_427,N_492);
or U740 (N_740,N_481,N_492);
or U741 (N_741,N_519,N_409);
nand U742 (N_742,N_539,N_480);
or U743 (N_743,N_523,N_538);
or U744 (N_744,N_482,N_421);
or U745 (N_745,N_418,N_496);
and U746 (N_746,N_491,N_452);
nor U747 (N_747,N_486,N_518);
nand U748 (N_748,N_577,N_563);
nor U749 (N_749,N_440,N_582);
and U750 (N_750,N_522,N_400);
nor U751 (N_751,N_428,N_561);
nand U752 (N_752,N_548,N_437);
nand U753 (N_753,N_416,N_422);
or U754 (N_754,N_593,N_513);
or U755 (N_755,N_499,N_543);
nor U756 (N_756,N_406,N_437);
nor U757 (N_757,N_451,N_437);
nand U758 (N_758,N_497,N_515);
and U759 (N_759,N_507,N_490);
and U760 (N_760,N_488,N_480);
and U761 (N_761,N_573,N_443);
nand U762 (N_762,N_513,N_482);
nand U763 (N_763,N_555,N_456);
nor U764 (N_764,N_460,N_404);
nand U765 (N_765,N_555,N_566);
and U766 (N_766,N_551,N_437);
and U767 (N_767,N_458,N_436);
and U768 (N_768,N_470,N_559);
and U769 (N_769,N_513,N_486);
or U770 (N_770,N_530,N_425);
and U771 (N_771,N_580,N_466);
or U772 (N_772,N_589,N_551);
nor U773 (N_773,N_549,N_408);
or U774 (N_774,N_438,N_418);
nor U775 (N_775,N_421,N_501);
or U776 (N_776,N_597,N_592);
and U777 (N_777,N_457,N_452);
nand U778 (N_778,N_447,N_433);
and U779 (N_779,N_518,N_550);
and U780 (N_780,N_525,N_438);
nor U781 (N_781,N_488,N_578);
or U782 (N_782,N_540,N_462);
and U783 (N_783,N_433,N_542);
and U784 (N_784,N_511,N_456);
and U785 (N_785,N_469,N_443);
and U786 (N_786,N_562,N_424);
nand U787 (N_787,N_554,N_449);
nand U788 (N_788,N_517,N_477);
nand U789 (N_789,N_563,N_428);
nand U790 (N_790,N_592,N_506);
nand U791 (N_791,N_556,N_416);
and U792 (N_792,N_539,N_474);
nor U793 (N_793,N_582,N_478);
nor U794 (N_794,N_560,N_407);
and U795 (N_795,N_505,N_412);
nand U796 (N_796,N_465,N_514);
nand U797 (N_797,N_450,N_500);
nand U798 (N_798,N_551,N_523);
or U799 (N_799,N_576,N_490);
and U800 (N_800,N_643,N_726);
or U801 (N_801,N_687,N_667);
and U802 (N_802,N_712,N_769);
or U803 (N_803,N_627,N_664);
and U804 (N_804,N_648,N_697);
and U805 (N_805,N_662,N_760);
and U806 (N_806,N_683,N_796);
or U807 (N_807,N_617,N_694);
nor U808 (N_808,N_693,N_671);
or U809 (N_809,N_729,N_636);
nand U810 (N_810,N_625,N_799);
or U811 (N_811,N_780,N_742);
nor U812 (N_812,N_758,N_727);
and U813 (N_813,N_637,N_656);
nand U814 (N_814,N_620,N_724);
or U815 (N_815,N_644,N_604);
nor U816 (N_816,N_794,N_791);
nand U817 (N_817,N_610,N_663);
nor U818 (N_818,N_673,N_650);
and U819 (N_819,N_642,N_657);
nand U820 (N_820,N_615,N_741);
xor U821 (N_821,N_661,N_764);
nor U822 (N_822,N_612,N_776);
nand U823 (N_823,N_613,N_665);
nand U824 (N_824,N_700,N_649);
nor U825 (N_825,N_715,N_768);
or U826 (N_826,N_708,N_606);
or U827 (N_827,N_737,N_631);
or U828 (N_828,N_679,N_674);
nand U829 (N_829,N_774,N_739);
nor U830 (N_830,N_713,N_785);
nor U831 (N_831,N_781,N_778);
nor U832 (N_832,N_702,N_755);
nand U833 (N_833,N_782,N_744);
xnor U834 (N_834,N_734,N_775);
nand U835 (N_835,N_784,N_777);
nand U836 (N_836,N_770,N_728);
or U837 (N_837,N_732,N_761);
nor U838 (N_838,N_668,N_669);
or U839 (N_839,N_685,N_771);
nor U840 (N_840,N_691,N_660);
nand U841 (N_841,N_624,N_719);
nor U842 (N_842,N_688,N_640);
nand U843 (N_843,N_720,N_692);
or U844 (N_844,N_754,N_705);
and U845 (N_845,N_709,N_628);
or U846 (N_846,N_797,N_696);
nor U847 (N_847,N_611,N_751);
and U848 (N_848,N_602,N_757);
or U849 (N_849,N_600,N_772);
or U850 (N_850,N_601,N_675);
nand U851 (N_851,N_701,N_786);
or U852 (N_852,N_623,N_635);
or U853 (N_853,N_767,N_733);
nor U854 (N_854,N_753,N_655);
and U855 (N_855,N_698,N_750);
nor U856 (N_856,N_722,N_630);
or U857 (N_857,N_618,N_795);
and U858 (N_858,N_735,N_680);
or U859 (N_859,N_638,N_629);
nor U860 (N_860,N_653,N_639);
and U861 (N_861,N_621,N_658);
nand U862 (N_862,N_607,N_756);
nand U863 (N_863,N_706,N_654);
and U864 (N_864,N_690,N_609);
nand U865 (N_865,N_689,N_633);
and U866 (N_866,N_740,N_787);
nor U867 (N_867,N_789,N_676);
or U868 (N_868,N_752,N_646);
nand U869 (N_869,N_783,N_717);
and U870 (N_870,N_632,N_721);
or U871 (N_871,N_603,N_614);
or U872 (N_872,N_619,N_762);
and U873 (N_873,N_793,N_641);
and U874 (N_874,N_792,N_798);
or U875 (N_875,N_616,N_677);
or U876 (N_876,N_704,N_743);
nor U877 (N_877,N_749,N_672);
nor U878 (N_878,N_634,N_647);
nor U879 (N_879,N_736,N_703);
nor U880 (N_880,N_686,N_684);
and U881 (N_881,N_725,N_605);
nand U882 (N_882,N_763,N_788);
nor U883 (N_883,N_746,N_608);
or U884 (N_884,N_659,N_716);
nand U885 (N_885,N_695,N_745);
or U886 (N_886,N_766,N_699);
nor U887 (N_887,N_626,N_765);
nand U888 (N_888,N_707,N_730);
nand U889 (N_889,N_773,N_759);
or U890 (N_890,N_747,N_779);
and U891 (N_891,N_670,N_748);
or U892 (N_892,N_714,N_645);
nand U893 (N_893,N_678,N_652);
or U894 (N_894,N_790,N_731);
nor U895 (N_895,N_718,N_723);
nor U896 (N_896,N_622,N_711);
nand U897 (N_897,N_666,N_681);
and U898 (N_898,N_682,N_710);
nor U899 (N_899,N_738,N_651);
nand U900 (N_900,N_629,N_667);
nor U901 (N_901,N_640,N_682);
nand U902 (N_902,N_605,N_748);
or U903 (N_903,N_613,N_755);
or U904 (N_904,N_755,N_785);
or U905 (N_905,N_699,N_688);
and U906 (N_906,N_732,N_645);
nor U907 (N_907,N_624,N_722);
nand U908 (N_908,N_626,N_796);
and U909 (N_909,N_685,N_659);
nor U910 (N_910,N_677,N_735);
or U911 (N_911,N_614,N_752);
nor U912 (N_912,N_750,N_628);
and U913 (N_913,N_728,N_636);
and U914 (N_914,N_734,N_776);
nand U915 (N_915,N_728,N_747);
or U916 (N_916,N_778,N_686);
nor U917 (N_917,N_725,N_744);
xor U918 (N_918,N_681,N_720);
nand U919 (N_919,N_627,N_753);
or U920 (N_920,N_670,N_717);
and U921 (N_921,N_745,N_723);
and U922 (N_922,N_699,N_682);
or U923 (N_923,N_622,N_638);
nand U924 (N_924,N_601,N_776);
or U925 (N_925,N_683,N_671);
and U926 (N_926,N_727,N_782);
nand U927 (N_927,N_649,N_705);
and U928 (N_928,N_692,N_693);
nand U929 (N_929,N_761,N_727);
nand U930 (N_930,N_719,N_725);
and U931 (N_931,N_682,N_730);
nor U932 (N_932,N_715,N_713);
or U933 (N_933,N_709,N_700);
nor U934 (N_934,N_685,N_775);
nor U935 (N_935,N_774,N_741);
and U936 (N_936,N_771,N_769);
and U937 (N_937,N_773,N_618);
nor U938 (N_938,N_721,N_601);
nor U939 (N_939,N_703,N_716);
nor U940 (N_940,N_645,N_767);
nor U941 (N_941,N_662,N_614);
and U942 (N_942,N_707,N_632);
nor U943 (N_943,N_606,N_650);
nor U944 (N_944,N_749,N_614);
nand U945 (N_945,N_673,N_705);
nor U946 (N_946,N_750,N_738);
nor U947 (N_947,N_786,N_620);
and U948 (N_948,N_648,N_601);
nor U949 (N_949,N_710,N_622);
nor U950 (N_950,N_727,N_604);
nand U951 (N_951,N_627,N_609);
nand U952 (N_952,N_773,N_626);
nand U953 (N_953,N_689,N_667);
nor U954 (N_954,N_721,N_692);
or U955 (N_955,N_745,N_799);
or U956 (N_956,N_775,N_776);
nand U957 (N_957,N_690,N_778);
and U958 (N_958,N_679,N_659);
nor U959 (N_959,N_648,N_768);
and U960 (N_960,N_770,N_694);
nand U961 (N_961,N_737,N_728);
or U962 (N_962,N_724,N_678);
and U963 (N_963,N_715,N_630);
nand U964 (N_964,N_742,N_673);
nor U965 (N_965,N_665,N_737);
nor U966 (N_966,N_645,N_602);
nor U967 (N_967,N_674,N_780);
nor U968 (N_968,N_669,N_630);
and U969 (N_969,N_703,N_628);
or U970 (N_970,N_614,N_610);
and U971 (N_971,N_694,N_771);
nor U972 (N_972,N_693,N_657);
or U973 (N_973,N_736,N_633);
nand U974 (N_974,N_793,N_686);
nor U975 (N_975,N_615,N_757);
nand U976 (N_976,N_644,N_665);
nand U977 (N_977,N_726,N_741);
and U978 (N_978,N_645,N_723);
or U979 (N_979,N_770,N_763);
nor U980 (N_980,N_651,N_647);
nor U981 (N_981,N_610,N_603);
or U982 (N_982,N_633,N_688);
and U983 (N_983,N_687,N_644);
and U984 (N_984,N_626,N_743);
or U985 (N_985,N_616,N_799);
nand U986 (N_986,N_724,N_706);
nand U987 (N_987,N_724,N_717);
and U988 (N_988,N_670,N_624);
nor U989 (N_989,N_794,N_772);
nor U990 (N_990,N_626,N_676);
or U991 (N_991,N_784,N_609);
nor U992 (N_992,N_712,N_608);
and U993 (N_993,N_640,N_697);
nor U994 (N_994,N_686,N_714);
or U995 (N_995,N_701,N_677);
nand U996 (N_996,N_747,N_611);
or U997 (N_997,N_675,N_795);
and U998 (N_998,N_648,N_776);
or U999 (N_999,N_703,N_733);
nand U1000 (N_1000,N_957,N_876);
nand U1001 (N_1001,N_882,N_858);
nor U1002 (N_1002,N_877,N_989);
and U1003 (N_1003,N_949,N_866);
nand U1004 (N_1004,N_856,N_948);
nor U1005 (N_1005,N_923,N_965);
and U1006 (N_1006,N_873,N_811);
and U1007 (N_1007,N_920,N_977);
or U1008 (N_1008,N_905,N_883);
or U1009 (N_1009,N_919,N_975);
nor U1010 (N_1010,N_937,N_821);
xor U1011 (N_1011,N_844,N_847);
and U1012 (N_1012,N_978,N_933);
nand U1013 (N_1013,N_820,N_888);
or U1014 (N_1014,N_834,N_867);
and U1015 (N_1015,N_988,N_926);
nor U1016 (N_1016,N_852,N_803);
nor U1017 (N_1017,N_947,N_941);
and U1018 (N_1018,N_857,N_804);
and U1019 (N_1019,N_816,N_909);
and U1020 (N_1020,N_936,N_906);
and U1021 (N_1021,N_964,N_907);
nand U1022 (N_1022,N_929,N_984);
and U1023 (N_1023,N_991,N_843);
nand U1024 (N_1024,N_939,N_963);
nand U1025 (N_1025,N_953,N_955);
nor U1026 (N_1026,N_841,N_951);
nand U1027 (N_1027,N_863,N_842);
nor U1028 (N_1028,N_887,N_818);
or U1029 (N_1029,N_924,N_826);
and U1030 (N_1030,N_854,N_845);
nand U1031 (N_1031,N_896,N_925);
or U1032 (N_1032,N_945,N_817);
or U1033 (N_1033,N_899,N_908);
or U1034 (N_1034,N_934,N_830);
or U1035 (N_1035,N_892,N_979);
or U1036 (N_1036,N_998,N_930);
nor U1037 (N_1037,N_806,N_808);
nand U1038 (N_1038,N_972,N_802);
or U1039 (N_1039,N_956,N_800);
nor U1040 (N_1040,N_827,N_838);
or U1041 (N_1041,N_864,N_801);
nor U1042 (N_1042,N_889,N_990);
nor U1043 (N_1043,N_961,N_822);
nand U1044 (N_1044,N_828,N_954);
nor U1045 (N_1045,N_996,N_879);
nor U1046 (N_1046,N_943,N_938);
or U1047 (N_1047,N_966,N_898);
and U1048 (N_1048,N_962,N_987);
nand U1049 (N_1049,N_950,N_895);
or U1050 (N_1050,N_922,N_983);
and U1051 (N_1051,N_809,N_851);
and U1052 (N_1052,N_805,N_917);
nand U1053 (N_1053,N_981,N_902);
nor U1054 (N_1054,N_940,N_969);
nor U1055 (N_1055,N_831,N_944);
or U1056 (N_1056,N_927,N_960);
and U1057 (N_1057,N_872,N_824);
or U1058 (N_1058,N_900,N_995);
or U1059 (N_1059,N_807,N_814);
nand U1060 (N_1060,N_985,N_835);
nand U1061 (N_1061,N_946,N_859);
nand U1062 (N_1062,N_994,N_846);
and U1063 (N_1063,N_819,N_986);
nor U1064 (N_1064,N_881,N_968);
nand U1065 (N_1065,N_942,N_973);
or U1066 (N_1066,N_880,N_980);
nand U1067 (N_1067,N_853,N_823);
and U1068 (N_1068,N_894,N_832);
or U1069 (N_1069,N_885,N_868);
nand U1070 (N_1070,N_901,N_976);
and U1071 (N_1071,N_903,N_836);
nor U1072 (N_1072,N_916,N_810);
nand U1073 (N_1073,N_850,N_959);
nor U1074 (N_1074,N_862,N_997);
or U1075 (N_1075,N_870,N_915);
and U1076 (N_1076,N_855,N_840);
nand U1077 (N_1077,N_865,N_974);
or U1078 (N_1078,N_837,N_829);
xor U1079 (N_1079,N_993,N_860);
and U1080 (N_1080,N_932,N_890);
or U1081 (N_1081,N_825,N_992);
and U1082 (N_1082,N_913,N_910);
or U1083 (N_1083,N_833,N_869);
or U1084 (N_1084,N_971,N_967);
and U1085 (N_1085,N_970,N_874);
xor U1086 (N_1086,N_812,N_813);
or U1087 (N_1087,N_886,N_931);
nor U1088 (N_1088,N_958,N_839);
nor U1089 (N_1089,N_935,N_952);
nand U1090 (N_1090,N_861,N_921);
nor U1091 (N_1091,N_912,N_911);
and U1092 (N_1092,N_914,N_893);
and U1093 (N_1093,N_884,N_871);
nand U1094 (N_1094,N_918,N_928);
or U1095 (N_1095,N_875,N_878);
nand U1096 (N_1096,N_999,N_848);
and U1097 (N_1097,N_904,N_815);
nand U1098 (N_1098,N_897,N_891);
or U1099 (N_1099,N_982,N_849);
nor U1100 (N_1100,N_978,N_822);
or U1101 (N_1101,N_902,N_810);
nor U1102 (N_1102,N_995,N_829);
or U1103 (N_1103,N_972,N_919);
or U1104 (N_1104,N_891,N_927);
or U1105 (N_1105,N_808,N_982);
nor U1106 (N_1106,N_962,N_986);
and U1107 (N_1107,N_966,N_942);
or U1108 (N_1108,N_864,N_937);
nor U1109 (N_1109,N_930,N_873);
nand U1110 (N_1110,N_990,N_972);
and U1111 (N_1111,N_945,N_806);
nand U1112 (N_1112,N_943,N_903);
nand U1113 (N_1113,N_969,N_945);
nand U1114 (N_1114,N_941,N_967);
nand U1115 (N_1115,N_809,N_998);
and U1116 (N_1116,N_961,N_972);
and U1117 (N_1117,N_805,N_869);
nor U1118 (N_1118,N_889,N_978);
nand U1119 (N_1119,N_947,N_882);
nand U1120 (N_1120,N_825,N_868);
nor U1121 (N_1121,N_915,N_837);
nand U1122 (N_1122,N_924,N_862);
nor U1123 (N_1123,N_967,N_954);
nor U1124 (N_1124,N_984,N_905);
or U1125 (N_1125,N_844,N_897);
and U1126 (N_1126,N_957,N_911);
or U1127 (N_1127,N_962,N_951);
and U1128 (N_1128,N_882,N_832);
nor U1129 (N_1129,N_894,N_991);
nand U1130 (N_1130,N_916,N_899);
nor U1131 (N_1131,N_903,N_941);
nor U1132 (N_1132,N_853,N_837);
nor U1133 (N_1133,N_857,N_973);
nand U1134 (N_1134,N_853,N_886);
nand U1135 (N_1135,N_977,N_982);
nand U1136 (N_1136,N_925,N_888);
or U1137 (N_1137,N_901,N_820);
or U1138 (N_1138,N_812,N_987);
nor U1139 (N_1139,N_892,N_824);
or U1140 (N_1140,N_985,N_943);
nand U1141 (N_1141,N_970,N_899);
nor U1142 (N_1142,N_860,N_887);
or U1143 (N_1143,N_975,N_992);
and U1144 (N_1144,N_898,N_954);
nand U1145 (N_1145,N_883,N_898);
nor U1146 (N_1146,N_888,N_916);
nor U1147 (N_1147,N_956,N_991);
nor U1148 (N_1148,N_839,N_837);
or U1149 (N_1149,N_832,N_862);
nand U1150 (N_1150,N_969,N_829);
nand U1151 (N_1151,N_975,N_815);
nand U1152 (N_1152,N_993,N_805);
nand U1153 (N_1153,N_804,N_915);
and U1154 (N_1154,N_840,N_815);
nor U1155 (N_1155,N_965,N_899);
or U1156 (N_1156,N_861,N_996);
nand U1157 (N_1157,N_998,N_979);
nor U1158 (N_1158,N_997,N_965);
and U1159 (N_1159,N_871,N_903);
or U1160 (N_1160,N_852,N_954);
and U1161 (N_1161,N_921,N_897);
nor U1162 (N_1162,N_871,N_977);
nor U1163 (N_1163,N_907,N_974);
and U1164 (N_1164,N_898,N_961);
nand U1165 (N_1165,N_892,N_883);
nand U1166 (N_1166,N_853,N_903);
and U1167 (N_1167,N_832,N_833);
nand U1168 (N_1168,N_909,N_898);
nor U1169 (N_1169,N_973,N_933);
or U1170 (N_1170,N_875,N_822);
nand U1171 (N_1171,N_924,N_819);
and U1172 (N_1172,N_927,N_931);
or U1173 (N_1173,N_811,N_976);
nand U1174 (N_1174,N_847,N_951);
or U1175 (N_1175,N_946,N_831);
and U1176 (N_1176,N_960,N_908);
nor U1177 (N_1177,N_996,N_824);
or U1178 (N_1178,N_928,N_817);
nor U1179 (N_1179,N_966,N_896);
or U1180 (N_1180,N_854,N_844);
nor U1181 (N_1181,N_821,N_957);
nand U1182 (N_1182,N_983,N_871);
nand U1183 (N_1183,N_948,N_880);
and U1184 (N_1184,N_974,N_870);
and U1185 (N_1185,N_829,N_883);
nand U1186 (N_1186,N_868,N_940);
nand U1187 (N_1187,N_800,N_824);
nor U1188 (N_1188,N_843,N_942);
nor U1189 (N_1189,N_811,N_858);
nand U1190 (N_1190,N_984,N_820);
nor U1191 (N_1191,N_814,N_810);
or U1192 (N_1192,N_834,N_908);
nor U1193 (N_1193,N_806,N_979);
and U1194 (N_1194,N_986,N_960);
nand U1195 (N_1195,N_896,N_843);
or U1196 (N_1196,N_973,N_882);
or U1197 (N_1197,N_801,N_853);
nor U1198 (N_1198,N_888,N_944);
or U1199 (N_1199,N_951,N_916);
nand U1200 (N_1200,N_1105,N_1013);
or U1201 (N_1201,N_1190,N_1044);
and U1202 (N_1202,N_1187,N_1090);
nor U1203 (N_1203,N_1134,N_1152);
or U1204 (N_1204,N_1102,N_1178);
and U1205 (N_1205,N_1151,N_1164);
and U1206 (N_1206,N_1149,N_1036);
and U1207 (N_1207,N_1162,N_1147);
or U1208 (N_1208,N_1086,N_1096);
or U1209 (N_1209,N_1006,N_1154);
nand U1210 (N_1210,N_1041,N_1046);
nand U1211 (N_1211,N_1167,N_1042);
and U1212 (N_1212,N_1195,N_1139);
nor U1213 (N_1213,N_1043,N_1197);
nand U1214 (N_1214,N_1170,N_1122);
or U1215 (N_1215,N_1072,N_1039);
nor U1216 (N_1216,N_1020,N_1131);
and U1217 (N_1217,N_1088,N_1063);
nor U1218 (N_1218,N_1113,N_1062);
nand U1219 (N_1219,N_1015,N_1185);
and U1220 (N_1220,N_1002,N_1057);
and U1221 (N_1221,N_1196,N_1128);
and U1222 (N_1222,N_1012,N_1172);
nor U1223 (N_1223,N_1125,N_1047);
nand U1224 (N_1224,N_1118,N_1037);
and U1225 (N_1225,N_1048,N_1153);
and U1226 (N_1226,N_1022,N_1000);
nand U1227 (N_1227,N_1021,N_1106);
nor U1228 (N_1228,N_1007,N_1191);
or U1229 (N_1229,N_1138,N_1065);
and U1230 (N_1230,N_1028,N_1142);
nor U1231 (N_1231,N_1155,N_1034);
and U1232 (N_1232,N_1010,N_1071);
and U1233 (N_1233,N_1101,N_1097);
nor U1234 (N_1234,N_1098,N_1176);
xnor U1235 (N_1235,N_1052,N_1011);
nand U1236 (N_1236,N_1112,N_1068);
nor U1237 (N_1237,N_1163,N_1144);
nor U1238 (N_1238,N_1005,N_1076);
and U1239 (N_1239,N_1182,N_1115);
nor U1240 (N_1240,N_1130,N_1018);
nand U1241 (N_1241,N_1129,N_1024);
nor U1242 (N_1242,N_1161,N_1014);
nand U1243 (N_1243,N_1188,N_1023);
and U1244 (N_1244,N_1059,N_1035);
or U1245 (N_1245,N_1078,N_1027);
nor U1246 (N_1246,N_1111,N_1119);
or U1247 (N_1247,N_1186,N_1140);
nand U1248 (N_1248,N_1133,N_1091);
and U1249 (N_1249,N_1089,N_1177);
or U1250 (N_1250,N_1087,N_1019);
nand U1251 (N_1251,N_1114,N_1031);
or U1252 (N_1252,N_1104,N_1120);
or U1253 (N_1253,N_1193,N_1171);
and U1254 (N_1254,N_1081,N_1169);
or U1255 (N_1255,N_1085,N_1137);
or U1256 (N_1256,N_1053,N_1054);
and U1257 (N_1257,N_1173,N_1074);
nor U1258 (N_1258,N_1030,N_1056);
nand U1259 (N_1259,N_1095,N_1159);
nor U1260 (N_1260,N_1073,N_1077);
nor U1261 (N_1261,N_1124,N_1156);
nor U1262 (N_1262,N_1029,N_1189);
or U1263 (N_1263,N_1108,N_1121);
and U1264 (N_1264,N_1079,N_1066);
and U1265 (N_1265,N_1168,N_1050);
nand U1266 (N_1266,N_1080,N_1003);
and U1267 (N_1267,N_1058,N_1145);
nor U1268 (N_1268,N_1051,N_1150);
nand U1269 (N_1269,N_1181,N_1148);
nor U1270 (N_1270,N_1067,N_1026);
nand U1271 (N_1271,N_1123,N_1157);
and U1272 (N_1272,N_1061,N_1146);
nand U1273 (N_1273,N_1117,N_1135);
and U1274 (N_1274,N_1001,N_1116);
or U1275 (N_1275,N_1017,N_1070);
nor U1276 (N_1276,N_1174,N_1192);
nand U1277 (N_1277,N_1016,N_1160);
nand U1278 (N_1278,N_1158,N_1045);
and U1279 (N_1279,N_1194,N_1055);
nor U1280 (N_1280,N_1075,N_1100);
and U1281 (N_1281,N_1141,N_1107);
or U1282 (N_1282,N_1184,N_1110);
nor U1283 (N_1283,N_1038,N_1166);
and U1284 (N_1284,N_1143,N_1099);
and U1285 (N_1285,N_1009,N_1127);
nand U1286 (N_1286,N_1132,N_1084);
and U1287 (N_1287,N_1092,N_1083);
and U1288 (N_1288,N_1109,N_1165);
nand U1289 (N_1289,N_1033,N_1093);
xnor U1290 (N_1290,N_1199,N_1069);
nand U1291 (N_1291,N_1008,N_1126);
nand U1292 (N_1292,N_1032,N_1179);
or U1293 (N_1293,N_1049,N_1025);
and U1294 (N_1294,N_1175,N_1082);
and U1295 (N_1295,N_1094,N_1183);
nor U1296 (N_1296,N_1060,N_1064);
nor U1297 (N_1297,N_1136,N_1103);
nor U1298 (N_1298,N_1004,N_1198);
nor U1299 (N_1299,N_1180,N_1040);
or U1300 (N_1300,N_1074,N_1158);
and U1301 (N_1301,N_1044,N_1053);
nor U1302 (N_1302,N_1018,N_1034);
nor U1303 (N_1303,N_1034,N_1156);
and U1304 (N_1304,N_1168,N_1104);
nor U1305 (N_1305,N_1159,N_1197);
or U1306 (N_1306,N_1063,N_1142);
and U1307 (N_1307,N_1196,N_1112);
and U1308 (N_1308,N_1009,N_1078);
nor U1309 (N_1309,N_1015,N_1057);
or U1310 (N_1310,N_1005,N_1188);
nand U1311 (N_1311,N_1126,N_1099);
and U1312 (N_1312,N_1183,N_1166);
or U1313 (N_1313,N_1057,N_1083);
nor U1314 (N_1314,N_1107,N_1083);
or U1315 (N_1315,N_1089,N_1108);
nor U1316 (N_1316,N_1030,N_1141);
nor U1317 (N_1317,N_1175,N_1049);
and U1318 (N_1318,N_1056,N_1109);
or U1319 (N_1319,N_1183,N_1040);
nand U1320 (N_1320,N_1148,N_1102);
nor U1321 (N_1321,N_1069,N_1173);
or U1322 (N_1322,N_1018,N_1023);
nor U1323 (N_1323,N_1135,N_1051);
or U1324 (N_1324,N_1195,N_1046);
nor U1325 (N_1325,N_1081,N_1182);
nand U1326 (N_1326,N_1178,N_1054);
or U1327 (N_1327,N_1083,N_1165);
nand U1328 (N_1328,N_1052,N_1156);
nor U1329 (N_1329,N_1157,N_1027);
or U1330 (N_1330,N_1197,N_1077);
nand U1331 (N_1331,N_1005,N_1102);
nand U1332 (N_1332,N_1019,N_1179);
and U1333 (N_1333,N_1042,N_1014);
nor U1334 (N_1334,N_1046,N_1044);
nor U1335 (N_1335,N_1073,N_1146);
or U1336 (N_1336,N_1116,N_1106);
nor U1337 (N_1337,N_1047,N_1101);
or U1338 (N_1338,N_1197,N_1093);
and U1339 (N_1339,N_1082,N_1152);
and U1340 (N_1340,N_1026,N_1096);
nand U1341 (N_1341,N_1080,N_1024);
or U1342 (N_1342,N_1000,N_1174);
nand U1343 (N_1343,N_1171,N_1126);
and U1344 (N_1344,N_1163,N_1002);
nor U1345 (N_1345,N_1195,N_1147);
and U1346 (N_1346,N_1144,N_1056);
nor U1347 (N_1347,N_1129,N_1128);
or U1348 (N_1348,N_1180,N_1079);
nand U1349 (N_1349,N_1123,N_1082);
nand U1350 (N_1350,N_1056,N_1075);
and U1351 (N_1351,N_1022,N_1109);
nor U1352 (N_1352,N_1022,N_1004);
or U1353 (N_1353,N_1026,N_1033);
and U1354 (N_1354,N_1114,N_1147);
or U1355 (N_1355,N_1027,N_1167);
or U1356 (N_1356,N_1096,N_1033);
and U1357 (N_1357,N_1032,N_1065);
nand U1358 (N_1358,N_1005,N_1149);
or U1359 (N_1359,N_1167,N_1029);
or U1360 (N_1360,N_1176,N_1188);
nor U1361 (N_1361,N_1065,N_1050);
or U1362 (N_1362,N_1044,N_1032);
nor U1363 (N_1363,N_1183,N_1020);
nand U1364 (N_1364,N_1022,N_1162);
and U1365 (N_1365,N_1162,N_1199);
or U1366 (N_1366,N_1085,N_1189);
or U1367 (N_1367,N_1138,N_1142);
and U1368 (N_1368,N_1017,N_1077);
nor U1369 (N_1369,N_1029,N_1009);
or U1370 (N_1370,N_1164,N_1097);
nor U1371 (N_1371,N_1142,N_1067);
and U1372 (N_1372,N_1043,N_1045);
nand U1373 (N_1373,N_1184,N_1020);
nor U1374 (N_1374,N_1095,N_1162);
or U1375 (N_1375,N_1071,N_1037);
and U1376 (N_1376,N_1025,N_1033);
nand U1377 (N_1377,N_1159,N_1173);
or U1378 (N_1378,N_1117,N_1072);
or U1379 (N_1379,N_1082,N_1159);
nor U1380 (N_1380,N_1180,N_1085);
and U1381 (N_1381,N_1088,N_1193);
and U1382 (N_1382,N_1067,N_1183);
nor U1383 (N_1383,N_1079,N_1076);
nor U1384 (N_1384,N_1076,N_1102);
and U1385 (N_1385,N_1157,N_1192);
and U1386 (N_1386,N_1079,N_1197);
nand U1387 (N_1387,N_1129,N_1025);
or U1388 (N_1388,N_1087,N_1163);
and U1389 (N_1389,N_1021,N_1017);
nand U1390 (N_1390,N_1193,N_1001);
nand U1391 (N_1391,N_1111,N_1034);
and U1392 (N_1392,N_1189,N_1098);
and U1393 (N_1393,N_1152,N_1018);
or U1394 (N_1394,N_1196,N_1182);
or U1395 (N_1395,N_1113,N_1151);
nand U1396 (N_1396,N_1179,N_1191);
or U1397 (N_1397,N_1142,N_1045);
or U1398 (N_1398,N_1091,N_1020);
and U1399 (N_1399,N_1094,N_1186);
and U1400 (N_1400,N_1204,N_1254);
nand U1401 (N_1401,N_1344,N_1206);
nor U1402 (N_1402,N_1336,N_1340);
nand U1403 (N_1403,N_1350,N_1239);
and U1404 (N_1404,N_1289,N_1379);
nand U1405 (N_1405,N_1361,N_1390);
nor U1406 (N_1406,N_1359,N_1322);
nand U1407 (N_1407,N_1243,N_1286);
and U1408 (N_1408,N_1365,N_1298);
and U1409 (N_1409,N_1266,N_1332);
and U1410 (N_1410,N_1217,N_1372);
or U1411 (N_1411,N_1326,N_1327);
and U1412 (N_1412,N_1224,N_1240);
and U1413 (N_1413,N_1395,N_1329);
and U1414 (N_1414,N_1354,N_1269);
and U1415 (N_1415,N_1393,N_1335);
nor U1416 (N_1416,N_1323,N_1290);
or U1417 (N_1417,N_1328,N_1397);
or U1418 (N_1418,N_1392,N_1312);
and U1419 (N_1419,N_1317,N_1315);
and U1420 (N_1420,N_1234,N_1325);
and U1421 (N_1421,N_1352,N_1351);
nor U1422 (N_1422,N_1292,N_1252);
or U1423 (N_1423,N_1238,N_1235);
or U1424 (N_1424,N_1376,N_1229);
or U1425 (N_1425,N_1313,N_1345);
or U1426 (N_1426,N_1341,N_1346);
nor U1427 (N_1427,N_1314,N_1246);
or U1428 (N_1428,N_1202,N_1384);
and U1429 (N_1429,N_1277,N_1241);
nand U1430 (N_1430,N_1226,N_1219);
nor U1431 (N_1431,N_1296,N_1330);
and U1432 (N_1432,N_1378,N_1220);
and U1433 (N_1433,N_1318,N_1270);
and U1434 (N_1434,N_1309,N_1380);
and U1435 (N_1435,N_1389,N_1360);
or U1436 (N_1436,N_1253,N_1256);
nor U1437 (N_1437,N_1310,N_1207);
nand U1438 (N_1438,N_1374,N_1237);
nand U1439 (N_1439,N_1259,N_1299);
and U1440 (N_1440,N_1334,N_1213);
and U1441 (N_1441,N_1348,N_1362);
and U1442 (N_1442,N_1337,N_1285);
nor U1443 (N_1443,N_1368,N_1386);
nand U1444 (N_1444,N_1225,N_1230);
or U1445 (N_1445,N_1331,N_1321);
or U1446 (N_1446,N_1281,N_1210);
and U1447 (N_1447,N_1342,N_1394);
nand U1448 (N_1448,N_1282,N_1244);
nor U1449 (N_1449,N_1358,N_1353);
nor U1450 (N_1450,N_1349,N_1320);
nand U1451 (N_1451,N_1221,N_1249);
and U1452 (N_1452,N_1355,N_1271);
and U1453 (N_1453,N_1261,N_1245);
nor U1454 (N_1454,N_1250,N_1232);
nand U1455 (N_1455,N_1264,N_1302);
or U1456 (N_1456,N_1223,N_1399);
nand U1457 (N_1457,N_1274,N_1248);
and U1458 (N_1458,N_1216,N_1279);
nand U1459 (N_1459,N_1201,N_1303);
nor U1460 (N_1460,N_1398,N_1366);
and U1461 (N_1461,N_1247,N_1257);
or U1462 (N_1462,N_1278,N_1295);
or U1463 (N_1463,N_1396,N_1227);
and U1464 (N_1464,N_1381,N_1242);
nor U1465 (N_1465,N_1275,N_1306);
or U1466 (N_1466,N_1311,N_1371);
and U1467 (N_1467,N_1258,N_1373);
nor U1468 (N_1468,N_1391,N_1215);
or U1469 (N_1469,N_1288,N_1367);
or U1470 (N_1470,N_1370,N_1388);
nand U1471 (N_1471,N_1338,N_1236);
or U1472 (N_1472,N_1297,N_1211);
or U1473 (N_1473,N_1375,N_1364);
nand U1474 (N_1474,N_1324,N_1233);
or U1475 (N_1475,N_1284,N_1304);
nand U1476 (N_1476,N_1356,N_1208);
nor U1477 (N_1477,N_1343,N_1333);
and U1478 (N_1478,N_1383,N_1251);
and U1479 (N_1479,N_1377,N_1205);
nand U1480 (N_1480,N_1260,N_1308);
or U1481 (N_1481,N_1267,N_1293);
and U1482 (N_1482,N_1357,N_1363);
and U1483 (N_1483,N_1200,N_1222);
nor U1484 (N_1484,N_1307,N_1231);
nor U1485 (N_1485,N_1294,N_1369);
or U1486 (N_1486,N_1291,N_1268);
nor U1487 (N_1487,N_1339,N_1214);
nand U1488 (N_1488,N_1203,N_1255);
and U1489 (N_1489,N_1276,N_1319);
and U1490 (N_1490,N_1218,N_1228);
or U1491 (N_1491,N_1212,N_1301);
or U1492 (N_1492,N_1385,N_1283);
and U1493 (N_1493,N_1263,N_1316);
or U1494 (N_1494,N_1347,N_1305);
nand U1495 (N_1495,N_1300,N_1280);
nor U1496 (N_1496,N_1273,N_1272);
nand U1497 (N_1497,N_1265,N_1387);
or U1498 (N_1498,N_1209,N_1382);
and U1499 (N_1499,N_1262,N_1287);
or U1500 (N_1500,N_1313,N_1280);
and U1501 (N_1501,N_1374,N_1299);
nand U1502 (N_1502,N_1218,N_1315);
nor U1503 (N_1503,N_1296,N_1300);
and U1504 (N_1504,N_1398,N_1275);
and U1505 (N_1505,N_1379,N_1345);
or U1506 (N_1506,N_1369,N_1334);
and U1507 (N_1507,N_1273,N_1209);
nor U1508 (N_1508,N_1314,N_1276);
nand U1509 (N_1509,N_1338,N_1377);
and U1510 (N_1510,N_1297,N_1248);
or U1511 (N_1511,N_1301,N_1365);
nand U1512 (N_1512,N_1241,N_1330);
and U1513 (N_1513,N_1333,N_1379);
nand U1514 (N_1514,N_1369,N_1212);
and U1515 (N_1515,N_1215,N_1220);
and U1516 (N_1516,N_1309,N_1335);
or U1517 (N_1517,N_1213,N_1352);
nor U1518 (N_1518,N_1358,N_1284);
or U1519 (N_1519,N_1296,N_1271);
or U1520 (N_1520,N_1235,N_1250);
and U1521 (N_1521,N_1322,N_1253);
nor U1522 (N_1522,N_1218,N_1375);
xor U1523 (N_1523,N_1357,N_1238);
or U1524 (N_1524,N_1281,N_1277);
and U1525 (N_1525,N_1287,N_1398);
nor U1526 (N_1526,N_1205,N_1291);
xnor U1527 (N_1527,N_1399,N_1326);
nand U1528 (N_1528,N_1210,N_1277);
and U1529 (N_1529,N_1298,N_1357);
nand U1530 (N_1530,N_1202,N_1224);
nor U1531 (N_1531,N_1298,N_1374);
and U1532 (N_1532,N_1334,N_1270);
nor U1533 (N_1533,N_1337,N_1340);
nand U1534 (N_1534,N_1360,N_1257);
nand U1535 (N_1535,N_1303,N_1246);
nor U1536 (N_1536,N_1212,N_1320);
and U1537 (N_1537,N_1329,N_1244);
nand U1538 (N_1538,N_1211,N_1336);
nor U1539 (N_1539,N_1318,N_1367);
and U1540 (N_1540,N_1233,N_1300);
xnor U1541 (N_1541,N_1267,N_1379);
nor U1542 (N_1542,N_1302,N_1348);
nor U1543 (N_1543,N_1307,N_1378);
and U1544 (N_1544,N_1320,N_1396);
and U1545 (N_1545,N_1248,N_1343);
nand U1546 (N_1546,N_1328,N_1376);
nor U1547 (N_1547,N_1216,N_1390);
nand U1548 (N_1548,N_1279,N_1352);
nor U1549 (N_1549,N_1328,N_1343);
and U1550 (N_1550,N_1388,N_1363);
nand U1551 (N_1551,N_1233,N_1251);
nand U1552 (N_1552,N_1214,N_1345);
nor U1553 (N_1553,N_1370,N_1393);
or U1554 (N_1554,N_1266,N_1294);
nand U1555 (N_1555,N_1374,N_1309);
and U1556 (N_1556,N_1341,N_1351);
or U1557 (N_1557,N_1251,N_1331);
and U1558 (N_1558,N_1293,N_1374);
or U1559 (N_1559,N_1398,N_1311);
nand U1560 (N_1560,N_1353,N_1207);
nand U1561 (N_1561,N_1259,N_1335);
or U1562 (N_1562,N_1210,N_1249);
or U1563 (N_1563,N_1354,N_1293);
or U1564 (N_1564,N_1327,N_1387);
nor U1565 (N_1565,N_1357,N_1342);
or U1566 (N_1566,N_1208,N_1390);
nor U1567 (N_1567,N_1217,N_1206);
nand U1568 (N_1568,N_1256,N_1358);
and U1569 (N_1569,N_1353,N_1209);
nor U1570 (N_1570,N_1225,N_1263);
and U1571 (N_1571,N_1301,N_1382);
nor U1572 (N_1572,N_1309,N_1320);
and U1573 (N_1573,N_1202,N_1227);
nor U1574 (N_1574,N_1371,N_1225);
or U1575 (N_1575,N_1202,N_1247);
nor U1576 (N_1576,N_1247,N_1377);
or U1577 (N_1577,N_1329,N_1304);
nor U1578 (N_1578,N_1288,N_1203);
or U1579 (N_1579,N_1202,N_1392);
nor U1580 (N_1580,N_1232,N_1251);
nand U1581 (N_1581,N_1309,N_1336);
nor U1582 (N_1582,N_1317,N_1325);
or U1583 (N_1583,N_1325,N_1267);
nand U1584 (N_1584,N_1297,N_1349);
nor U1585 (N_1585,N_1372,N_1202);
nor U1586 (N_1586,N_1244,N_1308);
nor U1587 (N_1587,N_1353,N_1377);
and U1588 (N_1588,N_1261,N_1212);
nor U1589 (N_1589,N_1258,N_1272);
nor U1590 (N_1590,N_1259,N_1275);
nand U1591 (N_1591,N_1336,N_1293);
or U1592 (N_1592,N_1306,N_1350);
or U1593 (N_1593,N_1387,N_1299);
and U1594 (N_1594,N_1207,N_1360);
or U1595 (N_1595,N_1254,N_1235);
nor U1596 (N_1596,N_1239,N_1351);
and U1597 (N_1597,N_1248,N_1216);
nand U1598 (N_1598,N_1219,N_1224);
nand U1599 (N_1599,N_1282,N_1365);
and U1600 (N_1600,N_1569,N_1424);
and U1601 (N_1601,N_1520,N_1438);
and U1602 (N_1602,N_1579,N_1589);
or U1603 (N_1603,N_1418,N_1431);
nor U1604 (N_1604,N_1477,N_1504);
or U1605 (N_1605,N_1456,N_1455);
nor U1606 (N_1606,N_1591,N_1468);
and U1607 (N_1607,N_1474,N_1543);
and U1608 (N_1608,N_1506,N_1580);
or U1609 (N_1609,N_1551,N_1471);
nor U1610 (N_1610,N_1414,N_1412);
nor U1611 (N_1611,N_1446,N_1406);
nor U1612 (N_1612,N_1531,N_1415);
or U1613 (N_1613,N_1411,N_1558);
nor U1614 (N_1614,N_1566,N_1593);
or U1615 (N_1615,N_1545,N_1473);
nand U1616 (N_1616,N_1501,N_1507);
and U1617 (N_1617,N_1428,N_1554);
and U1618 (N_1618,N_1434,N_1461);
nor U1619 (N_1619,N_1595,N_1518);
nor U1620 (N_1620,N_1459,N_1436);
nor U1621 (N_1621,N_1449,N_1466);
or U1622 (N_1622,N_1403,N_1492);
nor U1623 (N_1623,N_1464,N_1423);
or U1624 (N_1624,N_1481,N_1425);
nand U1625 (N_1625,N_1409,N_1485);
and U1626 (N_1626,N_1450,N_1581);
nor U1627 (N_1627,N_1557,N_1586);
and U1628 (N_1628,N_1478,N_1467);
or U1629 (N_1629,N_1494,N_1517);
nor U1630 (N_1630,N_1571,N_1493);
nor U1631 (N_1631,N_1496,N_1463);
nand U1632 (N_1632,N_1408,N_1479);
nor U1633 (N_1633,N_1439,N_1495);
nand U1634 (N_1634,N_1499,N_1500);
nor U1635 (N_1635,N_1437,N_1564);
and U1636 (N_1636,N_1556,N_1539);
nor U1637 (N_1637,N_1592,N_1510);
or U1638 (N_1638,N_1599,N_1516);
nor U1639 (N_1639,N_1427,N_1401);
or U1640 (N_1640,N_1410,N_1458);
nand U1641 (N_1641,N_1513,N_1553);
or U1642 (N_1642,N_1598,N_1542);
nand U1643 (N_1643,N_1572,N_1433);
and U1644 (N_1644,N_1451,N_1570);
nor U1645 (N_1645,N_1472,N_1470);
nor U1646 (N_1646,N_1452,N_1582);
nor U1647 (N_1647,N_1521,N_1441);
or U1648 (N_1648,N_1555,N_1594);
nand U1649 (N_1649,N_1597,N_1430);
nand U1650 (N_1650,N_1535,N_1541);
and U1651 (N_1651,N_1532,N_1469);
nand U1652 (N_1652,N_1562,N_1405);
and U1653 (N_1653,N_1560,N_1453);
or U1654 (N_1654,N_1443,N_1448);
and U1655 (N_1655,N_1419,N_1476);
or U1656 (N_1656,N_1578,N_1497);
or U1657 (N_1657,N_1422,N_1530);
nor U1658 (N_1658,N_1489,N_1511);
nand U1659 (N_1659,N_1421,N_1505);
nor U1660 (N_1660,N_1587,N_1462);
nor U1661 (N_1661,N_1527,N_1454);
nor U1662 (N_1662,N_1465,N_1546);
and U1663 (N_1663,N_1568,N_1460);
or U1664 (N_1664,N_1549,N_1512);
nand U1665 (N_1665,N_1577,N_1429);
xnor U1666 (N_1666,N_1565,N_1514);
nand U1667 (N_1667,N_1561,N_1435);
nand U1668 (N_1668,N_1420,N_1559);
or U1669 (N_1669,N_1503,N_1544);
or U1670 (N_1670,N_1400,N_1575);
nor U1671 (N_1671,N_1484,N_1402);
and U1672 (N_1672,N_1480,N_1585);
nor U1673 (N_1673,N_1444,N_1588);
or U1674 (N_1674,N_1413,N_1590);
nand U1675 (N_1675,N_1567,N_1573);
nand U1676 (N_1676,N_1529,N_1536);
and U1677 (N_1677,N_1525,N_1416);
or U1678 (N_1678,N_1482,N_1584);
and U1679 (N_1679,N_1442,N_1486);
nand U1680 (N_1680,N_1515,N_1488);
nor U1681 (N_1681,N_1417,N_1475);
nor U1682 (N_1682,N_1440,N_1596);
nor U1683 (N_1683,N_1583,N_1498);
nand U1684 (N_1684,N_1432,N_1540);
nand U1685 (N_1685,N_1508,N_1533);
nor U1686 (N_1686,N_1548,N_1547);
nand U1687 (N_1687,N_1483,N_1538);
and U1688 (N_1688,N_1523,N_1487);
or U1689 (N_1689,N_1537,N_1445);
and U1690 (N_1690,N_1447,N_1534);
nand U1691 (N_1691,N_1509,N_1490);
nor U1692 (N_1692,N_1491,N_1576);
and U1693 (N_1693,N_1528,N_1502);
and U1694 (N_1694,N_1519,N_1563);
nand U1695 (N_1695,N_1526,N_1457);
nor U1696 (N_1696,N_1426,N_1522);
or U1697 (N_1697,N_1407,N_1550);
or U1698 (N_1698,N_1404,N_1524);
nor U1699 (N_1699,N_1552,N_1574);
nor U1700 (N_1700,N_1427,N_1406);
nand U1701 (N_1701,N_1415,N_1518);
nand U1702 (N_1702,N_1557,N_1404);
and U1703 (N_1703,N_1492,N_1593);
or U1704 (N_1704,N_1473,N_1400);
or U1705 (N_1705,N_1477,N_1533);
nor U1706 (N_1706,N_1574,N_1550);
or U1707 (N_1707,N_1529,N_1555);
and U1708 (N_1708,N_1543,N_1560);
nand U1709 (N_1709,N_1578,N_1475);
nand U1710 (N_1710,N_1573,N_1589);
nor U1711 (N_1711,N_1423,N_1426);
and U1712 (N_1712,N_1589,N_1571);
or U1713 (N_1713,N_1528,N_1571);
and U1714 (N_1714,N_1561,N_1441);
nand U1715 (N_1715,N_1575,N_1553);
nand U1716 (N_1716,N_1483,N_1481);
nor U1717 (N_1717,N_1555,N_1547);
nand U1718 (N_1718,N_1562,N_1556);
nand U1719 (N_1719,N_1567,N_1542);
and U1720 (N_1720,N_1496,N_1449);
nor U1721 (N_1721,N_1551,N_1496);
and U1722 (N_1722,N_1515,N_1442);
nor U1723 (N_1723,N_1558,N_1575);
and U1724 (N_1724,N_1429,N_1519);
or U1725 (N_1725,N_1510,N_1428);
or U1726 (N_1726,N_1440,N_1457);
nand U1727 (N_1727,N_1583,N_1549);
and U1728 (N_1728,N_1432,N_1533);
nand U1729 (N_1729,N_1447,N_1576);
and U1730 (N_1730,N_1471,N_1448);
and U1731 (N_1731,N_1539,N_1596);
and U1732 (N_1732,N_1448,N_1422);
nand U1733 (N_1733,N_1550,N_1561);
and U1734 (N_1734,N_1482,N_1596);
and U1735 (N_1735,N_1578,N_1495);
and U1736 (N_1736,N_1568,N_1534);
and U1737 (N_1737,N_1436,N_1452);
and U1738 (N_1738,N_1500,N_1429);
nand U1739 (N_1739,N_1442,N_1446);
nor U1740 (N_1740,N_1473,N_1491);
or U1741 (N_1741,N_1485,N_1554);
nor U1742 (N_1742,N_1530,N_1511);
and U1743 (N_1743,N_1573,N_1522);
nor U1744 (N_1744,N_1567,N_1424);
nor U1745 (N_1745,N_1462,N_1504);
nand U1746 (N_1746,N_1548,N_1408);
or U1747 (N_1747,N_1427,N_1528);
or U1748 (N_1748,N_1540,N_1459);
or U1749 (N_1749,N_1584,N_1537);
and U1750 (N_1750,N_1500,N_1572);
or U1751 (N_1751,N_1482,N_1422);
nand U1752 (N_1752,N_1401,N_1470);
nor U1753 (N_1753,N_1578,N_1420);
nand U1754 (N_1754,N_1403,N_1557);
or U1755 (N_1755,N_1571,N_1509);
and U1756 (N_1756,N_1593,N_1516);
nor U1757 (N_1757,N_1483,N_1518);
and U1758 (N_1758,N_1593,N_1493);
or U1759 (N_1759,N_1504,N_1417);
nand U1760 (N_1760,N_1430,N_1402);
nand U1761 (N_1761,N_1598,N_1514);
nor U1762 (N_1762,N_1417,N_1494);
nand U1763 (N_1763,N_1514,N_1434);
or U1764 (N_1764,N_1575,N_1561);
nand U1765 (N_1765,N_1526,N_1453);
nor U1766 (N_1766,N_1598,N_1405);
nand U1767 (N_1767,N_1468,N_1445);
nand U1768 (N_1768,N_1455,N_1438);
or U1769 (N_1769,N_1545,N_1496);
and U1770 (N_1770,N_1529,N_1549);
nor U1771 (N_1771,N_1490,N_1412);
nand U1772 (N_1772,N_1542,N_1572);
nand U1773 (N_1773,N_1516,N_1465);
nor U1774 (N_1774,N_1522,N_1525);
or U1775 (N_1775,N_1425,N_1553);
nand U1776 (N_1776,N_1563,N_1558);
nand U1777 (N_1777,N_1586,N_1493);
and U1778 (N_1778,N_1521,N_1563);
and U1779 (N_1779,N_1417,N_1557);
nand U1780 (N_1780,N_1528,N_1457);
nand U1781 (N_1781,N_1474,N_1534);
nand U1782 (N_1782,N_1521,N_1432);
nand U1783 (N_1783,N_1470,N_1536);
xor U1784 (N_1784,N_1583,N_1432);
and U1785 (N_1785,N_1575,N_1492);
xnor U1786 (N_1786,N_1574,N_1577);
and U1787 (N_1787,N_1505,N_1473);
xor U1788 (N_1788,N_1524,N_1513);
nor U1789 (N_1789,N_1573,N_1453);
or U1790 (N_1790,N_1512,N_1426);
nor U1791 (N_1791,N_1515,N_1446);
nor U1792 (N_1792,N_1492,N_1540);
nor U1793 (N_1793,N_1436,N_1574);
nor U1794 (N_1794,N_1435,N_1442);
nand U1795 (N_1795,N_1491,N_1426);
or U1796 (N_1796,N_1584,N_1405);
or U1797 (N_1797,N_1432,N_1469);
and U1798 (N_1798,N_1411,N_1566);
nor U1799 (N_1799,N_1452,N_1483);
or U1800 (N_1800,N_1785,N_1653);
or U1801 (N_1801,N_1772,N_1774);
nand U1802 (N_1802,N_1790,N_1639);
nand U1803 (N_1803,N_1642,N_1725);
or U1804 (N_1804,N_1770,N_1650);
or U1805 (N_1805,N_1655,N_1706);
nor U1806 (N_1806,N_1730,N_1726);
and U1807 (N_1807,N_1767,N_1610);
or U1808 (N_1808,N_1608,N_1683);
nor U1809 (N_1809,N_1736,N_1702);
and U1810 (N_1810,N_1751,N_1648);
nand U1811 (N_1811,N_1737,N_1668);
and U1812 (N_1812,N_1742,N_1631);
or U1813 (N_1813,N_1606,N_1659);
nand U1814 (N_1814,N_1618,N_1636);
nor U1815 (N_1815,N_1629,N_1695);
nor U1816 (N_1816,N_1732,N_1614);
nand U1817 (N_1817,N_1753,N_1764);
nand U1818 (N_1818,N_1626,N_1784);
nor U1819 (N_1819,N_1691,N_1722);
nor U1820 (N_1820,N_1609,N_1689);
and U1821 (N_1821,N_1690,N_1778);
and U1822 (N_1822,N_1611,N_1723);
nor U1823 (N_1823,N_1763,N_1708);
nor U1824 (N_1824,N_1715,N_1787);
nor U1825 (N_1825,N_1647,N_1757);
or U1826 (N_1826,N_1782,N_1605);
and U1827 (N_1827,N_1602,N_1781);
and U1828 (N_1828,N_1777,N_1704);
and U1829 (N_1829,N_1749,N_1612);
or U1830 (N_1830,N_1769,N_1638);
nand U1831 (N_1831,N_1740,N_1795);
nand U1832 (N_1832,N_1613,N_1646);
and U1833 (N_1833,N_1640,N_1630);
and U1834 (N_1834,N_1676,N_1745);
or U1835 (N_1835,N_1697,N_1643);
and U1836 (N_1836,N_1700,N_1645);
or U1837 (N_1837,N_1601,N_1658);
nor U1838 (N_1838,N_1665,N_1771);
or U1839 (N_1839,N_1661,N_1705);
or U1840 (N_1840,N_1780,N_1796);
nor U1841 (N_1841,N_1709,N_1733);
nor U1842 (N_1842,N_1670,N_1701);
nand U1843 (N_1843,N_1607,N_1652);
nor U1844 (N_1844,N_1651,N_1622);
nor U1845 (N_1845,N_1750,N_1746);
nor U1846 (N_1846,N_1687,N_1710);
nor U1847 (N_1847,N_1714,N_1776);
and U1848 (N_1848,N_1671,N_1719);
nor U1849 (N_1849,N_1624,N_1634);
nor U1850 (N_1850,N_1788,N_1698);
and U1851 (N_1851,N_1684,N_1762);
or U1852 (N_1852,N_1672,N_1669);
nand U1853 (N_1853,N_1625,N_1656);
nand U1854 (N_1854,N_1756,N_1734);
nand U1855 (N_1855,N_1724,N_1688);
nor U1856 (N_1856,N_1673,N_1752);
or U1857 (N_1857,N_1662,N_1693);
and U1858 (N_1858,N_1720,N_1616);
nor U1859 (N_1859,N_1694,N_1681);
or U1860 (N_1860,N_1677,N_1761);
nor U1861 (N_1861,N_1679,N_1604);
nand U1862 (N_1862,N_1786,N_1644);
and U1863 (N_1863,N_1703,N_1603);
nor U1864 (N_1864,N_1739,N_1664);
or U1865 (N_1865,N_1635,N_1741);
nor U1866 (N_1866,N_1711,N_1789);
and U1867 (N_1867,N_1729,N_1663);
and U1868 (N_1868,N_1727,N_1678);
nor U1869 (N_1869,N_1791,N_1798);
and U1870 (N_1870,N_1779,N_1696);
nor U1871 (N_1871,N_1738,N_1654);
or U1872 (N_1872,N_1660,N_1675);
xnor U1873 (N_1873,N_1667,N_1632);
or U1874 (N_1874,N_1773,N_1685);
or U1875 (N_1875,N_1623,N_1682);
nor U1876 (N_1876,N_1758,N_1619);
and U1877 (N_1877,N_1754,N_1657);
or U1878 (N_1878,N_1775,N_1759);
nand U1879 (N_1879,N_1600,N_1680);
or U1880 (N_1880,N_1755,N_1674);
or U1881 (N_1881,N_1686,N_1768);
and U1882 (N_1882,N_1721,N_1717);
nand U1883 (N_1883,N_1731,N_1743);
or U1884 (N_1884,N_1718,N_1707);
nand U1885 (N_1885,N_1628,N_1744);
and U1886 (N_1886,N_1783,N_1666);
or U1887 (N_1887,N_1627,N_1799);
nand U1888 (N_1888,N_1793,N_1712);
nor U1889 (N_1889,N_1641,N_1728);
nor U1890 (N_1890,N_1692,N_1699);
and U1891 (N_1891,N_1760,N_1620);
nand U1892 (N_1892,N_1713,N_1797);
or U1893 (N_1893,N_1637,N_1615);
nand U1894 (N_1894,N_1621,N_1792);
nor U1895 (N_1895,N_1735,N_1748);
nand U1896 (N_1896,N_1633,N_1649);
or U1897 (N_1897,N_1794,N_1747);
or U1898 (N_1898,N_1765,N_1716);
nand U1899 (N_1899,N_1617,N_1766);
and U1900 (N_1900,N_1634,N_1769);
nor U1901 (N_1901,N_1706,N_1623);
nor U1902 (N_1902,N_1656,N_1645);
nor U1903 (N_1903,N_1770,N_1632);
nand U1904 (N_1904,N_1655,N_1657);
nand U1905 (N_1905,N_1659,N_1645);
nor U1906 (N_1906,N_1767,N_1693);
and U1907 (N_1907,N_1771,N_1704);
nor U1908 (N_1908,N_1782,N_1700);
nand U1909 (N_1909,N_1713,N_1696);
nand U1910 (N_1910,N_1640,N_1780);
and U1911 (N_1911,N_1756,N_1626);
or U1912 (N_1912,N_1610,N_1772);
or U1913 (N_1913,N_1717,N_1757);
and U1914 (N_1914,N_1719,N_1658);
nand U1915 (N_1915,N_1677,N_1732);
nor U1916 (N_1916,N_1725,N_1616);
and U1917 (N_1917,N_1693,N_1710);
and U1918 (N_1918,N_1700,N_1704);
nand U1919 (N_1919,N_1783,N_1621);
nor U1920 (N_1920,N_1711,N_1753);
nand U1921 (N_1921,N_1668,N_1698);
and U1922 (N_1922,N_1718,N_1692);
and U1923 (N_1923,N_1748,N_1685);
nor U1924 (N_1924,N_1736,N_1783);
or U1925 (N_1925,N_1605,N_1669);
and U1926 (N_1926,N_1763,N_1797);
and U1927 (N_1927,N_1744,N_1634);
nor U1928 (N_1928,N_1680,N_1677);
nand U1929 (N_1929,N_1794,N_1781);
or U1930 (N_1930,N_1726,N_1671);
nand U1931 (N_1931,N_1788,N_1739);
or U1932 (N_1932,N_1694,N_1668);
nor U1933 (N_1933,N_1770,N_1691);
or U1934 (N_1934,N_1763,N_1706);
nor U1935 (N_1935,N_1684,N_1704);
and U1936 (N_1936,N_1667,N_1621);
nor U1937 (N_1937,N_1794,N_1664);
nand U1938 (N_1938,N_1630,N_1751);
nand U1939 (N_1939,N_1625,N_1714);
or U1940 (N_1940,N_1797,N_1777);
xnor U1941 (N_1941,N_1649,N_1640);
nand U1942 (N_1942,N_1788,N_1670);
nand U1943 (N_1943,N_1786,N_1626);
and U1944 (N_1944,N_1600,N_1621);
and U1945 (N_1945,N_1607,N_1773);
or U1946 (N_1946,N_1668,N_1742);
nand U1947 (N_1947,N_1670,N_1615);
and U1948 (N_1948,N_1613,N_1626);
or U1949 (N_1949,N_1706,N_1691);
and U1950 (N_1950,N_1737,N_1742);
nor U1951 (N_1951,N_1674,N_1757);
nor U1952 (N_1952,N_1657,N_1743);
and U1953 (N_1953,N_1614,N_1745);
or U1954 (N_1954,N_1755,N_1607);
and U1955 (N_1955,N_1726,N_1775);
nand U1956 (N_1956,N_1784,N_1719);
nand U1957 (N_1957,N_1627,N_1687);
nor U1958 (N_1958,N_1698,N_1740);
and U1959 (N_1959,N_1748,N_1614);
or U1960 (N_1960,N_1643,N_1640);
or U1961 (N_1961,N_1612,N_1619);
or U1962 (N_1962,N_1788,N_1718);
nand U1963 (N_1963,N_1652,N_1772);
and U1964 (N_1964,N_1723,N_1641);
nor U1965 (N_1965,N_1726,N_1780);
or U1966 (N_1966,N_1797,N_1678);
nand U1967 (N_1967,N_1760,N_1748);
nor U1968 (N_1968,N_1678,N_1734);
nand U1969 (N_1969,N_1709,N_1617);
or U1970 (N_1970,N_1703,N_1753);
or U1971 (N_1971,N_1685,N_1720);
nand U1972 (N_1972,N_1769,N_1619);
nand U1973 (N_1973,N_1638,N_1784);
or U1974 (N_1974,N_1602,N_1736);
or U1975 (N_1975,N_1641,N_1760);
and U1976 (N_1976,N_1753,N_1761);
nand U1977 (N_1977,N_1676,N_1604);
xor U1978 (N_1978,N_1709,N_1742);
and U1979 (N_1979,N_1733,N_1790);
or U1980 (N_1980,N_1617,N_1788);
nor U1981 (N_1981,N_1653,N_1752);
or U1982 (N_1982,N_1784,N_1662);
nand U1983 (N_1983,N_1699,N_1603);
or U1984 (N_1984,N_1600,N_1648);
and U1985 (N_1985,N_1782,N_1729);
nand U1986 (N_1986,N_1741,N_1757);
nand U1987 (N_1987,N_1711,N_1664);
or U1988 (N_1988,N_1743,N_1733);
xor U1989 (N_1989,N_1723,N_1634);
or U1990 (N_1990,N_1734,N_1680);
or U1991 (N_1991,N_1774,N_1633);
nor U1992 (N_1992,N_1722,N_1791);
nor U1993 (N_1993,N_1789,N_1670);
nand U1994 (N_1994,N_1614,N_1774);
and U1995 (N_1995,N_1789,N_1663);
and U1996 (N_1996,N_1689,N_1690);
nand U1997 (N_1997,N_1743,N_1709);
nand U1998 (N_1998,N_1647,N_1730);
or U1999 (N_1999,N_1679,N_1613);
nand U2000 (N_2000,N_1960,N_1995);
nand U2001 (N_2001,N_1868,N_1831);
nand U2002 (N_2002,N_1977,N_1805);
nand U2003 (N_2003,N_1850,N_1934);
nand U2004 (N_2004,N_1871,N_1908);
nand U2005 (N_2005,N_1856,N_1949);
nand U2006 (N_2006,N_1833,N_1828);
nor U2007 (N_2007,N_1975,N_1984);
and U2008 (N_2008,N_1978,N_1881);
and U2009 (N_2009,N_1826,N_1943);
nor U2010 (N_2010,N_1937,N_1815);
nor U2011 (N_2011,N_1955,N_1914);
or U2012 (N_2012,N_1883,N_1879);
nand U2013 (N_2013,N_1877,N_1812);
and U2014 (N_2014,N_1823,N_1911);
nor U2015 (N_2015,N_1971,N_1819);
or U2016 (N_2016,N_1865,N_1816);
nand U2017 (N_2017,N_1836,N_1994);
or U2018 (N_2018,N_1809,N_1966);
nor U2019 (N_2019,N_1933,N_1834);
nand U2020 (N_2020,N_1848,N_1800);
xnor U2021 (N_2021,N_1860,N_1974);
or U2022 (N_2022,N_1885,N_1916);
nand U2023 (N_2023,N_1876,N_1987);
nor U2024 (N_2024,N_1981,N_1963);
nor U2025 (N_2025,N_1982,N_1895);
and U2026 (N_2026,N_1864,N_1991);
or U2027 (N_2027,N_1878,N_1867);
nor U2028 (N_2028,N_1983,N_1938);
nor U2029 (N_2029,N_1939,N_1925);
nand U2030 (N_2030,N_1844,N_1909);
and U2031 (N_2031,N_1808,N_1958);
nand U2032 (N_2032,N_1891,N_1959);
or U2033 (N_2033,N_1892,N_1968);
and U2034 (N_2034,N_1967,N_1854);
nand U2035 (N_2035,N_1972,N_1957);
or U2036 (N_2036,N_1920,N_1946);
nand U2037 (N_2037,N_1950,N_1875);
nand U2038 (N_2038,N_1843,N_1842);
nand U2039 (N_2039,N_1952,N_1870);
nand U2040 (N_2040,N_1897,N_1874);
nor U2041 (N_2041,N_1979,N_1969);
nor U2042 (N_2042,N_1947,N_1830);
and U2043 (N_2043,N_1896,N_1941);
nand U2044 (N_2044,N_1917,N_1962);
nor U2045 (N_2045,N_1861,N_1820);
nor U2046 (N_2046,N_1999,N_1845);
nand U2047 (N_2047,N_1902,N_1997);
and U2048 (N_2048,N_1901,N_1998);
or U2049 (N_2049,N_1989,N_1829);
nand U2050 (N_2050,N_1910,N_1980);
or U2051 (N_2051,N_1927,N_1803);
nor U2052 (N_2052,N_1832,N_1898);
nor U2053 (N_2053,N_1930,N_1847);
or U2054 (N_2054,N_1890,N_1922);
and U2055 (N_2055,N_1837,N_1863);
and U2056 (N_2056,N_1900,N_1986);
nor U2057 (N_2057,N_1857,N_1818);
nor U2058 (N_2058,N_1841,N_1846);
nand U2059 (N_2059,N_1905,N_1953);
and U2060 (N_2060,N_1821,N_1906);
nand U2061 (N_2061,N_1965,N_1929);
nand U2062 (N_2062,N_1918,N_1976);
and U2063 (N_2063,N_1822,N_1804);
or U2064 (N_2064,N_1990,N_1899);
or U2065 (N_2065,N_1882,N_1889);
or U2066 (N_2066,N_1945,N_1907);
nor U2067 (N_2067,N_1942,N_1931);
nand U2068 (N_2068,N_1961,N_1807);
or U2069 (N_2069,N_1817,N_1887);
or U2070 (N_2070,N_1884,N_1851);
nand U2071 (N_2071,N_1964,N_1835);
nor U2072 (N_2072,N_1985,N_1888);
nor U2073 (N_2073,N_1903,N_1948);
and U2074 (N_2074,N_1810,N_1849);
nand U2075 (N_2075,N_1915,N_1919);
and U2076 (N_2076,N_1970,N_1904);
and U2077 (N_2077,N_1923,N_1813);
nor U2078 (N_2078,N_1973,N_1921);
nor U2079 (N_2079,N_1913,N_1924);
nand U2080 (N_2080,N_1802,N_1940);
nor U2081 (N_2081,N_1954,N_1839);
nor U2082 (N_2082,N_1806,N_1932);
nor U2083 (N_2083,N_1869,N_1853);
nand U2084 (N_2084,N_1951,N_1814);
nor U2085 (N_2085,N_1838,N_1893);
nand U2086 (N_2086,N_1956,N_1872);
or U2087 (N_2087,N_1912,N_1996);
or U2088 (N_2088,N_1825,N_1880);
nor U2089 (N_2089,N_1936,N_1840);
or U2090 (N_2090,N_1992,N_1859);
nand U2091 (N_2091,N_1827,N_1894);
and U2092 (N_2092,N_1886,N_1928);
nor U2093 (N_2093,N_1944,N_1858);
nor U2094 (N_2094,N_1855,N_1866);
or U2095 (N_2095,N_1811,N_1852);
nand U2096 (N_2096,N_1988,N_1824);
or U2097 (N_2097,N_1801,N_1862);
and U2098 (N_2098,N_1993,N_1926);
nand U2099 (N_2099,N_1873,N_1935);
and U2100 (N_2100,N_1964,N_1879);
and U2101 (N_2101,N_1993,N_1984);
or U2102 (N_2102,N_1820,N_1889);
nand U2103 (N_2103,N_1883,N_1816);
and U2104 (N_2104,N_1931,N_1973);
and U2105 (N_2105,N_1978,N_1970);
and U2106 (N_2106,N_1882,N_1916);
xnor U2107 (N_2107,N_1823,N_1920);
or U2108 (N_2108,N_1839,N_1901);
or U2109 (N_2109,N_1893,N_1843);
or U2110 (N_2110,N_1931,N_1856);
or U2111 (N_2111,N_1800,N_1833);
xnor U2112 (N_2112,N_1995,N_1848);
or U2113 (N_2113,N_1957,N_1909);
and U2114 (N_2114,N_1800,N_1858);
or U2115 (N_2115,N_1926,N_1880);
and U2116 (N_2116,N_1903,N_1829);
nor U2117 (N_2117,N_1978,N_1920);
nand U2118 (N_2118,N_1801,N_1934);
xor U2119 (N_2119,N_1893,N_1872);
and U2120 (N_2120,N_1897,N_1963);
or U2121 (N_2121,N_1844,N_1904);
nand U2122 (N_2122,N_1932,N_1877);
nor U2123 (N_2123,N_1887,N_1906);
nor U2124 (N_2124,N_1948,N_1832);
nand U2125 (N_2125,N_1892,N_1885);
nand U2126 (N_2126,N_1909,N_1867);
and U2127 (N_2127,N_1884,N_1855);
and U2128 (N_2128,N_1859,N_1996);
and U2129 (N_2129,N_1923,N_1836);
nor U2130 (N_2130,N_1820,N_1821);
and U2131 (N_2131,N_1849,N_1982);
nor U2132 (N_2132,N_1832,N_1859);
nor U2133 (N_2133,N_1993,N_1972);
nor U2134 (N_2134,N_1888,N_1828);
nand U2135 (N_2135,N_1884,N_1889);
nor U2136 (N_2136,N_1865,N_1982);
and U2137 (N_2137,N_1973,N_1883);
and U2138 (N_2138,N_1954,N_1983);
and U2139 (N_2139,N_1836,N_1870);
nand U2140 (N_2140,N_1981,N_1957);
and U2141 (N_2141,N_1851,N_1956);
or U2142 (N_2142,N_1982,N_1874);
or U2143 (N_2143,N_1973,N_1830);
or U2144 (N_2144,N_1959,N_1873);
nor U2145 (N_2145,N_1949,N_1867);
nor U2146 (N_2146,N_1925,N_1905);
or U2147 (N_2147,N_1821,N_1847);
and U2148 (N_2148,N_1955,N_1805);
nor U2149 (N_2149,N_1858,N_1940);
or U2150 (N_2150,N_1891,N_1923);
nand U2151 (N_2151,N_1984,N_1844);
nand U2152 (N_2152,N_1933,N_1884);
or U2153 (N_2153,N_1899,N_1840);
and U2154 (N_2154,N_1945,N_1993);
nand U2155 (N_2155,N_1867,N_1858);
and U2156 (N_2156,N_1899,N_1801);
and U2157 (N_2157,N_1992,N_1902);
or U2158 (N_2158,N_1898,N_1943);
nand U2159 (N_2159,N_1898,N_1937);
or U2160 (N_2160,N_1850,N_1835);
or U2161 (N_2161,N_1947,N_1951);
nand U2162 (N_2162,N_1999,N_1934);
or U2163 (N_2163,N_1870,N_1886);
nor U2164 (N_2164,N_1873,N_1842);
nor U2165 (N_2165,N_1863,N_1919);
and U2166 (N_2166,N_1905,N_1962);
or U2167 (N_2167,N_1948,N_1814);
nand U2168 (N_2168,N_1818,N_1884);
and U2169 (N_2169,N_1847,N_1882);
and U2170 (N_2170,N_1854,N_1881);
nand U2171 (N_2171,N_1842,N_1912);
or U2172 (N_2172,N_1820,N_1810);
nor U2173 (N_2173,N_1818,N_1805);
nand U2174 (N_2174,N_1999,N_1855);
xnor U2175 (N_2175,N_1900,N_1875);
nand U2176 (N_2176,N_1829,N_1863);
nor U2177 (N_2177,N_1915,N_1935);
nand U2178 (N_2178,N_1925,N_1864);
or U2179 (N_2179,N_1918,N_1940);
and U2180 (N_2180,N_1962,N_1845);
nor U2181 (N_2181,N_1916,N_1914);
nand U2182 (N_2182,N_1930,N_1953);
nand U2183 (N_2183,N_1975,N_1902);
or U2184 (N_2184,N_1835,N_1935);
and U2185 (N_2185,N_1857,N_1929);
nand U2186 (N_2186,N_1946,N_1931);
and U2187 (N_2187,N_1839,N_1917);
and U2188 (N_2188,N_1909,N_1913);
nor U2189 (N_2189,N_1898,N_1954);
or U2190 (N_2190,N_1978,N_1876);
nor U2191 (N_2191,N_1805,N_1857);
or U2192 (N_2192,N_1877,N_1996);
nand U2193 (N_2193,N_1899,N_1880);
nand U2194 (N_2194,N_1840,N_1950);
nand U2195 (N_2195,N_1971,N_1860);
nor U2196 (N_2196,N_1823,N_1928);
and U2197 (N_2197,N_1937,N_1916);
nor U2198 (N_2198,N_1809,N_1841);
nand U2199 (N_2199,N_1845,N_1924);
and U2200 (N_2200,N_2148,N_2077);
nor U2201 (N_2201,N_2033,N_2057);
nor U2202 (N_2202,N_2039,N_2037);
nor U2203 (N_2203,N_2147,N_2197);
nand U2204 (N_2204,N_2075,N_2023);
nand U2205 (N_2205,N_2119,N_2118);
nor U2206 (N_2206,N_2173,N_2103);
or U2207 (N_2207,N_2133,N_2064);
nor U2208 (N_2208,N_2088,N_2116);
nor U2209 (N_2209,N_2168,N_2069);
nand U2210 (N_2210,N_2150,N_2025);
and U2211 (N_2211,N_2007,N_2092);
nor U2212 (N_2212,N_2123,N_2099);
and U2213 (N_2213,N_2107,N_2014);
nor U2214 (N_2214,N_2142,N_2018);
nand U2215 (N_2215,N_2079,N_2054);
nand U2216 (N_2216,N_2113,N_2029);
nand U2217 (N_2217,N_2073,N_2026);
nor U2218 (N_2218,N_2082,N_2106);
or U2219 (N_2219,N_2078,N_2165);
nand U2220 (N_2220,N_2162,N_2087);
or U2221 (N_2221,N_2085,N_2108);
nor U2222 (N_2222,N_2056,N_2171);
nand U2223 (N_2223,N_2180,N_2086);
nand U2224 (N_2224,N_2098,N_2009);
nor U2225 (N_2225,N_2070,N_2144);
nor U2226 (N_2226,N_2112,N_2058);
and U2227 (N_2227,N_2021,N_2061);
nand U2228 (N_2228,N_2186,N_2158);
or U2229 (N_2229,N_2084,N_2024);
or U2230 (N_2230,N_2149,N_2019);
nand U2231 (N_2231,N_2076,N_2128);
nand U2232 (N_2232,N_2141,N_2050);
nor U2233 (N_2233,N_2028,N_2072);
nand U2234 (N_2234,N_2191,N_2071);
nor U2235 (N_2235,N_2174,N_2059);
and U2236 (N_2236,N_2164,N_2111);
nand U2237 (N_2237,N_2110,N_2109);
nand U2238 (N_2238,N_2187,N_2134);
nor U2239 (N_2239,N_2005,N_2089);
and U2240 (N_2240,N_2065,N_2042);
nor U2241 (N_2241,N_2045,N_2012);
nand U2242 (N_2242,N_2008,N_2146);
nor U2243 (N_2243,N_2167,N_2083);
or U2244 (N_2244,N_2135,N_2176);
nand U2245 (N_2245,N_2169,N_2055);
nor U2246 (N_2246,N_2184,N_2105);
or U2247 (N_2247,N_2122,N_2038);
or U2248 (N_2248,N_2027,N_2049);
nand U2249 (N_2249,N_2172,N_2091);
xor U2250 (N_2250,N_2017,N_2129);
nor U2251 (N_2251,N_2190,N_2137);
and U2252 (N_2252,N_2153,N_2094);
nor U2253 (N_2253,N_2003,N_2127);
or U2254 (N_2254,N_2192,N_2011);
nor U2255 (N_2255,N_2062,N_2080);
or U2256 (N_2256,N_2090,N_2124);
or U2257 (N_2257,N_2048,N_2081);
nor U2258 (N_2258,N_2178,N_2117);
and U2259 (N_2259,N_2068,N_2053);
and U2260 (N_2260,N_2160,N_2036);
or U2261 (N_2261,N_2022,N_2004);
and U2262 (N_2262,N_2161,N_2030);
nor U2263 (N_2263,N_2002,N_2035);
nor U2264 (N_2264,N_2047,N_2031);
or U2265 (N_2265,N_2051,N_2060);
nor U2266 (N_2266,N_2183,N_2126);
and U2267 (N_2267,N_2163,N_2015);
or U2268 (N_2268,N_2151,N_2010);
or U2269 (N_2269,N_2114,N_2074);
and U2270 (N_2270,N_2120,N_2121);
nand U2271 (N_2271,N_2188,N_2181);
nand U2272 (N_2272,N_2041,N_2020);
and U2273 (N_2273,N_2189,N_2034);
or U2274 (N_2274,N_2140,N_2096);
nand U2275 (N_2275,N_2177,N_2155);
nor U2276 (N_2276,N_2199,N_2066);
or U2277 (N_2277,N_2138,N_2166);
nand U2278 (N_2278,N_2040,N_2093);
nor U2279 (N_2279,N_2139,N_2154);
and U2280 (N_2280,N_2179,N_2193);
or U2281 (N_2281,N_2195,N_2046);
or U2282 (N_2282,N_2016,N_2063);
or U2283 (N_2283,N_2001,N_2157);
or U2284 (N_2284,N_2013,N_2175);
nor U2285 (N_2285,N_2143,N_2104);
nand U2286 (N_2286,N_2136,N_2156);
and U2287 (N_2287,N_2044,N_2067);
nand U2288 (N_2288,N_2097,N_2170);
or U2289 (N_2289,N_2125,N_2100);
or U2290 (N_2290,N_2130,N_2198);
and U2291 (N_2291,N_2052,N_2132);
or U2292 (N_2292,N_2131,N_2152);
or U2293 (N_2293,N_2182,N_2101);
or U2294 (N_2294,N_2194,N_2159);
nor U2295 (N_2295,N_2102,N_2000);
nor U2296 (N_2296,N_2095,N_2196);
and U2297 (N_2297,N_2145,N_2032);
nor U2298 (N_2298,N_2043,N_2006);
or U2299 (N_2299,N_2185,N_2115);
and U2300 (N_2300,N_2168,N_2013);
nand U2301 (N_2301,N_2101,N_2160);
nand U2302 (N_2302,N_2119,N_2124);
nor U2303 (N_2303,N_2015,N_2017);
nor U2304 (N_2304,N_2133,N_2124);
nor U2305 (N_2305,N_2167,N_2088);
and U2306 (N_2306,N_2024,N_2131);
and U2307 (N_2307,N_2053,N_2149);
nand U2308 (N_2308,N_2143,N_2004);
or U2309 (N_2309,N_2160,N_2078);
or U2310 (N_2310,N_2042,N_2106);
and U2311 (N_2311,N_2070,N_2028);
and U2312 (N_2312,N_2186,N_2119);
or U2313 (N_2313,N_2177,N_2018);
or U2314 (N_2314,N_2184,N_2147);
nor U2315 (N_2315,N_2003,N_2171);
or U2316 (N_2316,N_2174,N_2070);
nand U2317 (N_2317,N_2088,N_2053);
nor U2318 (N_2318,N_2042,N_2165);
nor U2319 (N_2319,N_2166,N_2160);
nor U2320 (N_2320,N_2006,N_2020);
nand U2321 (N_2321,N_2073,N_2133);
nand U2322 (N_2322,N_2104,N_2176);
or U2323 (N_2323,N_2044,N_2122);
or U2324 (N_2324,N_2125,N_2108);
nand U2325 (N_2325,N_2054,N_2101);
nor U2326 (N_2326,N_2033,N_2122);
nand U2327 (N_2327,N_2050,N_2022);
and U2328 (N_2328,N_2010,N_2020);
xor U2329 (N_2329,N_2130,N_2181);
and U2330 (N_2330,N_2189,N_2156);
nand U2331 (N_2331,N_2147,N_2082);
and U2332 (N_2332,N_2047,N_2104);
nor U2333 (N_2333,N_2056,N_2015);
or U2334 (N_2334,N_2063,N_2159);
or U2335 (N_2335,N_2171,N_2080);
nand U2336 (N_2336,N_2031,N_2139);
nand U2337 (N_2337,N_2103,N_2078);
and U2338 (N_2338,N_2113,N_2151);
nor U2339 (N_2339,N_2162,N_2067);
or U2340 (N_2340,N_2018,N_2006);
and U2341 (N_2341,N_2055,N_2130);
and U2342 (N_2342,N_2173,N_2185);
nor U2343 (N_2343,N_2109,N_2028);
and U2344 (N_2344,N_2158,N_2031);
and U2345 (N_2345,N_2036,N_2129);
nor U2346 (N_2346,N_2133,N_2027);
or U2347 (N_2347,N_2135,N_2154);
nor U2348 (N_2348,N_2036,N_2166);
or U2349 (N_2349,N_2028,N_2107);
nor U2350 (N_2350,N_2088,N_2015);
nor U2351 (N_2351,N_2091,N_2157);
nand U2352 (N_2352,N_2155,N_2169);
nand U2353 (N_2353,N_2118,N_2071);
nor U2354 (N_2354,N_2036,N_2183);
nand U2355 (N_2355,N_2048,N_2112);
nand U2356 (N_2356,N_2017,N_2135);
nor U2357 (N_2357,N_2094,N_2125);
or U2358 (N_2358,N_2084,N_2160);
or U2359 (N_2359,N_2157,N_2190);
nand U2360 (N_2360,N_2159,N_2184);
nand U2361 (N_2361,N_2076,N_2139);
nor U2362 (N_2362,N_2025,N_2160);
nor U2363 (N_2363,N_2148,N_2110);
nand U2364 (N_2364,N_2125,N_2191);
or U2365 (N_2365,N_2018,N_2044);
nor U2366 (N_2366,N_2119,N_2097);
and U2367 (N_2367,N_2139,N_2185);
and U2368 (N_2368,N_2072,N_2088);
nor U2369 (N_2369,N_2076,N_2037);
or U2370 (N_2370,N_2198,N_2140);
nor U2371 (N_2371,N_2125,N_2091);
or U2372 (N_2372,N_2106,N_2091);
nand U2373 (N_2373,N_2080,N_2020);
nand U2374 (N_2374,N_2016,N_2111);
and U2375 (N_2375,N_2057,N_2114);
nor U2376 (N_2376,N_2155,N_2140);
and U2377 (N_2377,N_2054,N_2063);
nor U2378 (N_2378,N_2063,N_2013);
or U2379 (N_2379,N_2149,N_2087);
nand U2380 (N_2380,N_2164,N_2024);
nand U2381 (N_2381,N_2042,N_2067);
or U2382 (N_2382,N_2081,N_2117);
nand U2383 (N_2383,N_2038,N_2053);
nand U2384 (N_2384,N_2067,N_2007);
or U2385 (N_2385,N_2121,N_2073);
and U2386 (N_2386,N_2033,N_2025);
nand U2387 (N_2387,N_2087,N_2056);
and U2388 (N_2388,N_2059,N_2073);
and U2389 (N_2389,N_2143,N_2181);
and U2390 (N_2390,N_2184,N_2055);
or U2391 (N_2391,N_2005,N_2049);
and U2392 (N_2392,N_2150,N_2006);
xor U2393 (N_2393,N_2160,N_2070);
or U2394 (N_2394,N_2183,N_2068);
and U2395 (N_2395,N_2192,N_2151);
nor U2396 (N_2396,N_2114,N_2166);
and U2397 (N_2397,N_2051,N_2097);
or U2398 (N_2398,N_2147,N_2056);
and U2399 (N_2399,N_2194,N_2167);
and U2400 (N_2400,N_2254,N_2389);
xnor U2401 (N_2401,N_2352,N_2358);
and U2402 (N_2402,N_2342,N_2206);
nor U2403 (N_2403,N_2256,N_2375);
or U2404 (N_2404,N_2399,N_2397);
nand U2405 (N_2405,N_2211,N_2380);
or U2406 (N_2406,N_2229,N_2286);
nand U2407 (N_2407,N_2393,N_2388);
nor U2408 (N_2408,N_2290,N_2232);
and U2409 (N_2409,N_2316,N_2268);
and U2410 (N_2410,N_2287,N_2249);
or U2411 (N_2411,N_2215,N_2225);
nand U2412 (N_2412,N_2362,N_2324);
or U2413 (N_2413,N_2282,N_2213);
nand U2414 (N_2414,N_2207,N_2216);
and U2415 (N_2415,N_2212,N_2303);
nand U2416 (N_2416,N_2340,N_2251);
nor U2417 (N_2417,N_2291,N_2366);
and U2418 (N_2418,N_2355,N_2265);
nand U2419 (N_2419,N_2387,N_2244);
or U2420 (N_2420,N_2293,N_2237);
and U2421 (N_2421,N_2261,N_2264);
and U2422 (N_2422,N_2329,N_2377);
or U2423 (N_2423,N_2337,N_2271);
and U2424 (N_2424,N_2378,N_2334);
and U2425 (N_2425,N_2279,N_2349);
nand U2426 (N_2426,N_2273,N_2353);
nand U2427 (N_2427,N_2319,N_2208);
nand U2428 (N_2428,N_2392,N_2347);
nor U2429 (N_2429,N_2336,N_2344);
nand U2430 (N_2430,N_2266,N_2236);
or U2431 (N_2431,N_2361,N_2385);
or U2432 (N_2432,N_2328,N_2354);
nor U2433 (N_2433,N_2220,N_2257);
and U2434 (N_2434,N_2255,N_2322);
nand U2435 (N_2435,N_2373,N_2310);
or U2436 (N_2436,N_2226,N_2368);
and U2437 (N_2437,N_2351,N_2267);
nor U2438 (N_2438,N_2296,N_2292);
nand U2439 (N_2439,N_2314,N_2350);
nand U2440 (N_2440,N_2395,N_2396);
and U2441 (N_2441,N_2201,N_2248);
and U2442 (N_2442,N_2218,N_2259);
and U2443 (N_2443,N_2348,N_2357);
and U2444 (N_2444,N_2363,N_2243);
nor U2445 (N_2445,N_2376,N_2203);
and U2446 (N_2446,N_2384,N_2302);
or U2447 (N_2447,N_2240,N_2394);
xnor U2448 (N_2448,N_2332,N_2305);
xnor U2449 (N_2449,N_2230,N_2253);
nor U2450 (N_2450,N_2325,N_2200);
nor U2451 (N_2451,N_2374,N_2239);
nor U2452 (N_2452,N_2383,N_2234);
or U2453 (N_2453,N_2227,N_2306);
and U2454 (N_2454,N_2275,N_2326);
or U2455 (N_2455,N_2263,N_2204);
and U2456 (N_2456,N_2331,N_2258);
nor U2457 (N_2457,N_2221,N_2307);
or U2458 (N_2458,N_2346,N_2369);
nor U2459 (N_2459,N_2311,N_2330);
nor U2460 (N_2460,N_2224,N_2360);
nand U2461 (N_2461,N_2245,N_2323);
nor U2462 (N_2462,N_2301,N_2294);
nor U2463 (N_2463,N_2313,N_2338);
or U2464 (N_2464,N_2210,N_2214);
nor U2465 (N_2465,N_2315,N_2231);
nand U2466 (N_2466,N_2367,N_2308);
nand U2467 (N_2467,N_2382,N_2235);
and U2468 (N_2468,N_2284,N_2247);
and U2469 (N_2469,N_2312,N_2327);
and U2470 (N_2470,N_2223,N_2285);
nor U2471 (N_2471,N_2370,N_2379);
nor U2472 (N_2472,N_2297,N_2242);
and U2473 (N_2473,N_2250,N_2217);
nand U2474 (N_2474,N_2298,N_2365);
nand U2475 (N_2475,N_2278,N_2364);
or U2476 (N_2476,N_2280,N_2391);
nand U2477 (N_2477,N_2289,N_2345);
and U2478 (N_2478,N_2241,N_2343);
or U2479 (N_2479,N_2269,N_2317);
nand U2480 (N_2480,N_2288,N_2277);
nand U2481 (N_2481,N_2270,N_2274);
and U2482 (N_2482,N_2276,N_2262);
nand U2483 (N_2483,N_2335,N_2246);
or U2484 (N_2484,N_2372,N_2295);
and U2485 (N_2485,N_2381,N_2386);
nand U2486 (N_2486,N_2371,N_2333);
or U2487 (N_2487,N_2205,N_2252);
nand U2488 (N_2488,N_2272,N_2321);
and U2489 (N_2489,N_2356,N_2320);
or U2490 (N_2490,N_2309,N_2304);
and U2491 (N_2491,N_2209,N_2390);
nor U2492 (N_2492,N_2339,N_2398);
and U2493 (N_2493,N_2283,N_2300);
or U2494 (N_2494,N_2219,N_2318);
nand U2495 (N_2495,N_2228,N_2202);
nor U2496 (N_2496,N_2222,N_2281);
nor U2497 (N_2497,N_2233,N_2238);
and U2498 (N_2498,N_2260,N_2299);
nand U2499 (N_2499,N_2341,N_2359);
or U2500 (N_2500,N_2220,N_2328);
nor U2501 (N_2501,N_2380,N_2254);
nor U2502 (N_2502,N_2272,N_2279);
nand U2503 (N_2503,N_2395,N_2397);
nor U2504 (N_2504,N_2311,N_2203);
or U2505 (N_2505,N_2215,N_2337);
and U2506 (N_2506,N_2284,N_2299);
or U2507 (N_2507,N_2339,N_2305);
or U2508 (N_2508,N_2253,N_2373);
or U2509 (N_2509,N_2378,N_2344);
and U2510 (N_2510,N_2379,N_2345);
and U2511 (N_2511,N_2368,N_2209);
and U2512 (N_2512,N_2206,N_2345);
and U2513 (N_2513,N_2288,N_2387);
nand U2514 (N_2514,N_2362,N_2260);
nand U2515 (N_2515,N_2388,N_2337);
nand U2516 (N_2516,N_2282,N_2311);
and U2517 (N_2517,N_2224,N_2257);
or U2518 (N_2518,N_2296,N_2368);
nand U2519 (N_2519,N_2237,N_2300);
or U2520 (N_2520,N_2393,N_2230);
nand U2521 (N_2521,N_2208,N_2355);
and U2522 (N_2522,N_2288,N_2385);
nand U2523 (N_2523,N_2363,N_2220);
or U2524 (N_2524,N_2334,N_2336);
nor U2525 (N_2525,N_2393,N_2383);
nand U2526 (N_2526,N_2381,N_2266);
nor U2527 (N_2527,N_2394,N_2389);
and U2528 (N_2528,N_2250,N_2316);
and U2529 (N_2529,N_2229,N_2206);
nor U2530 (N_2530,N_2377,N_2245);
and U2531 (N_2531,N_2389,N_2369);
nand U2532 (N_2532,N_2252,N_2340);
or U2533 (N_2533,N_2334,N_2343);
nor U2534 (N_2534,N_2265,N_2288);
nand U2535 (N_2535,N_2218,N_2241);
and U2536 (N_2536,N_2376,N_2347);
or U2537 (N_2537,N_2355,N_2224);
or U2538 (N_2538,N_2230,N_2269);
nand U2539 (N_2539,N_2392,N_2201);
nor U2540 (N_2540,N_2355,N_2322);
and U2541 (N_2541,N_2387,N_2245);
nand U2542 (N_2542,N_2252,N_2282);
and U2543 (N_2543,N_2349,N_2252);
nor U2544 (N_2544,N_2207,N_2274);
or U2545 (N_2545,N_2237,N_2295);
nor U2546 (N_2546,N_2348,N_2242);
nor U2547 (N_2547,N_2377,N_2242);
xor U2548 (N_2548,N_2344,N_2241);
nand U2549 (N_2549,N_2265,N_2247);
and U2550 (N_2550,N_2368,N_2373);
nor U2551 (N_2551,N_2266,N_2394);
nor U2552 (N_2552,N_2261,N_2343);
or U2553 (N_2553,N_2244,N_2243);
and U2554 (N_2554,N_2248,N_2242);
nand U2555 (N_2555,N_2208,N_2266);
xnor U2556 (N_2556,N_2274,N_2243);
nor U2557 (N_2557,N_2229,N_2310);
nand U2558 (N_2558,N_2295,N_2210);
and U2559 (N_2559,N_2370,N_2323);
nand U2560 (N_2560,N_2305,N_2341);
or U2561 (N_2561,N_2231,N_2299);
nor U2562 (N_2562,N_2372,N_2344);
or U2563 (N_2563,N_2368,N_2221);
and U2564 (N_2564,N_2393,N_2216);
nor U2565 (N_2565,N_2289,N_2208);
and U2566 (N_2566,N_2337,N_2206);
nor U2567 (N_2567,N_2374,N_2244);
or U2568 (N_2568,N_2378,N_2370);
or U2569 (N_2569,N_2298,N_2261);
and U2570 (N_2570,N_2392,N_2397);
xor U2571 (N_2571,N_2369,N_2342);
nand U2572 (N_2572,N_2370,N_2207);
and U2573 (N_2573,N_2229,N_2232);
and U2574 (N_2574,N_2333,N_2313);
or U2575 (N_2575,N_2284,N_2313);
nor U2576 (N_2576,N_2244,N_2335);
nor U2577 (N_2577,N_2341,N_2387);
nand U2578 (N_2578,N_2397,N_2375);
nand U2579 (N_2579,N_2296,N_2384);
and U2580 (N_2580,N_2201,N_2236);
nand U2581 (N_2581,N_2293,N_2372);
and U2582 (N_2582,N_2215,N_2270);
or U2583 (N_2583,N_2272,N_2244);
or U2584 (N_2584,N_2368,N_2281);
nand U2585 (N_2585,N_2394,N_2235);
or U2586 (N_2586,N_2286,N_2320);
nor U2587 (N_2587,N_2312,N_2344);
and U2588 (N_2588,N_2215,N_2258);
and U2589 (N_2589,N_2323,N_2281);
and U2590 (N_2590,N_2298,N_2381);
and U2591 (N_2591,N_2389,N_2251);
or U2592 (N_2592,N_2399,N_2280);
nor U2593 (N_2593,N_2345,N_2396);
nor U2594 (N_2594,N_2388,N_2336);
and U2595 (N_2595,N_2243,N_2380);
or U2596 (N_2596,N_2308,N_2239);
or U2597 (N_2597,N_2200,N_2331);
nor U2598 (N_2598,N_2324,N_2281);
nand U2599 (N_2599,N_2207,N_2259);
or U2600 (N_2600,N_2450,N_2456);
nand U2601 (N_2601,N_2493,N_2571);
nand U2602 (N_2602,N_2479,N_2464);
nor U2603 (N_2603,N_2512,N_2484);
or U2604 (N_2604,N_2596,N_2449);
nand U2605 (N_2605,N_2532,N_2429);
or U2606 (N_2606,N_2516,N_2415);
or U2607 (N_2607,N_2416,N_2508);
nor U2608 (N_2608,N_2530,N_2547);
nand U2609 (N_2609,N_2550,N_2436);
nand U2610 (N_2610,N_2579,N_2455);
nand U2611 (N_2611,N_2564,N_2406);
or U2612 (N_2612,N_2466,N_2561);
and U2613 (N_2613,N_2536,N_2457);
and U2614 (N_2614,N_2551,N_2408);
and U2615 (N_2615,N_2409,N_2447);
and U2616 (N_2616,N_2446,N_2510);
nand U2617 (N_2617,N_2505,N_2474);
or U2618 (N_2618,N_2437,N_2475);
or U2619 (N_2619,N_2470,N_2595);
or U2620 (N_2620,N_2472,N_2435);
and U2621 (N_2621,N_2578,N_2552);
nand U2622 (N_2622,N_2545,N_2478);
nand U2623 (N_2623,N_2507,N_2423);
nor U2624 (N_2624,N_2485,N_2468);
nor U2625 (N_2625,N_2521,N_2407);
nand U2626 (N_2626,N_2525,N_2534);
nor U2627 (N_2627,N_2402,N_2425);
and U2628 (N_2628,N_2588,N_2556);
nand U2629 (N_2629,N_2565,N_2494);
and U2630 (N_2630,N_2569,N_2433);
and U2631 (N_2631,N_2482,N_2465);
and U2632 (N_2632,N_2483,N_2454);
or U2633 (N_2633,N_2487,N_2517);
or U2634 (N_2634,N_2555,N_2461);
nor U2635 (N_2635,N_2424,N_2419);
and U2636 (N_2636,N_2497,N_2524);
nor U2637 (N_2637,N_2543,N_2528);
or U2638 (N_2638,N_2432,N_2553);
nor U2639 (N_2639,N_2593,N_2502);
nor U2640 (N_2640,N_2498,N_2513);
or U2641 (N_2641,N_2583,N_2486);
nor U2642 (N_2642,N_2539,N_2599);
or U2643 (N_2643,N_2591,N_2412);
nor U2644 (N_2644,N_2538,N_2434);
nor U2645 (N_2645,N_2480,N_2584);
or U2646 (N_2646,N_2560,N_2557);
and U2647 (N_2647,N_2469,N_2404);
and U2648 (N_2648,N_2540,N_2506);
nor U2649 (N_2649,N_2413,N_2535);
or U2650 (N_2650,N_2411,N_2541);
or U2651 (N_2651,N_2586,N_2581);
and U2652 (N_2652,N_2471,N_2439);
or U2653 (N_2653,N_2488,N_2597);
or U2654 (N_2654,N_2577,N_2430);
nor U2655 (N_2655,N_2421,N_2589);
nand U2656 (N_2656,N_2573,N_2438);
or U2657 (N_2657,N_2458,N_2473);
xor U2658 (N_2658,N_2522,N_2549);
nor U2659 (N_2659,N_2527,N_2417);
nand U2660 (N_2660,N_2533,N_2453);
nor U2661 (N_2661,N_2598,N_2537);
and U2662 (N_2662,N_2567,N_2519);
and U2663 (N_2663,N_2520,N_2570);
or U2664 (N_2664,N_2448,N_2499);
and U2665 (N_2665,N_2559,N_2492);
or U2666 (N_2666,N_2529,N_2503);
xnor U2667 (N_2667,N_2490,N_2477);
or U2668 (N_2668,N_2544,N_2428);
nor U2669 (N_2669,N_2427,N_2523);
nand U2670 (N_2670,N_2509,N_2476);
xor U2671 (N_2671,N_2426,N_2500);
nor U2672 (N_2672,N_2592,N_2548);
or U2673 (N_2673,N_2400,N_2442);
or U2674 (N_2674,N_2460,N_2403);
nor U2675 (N_2675,N_2459,N_2414);
or U2676 (N_2676,N_2568,N_2518);
and U2677 (N_2677,N_2531,N_2580);
nor U2678 (N_2678,N_2467,N_2572);
nor U2679 (N_2679,N_2590,N_2511);
or U2680 (N_2680,N_2422,N_2431);
and U2681 (N_2681,N_2587,N_2576);
nor U2682 (N_2682,N_2481,N_2582);
or U2683 (N_2683,N_2566,N_2526);
nand U2684 (N_2684,N_2405,N_2444);
or U2685 (N_2685,N_2445,N_2441);
or U2686 (N_2686,N_2410,N_2575);
nand U2687 (N_2687,N_2443,N_2585);
or U2688 (N_2688,N_2515,N_2420);
nor U2689 (N_2689,N_2554,N_2451);
or U2690 (N_2690,N_2440,N_2491);
and U2691 (N_2691,N_2563,N_2594);
and U2692 (N_2692,N_2452,N_2558);
nor U2693 (N_2693,N_2501,N_2401);
nand U2694 (N_2694,N_2463,N_2574);
and U2695 (N_2695,N_2504,N_2514);
nand U2696 (N_2696,N_2489,N_2546);
nor U2697 (N_2697,N_2542,N_2462);
nor U2698 (N_2698,N_2562,N_2418);
and U2699 (N_2699,N_2495,N_2496);
and U2700 (N_2700,N_2592,N_2572);
and U2701 (N_2701,N_2487,N_2568);
and U2702 (N_2702,N_2534,N_2477);
nor U2703 (N_2703,N_2427,N_2518);
and U2704 (N_2704,N_2483,N_2460);
nand U2705 (N_2705,N_2495,N_2515);
nand U2706 (N_2706,N_2523,N_2570);
nor U2707 (N_2707,N_2522,N_2562);
or U2708 (N_2708,N_2483,N_2427);
or U2709 (N_2709,N_2571,N_2551);
and U2710 (N_2710,N_2562,N_2421);
or U2711 (N_2711,N_2492,N_2411);
nor U2712 (N_2712,N_2539,N_2591);
nand U2713 (N_2713,N_2400,N_2424);
nand U2714 (N_2714,N_2448,N_2487);
nor U2715 (N_2715,N_2413,N_2426);
nor U2716 (N_2716,N_2437,N_2503);
and U2717 (N_2717,N_2472,N_2509);
nor U2718 (N_2718,N_2547,N_2470);
or U2719 (N_2719,N_2500,N_2586);
nand U2720 (N_2720,N_2478,N_2495);
nand U2721 (N_2721,N_2479,N_2550);
and U2722 (N_2722,N_2590,N_2562);
nand U2723 (N_2723,N_2477,N_2467);
nor U2724 (N_2724,N_2573,N_2542);
or U2725 (N_2725,N_2579,N_2421);
nor U2726 (N_2726,N_2453,N_2558);
and U2727 (N_2727,N_2471,N_2566);
and U2728 (N_2728,N_2511,N_2457);
nand U2729 (N_2729,N_2512,N_2446);
nand U2730 (N_2730,N_2587,N_2491);
and U2731 (N_2731,N_2593,N_2503);
nor U2732 (N_2732,N_2418,N_2497);
nand U2733 (N_2733,N_2502,N_2420);
nor U2734 (N_2734,N_2421,N_2451);
nor U2735 (N_2735,N_2463,N_2515);
nand U2736 (N_2736,N_2499,N_2566);
nand U2737 (N_2737,N_2489,N_2419);
nor U2738 (N_2738,N_2488,N_2529);
nor U2739 (N_2739,N_2443,N_2404);
or U2740 (N_2740,N_2447,N_2415);
nand U2741 (N_2741,N_2596,N_2401);
nand U2742 (N_2742,N_2502,N_2531);
nor U2743 (N_2743,N_2563,N_2560);
and U2744 (N_2744,N_2599,N_2579);
nor U2745 (N_2745,N_2429,N_2489);
or U2746 (N_2746,N_2559,N_2570);
nor U2747 (N_2747,N_2483,N_2580);
nor U2748 (N_2748,N_2495,N_2570);
and U2749 (N_2749,N_2424,N_2576);
nor U2750 (N_2750,N_2584,N_2436);
or U2751 (N_2751,N_2553,N_2582);
and U2752 (N_2752,N_2583,N_2498);
nor U2753 (N_2753,N_2416,N_2503);
nor U2754 (N_2754,N_2472,N_2565);
or U2755 (N_2755,N_2572,N_2492);
and U2756 (N_2756,N_2430,N_2567);
nand U2757 (N_2757,N_2476,N_2424);
nor U2758 (N_2758,N_2402,N_2479);
nand U2759 (N_2759,N_2595,N_2542);
or U2760 (N_2760,N_2474,N_2478);
xnor U2761 (N_2761,N_2463,N_2504);
and U2762 (N_2762,N_2499,N_2581);
nor U2763 (N_2763,N_2563,N_2491);
nor U2764 (N_2764,N_2446,N_2562);
or U2765 (N_2765,N_2478,N_2590);
and U2766 (N_2766,N_2454,N_2400);
nor U2767 (N_2767,N_2556,N_2443);
nand U2768 (N_2768,N_2582,N_2402);
and U2769 (N_2769,N_2412,N_2567);
nand U2770 (N_2770,N_2539,N_2433);
and U2771 (N_2771,N_2553,N_2450);
or U2772 (N_2772,N_2415,N_2502);
nand U2773 (N_2773,N_2465,N_2546);
or U2774 (N_2774,N_2566,N_2451);
or U2775 (N_2775,N_2447,N_2595);
nand U2776 (N_2776,N_2557,N_2542);
or U2777 (N_2777,N_2525,N_2475);
or U2778 (N_2778,N_2560,N_2439);
and U2779 (N_2779,N_2444,N_2542);
nor U2780 (N_2780,N_2550,N_2445);
or U2781 (N_2781,N_2444,N_2410);
nand U2782 (N_2782,N_2422,N_2560);
nor U2783 (N_2783,N_2544,N_2465);
nand U2784 (N_2784,N_2553,N_2504);
or U2785 (N_2785,N_2425,N_2595);
nor U2786 (N_2786,N_2401,N_2595);
nor U2787 (N_2787,N_2599,N_2418);
or U2788 (N_2788,N_2441,N_2403);
or U2789 (N_2789,N_2547,N_2450);
or U2790 (N_2790,N_2555,N_2409);
nand U2791 (N_2791,N_2423,N_2445);
or U2792 (N_2792,N_2533,N_2413);
or U2793 (N_2793,N_2513,N_2441);
and U2794 (N_2794,N_2578,N_2448);
nand U2795 (N_2795,N_2484,N_2416);
and U2796 (N_2796,N_2527,N_2588);
nor U2797 (N_2797,N_2458,N_2447);
and U2798 (N_2798,N_2451,N_2490);
nor U2799 (N_2799,N_2485,N_2546);
or U2800 (N_2800,N_2783,N_2647);
nand U2801 (N_2801,N_2685,N_2778);
and U2802 (N_2802,N_2747,N_2788);
nor U2803 (N_2803,N_2682,N_2694);
nand U2804 (N_2804,N_2710,N_2611);
or U2805 (N_2805,N_2753,N_2626);
nor U2806 (N_2806,N_2603,N_2708);
nand U2807 (N_2807,N_2734,N_2727);
nor U2808 (N_2808,N_2616,N_2619);
nor U2809 (N_2809,N_2777,N_2683);
or U2810 (N_2810,N_2772,N_2787);
or U2811 (N_2811,N_2775,N_2608);
and U2812 (N_2812,N_2666,N_2638);
nor U2813 (N_2813,N_2659,N_2706);
nand U2814 (N_2814,N_2718,N_2670);
or U2815 (N_2815,N_2711,N_2679);
or U2816 (N_2816,N_2776,N_2764);
or U2817 (N_2817,N_2742,N_2672);
or U2818 (N_2818,N_2652,N_2690);
and U2819 (N_2819,N_2739,N_2761);
or U2820 (N_2820,N_2635,N_2600);
nand U2821 (N_2821,N_2766,N_2741);
nand U2822 (N_2822,N_2673,N_2634);
nand U2823 (N_2823,N_2760,N_2722);
nor U2824 (N_2824,N_2693,N_2724);
nand U2825 (N_2825,N_2657,N_2612);
xor U2826 (N_2826,N_2756,N_2779);
and U2827 (N_2827,N_2643,N_2656);
nand U2828 (N_2828,N_2660,N_2786);
and U2829 (N_2829,N_2709,N_2618);
nand U2830 (N_2830,N_2642,N_2798);
nand U2831 (N_2831,N_2719,N_2607);
and U2832 (N_2832,N_2799,N_2781);
or U2833 (N_2833,N_2624,N_2684);
nand U2834 (N_2834,N_2645,N_2767);
and U2835 (N_2835,N_2692,N_2791);
or U2836 (N_2836,N_2629,N_2630);
nor U2837 (N_2837,N_2768,N_2697);
nand U2838 (N_2838,N_2644,N_2623);
or U2839 (N_2839,N_2758,N_2707);
nor U2840 (N_2840,N_2733,N_2649);
nor U2841 (N_2841,N_2646,N_2754);
or U2842 (N_2842,N_2606,N_2789);
and U2843 (N_2843,N_2704,N_2723);
or U2844 (N_2844,N_2633,N_2691);
or U2845 (N_2845,N_2662,N_2701);
or U2846 (N_2846,N_2762,N_2713);
or U2847 (N_2847,N_2625,N_2726);
or U2848 (N_2848,N_2628,N_2774);
or U2849 (N_2849,N_2702,N_2757);
nand U2850 (N_2850,N_2636,N_2716);
nand U2851 (N_2851,N_2770,N_2627);
nand U2852 (N_2852,N_2655,N_2769);
nand U2853 (N_2853,N_2720,N_2780);
nor U2854 (N_2854,N_2700,N_2740);
or U2855 (N_2855,N_2792,N_2759);
nor U2856 (N_2856,N_2632,N_2746);
or U2857 (N_2857,N_2677,N_2782);
nand U2858 (N_2858,N_2639,N_2689);
nor U2859 (N_2859,N_2668,N_2663);
nand U2860 (N_2860,N_2745,N_2640);
and U2861 (N_2861,N_2650,N_2654);
and U2862 (N_2862,N_2771,N_2610);
or U2863 (N_2863,N_2744,N_2653);
and U2864 (N_2864,N_2658,N_2750);
or U2865 (N_2865,N_2614,N_2617);
nor U2866 (N_2866,N_2748,N_2631);
or U2867 (N_2867,N_2669,N_2696);
nor U2868 (N_2868,N_2687,N_2797);
nand U2869 (N_2869,N_2695,N_2763);
nand U2870 (N_2870,N_2728,N_2648);
and U2871 (N_2871,N_2731,N_2736);
and U2872 (N_2872,N_2605,N_2686);
and U2873 (N_2873,N_2671,N_2681);
nand U2874 (N_2874,N_2680,N_2637);
and U2875 (N_2875,N_2609,N_2621);
nand U2876 (N_2876,N_2651,N_2712);
nor U2877 (N_2877,N_2604,N_2773);
or U2878 (N_2878,N_2676,N_2743);
xnor U2879 (N_2879,N_2674,N_2738);
or U2880 (N_2880,N_2749,N_2675);
nand U2881 (N_2881,N_2732,N_2667);
nand U2882 (N_2882,N_2703,N_2735);
and U2883 (N_2883,N_2665,N_2698);
or U2884 (N_2884,N_2622,N_2794);
or U2885 (N_2885,N_2790,N_2688);
nor U2886 (N_2886,N_2601,N_2784);
nor U2887 (N_2887,N_2714,N_2678);
or U2888 (N_2888,N_2661,N_2699);
nor U2889 (N_2889,N_2729,N_2751);
and U2890 (N_2890,N_2705,N_2795);
or U2891 (N_2891,N_2725,N_2793);
and U2892 (N_2892,N_2715,N_2615);
nand U2893 (N_2893,N_2752,N_2755);
nor U2894 (N_2894,N_2730,N_2765);
or U2895 (N_2895,N_2613,N_2641);
or U2896 (N_2896,N_2664,N_2602);
nor U2897 (N_2897,N_2717,N_2620);
nor U2898 (N_2898,N_2796,N_2721);
or U2899 (N_2899,N_2737,N_2785);
or U2900 (N_2900,N_2669,N_2605);
or U2901 (N_2901,N_2657,N_2772);
and U2902 (N_2902,N_2744,N_2752);
and U2903 (N_2903,N_2779,N_2612);
nor U2904 (N_2904,N_2691,N_2690);
or U2905 (N_2905,N_2679,N_2752);
and U2906 (N_2906,N_2783,N_2689);
nor U2907 (N_2907,N_2755,N_2799);
nand U2908 (N_2908,N_2782,N_2649);
nand U2909 (N_2909,N_2633,N_2652);
nand U2910 (N_2910,N_2620,N_2694);
or U2911 (N_2911,N_2700,N_2647);
nor U2912 (N_2912,N_2605,N_2798);
nor U2913 (N_2913,N_2679,N_2773);
or U2914 (N_2914,N_2615,N_2690);
nand U2915 (N_2915,N_2753,N_2762);
nand U2916 (N_2916,N_2615,N_2737);
nand U2917 (N_2917,N_2637,N_2796);
or U2918 (N_2918,N_2654,N_2625);
nand U2919 (N_2919,N_2691,N_2642);
or U2920 (N_2920,N_2659,N_2703);
nor U2921 (N_2921,N_2617,N_2686);
and U2922 (N_2922,N_2636,N_2602);
nor U2923 (N_2923,N_2789,N_2735);
nand U2924 (N_2924,N_2740,N_2798);
nor U2925 (N_2925,N_2766,N_2795);
nor U2926 (N_2926,N_2787,N_2668);
nand U2927 (N_2927,N_2705,N_2675);
nor U2928 (N_2928,N_2754,N_2641);
nand U2929 (N_2929,N_2690,N_2637);
nor U2930 (N_2930,N_2626,N_2645);
and U2931 (N_2931,N_2769,N_2760);
or U2932 (N_2932,N_2771,N_2659);
nor U2933 (N_2933,N_2614,N_2682);
nor U2934 (N_2934,N_2674,N_2711);
nor U2935 (N_2935,N_2791,N_2734);
nand U2936 (N_2936,N_2611,N_2627);
nor U2937 (N_2937,N_2645,N_2654);
and U2938 (N_2938,N_2642,N_2641);
nand U2939 (N_2939,N_2690,N_2728);
nor U2940 (N_2940,N_2606,N_2758);
nor U2941 (N_2941,N_2766,N_2698);
nand U2942 (N_2942,N_2668,N_2732);
nand U2943 (N_2943,N_2608,N_2633);
and U2944 (N_2944,N_2621,N_2699);
nor U2945 (N_2945,N_2798,N_2705);
or U2946 (N_2946,N_2671,N_2678);
nand U2947 (N_2947,N_2706,N_2709);
and U2948 (N_2948,N_2675,N_2695);
nor U2949 (N_2949,N_2616,N_2728);
or U2950 (N_2950,N_2640,N_2671);
nand U2951 (N_2951,N_2733,N_2706);
or U2952 (N_2952,N_2669,N_2651);
nor U2953 (N_2953,N_2714,N_2690);
nand U2954 (N_2954,N_2634,N_2639);
and U2955 (N_2955,N_2652,N_2636);
nand U2956 (N_2956,N_2701,N_2787);
nor U2957 (N_2957,N_2781,N_2735);
nand U2958 (N_2958,N_2704,N_2677);
and U2959 (N_2959,N_2725,N_2792);
xor U2960 (N_2960,N_2748,N_2688);
nor U2961 (N_2961,N_2642,N_2647);
and U2962 (N_2962,N_2728,N_2766);
nor U2963 (N_2963,N_2652,N_2638);
and U2964 (N_2964,N_2634,N_2628);
nand U2965 (N_2965,N_2744,N_2773);
nand U2966 (N_2966,N_2775,N_2635);
nand U2967 (N_2967,N_2759,N_2777);
nor U2968 (N_2968,N_2715,N_2683);
or U2969 (N_2969,N_2702,N_2639);
or U2970 (N_2970,N_2798,N_2661);
nor U2971 (N_2971,N_2638,N_2663);
and U2972 (N_2972,N_2668,N_2616);
or U2973 (N_2973,N_2786,N_2621);
or U2974 (N_2974,N_2667,N_2703);
nand U2975 (N_2975,N_2705,N_2625);
xor U2976 (N_2976,N_2786,N_2666);
nand U2977 (N_2977,N_2789,N_2675);
or U2978 (N_2978,N_2669,N_2600);
and U2979 (N_2979,N_2661,N_2712);
and U2980 (N_2980,N_2783,N_2687);
nand U2981 (N_2981,N_2741,N_2610);
or U2982 (N_2982,N_2658,N_2798);
or U2983 (N_2983,N_2702,N_2631);
nor U2984 (N_2984,N_2653,N_2703);
nor U2985 (N_2985,N_2615,N_2679);
nor U2986 (N_2986,N_2654,N_2600);
nor U2987 (N_2987,N_2747,N_2783);
nor U2988 (N_2988,N_2744,N_2759);
nor U2989 (N_2989,N_2736,N_2605);
nand U2990 (N_2990,N_2624,N_2751);
nor U2991 (N_2991,N_2660,N_2626);
nand U2992 (N_2992,N_2712,N_2792);
nor U2993 (N_2993,N_2672,N_2604);
nand U2994 (N_2994,N_2714,N_2780);
nor U2995 (N_2995,N_2650,N_2776);
and U2996 (N_2996,N_2637,N_2730);
nor U2997 (N_2997,N_2664,N_2748);
nand U2998 (N_2998,N_2669,N_2719);
and U2999 (N_2999,N_2609,N_2643);
or UO_0 (O_0,N_2945,N_2879);
or UO_1 (O_1,N_2955,N_2963);
nor UO_2 (O_2,N_2834,N_2915);
nand UO_3 (O_3,N_2953,N_2921);
nand UO_4 (O_4,N_2992,N_2925);
or UO_5 (O_5,N_2987,N_2971);
and UO_6 (O_6,N_2996,N_2979);
nand UO_7 (O_7,N_2844,N_2958);
nand UO_8 (O_8,N_2899,N_2885);
or UO_9 (O_9,N_2954,N_2962);
and UO_10 (O_10,N_2824,N_2827);
and UO_11 (O_11,N_2914,N_2803);
nand UO_12 (O_12,N_2883,N_2820);
nor UO_13 (O_13,N_2943,N_2970);
nand UO_14 (O_14,N_2822,N_2946);
nand UO_15 (O_15,N_2806,N_2852);
and UO_16 (O_16,N_2947,N_2931);
and UO_17 (O_17,N_2912,N_2810);
nand UO_18 (O_18,N_2805,N_2850);
and UO_19 (O_19,N_2841,N_2929);
nor UO_20 (O_20,N_2981,N_2892);
nor UO_21 (O_21,N_2870,N_2895);
and UO_22 (O_22,N_2887,N_2873);
nand UO_23 (O_23,N_2864,N_2871);
nand UO_24 (O_24,N_2878,N_2817);
or UO_25 (O_25,N_2994,N_2837);
or UO_26 (O_26,N_2959,N_2869);
or UO_27 (O_27,N_2927,N_2934);
nor UO_28 (O_28,N_2818,N_2941);
and UO_29 (O_29,N_2865,N_2966);
nor UO_30 (O_30,N_2976,N_2831);
and UO_31 (O_31,N_2825,N_2889);
nor UO_32 (O_32,N_2975,N_2893);
nand UO_33 (O_33,N_2863,N_2972);
nand UO_34 (O_34,N_2967,N_2860);
or UO_35 (O_35,N_2986,N_2876);
or UO_36 (O_36,N_2957,N_2922);
and UO_37 (O_37,N_2882,N_2886);
or UO_38 (O_38,N_2830,N_2872);
nand UO_39 (O_39,N_2916,N_2801);
and UO_40 (O_40,N_2853,N_2989);
or UO_41 (O_41,N_2815,N_2884);
or UO_42 (O_42,N_2898,N_2950);
nor UO_43 (O_43,N_2812,N_2874);
nor UO_44 (O_44,N_2948,N_2867);
and UO_45 (O_45,N_2926,N_2999);
nor UO_46 (O_46,N_2909,N_2951);
nor UO_47 (O_47,N_2988,N_2908);
nor UO_48 (O_48,N_2930,N_2832);
or UO_49 (O_49,N_2888,N_2849);
or UO_50 (O_50,N_2845,N_2932);
or UO_51 (O_51,N_2809,N_2969);
and UO_52 (O_52,N_2851,N_2983);
nor UO_53 (O_53,N_2814,N_2942);
nand UO_54 (O_54,N_2808,N_2890);
nand UO_55 (O_55,N_2924,N_2859);
and UO_56 (O_56,N_2990,N_2843);
or UO_57 (O_57,N_2868,N_2855);
nor UO_58 (O_58,N_2928,N_2984);
or UO_59 (O_59,N_2811,N_2866);
and UO_60 (O_60,N_2857,N_2802);
nor UO_61 (O_61,N_2816,N_2939);
or UO_62 (O_62,N_2875,N_2901);
nor UO_63 (O_63,N_2919,N_2840);
xor UO_64 (O_64,N_2842,N_2880);
nand UO_65 (O_65,N_2847,N_2923);
and UO_66 (O_66,N_2833,N_2935);
or UO_67 (O_67,N_2861,N_2897);
and UO_68 (O_68,N_2985,N_2968);
nand UO_69 (O_69,N_2913,N_2838);
xnor UO_70 (O_70,N_2804,N_2944);
nand UO_71 (O_71,N_2911,N_2839);
nand UO_72 (O_72,N_2993,N_2961);
nor UO_73 (O_73,N_2906,N_2991);
nand UO_74 (O_74,N_2854,N_2862);
and UO_75 (O_75,N_2938,N_2918);
nand UO_76 (O_76,N_2982,N_2933);
nand UO_77 (O_77,N_2952,N_2836);
nor UO_78 (O_78,N_2905,N_2917);
and UO_79 (O_79,N_2826,N_2856);
or UO_80 (O_80,N_2960,N_2846);
nand UO_81 (O_81,N_2813,N_2964);
and UO_82 (O_82,N_2800,N_2907);
and UO_83 (O_83,N_2823,N_2891);
or UO_84 (O_84,N_2858,N_2910);
and UO_85 (O_85,N_2903,N_2877);
nor UO_86 (O_86,N_2936,N_2904);
or UO_87 (O_87,N_2965,N_2900);
or UO_88 (O_88,N_2819,N_2973);
and UO_89 (O_89,N_2835,N_2920);
or UO_90 (O_90,N_2974,N_2881);
nand UO_91 (O_91,N_2997,N_2894);
and UO_92 (O_92,N_2995,N_2949);
and UO_93 (O_93,N_2978,N_2807);
nand UO_94 (O_94,N_2977,N_2829);
and UO_95 (O_95,N_2998,N_2821);
or UO_96 (O_96,N_2940,N_2980);
nor UO_97 (O_97,N_2896,N_2848);
nor UO_98 (O_98,N_2902,N_2956);
or UO_99 (O_99,N_2828,N_2937);
or UO_100 (O_100,N_2813,N_2961);
nand UO_101 (O_101,N_2857,N_2897);
nor UO_102 (O_102,N_2998,N_2879);
nor UO_103 (O_103,N_2926,N_2854);
nor UO_104 (O_104,N_2916,N_2984);
or UO_105 (O_105,N_2822,N_2947);
nor UO_106 (O_106,N_2820,N_2918);
nand UO_107 (O_107,N_2897,N_2864);
or UO_108 (O_108,N_2858,N_2808);
nor UO_109 (O_109,N_2840,N_2987);
nor UO_110 (O_110,N_2913,N_2887);
nor UO_111 (O_111,N_2872,N_2996);
or UO_112 (O_112,N_2953,N_2843);
and UO_113 (O_113,N_2822,N_2802);
nor UO_114 (O_114,N_2945,N_2871);
or UO_115 (O_115,N_2911,N_2807);
and UO_116 (O_116,N_2867,N_2889);
nor UO_117 (O_117,N_2844,N_2863);
xor UO_118 (O_118,N_2875,N_2915);
or UO_119 (O_119,N_2901,N_2802);
or UO_120 (O_120,N_2977,N_2868);
or UO_121 (O_121,N_2949,N_2903);
nand UO_122 (O_122,N_2829,N_2951);
or UO_123 (O_123,N_2927,N_2999);
and UO_124 (O_124,N_2828,N_2947);
and UO_125 (O_125,N_2888,N_2997);
nor UO_126 (O_126,N_2860,N_2824);
nor UO_127 (O_127,N_2935,N_2898);
or UO_128 (O_128,N_2986,N_2920);
or UO_129 (O_129,N_2933,N_2950);
nand UO_130 (O_130,N_2873,N_2998);
or UO_131 (O_131,N_2957,N_2978);
nand UO_132 (O_132,N_2889,N_2863);
nand UO_133 (O_133,N_2881,N_2834);
nor UO_134 (O_134,N_2825,N_2856);
and UO_135 (O_135,N_2918,N_2969);
nor UO_136 (O_136,N_2914,N_2875);
or UO_137 (O_137,N_2880,N_2910);
nor UO_138 (O_138,N_2826,N_2985);
nor UO_139 (O_139,N_2978,N_2928);
and UO_140 (O_140,N_2825,N_2822);
and UO_141 (O_141,N_2891,N_2852);
and UO_142 (O_142,N_2824,N_2972);
and UO_143 (O_143,N_2974,N_2891);
or UO_144 (O_144,N_2901,N_2864);
nand UO_145 (O_145,N_2815,N_2835);
and UO_146 (O_146,N_2902,N_2853);
nand UO_147 (O_147,N_2979,N_2988);
or UO_148 (O_148,N_2860,N_2960);
or UO_149 (O_149,N_2910,N_2987);
and UO_150 (O_150,N_2951,N_2927);
and UO_151 (O_151,N_2970,N_2917);
and UO_152 (O_152,N_2834,N_2957);
and UO_153 (O_153,N_2851,N_2964);
and UO_154 (O_154,N_2884,N_2928);
or UO_155 (O_155,N_2818,N_2963);
nor UO_156 (O_156,N_2898,N_2926);
nor UO_157 (O_157,N_2928,N_2802);
and UO_158 (O_158,N_2920,N_2829);
or UO_159 (O_159,N_2812,N_2933);
nand UO_160 (O_160,N_2927,N_2970);
nor UO_161 (O_161,N_2900,N_2850);
nor UO_162 (O_162,N_2919,N_2888);
nand UO_163 (O_163,N_2915,N_2910);
or UO_164 (O_164,N_2814,N_2906);
nand UO_165 (O_165,N_2981,N_2898);
nand UO_166 (O_166,N_2883,N_2870);
and UO_167 (O_167,N_2927,N_2980);
nand UO_168 (O_168,N_2973,N_2967);
or UO_169 (O_169,N_2936,N_2991);
nor UO_170 (O_170,N_2955,N_2826);
and UO_171 (O_171,N_2991,N_2959);
and UO_172 (O_172,N_2871,N_2805);
nand UO_173 (O_173,N_2900,N_2877);
or UO_174 (O_174,N_2954,N_2993);
nor UO_175 (O_175,N_2995,N_2885);
nand UO_176 (O_176,N_2809,N_2886);
nor UO_177 (O_177,N_2838,N_2963);
and UO_178 (O_178,N_2853,N_2830);
or UO_179 (O_179,N_2845,N_2934);
xnor UO_180 (O_180,N_2932,N_2999);
and UO_181 (O_181,N_2812,N_2851);
and UO_182 (O_182,N_2953,N_2830);
or UO_183 (O_183,N_2914,N_2804);
or UO_184 (O_184,N_2865,N_2963);
nand UO_185 (O_185,N_2837,N_2875);
and UO_186 (O_186,N_2833,N_2888);
or UO_187 (O_187,N_2878,N_2970);
and UO_188 (O_188,N_2894,N_2963);
and UO_189 (O_189,N_2886,N_2822);
nor UO_190 (O_190,N_2983,N_2986);
or UO_191 (O_191,N_2945,N_2844);
xnor UO_192 (O_192,N_2872,N_2896);
nand UO_193 (O_193,N_2877,N_2994);
nand UO_194 (O_194,N_2864,N_2982);
nor UO_195 (O_195,N_2870,N_2882);
nand UO_196 (O_196,N_2896,N_2941);
and UO_197 (O_197,N_2807,N_2810);
nand UO_198 (O_198,N_2833,N_2934);
nor UO_199 (O_199,N_2990,N_2880);
or UO_200 (O_200,N_2875,N_2831);
and UO_201 (O_201,N_2917,N_2857);
or UO_202 (O_202,N_2962,N_2859);
and UO_203 (O_203,N_2946,N_2943);
nand UO_204 (O_204,N_2942,N_2863);
or UO_205 (O_205,N_2831,N_2898);
nor UO_206 (O_206,N_2845,N_2858);
or UO_207 (O_207,N_2886,N_2954);
or UO_208 (O_208,N_2978,N_2832);
and UO_209 (O_209,N_2974,N_2933);
nor UO_210 (O_210,N_2865,N_2933);
nand UO_211 (O_211,N_2992,N_2958);
nor UO_212 (O_212,N_2804,N_2893);
nor UO_213 (O_213,N_2808,N_2896);
and UO_214 (O_214,N_2990,N_2955);
nor UO_215 (O_215,N_2866,N_2948);
nor UO_216 (O_216,N_2985,N_2863);
and UO_217 (O_217,N_2907,N_2936);
and UO_218 (O_218,N_2800,N_2848);
or UO_219 (O_219,N_2800,N_2951);
or UO_220 (O_220,N_2858,N_2824);
or UO_221 (O_221,N_2990,N_2807);
or UO_222 (O_222,N_2958,N_2987);
nand UO_223 (O_223,N_2922,N_2832);
nor UO_224 (O_224,N_2822,N_2972);
nor UO_225 (O_225,N_2933,N_2921);
nor UO_226 (O_226,N_2992,N_2853);
and UO_227 (O_227,N_2926,N_2864);
nor UO_228 (O_228,N_2924,N_2978);
and UO_229 (O_229,N_2933,N_2996);
and UO_230 (O_230,N_2905,N_2873);
or UO_231 (O_231,N_2935,N_2861);
and UO_232 (O_232,N_2811,N_2996);
nor UO_233 (O_233,N_2924,N_2833);
nand UO_234 (O_234,N_2862,N_2859);
nand UO_235 (O_235,N_2976,N_2827);
nand UO_236 (O_236,N_2888,N_2975);
and UO_237 (O_237,N_2966,N_2891);
and UO_238 (O_238,N_2814,N_2929);
nand UO_239 (O_239,N_2886,N_2837);
and UO_240 (O_240,N_2907,N_2856);
xor UO_241 (O_241,N_2834,N_2826);
or UO_242 (O_242,N_2862,N_2967);
and UO_243 (O_243,N_2818,N_2893);
nand UO_244 (O_244,N_2920,N_2850);
nor UO_245 (O_245,N_2829,N_2891);
or UO_246 (O_246,N_2909,N_2948);
and UO_247 (O_247,N_2932,N_2974);
and UO_248 (O_248,N_2881,N_2938);
and UO_249 (O_249,N_2847,N_2858);
or UO_250 (O_250,N_2917,N_2937);
nor UO_251 (O_251,N_2827,N_2902);
nand UO_252 (O_252,N_2870,N_2913);
or UO_253 (O_253,N_2938,N_2877);
nand UO_254 (O_254,N_2812,N_2925);
or UO_255 (O_255,N_2985,N_2825);
nand UO_256 (O_256,N_2801,N_2964);
nor UO_257 (O_257,N_2853,N_2969);
and UO_258 (O_258,N_2948,N_2933);
nand UO_259 (O_259,N_2920,N_2839);
or UO_260 (O_260,N_2895,N_2968);
nand UO_261 (O_261,N_2904,N_2881);
or UO_262 (O_262,N_2800,N_2908);
nor UO_263 (O_263,N_2991,N_2954);
or UO_264 (O_264,N_2911,N_2930);
nand UO_265 (O_265,N_2836,N_2810);
nor UO_266 (O_266,N_2985,N_2883);
or UO_267 (O_267,N_2942,N_2977);
nor UO_268 (O_268,N_2869,N_2858);
nand UO_269 (O_269,N_2819,N_2927);
nor UO_270 (O_270,N_2937,N_2986);
nand UO_271 (O_271,N_2844,N_2999);
nor UO_272 (O_272,N_2863,N_2869);
or UO_273 (O_273,N_2910,N_2888);
and UO_274 (O_274,N_2888,N_2809);
and UO_275 (O_275,N_2945,N_2878);
nor UO_276 (O_276,N_2833,N_2979);
and UO_277 (O_277,N_2987,N_2983);
or UO_278 (O_278,N_2850,N_2871);
and UO_279 (O_279,N_2819,N_2995);
or UO_280 (O_280,N_2809,N_2808);
and UO_281 (O_281,N_2935,N_2966);
or UO_282 (O_282,N_2868,N_2982);
and UO_283 (O_283,N_2965,N_2888);
and UO_284 (O_284,N_2837,N_2825);
or UO_285 (O_285,N_2966,N_2862);
or UO_286 (O_286,N_2899,N_2862);
nand UO_287 (O_287,N_2867,N_2947);
or UO_288 (O_288,N_2809,N_2821);
xnor UO_289 (O_289,N_2946,N_2804);
or UO_290 (O_290,N_2903,N_2848);
nand UO_291 (O_291,N_2963,N_2851);
xnor UO_292 (O_292,N_2865,N_2914);
or UO_293 (O_293,N_2974,N_2840);
or UO_294 (O_294,N_2830,N_2963);
and UO_295 (O_295,N_2819,N_2980);
nand UO_296 (O_296,N_2963,N_2959);
or UO_297 (O_297,N_2912,N_2852);
or UO_298 (O_298,N_2810,N_2986);
or UO_299 (O_299,N_2886,N_2834);
and UO_300 (O_300,N_2869,N_2829);
or UO_301 (O_301,N_2991,N_2824);
nand UO_302 (O_302,N_2945,N_2896);
nor UO_303 (O_303,N_2942,N_2837);
nor UO_304 (O_304,N_2860,N_2977);
nor UO_305 (O_305,N_2899,N_2916);
nand UO_306 (O_306,N_2974,N_2909);
and UO_307 (O_307,N_2938,N_2855);
or UO_308 (O_308,N_2935,N_2997);
nor UO_309 (O_309,N_2931,N_2803);
and UO_310 (O_310,N_2849,N_2901);
and UO_311 (O_311,N_2894,N_2942);
nor UO_312 (O_312,N_2924,N_2820);
nor UO_313 (O_313,N_2948,N_2860);
nor UO_314 (O_314,N_2963,N_2987);
or UO_315 (O_315,N_2877,N_2817);
nand UO_316 (O_316,N_2858,N_2948);
or UO_317 (O_317,N_2881,N_2948);
or UO_318 (O_318,N_2845,N_2989);
nand UO_319 (O_319,N_2898,N_2914);
nor UO_320 (O_320,N_2860,N_2922);
nand UO_321 (O_321,N_2848,N_2997);
and UO_322 (O_322,N_2928,N_2971);
nand UO_323 (O_323,N_2876,N_2912);
nor UO_324 (O_324,N_2853,N_2893);
and UO_325 (O_325,N_2975,N_2897);
nand UO_326 (O_326,N_2965,N_2892);
or UO_327 (O_327,N_2815,N_2933);
and UO_328 (O_328,N_2983,N_2919);
nand UO_329 (O_329,N_2847,N_2974);
or UO_330 (O_330,N_2976,N_2912);
and UO_331 (O_331,N_2902,N_2849);
nand UO_332 (O_332,N_2852,N_2913);
or UO_333 (O_333,N_2915,N_2840);
or UO_334 (O_334,N_2959,N_2835);
and UO_335 (O_335,N_2894,N_2981);
and UO_336 (O_336,N_2833,N_2906);
nor UO_337 (O_337,N_2903,N_2952);
nor UO_338 (O_338,N_2854,N_2847);
or UO_339 (O_339,N_2916,N_2811);
nor UO_340 (O_340,N_2898,N_2822);
nand UO_341 (O_341,N_2807,N_2983);
nor UO_342 (O_342,N_2877,N_2929);
or UO_343 (O_343,N_2972,N_2939);
nand UO_344 (O_344,N_2978,N_2947);
and UO_345 (O_345,N_2949,N_2864);
nand UO_346 (O_346,N_2982,N_2889);
nand UO_347 (O_347,N_2855,N_2964);
nor UO_348 (O_348,N_2902,N_2840);
and UO_349 (O_349,N_2898,N_2909);
or UO_350 (O_350,N_2967,N_2947);
nor UO_351 (O_351,N_2958,N_2921);
and UO_352 (O_352,N_2878,N_2956);
and UO_353 (O_353,N_2802,N_2801);
or UO_354 (O_354,N_2831,N_2868);
and UO_355 (O_355,N_2857,N_2852);
or UO_356 (O_356,N_2971,N_2804);
nor UO_357 (O_357,N_2850,N_2951);
and UO_358 (O_358,N_2991,N_2849);
or UO_359 (O_359,N_2939,N_2959);
nor UO_360 (O_360,N_2839,N_2975);
nor UO_361 (O_361,N_2991,N_2974);
nand UO_362 (O_362,N_2859,N_2917);
nor UO_363 (O_363,N_2935,N_2924);
nand UO_364 (O_364,N_2941,N_2856);
nor UO_365 (O_365,N_2895,N_2962);
nand UO_366 (O_366,N_2956,N_2830);
nor UO_367 (O_367,N_2937,N_2898);
and UO_368 (O_368,N_2819,N_2803);
nor UO_369 (O_369,N_2897,N_2840);
or UO_370 (O_370,N_2964,N_2937);
nand UO_371 (O_371,N_2975,N_2986);
nor UO_372 (O_372,N_2949,N_2931);
and UO_373 (O_373,N_2890,N_2957);
nor UO_374 (O_374,N_2881,N_2871);
nor UO_375 (O_375,N_2969,N_2929);
or UO_376 (O_376,N_2923,N_2872);
nor UO_377 (O_377,N_2976,N_2925);
nor UO_378 (O_378,N_2893,N_2908);
and UO_379 (O_379,N_2822,N_2851);
or UO_380 (O_380,N_2959,N_2867);
nor UO_381 (O_381,N_2867,N_2844);
nand UO_382 (O_382,N_2976,N_2870);
nor UO_383 (O_383,N_2965,N_2905);
nand UO_384 (O_384,N_2866,N_2951);
or UO_385 (O_385,N_2863,N_2807);
and UO_386 (O_386,N_2889,N_2994);
or UO_387 (O_387,N_2963,N_2864);
and UO_388 (O_388,N_2882,N_2917);
nand UO_389 (O_389,N_2896,N_2865);
or UO_390 (O_390,N_2920,N_2802);
or UO_391 (O_391,N_2800,N_2865);
or UO_392 (O_392,N_2854,N_2831);
nand UO_393 (O_393,N_2946,N_2936);
nor UO_394 (O_394,N_2825,N_2964);
nand UO_395 (O_395,N_2936,N_2842);
and UO_396 (O_396,N_2801,N_2941);
nor UO_397 (O_397,N_2847,N_2916);
and UO_398 (O_398,N_2862,N_2888);
nor UO_399 (O_399,N_2938,N_2998);
nor UO_400 (O_400,N_2961,N_2850);
and UO_401 (O_401,N_2904,N_2947);
nand UO_402 (O_402,N_2816,N_2990);
nand UO_403 (O_403,N_2889,N_2910);
nor UO_404 (O_404,N_2932,N_2956);
and UO_405 (O_405,N_2874,N_2859);
nand UO_406 (O_406,N_2985,N_2974);
and UO_407 (O_407,N_2800,N_2963);
nand UO_408 (O_408,N_2980,N_2903);
and UO_409 (O_409,N_2876,N_2874);
or UO_410 (O_410,N_2893,N_2868);
and UO_411 (O_411,N_2830,N_2974);
and UO_412 (O_412,N_2883,N_2981);
nor UO_413 (O_413,N_2846,N_2946);
nor UO_414 (O_414,N_2949,N_2871);
nor UO_415 (O_415,N_2987,N_2850);
nor UO_416 (O_416,N_2864,N_2878);
and UO_417 (O_417,N_2834,N_2945);
or UO_418 (O_418,N_2974,N_2837);
or UO_419 (O_419,N_2948,N_2942);
nand UO_420 (O_420,N_2899,N_2841);
nor UO_421 (O_421,N_2937,N_2877);
nand UO_422 (O_422,N_2898,N_2953);
nor UO_423 (O_423,N_2885,N_2803);
nor UO_424 (O_424,N_2861,N_2927);
nor UO_425 (O_425,N_2889,N_2829);
and UO_426 (O_426,N_2858,N_2984);
nor UO_427 (O_427,N_2945,N_2960);
nand UO_428 (O_428,N_2986,N_2823);
or UO_429 (O_429,N_2835,N_2901);
xnor UO_430 (O_430,N_2987,N_2970);
and UO_431 (O_431,N_2962,N_2975);
nand UO_432 (O_432,N_2981,N_2905);
nor UO_433 (O_433,N_2828,N_2948);
or UO_434 (O_434,N_2823,N_2966);
or UO_435 (O_435,N_2988,N_2971);
and UO_436 (O_436,N_2912,N_2948);
and UO_437 (O_437,N_2931,N_2878);
or UO_438 (O_438,N_2970,N_2895);
nor UO_439 (O_439,N_2827,N_2826);
nor UO_440 (O_440,N_2940,N_2955);
and UO_441 (O_441,N_2883,N_2887);
or UO_442 (O_442,N_2819,N_2829);
nand UO_443 (O_443,N_2893,N_2841);
and UO_444 (O_444,N_2962,N_2868);
nor UO_445 (O_445,N_2930,N_2917);
or UO_446 (O_446,N_2886,N_2875);
and UO_447 (O_447,N_2968,N_2990);
nor UO_448 (O_448,N_2970,N_2888);
nor UO_449 (O_449,N_2809,N_2908);
and UO_450 (O_450,N_2868,N_2921);
nand UO_451 (O_451,N_2853,N_2925);
or UO_452 (O_452,N_2930,N_2876);
or UO_453 (O_453,N_2973,N_2906);
nand UO_454 (O_454,N_2887,N_2961);
nand UO_455 (O_455,N_2865,N_2875);
and UO_456 (O_456,N_2975,N_2836);
nand UO_457 (O_457,N_2903,N_2982);
nand UO_458 (O_458,N_2865,N_2822);
and UO_459 (O_459,N_2847,N_2952);
nor UO_460 (O_460,N_2959,N_2853);
nand UO_461 (O_461,N_2802,N_2881);
and UO_462 (O_462,N_2885,N_2938);
nor UO_463 (O_463,N_2903,N_2962);
and UO_464 (O_464,N_2845,N_2895);
nor UO_465 (O_465,N_2948,N_2931);
nand UO_466 (O_466,N_2936,N_2848);
and UO_467 (O_467,N_2986,N_2927);
or UO_468 (O_468,N_2838,N_2860);
nor UO_469 (O_469,N_2837,N_2816);
or UO_470 (O_470,N_2808,N_2879);
nand UO_471 (O_471,N_2971,N_2828);
or UO_472 (O_472,N_2801,N_2808);
nor UO_473 (O_473,N_2833,N_2896);
and UO_474 (O_474,N_2957,N_2821);
nor UO_475 (O_475,N_2878,N_2851);
and UO_476 (O_476,N_2983,N_2841);
and UO_477 (O_477,N_2802,N_2979);
nand UO_478 (O_478,N_2981,N_2986);
and UO_479 (O_479,N_2865,N_2942);
and UO_480 (O_480,N_2891,N_2840);
nand UO_481 (O_481,N_2827,N_2874);
and UO_482 (O_482,N_2903,N_2800);
nand UO_483 (O_483,N_2871,N_2927);
and UO_484 (O_484,N_2999,N_2889);
or UO_485 (O_485,N_2822,N_2963);
or UO_486 (O_486,N_2841,N_2925);
or UO_487 (O_487,N_2932,N_2850);
or UO_488 (O_488,N_2962,N_2899);
or UO_489 (O_489,N_2811,N_2853);
or UO_490 (O_490,N_2827,N_2877);
nor UO_491 (O_491,N_2804,N_2979);
nand UO_492 (O_492,N_2812,N_2990);
or UO_493 (O_493,N_2913,N_2979);
or UO_494 (O_494,N_2962,N_2881);
nor UO_495 (O_495,N_2964,N_2804);
and UO_496 (O_496,N_2972,N_2880);
nor UO_497 (O_497,N_2894,N_2896);
and UO_498 (O_498,N_2840,N_2958);
and UO_499 (O_499,N_2980,N_2865);
endmodule