module basic_500_3000_500_4_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_133,In_146);
or U1 (N_1,In_391,In_167);
nand U2 (N_2,In_305,In_462);
xor U3 (N_3,In_404,In_3);
nand U4 (N_4,In_148,In_439);
or U5 (N_5,In_378,In_414);
and U6 (N_6,In_301,In_231);
xnor U7 (N_7,In_111,In_260);
nand U8 (N_8,In_356,In_43);
and U9 (N_9,In_273,In_358);
and U10 (N_10,In_71,In_7);
or U11 (N_11,In_15,In_251);
nor U12 (N_12,In_426,In_469);
and U13 (N_13,In_11,In_61);
nand U14 (N_14,In_152,In_267);
and U15 (N_15,In_178,In_31);
nor U16 (N_16,In_52,In_198);
and U17 (N_17,In_176,In_406);
or U18 (N_18,In_286,In_241);
or U19 (N_19,In_367,In_242);
or U20 (N_20,In_27,In_486);
or U21 (N_21,In_172,In_475);
xnor U22 (N_22,In_262,In_185);
or U23 (N_23,In_177,In_62);
or U24 (N_24,In_168,In_42);
nand U25 (N_25,In_6,In_73);
and U26 (N_26,In_104,In_129);
and U27 (N_27,In_332,In_463);
nor U28 (N_28,In_153,In_25);
nor U29 (N_29,In_481,In_65);
and U30 (N_30,In_388,In_109);
nor U31 (N_31,In_54,In_105);
nand U32 (N_32,In_280,In_409);
and U33 (N_33,In_239,In_100);
nand U34 (N_34,In_429,In_490);
xor U35 (N_35,In_103,In_413);
nor U36 (N_36,In_284,In_106);
and U37 (N_37,In_383,In_59);
and U38 (N_38,In_304,In_44);
xnor U39 (N_39,In_214,In_279);
xnor U40 (N_40,In_194,In_86);
nor U41 (N_41,In_425,In_182);
nand U42 (N_42,In_88,In_67);
and U43 (N_43,In_10,In_116);
or U44 (N_44,In_16,In_258);
or U45 (N_45,In_164,In_226);
and U46 (N_46,In_477,In_157);
and U47 (N_47,In_181,In_322);
nor U48 (N_48,In_2,In_76);
and U49 (N_49,In_47,In_115);
nand U50 (N_50,In_455,In_63);
or U51 (N_51,In_319,In_366);
and U52 (N_52,In_89,In_350);
and U53 (N_53,In_126,In_271);
nand U54 (N_54,In_252,In_184);
and U55 (N_55,In_277,In_438);
or U56 (N_56,In_220,In_158);
or U57 (N_57,In_345,In_134);
or U58 (N_58,In_99,In_308);
and U59 (N_59,In_323,In_432);
nor U60 (N_60,In_493,In_142);
and U61 (N_61,In_349,In_183);
or U62 (N_62,In_472,In_238);
nand U63 (N_63,In_246,In_180);
nand U64 (N_64,In_447,In_492);
nand U65 (N_65,In_56,In_163);
nor U66 (N_66,In_327,In_21);
xor U67 (N_67,In_313,In_204);
or U68 (N_68,In_140,In_309);
and U69 (N_69,In_36,In_57);
nor U70 (N_70,In_297,In_84);
xor U71 (N_71,In_159,In_17);
or U72 (N_72,In_113,In_147);
or U73 (N_73,In_41,In_173);
nand U74 (N_74,In_371,In_321);
or U75 (N_75,In_179,In_390);
nand U76 (N_76,In_411,In_424);
xnor U77 (N_77,In_131,In_22);
xnor U78 (N_78,In_275,In_225);
or U79 (N_79,In_255,In_200);
nor U80 (N_80,In_249,In_488);
and U81 (N_81,In_289,In_49);
or U82 (N_82,In_110,In_368);
xnor U83 (N_83,In_64,In_376);
nand U84 (N_84,In_456,In_94);
and U85 (N_85,In_34,In_5);
nand U86 (N_86,In_274,In_46);
or U87 (N_87,In_58,In_160);
and U88 (N_88,In_174,In_290);
or U89 (N_89,In_359,In_81);
nand U90 (N_90,In_276,In_235);
nor U91 (N_91,In_269,In_278);
nand U92 (N_92,In_195,In_29);
nor U93 (N_93,In_418,In_362);
nand U94 (N_94,In_26,In_270);
and U95 (N_95,In_398,In_282);
nand U96 (N_96,In_8,In_123);
nor U97 (N_97,In_303,In_407);
nor U98 (N_98,In_395,In_449);
and U99 (N_99,In_292,In_487);
or U100 (N_100,In_291,In_340);
or U101 (N_101,In_234,In_468);
nand U102 (N_102,In_119,In_82);
or U103 (N_103,In_364,In_474);
or U104 (N_104,In_320,In_460);
nor U105 (N_105,In_445,In_387);
and U106 (N_106,In_216,In_93);
or U107 (N_107,In_466,In_85);
or U108 (N_108,In_192,In_318);
and U109 (N_109,In_221,In_331);
xnor U110 (N_110,In_248,In_431);
xnor U111 (N_111,In_373,In_312);
xor U112 (N_112,In_259,In_441);
and U113 (N_113,In_66,In_35);
nand U114 (N_114,In_434,In_50);
and U115 (N_115,In_324,In_410);
or U116 (N_116,In_154,In_202);
nor U117 (N_117,In_298,In_268);
nor U118 (N_118,In_346,In_296);
nand U119 (N_119,In_243,In_55);
and U120 (N_120,In_400,In_405);
and U121 (N_121,In_219,In_263);
and U122 (N_122,In_139,In_394);
and U123 (N_123,In_28,In_496);
and U124 (N_124,In_333,In_471);
and U125 (N_125,In_162,In_156);
nor U126 (N_126,In_402,In_326);
nor U127 (N_127,In_261,In_385);
nand U128 (N_128,In_87,In_299);
nand U129 (N_129,In_347,In_440);
or U130 (N_130,In_92,In_215);
nand U131 (N_131,In_257,In_452);
or U132 (N_132,In_265,In_196);
and U133 (N_133,In_75,In_232);
nand U134 (N_134,In_342,In_121);
nor U135 (N_135,In_341,In_130);
nand U136 (N_136,In_302,In_69);
nor U137 (N_137,In_428,In_498);
and U138 (N_138,In_166,In_485);
nand U139 (N_139,In_461,In_442);
and U140 (N_140,In_101,In_499);
nor U141 (N_141,In_91,In_392);
or U142 (N_142,In_209,In_375);
nor U143 (N_143,In_1,In_132);
nand U144 (N_144,In_479,In_287);
nand U145 (N_145,In_408,In_430);
and U146 (N_146,In_495,In_14);
nor U147 (N_147,In_13,In_169);
or U148 (N_148,In_186,In_476);
nor U149 (N_149,In_328,In_144);
nor U150 (N_150,In_337,In_236);
xor U151 (N_151,In_12,In_427);
nor U152 (N_152,In_330,In_199);
nand U153 (N_153,In_306,In_165);
and U154 (N_154,In_372,In_229);
or U155 (N_155,In_230,In_416);
nor U156 (N_156,In_124,In_102);
and U157 (N_157,In_83,In_206);
nor U158 (N_158,In_141,In_228);
or U159 (N_159,In_150,In_191);
nand U160 (N_160,In_51,In_369);
nor U161 (N_161,In_421,In_448);
or U162 (N_162,In_70,In_77);
or U163 (N_163,In_40,In_117);
xnor U164 (N_164,In_253,In_415);
nand U165 (N_165,In_193,In_227);
nor U166 (N_166,In_454,In_108);
xnor U167 (N_167,In_363,In_125);
nor U168 (N_168,In_213,In_365);
and U169 (N_169,In_171,In_38);
nand U170 (N_170,In_444,In_112);
or U171 (N_171,In_436,In_33);
and U172 (N_172,In_128,In_433);
nand U173 (N_173,In_233,In_453);
nand U174 (N_174,In_329,In_310);
nor U175 (N_175,In_201,In_355);
nor U176 (N_176,In_380,In_491);
nor U177 (N_177,In_325,In_457);
nor U178 (N_178,In_357,In_4);
xor U179 (N_179,In_352,In_18);
nor U180 (N_180,In_207,In_19);
nand U181 (N_181,In_212,In_294);
and U182 (N_182,In_422,In_339);
nand U183 (N_183,In_283,In_118);
xor U184 (N_184,In_343,In_211);
nor U185 (N_185,In_272,In_403);
nand U186 (N_186,In_161,In_264);
nor U187 (N_187,In_107,In_483);
nand U188 (N_188,In_353,In_437);
or U189 (N_189,In_23,In_203);
or U190 (N_190,In_401,In_417);
nand U191 (N_191,In_467,In_90);
or U192 (N_192,In_300,In_247);
nand U193 (N_193,In_237,In_489);
nand U194 (N_194,In_240,In_170);
and U195 (N_195,In_32,In_217);
nor U196 (N_196,In_374,In_381);
and U197 (N_197,In_143,In_480);
and U198 (N_198,In_149,In_151);
nand U199 (N_199,In_311,In_79);
and U200 (N_200,In_458,In_338);
and U201 (N_201,In_208,In_473);
nor U202 (N_202,In_497,In_443);
nor U203 (N_203,In_396,In_335);
or U204 (N_204,In_354,In_95);
nor U205 (N_205,In_389,In_254);
nand U206 (N_206,In_188,In_114);
nand U207 (N_207,In_397,In_24);
nor U208 (N_208,In_360,In_37);
xor U209 (N_209,In_446,In_478);
and U210 (N_210,In_465,In_293);
nor U211 (N_211,In_210,In_316);
xnor U212 (N_212,In_53,In_60);
nand U213 (N_213,In_399,In_9);
nand U214 (N_214,In_74,In_98);
nor U215 (N_215,In_30,In_245);
nor U216 (N_216,In_423,In_334);
or U217 (N_217,In_351,In_484);
nor U218 (N_218,In_175,In_379);
nand U219 (N_219,In_0,In_155);
xnor U220 (N_220,In_288,In_120);
or U221 (N_221,In_122,In_419);
or U222 (N_222,In_370,In_459);
and U223 (N_223,In_344,In_382);
xor U224 (N_224,In_223,In_224);
or U225 (N_225,In_138,In_295);
nand U226 (N_226,In_361,In_197);
xor U227 (N_227,In_68,In_464);
nor U228 (N_228,In_482,In_48);
nand U229 (N_229,In_145,In_78);
or U230 (N_230,In_20,In_451);
or U231 (N_231,In_189,In_187);
nor U232 (N_232,In_307,In_494);
nor U233 (N_233,In_205,In_412);
xnor U234 (N_234,In_450,In_470);
nor U235 (N_235,In_97,In_281);
and U236 (N_236,In_96,In_222);
nand U237 (N_237,In_285,In_250);
and U238 (N_238,In_336,In_420);
nor U239 (N_239,In_45,In_39);
or U240 (N_240,In_266,In_386);
or U241 (N_241,In_127,In_377);
nand U242 (N_242,In_256,In_135);
and U243 (N_243,In_314,In_80);
nor U244 (N_244,In_137,In_244);
and U245 (N_245,In_435,In_317);
nand U246 (N_246,In_384,In_393);
or U247 (N_247,In_218,In_348);
nor U248 (N_248,In_136,In_72);
nor U249 (N_249,In_315,In_190);
nor U250 (N_250,In_268,In_302);
nor U251 (N_251,In_274,In_32);
nor U252 (N_252,In_464,In_189);
xor U253 (N_253,In_92,In_341);
nor U254 (N_254,In_481,In_391);
and U255 (N_255,In_297,In_92);
nor U256 (N_256,In_74,In_51);
nor U257 (N_257,In_114,In_33);
or U258 (N_258,In_93,In_14);
or U259 (N_259,In_276,In_44);
and U260 (N_260,In_301,In_354);
and U261 (N_261,In_96,In_206);
and U262 (N_262,In_492,In_380);
nand U263 (N_263,In_356,In_260);
nand U264 (N_264,In_137,In_494);
nand U265 (N_265,In_241,In_294);
nand U266 (N_266,In_218,In_363);
nor U267 (N_267,In_410,In_221);
and U268 (N_268,In_433,In_410);
or U269 (N_269,In_422,In_328);
nor U270 (N_270,In_63,In_387);
nor U271 (N_271,In_116,In_318);
nand U272 (N_272,In_281,In_409);
and U273 (N_273,In_351,In_387);
nand U274 (N_274,In_24,In_435);
nor U275 (N_275,In_391,In_340);
xor U276 (N_276,In_302,In_200);
and U277 (N_277,In_193,In_206);
and U278 (N_278,In_469,In_11);
nand U279 (N_279,In_218,In_320);
nand U280 (N_280,In_18,In_300);
nor U281 (N_281,In_397,In_371);
xnor U282 (N_282,In_456,In_141);
nor U283 (N_283,In_129,In_480);
xor U284 (N_284,In_44,In_446);
or U285 (N_285,In_225,In_329);
nand U286 (N_286,In_103,In_440);
or U287 (N_287,In_369,In_194);
and U288 (N_288,In_97,In_335);
xor U289 (N_289,In_404,In_276);
nand U290 (N_290,In_498,In_350);
and U291 (N_291,In_50,In_402);
and U292 (N_292,In_343,In_288);
xnor U293 (N_293,In_263,In_283);
or U294 (N_294,In_306,In_352);
xnor U295 (N_295,In_226,In_309);
nor U296 (N_296,In_56,In_371);
nor U297 (N_297,In_254,In_24);
and U298 (N_298,In_255,In_475);
nand U299 (N_299,In_419,In_322);
xnor U300 (N_300,In_231,In_173);
nor U301 (N_301,In_234,In_445);
nand U302 (N_302,In_91,In_129);
or U303 (N_303,In_335,In_460);
or U304 (N_304,In_48,In_443);
or U305 (N_305,In_115,In_331);
and U306 (N_306,In_368,In_488);
or U307 (N_307,In_119,In_35);
nor U308 (N_308,In_297,In_10);
xor U309 (N_309,In_440,In_408);
or U310 (N_310,In_182,In_480);
nand U311 (N_311,In_461,In_462);
xnor U312 (N_312,In_103,In_374);
nand U313 (N_313,In_135,In_344);
and U314 (N_314,In_213,In_392);
and U315 (N_315,In_383,In_322);
or U316 (N_316,In_170,In_374);
nand U317 (N_317,In_261,In_3);
nor U318 (N_318,In_320,In_377);
nor U319 (N_319,In_245,In_266);
nand U320 (N_320,In_22,In_316);
or U321 (N_321,In_39,In_286);
xnor U322 (N_322,In_165,In_249);
and U323 (N_323,In_325,In_149);
or U324 (N_324,In_242,In_64);
nor U325 (N_325,In_75,In_81);
nor U326 (N_326,In_140,In_499);
and U327 (N_327,In_287,In_443);
nor U328 (N_328,In_230,In_349);
nand U329 (N_329,In_295,In_211);
and U330 (N_330,In_307,In_474);
and U331 (N_331,In_131,In_264);
nor U332 (N_332,In_292,In_326);
or U333 (N_333,In_359,In_462);
nor U334 (N_334,In_347,In_30);
and U335 (N_335,In_369,In_69);
nor U336 (N_336,In_407,In_231);
nor U337 (N_337,In_189,In_287);
nand U338 (N_338,In_162,In_228);
nand U339 (N_339,In_459,In_134);
nand U340 (N_340,In_91,In_383);
xnor U341 (N_341,In_249,In_368);
nor U342 (N_342,In_368,In_50);
and U343 (N_343,In_447,In_127);
nor U344 (N_344,In_487,In_289);
xnor U345 (N_345,In_147,In_86);
and U346 (N_346,In_276,In_185);
nand U347 (N_347,In_271,In_88);
and U348 (N_348,In_1,In_364);
xor U349 (N_349,In_224,In_394);
or U350 (N_350,In_33,In_118);
and U351 (N_351,In_356,In_169);
nand U352 (N_352,In_328,In_86);
nand U353 (N_353,In_16,In_218);
or U354 (N_354,In_40,In_13);
or U355 (N_355,In_68,In_35);
nor U356 (N_356,In_163,In_387);
nand U357 (N_357,In_440,In_349);
and U358 (N_358,In_266,In_362);
and U359 (N_359,In_343,In_230);
nand U360 (N_360,In_129,In_26);
nor U361 (N_361,In_79,In_229);
and U362 (N_362,In_178,In_431);
and U363 (N_363,In_286,In_270);
or U364 (N_364,In_84,In_366);
and U365 (N_365,In_25,In_397);
nor U366 (N_366,In_209,In_373);
nand U367 (N_367,In_217,In_155);
or U368 (N_368,In_10,In_416);
nand U369 (N_369,In_380,In_263);
or U370 (N_370,In_184,In_84);
and U371 (N_371,In_216,In_225);
or U372 (N_372,In_368,In_181);
nand U373 (N_373,In_258,In_346);
and U374 (N_374,In_1,In_312);
and U375 (N_375,In_425,In_157);
or U376 (N_376,In_230,In_293);
nand U377 (N_377,In_428,In_239);
and U378 (N_378,In_207,In_307);
nand U379 (N_379,In_101,In_345);
or U380 (N_380,In_207,In_454);
nor U381 (N_381,In_483,In_492);
nand U382 (N_382,In_61,In_2);
or U383 (N_383,In_153,In_263);
nand U384 (N_384,In_140,In_458);
nand U385 (N_385,In_107,In_10);
or U386 (N_386,In_338,In_497);
nor U387 (N_387,In_167,In_438);
nor U388 (N_388,In_407,In_388);
and U389 (N_389,In_382,In_200);
nor U390 (N_390,In_28,In_116);
or U391 (N_391,In_378,In_75);
nand U392 (N_392,In_131,In_102);
nand U393 (N_393,In_141,In_166);
or U394 (N_394,In_114,In_35);
nor U395 (N_395,In_79,In_213);
nor U396 (N_396,In_177,In_361);
nor U397 (N_397,In_457,In_64);
nor U398 (N_398,In_254,In_425);
and U399 (N_399,In_206,In_282);
or U400 (N_400,In_426,In_365);
nor U401 (N_401,In_60,In_56);
and U402 (N_402,In_73,In_495);
and U403 (N_403,In_332,In_5);
and U404 (N_404,In_97,In_424);
nor U405 (N_405,In_359,In_167);
nor U406 (N_406,In_183,In_173);
nand U407 (N_407,In_139,In_161);
nand U408 (N_408,In_212,In_155);
xnor U409 (N_409,In_218,In_195);
nand U410 (N_410,In_317,In_456);
nand U411 (N_411,In_106,In_463);
nand U412 (N_412,In_21,In_110);
nor U413 (N_413,In_91,In_107);
nor U414 (N_414,In_370,In_3);
nand U415 (N_415,In_194,In_47);
or U416 (N_416,In_4,In_249);
xnor U417 (N_417,In_204,In_134);
and U418 (N_418,In_255,In_52);
nand U419 (N_419,In_269,In_344);
nand U420 (N_420,In_114,In_18);
nor U421 (N_421,In_253,In_18);
or U422 (N_422,In_486,In_68);
nand U423 (N_423,In_246,In_87);
nor U424 (N_424,In_367,In_21);
and U425 (N_425,In_215,In_52);
nor U426 (N_426,In_29,In_147);
xnor U427 (N_427,In_142,In_140);
and U428 (N_428,In_384,In_178);
and U429 (N_429,In_56,In_292);
and U430 (N_430,In_284,In_25);
nand U431 (N_431,In_429,In_228);
or U432 (N_432,In_28,In_227);
or U433 (N_433,In_170,In_421);
or U434 (N_434,In_484,In_275);
nand U435 (N_435,In_184,In_34);
nand U436 (N_436,In_417,In_356);
xor U437 (N_437,In_240,In_10);
and U438 (N_438,In_356,In_484);
or U439 (N_439,In_208,In_153);
nor U440 (N_440,In_50,In_414);
nor U441 (N_441,In_224,In_471);
and U442 (N_442,In_416,In_162);
nor U443 (N_443,In_412,In_91);
nand U444 (N_444,In_53,In_364);
nor U445 (N_445,In_347,In_375);
nand U446 (N_446,In_338,In_405);
nand U447 (N_447,In_111,In_197);
nor U448 (N_448,In_191,In_455);
or U449 (N_449,In_316,In_26);
nor U450 (N_450,In_322,In_298);
or U451 (N_451,In_11,In_231);
nor U452 (N_452,In_315,In_157);
or U453 (N_453,In_273,In_217);
or U454 (N_454,In_23,In_15);
and U455 (N_455,In_99,In_319);
and U456 (N_456,In_193,In_172);
nor U457 (N_457,In_379,In_470);
or U458 (N_458,In_176,In_205);
or U459 (N_459,In_409,In_28);
and U460 (N_460,In_276,In_129);
xnor U461 (N_461,In_324,In_289);
and U462 (N_462,In_498,In_446);
and U463 (N_463,In_89,In_367);
or U464 (N_464,In_98,In_202);
or U465 (N_465,In_203,In_221);
nand U466 (N_466,In_343,In_232);
xnor U467 (N_467,In_467,In_256);
xor U468 (N_468,In_140,In_64);
nand U469 (N_469,In_110,In_345);
or U470 (N_470,In_190,In_434);
or U471 (N_471,In_415,In_64);
or U472 (N_472,In_173,In_475);
nor U473 (N_473,In_133,In_366);
xor U474 (N_474,In_275,In_316);
nor U475 (N_475,In_2,In_472);
nand U476 (N_476,In_122,In_207);
or U477 (N_477,In_346,In_180);
and U478 (N_478,In_443,In_178);
nor U479 (N_479,In_36,In_44);
and U480 (N_480,In_244,In_192);
and U481 (N_481,In_291,In_99);
and U482 (N_482,In_414,In_490);
and U483 (N_483,In_499,In_114);
nor U484 (N_484,In_90,In_300);
and U485 (N_485,In_108,In_399);
and U486 (N_486,In_267,In_483);
or U487 (N_487,In_164,In_318);
or U488 (N_488,In_340,In_463);
and U489 (N_489,In_60,In_440);
and U490 (N_490,In_78,In_129);
nor U491 (N_491,In_416,In_293);
nand U492 (N_492,In_116,In_9);
nor U493 (N_493,In_331,In_96);
nor U494 (N_494,In_365,In_437);
nor U495 (N_495,In_266,In_220);
nand U496 (N_496,In_364,In_489);
or U497 (N_497,In_399,In_0);
and U498 (N_498,In_344,In_442);
xnor U499 (N_499,In_270,In_334);
or U500 (N_500,In_416,In_40);
nand U501 (N_501,In_213,In_59);
nand U502 (N_502,In_83,In_22);
or U503 (N_503,In_428,In_79);
and U504 (N_504,In_367,In_40);
and U505 (N_505,In_376,In_235);
and U506 (N_506,In_309,In_365);
xor U507 (N_507,In_79,In_202);
or U508 (N_508,In_43,In_485);
nor U509 (N_509,In_438,In_443);
nand U510 (N_510,In_272,In_62);
nand U511 (N_511,In_398,In_325);
nand U512 (N_512,In_18,In_14);
and U513 (N_513,In_130,In_274);
or U514 (N_514,In_65,In_123);
nor U515 (N_515,In_329,In_176);
nor U516 (N_516,In_184,In_388);
nand U517 (N_517,In_199,In_459);
nand U518 (N_518,In_196,In_334);
nor U519 (N_519,In_247,In_458);
or U520 (N_520,In_215,In_151);
nand U521 (N_521,In_84,In_167);
xnor U522 (N_522,In_68,In_381);
nand U523 (N_523,In_259,In_90);
or U524 (N_524,In_410,In_137);
and U525 (N_525,In_418,In_62);
nand U526 (N_526,In_438,In_414);
or U527 (N_527,In_116,In_319);
nor U528 (N_528,In_31,In_169);
nor U529 (N_529,In_120,In_275);
xor U530 (N_530,In_5,In_45);
or U531 (N_531,In_461,In_492);
nor U532 (N_532,In_70,In_12);
nor U533 (N_533,In_23,In_176);
nand U534 (N_534,In_148,In_493);
or U535 (N_535,In_199,In_487);
and U536 (N_536,In_123,In_20);
nand U537 (N_537,In_15,In_201);
nor U538 (N_538,In_282,In_454);
or U539 (N_539,In_123,In_467);
xor U540 (N_540,In_232,In_234);
nand U541 (N_541,In_233,In_451);
nand U542 (N_542,In_58,In_6);
nand U543 (N_543,In_95,In_40);
and U544 (N_544,In_353,In_55);
nor U545 (N_545,In_152,In_66);
or U546 (N_546,In_148,In_402);
or U547 (N_547,In_196,In_437);
or U548 (N_548,In_348,In_43);
nand U549 (N_549,In_467,In_275);
nor U550 (N_550,In_462,In_365);
xor U551 (N_551,In_88,In_243);
nor U552 (N_552,In_331,In_8);
and U553 (N_553,In_38,In_458);
nand U554 (N_554,In_30,In_65);
nand U555 (N_555,In_179,In_70);
or U556 (N_556,In_334,In_420);
and U557 (N_557,In_207,In_203);
and U558 (N_558,In_138,In_308);
nand U559 (N_559,In_353,In_400);
or U560 (N_560,In_32,In_387);
xnor U561 (N_561,In_15,In_402);
and U562 (N_562,In_348,In_372);
nor U563 (N_563,In_400,In_231);
nand U564 (N_564,In_478,In_433);
or U565 (N_565,In_326,In_134);
xor U566 (N_566,In_196,In_220);
or U567 (N_567,In_96,In_265);
or U568 (N_568,In_409,In_414);
xnor U569 (N_569,In_101,In_378);
or U570 (N_570,In_210,In_240);
or U571 (N_571,In_370,In_396);
nand U572 (N_572,In_195,In_342);
and U573 (N_573,In_184,In_9);
nand U574 (N_574,In_254,In_75);
or U575 (N_575,In_198,In_498);
xnor U576 (N_576,In_288,In_31);
and U577 (N_577,In_480,In_201);
xnor U578 (N_578,In_455,In_293);
nor U579 (N_579,In_302,In_87);
or U580 (N_580,In_442,In_414);
nand U581 (N_581,In_478,In_320);
nor U582 (N_582,In_229,In_185);
and U583 (N_583,In_394,In_59);
nand U584 (N_584,In_486,In_340);
and U585 (N_585,In_481,In_274);
and U586 (N_586,In_411,In_451);
or U587 (N_587,In_379,In_413);
nand U588 (N_588,In_365,In_121);
or U589 (N_589,In_31,In_329);
or U590 (N_590,In_136,In_397);
or U591 (N_591,In_234,In_287);
nor U592 (N_592,In_48,In_143);
and U593 (N_593,In_288,In_375);
and U594 (N_594,In_296,In_281);
nand U595 (N_595,In_488,In_413);
and U596 (N_596,In_171,In_378);
and U597 (N_597,In_442,In_333);
nor U598 (N_598,In_478,In_189);
nor U599 (N_599,In_281,In_67);
nor U600 (N_600,In_344,In_498);
nor U601 (N_601,In_417,In_382);
and U602 (N_602,In_2,In_206);
nand U603 (N_603,In_36,In_429);
or U604 (N_604,In_218,In_204);
xnor U605 (N_605,In_387,In_306);
and U606 (N_606,In_257,In_339);
nand U607 (N_607,In_412,In_175);
or U608 (N_608,In_66,In_247);
nand U609 (N_609,In_13,In_217);
xnor U610 (N_610,In_418,In_387);
nor U611 (N_611,In_159,In_318);
or U612 (N_612,In_265,In_226);
nor U613 (N_613,In_112,In_181);
or U614 (N_614,In_50,In_365);
nor U615 (N_615,In_294,In_108);
or U616 (N_616,In_88,In_223);
and U617 (N_617,In_493,In_60);
and U618 (N_618,In_441,In_131);
nor U619 (N_619,In_464,In_35);
and U620 (N_620,In_54,In_341);
nand U621 (N_621,In_477,In_247);
nand U622 (N_622,In_322,In_15);
or U623 (N_623,In_75,In_344);
nand U624 (N_624,In_93,In_452);
nor U625 (N_625,In_62,In_98);
or U626 (N_626,In_452,In_285);
or U627 (N_627,In_208,In_166);
xnor U628 (N_628,In_118,In_158);
nand U629 (N_629,In_30,In_415);
nor U630 (N_630,In_92,In_482);
nand U631 (N_631,In_419,In_382);
and U632 (N_632,In_229,In_162);
and U633 (N_633,In_377,In_17);
or U634 (N_634,In_302,In_420);
or U635 (N_635,In_295,In_423);
xnor U636 (N_636,In_445,In_449);
nand U637 (N_637,In_171,In_259);
or U638 (N_638,In_393,In_409);
nand U639 (N_639,In_450,In_42);
or U640 (N_640,In_57,In_173);
xor U641 (N_641,In_315,In_177);
and U642 (N_642,In_417,In_89);
nor U643 (N_643,In_366,In_430);
nor U644 (N_644,In_328,In_456);
and U645 (N_645,In_401,In_265);
nand U646 (N_646,In_185,In_41);
nand U647 (N_647,In_239,In_202);
nor U648 (N_648,In_493,In_252);
and U649 (N_649,In_261,In_394);
nand U650 (N_650,In_159,In_475);
and U651 (N_651,In_457,In_296);
or U652 (N_652,In_261,In_94);
and U653 (N_653,In_333,In_252);
and U654 (N_654,In_287,In_382);
or U655 (N_655,In_33,In_373);
or U656 (N_656,In_374,In_218);
and U657 (N_657,In_7,In_151);
nor U658 (N_658,In_346,In_466);
nand U659 (N_659,In_73,In_164);
and U660 (N_660,In_351,In_111);
nand U661 (N_661,In_286,In_485);
xor U662 (N_662,In_115,In_285);
nor U663 (N_663,In_156,In_69);
or U664 (N_664,In_125,In_285);
or U665 (N_665,In_130,In_153);
xor U666 (N_666,In_43,In_235);
and U667 (N_667,In_460,In_11);
nor U668 (N_668,In_257,In_298);
xor U669 (N_669,In_341,In_226);
nor U670 (N_670,In_179,In_111);
or U671 (N_671,In_46,In_474);
and U672 (N_672,In_100,In_162);
and U673 (N_673,In_190,In_272);
nor U674 (N_674,In_170,In_107);
nor U675 (N_675,In_264,In_191);
xnor U676 (N_676,In_459,In_393);
and U677 (N_677,In_389,In_295);
nor U678 (N_678,In_239,In_480);
and U679 (N_679,In_23,In_464);
nor U680 (N_680,In_213,In_458);
nand U681 (N_681,In_20,In_444);
xor U682 (N_682,In_396,In_443);
nand U683 (N_683,In_8,In_172);
or U684 (N_684,In_232,In_123);
nand U685 (N_685,In_38,In_14);
nor U686 (N_686,In_110,In_317);
or U687 (N_687,In_72,In_46);
nor U688 (N_688,In_134,In_172);
xor U689 (N_689,In_230,In_34);
nand U690 (N_690,In_169,In_323);
and U691 (N_691,In_117,In_232);
nor U692 (N_692,In_44,In_338);
or U693 (N_693,In_324,In_62);
nor U694 (N_694,In_438,In_276);
nand U695 (N_695,In_443,In_402);
nand U696 (N_696,In_196,In_94);
or U697 (N_697,In_140,In_202);
and U698 (N_698,In_61,In_412);
nor U699 (N_699,In_273,In_223);
or U700 (N_700,In_492,In_399);
nor U701 (N_701,In_369,In_261);
or U702 (N_702,In_274,In_257);
and U703 (N_703,In_166,In_24);
xor U704 (N_704,In_267,In_373);
nor U705 (N_705,In_279,In_63);
or U706 (N_706,In_65,In_69);
nor U707 (N_707,In_126,In_239);
nand U708 (N_708,In_345,In_94);
or U709 (N_709,In_479,In_345);
xor U710 (N_710,In_19,In_38);
nand U711 (N_711,In_189,In_393);
nor U712 (N_712,In_130,In_6);
or U713 (N_713,In_108,In_102);
nand U714 (N_714,In_169,In_234);
nor U715 (N_715,In_289,In_166);
nor U716 (N_716,In_325,In_258);
xor U717 (N_717,In_34,In_47);
nand U718 (N_718,In_220,In_25);
and U719 (N_719,In_342,In_30);
nand U720 (N_720,In_75,In_464);
nor U721 (N_721,In_305,In_275);
xnor U722 (N_722,In_456,In_440);
and U723 (N_723,In_128,In_424);
xnor U724 (N_724,In_10,In_367);
nor U725 (N_725,In_15,In_6);
and U726 (N_726,In_193,In_129);
or U727 (N_727,In_10,In_496);
or U728 (N_728,In_424,In_306);
or U729 (N_729,In_490,In_90);
or U730 (N_730,In_197,In_39);
or U731 (N_731,In_57,In_275);
xnor U732 (N_732,In_350,In_239);
nand U733 (N_733,In_129,In_490);
nor U734 (N_734,In_238,In_468);
nor U735 (N_735,In_166,In_213);
nor U736 (N_736,In_325,In_383);
nor U737 (N_737,In_29,In_364);
nor U738 (N_738,In_157,In_164);
nor U739 (N_739,In_394,In_187);
and U740 (N_740,In_136,In_212);
xor U741 (N_741,In_82,In_115);
or U742 (N_742,In_27,In_143);
nand U743 (N_743,In_306,In_444);
or U744 (N_744,In_227,In_189);
or U745 (N_745,In_68,In_17);
nor U746 (N_746,In_402,In_41);
nand U747 (N_747,In_250,In_134);
and U748 (N_748,In_59,In_325);
and U749 (N_749,In_8,In_495);
or U750 (N_750,N_477,N_613);
xnor U751 (N_751,N_211,N_498);
or U752 (N_752,N_516,N_259);
and U753 (N_753,N_744,N_73);
or U754 (N_754,N_324,N_658);
and U755 (N_755,N_708,N_473);
or U756 (N_756,N_688,N_695);
and U757 (N_757,N_65,N_33);
nor U758 (N_758,N_86,N_639);
and U759 (N_759,N_712,N_574);
nor U760 (N_760,N_589,N_623);
nand U761 (N_761,N_145,N_631);
nor U762 (N_762,N_434,N_601);
xnor U763 (N_763,N_442,N_20);
nand U764 (N_764,N_437,N_647);
or U765 (N_765,N_611,N_171);
nor U766 (N_766,N_528,N_375);
nor U767 (N_767,N_285,N_167);
or U768 (N_768,N_3,N_519);
or U769 (N_769,N_316,N_311);
and U770 (N_770,N_597,N_274);
and U771 (N_771,N_263,N_487);
xor U772 (N_772,N_677,N_642);
nand U773 (N_773,N_42,N_691);
nor U774 (N_774,N_247,N_585);
or U775 (N_775,N_441,N_321);
or U776 (N_776,N_50,N_340);
or U777 (N_777,N_128,N_665);
or U778 (N_778,N_191,N_686);
nor U779 (N_779,N_29,N_55);
xor U780 (N_780,N_350,N_370);
nor U781 (N_781,N_135,N_2);
xnor U782 (N_782,N_439,N_233);
and U783 (N_783,N_396,N_231);
and U784 (N_784,N_275,N_619);
or U785 (N_785,N_666,N_300);
nand U786 (N_786,N_577,N_292);
or U787 (N_787,N_355,N_314);
nand U788 (N_788,N_440,N_12);
nor U789 (N_789,N_322,N_599);
and U790 (N_790,N_289,N_36);
and U791 (N_791,N_667,N_297);
and U792 (N_792,N_70,N_106);
nor U793 (N_793,N_312,N_409);
or U794 (N_794,N_572,N_200);
nand U795 (N_795,N_232,N_557);
nand U796 (N_796,N_150,N_172);
nand U797 (N_797,N_747,N_290);
and U798 (N_798,N_710,N_626);
and U799 (N_799,N_410,N_347);
nor U800 (N_800,N_715,N_124);
nand U801 (N_801,N_485,N_662);
nand U802 (N_802,N_672,N_122);
and U803 (N_803,N_668,N_532);
or U804 (N_804,N_0,N_587);
or U805 (N_805,N_117,N_227);
nand U806 (N_806,N_168,N_353);
nand U807 (N_807,N_371,N_652);
or U808 (N_808,N_146,N_228);
nand U809 (N_809,N_511,N_335);
nand U810 (N_810,N_35,N_278);
nor U811 (N_811,N_664,N_286);
and U812 (N_812,N_205,N_709);
nor U813 (N_813,N_418,N_236);
and U814 (N_814,N_305,N_447);
or U815 (N_815,N_663,N_749);
nor U816 (N_816,N_424,N_154);
and U817 (N_817,N_66,N_414);
nand U818 (N_818,N_451,N_25);
xnor U819 (N_819,N_184,N_326);
and U820 (N_820,N_4,N_593);
nand U821 (N_821,N_416,N_68);
and U822 (N_822,N_294,N_334);
and U823 (N_823,N_500,N_617);
nand U824 (N_824,N_563,N_746);
nor U825 (N_825,N_210,N_644);
nand U826 (N_826,N_108,N_295);
xnor U827 (N_827,N_185,N_384);
nand U828 (N_828,N_397,N_555);
nand U829 (N_829,N_320,N_576);
or U830 (N_830,N_8,N_507);
nand U831 (N_831,N_367,N_160);
or U832 (N_832,N_391,N_678);
or U833 (N_833,N_607,N_645);
or U834 (N_834,N_304,N_43);
and U835 (N_835,N_554,N_521);
or U836 (N_836,N_279,N_583);
xor U837 (N_837,N_85,N_685);
nand U838 (N_838,N_470,N_573);
and U839 (N_839,N_248,N_482);
or U840 (N_840,N_386,N_129);
nand U841 (N_841,N_579,N_338);
nand U842 (N_842,N_348,N_54);
nor U843 (N_843,N_635,N_229);
nand U844 (N_844,N_45,N_354);
or U845 (N_845,N_313,N_458);
or U846 (N_846,N_656,N_392);
or U847 (N_847,N_343,N_330);
nand U848 (N_848,N_430,N_540);
and U849 (N_849,N_121,N_132);
nand U850 (N_850,N_366,N_280);
or U851 (N_851,N_520,N_360);
xnor U852 (N_852,N_475,N_98);
nor U853 (N_853,N_649,N_147);
or U854 (N_854,N_69,N_468);
or U855 (N_855,N_249,N_49);
nand U856 (N_856,N_676,N_78);
and U857 (N_857,N_443,N_284);
or U858 (N_858,N_199,N_553);
nand U859 (N_859,N_632,N_131);
nor U860 (N_860,N_533,N_161);
and U861 (N_861,N_244,N_408);
nand U862 (N_862,N_515,N_17);
and U863 (N_863,N_163,N_454);
nor U864 (N_864,N_361,N_213);
nand U865 (N_865,N_499,N_389);
and U866 (N_866,N_88,N_153);
or U867 (N_867,N_245,N_183);
xor U868 (N_868,N_719,N_188);
xnor U869 (N_869,N_272,N_201);
nand U870 (N_870,N_738,N_522);
or U871 (N_871,N_552,N_735);
nor U872 (N_872,N_693,N_123);
nand U873 (N_873,N_365,N_143);
or U874 (N_874,N_92,N_568);
or U875 (N_875,N_125,N_219);
nor U876 (N_876,N_192,N_400);
nor U877 (N_877,N_683,N_653);
and U878 (N_878,N_378,N_701);
and U879 (N_879,N_637,N_264);
nand U880 (N_880,N_369,N_336);
xnor U881 (N_881,N_291,N_591);
and U882 (N_882,N_260,N_100);
and U883 (N_883,N_598,N_559);
nand U884 (N_884,N_425,N_620);
nor U885 (N_885,N_446,N_327);
and U886 (N_886,N_26,N_342);
xor U887 (N_887,N_716,N_699);
nor U888 (N_888,N_536,N_376);
and U889 (N_889,N_718,N_696);
nand U890 (N_890,N_256,N_159);
nor U891 (N_891,N_670,N_692);
or U892 (N_892,N_339,N_673);
and U893 (N_893,N_594,N_571);
or U894 (N_894,N_212,N_257);
or U895 (N_895,N_242,N_281);
nand U896 (N_896,N_195,N_243);
nor U897 (N_897,N_506,N_99);
nand U898 (N_898,N_208,N_303);
nor U899 (N_899,N_445,N_251);
nand U900 (N_900,N_372,N_234);
nand U901 (N_901,N_58,N_721);
or U902 (N_902,N_112,N_44);
xnor U903 (N_903,N_514,N_728);
and U904 (N_904,N_467,N_651);
and U905 (N_905,N_187,N_287);
or U906 (N_906,N_592,N_733);
and U907 (N_907,N_302,N_341);
nor U908 (N_908,N_93,N_64);
or U909 (N_909,N_116,N_407);
or U910 (N_910,N_429,N_346);
or U911 (N_911,N_282,N_262);
xor U912 (N_912,N_513,N_222);
xnor U913 (N_913,N_11,N_450);
nor U914 (N_914,N_155,N_241);
or U915 (N_915,N_398,N_5);
and U916 (N_916,N_464,N_406);
nor U917 (N_917,N_518,N_165);
nor U918 (N_918,N_13,N_615);
xnor U919 (N_919,N_586,N_89);
or U920 (N_920,N_215,N_255);
or U921 (N_921,N_436,N_83);
nand U922 (N_922,N_104,N_603);
nand U923 (N_923,N_469,N_741);
or U924 (N_924,N_81,N_551);
nor U925 (N_925,N_137,N_114);
xor U926 (N_926,N_486,N_307);
nor U927 (N_927,N_344,N_140);
nand U928 (N_928,N_399,N_456);
nand U929 (N_929,N_10,N_494);
nand U930 (N_930,N_731,N_660);
and U931 (N_931,N_734,N_197);
and U932 (N_932,N_748,N_95);
nand U933 (N_933,N_56,N_562);
nand U934 (N_934,N_684,N_462);
nand U935 (N_935,N_503,N_30);
and U936 (N_936,N_37,N_657);
nand U937 (N_937,N_61,N_564);
nand U938 (N_938,N_432,N_561);
nor U939 (N_939,N_411,N_534);
or U940 (N_940,N_180,N_537);
nand U941 (N_941,N_141,N_535);
and U942 (N_942,N_704,N_202);
or U943 (N_943,N_48,N_101);
nor U944 (N_944,N_722,N_523);
and U945 (N_945,N_390,N_214);
nor U946 (N_946,N_428,N_190);
nand U947 (N_947,N_707,N_359);
and U948 (N_948,N_169,N_438);
and U949 (N_949,N_727,N_266);
or U950 (N_950,N_345,N_46);
and U951 (N_951,N_674,N_84);
or U952 (N_952,N_459,N_633);
nand U953 (N_953,N_136,N_706);
nand U954 (N_954,N_182,N_526);
nand U955 (N_955,N_694,N_690);
nor U956 (N_956,N_230,N_541);
nor U957 (N_957,N_157,N_74);
or U958 (N_958,N_725,N_119);
xnor U959 (N_959,N_253,N_550);
and U960 (N_960,N_40,N_698);
nor U961 (N_961,N_318,N_618);
nand U962 (N_962,N_268,N_393);
nor U963 (N_963,N_655,N_596);
nand U964 (N_964,N_134,N_269);
and U965 (N_965,N_39,N_118);
nand U966 (N_966,N_648,N_224);
xor U967 (N_967,N_501,N_90);
or U968 (N_968,N_363,N_705);
and U969 (N_969,N_349,N_700);
and U970 (N_970,N_388,N_53);
or U971 (N_971,N_544,N_337);
nand U972 (N_972,N_736,N_567);
nor U973 (N_973,N_558,N_193);
or U974 (N_974,N_356,N_588);
nand U975 (N_975,N_493,N_745);
nand U976 (N_976,N_556,N_276);
or U977 (N_977,N_237,N_604);
nor U978 (N_978,N_298,N_614);
or U979 (N_979,N_174,N_570);
and U980 (N_980,N_130,N_608);
nor U981 (N_981,N_332,N_270);
nor U982 (N_982,N_600,N_273);
nor U983 (N_983,N_629,N_739);
or U984 (N_984,N_524,N_323);
nor U985 (N_985,N_301,N_252);
and U986 (N_986,N_109,N_480);
xor U987 (N_987,N_527,N_622);
nand U988 (N_988,N_385,N_463);
nand U989 (N_989,N_82,N_415);
nand U990 (N_990,N_394,N_283);
nor U991 (N_991,N_457,N_606);
or U992 (N_992,N_203,N_403);
or U993 (N_993,N_206,N_261);
xor U994 (N_994,N_401,N_640);
and U995 (N_995,N_479,N_226);
and U996 (N_996,N_510,N_723);
nand U997 (N_997,N_584,N_529);
and U998 (N_998,N_546,N_650);
nand U999 (N_999,N_246,N_357);
nand U1000 (N_1000,N_60,N_669);
nor U1001 (N_1001,N_94,N_115);
nor U1002 (N_1002,N_627,N_308);
nand U1003 (N_1003,N_221,N_198);
nor U1004 (N_1004,N_138,N_460);
nand U1005 (N_1005,N_542,N_328);
nor U1006 (N_1006,N_176,N_713);
nor U1007 (N_1007,N_235,N_702);
nor U1008 (N_1008,N_51,N_413);
xnor U1009 (N_1009,N_654,N_164);
or U1010 (N_1010,N_267,N_15);
xor U1011 (N_1011,N_508,N_489);
or U1012 (N_1012,N_382,N_448);
and U1013 (N_1013,N_580,N_126);
nor U1014 (N_1014,N_638,N_525);
and U1015 (N_1015,N_220,N_315);
nand U1016 (N_1016,N_681,N_502);
xnor U1017 (N_1017,N_680,N_720);
xnor U1018 (N_1018,N_545,N_310);
nand U1019 (N_1019,N_148,N_377);
nor U1020 (N_1020,N_111,N_703);
nor U1021 (N_1021,N_582,N_52);
or U1022 (N_1022,N_31,N_530);
nand U1023 (N_1023,N_481,N_196);
xor U1024 (N_1024,N_621,N_417);
xnor U1025 (N_1025,N_250,N_110);
nand U1026 (N_1026,N_387,N_364);
xor U1027 (N_1027,N_726,N_488);
nand U1028 (N_1028,N_509,N_333);
nor U1029 (N_1029,N_299,N_277);
nand U1030 (N_1030,N_331,N_306);
nor U1031 (N_1031,N_610,N_549);
or U1032 (N_1032,N_62,N_402);
and U1033 (N_1033,N_547,N_566);
xnor U1034 (N_1034,N_609,N_543);
nor U1035 (N_1035,N_697,N_223);
and U1036 (N_1036,N_379,N_194);
and U1037 (N_1037,N_151,N_724);
nand U1038 (N_1038,N_166,N_158);
and U1039 (N_1039,N_9,N_675);
nand U1040 (N_1040,N_170,N_218);
nand U1041 (N_1041,N_127,N_431);
nand U1042 (N_1042,N_21,N_512);
or U1043 (N_1043,N_87,N_373);
or U1044 (N_1044,N_740,N_24);
or U1045 (N_1045,N_156,N_216);
nor U1046 (N_1046,N_538,N_565);
nor U1047 (N_1047,N_139,N_368);
or U1048 (N_1048,N_453,N_317);
nor U1049 (N_1049,N_6,N_319);
nand U1050 (N_1050,N_465,N_293);
nand U1051 (N_1051,N_149,N_22);
and U1052 (N_1052,N_7,N_497);
nor U1053 (N_1053,N_496,N_420);
nor U1054 (N_1054,N_76,N_225);
xor U1055 (N_1055,N_217,N_362);
nand U1056 (N_1056,N_605,N_419);
nor U1057 (N_1057,N_177,N_144);
nand U1058 (N_1058,N_57,N_186);
or U1059 (N_1059,N_423,N_67);
nand U1060 (N_1060,N_483,N_309);
and U1061 (N_1061,N_484,N_258);
nor U1062 (N_1062,N_120,N_581);
or U1063 (N_1063,N_133,N_113);
nor U1064 (N_1064,N_102,N_271);
nor U1065 (N_1065,N_27,N_91);
nand U1066 (N_1066,N_444,N_422);
nor U1067 (N_1067,N_624,N_238);
and U1068 (N_1068,N_351,N_449);
and U1069 (N_1069,N_630,N_472);
and U1070 (N_1070,N_28,N_296);
and U1071 (N_1071,N_178,N_732);
nor U1072 (N_1072,N_19,N_661);
nor U1073 (N_1073,N_602,N_152);
nand U1074 (N_1074,N_175,N_679);
nand U1075 (N_1075,N_590,N_717);
nand U1076 (N_1076,N_517,N_1);
nor U1077 (N_1077,N_730,N_358);
nor U1078 (N_1078,N_59,N_671);
nand U1079 (N_1079,N_288,N_471);
and U1080 (N_1080,N_103,N_531);
or U1081 (N_1081,N_23,N_492);
and U1082 (N_1082,N_569,N_41);
or U1083 (N_1083,N_239,N_714);
and U1084 (N_1084,N_173,N_404);
nand U1085 (N_1085,N_505,N_265);
nor U1086 (N_1086,N_325,N_162);
xnor U1087 (N_1087,N_179,N_374);
nor U1088 (N_1088,N_16,N_381);
nand U1089 (N_1089,N_14,N_466);
nor U1090 (N_1090,N_38,N_737);
and U1091 (N_1091,N_107,N_742);
xnor U1092 (N_1092,N_18,N_474);
nor U1093 (N_1093,N_491,N_504);
nand U1094 (N_1094,N_539,N_75);
or U1095 (N_1095,N_80,N_412);
and U1096 (N_1096,N_461,N_405);
or U1097 (N_1097,N_455,N_142);
and U1098 (N_1098,N_352,N_421);
nor U1099 (N_1099,N_96,N_77);
xor U1100 (N_1100,N_641,N_433);
nor U1101 (N_1101,N_476,N_435);
or U1102 (N_1102,N_72,N_204);
or U1103 (N_1103,N_490,N_63);
or U1104 (N_1104,N_729,N_79);
nor U1105 (N_1105,N_47,N_105);
or U1106 (N_1106,N_578,N_34);
nor U1107 (N_1107,N_612,N_616);
xor U1108 (N_1108,N_575,N_383);
nand U1109 (N_1109,N_478,N_634);
nor U1110 (N_1110,N_687,N_71);
or U1111 (N_1111,N_209,N_659);
or U1112 (N_1112,N_395,N_595);
and U1113 (N_1113,N_682,N_560);
nand U1114 (N_1114,N_380,N_689);
and U1115 (N_1115,N_711,N_426);
nand U1116 (N_1116,N_181,N_427);
nor U1117 (N_1117,N_743,N_240);
and U1118 (N_1118,N_329,N_207);
nor U1119 (N_1119,N_452,N_646);
and U1120 (N_1120,N_495,N_97);
or U1121 (N_1121,N_32,N_189);
and U1122 (N_1122,N_625,N_643);
nand U1123 (N_1123,N_636,N_548);
and U1124 (N_1124,N_254,N_628);
and U1125 (N_1125,N_699,N_379);
or U1126 (N_1126,N_568,N_346);
nor U1127 (N_1127,N_708,N_184);
or U1128 (N_1128,N_749,N_556);
nand U1129 (N_1129,N_551,N_526);
and U1130 (N_1130,N_53,N_532);
nand U1131 (N_1131,N_107,N_628);
nand U1132 (N_1132,N_665,N_629);
and U1133 (N_1133,N_540,N_695);
nor U1134 (N_1134,N_78,N_405);
nor U1135 (N_1135,N_558,N_360);
nand U1136 (N_1136,N_617,N_79);
nor U1137 (N_1137,N_78,N_462);
nor U1138 (N_1138,N_355,N_560);
and U1139 (N_1139,N_31,N_336);
nand U1140 (N_1140,N_673,N_337);
nand U1141 (N_1141,N_465,N_622);
and U1142 (N_1142,N_21,N_379);
and U1143 (N_1143,N_404,N_35);
nor U1144 (N_1144,N_583,N_568);
nor U1145 (N_1145,N_220,N_4);
or U1146 (N_1146,N_494,N_449);
and U1147 (N_1147,N_517,N_190);
nand U1148 (N_1148,N_428,N_159);
nand U1149 (N_1149,N_61,N_464);
and U1150 (N_1150,N_374,N_366);
nand U1151 (N_1151,N_132,N_73);
nor U1152 (N_1152,N_235,N_629);
nor U1153 (N_1153,N_680,N_609);
or U1154 (N_1154,N_604,N_538);
nor U1155 (N_1155,N_416,N_74);
and U1156 (N_1156,N_101,N_334);
nor U1157 (N_1157,N_56,N_438);
nor U1158 (N_1158,N_145,N_327);
nand U1159 (N_1159,N_701,N_747);
xor U1160 (N_1160,N_146,N_455);
nand U1161 (N_1161,N_738,N_305);
or U1162 (N_1162,N_504,N_450);
and U1163 (N_1163,N_652,N_445);
nor U1164 (N_1164,N_304,N_116);
nor U1165 (N_1165,N_257,N_45);
nand U1166 (N_1166,N_537,N_195);
or U1167 (N_1167,N_253,N_385);
and U1168 (N_1168,N_736,N_692);
nor U1169 (N_1169,N_342,N_445);
nand U1170 (N_1170,N_154,N_325);
nand U1171 (N_1171,N_4,N_400);
nand U1172 (N_1172,N_22,N_217);
nand U1173 (N_1173,N_395,N_540);
nand U1174 (N_1174,N_560,N_338);
and U1175 (N_1175,N_702,N_694);
nor U1176 (N_1176,N_102,N_466);
nand U1177 (N_1177,N_284,N_719);
and U1178 (N_1178,N_183,N_289);
nor U1179 (N_1179,N_74,N_145);
or U1180 (N_1180,N_713,N_462);
nor U1181 (N_1181,N_390,N_661);
or U1182 (N_1182,N_723,N_684);
nor U1183 (N_1183,N_200,N_506);
and U1184 (N_1184,N_117,N_608);
nor U1185 (N_1185,N_195,N_32);
or U1186 (N_1186,N_248,N_488);
or U1187 (N_1187,N_86,N_737);
or U1188 (N_1188,N_95,N_319);
nand U1189 (N_1189,N_45,N_459);
xnor U1190 (N_1190,N_392,N_201);
nand U1191 (N_1191,N_670,N_15);
nor U1192 (N_1192,N_18,N_264);
nand U1193 (N_1193,N_593,N_107);
or U1194 (N_1194,N_23,N_65);
xor U1195 (N_1195,N_162,N_421);
nor U1196 (N_1196,N_429,N_7);
and U1197 (N_1197,N_203,N_594);
nor U1198 (N_1198,N_429,N_232);
nand U1199 (N_1199,N_441,N_491);
nand U1200 (N_1200,N_438,N_447);
nand U1201 (N_1201,N_104,N_355);
and U1202 (N_1202,N_646,N_198);
nand U1203 (N_1203,N_732,N_702);
and U1204 (N_1204,N_41,N_237);
nand U1205 (N_1205,N_454,N_110);
nor U1206 (N_1206,N_391,N_614);
nand U1207 (N_1207,N_538,N_496);
and U1208 (N_1208,N_354,N_39);
or U1209 (N_1209,N_675,N_734);
xor U1210 (N_1210,N_454,N_530);
and U1211 (N_1211,N_297,N_175);
nand U1212 (N_1212,N_637,N_212);
or U1213 (N_1213,N_567,N_579);
xnor U1214 (N_1214,N_30,N_734);
or U1215 (N_1215,N_552,N_235);
nand U1216 (N_1216,N_729,N_33);
and U1217 (N_1217,N_322,N_722);
xnor U1218 (N_1218,N_531,N_33);
nand U1219 (N_1219,N_675,N_440);
or U1220 (N_1220,N_560,N_480);
nor U1221 (N_1221,N_136,N_309);
or U1222 (N_1222,N_622,N_573);
nand U1223 (N_1223,N_145,N_456);
nor U1224 (N_1224,N_246,N_109);
and U1225 (N_1225,N_457,N_67);
and U1226 (N_1226,N_495,N_218);
nand U1227 (N_1227,N_396,N_720);
nor U1228 (N_1228,N_147,N_5);
nand U1229 (N_1229,N_420,N_170);
and U1230 (N_1230,N_600,N_128);
and U1231 (N_1231,N_515,N_601);
xnor U1232 (N_1232,N_154,N_445);
or U1233 (N_1233,N_259,N_479);
and U1234 (N_1234,N_115,N_282);
or U1235 (N_1235,N_152,N_50);
nor U1236 (N_1236,N_146,N_247);
nand U1237 (N_1237,N_355,N_89);
nand U1238 (N_1238,N_14,N_182);
nand U1239 (N_1239,N_312,N_552);
nand U1240 (N_1240,N_185,N_288);
or U1241 (N_1241,N_35,N_593);
nand U1242 (N_1242,N_175,N_380);
xor U1243 (N_1243,N_240,N_664);
and U1244 (N_1244,N_698,N_48);
and U1245 (N_1245,N_406,N_58);
and U1246 (N_1246,N_417,N_546);
and U1247 (N_1247,N_308,N_423);
and U1248 (N_1248,N_252,N_647);
and U1249 (N_1249,N_477,N_326);
or U1250 (N_1250,N_485,N_303);
or U1251 (N_1251,N_409,N_345);
nor U1252 (N_1252,N_654,N_0);
nand U1253 (N_1253,N_530,N_40);
or U1254 (N_1254,N_684,N_678);
nand U1255 (N_1255,N_24,N_603);
or U1256 (N_1256,N_233,N_605);
nor U1257 (N_1257,N_172,N_320);
nand U1258 (N_1258,N_96,N_512);
nand U1259 (N_1259,N_78,N_519);
nand U1260 (N_1260,N_494,N_95);
nor U1261 (N_1261,N_321,N_299);
or U1262 (N_1262,N_410,N_387);
and U1263 (N_1263,N_618,N_329);
nor U1264 (N_1264,N_442,N_195);
nand U1265 (N_1265,N_524,N_82);
and U1266 (N_1266,N_387,N_274);
and U1267 (N_1267,N_261,N_416);
nor U1268 (N_1268,N_678,N_452);
nand U1269 (N_1269,N_665,N_205);
nor U1270 (N_1270,N_418,N_86);
xnor U1271 (N_1271,N_266,N_304);
or U1272 (N_1272,N_358,N_656);
and U1273 (N_1273,N_473,N_517);
nor U1274 (N_1274,N_130,N_629);
nand U1275 (N_1275,N_418,N_504);
nor U1276 (N_1276,N_436,N_390);
nand U1277 (N_1277,N_431,N_697);
xor U1278 (N_1278,N_212,N_714);
and U1279 (N_1279,N_137,N_290);
nand U1280 (N_1280,N_91,N_335);
or U1281 (N_1281,N_481,N_19);
nor U1282 (N_1282,N_545,N_199);
and U1283 (N_1283,N_88,N_348);
and U1284 (N_1284,N_303,N_636);
or U1285 (N_1285,N_671,N_117);
and U1286 (N_1286,N_295,N_190);
nor U1287 (N_1287,N_442,N_632);
and U1288 (N_1288,N_128,N_673);
and U1289 (N_1289,N_577,N_258);
and U1290 (N_1290,N_118,N_481);
xor U1291 (N_1291,N_746,N_493);
or U1292 (N_1292,N_588,N_413);
nand U1293 (N_1293,N_399,N_650);
nor U1294 (N_1294,N_150,N_672);
or U1295 (N_1295,N_37,N_661);
or U1296 (N_1296,N_302,N_116);
or U1297 (N_1297,N_232,N_202);
or U1298 (N_1298,N_536,N_341);
xor U1299 (N_1299,N_649,N_262);
or U1300 (N_1300,N_282,N_108);
nand U1301 (N_1301,N_636,N_401);
nor U1302 (N_1302,N_149,N_98);
nand U1303 (N_1303,N_92,N_86);
xor U1304 (N_1304,N_437,N_269);
nand U1305 (N_1305,N_575,N_399);
and U1306 (N_1306,N_233,N_163);
nand U1307 (N_1307,N_527,N_404);
or U1308 (N_1308,N_592,N_251);
nor U1309 (N_1309,N_53,N_363);
or U1310 (N_1310,N_298,N_744);
xnor U1311 (N_1311,N_278,N_654);
nor U1312 (N_1312,N_103,N_280);
nor U1313 (N_1313,N_590,N_400);
nand U1314 (N_1314,N_272,N_122);
nor U1315 (N_1315,N_682,N_73);
nor U1316 (N_1316,N_156,N_72);
xnor U1317 (N_1317,N_93,N_462);
xnor U1318 (N_1318,N_547,N_200);
xnor U1319 (N_1319,N_120,N_78);
nor U1320 (N_1320,N_647,N_450);
nor U1321 (N_1321,N_159,N_724);
nand U1322 (N_1322,N_447,N_681);
nand U1323 (N_1323,N_393,N_40);
nand U1324 (N_1324,N_736,N_715);
nor U1325 (N_1325,N_61,N_42);
and U1326 (N_1326,N_481,N_604);
nand U1327 (N_1327,N_110,N_106);
nand U1328 (N_1328,N_347,N_145);
nor U1329 (N_1329,N_197,N_328);
or U1330 (N_1330,N_162,N_427);
nor U1331 (N_1331,N_77,N_177);
nand U1332 (N_1332,N_18,N_207);
or U1333 (N_1333,N_512,N_453);
and U1334 (N_1334,N_192,N_168);
or U1335 (N_1335,N_189,N_124);
nand U1336 (N_1336,N_607,N_688);
and U1337 (N_1337,N_603,N_434);
nand U1338 (N_1338,N_232,N_226);
nor U1339 (N_1339,N_608,N_725);
nor U1340 (N_1340,N_490,N_82);
nand U1341 (N_1341,N_579,N_621);
nand U1342 (N_1342,N_560,N_267);
nand U1343 (N_1343,N_620,N_124);
or U1344 (N_1344,N_29,N_513);
nand U1345 (N_1345,N_177,N_284);
nand U1346 (N_1346,N_473,N_9);
or U1347 (N_1347,N_627,N_501);
nand U1348 (N_1348,N_263,N_88);
xnor U1349 (N_1349,N_726,N_359);
and U1350 (N_1350,N_444,N_651);
nor U1351 (N_1351,N_732,N_495);
nand U1352 (N_1352,N_437,N_336);
nor U1353 (N_1353,N_482,N_332);
nand U1354 (N_1354,N_455,N_357);
or U1355 (N_1355,N_35,N_110);
or U1356 (N_1356,N_409,N_536);
xnor U1357 (N_1357,N_522,N_643);
and U1358 (N_1358,N_381,N_342);
nand U1359 (N_1359,N_124,N_222);
nand U1360 (N_1360,N_635,N_744);
and U1361 (N_1361,N_217,N_428);
nor U1362 (N_1362,N_174,N_178);
nor U1363 (N_1363,N_379,N_228);
and U1364 (N_1364,N_448,N_103);
or U1365 (N_1365,N_351,N_574);
xnor U1366 (N_1366,N_122,N_254);
or U1367 (N_1367,N_293,N_45);
or U1368 (N_1368,N_688,N_745);
or U1369 (N_1369,N_493,N_354);
nand U1370 (N_1370,N_275,N_446);
nor U1371 (N_1371,N_213,N_39);
nor U1372 (N_1372,N_382,N_481);
nand U1373 (N_1373,N_495,N_502);
nor U1374 (N_1374,N_254,N_336);
or U1375 (N_1375,N_630,N_536);
nor U1376 (N_1376,N_727,N_274);
or U1377 (N_1377,N_319,N_520);
nor U1378 (N_1378,N_123,N_691);
or U1379 (N_1379,N_188,N_735);
nand U1380 (N_1380,N_703,N_146);
nor U1381 (N_1381,N_305,N_362);
and U1382 (N_1382,N_376,N_611);
nand U1383 (N_1383,N_241,N_372);
nand U1384 (N_1384,N_537,N_71);
nor U1385 (N_1385,N_729,N_568);
nor U1386 (N_1386,N_610,N_32);
nor U1387 (N_1387,N_311,N_551);
nor U1388 (N_1388,N_403,N_465);
nand U1389 (N_1389,N_453,N_687);
and U1390 (N_1390,N_387,N_681);
nor U1391 (N_1391,N_502,N_111);
or U1392 (N_1392,N_279,N_319);
nor U1393 (N_1393,N_412,N_323);
xor U1394 (N_1394,N_536,N_31);
and U1395 (N_1395,N_133,N_533);
or U1396 (N_1396,N_255,N_282);
or U1397 (N_1397,N_160,N_569);
nor U1398 (N_1398,N_217,N_250);
or U1399 (N_1399,N_295,N_80);
nand U1400 (N_1400,N_161,N_580);
or U1401 (N_1401,N_635,N_636);
and U1402 (N_1402,N_699,N_267);
or U1403 (N_1403,N_18,N_466);
nor U1404 (N_1404,N_680,N_411);
or U1405 (N_1405,N_603,N_324);
nor U1406 (N_1406,N_632,N_88);
or U1407 (N_1407,N_37,N_410);
xor U1408 (N_1408,N_126,N_470);
and U1409 (N_1409,N_206,N_300);
and U1410 (N_1410,N_562,N_89);
nand U1411 (N_1411,N_422,N_19);
xnor U1412 (N_1412,N_680,N_24);
and U1413 (N_1413,N_358,N_232);
and U1414 (N_1414,N_502,N_546);
or U1415 (N_1415,N_122,N_173);
nor U1416 (N_1416,N_722,N_156);
and U1417 (N_1417,N_195,N_624);
nand U1418 (N_1418,N_534,N_66);
nand U1419 (N_1419,N_451,N_195);
nand U1420 (N_1420,N_681,N_5);
nor U1421 (N_1421,N_234,N_550);
and U1422 (N_1422,N_527,N_304);
and U1423 (N_1423,N_656,N_359);
nand U1424 (N_1424,N_666,N_441);
nor U1425 (N_1425,N_702,N_441);
nand U1426 (N_1426,N_160,N_2);
or U1427 (N_1427,N_220,N_612);
nand U1428 (N_1428,N_624,N_571);
and U1429 (N_1429,N_24,N_307);
nand U1430 (N_1430,N_412,N_38);
nor U1431 (N_1431,N_177,N_242);
nor U1432 (N_1432,N_591,N_494);
and U1433 (N_1433,N_89,N_676);
nor U1434 (N_1434,N_271,N_46);
and U1435 (N_1435,N_741,N_739);
nand U1436 (N_1436,N_333,N_178);
and U1437 (N_1437,N_661,N_33);
and U1438 (N_1438,N_567,N_622);
or U1439 (N_1439,N_214,N_558);
and U1440 (N_1440,N_452,N_565);
and U1441 (N_1441,N_332,N_231);
nor U1442 (N_1442,N_599,N_185);
or U1443 (N_1443,N_654,N_268);
nor U1444 (N_1444,N_475,N_612);
nand U1445 (N_1445,N_252,N_253);
and U1446 (N_1446,N_489,N_539);
nand U1447 (N_1447,N_280,N_155);
or U1448 (N_1448,N_379,N_544);
and U1449 (N_1449,N_733,N_344);
or U1450 (N_1450,N_243,N_194);
nor U1451 (N_1451,N_414,N_440);
nand U1452 (N_1452,N_502,N_304);
xnor U1453 (N_1453,N_545,N_147);
or U1454 (N_1454,N_436,N_295);
or U1455 (N_1455,N_69,N_334);
or U1456 (N_1456,N_41,N_725);
nor U1457 (N_1457,N_201,N_294);
xnor U1458 (N_1458,N_543,N_349);
nor U1459 (N_1459,N_602,N_66);
or U1460 (N_1460,N_630,N_692);
xnor U1461 (N_1461,N_121,N_42);
and U1462 (N_1462,N_657,N_331);
nand U1463 (N_1463,N_341,N_700);
and U1464 (N_1464,N_384,N_416);
or U1465 (N_1465,N_348,N_275);
or U1466 (N_1466,N_618,N_163);
nand U1467 (N_1467,N_453,N_476);
and U1468 (N_1468,N_72,N_288);
and U1469 (N_1469,N_256,N_156);
and U1470 (N_1470,N_529,N_289);
and U1471 (N_1471,N_662,N_434);
nor U1472 (N_1472,N_340,N_135);
or U1473 (N_1473,N_611,N_104);
nor U1474 (N_1474,N_385,N_530);
and U1475 (N_1475,N_218,N_570);
and U1476 (N_1476,N_372,N_36);
nor U1477 (N_1477,N_194,N_56);
or U1478 (N_1478,N_404,N_356);
nand U1479 (N_1479,N_132,N_104);
nor U1480 (N_1480,N_396,N_170);
and U1481 (N_1481,N_219,N_235);
nor U1482 (N_1482,N_294,N_280);
and U1483 (N_1483,N_158,N_635);
and U1484 (N_1484,N_257,N_220);
xor U1485 (N_1485,N_604,N_101);
nand U1486 (N_1486,N_132,N_660);
nand U1487 (N_1487,N_641,N_465);
nand U1488 (N_1488,N_10,N_679);
or U1489 (N_1489,N_680,N_409);
nor U1490 (N_1490,N_170,N_709);
nor U1491 (N_1491,N_205,N_10);
and U1492 (N_1492,N_173,N_95);
or U1493 (N_1493,N_712,N_725);
nor U1494 (N_1494,N_39,N_79);
nor U1495 (N_1495,N_140,N_84);
nor U1496 (N_1496,N_74,N_385);
nand U1497 (N_1497,N_76,N_563);
nand U1498 (N_1498,N_219,N_126);
or U1499 (N_1499,N_305,N_184);
or U1500 (N_1500,N_1161,N_1025);
xnor U1501 (N_1501,N_849,N_783);
nand U1502 (N_1502,N_1198,N_1176);
or U1503 (N_1503,N_808,N_1345);
nor U1504 (N_1504,N_768,N_934);
nor U1505 (N_1505,N_1071,N_1319);
and U1506 (N_1506,N_1196,N_840);
xnor U1507 (N_1507,N_1094,N_805);
and U1508 (N_1508,N_886,N_1290);
xor U1509 (N_1509,N_1070,N_1254);
nand U1510 (N_1510,N_809,N_833);
nand U1511 (N_1511,N_967,N_1495);
and U1512 (N_1512,N_1143,N_1440);
and U1513 (N_1513,N_1314,N_1037);
nor U1514 (N_1514,N_885,N_859);
nand U1515 (N_1515,N_1115,N_831);
nand U1516 (N_1516,N_865,N_1239);
and U1517 (N_1517,N_1077,N_1051);
or U1518 (N_1518,N_1043,N_1388);
or U1519 (N_1519,N_829,N_998);
nor U1520 (N_1520,N_837,N_1179);
xnor U1521 (N_1521,N_867,N_1112);
xnor U1522 (N_1522,N_1018,N_1020);
xor U1523 (N_1523,N_1191,N_1142);
and U1524 (N_1524,N_1318,N_1009);
nor U1525 (N_1525,N_1230,N_1151);
nand U1526 (N_1526,N_1412,N_1086);
or U1527 (N_1527,N_980,N_990);
nor U1528 (N_1528,N_1117,N_1288);
nor U1529 (N_1529,N_917,N_1247);
xnor U1530 (N_1530,N_1449,N_931);
nor U1531 (N_1531,N_1425,N_1453);
xnor U1532 (N_1532,N_1457,N_858);
nand U1533 (N_1533,N_1067,N_1418);
and U1534 (N_1534,N_1478,N_1378);
and U1535 (N_1535,N_924,N_1262);
nand U1536 (N_1536,N_825,N_1365);
xnor U1537 (N_1537,N_1178,N_1032);
nor U1538 (N_1538,N_894,N_1058);
and U1539 (N_1539,N_953,N_977);
and U1540 (N_1540,N_943,N_1344);
nand U1541 (N_1541,N_1061,N_817);
or U1542 (N_1542,N_951,N_1012);
nor U1543 (N_1543,N_772,N_1223);
nor U1544 (N_1544,N_1097,N_1141);
and U1545 (N_1545,N_1225,N_972);
nand U1546 (N_1546,N_1181,N_1099);
nand U1547 (N_1547,N_1232,N_1209);
nand U1548 (N_1548,N_1486,N_1108);
nor U1549 (N_1549,N_1039,N_774);
nand U1550 (N_1550,N_845,N_1040);
xor U1551 (N_1551,N_781,N_856);
xor U1552 (N_1552,N_1121,N_920);
and U1553 (N_1553,N_1361,N_1407);
nor U1554 (N_1554,N_810,N_806);
and U1555 (N_1555,N_1304,N_1217);
and U1556 (N_1556,N_1251,N_1311);
nor U1557 (N_1557,N_933,N_1190);
nor U1558 (N_1558,N_1171,N_974);
or U1559 (N_1559,N_1122,N_883);
and U1560 (N_1560,N_893,N_841);
xnor U1561 (N_1561,N_1477,N_759);
nand U1562 (N_1562,N_1134,N_982);
nand U1563 (N_1563,N_1085,N_821);
and U1564 (N_1564,N_1158,N_1422);
or U1565 (N_1565,N_1283,N_1308);
and U1566 (N_1566,N_1256,N_1253);
nor U1567 (N_1567,N_1342,N_964);
or U1568 (N_1568,N_1332,N_873);
or U1569 (N_1569,N_1033,N_1102);
nor U1570 (N_1570,N_1474,N_1348);
nor U1571 (N_1571,N_1073,N_877);
nand U1572 (N_1572,N_1007,N_1420);
xor U1573 (N_1573,N_1464,N_1231);
and U1574 (N_1574,N_1056,N_1369);
and U1575 (N_1575,N_1416,N_756);
nor U1576 (N_1576,N_1368,N_1060);
or U1577 (N_1577,N_1057,N_1078);
nor U1578 (N_1578,N_887,N_947);
and U1579 (N_1579,N_1444,N_1303);
xnor U1580 (N_1580,N_970,N_1170);
and U1581 (N_1581,N_1499,N_1350);
nand U1582 (N_1582,N_969,N_1207);
and U1583 (N_1583,N_1343,N_1458);
and U1584 (N_1584,N_814,N_860);
nand U1585 (N_1585,N_959,N_1364);
or U1586 (N_1586,N_1356,N_1131);
and U1587 (N_1587,N_1355,N_767);
nand U1588 (N_1588,N_1116,N_1469);
or U1589 (N_1589,N_762,N_1245);
and U1590 (N_1590,N_765,N_1392);
nor U1591 (N_1591,N_1016,N_1448);
nor U1592 (N_1592,N_1295,N_1341);
and U1593 (N_1593,N_1307,N_1405);
nor U1594 (N_1594,N_985,N_863);
xnor U1595 (N_1595,N_1320,N_1049);
nor U1596 (N_1596,N_791,N_854);
nor U1597 (N_1597,N_1358,N_950);
nand U1598 (N_1598,N_798,N_1235);
nor U1599 (N_1599,N_789,N_991);
or U1600 (N_1600,N_761,N_1466);
nor U1601 (N_1601,N_866,N_1136);
nand U1602 (N_1602,N_935,N_842);
or U1603 (N_1603,N_1296,N_1492);
nand U1604 (N_1604,N_1434,N_1423);
nand U1605 (N_1605,N_1278,N_910);
and U1606 (N_1606,N_989,N_795);
and U1607 (N_1607,N_790,N_1447);
or U1608 (N_1608,N_1175,N_846);
or U1609 (N_1609,N_1010,N_1273);
nor U1610 (N_1610,N_1059,N_1024);
nor U1611 (N_1611,N_1221,N_952);
and U1612 (N_1612,N_1274,N_981);
or U1613 (N_1613,N_1306,N_876);
xnor U1614 (N_1614,N_1322,N_1242);
or U1615 (N_1615,N_927,N_912);
nor U1616 (N_1616,N_1383,N_929);
nor U1617 (N_1617,N_1427,N_1252);
and U1618 (N_1618,N_1475,N_1431);
and U1619 (N_1619,N_1334,N_987);
and U1620 (N_1620,N_1488,N_1233);
or U1621 (N_1621,N_1485,N_1321);
nor U1622 (N_1622,N_822,N_1005);
and U1623 (N_1623,N_1271,N_764);
nand U1624 (N_1624,N_971,N_1026);
or U1625 (N_1625,N_913,N_1132);
and U1626 (N_1626,N_1015,N_1034);
nor U1627 (N_1627,N_948,N_1200);
nand U1628 (N_1628,N_1091,N_797);
and U1629 (N_1629,N_1272,N_757);
and U1630 (N_1630,N_1479,N_1194);
nand U1631 (N_1631,N_1301,N_1246);
and U1632 (N_1632,N_1030,N_1443);
or U1633 (N_1633,N_1195,N_1244);
nor U1634 (N_1634,N_796,N_996);
xor U1635 (N_1635,N_1206,N_1090);
nand U1636 (N_1636,N_1236,N_1397);
nor U1637 (N_1637,N_1384,N_1381);
nand U1638 (N_1638,N_1192,N_1144);
and U1639 (N_1639,N_1360,N_961);
nand U1640 (N_1640,N_1048,N_1113);
or U1641 (N_1641,N_864,N_1315);
and U1642 (N_1642,N_1385,N_901);
nand U1643 (N_1643,N_1297,N_1075);
nor U1644 (N_1644,N_1014,N_1154);
and U1645 (N_1645,N_1261,N_1180);
nor U1646 (N_1646,N_1399,N_750);
nand U1647 (N_1647,N_823,N_1463);
xor U1648 (N_1648,N_811,N_1237);
nor U1649 (N_1649,N_1001,N_992);
nand U1650 (N_1650,N_1189,N_1064);
nor U1651 (N_1651,N_786,N_1337);
nor U1652 (N_1652,N_1096,N_1489);
nand U1653 (N_1653,N_1177,N_1352);
nor U1654 (N_1654,N_1011,N_1027);
nand U1655 (N_1655,N_843,N_1199);
xor U1656 (N_1656,N_1211,N_919);
nor U1657 (N_1657,N_1159,N_1260);
nand U1658 (N_1658,N_1228,N_1292);
or U1659 (N_1659,N_1462,N_1240);
and U1660 (N_1660,N_1339,N_780);
nand U1661 (N_1661,N_986,N_1391);
or U1662 (N_1662,N_874,N_1327);
xnor U1663 (N_1663,N_1249,N_1490);
or U1664 (N_1664,N_1476,N_1081);
and U1665 (N_1665,N_872,N_1417);
and U1666 (N_1666,N_1493,N_1413);
xnor U1667 (N_1667,N_949,N_1268);
nand U1668 (N_1668,N_1351,N_1193);
nor U1669 (N_1669,N_835,N_1266);
xnor U1670 (N_1670,N_1347,N_1396);
or U1671 (N_1671,N_1286,N_1394);
nand U1672 (N_1672,N_923,N_1287);
xnor U1673 (N_1673,N_1335,N_1269);
or U1674 (N_1674,N_1386,N_1205);
nor U1675 (N_1675,N_1038,N_1021);
and U1676 (N_1676,N_928,N_1291);
and U1677 (N_1677,N_1183,N_1432);
or U1678 (N_1678,N_1101,N_936);
nor U1679 (N_1679,N_994,N_1324);
nor U1680 (N_1680,N_875,N_1002);
or U1681 (N_1681,N_1069,N_1046);
or U1682 (N_1682,N_851,N_1155);
nand U1683 (N_1683,N_784,N_1338);
nor U1684 (N_1684,N_899,N_1241);
nor U1685 (N_1685,N_1406,N_1461);
nor U1686 (N_1686,N_1250,N_881);
or U1687 (N_1687,N_1215,N_1340);
nor U1688 (N_1688,N_1293,N_914);
and U1689 (N_1689,N_1050,N_778);
nor U1690 (N_1690,N_787,N_1367);
nand U1691 (N_1691,N_1036,N_1052);
and U1692 (N_1692,N_1310,N_946);
nand U1693 (N_1693,N_1389,N_869);
and U1694 (N_1694,N_1202,N_960);
xor U1695 (N_1695,N_853,N_1390);
and U1696 (N_1696,N_1210,N_1088);
or U1697 (N_1697,N_938,N_1277);
and U1698 (N_1698,N_1430,N_820);
nor U1699 (N_1699,N_847,N_1387);
nor U1700 (N_1700,N_1325,N_1095);
nand U1701 (N_1701,N_1238,N_1234);
nand U1702 (N_1702,N_816,N_1186);
nor U1703 (N_1703,N_1465,N_1068);
and U1704 (N_1704,N_1008,N_802);
xnor U1705 (N_1705,N_1197,N_1300);
or U1706 (N_1706,N_1433,N_1137);
or U1707 (N_1707,N_1316,N_1375);
nand U1708 (N_1708,N_1126,N_1135);
nand U1709 (N_1709,N_1395,N_1419);
nand U1710 (N_1710,N_958,N_978);
or U1711 (N_1711,N_1006,N_1333);
nor U1712 (N_1712,N_1227,N_909);
nor U1713 (N_1713,N_1129,N_1166);
nand U1714 (N_1714,N_1243,N_1082);
or U1715 (N_1715,N_1289,N_1302);
or U1716 (N_1716,N_1019,N_792);
nor U1717 (N_1717,N_776,N_888);
nand U1718 (N_1718,N_1362,N_896);
nand U1719 (N_1719,N_771,N_838);
nor U1720 (N_1720,N_1226,N_1029);
and U1721 (N_1721,N_779,N_1424);
and U1722 (N_1722,N_1473,N_1281);
or U1723 (N_1723,N_1372,N_782);
and U1724 (N_1724,N_1053,N_908);
and U1725 (N_1725,N_916,N_1214);
and U1726 (N_1726,N_1363,N_1164);
and U1727 (N_1727,N_1063,N_1089);
or U1728 (N_1728,N_1098,N_1201);
or U1729 (N_1729,N_1437,N_1258);
and U1730 (N_1730,N_1248,N_1468);
and U1731 (N_1731,N_1152,N_836);
nand U1732 (N_1732,N_769,N_882);
xor U1733 (N_1733,N_1275,N_1328);
nor U1734 (N_1734,N_852,N_1376);
nand U1735 (N_1735,N_1471,N_1280);
or U1736 (N_1736,N_1054,N_754);
or U1737 (N_1737,N_1435,N_1371);
xor U1738 (N_1738,N_1087,N_1445);
and U1739 (N_1739,N_1487,N_1401);
and U1740 (N_1740,N_760,N_925);
nand U1741 (N_1741,N_1162,N_1213);
or U1742 (N_1742,N_1467,N_889);
and U1743 (N_1743,N_944,N_1373);
or U1744 (N_1744,N_1284,N_812);
nor U1745 (N_1745,N_1188,N_1150);
and U1746 (N_1746,N_857,N_1497);
or U1747 (N_1747,N_1279,N_1404);
nand U1748 (N_1748,N_1106,N_895);
and U1749 (N_1749,N_1374,N_1276);
and U1750 (N_1750,N_844,N_879);
or U1751 (N_1751,N_1346,N_751);
and U1752 (N_1752,N_1400,N_1439);
xor U1753 (N_1753,N_907,N_1402);
or U1754 (N_1754,N_1168,N_1204);
nand U1755 (N_1755,N_997,N_870);
and U1756 (N_1756,N_1042,N_1124);
nor U1757 (N_1757,N_1379,N_1410);
nor U1758 (N_1758,N_1366,N_1072);
and U1759 (N_1759,N_880,N_800);
xnor U1760 (N_1760,N_1481,N_1173);
nand U1761 (N_1761,N_1045,N_1357);
nand U1762 (N_1762,N_1265,N_1031);
and U1763 (N_1763,N_1496,N_1083);
and U1764 (N_1764,N_956,N_1110);
and U1765 (N_1765,N_1222,N_1153);
or U1766 (N_1766,N_1047,N_973);
nand U1767 (N_1767,N_890,N_884);
nand U1768 (N_1768,N_794,N_1294);
and U1769 (N_1769,N_1455,N_1148);
and U1770 (N_1770,N_1174,N_1220);
or U1771 (N_1771,N_1156,N_945);
xor U1772 (N_1772,N_1118,N_1403);
and U1773 (N_1773,N_1013,N_1359);
or U1774 (N_1774,N_1330,N_1123);
nand U1775 (N_1775,N_1229,N_1442);
or U1776 (N_1776,N_1000,N_993);
or U1777 (N_1777,N_1336,N_891);
nor U1778 (N_1778,N_1218,N_1128);
and U1779 (N_1779,N_1264,N_1105);
and U1780 (N_1780,N_892,N_932);
and U1781 (N_1781,N_1120,N_1414);
nor U1782 (N_1782,N_1160,N_1035);
nand U1783 (N_1783,N_1323,N_1259);
nor U1784 (N_1784,N_1454,N_753);
or U1785 (N_1785,N_1329,N_966);
nand U1786 (N_1786,N_1100,N_1257);
xor U1787 (N_1787,N_1149,N_801);
nor U1788 (N_1788,N_871,N_1103);
nor U1789 (N_1789,N_770,N_826);
nor U1790 (N_1790,N_1139,N_1353);
nor U1791 (N_1791,N_1393,N_1456);
nand U1792 (N_1792,N_1438,N_1411);
or U1793 (N_1793,N_1145,N_1023);
nand U1794 (N_1794,N_1165,N_1426);
nand U1795 (N_1795,N_1182,N_905);
or U1796 (N_1796,N_1298,N_775);
or U1797 (N_1797,N_773,N_1219);
nor U1798 (N_1798,N_855,N_902);
or U1799 (N_1799,N_1498,N_1451);
and U1800 (N_1800,N_955,N_979);
and U1801 (N_1801,N_1491,N_1157);
and U1802 (N_1802,N_1109,N_1133);
or U1803 (N_1803,N_1354,N_832);
nand U1804 (N_1804,N_861,N_807);
nor U1805 (N_1805,N_954,N_939);
and U1806 (N_1806,N_763,N_1460);
nand U1807 (N_1807,N_819,N_926);
nand U1808 (N_1808,N_799,N_1080);
xor U1809 (N_1809,N_1107,N_999);
xor U1810 (N_1810,N_1470,N_1494);
nor U1811 (N_1811,N_1065,N_868);
and U1812 (N_1812,N_975,N_1282);
or U1813 (N_1813,N_1267,N_906);
and U1814 (N_1814,N_1169,N_1482);
and U1815 (N_1815,N_1111,N_1185);
or U1816 (N_1816,N_755,N_827);
and U1817 (N_1817,N_1119,N_828);
xnor U1818 (N_1818,N_1472,N_1450);
nand U1819 (N_1819,N_793,N_1044);
nor U1820 (N_1820,N_1312,N_1066);
nor U1821 (N_1821,N_777,N_1125);
nor U1822 (N_1822,N_1184,N_1428);
nor U1823 (N_1823,N_1130,N_1299);
or U1824 (N_1824,N_1409,N_1140);
and U1825 (N_1825,N_1483,N_1421);
nor U1826 (N_1826,N_1446,N_1041);
and U1827 (N_1827,N_862,N_1370);
nor U1828 (N_1828,N_803,N_1441);
or U1829 (N_1829,N_1212,N_1146);
nand U1830 (N_1830,N_976,N_850);
nand U1831 (N_1831,N_1084,N_988);
or U1832 (N_1832,N_1377,N_900);
xnor U1833 (N_1833,N_1216,N_824);
nand U1834 (N_1834,N_1452,N_965);
nor U1835 (N_1835,N_940,N_1429);
nand U1836 (N_1836,N_942,N_1167);
nor U1837 (N_1837,N_1459,N_834);
nor U1838 (N_1838,N_1092,N_1255);
or U1839 (N_1839,N_1172,N_962);
or U1840 (N_1840,N_1309,N_941);
nand U1841 (N_1841,N_922,N_937);
and U1842 (N_1842,N_1076,N_1127);
and U1843 (N_1843,N_1331,N_1163);
and U1844 (N_1844,N_1436,N_804);
nand U1845 (N_1845,N_1022,N_957);
and U1846 (N_1846,N_1263,N_1003);
and U1847 (N_1847,N_1104,N_815);
or U1848 (N_1848,N_1055,N_758);
or U1849 (N_1849,N_1203,N_878);
or U1850 (N_1850,N_904,N_1017);
nor U1851 (N_1851,N_1398,N_911);
nand U1852 (N_1852,N_918,N_1349);
or U1853 (N_1853,N_898,N_1028);
nor U1854 (N_1854,N_818,N_897);
nand U1855 (N_1855,N_983,N_921);
or U1856 (N_1856,N_1484,N_984);
and U1857 (N_1857,N_1147,N_968);
nand U1858 (N_1858,N_785,N_1380);
and U1859 (N_1859,N_1313,N_1326);
and U1860 (N_1860,N_766,N_1270);
nand U1861 (N_1861,N_1079,N_1317);
xor U1862 (N_1862,N_1062,N_1187);
or U1863 (N_1863,N_788,N_752);
nand U1864 (N_1864,N_1480,N_1285);
nor U1865 (N_1865,N_839,N_1114);
or U1866 (N_1866,N_830,N_963);
nor U1867 (N_1867,N_1004,N_915);
or U1868 (N_1868,N_1093,N_1224);
and U1869 (N_1869,N_1305,N_1074);
nor U1870 (N_1870,N_1382,N_1408);
and U1871 (N_1871,N_1138,N_995);
xor U1872 (N_1872,N_1208,N_930);
nor U1873 (N_1873,N_848,N_1415);
or U1874 (N_1874,N_813,N_903);
or U1875 (N_1875,N_814,N_1387);
nor U1876 (N_1876,N_1108,N_1294);
or U1877 (N_1877,N_851,N_1175);
xnor U1878 (N_1878,N_1307,N_1299);
nand U1879 (N_1879,N_931,N_1434);
or U1880 (N_1880,N_1317,N_882);
and U1881 (N_1881,N_1478,N_1091);
nor U1882 (N_1882,N_1452,N_1481);
or U1883 (N_1883,N_870,N_1332);
nand U1884 (N_1884,N_799,N_1349);
and U1885 (N_1885,N_1227,N_1329);
nor U1886 (N_1886,N_789,N_1289);
nand U1887 (N_1887,N_1084,N_1351);
xor U1888 (N_1888,N_1086,N_1480);
or U1889 (N_1889,N_1366,N_1143);
nor U1890 (N_1890,N_1065,N_840);
and U1891 (N_1891,N_1078,N_1499);
nand U1892 (N_1892,N_1013,N_1118);
nand U1893 (N_1893,N_1035,N_753);
and U1894 (N_1894,N_967,N_979);
and U1895 (N_1895,N_1476,N_871);
and U1896 (N_1896,N_824,N_1259);
and U1897 (N_1897,N_1116,N_1496);
nor U1898 (N_1898,N_1378,N_1358);
xor U1899 (N_1899,N_1369,N_1066);
nor U1900 (N_1900,N_1025,N_1353);
or U1901 (N_1901,N_1185,N_1287);
nor U1902 (N_1902,N_867,N_877);
nand U1903 (N_1903,N_1411,N_1467);
xnor U1904 (N_1904,N_1252,N_914);
nor U1905 (N_1905,N_1046,N_845);
or U1906 (N_1906,N_1074,N_1211);
nor U1907 (N_1907,N_1205,N_1127);
and U1908 (N_1908,N_1157,N_970);
nand U1909 (N_1909,N_775,N_1044);
xnor U1910 (N_1910,N_864,N_1004);
xnor U1911 (N_1911,N_892,N_1146);
or U1912 (N_1912,N_1349,N_1028);
nor U1913 (N_1913,N_1422,N_803);
or U1914 (N_1914,N_1295,N_1167);
or U1915 (N_1915,N_857,N_880);
nor U1916 (N_1916,N_807,N_1195);
or U1917 (N_1917,N_954,N_1121);
or U1918 (N_1918,N_1119,N_959);
xor U1919 (N_1919,N_1206,N_1039);
and U1920 (N_1920,N_1424,N_863);
nand U1921 (N_1921,N_1307,N_1206);
and U1922 (N_1922,N_1257,N_859);
nand U1923 (N_1923,N_1397,N_1048);
nor U1924 (N_1924,N_1024,N_1251);
and U1925 (N_1925,N_920,N_1151);
nand U1926 (N_1926,N_1267,N_1243);
and U1927 (N_1927,N_1173,N_1189);
or U1928 (N_1928,N_1409,N_1172);
and U1929 (N_1929,N_852,N_1292);
and U1930 (N_1930,N_1345,N_1080);
or U1931 (N_1931,N_773,N_1372);
nor U1932 (N_1932,N_1251,N_1135);
nor U1933 (N_1933,N_1160,N_802);
nand U1934 (N_1934,N_1251,N_1488);
or U1935 (N_1935,N_872,N_1057);
nor U1936 (N_1936,N_1396,N_1129);
or U1937 (N_1937,N_1060,N_1135);
nor U1938 (N_1938,N_1497,N_761);
nor U1939 (N_1939,N_1360,N_1206);
nor U1940 (N_1940,N_944,N_1244);
nor U1941 (N_1941,N_1263,N_989);
nand U1942 (N_1942,N_771,N_785);
and U1943 (N_1943,N_1385,N_1052);
nor U1944 (N_1944,N_1197,N_1344);
nand U1945 (N_1945,N_1416,N_1188);
or U1946 (N_1946,N_973,N_1154);
nand U1947 (N_1947,N_1050,N_1314);
xor U1948 (N_1948,N_808,N_964);
xor U1949 (N_1949,N_1125,N_1088);
nand U1950 (N_1950,N_917,N_1303);
nand U1951 (N_1951,N_912,N_960);
xnor U1952 (N_1952,N_777,N_1253);
nand U1953 (N_1953,N_1202,N_922);
nand U1954 (N_1954,N_1392,N_1208);
or U1955 (N_1955,N_754,N_1297);
or U1956 (N_1956,N_950,N_1475);
and U1957 (N_1957,N_1295,N_1498);
and U1958 (N_1958,N_1226,N_882);
and U1959 (N_1959,N_1198,N_788);
nand U1960 (N_1960,N_1384,N_1130);
or U1961 (N_1961,N_1315,N_1128);
and U1962 (N_1962,N_1353,N_1054);
or U1963 (N_1963,N_1010,N_1114);
and U1964 (N_1964,N_807,N_1298);
and U1965 (N_1965,N_1404,N_954);
nor U1966 (N_1966,N_1036,N_1336);
xnor U1967 (N_1967,N_820,N_1491);
and U1968 (N_1968,N_907,N_1166);
nor U1969 (N_1969,N_1486,N_1364);
nor U1970 (N_1970,N_1050,N_1372);
xnor U1971 (N_1971,N_969,N_899);
xor U1972 (N_1972,N_1283,N_870);
or U1973 (N_1973,N_1347,N_1009);
or U1974 (N_1974,N_955,N_812);
xor U1975 (N_1975,N_1221,N_781);
xnor U1976 (N_1976,N_1036,N_1106);
nor U1977 (N_1977,N_921,N_1026);
nand U1978 (N_1978,N_866,N_885);
or U1979 (N_1979,N_996,N_1493);
nor U1980 (N_1980,N_775,N_1435);
xor U1981 (N_1981,N_1416,N_1054);
nor U1982 (N_1982,N_859,N_1223);
nand U1983 (N_1983,N_1079,N_1217);
nor U1984 (N_1984,N_929,N_815);
xor U1985 (N_1985,N_1475,N_1241);
nand U1986 (N_1986,N_1319,N_1152);
nand U1987 (N_1987,N_1369,N_1256);
nor U1988 (N_1988,N_952,N_782);
nor U1989 (N_1989,N_1397,N_750);
nand U1990 (N_1990,N_1465,N_1310);
nand U1991 (N_1991,N_933,N_1159);
xor U1992 (N_1992,N_966,N_1487);
and U1993 (N_1993,N_753,N_1040);
and U1994 (N_1994,N_821,N_1165);
xor U1995 (N_1995,N_1349,N_1436);
and U1996 (N_1996,N_999,N_1203);
or U1997 (N_1997,N_931,N_1353);
nor U1998 (N_1998,N_924,N_1061);
nor U1999 (N_1999,N_1392,N_904);
nor U2000 (N_2000,N_882,N_786);
xor U2001 (N_2001,N_1441,N_1393);
and U2002 (N_2002,N_1031,N_1121);
or U2003 (N_2003,N_861,N_1449);
or U2004 (N_2004,N_1244,N_975);
nor U2005 (N_2005,N_1339,N_1463);
nand U2006 (N_2006,N_1052,N_1434);
xor U2007 (N_2007,N_1357,N_1386);
nand U2008 (N_2008,N_1356,N_1005);
nor U2009 (N_2009,N_1303,N_1126);
nor U2010 (N_2010,N_1005,N_1318);
nand U2011 (N_2011,N_1095,N_873);
or U2012 (N_2012,N_1376,N_1158);
and U2013 (N_2013,N_1197,N_800);
or U2014 (N_2014,N_1095,N_832);
or U2015 (N_2015,N_933,N_1015);
or U2016 (N_2016,N_1210,N_1317);
xnor U2017 (N_2017,N_842,N_1269);
nand U2018 (N_2018,N_1043,N_947);
nor U2019 (N_2019,N_1179,N_896);
nand U2020 (N_2020,N_805,N_944);
or U2021 (N_2021,N_1488,N_1146);
and U2022 (N_2022,N_1117,N_1402);
xnor U2023 (N_2023,N_1042,N_953);
or U2024 (N_2024,N_1251,N_905);
nand U2025 (N_2025,N_1143,N_1362);
nor U2026 (N_2026,N_1217,N_1127);
or U2027 (N_2027,N_1297,N_1060);
or U2028 (N_2028,N_882,N_1305);
nor U2029 (N_2029,N_1486,N_1087);
and U2030 (N_2030,N_1164,N_808);
nand U2031 (N_2031,N_898,N_1144);
nor U2032 (N_2032,N_1092,N_1149);
nand U2033 (N_2033,N_1204,N_836);
or U2034 (N_2034,N_992,N_1135);
and U2035 (N_2035,N_754,N_1047);
and U2036 (N_2036,N_896,N_1233);
nand U2037 (N_2037,N_754,N_1384);
xnor U2038 (N_2038,N_1268,N_895);
or U2039 (N_2039,N_1007,N_1042);
xnor U2040 (N_2040,N_901,N_1370);
and U2041 (N_2041,N_1005,N_1189);
or U2042 (N_2042,N_1166,N_1250);
xor U2043 (N_2043,N_1082,N_796);
nand U2044 (N_2044,N_760,N_989);
nand U2045 (N_2045,N_1235,N_792);
or U2046 (N_2046,N_881,N_1369);
or U2047 (N_2047,N_1446,N_1259);
or U2048 (N_2048,N_1467,N_1101);
nor U2049 (N_2049,N_1362,N_868);
nand U2050 (N_2050,N_1449,N_1324);
nor U2051 (N_2051,N_1084,N_1311);
nor U2052 (N_2052,N_1023,N_1230);
xnor U2053 (N_2053,N_916,N_1390);
and U2054 (N_2054,N_1018,N_995);
and U2055 (N_2055,N_824,N_1128);
nor U2056 (N_2056,N_1278,N_1402);
nor U2057 (N_2057,N_833,N_1292);
nor U2058 (N_2058,N_1291,N_933);
or U2059 (N_2059,N_925,N_753);
xnor U2060 (N_2060,N_838,N_1411);
nand U2061 (N_2061,N_1284,N_1402);
and U2062 (N_2062,N_1266,N_1012);
nor U2063 (N_2063,N_909,N_849);
and U2064 (N_2064,N_1403,N_1214);
and U2065 (N_2065,N_1126,N_1208);
or U2066 (N_2066,N_1485,N_1303);
nand U2067 (N_2067,N_828,N_1499);
nand U2068 (N_2068,N_1299,N_1335);
nor U2069 (N_2069,N_1106,N_926);
and U2070 (N_2070,N_1410,N_1023);
and U2071 (N_2071,N_1018,N_1418);
nand U2072 (N_2072,N_981,N_937);
nor U2073 (N_2073,N_1396,N_817);
nand U2074 (N_2074,N_969,N_1365);
xnor U2075 (N_2075,N_893,N_1022);
nand U2076 (N_2076,N_895,N_848);
xor U2077 (N_2077,N_1236,N_861);
and U2078 (N_2078,N_1090,N_1322);
nor U2079 (N_2079,N_1286,N_1200);
nand U2080 (N_2080,N_1190,N_1067);
nor U2081 (N_2081,N_1255,N_1247);
nor U2082 (N_2082,N_1406,N_1285);
nand U2083 (N_2083,N_1157,N_1268);
nor U2084 (N_2084,N_1427,N_1366);
nand U2085 (N_2085,N_1012,N_1327);
or U2086 (N_2086,N_1239,N_1007);
and U2087 (N_2087,N_1051,N_1385);
xor U2088 (N_2088,N_984,N_781);
nor U2089 (N_2089,N_844,N_1473);
nor U2090 (N_2090,N_1456,N_1374);
nand U2091 (N_2091,N_1246,N_1094);
nand U2092 (N_2092,N_1445,N_1116);
or U2093 (N_2093,N_1283,N_794);
nand U2094 (N_2094,N_933,N_883);
nand U2095 (N_2095,N_941,N_1054);
nor U2096 (N_2096,N_862,N_1393);
or U2097 (N_2097,N_794,N_1077);
and U2098 (N_2098,N_1393,N_786);
nand U2099 (N_2099,N_1341,N_903);
and U2100 (N_2100,N_1169,N_1230);
nand U2101 (N_2101,N_1123,N_1055);
nand U2102 (N_2102,N_1166,N_1373);
nor U2103 (N_2103,N_1053,N_1274);
nand U2104 (N_2104,N_1031,N_1442);
and U2105 (N_2105,N_1097,N_821);
or U2106 (N_2106,N_1351,N_1118);
and U2107 (N_2107,N_1496,N_887);
nor U2108 (N_2108,N_1333,N_984);
nor U2109 (N_2109,N_1055,N_1256);
nand U2110 (N_2110,N_1346,N_1316);
nor U2111 (N_2111,N_774,N_1253);
nand U2112 (N_2112,N_1078,N_1495);
nand U2113 (N_2113,N_1084,N_1256);
nand U2114 (N_2114,N_1445,N_1193);
or U2115 (N_2115,N_1005,N_1263);
nand U2116 (N_2116,N_1035,N_793);
and U2117 (N_2117,N_1040,N_762);
nor U2118 (N_2118,N_1286,N_752);
nor U2119 (N_2119,N_1265,N_790);
or U2120 (N_2120,N_1422,N_979);
nand U2121 (N_2121,N_1431,N_1082);
or U2122 (N_2122,N_1336,N_1061);
or U2123 (N_2123,N_906,N_1107);
and U2124 (N_2124,N_761,N_1165);
nor U2125 (N_2125,N_991,N_1498);
or U2126 (N_2126,N_971,N_894);
and U2127 (N_2127,N_844,N_1319);
or U2128 (N_2128,N_838,N_1146);
and U2129 (N_2129,N_976,N_975);
or U2130 (N_2130,N_794,N_1263);
nand U2131 (N_2131,N_1472,N_1169);
xor U2132 (N_2132,N_832,N_1149);
nor U2133 (N_2133,N_832,N_811);
nand U2134 (N_2134,N_1383,N_1145);
nand U2135 (N_2135,N_811,N_1039);
nand U2136 (N_2136,N_1337,N_1421);
xor U2137 (N_2137,N_1436,N_1046);
xor U2138 (N_2138,N_1388,N_1115);
nand U2139 (N_2139,N_1267,N_1260);
and U2140 (N_2140,N_1173,N_1272);
and U2141 (N_2141,N_770,N_1423);
or U2142 (N_2142,N_1466,N_1422);
nand U2143 (N_2143,N_1293,N_1218);
or U2144 (N_2144,N_1229,N_1169);
nor U2145 (N_2145,N_1383,N_1311);
or U2146 (N_2146,N_864,N_1492);
nand U2147 (N_2147,N_1043,N_1181);
nor U2148 (N_2148,N_1189,N_762);
and U2149 (N_2149,N_1087,N_1276);
nor U2150 (N_2150,N_1370,N_1401);
xnor U2151 (N_2151,N_813,N_759);
xor U2152 (N_2152,N_937,N_1155);
nor U2153 (N_2153,N_814,N_943);
nor U2154 (N_2154,N_924,N_1169);
and U2155 (N_2155,N_1290,N_756);
nor U2156 (N_2156,N_1158,N_1055);
nor U2157 (N_2157,N_1338,N_1099);
or U2158 (N_2158,N_1181,N_1230);
nor U2159 (N_2159,N_877,N_1191);
or U2160 (N_2160,N_1283,N_1237);
and U2161 (N_2161,N_1053,N_916);
or U2162 (N_2162,N_960,N_924);
nand U2163 (N_2163,N_1470,N_1232);
nand U2164 (N_2164,N_932,N_1068);
nor U2165 (N_2165,N_904,N_1188);
nand U2166 (N_2166,N_1310,N_1376);
nand U2167 (N_2167,N_1314,N_786);
and U2168 (N_2168,N_945,N_899);
nand U2169 (N_2169,N_996,N_978);
nand U2170 (N_2170,N_1379,N_1109);
or U2171 (N_2171,N_1321,N_1108);
or U2172 (N_2172,N_982,N_1099);
nor U2173 (N_2173,N_1009,N_1407);
xnor U2174 (N_2174,N_1455,N_785);
xnor U2175 (N_2175,N_885,N_1197);
nor U2176 (N_2176,N_1461,N_1419);
nor U2177 (N_2177,N_794,N_832);
nor U2178 (N_2178,N_914,N_1409);
or U2179 (N_2179,N_1340,N_1191);
xnor U2180 (N_2180,N_1384,N_1204);
or U2181 (N_2181,N_1495,N_1064);
and U2182 (N_2182,N_1055,N_1085);
nor U2183 (N_2183,N_1084,N_878);
and U2184 (N_2184,N_1092,N_1258);
nand U2185 (N_2185,N_1262,N_818);
nand U2186 (N_2186,N_1395,N_914);
or U2187 (N_2187,N_801,N_1290);
nor U2188 (N_2188,N_928,N_833);
nand U2189 (N_2189,N_1268,N_939);
or U2190 (N_2190,N_1272,N_1103);
nor U2191 (N_2191,N_827,N_1233);
nand U2192 (N_2192,N_832,N_752);
nand U2193 (N_2193,N_1398,N_910);
nand U2194 (N_2194,N_1356,N_1151);
or U2195 (N_2195,N_917,N_1408);
or U2196 (N_2196,N_943,N_1444);
and U2197 (N_2197,N_940,N_1027);
nand U2198 (N_2198,N_1256,N_851);
nand U2199 (N_2199,N_1235,N_902);
nand U2200 (N_2200,N_1421,N_1280);
and U2201 (N_2201,N_1204,N_1005);
nand U2202 (N_2202,N_1395,N_1154);
nor U2203 (N_2203,N_1053,N_1449);
nand U2204 (N_2204,N_1017,N_1216);
nand U2205 (N_2205,N_951,N_1284);
or U2206 (N_2206,N_1003,N_915);
and U2207 (N_2207,N_750,N_1265);
nor U2208 (N_2208,N_1011,N_1037);
or U2209 (N_2209,N_1421,N_981);
nand U2210 (N_2210,N_1474,N_1013);
or U2211 (N_2211,N_1296,N_1279);
nor U2212 (N_2212,N_852,N_1245);
and U2213 (N_2213,N_927,N_1149);
nor U2214 (N_2214,N_1298,N_1343);
nor U2215 (N_2215,N_800,N_1249);
nand U2216 (N_2216,N_1189,N_1002);
nand U2217 (N_2217,N_1371,N_1266);
nand U2218 (N_2218,N_1021,N_917);
or U2219 (N_2219,N_1477,N_1495);
nor U2220 (N_2220,N_794,N_1238);
nand U2221 (N_2221,N_1354,N_1355);
and U2222 (N_2222,N_1300,N_1145);
or U2223 (N_2223,N_950,N_896);
or U2224 (N_2224,N_1257,N_983);
nand U2225 (N_2225,N_1057,N_1392);
or U2226 (N_2226,N_1213,N_947);
and U2227 (N_2227,N_922,N_1398);
and U2228 (N_2228,N_1379,N_1107);
nor U2229 (N_2229,N_1372,N_766);
and U2230 (N_2230,N_996,N_859);
nand U2231 (N_2231,N_1310,N_1481);
and U2232 (N_2232,N_793,N_1456);
xnor U2233 (N_2233,N_845,N_1383);
nor U2234 (N_2234,N_1023,N_809);
or U2235 (N_2235,N_1243,N_1205);
or U2236 (N_2236,N_862,N_1217);
or U2237 (N_2237,N_1006,N_978);
xor U2238 (N_2238,N_1177,N_1401);
nor U2239 (N_2239,N_1440,N_1254);
nand U2240 (N_2240,N_1183,N_1267);
nand U2241 (N_2241,N_801,N_1045);
or U2242 (N_2242,N_1244,N_795);
nor U2243 (N_2243,N_1425,N_1492);
xor U2244 (N_2244,N_921,N_1369);
nand U2245 (N_2245,N_1203,N_824);
xnor U2246 (N_2246,N_1479,N_930);
nand U2247 (N_2247,N_1199,N_1156);
and U2248 (N_2248,N_978,N_1253);
nand U2249 (N_2249,N_781,N_780);
or U2250 (N_2250,N_1651,N_1959);
xnor U2251 (N_2251,N_1980,N_1521);
nor U2252 (N_2252,N_2163,N_1695);
or U2253 (N_2253,N_2037,N_1592);
nor U2254 (N_2254,N_2109,N_1953);
or U2255 (N_2255,N_1863,N_1687);
and U2256 (N_2256,N_2117,N_1560);
nor U2257 (N_2257,N_1729,N_1799);
or U2258 (N_2258,N_1828,N_2173);
nand U2259 (N_2259,N_1827,N_1735);
and U2260 (N_2260,N_1787,N_2123);
and U2261 (N_2261,N_2116,N_1619);
or U2262 (N_2262,N_1842,N_2039);
and U2263 (N_2263,N_2023,N_1839);
and U2264 (N_2264,N_1565,N_1768);
nand U2265 (N_2265,N_1722,N_1831);
nor U2266 (N_2266,N_1769,N_1870);
nand U2267 (N_2267,N_1671,N_2158);
and U2268 (N_2268,N_2206,N_2111);
xor U2269 (N_2269,N_1856,N_1534);
nor U2270 (N_2270,N_1784,N_1541);
nand U2271 (N_2271,N_1869,N_1855);
or U2272 (N_2272,N_1589,N_2075);
or U2273 (N_2273,N_1653,N_1615);
nand U2274 (N_2274,N_1824,N_1758);
xor U2275 (N_2275,N_1810,N_2017);
xnor U2276 (N_2276,N_1938,N_1871);
and U2277 (N_2277,N_1701,N_2180);
or U2278 (N_2278,N_1976,N_2129);
nand U2279 (N_2279,N_2221,N_2024);
nand U2280 (N_2280,N_1952,N_1584);
or U2281 (N_2281,N_1508,N_2095);
or U2282 (N_2282,N_1984,N_1776);
and U2283 (N_2283,N_2190,N_2201);
or U2284 (N_2284,N_1928,N_1807);
or U2285 (N_2285,N_2072,N_2004);
nor U2286 (N_2286,N_1647,N_1524);
or U2287 (N_2287,N_1836,N_1595);
nor U2288 (N_2288,N_1689,N_2053);
and U2289 (N_2289,N_2038,N_1732);
and U2290 (N_2290,N_1992,N_1533);
or U2291 (N_2291,N_1755,N_1895);
or U2292 (N_2292,N_1585,N_1969);
and U2293 (N_2293,N_1756,N_2169);
and U2294 (N_2294,N_2167,N_2064);
nor U2295 (N_2295,N_2210,N_1819);
nand U2296 (N_2296,N_1929,N_1553);
nor U2297 (N_2297,N_1557,N_2226);
or U2298 (N_2298,N_1919,N_1935);
nor U2299 (N_2299,N_2199,N_1670);
or U2300 (N_2300,N_2026,N_1901);
nor U2301 (N_2301,N_2040,N_1883);
or U2302 (N_2302,N_1958,N_1593);
nor U2303 (N_2303,N_1598,N_2203);
or U2304 (N_2304,N_1973,N_1970);
nor U2305 (N_2305,N_1606,N_1994);
or U2306 (N_2306,N_2029,N_1632);
nor U2307 (N_2307,N_1679,N_1878);
or U2308 (N_2308,N_1536,N_1968);
nand U2309 (N_2309,N_2014,N_1607);
or U2310 (N_2310,N_1767,N_1682);
xnor U2311 (N_2311,N_2022,N_1946);
nor U2312 (N_2312,N_1520,N_1597);
and U2313 (N_2313,N_1507,N_1617);
or U2314 (N_2314,N_1932,N_1691);
xor U2315 (N_2315,N_1724,N_2178);
nor U2316 (N_2316,N_2225,N_1730);
and U2317 (N_2317,N_1900,N_1568);
xor U2318 (N_2318,N_2223,N_1849);
nor U2319 (N_2319,N_2013,N_1539);
or U2320 (N_2320,N_1550,N_2010);
nand U2321 (N_2321,N_1942,N_2165);
xnor U2322 (N_2322,N_2197,N_2103);
or U2323 (N_2323,N_1821,N_2020);
nand U2324 (N_2324,N_1795,N_1800);
nor U2325 (N_2325,N_1504,N_1741);
nor U2326 (N_2326,N_1841,N_2045);
nor U2327 (N_2327,N_1634,N_2241);
nand U2328 (N_2328,N_1678,N_1788);
nor U2329 (N_2329,N_1751,N_1727);
or U2330 (N_2330,N_1552,N_1752);
xor U2331 (N_2331,N_1840,N_1509);
and U2332 (N_2332,N_1979,N_2133);
and U2333 (N_2333,N_1638,N_2106);
xor U2334 (N_2334,N_2021,N_2157);
nand U2335 (N_2335,N_1914,N_1710);
nand U2336 (N_2336,N_2125,N_1746);
and U2337 (N_2337,N_2249,N_1889);
nor U2338 (N_2338,N_2036,N_1982);
xnor U2339 (N_2339,N_1618,N_1581);
and U2340 (N_2340,N_1657,N_2175);
nand U2341 (N_2341,N_1545,N_1714);
nor U2342 (N_2342,N_2148,N_2061);
nor U2343 (N_2343,N_1640,N_1720);
nor U2344 (N_2344,N_2142,N_1894);
nand U2345 (N_2345,N_2028,N_1542);
nand U2346 (N_2346,N_1853,N_1793);
or U2347 (N_2347,N_2149,N_1804);
and U2348 (N_2348,N_1556,N_2110);
or U2349 (N_2349,N_2016,N_1780);
nand U2350 (N_2350,N_1912,N_2008);
and U2351 (N_2351,N_1896,N_1728);
and U2352 (N_2352,N_1558,N_1674);
or U2353 (N_2353,N_2091,N_2235);
xnor U2354 (N_2354,N_2087,N_2236);
or U2355 (N_2355,N_2162,N_1676);
or U2356 (N_2356,N_1708,N_1566);
and U2357 (N_2357,N_1621,N_2208);
or U2358 (N_2358,N_2047,N_1846);
or U2359 (N_2359,N_1677,N_1660);
xor U2360 (N_2360,N_1759,N_2056);
nor U2361 (N_2361,N_1683,N_1988);
nand U2362 (N_2362,N_2219,N_2182);
nand U2363 (N_2363,N_1939,N_1622);
or U2364 (N_2364,N_1656,N_1705);
nand U2365 (N_2365,N_1884,N_2009);
nand U2366 (N_2366,N_1949,N_1512);
nor U2367 (N_2367,N_1610,N_2082);
nor U2368 (N_2368,N_2071,N_1789);
nor U2369 (N_2369,N_1662,N_1882);
nand U2370 (N_2370,N_2172,N_1774);
or U2371 (N_2371,N_1818,N_1986);
xor U2372 (N_2372,N_1835,N_2243);
nand U2373 (N_2373,N_1765,N_1697);
nand U2374 (N_2374,N_1590,N_2033);
nor U2375 (N_2375,N_2198,N_2239);
or U2376 (N_2376,N_1916,N_2151);
or U2377 (N_2377,N_1663,N_1899);
nand U2378 (N_2378,N_1950,N_2212);
and U2379 (N_2379,N_1685,N_1675);
or U2380 (N_2380,N_1829,N_1904);
nor U2381 (N_2381,N_1918,N_2060);
or U2382 (N_2382,N_1974,N_2119);
nor U2383 (N_2383,N_1530,N_1844);
nor U2384 (N_2384,N_1833,N_1599);
or U2385 (N_2385,N_2126,N_1813);
and U2386 (N_2386,N_1930,N_2144);
nand U2387 (N_2387,N_2193,N_1785);
nor U2388 (N_2388,N_2205,N_1718);
nand U2389 (N_2389,N_1514,N_1978);
or U2390 (N_2390,N_2011,N_2244);
nand U2391 (N_2391,N_2114,N_1587);
xor U2392 (N_2392,N_1888,N_2130);
nand U2393 (N_2393,N_2050,N_2231);
nor U2394 (N_2394,N_1713,N_1910);
or U2395 (N_2395,N_1612,N_1551);
or U2396 (N_2396,N_2000,N_2015);
xor U2397 (N_2397,N_1931,N_2120);
xor U2398 (N_2398,N_1965,N_1649);
and U2399 (N_2399,N_1602,N_1913);
nand U2400 (N_2400,N_2058,N_1731);
nor U2401 (N_2401,N_1519,N_1549);
nand U2402 (N_2402,N_2183,N_2030);
nand U2403 (N_2403,N_1905,N_1567);
nor U2404 (N_2404,N_1951,N_2138);
nor U2405 (N_2405,N_1594,N_1528);
nor U2406 (N_2406,N_1891,N_1754);
nand U2407 (N_2407,N_2143,N_1936);
or U2408 (N_2408,N_2032,N_1806);
nand U2409 (N_2409,N_1652,N_1583);
nand U2410 (N_2410,N_1921,N_2211);
xnor U2411 (N_2411,N_2090,N_1515);
or U2412 (N_2412,N_2153,N_1817);
and U2413 (N_2413,N_1977,N_2080);
nor U2414 (N_2414,N_1516,N_2139);
nor U2415 (N_2415,N_1502,N_1700);
xnor U2416 (N_2416,N_2077,N_1865);
and U2417 (N_2417,N_2248,N_2122);
and U2418 (N_2418,N_2222,N_1760);
nand U2419 (N_2419,N_1803,N_1911);
or U2420 (N_2420,N_1966,N_1559);
and U2421 (N_2421,N_1538,N_2207);
or U2422 (N_2422,N_1748,N_1673);
nor U2423 (N_2423,N_1954,N_2066);
nand U2424 (N_2424,N_1802,N_1847);
nor U2425 (N_2425,N_2127,N_1537);
and U2426 (N_2426,N_2229,N_1922);
and U2427 (N_2427,N_1555,N_2228);
nor U2428 (N_2428,N_1535,N_1838);
and U2429 (N_2429,N_2048,N_1843);
nand U2430 (N_2430,N_1991,N_1624);
and U2431 (N_2431,N_1655,N_1503);
or U2432 (N_2432,N_1642,N_2107);
and U2433 (N_2433,N_1650,N_1775);
nor U2434 (N_2434,N_1805,N_1646);
nand U2435 (N_2435,N_1955,N_1906);
or U2436 (N_2436,N_2078,N_1811);
nor U2437 (N_2437,N_1540,N_2131);
nand U2438 (N_2438,N_1860,N_1639);
xor U2439 (N_2439,N_2186,N_1750);
and U2440 (N_2440,N_2135,N_1517);
or U2441 (N_2441,N_2217,N_2192);
and U2442 (N_2442,N_1688,N_1690);
nand U2443 (N_2443,N_1572,N_1845);
or U2444 (N_2444,N_2108,N_2220);
nand U2445 (N_2445,N_2202,N_1588);
and U2446 (N_2446,N_1511,N_2044);
and U2447 (N_2447,N_2073,N_1825);
and U2448 (N_2448,N_2034,N_1814);
and U2449 (N_2449,N_1961,N_1770);
or U2450 (N_2450,N_1791,N_2046);
nor U2451 (N_2451,N_2164,N_1993);
and U2452 (N_2452,N_1763,N_1726);
or U2453 (N_2453,N_1664,N_1715);
nand U2454 (N_2454,N_1893,N_1880);
nor U2455 (N_2455,N_1609,N_1658);
nand U2456 (N_2456,N_1945,N_1852);
or U2457 (N_2457,N_1987,N_1696);
nand U2458 (N_2458,N_1586,N_2132);
or U2459 (N_2459,N_2240,N_1591);
nor U2460 (N_2460,N_2184,N_1518);
nand U2461 (N_2461,N_1500,N_1578);
xor U2462 (N_2462,N_2200,N_2003);
or U2463 (N_2463,N_1563,N_1749);
nor U2464 (N_2464,N_1531,N_1872);
nor U2465 (N_2465,N_1779,N_1794);
or U2466 (N_2466,N_1686,N_2237);
nand U2467 (N_2467,N_1908,N_1757);
and U2468 (N_2468,N_2213,N_1554);
and U2469 (N_2469,N_2019,N_2096);
nor U2470 (N_2470,N_1781,N_1698);
and U2471 (N_2471,N_1620,N_1734);
nor U2472 (N_2472,N_2089,N_2067);
nor U2473 (N_2473,N_2059,N_1740);
and U2474 (N_2474,N_1628,N_1564);
or U2475 (N_2475,N_2156,N_1867);
and U2476 (N_2476,N_1873,N_2227);
nor U2477 (N_2477,N_2042,N_2031);
nor U2478 (N_2478,N_1739,N_2238);
or U2479 (N_2479,N_1963,N_1772);
or U2480 (N_2480,N_1857,N_1903);
nand U2481 (N_2481,N_2025,N_1926);
xnor U2482 (N_2482,N_2115,N_2145);
and U2483 (N_2483,N_1861,N_1995);
nand U2484 (N_2484,N_2191,N_2194);
xor U2485 (N_2485,N_1964,N_2188);
nand U2486 (N_2486,N_1522,N_1637);
or U2487 (N_2487,N_1577,N_1782);
xor U2488 (N_2488,N_1762,N_2242);
nand U2489 (N_2489,N_1956,N_1771);
and U2490 (N_2490,N_1877,N_2214);
nand U2491 (N_2491,N_2035,N_1645);
and U2492 (N_2492,N_1672,N_2176);
xnor U2493 (N_2493,N_1601,N_1796);
and U2494 (N_2494,N_1625,N_1773);
and U2495 (N_2495,N_2185,N_1943);
nor U2496 (N_2496,N_1742,N_1854);
or U2497 (N_2497,N_1989,N_1786);
nor U2498 (N_2498,N_1631,N_1834);
and U2499 (N_2499,N_1764,N_1874);
xnor U2500 (N_2500,N_1902,N_1630);
nand U2501 (N_2501,N_2121,N_2204);
xnor U2502 (N_2502,N_1546,N_1527);
nand U2503 (N_2503,N_2189,N_2088);
nand U2504 (N_2504,N_1526,N_1736);
and U2505 (N_2505,N_1699,N_1915);
and U2506 (N_2506,N_2136,N_1960);
and U2507 (N_2507,N_1702,N_1830);
or U2508 (N_2508,N_1603,N_2068);
nor U2509 (N_2509,N_1934,N_2166);
nor U2510 (N_2510,N_2170,N_1801);
and U2511 (N_2511,N_1909,N_1711);
nand U2512 (N_2512,N_2152,N_1626);
or U2513 (N_2513,N_1745,N_1571);
xnor U2514 (N_2514,N_2002,N_1669);
and U2515 (N_2515,N_1641,N_1957);
or U2516 (N_2516,N_1820,N_1850);
nor U2517 (N_2517,N_2027,N_1999);
and U2518 (N_2518,N_2150,N_1614);
or U2519 (N_2519,N_1665,N_2093);
and U2520 (N_2520,N_1975,N_2146);
xor U2521 (N_2521,N_2018,N_2112);
nand U2522 (N_2522,N_1937,N_1738);
nand U2523 (N_2523,N_2099,N_1629);
nor U2524 (N_2524,N_1823,N_1998);
nand U2525 (N_2525,N_1666,N_2196);
nor U2526 (N_2526,N_1707,N_2195);
nor U2527 (N_2527,N_1579,N_2159);
nand U2528 (N_2528,N_2006,N_1815);
xor U2529 (N_2529,N_2094,N_1744);
nand U2530 (N_2530,N_1562,N_1897);
nor U2531 (N_2531,N_1737,N_1887);
nand U2532 (N_2532,N_1920,N_1643);
nor U2533 (N_2533,N_1709,N_1668);
nor U2534 (N_2534,N_2001,N_2083);
nand U2535 (N_2535,N_2085,N_2179);
or U2536 (N_2536,N_1627,N_1575);
xor U2537 (N_2537,N_1616,N_1721);
or U2538 (N_2538,N_2104,N_2154);
nor U2539 (N_2539,N_1885,N_2070);
and U2540 (N_2540,N_1792,N_1809);
xor U2541 (N_2541,N_1967,N_1654);
nand U2542 (N_2542,N_1747,N_2100);
xnor U2543 (N_2543,N_1543,N_1693);
or U2544 (N_2544,N_1766,N_2069);
and U2545 (N_2545,N_2174,N_2181);
nand U2546 (N_2546,N_1611,N_1723);
or U2547 (N_2547,N_2012,N_1866);
or U2548 (N_2548,N_1608,N_2076);
and U2549 (N_2549,N_1600,N_2074);
and U2550 (N_2550,N_1983,N_2216);
nand U2551 (N_2551,N_1875,N_1703);
and U2552 (N_2552,N_1862,N_1777);
or U2553 (N_2553,N_1941,N_2218);
or U2554 (N_2554,N_1525,N_1694);
and U2555 (N_2555,N_1851,N_1925);
and U2556 (N_2556,N_1681,N_2043);
nand U2557 (N_2557,N_1890,N_2049);
or U2558 (N_2558,N_1990,N_1981);
or U2559 (N_2559,N_1570,N_2247);
xor U2560 (N_2560,N_1644,N_2168);
and U2561 (N_2561,N_2052,N_2007);
or U2562 (N_2562,N_2215,N_2224);
xor U2563 (N_2563,N_1633,N_1948);
nor U2564 (N_2564,N_2234,N_1706);
xor U2565 (N_2565,N_1907,N_1661);
or U2566 (N_2566,N_2054,N_1501);
or U2567 (N_2567,N_1924,N_1725);
xnor U2568 (N_2568,N_2246,N_1790);
and U2569 (N_2569,N_1881,N_2118);
and U2570 (N_2570,N_1927,N_1944);
xnor U2571 (N_2571,N_2209,N_2057);
nand U2572 (N_2572,N_1996,N_2141);
nand U2573 (N_2573,N_1864,N_1797);
nor U2574 (N_2574,N_1574,N_1761);
and U2575 (N_2575,N_1783,N_2134);
and U2576 (N_2576,N_2187,N_1604);
and U2577 (N_2577,N_1532,N_1547);
and U2578 (N_2578,N_1648,N_2177);
or U2579 (N_2579,N_1837,N_2055);
or U2580 (N_2580,N_1623,N_1513);
or U2581 (N_2581,N_2041,N_1997);
nor U2582 (N_2582,N_2128,N_2155);
nand U2583 (N_2583,N_1635,N_1778);
nand U2584 (N_2584,N_2245,N_1712);
xor U2585 (N_2585,N_1596,N_2140);
or U2586 (N_2586,N_2101,N_1933);
xor U2587 (N_2587,N_1985,N_2124);
and U2588 (N_2588,N_1506,N_1972);
and U2589 (N_2589,N_1962,N_1798);
nand U2590 (N_2590,N_1548,N_2065);
nand U2591 (N_2591,N_1659,N_1529);
and U2592 (N_2592,N_2092,N_2232);
nor U2593 (N_2593,N_1733,N_2105);
nor U2594 (N_2594,N_2161,N_2051);
nand U2595 (N_2595,N_1858,N_1605);
and U2596 (N_2596,N_2063,N_1582);
xnor U2597 (N_2597,N_1580,N_1717);
or U2598 (N_2598,N_1680,N_2230);
and U2599 (N_2599,N_1753,N_1573);
and U2600 (N_2600,N_1848,N_1505);
nand U2601 (N_2601,N_2160,N_1923);
xnor U2602 (N_2602,N_1886,N_1808);
and U2603 (N_2603,N_1971,N_2147);
xor U2604 (N_2604,N_1743,N_1719);
or U2605 (N_2605,N_2113,N_2097);
nor U2606 (N_2606,N_1613,N_2137);
nor U2607 (N_2607,N_2098,N_2005);
nor U2608 (N_2608,N_1667,N_1859);
nor U2609 (N_2609,N_1832,N_1947);
and U2610 (N_2610,N_1561,N_2084);
and U2611 (N_2611,N_1684,N_1917);
nor U2612 (N_2612,N_1636,N_1812);
and U2613 (N_2613,N_1704,N_2102);
and U2614 (N_2614,N_1892,N_1879);
and U2615 (N_2615,N_2233,N_1544);
xnor U2616 (N_2616,N_1692,N_1576);
nand U2617 (N_2617,N_1876,N_1826);
or U2618 (N_2618,N_1898,N_2171);
and U2619 (N_2619,N_2062,N_1510);
and U2620 (N_2620,N_1868,N_1816);
and U2621 (N_2621,N_1716,N_2086);
and U2622 (N_2622,N_1822,N_1940);
nor U2623 (N_2623,N_1569,N_2079);
and U2624 (N_2624,N_1523,N_2081);
nor U2625 (N_2625,N_2096,N_1835);
and U2626 (N_2626,N_1734,N_2158);
nor U2627 (N_2627,N_1740,N_2227);
nand U2628 (N_2628,N_2006,N_1989);
and U2629 (N_2629,N_1610,N_2199);
or U2630 (N_2630,N_2111,N_2032);
or U2631 (N_2631,N_1879,N_1813);
nand U2632 (N_2632,N_1956,N_1739);
nor U2633 (N_2633,N_1542,N_1635);
nand U2634 (N_2634,N_2171,N_2153);
nand U2635 (N_2635,N_1780,N_2088);
xnor U2636 (N_2636,N_1931,N_1729);
xnor U2637 (N_2637,N_2144,N_1997);
xnor U2638 (N_2638,N_1951,N_1673);
xor U2639 (N_2639,N_1725,N_1680);
nand U2640 (N_2640,N_1621,N_1820);
nor U2641 (N_2641,N_1830,N_1974);
or U2642 (N_2642,N_1521,N_1755);
and U2643 (N_2643,N_1823,N_1667);
or U2644 (N_2644,N_1711,N_2114);
and U2645 (N_2645,N_1500,N_2170);
nor U2646 (N_2646,N_2242,N_1512);
or U2647 (N_2647,N_1996,N_1791);
and U2648 (N_2648,N_2062,N_1922);
nand U2649 (N_2649,N_1804,N_1959);
and U2650 (N_2650,N_1551,N_2088);
nand U2651 (N_2651,N_2200,N_1897);
nor U2652 (N_2652,N_1751,N_1810);
and U2653 (N_2653,N_2156,N_1522);
or U2654 (N_2654,N_1797,N_1838);
and U2655 (N_2655,N_1776,N_1955);
nor U2656 (N_2656,N_1605,N_1534);
and U2657 (N_2657,N_1576,N_1930);
nand U2658 (N_2658,N_1727,N_1710);
nor U2659 (N_2659,N_2128,N_1896);
nand U2660 (N_2660,N_1549,N_2075);
nor U2661 (N_2661,N_1702,N_1694);
or U2662 (N_2662,N_2149,N_2006);
or U2663 (N_2663,N_1968,N_2009);
nand U2664 (N_2664,N_1904,N_2163);
and U2665 (N_2665,N_2141,N_1835);
nand U2666 (N_2666,N_1702,N_2049);
xnor U2667 (N_2667,N_2025,N_1934);
and U2668 (N_2668,N_1619,N_1838);
nand U2669 (N_2669,N_1745,N_1724);
nand U2670 (N_2670,N_1856,N_1736);
nand U2671 (N_2671,N_1530,N_1924);
and U2672 (N_2672,N_1839,N_1608);
and U2673 (N_2673,N_1712,N_2071);
and U2674 (N_2674,N_1872,N_1880);
xnor U2675 (N_2675,N_1506,N_1542);
xor U2676 (N_2676,N_1579,N_1760);
nand U2677 (N_2677,N_2057,N_1603);
or U2678 (N_2678,N_2197,N_1654);
or U2679 (N_2679,N_1556,N_1605);
nand U2680 (N_2680,N_1890,N_1579);
nor U2681 (N_2681,N_2235,N_1695);
or U2682 (N_2682,N_2153,N_2150);
or U2683 (N_2683,N_2077,N_1738);
nand U2684 (N_2684,N_2195,N_1981);
nor U2685 (N_2685,N_1763,N_2034);
and U2686 (N_2686,N_2027,N_2093);
nor U2687 (N_2687,N_1874,N_1618);
and U2688 (N_2688,N_1740,N_1929);
nand U2689 (N_2689,N_1962,N_1796);
and U2690 (N_2690,N_1540,N_1961);
nor U2691 (N_2691,N_1561,N_1735);
nor U2692 (N_2692,N_2228,N_1933);
xnor U2693 (N_2693,N_1622,N_1584);
and U2694 (N_2694,N_1900,N_1736);
xor U2695 (N_2695,N_2208,N_1973);
nor U2696 (N_2696,N_1905,N_1984);
nor U2697 (N_2697,N_1762,N_1517);
and U2698 (N_2698,N_1576,N_1590);
or U2699 (N_2699,N_2100,N_1628);
nor U2700 (N_2700,N_1517,N_1858);
and U2701 (N_2701,N_1901,N_1681);
nand U2702 (N_2702,N_1940,N_1894);
or U2703 (N_2703,N_2006,N_1702);
nor U2704 (N_2704,N_2077,N_2105);
nand U2705 (N_2705,N_1574,N_2027);
nand U2706 (N_2706,N_2147,N_2195);
and U2707 (N_2707,N_1770,N_2127);
and U2708 (N_2708,N_2193,N_1835);
xor U2709 (N_2709,N_2082,N_1666);
nor U2710 (N_2710,N_2025,N_1919);
nor U2711 (N_2711,N_1508,N_1689);
xor U2712 (N_2712,N_2031,N_2130);
or U2713 (N_2713,N_1974,N_2028);
nand U2714 (N_2714,N_2051,N_1749);
and U2715 (N_2715,N_1756,N_2132);
nand U2716 (N_2716,N_2136,N_1828);
xor U2717 (N_2717,N_1843,N_2149);
and U2718 (N_2718,N_2123,N_2193);
nor U2719 (N_2719,N_2029,N_1584);
or U2720 (N_2720,N_1799,N_2222);
nand U2721 (N_2721,N_1757,N_1958);
and U2722 (N_2722,N_1980,N_1900);
xnor U2723 (N_2723,N_1815,N_2066);
or U2724 (N_2724,N_1598,N_2235);
and U2725 (N_2725,N_1609,N_1966);
xnor U2726 (N_2726,N_1589,N_1957);
nor U2727 (N_2727,N_2231,N_1515);
and U2728 (N_2728,N_1534,N_1541);
and U2729 (N_2729,N_2109,N_1684);
nor U2730 (N_2730,N_2110,N_1504);
or U2731 (N_2731,N_1852,N_1766);
or U2732 (N_2732,N_1504,N_2224);
nand U2733 (N_2733,N_2016,N_1756);
and U2734 (N_2734,N_1773,N_2245);
or U2735 (N_2735,N_1873,N_1682);
or U2736 (N_2736,N_2106,N_1764);
nor U2737 (N_2737,N_2129,N_1844);
and U2738 (N_2738,N_1867,N_1544);
nand U2739 (N_2739,N_2078,N_1545);
or U2740 (N_2740,N_1605,N_2164);
and U2741 (N_2741,N_1847,N_1707);
and U2742 (N_2742,N_1500,N_1553);
or U2743 (N_2743,N_1582,N_1636);
and U2744 (N_2744,N_2134,N_1924);
nor U2745 (N_2745,N_1788,N_1997);
and U2746 (N_2746,N_1520,N_1549);
nor U2747 (N_2747,N_1538,N_1722);
nand U2748 (N_2748,N_1555,N_1831);
nor U2749 (N_2749,N_1775,N_1968);
nand U2750 (N_2750,N_1546,N_1622);
xor U2751 (N_2751,N_1972,N_1626);
and U2752 (N_2752,N_1775,N_1601);
and U2753 (N_2753,N_2144,N_2016);
or U2754 (N_2754,N_2083,N_1919);
xnor U2755 (N_2755,N_1686,N_1991);
and U2756 (N_2756,N_2113,N_1613);
or U2757 (N_2757,N_1584,N_2070);
nand U2758 (N_2758,N_1659,N_1861);
nand U2759 (N_2759,N_1602,N_1593);
nor U2760 (N_2760,N_1729,N_2208);
and U2761 (N_2761,N_1527,N_2098);
and U2762 (N_2762,N_2227,N_1515);
nand U2763 (N_2763,N_1529,N_2233);
and U2764 (N_2764,N_1638,N_1764);
xnor U2765 (N_2765,N_2021,N_1923);
or U2766 (N_2766,N_2110,N_2087);
nand U2767 (N_2767,N_1989,N_2015);
nor U2768 (N_2768,N_1998,N_2190);
and U2769 (N_2769,N_2085,N_1886);
nand U2770 (N_2770,N_1826,N_1865);
nor U2771 (N_2771,N_1553,N_1831);
nand U2772 (N_2772,N_2147,N_1507);
nand U2773 (N_2773,N_2022,N_1656);
or U2774 (N_2774,N_1521,N_2182);
nand U2775 (N_2775,N_1562,N_2198);
nand U2776 (N_2776,N_1612,N_1729);
or U2777 (N_2777,N_1534,N_2134);
and U2778 (N_2778,N_2154,N_1670);
nand U2779 (N_2779,N_1903,N_1821);
and U2780 (N_2780,N_2059,N_1667);
xor U2781 (N_2781,N_2153,N_1518);
nand U2782 (N_2782,N_1603,N_2195);
nand U2783 (N_2783,N_2057,N_2234);
or U2784 (N_2784,N_1513,N_1521);
and U2785 (N_2785,N_1906,N_2122);
and U2786 (N_2786,N_2217,N_1841);
or U2787 (N_2787,N_1917,N_1744);
nor U2788 (N_2788,N_1800,N_1916);
and U2789 (N_2789,N_2043,N_1822);
nor U2790 (N_2790,N_1527,N_2168);
and U2791 (N_2791,N_1575,N_1866);
nand U2792 (N_2792,N_1794,N_2036);
or U2793 (N_2793,N_2195,N_1525);
nand U2794 (N_2794,N_2101,N_2149);
nand U2795 (N_2795,N_1985,N_1714);
nand U2796 (N_2796,N_2162,N_1689);
and U2797 (N_2797,N_1649,N_1986);
and U2798 (N_2798,N_1524,N_1892);
or U2799 (N_2799,N_1825,N_2240);
and U2800 (N_2800,N_1996,N_1780);
or U2801 (N_2801,N_2000,N_2098);
nand U2802 (N_2802,N_2146,N_1554);
nor U2803 (N_2803,N_2095,N_1676);
nor U2804 (N_2804,N_1616,N_2047);
nand U2805 (N_2805,N_1550,N_1724);
and U2806 (N_2806,N_2068,N_1555);
and U2807 (N_2807,N_1705,N_1917);
nor U2808 (N_2808,N_2105,N_1874);
nor U2809 (N_2809,N_1673,N_1823);
nand U2810 (N_2810,N_1786,N_2174);
or U2811 (N_2811,N_1579,N_2182);
or U2812 (N_2812,N_1946,N_1777);
nand U2813 (N_2813,N_1608,N_1944);
nand U2814 (N_2814,N_1952,N_1757);
nand U2815 (N_2815,N_2080,N_2137);
or U2816 (N_2816,N_1949,N_1596);
nor U2817 (N_2817,N_1717,N_2128);
nand U2818 (N_2818,N_1788,N_1504);
and U2819 (N_2819,N_1528,N_2019);
nor U2820 (N_2820,N_1806,N_1810);
nor U2821 (N_2821,N_1767,N_2077);
nor U2822 (N_2822,N_1810,N_1714);
and U2823 (N_2823,N_1585,N_2156);
nor U2824 (N_2824,N_1586,N_1717);
nand U2825 (N_2825,N_2203,N_1621);
and U2826 (N_2826,N_2192,N_1997);
and U2827 (N_2827,N_2036,N_1665);
nor U2828 (N_2828,N_1896,N_1702);
nor U2829 (N_2829,N_1861,N_1919);
nor U2830 (N_2830,N_2042,N_1700);
and U2831 (N_2831,N_1821,N_1795);
or U2832 (N_2832,N_1715,N_1876);
nor U2833 (N_2833,N_2096,N_1547);
or U2834 (N_2834,N_1983,N_2193);
nor U2835 (N_2835,N_1577,N_1594);
nand U2836 (N_2836,N_1882,N_2176);
nand U2837 (N_2837,N_1966,N_1706);
xnor U2838 (N_2838,N_1886,N_2198);
xnor U2839 (N_2839,N_2102,N_1591);
nor U2840 (N_2840,N_2098,N_1990);
nand U2841 (N_2841,N_1607,N_1947);
nor U2842 (N_2842,N_1602,N_2081);
or U2843 (N_2843,N_1614,N_1541);
xnor U2844 (N_2844,N_1825,N_1554);
nand U2845 (N_2845,N_2215,N_1753);
xor U2846 (N_2846,N_1693,N_2013);
or U2847 (N_2847,N_2130,N_1756);
nor U2848 (N_2848,N_1522,N_2164);
nand U2849 (N_2849,N_2211,N_1562);
nand U2850 (N_2850,N_1861,N_2017);
nand U2851 (N_2851,N_1559,N_2018);
and U2852 (N_2852,N_1794,N_1636);
xnor U2853 (N_2853,N_2139,N_2028);
nand U2854 (N_2854,N_1596,N_1644);
and U2855 (N_2855,N_2088,N_1767);
nor U2856 (N_2856,N_2176,N_1828);
and U2857 (N_2857,N_1720,N_2228);
xnor U2858 (N_2858,N_1614,N_1709);
xor U2859 (N_2859,N_1962,N_2128);
nor U2860 (N_2860,N_1538,N_1509);
nor U2861 (N_2861,N_2166,N_1798);
xnor U2862 (N_2862,N_2229,N_1864);
nand U2863 (N_2863,N_2074,N_2080);
nor U2864 (N_2864,N_2122,N_2128);
nand U2865 (N_2865,N_1992,N_1704);
nor U2866 (N_2866,N_1638,N_1886);
nor U2867 (N_2867,N_2027,N_1587);
or U2868 (N_2868,N_1782,N_1705);
nand U2869 (N_2869,N_2065,N_1780);
nand U2870 (N_2870,N_1773,N_1750);
nand U2871 (N_2871,N_2132,N_1751);
xnor U2872 (N_2872,N_1826,N_1568);
xor U2873 (N_2873,N_2105,N_1566);
nand U2874 (N_2874,N_2082,N_2023);
nand U2875 (N_2875,N_1564,N_2029);
or U2876 (N_2876,N_1857,N_2180);
and U2877 (N_2877,N_1625,N_1654);
and U2878 (N_2878,N_1867,N_2237);
or U2879 (N_2879,N_1865,N_1811);
nand U2880 (N_2880,N_2182,N_1924);
or U2881 (N_2881,N_2132,N_1520);
or U2882 (N_2882,N_1773,N_1859);
nor U2883 (N_2883,N_1697,N_1565);
xor U2884 (N_2884,N_2043,N_1725);
nor U2885 (N_2885,N_2166,N_2225);
or U2886 (N_2886,N_1654,N_1619);
nor U2887 (N_2887,N_2148,N_1752);
nor U2888 (N_2888,N_2157,N_1946);
nand U2889 (N_2889,N_1595,N_1884);
nand U2890 (N_2890,N_1988,N_1534);
or U2891 (N_2891,N_1679,N_2194);
xor U2892 (N_2892,N_1843,N_2058);
or U2893 (N_2893,N_1726,N_1529);
or U2894 (N_2894,N_2222,N_1966);
or U2895 (N_2895,N_1818,N_1876);
nand U2896 (N_2896,N_2067,N_2035);
and U2897 (N_2897,N_2011,N_1842);
and U2898 (N_2898,N_1738,N_1948);
nand U2899 (N_2899,N_1838,N_1874);
nand U2900 (N_2900,N_1527,N_1839);
nand U2901 (N_2901,N_1616,N_2240);
nor U2902 (N_2902,N_1776,N_1856);
nand U2903 (N_2903,N_2200,N_2229);
nand U2904 (N_2904,N_1906,N_1932);
or U2905 (N_2905,N_2096,N_1534);
xnor U2906 (N_2906,N_1861,N_2234);
nand U2907 (N_2907,N_2100,N_1539);
xor U2908 (N_2908,N_1544,N_1814);
or U2909 (N_2909,N_1916,N_1901);
and U2910 (N_2910,N_1819,N_1802);
or U2911 (N_2911,N_1803,N_2017);
and U2912 (N_2912,N_2069,N_2082);
or U2913 (N_2913,N_2040,N_1833);
or U2914 (N_2914,N_2101,N_2224);
and U2915 (N_2915,N_2017,N_2135);
or U2916 (N_2916,N_2248,N_2040);
nand U2917 (N_2917,N_1729,N_1981);
and U2918 (N_2918,N_1792,N_2006);
nor U2919 (N_2919,N_1546,N_1829);
nor U2920 (N_2920,N_2236,N_1684);
or U2921 (N_2921,N_1875,N_1960);
and U2922 (N_2922,N_1687,N_1633);
or U2923 (N_2923,N_1631,N_1816);
and U2924 (N_2924,N_2031,N_2210);
nor U2925 (N_2925,N_2160,N_1506);
nor U2926 (N_2926,N_1724,N_1860);
or U2927 (N_2927,N_1519,N_1769);
xnor U2928 (N_2928,N_1533,N_1694);
nand U2929 (N_2929,N_2075,N_1681);
nor U2930 (N_2930,N_2052,N_2087);
or U2931 (N_2931,N_1854,N_1903);
nor U2932 (N_2932,N_1804,N_1773);
or U2933 (N_2933,N_1770,N_2181);
nand U2934 (N_2934,N_1794,N_2175);
nand U2935 (N_2935,N_2039,N_2195);
and U2936 (N_2936,N_1845,N_2211);
and U2937 (N_2937,N_1931,N_2041);
or U2938 (N_2938,N_2009,N_2033);
nand U2939 (N_2939,N_1737,N_1687);
xor U2940 (N_2940,N_1968,N_1674);
nor U2941 (N_2941,N_2104,N_1958);
and U2942 (N_2942,N_1517,N_1664);
nor U2943 (N_2943,N_2180,N_2220);
nor U2944 (N_2944,N_1603,N_1841);
nor U2945 (N_2945,N_2129,N_1631);
nor U2946 (N_2946,N_2136,N_1652);
nor U2947 (N_2947,N_1692,N_1776);
and U2948 (N_2948,N_2038,N_1685);
and U2949 (N_2949,N_2172,N_1594);
nor U2950 (N_2950,N_1875,N_1557);
nand U2951 (N_2951,N_1551,N_1877);
nor U2952 (N_2952,N_1925,N_1920);
nand U2953 (N_2953,N_1814,N_2245);
xnor U2954 (N_2954,N_1931,N_1821);
or U2955 (N_2955,N_1840,N_1776);
nand U2956 (N_2956,N_1890,N_2192);
nand U2957 (N_2957,N_2218,N_1746);
nor U2958 (N_2958,N_2045,N_1864);
nand U2959 (N_2959,N_1928,N_2197);
nand U2960 (N_2960,N_1550,N_2061);
nor U2961 (N_2961,N_1841,N_1561);
or U2962 (N_2962,N_1943,N_1863);
nor U2963 (N_2963,N_1965,N_1580);
or U2964 (N_2964,N_1719,N_2212);
nor U2965 (N_2965,N_2199,N_2212);
nor U2966 (N_2966,N_1625,N_1610);
or U2967 (N_2967,N_1874,N_1603);
xnor U2968 (N_2968,N_1573,N_2175);
and U2969 (N_2969,N_2241,N_2178);
nand U2970 (N_2970,N_2229,N_1822);
or U2971 (N_2971,N_2246,N_1983);
xnor U2972 (N_2972,N_1806,N_1521);
or U2973 (N_2973,N_2156,N_1931);
xor U2974 (N_2974,N_1848,N_1678);
nand U2975 (N_2975,N_1741,N_1945);
nand U2976 (N_2976,N_2249,N_1751);
or U2977 (N_2977,N_2028,N_1678);
nand U2978 (N_2978,N_1780,N_1852);
and U2979 (N_2979,N_1539,N_2209);
or U2980 (N_2980,N_1857,N_1745);
xor U2981 (N_2981,N_1796,N_2171);
or U2982 (N_2982,N_1761,N_2232);
or U2983 (N_2983,N_1973,N_2227);
nor U2984 (N_2984,N_2198,N_2141);
nor U2985 (N_2985,N_2096,N_1561);
nor U2986 (N_2986,N_2058,N_2032);
and U2987 (N_2987,N_1619,N_1855);
or U2988 (N_2988,N_1633,N_1983);
nand U2989 (N_2989,N_2181,N_1511);
or U2990 (N_2990,N_1595,N_1598);
nor U2991 (N_2991,N_2050,N_1980);
nand U2992 (N_2992,N_1693,N_1964);
and U2993 (N_2993,N_2225,N_1678);
and U2994 (N_2994,N_2072,N_1777);
nand U2995 (N_2995,N_2214,N_1691);
and U2996 (N_2996,N_1785,N_2246);
or U2997 (N_2997,N_1808,N_1529);
nand U2998 (N_2998,N_1558,N_1611);
nand U2999 (N_2999,N_1510,N_2093);
nand UO_0 (O_0,N_2360,N_2743);
or UO_1 (O_1,N_2261,N_2418);
nor UO_2 (O_2,N_2751,N_2706);
and UO_3 (O_3,N_2495,N_2972);
nor UO_4 (O_4,N_2799,N_2894);
nand UO_5 (O_5,N_2762,N_2359);
xnor UO_6 (O_6,N_2756,N_2338);
and UO_7 (O_7,N_2708,N_2624);
nand UO_8 (O_8,N_2333,N_2672);
or UO_9 (O_9,N_2876,N_2608);
nand UO_10 (O_10,N_2330,N_2365);
or UO_11 (O_11,N_2677,N_2473);
nor UO_12 (O_12,N_2993,N_2652);
and UO_13 (O_13,N_2783,N_2325);
xnor UO_14 (O_14,N_2545,N_2503);
nand UO_15 (O_15,N_2324,N_2619);
nor UO_16 (O_16,N_2782,N_2784);
and UO_17 (O_17,N_2479,N_2753);
and UO_18 (O_18,N_2502,N_2494);
xnor UO_19 (O_19,N_2583,N_2530);
or UO_20 (O_20,N_2485,N_2565);
and UO_21 (O_21,N_2881,N_2446);
nand UO_22 (O_22,N_2486,N_2880);
nor UO_23 (O_23,N_2658,N_2251);
or UO_24 (O_24,N_2424,N_2576);
nor UO_25 (O_25,N_2728,N_2432);
and UO_26 (O_26,N_2308,N_2686);
and UO_27 (O_27,N_2295,N_2529);
nand UO_28 (O_28,N_2269,N_2638);
xnor UO_29 (O_29,N_2488,N_2430);
or UO_30 (O_30,N_2331,N_2605);
xor UO_31 (O_31,N_2755,N_2604);
xnor UO_32 (O_32,N_2673,N_2824);
nor UO_33 (O_33,N_2433,N_2662);
nand UO_34 (O_34,N_2777,N_2719);
and UO_35 (O_35,N_2519,N_2265);
and UO_36 (O_36,N_2748,N_2566);
or UO_37 (O_37,N_2795,N_2747);
nand UO_38 (O_38,N_2811,N_2959);
nand UO_39 (O_39,N_2855,N_2457);
nor UO_40 (O_40,N_2538,N_2685);
nor UO_41 (O_41,N_2438,N_2864);
nand UO_42 (O_42,N_2944,N_2649);
nor UO_43 (O_43,N_2459,N_2885);
nor UO_44 (O_44,N_2882,N_2287);
nor UO_45 (O_45,N_2981,N_2584);
nand UO_46 (O_46,N_2366,N_2839);
nand UO_47 (O_47,N_2384,N_2901);
and UO_48 (O_48,N_2840,N_2847);
nand UO_49 (O_49,N_2536,N_2588);
nand UO_50 (O_50,N_2443,N_2328);
nand UO_51 (O_51,N_2773,N_2460);
xnor UO_52 (O_52,N_2992,N_2377);
or UO_53 (O_53,N_2913,N_2655);
nor UO_54 (O_54,N_2822,N_2956);
nand UO_55 (O_55,N_2760,N_2872);
and UO_56 (O_56,N_2732,N_2408);
nor UO_57 (O_57,N_2970,N_2752);
or UO_58 (O_58,N_2998,N_2600);
or UO_59 (O_59,N_2742,N_2806);
nand UO_60 (O_60,N_2848,N_2632);
or UO_61 (O_61,N_2978,N_2267);
nand UO_62 (O_62,N_2317,N_2785);
and UO_63 (O_63,N_2830,N_2578);
nand UO_64 (O_64,N_2506,N_2634);
nor UO_65 (O_65,N_2362,N_2767);
nor UO_66 (O_66,N_2447,N_2387);
xor UO_67 (O_67,N_2699,N_2793);
nor UO_68 (O_68,N_2965,N_2818);
xor UO_69 (O_69,N_2252,N_2590);
nor UO_70 (O_70,N_2698,N_2680);
or UO_71 (O_71,N_2994,N_2513);
xnor UO_72 (O_72,N_2976,N_2693);
and UO_73 (O_73,N_2772,N_2311);
and UO_74 (O_74,N_2664,N_2466);
nand UO_75 (O_75,N_2585,N_2304);
nand UO_76 (O_76,N_2392,N_2904);
nor UO_77 (O_77,N_2544,N_2532);
or UO_78 (O_78,N_2442,N_2665);
nor UO_79 (O_79,N_2531,N_2819);
nor UO_80 (O_80,N_2758,N_2735);
xnor UO_81 (O_81,N_2650,N_2514);
nor UO_82 (O_82,N_2471,N_2508);
xnor UO_83 (O_83,N_2713,N_2381);
xor UO_84 (O_84,N_2862,N_2598);
nand UO_85 (O_85,N_2809,N_2716);
nand UO_86 (O_86,N_2254,N_2854);
nor UO_87 (O_87,N_2835,N_2397);
nor UO_88 (O_88,N_2937,N_2451);
and UO_89 (O_89,N_2358,N_2852);
nor UO_90 (O_90,N_2474,N_2524);
nor UO_91 (O_91,N_2946,N_2846);
or UO_92 (O_92,N_2765,N_2552);
or UO_93 (O_93,N_2285,N_2733);
nand UO_94 (O_94,N_2947,N_2964);
and UO_95 (O_95,N_2884,N_2292);
xor UO_96 (O_96,N_2606,N_2329);
xnor UO_97 (O_97,N_2450,N_2300);
nand UO_98 (O_98,N_2492,N_2873);
nor UO_99 (O_99,N_2663,N_2468);
or UO_100 (O_100,N_2682,N_2476);
or UO_101 (O_101,N_2501,N_2929);
nand UO_102 (O_102,N_2429,N_2568);
or UO_103 (O_103,N_2428,N_2660);
or UO_104 (O_104,N_2775,N_2934);
nand UO_105 (O_105,N_2412,N_2581);
xor UO_106 (O_106,N_2382,N_2940);
nand UO_107 (O_107,N_2286,N_2942);
or UO_108 (O_108,N_2787,N_2572);
and UO_109 (O_109,N_2990,N_2390);
or UO_110 (O_110,N_2487,N_2774);
or UO_111 (O_111,N_2518,N_2439);
or UO_112 (O_112,N_2816,N_2737);
nor UO_113 (O_113,N_2941,N_2813);
nor UO_114 (O_114,N_2607,N_2781);
xor UO_115 (O_115,N_2435,N_2293);
or UO_116 (O_116,N_2919,N_2420);
nand UO_117 (O_117,N_2354,N_2776);
and UO_118 (O_118,N_2410,N_2391);
and UO_119 (O_119,N_2804,N_2422);
and UO_120 (O_120,N_2689,N_2550);
and UO_121 (O_121,N_2385,N_2794);
or UO_122 (O_122,N_2915,N_2925);
and UO_123 (O_123,N_2761,N_2749);
and UO_124 (O_124,N_2388,N_2995);
or UO_125 (O_125,N_2419,N_2654);
nand UO_126 (O_126,N_2551,N_2714);
or UO_127 (O_127,N_2613,N_2979);
nor UO_128 (O_128,N_2938,N_2865);
nor UO_129 (O_129,N_2403,N_2296);
nand UO_130 (O_130,N_2564,N_2715);
nand UO_131 (O_131,N_2323,N_2879);
xor UO_132 (O_132,N_2920,N_2736);
or UO_133 (O_133,N_2386,N_2861);
or UO_134 (O_134,N_2945,N_2641);
and UO_135 (O_135,N_2691,N_2534);
nor UO_136 (O_136,N_2724,N_2630);
nand UO_137 (O_137,N_2356,N_2790);
nor UO_138 (O_138,N_2657,N_2318);
nand UO_139 (O_139,N_2725,N_2260);
or UO_140 (O_140,N_2368,N_2490);
xnor UO_141 (O_141,N_2951,N_2668);
or UO_142 (O_142,N_2599,N_2376);
xor UO_143 (O_143,N_2643,N_2969);
and UO_144 (O_144,N_2593,N_2561);
or UO_145 (O_145,N_2504,N_2288);
xnor UO_146 (O_146,N_2887,N_2859);
or UO_147 (O_147,N_2294,N_2922);
and UO_148 (O_148,N_2573,N_2921);
nor UO_149 (O_149,N_2797,N_2321);
or UO_150 (O_150,N_2319,N_2505);
or UO_151 (O_151,N_2923,N_2631);
nor UO_152 (O_152,N_2924,N_2526);
nor UO_153 (O_153,N_2842,N_2274);
or UO_154 (O_154,N_2931,N_2834);
nor UO_155 (O_155,N_2414,N_2263);
nor UO_156 (O_156,N_2905,N_2950);
and UO_157 (O_157,N_2477,N_2349);
nand UO_158 (O_158,N_2759,N_2290);
or UO_159 (O_159,N_2582,N_2374);
xnor UO_160 (O_160,N_2344,N_2498);
nor UO_161 (O_161,N_2579,N_2256);
and UO_162 (O_162,N_2509,N_2789);
or UO_163 (O_163,N_2301,N_2763);
xor UO_164 (O_164,N_2647,N_2516);
and UO_165 (O_165,N_2997,N_2826);
nand UO_166 (O_166,N_2908,N_2255);
nor UO_167 (O_167,N_2702,N_2710);
nand UO_168 (O_168,N_2455,N_2394);
nor UO_169 (O_169,N_2327,N_2957);
or UO_170 (O_170,N_2404,N_2609);
xnor UO_171 (O_171,N_2423,N_2540);
and UO_172 (O_172,N_2820,N_2461);
or UO_173 (O_173,N_2770,N_2268);
or UO_174 (O_174,N_2731,N_2548);
nand UO_175 (O_175,N_2895,N_2335);
and UO_176 (O_176,N_2483,N_2316);
or UO_177 (O_177,N_2517,N_2723);
or UO_178 (O_178,N_2684,N_2636);
nand UO_179 (O_179,N_2875,N_2543);
nand UO_180 (O_180,N_2987,N_2306);
or UO_181 (O_181,N_2798,N_2871);
and UO_182 (O_182,N_2371,N_2346);
or UO_183 (O_183,N_2900,N_2802);
and UO_184 (O_184,N_2982,N_2918);
nor UO_185 (O_185,N_2720,N_2928);
or UO_186 (O_186,N_2744,N_2332);
nand UO_187 (O_187,N_2322,N_2603);
and UO_188 (O_188,N_2930,N_2627);
or UO_189 (O_189,N_2955,N_2838);
or UO_190 (O_190,N_2963,N_2337);
or UO_191 (O_191,N_2464,N_2690);
nand UO_192 (O_192,N_2659,N_2717);
or UO_193 (O_193,N_2284,N_2860);
or UO_194 (O_194,N_2899,N_2431);
nor UO_195 (O_195,N_2546,N_2870);
nand UO_196 (O_196,N_2779,N_2766);
nor UO_197 (O_197,N_2857,N_2264);
and UO_198 (O_198,N_2314,N_2482);
nor UO_199 (O_199,N_2623,N_2470);
nand UO_200 (O_200,N_2746,N_2741);
xnor UO_201 (O_201,N_2910,N_2511);
xnor UO_202 (O_202,N_2449,N_2484);
nor UO_203 (O_203,N_2851,N_2591);
xnor UO_204 (O_204,N_2270,N_2537);
and UO_205 (O_205,N_2771,N_2694);
nor UO_206 (O_206,N_2253,N_2812);
nand UO_207 (O_207,N_2628,N_2909);
nor UO_208 (O_208,N_2258,N_2985);
or UO_209 (O_209,N_2521,N_2289);
and UO_210 (O_210,N_2415,N_2615);
nand UO_211 (O_211,N_2273,N_2475);
xor UO_212 (O_212,N_2640,N_2364);
or UO_213 (O_213,N_2307,N_2696);
or UO_214 (O_214,N_2991,N_2954);
nor UO_215 (O_215,N_2528,N_2653);
or UO_216 (O_216,N_2357,N_2850);
xnor UO_217 (O_217,N_2817,N_2786);
or UO_218 (O_218,N_2396,N_2952);
or UO_219 (O_219,N_2574,N_2988);
xor UO_220 (O_220,N_2712,N_2888);
nor UO_221 (O_221,N_2436,N_2278);
and UO_222 (O_222,N_2497,N_2589);
nand UO_223 (O_223,N_2629,N_2553);
and UO_224 (O_224,N_2315,N_2395);
nor UO_225 (O_225,N_2409,N_2932);
nand UO_226 (O_226,N_2869,N_2535);
nand UO_227 (O_227,N_2305,N_2935);
and UO_228 (O_228,N_2845,N_2454);
or UO_229 (O_229,N_2916,N_2788);
and UO_230 (O_230,N_2626,N_2562);
or UO_231 (O_231,N_2592,N_2507);
nor UO_232 (O_232,N_2764,N_2378);
nor UO_233 (O_233,N_2701,N_2907);
nor UO_234 (O_234,N_2823,N_2389);
nor UO_235 (O_235,N_2821,N_2625);
and UO_236 (O_236,N_2276,N_2676);
and UO_237 (O_237,N_2989,N_2542);
nor UO_238 (O_238,N_2815,N_2343);
or UO_239 (O_239,N_2666,N_2527);
nor UO_240 (O_240,N_2730,N_2577);
and UO_241 (O_241,N_2961,N_2596);
xor UO_242 (O_242,N_2645,N_2983);
nor UO_243 (O_243,N_2411,N_2383);
nand UO_244 (O_244,N_2996,N_2718);
and UO_245 (O_245,N_2275,N_2575);
xnor UO_246 (O_246,N_2547,N_2791);
and UO_247 (O_247,N_2858,N_2405);
and UO_248 (O_248,N_2656,N_2734);
nor UO_249 (O_249,N_2441,N_2635);
and UO_250 (O_250,N_2739,N_2571);
xnor UO_251 (O_251,N_2711,N_2469);
and UO_252 (O_252,N_2943,N_2310);
and UO_253 (O_253,N_2340,N_2803);
nor UO_254 (O_254,N_2974,N_2370);
and UO_255 (O_255,N_2646,N_2320);
nor UO_256 (O_256,N_2351,N_2448);
nand UO_257 (O_257,N_2611,N_2303);
nor UO_258 (O_258,N_2539,N_2651);
nand UO_259 (O_259,N_2525,N_2369);
and UO_260 (O_260,N_2695,N_2481);
nand UO_261 (O_261,N_2727,N_2678);
and UO_262 (O_262,N_2707,N_2363);
xor UO_263 (O_263,N_2867,N_2927);
nand UO_264 (O_264,N_2644,N_2836);
nand UO_265 (O_265,N_2282,N_2939);
or UO_266 (O_266,N_2480,N_2949);
nand UO_267 (O_267,N_2810,N_2266);
nand UO_268 (O_268,N_2444,N_2309);
and UO_269 (O_269,N_2704,N_2299);
xor UO_270 (O_270,N_2999,N_2866);
xor UO_271 (O_271,N_2661,N_2675);
or UO_272 (O_272,N_2407,N_2612);
nor UO_273 (O_273,N_2958,N_2906);
or UO_274 (O_274,N_2953,N_2533);
xor UO_275 (O_275,N_2973,N_2688);
or UO_276 (O_276,N_2515,N_2828);
xnor UO_277 (O_277,N_2971,N_2768);
xor UO_278 (O_278,N_2903,N_2347);
nor UO_279 (O_279,N_2610,N_2496);
nor UO_280 (O_280,N_2681,N_2355);
or UO_281 (O_281,N_2462,N_2421);
nand UO_282 (O_282,N_2456,N_2738);
nand UO_283 (O_283,N_2595,N_2345);
xnor UO_284 (O_284,N_2637,N_2825);
nor UO_285 (O_285,N_2336,N_2399);
or UO_286 (O_286,N_2570,N_2980);
nand UO_287 (O_287,N_2769,N_2620);
nand UO_288 (O_288,N_2780,N_2298);
nand UO_289 (O_289,N_2843,N_2440);
nand UO_290 (O_290,N_2878,N_2745);
or UO_291 (O_291,N_2465,N_2792);
xor UO_292 (O_292,N_2372,N_2499);
nand UO_293 (O_293,N_2297,N_2671);
nand UO_294 (O_294,N_2554,N_2601);
xor UO_295 (O_295,N_2902,N_2452);
nor UO_296 (O_296,N_2703,N_2962);
or UO_297 (O_297,N_2425,N_2281);
and UO_298 (O_298,N_2523,N_2401);
xnor UO_299 (O_299,N_2975,N_2912);
nand UO_300 (O_300,N_2594,N_2679);
nor UO_301 (O_301,N_2968,N_2639);
and UO_302 (O_302,N_2379,N_2402);
nand UO_303 (O_303,N_2709,N_2367);
nand UO_304 (O_304,N_2478,N_2966);
nor UO_305 (O_305,N_2986,N_2416);
xnor UO_306 (O_306,N_2602,N_2729);
nand UO_307 (O_307,N_2796,N_2896);
and UO_308 (O_308,N_2353,N_2334);
or UO_309 (O_309,N_2580,N_2726);
nand UO_310 (O_310,N_2807,N_2493);
or UO_311 (O_311,N_2642,N_2341);
xnor UO_312 (O_312,N_2348,N_2563);
nand UO_313 (O_313,N_2597,N_2890);
nor UO_314 (O_314,N_2467,N_2827);
nand UO_315 (O_315,N_2326,N_2617);
xor UO_316 (O_316,N_2250,N_2559);
and UO_317 (O_317,N_2437,N_2960);
nor UO_318 (O_318,N_2936,N_2808);
and UO_319 (O_319,N_2831,N_2555);
and UO_320 (O_320,N_2380,N_2445);
nor UO_321 (O_321,N_2863,N_2697);
nand UO_322 (O_322,N_2683,N_2841);
nand UO_323 (O_323,N_2754,N_2914);
nor UO_324 (O_324,N_2648,N_2883);
nand UO_325 (O_325,N_2977,N_2687);
nand UO_326 (O_326,N_2853,N_2614);
nand UO_327 (O_327,N_2586,N_2417);
nor UO_328 (O_328,N_2622,N_2453);
and UO_329 (O_329,N_2874,N_2560);
xor UO_330 (O_330,N_2283,N_2587);
nand UO_331 (O_331,N_2814,N_2434);
nand UO_332 (O_332,N_2279,N_2621);
nand UO_333 (O_333,N_2801,N_2721);
nor UO_334 (O_334,N_2398,N_2373);
nand UO_335 (O_335,N_2271,N_2911);
xor UO_336 (O_336,N_2800,N_2257);
and UO_337 (O_337,N_2413,N_2350);
nand UO_338 (O_338,N_2280,N_2569);
or UO_339 (O_339,N_2491,N_2926);
nand UO_340 (O_340,N_2891,N_2692);
nor UO_341 (O_341,N_2557,N_2272);
nor UO_342 (O_342,N_2618,N_2361);
or UO_343 (O_343,N_2674,N_2262);
and UO_344 (O_344,N_2556,N_2633);
xnor UO_345 (O_345,N_2849,N_2705);
xnor UO_346 (O_346,N_2520,N_2757);
xor UO_347 (O_347,N_2549,N_2700);
nor UO_348 (O_348,N_2277,N_2669);
or UO_349 (O_349,N_2500,N_2897);
nor UO_350 (O_350,N_2670,N_2458);
or UO_351 (O_351,N_2892,N_2837);
nand UO_352 (O_352,N_2868,N_2406);
nand UO_353 (O_353,N_2886,N_2375);
or UO_354 (O_354,N_2510,N_2948);
nor UO_355 (O_355,N_2567,N_2489);
xor UO_356 (O_356,N_2722,N_2558);
nor UO_357 (O_357,N_2259,N_2302);
nor UO_358 (O_358,N_2832,N_2393);
or UO_359 (O_359,N_2541,N_2339);
nand UO_360 (O_360,N_2898,N_2917);
or UO_361 (O_361,N_2805,N_2312);
and UO_362 (O_362,N_2463,N_2844);
or UO_363 (O_363,N_2400,N_2967);
nor UO_364 (O_364,N_2984,N_2616);
nand UO_365 (O_365,N_2426,N_2512);
nand UO_366 (O_366,N_2522,N_2933);
and UO_367 (O_367,N_2291,N_2778);
or UO_368 (O_368,N_2893,N_2833);
or UO_369 (O_369,N_2472,N_2427);
or UO_370 (O_370,N_2829,N_2856);
and UO_371 (O_371,N_2889,N_2667);
or UO_372 (O_372,N_2342,N_2740);
or UO_373 (O_373,N_2750,N_2352);
or UO_374 (O_374,N_2313,N_2877);
or UO_375 (O_375,N_2397,N_2765);
nor UO_376 (O_376,N_2542,N_2517);
nor UO_377 (O_377,N_2669,N_2691);
and UO_378 (O_378,N_2541,N_2493);
and UO_379 (O_379,N_2480,N_2823);
or UO_380 (O_380,N_2421,N_2638);
nand UO_381 (O_381,N_2309,N_2760);
nor UO_382 (O_382,N_2266,N_2809);
nor UO_383 (O_383,N_2340,N_2679);
nor UO_384 (O_384,N_2662,N_2925);
nor UO_385 (O_385,N_2410,N_2539);
nand UO_386 (O_386,N_2925,N_2871);
nand UO_387 (O_387,N_2497,N_2436);
and UO_388 (O_388,N_2582,N_2418);
nor UO_389 (O_389,N_2747,N_2278);
xor UO_390 (O_390,N_2487,N_2604);
or UO_391 (O_391,N_2700,N_2677);
or UO_392 (O_392,N_2534,N_2427);
or UO_393 (O_393,N_2907,N_2290);
and UO_394 (O_394,N_2822,N_2282);
and UO_395 (O_395,N_2358,N_2570);
and UO_396 (O_396,N_2859,N_2295);
xnor UO_397 (O_397,N_2304,N_2591);
or UO_398 (O_398,N_2488,N_2307);
nor UO_399 (O_399,N_2628,N_2479);
nand UO_400 (O_400,N_2372,N_2948);
and UO_401 (O_401,N_2846,N_2622);
and UO_402 (O_402,N_2353,N_2421);
or UO_403 (O_403,N_2629,N_2509);
or UO_404 (O_404,N_2488,N_2738);
nor UO_405 (O_405,N_2443,N_2367);
nor UO_406 (O_406,N_2981,N_2498);
nand UO_407 (O_407,N_2468,N_2507);
nor UO_408 (O_408,N_2428,N_2285);
nand UO_409 (O_409,N_2259,N_2945);
xnor UO_410 (O_410,N_2840,N_2926);
nor UO_411 (O_411,N_2655,N_2504);
or UO_412 (O_412,N_2830,N_2428);
and UO_413 (O_413,N_2563,N_2257);
or UO_414 (O_414,N_2647,N_2428);
or UO_415 (O_415,N_2339,N_2535);
nor UO_416 (O_416,N_2449,N_2687);
nor UO_417 (O_417,N_2710,N_2546);
and UO_418 (O_418,N_2419,N_2628);
nor UO_419 (O_419,N_2394,N_2520);
and UO_420 (O_420,N_2763,N_2611);
or UO_421 (O_421,N_2389,N_2977);
xor UO_422 (O_422,N_2922,N_2329);
nand UO_423 (O_423,N_2631,N_2670);
and UO_424 (O_424,N_2933,N_2334);
or UO_425 (O_425,N_2554,N_2308);
and UO_426 (O_426,N_2298,N_2803);
nand UO_427 (O_427,N_2310,N_2680);
nor UO_428 (O_428,N_2836,N_2463);
nand UO_429 (O_429,N_2398,N_2907);
nand UO_430 (O_430,N_2953,N_2524);
and UO_431 (O_431,N_2790,N_2688);
nor UO_432 (O_432,N_2352,N_2873);
xor UO_433 (O_433,N_2607,N_2710);
nand UO_434 (O_434,N_2886,N_2663);
nand UO_435 (O_435,N_2647,N_2937);
or UO_436 (O_436,N_2877,N_2995);
and UO_437 (O_437,N_2400,N_2542);
nor UO_438 (O_438,N_2326,N_2707);
nand UO_439 (O_439,N_2879,N_2641);
nor UO_440 (O_440,N_2329,N_2776);
xor UO_441 (O_441,N_2341,N_2314);
nor UO_442 (O_442,N_2817,N_2494);
or UO_443 (O_443,N_2400,N_2935);
nor UO_444 (O_444,N_2919,N_2715);
or UO_445 (O_445,N_2833,N_2313);
or UO_446 (O_446,N_2928,N_2684);
and UO_447 (O_447,N_2589,N_2727);
or UO_448 (O_448,N_2389,N_2526);
xnor UO_449 (O_449,N_2293,N_2583);
or UO_450 (O_450,N_2917,N_2621);
nand UO_451 (O_451,N_2254,N_2635);
nor UO_452 (O_452,N_2945,N_2726);
nor UO_453 (O_453,N_2396,N_2661);
and UO_454 (O_454,N_2440,N_2324);
nand UO_455 (O_455,N_2781,N_2383);
nand UO_456 (O_456,N_2908,N_2645);
and UO_457 (O_457,N_2451,N_2624);
and UO_458 (O_458,N_2254,N_2917);
or UO_459 (O_459,N_2329,N_2699);
or UO_460 (O_460,N_2500,N_2367);
nand UO_461 (O_461,N_2417,N_2871);
xor UO_462 (O_462,N_2293,N_2912);
or UO_463 (O_463,N_2949,N_2527);
nand UO_464 (O_464,N_2761,N_2933);
and UO_465 (O_465,N_2954,N_2405);
or UO_466 (O_466,N_2271,N_2671);
and UO_467 (O_467,N_2263,N_2642);
xnor UO_468 (O_468,N_2423,N_2690);
xnor UO_469 (O_469,N_2619,N_2794);
xor UO_470 (O_470,N_2808,N_2881);
nor UO_471 (O_471,N_2335,N_2308);
nand UO_472 (O_472,N_2647,N_2294);
nor UO_473 (O_473,N_2595,N_2359);
xor UO_474 (O_474,N_2854,N_2260);
and UO_475 (O_475,N_2287,N_2656);
or UO_476 (O_476,N_2347,N_2922);
xor UO_477 (O_477,N_2291,N_2724);
and UO_478 (O_478,N_2380,N_2758);
and UO_479 (O_479,N_2525,N_2407);
and UO_480 (O_480,N_2963,N_2761);
and UO_481 (O_481,N_2704,N_2421);
xnor UO_482 (O_482,N_2376,N_2277);
and UO_483 (O_483,N_2694,N_2799);
or UO_484 (O_484,N_2302,N_2601);
xor UO_485 (O_485,N_2542,N_2996);
nand UO_486 (O_486,N_2812,N_2335);
nor UO_487 (O_487,N_2300,N_2504);
or UO_488 (O_488,N_2595,N_2385);
and UO_489 (O_489,N_2298,N_2790);
or UO_490 (O_490,N_2974,N_2482);
nor UO_491 (O_491,N_2729,N_2293);
xor UO_492 (O_492,N_2801,N_2791);
or UO_493 (O_493,N_2544,N_2832);
or UO_494 (O_494,N_2328,N_2696);
or UO_495 (O_495,N_2726,N_2308);
xor UO_496 (O_496,N_2507,N_2947);
nand UO_497 (O_497,N_2873,N_2857);
nand UO_498 (O_498,N_2697,N_2995);
or UO_499 (O_499,N_2614,N_2522);
endmodule