module basic_500_3000_500_40_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_20,In_399);
and U1 (N_1,In_371,In_406);
nor U2 (N_2,In_263,In_90);
and U3 (N_3,In_13,In_264);
nor U4 (N_4,In_292,In_176);
nand U5 (N_5,In_380,In_425);
or U6 (N_6,In_312,In_342);
nor U7 (N_7,In_415,In_246);
and U8 (N_8,In_44,In_16);
nor U9 (N_9,In_444,In_430);
nor U10 (N_10,In_142,In_321);
xnor U11 (N_11,In_141,In_488);
nand U12 (N_12,In_148,In_432);
nand U13 (N_13,In_319,In_139);
xnor U14 (N_14,In_201,In_78);
or U15 (N_15,In_58,In_125);
and U16 (N_16,In_205,In_39);
or U17 (N_17,In_405,In_452);
xnor U18 (N_18,In_393,In_93);
nand U19 (N_19,In_208,In_314);
nand U20 (N_20,In_287,In_269);
xor U21 (N_21,In_57,In_127);
nor U22 (N_22,In_85,In_333);
nand U23 (N_23,In_449,In_423);
and U24 (N_24,In_222,In_219);
and U25 (N_25,In_402,In_99);
xnor U26 (N_26,In_355,In_153);
nand U27 (N_27,In_110,In_72);
or U28 (N_28,In_128,In_495);
xnor U29 (N_29,In_416,In_42);
nand U30 (N_30,In_181,In_216);
or U31 (N_31,In_56,In_112);
nand U32 (N_32,In_420,In_129);
and U33 (N_33,In_440,In_175);
nand U34 (N_34,In_28,In_316);
and U35 (N_35,In_29,In_436);
and U36 (N_36,In_100,In_298);
nor U37 (N_37,In_51,In_340);
xnor U38 (N_38,In_255,In_372);
nand U39 (N_39,In_41,In_233);
nand U40 (N_40,In_31,In_185);
and U41 (N_41,In_102,In_61);
nand U42 (N_42,In_464,In_326);
and U43 (N_43,In_207,In_266);
nor U44 (N_44,In_352,In_244);
and U45 (N_45,In_52,In_190);
nor U46 (N_46,In_426,In_170);
or U47 (N_47,In_294,In_45);
nor U48 (N_48,In_336,In_360);
or U49 (N_49,In_383,In_482);
nor U50 (N_50,In_435,In_22);
nor U51 (N_51,In_304,In_247);
nand U52 (N_52,In_50,In_103);
or U53 (N_53,In_136,In_106);
xnor U54 (N_54,In_4,In_53);
and U55 (N_55,In_446,In_450);
nand U56 (N_56,In_81,In_456);
xor U57 (N_57,In_356,In_282);
or U58 (N_58,In_289,In_487);
xnor U59 (N_59,In_6,In_178);
nor U60 (N_60,In_492,In_10);
xnor U61 (N_61,In_252,In_318);
nand U62 (N_62,In_109,In_241);
nor U63 (N_63,In_69,In_334);
xor U64 (N_64,In_145,In_479);
or U65 (N_65,In_218,In_92);
or U66 (N_66,In_468,In_21);
and U67 (N_67,In_150,In_83);
and U68 (N_68,In_418,In_443);
or U69 (N_69,In_410,In_79);
nand U70 (N_70,In_431,In_82);
xor U71 (N_71,In_439,In_121);
nor U72 (N_72,In_173,In_283);
and U73 (N_73,In_163,In_350);
nand U74 (N_74,In_303,In_276);
nor U75 (N_75,In_398,In_413);
and U76 (N_76,In_260,In_80);
xor U77 (N_77,In_373,In_235);
nor U78 (N_78,In_273,In_249);
or U79 (N_79,In_367,N_5);
and U80 (N_80,In_293,In_137);
and U81 (N_81,In_461,In_354);
nor U82 (N_82,In_242,In_95);
nand U83 (N_83,In_167,In_89);
nor U84 (N_84,In_258,In_169);
nand U85 (N_85,In_328,In_284);
xor U86 (N_86,In_23,In_183);
xor U87 (N_87,In_458,In_338);
nor U88 (N_88,In_113,N_60);
nand U89 (N_89,N_6,In_400);
or U90 (N_90,N_65,In_97);
nor U91 (N_91,In_147,In_359);
xnor U92 (N_92,N_14,N_0);
xnor U93 (N_93,In_265,In_476);
nand U94 (N_94,In_392,In_25);
or U95 (N_95,N_47,In_301);
xor U96 (N_96,N_72,In_346);
or U97 (N_97,In_119,In_236);
and U98 (N_98,In_451,N_4);
nand U99 (N_99,In_317,N_44);
xor U100 (N_100,In_489,N_18);
nand U101 (N_101,In_256,In_162);
and U102 (N_102,In_203,In_475);
and U103 (N_103,In_254,In_391);
and U104 (N_104,N_31,In_38);
nor U105 (N_105,In_417,In_123);
xnor U106 (N_106,In_124,In_310);
xor U107 (N_107,In_409,In_240);
and U108 (N_108,In_389,N_48);
or U109 (N_109,In_463,In_427);
nor U110 (N_110,In_49,In_313);
xnor U111 (N_111,N_39,In_447);
nand U112 (N_112,In_174,In_114);
and U113 (N_113,In_243,In_323);
xor U114 (N_114,In_480,In_473);
and U115 (N_115,N_36,N_35);
xnor U116 (N_116,In_362,In_324);
nor U117 (N_117,In_157,In_126);
xor U118 (N_118,N_24,In_143);
or U119 (N_119,In_344,In_101);
nand U120 (N_120,In_130,In_198);
and U121 (N_121,N_52,In_281);
or U122 (N_122,In_34,In_9);
or U123 (N_123,In_172,In_343);
nand U124 (N_124,In_339,In_193);
nor U125 (N_125,In_345,N_67);
or U126 (N_126,In_15,In_378);
or U127 (N_127,In_168,In_442);
or U128 (N_128,In_382,In_47);
and U129 (N_129,In_108,N_32);
nor U130 (N_130,In_248,In_472);
or U131 (N_131,In_98,In_295);
and U132 (N_132,In_33,In_306);
or U133 (N_133,In_151,In_88);
nand U134 (N_134,In_498,In_197);
xor U135 (N_135,In_74,In_275);
and U136 (N_136,N_56,In_94);
and U137 (N_137,In_3,In_84);
xor U138 (N_138,In_166,N_42);
and U139 (N_139,In_225,In_171);
or U140 (N_140,In_335,In_404);
xor U141 (N_141,N_29,In_285);
nand U142 (N_142,In_186,In_421);
nor U143 (N_143,In_238,In_348);
or U144 (N_144,In_386,In_154);
and U145 (N_145,In_55,In_374);
xor U146 (N_146,In_351,In_192);
nand U147 (N_147,In_327,In_332);
or U148 (N_148,In_361,N_49);
xor U149 (N_149,In_111,In_204);
nor U150 (N_150,N_143,N_103);
nor U151 (N_151,In_0,N_137);
and U152 (N_152,In_407,In_159);
xor U153 (N_153,In_272,In_457);
nand U154 (N_154,In_363,In_459);
nor U155 (N_155,In_239,In_140);
xor U156 (N_156,In_146,N_45);
xnor U157 (N_157,In_471,N_22);
nand U158 (N_158,N_130,N_11);
nor U159 (N_159,N_108,In_376);
or U160 (N_160,In_470,In_364);
or U161 (N_161,N_135,In_104);
xor U162 (N_162,N_126,N_140);
or U163 (N_163,N_77,N_97);
nor U164 (N_164,In_118,In_337);
or U165 (N_165,N_71,In_395);
xor U166 (N_166,In_271,In_237);
nand U167 (N_167,In_64,N_20);
nand U168 (N_168,In_215,In_230);
xnor U169 (N_169,N_85,In_202);
or U170 (N_170,In_408,In_330);
nand U171 (N_171,In_434,In_465);
xnor U172 (N_172,N_59,N_98);
nor U173 (N_173,In_368,N_12);
or U174 (N_174,In_220,In_76);
and U175 (N_175,In_296,In_499);
xor U176 (N_176,In_474,N_63);
or U177 (N_177,In_331,In_394);
and U178 (N_178,In_358,In_221);
nor U179 (N_179,N_61,N_142);
xor U180 (N_180,N_62,In_422);
and U181 (N_181,N_121,In_182);
xor U182 (N_182,N_120,In_187);
xor U183 (N_183,In_309,In_462);
xnor U184 (N_184,N_131,In_429);
nor U185 (N_185,N_128,N_1);
nor U186 (N_186,N_53,In_370);
nor U187 (N_187,N_84,In_412);
nand U188 (N_188,In_36,N_87);
nor U189 (N_189,In_477,N_148);
or U190 (N_190,In_86,In_48);
nand U191 (N_191,In_274,N_115);
or U192 (N_192,In_188,N_93);
or U193 (N_193,In_305,In_419);
nor U194 (N_194,In_60,N_2);
xor U195 (N_195,In_300,In_67);
nand U196 (N_196,N_43,In_17);
nand U197 (N_197,In_453,In_12);
xor U198 (N_198,In_2,N_78);
xnor U199 (N_199,In_245,In_26);
or U200 (N_200,In_325,In_68);
nor U201 (N_201,N_92,In_8);
nor U202 (N_202,N_25,In_164);
nor U203 (N_203,In_5,In_448);
nor U204 (N_204,N_118,N_58);
or U205 (N_205,In_497,In_437);
or U206 (N_206,N_109,In_441);
nor U207 (N_207,In_259,In_329);
xnor U208 (N_208,In_155,In_91);
nor U209 (N_209,N_37,In_18);
nand U210 (N_210,In_156,In_445);
and U211 (N_211,In_438,In_227);
or U212 (N_212,In_280,In_307);
xnor U213 (N_213,In_206,N_41);
xor U214 (N_214,In_70,N_134);
nor U215 (N_215,In_414,N_106);
nand U216 (N_216,N_111,In_234);
and U217 (N_217,In_231,In_308);
or U218 (N_218,In_286,In_214);
or U219 (N_219,In_117,In_66);
nor U220 (N_220,N_80,In_388);
xor U221 (N_221,In_132,In_387);
nand U222 (N_222,N_82,In_160);
nor U223 (N_223,N_15,N_129);
nor U224 (N_224,N_89,In_1);
nor U225 (N_225,In_73,In_270);
and U226 (N_226,In_369,In_486);
or U227 (N_227,N_174,N_191);
or U228 (N_228,In_229,N_214);
xor U229 (N_229,In_460,In_161);
and U230 (N_230,N_76,N_74);
and U231 (N_231,In_466,N_114);
nand U232 (N_232,N_91,In_30);
nand U233 (N_233,N_178,In_481);
nand U234 (N_234,In_253,N_139);
xor U235 (N_235,N_127,In_251);
xor U236 (N_236,N_211,In_96);
xnor U237 (N_237,In_144,In_189);
nor U238 (N_238,In_491,N_38);
and U239 (N_239,In_32,N_169);
nand U240 (N_240,In_277,N_172);
nor U241 (N_241,N_197,In_483);
xnor U242 (N_242,N_99,In_65);
nand U243 (N_243,In_62,N_216);
nand U244 (N_244,In_77,In_210);
or U245 (N_245,In_397,N_66);
nand U246 (N_246,In_40,In_375);
and U247 (N_247,N_179,In_403);
nand U248 (N_248,N_164,N_185);
and U249 (N_249,In_349,N_112);
and U250 (N_250,N_157,N_220);
and U251 (N_251,N_136,N_95);
and U252 (N_252,In_184,N_51);
nand U253 (N_253,N_9,In_75);
nor U254 (N_254,In_320,In_131);
and U255 (N_255,N_155,N_224);
xor U256 (N_256,In_35,In_226);
xnor U257 (N_257,In_191,In_180);
nor U258 (N_258,In_37,N_46);
xor U259 (N_259,In_19,In_54);
nor U260 (N_260,N_203,N_119);
or U261 (N_261,In_390,N_88);
and U262 (N_262,In_315,N_175);
xnor U263 (N_263,In_384,N_199);
xnor U264 (N_264,In_43,In_257);
or U265 (N_265,N_68,N_167);
or U266 (N_266,In_211,N_162);
or U267 (N_267,N_30,N_123);
xnor U268 (N_268,In_120,In_223);
xor U269 (N_269,N_73,N_209);
and U270 (N_270,In_24,In_224);
and U271 (N_271,In_347,In_262);
nor U272 (N_272,In_46,In_212);
or U273 (N_273,N_198,In_357);
nor U274 (N_274,In_122,In_268);
nand U275 (N_275,N_146,N_138);
or U276 (N_276,In_469,N_150);
nor U277 (N_277,In_490,N_218);
or U278 (N_278,N_210,In_279);
nor U279 (N_279,N_171,In_250);
and U280 (N_280,N_113,N_141);
xnor U281 (N_281,In_7,N_110);
or U282 (N_282,N_212,N_34);
nor U283 (N_283,In_454,N_183);
nand U284 (N_284,N_90,N_102);
nand U285 (N_285,In_385,In_195);
xor U286 (N_286,N_116,N_64);
xor U287 (N_287,N_154,N_132);
or U288 (N_288,N_147,N_13);
or U289 (N_289,N_54,N_193);
nand U290 (N_290,In_152,N_202);
nand U291 (N_291,N_16,In_494);
and U292 (N_292,N_192,In_341);
or U293 (N_293,N_184,In_496);
xnor U294 (N_294,N_17,N_200);
or U295 (N_295,N_158,In_291);
and U296 (N_296,In_478,In_455);
and U297 (N_297,In_322,In_411);
nor U298 (N_298,In_381,N_75);
nand U299 (N_299,In_433,N_27);
xor U300 (N_300,N_261,N_295);
xor U301 (N_301,N_291,N_81);
nand U302 (N_302,In_105,N_107);
or U303 (N_303,In_194,N_57);
nor U304 (N_304,In_133,N_144);
or U305 (N_305,N_145,N_122);
or U306 (N_306,N_231,N_285);
and U307 (N_307,N_26,N_238);
nor U308 (N_308,N_124,N_284);
and U309 (N_309,N_8,N_70);
nand U310 (N_310,N_204,N_242);
xor U311 (N_311,In_217,N_149);
or U312 (N_312,N_298,N_264);
nor U313 (N_313,N_133,N_100);
nor U314 (N_314,N_260,In_135);
xnor U315 (N_315,N_265,N_266);
and U316 (N_316,N_249,N_257);
nand U317 (N_317,N_246,N_10);
xor U318 (N_318,N_276,N_21);
nand U319 (N_319,N_253,N_296);
nand U320 (N_320,N_235,In_366);
and U321 (N_321,In_467,N_288);
nand U322 (N_322,N_289,In_177);
and U323 (N_323,N_290,In_165);
or U324 (N_324,In_290,N_297);
xor U325 (N_325,N_280,N_256);
nor U326 (N_326,N_279,N_180);
xor U327 (N_327,N_236,N_94);
or U328 (N_328,N_161,N_195);
and U329 (N_329,N_173,N_259);
nand U330 (N_330,N_254,N_247);
nand U331 (N_331,In_116,N_101);
or U332 (N_332,In_261,N_232);
nor U333 (N_333,N_117,N_240);
or U334 (N_334,N_226,In_71);
or U335 (N_335,N_293,N_170);
nand U336 (N_336,In_11,N_176);
and U337 (N_337,In_424,N_292);
xnor U338 (N_338,In_485,N_159);
nor U339 (N_339,N_40,In_14);
nand U340 (N_340,N_250,N_251);
or U341 (N_341,N_294,N_201);
nor U342 (N_342,N_281,In_428);
xor U343 (N_343,In_87,In_396);
nor U344 (N_344,N_207,N_269);
or U345 (N_345,N_248,N_217);
nor U346 (N_346,N_221,N_215);
and U347 (N_347,N_229,N_262);
and U348 (N_348,N_50,N_28);
and U349 (N_349,N_177,In_365);
nor U350 (N_350,In_59,N_206);
nand U351 (N_351,N_273,N_283);
nand U352 (N_352,N_160,N_244);
or U353 (N_353,In_299,N_190);
xnor U354 (N_354,N_156,In_353);
nand U355 (N_355,In_379,N_55);
xor U356 (N_356,N_7,N_151);
nand U357 (N_357,N_194,In_302);
or U358 (N_358,N_19,N_168);
nor U359 (N_359,N_287,N_153);
or U360 (N_360,N_223,N_233);
and U361 (N_361,In_115,N_3);
nand U362 (N_362,In_158,N_234);
or U363 (N_363,N_275,N_282);
or U364 (N_364,N_196,N_271);
and U365 (N_365,In_134,N_252);
nor U366 (N_366,N_274,In_232);
nand U367 (N_367,In_179,N_219);
or U368 (N_368,N_86,N_270);
nor U369 (N_369,In_267,In_377);
nand U370 (N_370,N_188,N_182);
nor U371 (N_371,N_83,N_205);
nand U372 (N_372,N_267,N_33);
nand U373 (N_373,N_299,In_213);
nor U374 (N_374,N_165,In_493);
xor U375 (N_375,N_189,N_186);
nand U376 (N_376,N_303,N_338);
and U377 (N_377,N_263,In_401);
nor U378 (N_378,N_243,N_181);
and U379 (N_379,N_339,N_300);
nor U380 (N_380,N_327,N_346);
nor U381 (N_381,N_125,N_358);
xor U382 (N_382,N_341,In_209);
nor U383 (N_383,N_372,N_364);
and U384 (N_384,In_278,N_308);
xor U385 (N_385,N_96,N_360);
nor U386 (N_386,N_268,N_239);
and U387 (N_387,N_255,N_301);
nor U388 (N_388,N_329,N_366);
nor U389 (N_389,N_69,In_27);
or U390 (N_390,N_163,N_373);
xnor U391 (N_391,N_348,N_166);
nand U392 (N_392,N_325,In_200);
xor U393 (N_393,N_230,N_228);
nor U394 (N_394,N_152,N_352);
nor U395 (N_395,N_359,N_309);
nor U396 (N_396,N_187,N_237);
and U397 (N_397,N_353,N_347);
nor U398 (N_398,N_342,N_337);
and U399 (N_399,N_355,N_310);
or U400 (N_400,N_227,N_315);
nor U401 (N_401,In_107,N_272);
and U402 (N_402,N_369,N_374);
xnor U403 (N_403,N_258,N_305);
or U404 (N_404,In_149,N_356);
nand U405 (N_405,In_196,In_138);
and U406 (N_406,N_365,N_334);
nor U407 (N_407,N_208,N_331);
nor U408 (N_408,N_344,N_311);
nor U409 (N_409,N_318,N_104);
nor U410 (N_410,N_316,N_357);
nor U411 (N_411,In_297,N_313);
and U412 (N_412,N_241,N_336);
nand U413 (N_413,N_371,N_368);
or U414 (N_414,N_343,N_322);
nand U415 (N_415,N_350,N_354);
and U416 (N_416,N_367,N_245);
nand U417 (N_417,N_351,N_319);
nand U418 (N_418,N_323,N_317);
xor U419 (N_419,N_370,N_312);
xnor U420 (N_420,N_306,N_345);
nor U421 (N_421,In_288,N_79);
and U422 (N_422,N_362,In_484);
nand U423 (N_423,N_302,N_105);
nand U424 (N_424,N_320,N_321);
or U425 (N_425,N_363,N_332);
nor U426 (N_426,N_324,N_314);
and U427 (N_427,In_311,N_326);
nand U428 (N_428,N_307,N_361);
and U429 (N_429,N_340,N_278);
or U430 (N_430,In_228,N_213);
and U431 (N_431,N_286,In_63);
or U432 (N_432,N_23,N_225);
nand U433 (N_433,N_328,N_304);
and U434 (N_434,N_333,N_335);
and U435 (N_435,N_222,N_277);
nor U436 (N_436,N_349,In_199);
xor U437 (N_437,N_330,N_337);
or U438 (N_438,N_305,N_166);
nor U439 (N_439,N_339,N_349);
xnor U440 (N_440,N_340,N_329);
and U441 (N_441,N_349,N_351);
nand U442 (N_442,In_297,In_209);
nand U443 (N_443,N_330,N_186);
nor U444 (N_444,N_258,N_340);
xor U445 (N_445,N_372,N_333);
and U446 (N_446,In_200,N_327);
xnor U447 (N_447,N_163,N_327);
and U448 (N_448,N_314,N_228);
or U449 (N_449,N_363,N_321);
or U450 (N_450,N_377,N_397);
nand U451 (N_451,N_378,N_415);
and U452 (N_452,N_433,N_398);
xnor U453 (N_453,N_394,N_401);
and U454 (N_454,N_385,N_439);
and U455 (N_455,N_403,N_426);
xnor U456 (N_456,N_434,N_440);
nor U457 (N_457,N_384,N_423);
and U458 (N_458,N_445,N_446);
nor U459 (N_459,N_404,N_392);
xor U460 (N_460,N_443,N_422);
or U461 (N_461,N_387,N_391);
nor U462 (N_462,N_409,N_438);
and U463 (N_463,N_442,N_393);
nand U464 (N_464,N_413,N_379);
xor U465 (N_465,N_380,N_437);
nand U466 (N_466,N_389,N_382);
nor U467 (N_467,N_421,N_381);
xnor U468 (N_468,N_400,N_430);
or U469 (N_469,N_417,N_375);
or U470 (N_470,N_447,N_424);
or U471 (N_471,N_388,N_432);
nand U472 (N_472,N_402,N_431);
nor U473 (N_473,N_399,N_436);
nor U474 (N_474,N_405,N_414);
nor U475 (N_475,N_406,N_416);
xnor U476 (N_476,N_383,N_412);
nand U477 (N_477,N_420,N_425);
or U478 (N_478,N_418,N_444);
nand U479 (N_479,N_410,N_411);
nor U480 (N_480,N_428,N_427);
nand U481 (N_481,N_395,N_449);
and U482 (N_482,N_386,N_376);
nand U483 (N_483,N_441,N_448);
nor U484 (N_484,N_396,N_419);
nand U485 (N_485,N_435,N_407);
xor U486 (N_486,N_429,N_408);
and U487 (N_487,N_390,N_386);
xnor U488 (N_488,N_384,N_391);
or U489 (N_489,N_440,N_392);
nor U490 (N_490,N_428,N_385);
nand U491 (N_491,N_443,N_408);
xnor U492 (N_492,N_426,N_448);
nor U493 (N_493,N_406,N_386);
nand U494 (N_494,N_444,N_429);
nand U495 (N_495,N_400,N_394);
nor U496 (N_496,N_422,N_387);
and U497 (N_497,N_415,N_400);
and U498 (N_498,N_381,N_393);
xor U499 (N_499,N_415,N_401);
xor U500 (N_500,N_434,N_393);
and U501 (N_501,N_395,N_398);
and U502 (N_502,N_406,N_414);
nand U503 (N_503,N_440,N_384);
or U504 (N_504,N_441,N_428);
nand U505 (N_505,N_439,N_375);
nand U506 (N_506,N_427,N_417);
xor U507 (N_507,N_388,N_375);
xnor U508 (N_508,N_415,N_388);
nor U509 (N_509,N_445,N_441);
or U510 (N_510,N_442,N_403);
xor U511 (N_511,N_375,N_426);
nand U512 (N_512,N_436,N_392);
and U513 (N_513,N_424,N_389);
xnor U514 (N_514,N_388,N_409);
xor U515 (N_515,N_387,N_441);
nor U516 (N_516,N_423,N_388);
or U517 (N_517,N_400,N_405);
nand U518 (N_518,N_401,N_390);
and U519 (N_519,N_432,N_389);
nand U520 (N_520,N_416,N_428);
nand U521 (N_521,N_428,N_442);
nand U522 (N_522,N_385,N_389);
or U523 (N_523,N_398,N_439);
nor U524 (N_524,N_385,N_381);
nor U525 (N_525,N_503,N_455);
nor U526 (N_526,N_464,N_451);
and U527 (N_527,N_514,N_518);
nand U528 (N_528,N_459,N_493);
xnor U529 (N_529,N_521,N_462);
nand U530 (N_530,N_502,N_512);
xnor U531 (N_531,N_468,N_507);
xnor U532 (N_532,N_454,N_513);
and U533 (N_533,N_463,N_487);
or U534 (N_534,N_509,N_504);
nor U535 (N_535,N_480,N_465);
and U536 (N_536,N_467,N_510);
or U537 (N_537,N_479,N_469);
xnor U538 (N_538,N_453,N_488);
nand U539 (N_539,N_461,N_483);
nor U540 (N_540,N_499,N_520);
nand U541 (N_541,N_497,N_485);
or U542 (N_542,N_523,N_466);
or U543 (N_543,N_473,N_470);
nand U544 (N_544,N_489,N_492);
or U545 (N_545,N_478,N_495);
or U546 (N_546,N_458,N_474);
and U547 (N_547,N_494,N_472);
xnor U548 (N_548,N_475,N_498);
nand U549 (N_549,N_516,N_491);
xor U550 (N_550,N_477,N_501);
nor U551 (N_551,N_486,N_505);
or U552 (N_552,N_519,N_456);
nand U553 (N_553,N_515,N_522);
and U554 (N_554,N_471,N_508);
or U555 (N_555,N_517,N_482);
nand U556 (N_556,N_506,N_496);
xor U557 (N_557,N_452,N_460);
nor U558 (N_558,N_524,N_500);
or U559 (N_559,N_490,N_481);
nand U560 (N_560,N_476,N_484);
or U561 (N_561,N_511,N_450);
and U562 (N_562,N_457,N_491);
or U563 (N_563,N_509,N_511);
nor U564 (N_564,N_522,N_466);
nand U565 (N_565,N_460,N_514);
and U566 (N_566,N_474,N_522);
or U567 (N_567,N_486,N_465);
xor U568 (N_568,N_459,N_454);
or U569 (N_569,N_496,N_468);
and U570 (N_570,N_454,N_499);
nand U571 (N_571,N_509,N_517);
xor U572 (N_572,N_456,N_459);
nor U573 (N_573,N_456,N_472);
or U574 (N_574,N_494,N_503);
nor U575 (N_575,N_503,N_483);
or U576 (N_576,N_458,N_499);
nor U577 (N_577,N_500,N_451);
or U578 (N_578,N_464,N_509);
and U579 (N_579,N_461,N_511);
xor U580 (N_580,N_498,N_494);
xnor U581 (N_581,N_458,N_468);
and U582 (N_582,N_487,N_490);
or U583 (N_583,N_465,N_492);
and U584 (N_584,N_516,N_493);
nor U585 (N_585,N_498,N_478);
xor U586 (N_586,N_486,N_457);
or U587 (N_587,N_517,N_501);
nand U588 (N_588,N_486,N_493);
and U589 (N_589,N_521,N_490);
and U590 (N_590,N_485,N_524);
nand U591 (N_591,N_477,N_512);
xor U592 (N_592,N_513,N_521);
nor U593 (N_593,N_490,N_460);
nand U594 (N_594,N_452,N_468);
nand U595 (N_595,N_503,N_495);
and U596 (N_596,N_453,N_518);
and U597 (N_597,N_484,N_471);
or U598 (N_598,N_474,N_496);
nor U599 (N_599,N_466,N_462);
nand U600 (N_600,N_592,N_565);
nor U601 (N_601,N_552,N_580);
and U602 (N_602,N_582,N_590);
or U603 (N_603,N_527,N_526);
nor U604 (N_604,N_563,N_534);
xor U605 (N_605,N_569,N_573);
xor U606 (N_606,N_591,N_566);
or U607 (N_607,N_581,N_564);
and U608 (N_608,N_574,N_542);
and U609 (N_609,N_529,N_568);
and U610 (N_610,N_586,N_541);
nor U611 (N_611,N_560,N_567);
nor U612 (N_612,N_561,N_575);
nand U613 (N_613,N_555,N_543);
and U614 (N_614,N_539,N_597);
and U615 (N_615,N_593,N_595);
xor U616 (N_616,N_584,N_557);
or U617 (N_617,N_535,N_544);
nand U618 (N_618,N_545,N_559);
and U619 (N_619,N_598,N_525);
xor U620 (N_620,N_556,N_530);
or U621 (N_621,N_570,N_547);
and U622 (N_622,N_546,N_528);
nand U623 (N_623,N_579,N_576);
nor U624 (N_624,N_558,N_553);
and U625 (N_625,N_589,N_585);
nor U626 (N_626,N_562,N_588);
nor U627 (N_627,N_549,N_532);
nand U628 (N_628,N_578,N_554);
nor U629 (N_629,N_577,N_531);
nand U630 (N_630,N_536,N_551);
nand U631 (N_631,N_599,N_596);
nand U632 (N_632,N_571,N_533);
or U633 (N_633,N_587,N_538);
or U634 (N_634,N_540,N_583);
nor U635 (N_635,N_550,N_572);
or U636 (N_636,N_548,N_594);
or U637 (N_637,N_537,N_576);
and U638 (N_638,N_596,N_560);
nand U639 (N_639,N_543,N_529);
or U640 (N_640,N_557,N_533);
nor U641 (N_641,N_541,N_583);
or U642 (N_642,N_548,N_532);
xnor U643 (N_643,N_563,N_536);
xor U644 (N_644,N_549,N_531);
or U645 (N_645,N_598,N_568);
nand U646 (N_646,N_575,N_574);
and U647 (N_647,N_543,N_564);
or U648 (N_648,N_541,N_559);
nand U649 (N_649,N_560,N_590);
or U650 (N_650,N_532,N_563);
xnor U651 (N_651,N_568,N_587);
and U652 (N_652,N_551,N_578);
nand U653 (N_653,N_557,N_587);
nor U654 (N_654,N_533,N_551);
nor U655 (N_655,N_597,N_585);
xnor U656 (N_656,N_593,N_526);
xor U657 (N_657,N_584,N_542);
xnor U658 (N_658,N_575,N_538);
nand U659 (N_659,N_533,N_559);
and U660 (N_660,N_565,N_533);
nand U661 (N_661,N_567,N_571);
nor U662 (N_662,N_543,N_527);
xnor U663 (N_663,N_552,N_599);
nand U664 (N_664,N_587,N_539);
and U665 (N_665,N_575,N_589);
xor U666 (N_666,N_547,N_595);
nand U667 (N_667,N_576,N_544);
or U668 (N_668,N_598,N_554);
or U669 (N_669,N_561,N_539);
nor U670 (N_670,N_569,N_538);
and U671 (N_671,N_594,N_598);
xor U672 (N_672,N_534,N_570);
or U673 (N_673,N_563,N_554);
and U674 (N_674,N_531,N_589);
xor U675 (N_675,N_618,N_611);
nand U676 (N_676,N_652,N_644);
xor U677 (N_677,N_637,N_657);
nor U678 (N_678,N_669,N_602);
xor U679 (N_679,N_648,N_634);
nor U680 (N_680,N_667,N_638);
nand U681 (N_681,N_646,N_614);
nor U682 (N_682,N_641,N_615);
xor U683 (N_683,N_672,N_630);
xor U684 (N_684,N_651,N_640);
and U685 (N_685,N_655,N_619);
nor U686 (N_686,N_626,N_600);
or U687 (N_687,N_649,N_617);
xor U688 (N_688,N_665,N_662);
xor U689 (N_689,N_621,N_663);
and U690 (N_690,N_653,N_613);
or U691 (N_691,N_620,N_624);
xor U692 (N_692,N_609,N_606);
nor U693 (N_693,N_612,N_647);
or U694 (N_694,N_608,N_604);
or U695 (N_695,N_635,N_616);
xor U696 (N_696,N_636,N_656);
xor U697 (N_697,N_642,N_650);
xnor U698 (N_698,N_628,N_659);
xnor U699 (N_699,N_661,N_603);
nand U700 (N_700,N_632,N_610);
nand U701 (N_701,N_631,N_627);
nand U702 (N_702,N_668,N_622);
nand U703 (N_703,N_645,N_658);
and U704 (N_704,N_643,N_625);
and U705 (N_705,N_654,N_670);
nand U706 (N_706,N_633,N_639);
xnor U707 (N_707,N_664,N_629);
nor U708 (N_708,N_666,N_660);
nor U709 (N_709,N_607,N_601);
or U710 (N_710,N_673,N_605);
nand U711 (N_711,N_623,N_671);
nor U712 (N_712,N_674,N_652);
and U713 (N_713,N_620,N_654);
and U714 (N_714,N_630,N_673);
nor U715 (N_715,N_641,N_619);
and U716 (N_716,N_650,N_669);
nor U717 (N_717,N_635,N_646);
and U718 (N_718,N_639,N_608);
or U719 (N_719,N_640,N_672);
nand U720 (N_720,N_652,N_658);
nand U721 (N_721,N_613,N_612);
and U722 (N_722,N_673,N_645);
or U723 (N_723,N_610,N_668);
and U724 (N_724,N_630,N_620);
xnor U725 (N_725,N_635,N_673);
xor U726 (N_726,N_664,N_630);
xnor U727 (N_727,N_638,N_622);
or U728 (N_728,N_673,N_610);
nand U729 (N_729,N_652,N_649);
or U730 (N_730,N_672,N_673);
or U731 (N_731,N_663,N_623);
or U732 (N_732,N_615,N_668);
or U733 (N_733,N_600,N_601);
nor U734 (N_734,N_629,N_628);
nor U735 (N_735,N_632,N_648);
nor U736 (N_736,N_617,N_650);
nand U737 (N_737,N_610,N_671);
nand U738 (N_738,N_605,N_658);
or U739 (N_739,N_658,N_648);
or U740 (N_740,N_615,N_612);
xor U741 (N_741,N_667,N_670);
xnor U742 (N_742,N_640,N_673);
or U743 (N_743,N_618,N_649);
or U744 (N_744,N_649,N_645);
xnor U745 (N_745,N_609,N_626);
nand U746 (N_746,N_655,N_672);
nor U747 (N_747,N_602,N_667);
or U748 (N_748,N_671,N_618);
and U749 (N_749,N_668,N_650);
or U750 (N_750,N_707,N_682);
or U751 (N_751,N_700,N_701);
nor U752 (N_752,N_677,N_730);
xnor U753 (N_753,N_721,N_676);
nor U754 (N_754,N_708,N_729);
and U755 (N_755,N_732,N_741);
or U756 (N_756,N_749,N_702);
and U757 (N_757,N_726,N_713);
or U758 (N_758,N_740,N_716);
and U759 (N_759,N_699,N_748);
xor U760 (N_760,N_731,N_703);
xnor U761 (N_761,N_675,N_733);
and U762 (N_762,N_711,N_745);
xor U763 (N_763,N_697,N_693);
nand U764 (N_764,N_747,N_737);
or U765 (N_765,N_718,N_719);
nor U766 (N_766,N_717,N_685);
and U767 (N_767,N_678,N_690);
and U768 (N_768,N_680,N_743);
and U769 (N_769,N_738,N_728);
xnor U770 (N_770,N_710,N_709);
xor U771 (N_771,N_739,N_694);
and U772 (N_772,N_727,N_746);
and U773 (N_773,N_712,N_706);
and U774 (N_774,N_723,N_735);
and U775 (N_775,N_696,N_681);
and U776 (N_776,N_687,N_695);
and U777 (N_777,N_720,N_698);
or U778 (N_778,N_689,N_742);
or U779 (N_779,N_714,N_736);
xor U780 (N_780,N_715,N_724);
nor U781 (N_781,N_684,N_686);
or U782 (N_782,N_705,N_683);
or U783 (N_783,N_679,N_692);
xor U784 (N_784,N_744,N_691);
nand U785 (N_785,N_704,N_734);
or U786 (N_786,N_725,N_722);
xor U787 (N_787,N_688,N_680);
nand U788 (N_788,N_706,N_682);
or U789 (N_789,N_724,N_743);
or U790 (N_790,N_730,N_716);
nand U791 (N_791,N_695,N_724);
or U792 (N_792,N_680,N_679);
or U793 (N_793,N_690,N_698);
xor U794 (N_794,N_696,N_689);
nand U795 (N_795,N_677,N_682);
or U796 (N_796,N_716,N_737);
nor U797 (N_797,N_737,N_741);
nor U798 (N_798,N_692,N_697);
nand U799 (N_799,N_729,N_748);
xnor U800 (N_800,N_676,N_711);
nand U801 (N_801,N_706,N_691);
nor U802 (N_802,N_701,N_736);
nor U803 (N_803,N_719,N_724);
nand U804 (N_804,N_691,N_742);
xor U805 (N_805,N_717,N_733);
xnor U806 (N_806,N_686,N_685);
xnor U807 (N_807,N_732,N_733);
xor U808 (N_808,N_678,N_719);
and U809 (N_809,N_714,N_738);
nand U810 (N_810,N_707,N_722);
and U811 (N_811,N_690,N_722);
nand U812 (N_812,N_731,N_749);
and U813 (N_813,N_729,N_682);
and U814 (N_814,N_693,N_701);
nand U815 (N_815,N_732,N_712);
nor U816 (N_816,N_725,N_692);
nand U817 (N_817,N_707,N_744);
nor U818 (N_818,N_723,N_694);
nand U819 (N_819,N_698,N_721);
nand U820 (N_820,N_713,N_690);
nor U821 (N_821,N_741,N_730);
nor U822 (N_822,N_710,N_713);
nand U823 (N_823,N_731,N_724);
xnor U824 (N_824,N_699,N_697);
xor U825 (N_825,N_796,N_793);
and U826 (N_826,N_766,N_787);
xnor U827 (N_827,N_761,N_789);
xor U828 (N_828,N_801,N_790);
or U829 (N_829,N_763,N_803);
and U830 (N_830,N_802,N_795);
or U831 (N_831,N_778,N_797);
nand U832 (N_832,N_772,N_807);
xor U833 (N_833,N_794,N_819);
nor U834 (N_834,N_750,N_815);
xnor U835 (N_835,N_785,N_817);
or U836 (N_836,N_756,N_823);
nand U837 (N_837,N_820,N_800);
nand U838 (N_838,N_788,N_783);
nand U839 (N_839,N_768,N_755);
nand U840 (N_840,N_760,N_753);
nand U841 (N_841,N_792,N_799);
nand U842 (N_842,N_804,N_782);
or U843 (N_843,N_786,N_822);
nor U844 (N_844,N_821,N_816);
nand U845 (N_845,N_818,N_762);
nor U846 (N_846,N_777,N_805);
xnor U847 (N_847,N_813,N_764);
or U848 (N_848,N_770,N_798);
nand U849 (N_849,N_767,N_781);
xnor U850 (N_850,N_775,N_774);
nand U851 (N_851,N_752,N_776);
nand U852 (N_852,N_824,N_771);
nor U853 (N_853,N_784,N_759);
xor U854 (N_854,N_809,N_779);
or U855 (N_855,N_765,N_751);
and U856 (N_856,N_811,N_812);
nor U857 (N_857,N_769,N_791);
nand U858 (N_858,N_808,N_780);
xor U859 (N_859,N_773,N_810);
and U860 (N_860,N_814,N_754);
and U861 (N_861,N_758,N_757);
or U862 (N_862,N_806,N_801);
nor U863 (N_863,N_753,N_797);
or U864 (N_864,N_777,N_811);
xnor U865 (N_865,N_750,N_765);
xnor U866 (N_866,N_780,N_760);
nor U867 (N_867,N_808,N_784);
nand U868 (N_868,N_772,N_798);
nand U869 (N_869,N_792,N_806);
nor U870 (N_870,N_814,N_769);
or U871 (N_871,N_768,N_784);
or U872 (N_872,N_763,N_814);
xor U873 (N_873,N_815,N_756);
and U874 (N_874,N_822,N_797);
xnor U875 (N_875,N_794,N_795);
and U876 (N_876,N_818,N_785);
and U877 (N_877,N_814,N_813);
nand U878 (N_878,N_778,N_805);
xnor U879 (N_879,N_769,N_772);
nand U880 (N_880,N_772,N_809);
or U881 (N_881,N_769,N_765);
xnor U882 (N_882,N_750,N_812);
nor U883 (N_883,N_789,N_811);
or U884 (N_884,N_776,N_795);
or U885 (N_885,N_756,N_801);
and U886 (N_886,N_823,N_771);
and U887 (N_887,N_811,N_757);
nand U888 (N_888,N_815,N_773);
nor U889 (N_889,N_774,N_765);
nor U890 (N_890,N_758,N_819);
nand U891 (N_891,N_823,N_788);
nand U892 (N_892,N_800,N_770);
nor U893 (N_893,N_818,N_753);
or U894 (N_894,N_765,N_789);
and U895 (N_895,N_793,N_819);
nor U896 (N_896,N_813,N_803);
nand U897 (N_897,N_796,N_794);
or U898 (N_898,N_751,N_783);
or U899 (N_899,N_821,N_773);
nand U900 (N_900,N_897,N_862);
nor U901 (N_901,N_848,N_857);
or U902 (N_902,N_843,N_870);
or U903 (N_903,N_827,N_828);
xor U904 (N_904,N_888,N_837);
nand U905 (N_905,N_880,N_891);
nor U906 (N_906,N_833,N_853);
nand U907 (N_907,N_842,N_894);
and U908 (N_908,N_844,N_845);
and U909 (N_909,N_831,N_825);
or U910 (N_910,N_875,N_855);
and U911 (N_911,N_834,N_873);
or U912 (N_912,N_850,N_832);
nand U913 (N_913,N_858,N_830);
xnor U914 (N_914,N_866,N_841);
and U915 (N_915,N_881,N_892);
xor U916 (N_916,N_860,N_884);
and U917 (N_917,N_851,N_864);
and U918 (N_918,N_854,N_826);
nor U919 (N_919,N_836,N_871);
or U920 (N_920,N_869,N_876);
nor U921 (N_921,N_878,N_889);
or U922 (N_922,N_839,N_896);
and U923 (N_923,N_890,N_829);
and U924 (N_924,N_847,N_898);
nor U925 (N_925,N_879,N_887);
xnor U926 (N_926,N_861,N_874);
and U927 (N_927,N_886,N_846);
and U928 (N_928,N_840,N_872);
nand U929 (N_929,N_882,N_856);
and U930 (N_930,N_849,N_838);
nand U931 (N_931,N_852,N_893);
or U932 (N_932,N_885,N_895);
xor U933 (N_933,N_899,N_865);
nand U934 (N_934,N_863,N_877);
nor U935 (N_935,N_883,N_868);
and U936 (N_936,N_867,N_835);
nor U937 (N_937,N_859,N_852);
and U938 (N_938,N_894,N_858);
or U939 (N_939,N_881,N_829);
or U940 (N_940,N_891,N_855);
or U941 (N_941,N_826,N_831);
nor U942 (N_942,N_848,N_828);
xor U943 (N_943,N_836,N_860);
and U944 (N_944,N_876,N_843);
nor U945 (N_945,N_862,N_844);
or U946 (N_946,N_838,N_846);
nand U947 (N_947,N_878,N_868);
or U948 (N_948,N_880,N_860);
nand U949 (N_949,N_896,N_843);
or U950 (N_950,N_864,N_836);
nand U951 (N_951,N_852,N_854);
nand U952 (N_952,N_889,N_876);
xor U953 (N_953,N_895,N_890);
xor U954 (N_954,N_879,N_873);
and U955 (N_955,N_880,N_845);
nor U956 (N_956,N_856,N_843);
and U957 (N_957,N_875,N_831);
xnor U958 (N_958,N_872,N_826);
nor U959 (N_959,N_892,N_888);
and U960 (N_960,N_860,N_837);
xnor U961 (N_961,N_862,N_869);
nand U962 (N_962,N_845,N_825);
or U963 (N_963,N_873,N_897);
nor U964 (N_964,N_860,N_830);
nand U965 (N_965,N_827,N_834);
xor U966 (N_966,N_895,N_854);
or U967 (N_967,N_896,N_898);
nand U968 (N_968,N_853,N_844);
or U969 (N_969,N_848,N_861);
and U970 (N_970,N_826,N_849);
xor U971 (N_971,N_893,N_886);
nand U972 (N_972,N_850,N_873);
or U973 (N_973,N_841,N_838);
and U974 (N_974,N_847,N_825);
and U975 (N_975,N_969,N_923);
nand U976 (N_976,N_922,N_951);
nor U977 (N_977,N_971,N_943);
xor U978 (N_978,N_927,N_949);
nor U979 (N_979,N_937,N_954);
and U980 (N_980,N_941,N_912);
nor U981 (N_981,N_965,N_911);
xnor U982 (N_982,N_915,N_903);
xor U983 (N_983,N_914,N_945);
and U984 (N_984,N_913,N_935);
nor U985 (N_985,N_905,N_932);
nor U986 (N_986,N_936,N_955);
and U987 (N_987,N_973,N_925);
and U988 (N_988,N_956,N_916);
nand U989 (N_989,N_967,N_901);
or U990 (N_990,N_960,N_953);
nor U991 (N_991,N_972,N_940);
or U992 (N_992,N_946,N_910);
and U993 (N_993,N_963,N_902);
xor U994 (N_994,N_970,N_900);
nor U995 (N_995,N_928,N_944);
or U996 (N_996,N_966,N_924);
and U997 (N_997,N_952,N_919);
and U998 (N_998,N_930,N_920);
and U999 (N_999,N_947,N_948);
or U1000 (N_1000,N_909,N_934);
and U1001 (N_1001,N_964,N_950);
nand U1002 (N_1002,N_959,N_906);
xor U1003 (N_1003,N_908,N_974);
nand U1004 (N_1004,N_921,N_958);
nand U1005 (N_1005,N_942,N_918);
or U1006 (N_1006,N_907,N_926);
or U1007 (N_1007,N_962,N_938);
nand U1008 (N_1008,N_931,N_957);
or U1009 (N_1009,N_904,N_929);
xor U1010 (N_1010,N_961,N_968);
or U1011 (N_1011,N_933,N_917);
nor U1012 (N_1012,N_939,N_947);
and U1013 (N_1013,N_942,N_928);
nor U1014 (N_1014,N_952,N_947);
nor U1015 (N_1015,N_949,N_908);
or U1016 (N_1016,N_967,N_944);
and U1017 (N_1017,N_915,N_900);
xnor U1018 (N_1018,N_931,N_939);
nor U1019 (N_1019,N_934,N_910);
nor U1020 (N_1020,N_940,N_926);
or U1021 (N_1021,N_965,N_938);
nand U1022 (N_1022,N_915,N_910);
and U1023 (N_1023,N_935,N_902);
xnor U1024 (N_1024,N_916,N_904);
and U1025 (N_1025,N_932,N_963);
nor U1026 (N_1026,N_910,N_913);
and U1027 (N_1027,N_940,N_959);
and U1028 (N_1028,N_937,N_905);
and U1029 (N_1029,N_954,N_903);
xnor U1030 (N_1030,N_915,N_955);
and U1031 (N_1031,N_965,N_942);
nand U1032 (N_1032,N_966,N_923);
nor U1033 (N_1033,N_901,N_916);
nand U1034 (N_1034,N_969,N_904);
or U1035 (N_1035,N_950,N_968);
nor U1036 (N_1036,N_971,N_904);
nor U1037 (N_1037,N_938,N_923);
and U1038 (N_1038,N_955,N_928);
nor U1039 (N_1039,N_949,N_939);
or U1040 (N_1040,N_931,N_956);
and U1041 (N_1041,N_933,N_932);
and U1042 (N_1042,N_940,N_966);
and U1043 (N_1043,N_903,N_945);
nor U1044 (N_1044,N_926,N_958);
nand U1045 (N_1045,N_949,N_937);
and U1046 (N_1046,N_944,N_971);
nand U1047 (N_1047,N_934,N_942);
xor U1048 (N_1048,N_929,N_917);
xnor U1049 (N_1049,N_927,N_934);
nand U1050 (N_1050,N_1032,N_1010);
and U1051 (N_1051,N_1049,N_1019);
nand U1052 (N_1052,N_1044,N_1040);
nand U1053 (N_1053,N_1045,N_1025);
and U1054 (N_1054,N_994,N_1014);
nor U1055 (N_1055,N_990,N_1047);
or U1056 (N_1056,N_999,N_989);
and U1057 (N_1057,N_1018,N_1038);
xor U1058 (N_1058,N_991,N_975);
and U1059 (N_1059,N_1001,N_1024);
nand U1060 (N_1060,N_1016,N_1041);
or U1061 (N_1061,N_993,N_998);
nand U1062 (N_1062,N_1029,N_1026);
and U1063 (N_1063,N_1013,N_988);
nand U1064 (N_1064,N_981,N_1000);
nor U1065 (N_1065,N_1011,N_995);
xor U1066 (N_1066,N_986,N_1005);
nand U1067 (N_1067,N_1003,N_1035);
and U1068 (N_1068,N_992,N_1048);
xor U1069 (N_1069,N_977,N_1002);
nand U1070 (N_1070,N_984,N_1027);
xnor U1071 (N_1071,N_978,N_996);
nor U1072 (N_1072,N_1022,N_1008);
nand U1073 (N_1073,N_1043,N_987);
and U1074 (N_1074,N_1009,N_982);
nand U1075 (N_1075,N_1020,N_979);
or U1076 (N_1076,N_1023,N_1012);
nor U1077 (N_1077,N_997,N_1017);
xor U1078 (N_1078,N_1039,N_1006);
nor U1079 (N_1079,N_976,N_1034);
nand U1080 (N_1080,N_1007,N_1021);
xnor U1081 (N_1081,N_1046,N_1036);
xnor U1082 (N_1082,N_1031,N_1042);
and U1083 (N_1083,N_1015,N_1033);
nor U1084 (N_1084,N_1028,N_1037);
or U1085 (N_1085,N_983,N_1004);
xor U1086 (N_1086,N_985,N_980);
or U1087 (N_1087,N_1030,N_1036);
nor U1088 (N_1088,N_1043,N_1003);
or U1089 (N_1089,N_990,N_1027);
or U1090 (N_1090,N_998,N_979);
nor U1091 (N_1091,N_1040,N_977);
xor U1092 (N_1092,N_988,N_1017);
nor U1093 (N_1093,N_1015,N_1031);
or U1094 (N_1094,N_994,N_1006);
xor U1095 (N_1095,N_1002,N_990);
or U1096 (N_1096,N_978,N_1016);
nor U1097 (N_1097,N_1017,N_982);
and U1098 (N_1098,N_986,N_1022);
nand U1099 (N_1099,N_984,N_1023);
and U1100 (N_1100,N_1031,N_1037);
nor U1101 (N_1101,N_992,N_986);
xor U1102 (N_1102,N_1038,N_1031);
xor U1103 (N_1103,N_1016,N_1011);
and U1104 (N_1104,N_1048,N_1045);
xnor U1105 (N_1105,N_990,N_992);
nand U1106 (N_1106,N_985,N_992);
and U1107 (N_1107,N_1045,N_1024);
nor U1108 (N_1108,N_1002,N_1033);
or U1109 (N_1109,N_1011,N_1001);
and U1110 (N_1110,N_1041,N_1008);
nand U1111 (N_1111,N_995,N_997);
nand U1112 (N_1112,N_986,N_1001);
or U1113 (N_1113,N_1006,N_1027);
or U1114 (N_1114,N_1038,N_981);
xnor U1115 (N_1115,N_1016,N_1028);
or U1116 (N_1116,N_1027,N_977);
and U1117 (N_1117,N_1014,N_980);
xnor U1118 (N_1118,N_987,N_979);
and U1119 (N_1119,N_1003,N_1040);
and U1120 (N_1120,N_986,N_989);
xor U1121 (N_1121,N_978,N_1038);
xnor U1122 (N_1122,N_992,N_1017);
nand U1123 (N_1123,N_976,N_1010);
and U1124 (N_1124,N_1036,N_1016);
nand U1125 (N_1125,N_1111,N_1079);
xnor U1126 (N_1126,N_1063,N_1058);
or U1127 (N_1127,N_1100,N_1067);
or U1128 (N_1128,N_1066,N_1050);
nand U1129 (N_1129,N_1097,N_1084);
and U1130 (N_1130,N_1075,N_1052);
and U1131 (N_1131,N_1073,N_1062);
or U1132 (N_1132,N_1118,N_1057);
nor U1133 (N_1133,N_1103,N_1116);
or U1134 (N_1134,N_1101,N_1059);
nand U1135 (N_1135,N_1056,N_1053);
nand U1136 (N_1136,N_1077,N_1121);
or U1137 (N_1137,N_1081,N_1098);
and U1138 (N_1138,N_1089,N_1102);
nor U1139 (N_1139,N_1122,N_1068);
or U1140 (N_1140,N_1114,N_1124);
and U1141 (N_1141,N_1117,N_1120);
nand U1142 (N_1142,N_1123,N_1095);
nor U1143 (N_1143,N_1071,N_1106);
nor U1144 (N_1144,N_1107,N_1092);
and U1145 (N_1145,N_1096,N_1072);
nor U1146 (N_1146,N_1085,N_1115);
nand U1147 (N_1147,N_1108,N_1064);
nand U1148 (N_1148,N_1087,N_1113);
and U1149 (N_1149,N_1054,N_1086);
nor U1150 (N_1150,N_1104,N_1076);
or U1151 (N_1151,N_1055,N_1094);
and U1152 (N_1152,N_1083,N_1088);
and U1153 (N_1153,N_1069,N_1051);
nor U1154 (N_1154,N_1090,N_1093);
and U1155 (N_1155,N_1110,N_1109);
nand U1156 (N_1156,N_1060,N_1099);
nand U1157 (N_1157,N_1078,N_1091);
nor U1158 (N_1158,N_1080,N_1070);
nand U1159 (N_1159,N_1105,N_1119);
nand U1160 (N_1160,N_1074,N_1112);
or U1161 (N_1161,N_1065,N_1082);
nand U1162 (N_1162,N_1061,N_1122);
or U1163 (N_1163,N_1116,N_1083);
or U1164 (N_1164,N_1109,N_1092);
and U1165 (N_1165,N_1074,N_1075);
and U1166 (N_1166,N_1076,N_1111);
or U1167 (N_1167,N_1074,N_1050);
or U1168 (N_1168,N_1061,N_1066);
xor U1169 (N_1169,N_1124,N_1071);
xor U1170 (N_1170,N_1071,N_1076);
and U1171 (N_1171,N_1121,N_1115);
nand U1172 (N_1172,N_1111,N_1092);
or U1173 (N_1173,N_1121,N_1082);
nand U1174 (N_1174,N_1116,N_1070);
nand U1175 (N_1175,N_1107,N_1070);
and U1176 (N_1176,N_1096,N_1094);
and U1177 (N_1177,N_1105,N_1071);
and U1178 (N_1178,N_1086,N_1080);
or U1179 (N_1179,N_1050,N_1063);
and U1180 (N_1180,N_1060,N_1057);
nor U1181 (N_1181,N_1088,N_1103);
or U1182 (N_1182,N_1123,N_1055);
nor U1183 (N_1183,N_1059,N_1102);
xor U1184 (N_1184,N_1084,N_1103);
nor U1185 (N_1185,N_1064,N_1078);
or U1186 (N_1186,N_1119,N_1100);
xnor U1187 (N_1187,N_1094,N_1057);
or U1188 (N_1188,N_1070,N_1059);
and U1189 (N_1189,N_1116,N_1072);
nor U1190 (N_1190,N_1071,N_1117);
and U1191 (N_1191,N_1061,N_1089);
nand U1192 (N_1192,N_1099,N_1102);
or U1193 (N_1193,N_1078,N_1062);
and U1194 (N_1194,N_1106,N_1060);
or U1195 (N_1195,N_1055,N_1091);
xor U1196 (N_1196,N_1065,N_1073);
and U1197 (N_1197,N_1071,N_1065);
xnor U1198 (N_1198,N_1062,N_1113);
nor U1199 (N_1199,N_1068,N_1120);
or U1200 (N_1200,N_1141,N_1199);
nor U1201 (N_1201,N_1125,N_1182);
nand U1202 (N_1202,N_1173,N_1193);
nand U1203 (N_1203,N_1139,N_1161);
and U1204 (N_1204,N_1151,N_1190);
nand U1205 (N_1205,N_1138,N_1126);
nor U1206 (N_1206,N_1195,N_1169);
or U1207 (N_1207,N_1148,N_1127);
nor U1208 (N_1208,N_1189,N_1129);
nand U1209 (N_1209,N_1185,N_1156);
nand U1210 (N_1210,N_1130,N_1165);
and U1211 (N_1211,N_1191,N_1146);
nand U1212 (N_1212,N_1176,N_1132);
nor U1213 (N_1213,N_1168,N_1192);
or U1214 (N_1214,N_1147,N_1170);
and U1215 (N_1215,N_1162,N_1140);
xor U1216 (N_1216,N_1197,N_1143);
nand U1217 (N_1217,N_1167,N_1137);
nand U1218 (N_1218,N_1183,N_1184);
nor U1219 (N_1219,N_1135,N_1136);
and U1220 (N_1220,N_1166,N_1194);
nor U1221 (N_1221,N_1177,N_1154);
or U1222 (N_1222,N_1181,N_1198);
xor U1223 (N_1223,N_1128,N_1134);
or U1224 (N_1224,N_1164,N_1150);
or U1225 (N_1225,N_1155,N_1158);
nor U1226 (N_1226,N_1160,N_1188);
xnor U1227 (N_1227,N_1196,N_1174);
xor U1228 (N_1228,N_1153,N_1175);
and U1229 (N_1229,N_1159,N_1163);
xnor U1230 (N_1230,N_1172,N_1145);
and U1231 (N_1231,N_1144,N_1178);
and U1232 (N_1232,N_1179,N_1152);
or U1233 (N_1233,N_1171,N_1133);
and U1234 (N_1234,N_1187,N_1157);
nor U1235 (N_1235,N_1186,N_1180);
xnor U1236 (N_1236,N_1131,N_1149);
or U1237 (N_1237,N_1142,N_1181);
nand U1238 (N_1238,N_1198,N_1180);
nor U1239 (N_1239,N_1163,N_1149);
and U1240 (N_1240,N_1164,N_1183);
or U1241 (N_1241,N_1183,N_1180);
nor U1242 (N_1242,N_1177,N_1153);
nor U1243 (N_1243,N_1147,N_1171);
nor U1244 (N_1244,N_1134,N_1163);
nand U1245 (N_1245,N_1133,N_1185);
nand U1246 (N_1246,N_1163,N_1198);
xor U1247 (N_1247,N_1129,N_1152);
nand U1248 (N_1248,N_1162,N_1199);
nand U1249 (N_1249,N_1149,N_1197);
and U1250 (N_1250,N_1171,N_1130);
xor U1251 (N_1251,N_1170,N_1137);
and U1252 (N_1252,N_1145,N_1165);
or U1253 (N_1253,N_1182,N_1196);
xor U1254 (N_1254,N_1163,N_1169);
xor U1255 (N_1255,N_1165,N_1179);
and U1256 (N_1256,N_1180,N_1193);
nor U1257 (N_1257,N_1196,N_1139);
or U1258 (N_1258,N_1175,N_1150);
nand U1259 (N_1259,N_1136,N_1196);
nand U1260 (N_1260,N_1141,N_1176);
nand U1261 (N_1261,N_1148,N_1198);
nand U1262 (N_1262,N_1156,N_1139);
nor U1263 (N_1263,N_1179,N_1135);
nor U1264 (N_1264,N_1173,N_1151);
xor U1265 (N_1265,N_1155,N_1136);
or U1266 (N_1266,N_1176,N_1154);
xnor U1267 (N_1267,N_1146,N_1183);
nand U1268 (N_1268,N_1154,N_1157);
or U1269 (N_1269,N_1136,N_1141);
xor U1270 (N_1270,N_1192,N_1197);
nand U1271 (N_1271,N_1132,N_1199);
xnor U1272 (N_1272,N_1152,N_1153);
nand U1273 (N_1273,N_1188,N_1191);
or U1274 (N_1274,N_1196,N_1129);
or U1275 (N_1275,N_1246,N_1264);
nor U1276 (N_1276,N_1217,N_1238);
nor U1277 (N_1277,N_1207,N_1213);
and U1278 (N_1278,N_1253,N_1240);
and U1279 (N_1279,N_1204,N_1218);
nor U1280 (N_1280,N_1252,N_1258);
xor U1281 (N_1281,N_1248,N_1254);
nor U1282 (N_1282,N_1251,N_1268);
and U1283 (N_1283,N_1230,N_1249);
nor U1284 (N_1284,N_1242,N_1224);
nand U1285 (N_1285,N_1244,N_1260);
xnor U1286 (N_1286,N_1227,N_1209);
or U1287 (N_1287,N_1250,N_1234);
nor U1288 (N_1288,N_1257,N_1262);
or U1289 (N_1289,N_1226,N_1229);
xor U1290 (N_1290,N_1273,N_1236);
or U1291 (N_1291,N_1271,N_1266);
nand U1292 (N_1292,N_1272,N_1269);
xor U1293 (N_1293,N_1263,N_1200);
or U1294 (N_1294,N_1243,N_1232);
nor U1295 (N_1295,N_1208,N_1219);
xnor U1296 (N_1296,N_1203,N_1265);
nor U1297 (N_1297,N_1222,N_1274);
xor U1298 (N_1298,N_1235,N_1202);
and U1299 (N_1299,N_1259,N_1212);
nor U1300 (N_1300,N_1223,N_1211);
nor U1301 (N_1301,N_1237,N_1216);
nand U1302 (N_1302,N_1228,N_1245);
xor U1303 (N_1303,N_1261,N_1205);
or U1304 (N_1304,N_1206,N_1239);
or U1305 (N_1305,N_1233,N_1214);
nor U1306 (N_1306,N_1225,N_1247);
nand U1307 (N_1307,N_1215,N_1201);
or U1308 (N_1308,N_1220,N_1231);
nor U1309 (N_1309,N_1241,N_1270);
nor U1310 (N_1310,N_1256,N_1267);
or U1311 (N_1311,N_1255,N_1210);
or U1312 (N_1312,N_1221,N_1238);
xor U1313 (N_1313,N_1264,N_1203);
and U1314 (N_1314,N_1219,N_1261);
nor U1315 (N_1315,N_1216,N_1201);
and U1316 (N_1316,N_1213,N_1256);
nand U1317 (N_1317,N_1202,N_1237);
xnor U1318 (N_1318,N_1258,N_1233);
or U1319 (N_1319,N_1262,N_1213);
xor U1320 (N_1320,N_1269,N_1217);
nand U1321 (N_1321,N_1257,N_1240);
nand U1322 (N_1322,N_1237,N_1273);
or U1323 (N_1323,N_1250,N_1228);
nand U1324 (N_1324,N_1250,N_1264);
or U1325 (N_1325,N_1226,N_1253);
or U1326 (N_1326,N_1249,N_1264);
xnor U1327 (N_1327,N_1230,N_1225);
and U1328 (N_1328,N_1263,N_1235);
xor U1329 (N_1329,N_1249,N_1237);
nor U1330 (N_1330,N_1237,N_1212);
and U1331 (N_1331,N_1270,N_1200);
nor U1332 (N_1332,N_1221,N_1218);
nand U1333 (N_1333,N_1224,N_1248);
or U1334 (N_1334,N_1219,N_1233);
xnor U1335 (N_1335,N_1204,N_1248);
or U1336 (N_1336,N_1240,N_1213);
nand U1337 (N_1337,N_1234,N_1265);
or U1338 (N_1338,N_1247,N_1219);
nor U1339 (N_1339,N_1218,N_1259);
and U1340 (N_1340,N_1232,N_1268);
and U1341 (N_1341,N_1206,N_1227);
and U1342 (N_1342,N_1224,N_1250);
nor U1343 (N_1343,N_1222,N_1250);
nor U1344 (N_1344,N_1240,N_1246);
or U1345 (N_1345,N_1216,N_1240);
nand U1346 (N_1346,N_1241,N_1218);
nand U1347 (N_1347,N_1219,N_1210);
and U1348 (N_1348,N_1268,N_1201);
and U1349 (N_1349,N_1259,N_1247);
xor U1350 (N_1350,N_1295,N_1302);
xnor U1351 (N_1351,N_1313,N_1315);
and U1352 (N_1352,N_1312,N_1342);
or U1353 (N_1353,N_1277,N_1317);
and U1354 (N_1354,N_1328,N_1314);
nand U1355 (N_1355,N_1292,N_1300);
nor U1356 (N_1356,N_1288,N_1311);
nor U1357 (N_1357,N_1327,N_1289);
or U1358 (N_1358,N_1278,N_1275);
nor U1359 (N_1359,N_1337,N_1347);
xnor U1360 (N_1360,N_1299,N_1307);
xnor U1361 (N_1361,N_1285,N_1348);
nand U1362 (N_1362,N_1294,N_1304);
xor U1363 (N_1363,N_1301,N_1336);
and U1364 (N_1364,N_1343,N_1333);
nor U1365 (N_1365,N_1309,N_1284);
or U1366 (N_1366,N_1281,N_1310);
nor U1367 (N_1367,N_1344,N_1306);
nand U1368 (N_1368,N_1287,N_1282);
nor U1369 (N_1369,N_1279,N_1330);
nand U1370 (N_1370,N_1346,N_1325);
or U1371 (N_1371,N_1331,N_1276);
nand U1372 (N_1372,N_1323,N_1319);
or U1373 (N_1373,N_1349,N_1329);
or U1374 (N_1374,N_1283,N_1334);
and U1375 (N_1375,N_1320,N_1297);
or U1376 (N_1376,N_1296,N_1335);
nor U1377 (N_1377,N_1298,N_1316);
nand U1378 (N_1378,N_1326,N_1332);
nor U1379 (N_1379,N_1305,N_1291);
and U1380 (N_1380,N_1339,N_1290);
xor U1381 (N_1381,N_1318,N_1345);
or U1382 (N_1382,N_1324,N_1340);
nand U1383 (N_1383,N_1303,N_1286);
nand U1384 (N_1384,N_1321,N_1341);
nor U1385 (N_1385,N_1322,N_1280);
xnor U1386 (N_1386,N_1293,N_1338);
or U1387 (N_1387,N_1308,N_1340);
and U1388 (N_1388,N_1306,N_1313);
or U1389 (N_1389,N_1295,N_1301);
nand U1390 (N_1390,N_1342,N_1300);
nand U1391 (N_1391,N_1305,N_1318);
xnor U1392 (N_1392,N_1277,N_1345);
and U1393 (N_1393,N_1322,N_1297);
xnor U1394 (N_1394,N_1278,N_1297);
and U1395 (N_1395,N_1347,N_1289);
or U1396 (N_1396,N_1322,N_1328);
nor U1397 (N_1397,N_1341,N_1331);
or U1398 (N_1398,N_1310,N_1284);
xor U1399 (N_1399,N_1341,N_1308);
xor U1400 (N_1400,N_1293,N_1322);
nor U1401 (N_1401,N_1285,N_1337);
and U1402 (N_1402,N_1319,N_1309);
and U1403 (N_1403,N_1311,N_1314);
xor U1404 (N_1404,N_1315,N_1301);
nor U1405 (N_1405,N_1315,N_1287);
or U1406 (N_1406,N_1309,N_1288);
xnor U1407 (N_1407,N_1326,N_1337);
and U1408 (N_1408,N_1321,N_1331);
or U1409 (N_1409,N_1311,N_1286);
xor U1410 (N_1410,N_1312,N_1276);
nor U1411 (N_1411,N_1298,N_1302);
nor U1412 (N_1412,N_1290,N_1305);
and U1413 (N_1413,N_1301,N_1323);
nor U1414 (N_1414,N_1294,N_1332);
nor U1415 (N_1415,N_1320,N_1305);
nand U1416 (N_1416,N_1307,N_1348);
nor U1417 (N_1417,N_1348,N_1318);
and U1418 (N_1418,N_1319,N_1347);
nand U1419 (N_1419,N_1315,N_1337);
or U1420 (N_1420,N_1293,N_1324);
nor U1421 (N_1421,N_1335,N_1284);
xor U1422 (N_1422,N_1322,N_1343);
and U1423 (N_1423,N_1339,N_1345);
nand U1424 (N_1424,N_1308,N_1329);
xnor U1425 (N_1425,N_1408,N_1379);
xnor U1426 (N_1426,N_1352,N_1364);
or U1427 (N_1427,N_1413,N_1367);
nand U1428 (N_1428,N_1392,N_1383);
or U1429 (N_1429,N_1409,N_1400);
or U1430 (N_1430,N_1376,N_1398);
nand U1431 (N_1431,N_1412,N_1422);
xnor U1432 (N_1432,N_1380,N_1378);
or U1433 (N_1433,N_1423,N_1401);
and U1434 (N_1434,N_1365,N_1357);
nand U1435 (N_1435,N_1411,N_1350);
nand U1436 (N_1436,N_1419,N_1372);
nand U1437 (N_1437,N_1358,N_1388);
or U1438 (N_1438,N_1396,N_1390);
and U1439 (N_1439,N_1402,N_1362);
and U1440 (N_1440,N_1377,N_1394);
nand U1441 (N_1441,N_1366,N_1405);
or U1442 (N_1442,N_1355,N_1393);
nand U1443 (N_1443,N_1351,N_1374);
nand U1444 (N_1444,N_1387,N_1415);
nand U1445 (N_1445,N_1397,N_1418);
or U1446 (N_1446,N_1354,N_1421);
xnor U1447 (N_1447,N_1403,N_1407);
or U1448 (N_1448,N_1381,N_1404);
nand U1449 (N_1449,N_1370,N_1417);
nor U1450 (N_1450,N_1373,N_1359);
nand U1451 (N_1451,N_1414,N_1363);
or U1452 (N_1452,N_1420,N_1395);
nand U1453 (N_1453,N_1360,N_1386);
nor U1454 (N_1454,N_1389,N_1424);
xnor U1455 (N_1455,N_1368,N_1371);
or U1456 (N_1456,N_1375,N_1399);
or U1457 (N_1457,N_1385,N_1353);
xnor U1458 (N_1458,N_1361,N_1391);
and U1459 (N_1459,N_1416,N_1369);
and U1460 (N_1460,N_1406,N_1382);
or U1461 (N_1461,N_1356,N_1384);
xor U1462 (N_1462,N_1410,N_1415);
or U1463 (N_1463,N_1387,N_1372);
xor U1464 (N_1464,N_1402,N_1424);
or U1465 (N_1465,N_1359,N_1402);
or U1466 (N_1466,N_1373,N_1393);
nor U1467 (N_1467,N_1350,N_1414);
or U1468 (N_1468,N_1352,N_1408);
and U1469 (N_1469,N_1384,N_1373);
and U1470 (N_1470,N_1389,N_1360);
nor U1471 (N_1471,N_1392,N_1404);
and U1472 (N_1472,N_1408,N_1357);
nand U1473 (N_1473,N_1351,N_1391);
nand U1474 (N_1474,N_1419,N_1382);
xor U1475 (N_1475,N_1422,N_1391);
or U1476 (N_1476,N_1364,N_1350);
xor U1477 (N_1477,N_1362,N_1406);
xnor U1478 (N_1478,N_1403,N_1369);
xnor U1479 (N_1479,N_1380,N_1387);
xor U1480 (N_1480,N_1392,N_1365);
xor U1481 (N_1481,N_1352,N_1367);
and U1482 (N_1482,N_1405,N_1370);
and U1483 (N_1483,N_1394,N_1361);
and U1484 (N_1484,N_1410,N_1419);
and U1485 (N_1485,N_1424,N_1352);
nor U1486 (N_1486,N_1370,N_1407);
nand U1487 (N_1487,N_1359,N_1382);
nor U1488 (N_1488,N_1407,N_1360);
and U1489 (N_1489,N_1374,N_1369);
or U1490 (N_1490,N_1390,N_1364);
nand U1491 (N_1491,N_1397,N_1384);
nand U1492 (N_1492,N_1416,N_1423);
and U1493 (N_1493,N_1423,N_1377);
or U1494 (N_1494,N_1415,N_1356);
or U1495 (N_1495,N_1420,N_1373);
or U1496 (N_1496,N_1361,N_1384);
and U1497 (N_1497,N_1358,N_1369);
nand U1498 (N_1498,N_1407,N_1351);
nand U1499 (N_1499,N_1414,N_1386);
xnor U1500 (N_1500,N_1477,N_1496);
or U1501 (N_1501,N_1442,N_1430);
nand U1502 (N_1502,N_1440,N_1478);
or U1503 (N_1503,N_1476,N_1454);
or U1504 (N_1504,N_1475,N_1453);
and U1505 (N_1505,N_1469,N_1481);
and U1506 (N_1506,N_1494,N_1450);
nand U1507 (N_1507,N_1493,N_1433);
or U1508 (N_1508,N_1426,N_1480);
or U1509 (N_1509,N_1487,N_1467);
nand U1510 (N_1510,N_1439,N_1495);
xor U1511 (N_1511,N_1443,N_1465);
or U1512 (N_1512,N_1451,N_1436);
and U1513 (N_1513,N_1489,N_1459);
xnor U1514 (N_1514,N_1435,N_1437);
or U1515 (N_1515,N_1427,N_1457);
xor U1516 (N_1516,N_1448,N_1463);
or U1517 (N_1517,N_1470,N_1441);
and U1518 (N_1518,N_1483,N_1485);
or U1519 (N_1519,N_1446,N_1474);
or U1520 (N_1520,N_1492,N_1473);
xor U1521 (N_1521,N_1486,N_1462);
xor U1522 (N_1522,N_1499,N_1490);
and U1523 (N_1523,N_1449,N_1452);
nand U1524 (N_1524,N_1447,N_1491);
xnor U1525 (N_1525,N_1471,N_1432);
or U1526 (N_1526,N_1466,N_1456);
and U1527 (N_1527,N_1455,N_1488);
or U1528 (N_1528,N_1444,N_1458);
nand U1529 (N_1529,N_1464,N_1431);
or U1530 (N_1530,N_1479,N_1438);
and U1531 (N_1531,N_1498,N_1428);
nor U1532 (N_1532,N_1434,N_1425);
nand U1533 (N_1533,N_1468,N_1429);
and U1534 (N_1534,N_1445,N_1461);
and U1535 (N_1535,N_1472,N_1497);
nand U1536 (N_1536,N_1482,N_1460);
nor U1537 (N_1537,N_1484,N_1492);
and U1538 (N_1538,N_1458,N_1487);
nand U1539 (N_1539,N_1467,N_1474);
nor U1540 (N_1540,N_1473,N_1499);
nand U1541 (N_1541,N_1499,N_1454);
and U1542 (N_1542,N_1471,N_1469);
or U1543 (N_1543,N_1430,N_1449);
and U1544 (N_1544,N_1492,N_1480);
xor U1545 (N_1545,N_1430,N_1486);
xor U1546 (N_1546,N_1442,N_1493);
and U1547 (N_1547,N_1425,N_1494);
or U1548 (N_1548,N_1495,N_1479);
nand U1549 (N_1549,N_1498,N_1451);
xnor U1550 (N_1550,N_1456,N_1438);
or U1551 (N_1551,N_1437,N_1427);
xor U1552 (N_1552,N_1470,N_1440);
and U1553 (N_1553,N_1470,N_1483);
xnor U1554 (N_1554,N_1482,N_1434);
xnor U1555 (N_1555,N_1458,N_1496);
and U1556 (N_1556,N_1434,N_1456);
and U1557 (N_1557,N_1427,N_1473);
or U1558 (N_1558,N_1471,N_1459);
or U1559 (N_1559,N_1497,N_1473);
or U1560 (N_1560,N_1426,N_1449);
nor U1561 (N_1561,N_1445,N_1494);
nor U1562 (N_1562,N_1436,N_1499);
and U1563 (N_1563,N_1469,N_1433);
and U1564 (N_1564,N_1432,N_1490);
or U1565 (N_1565,N_1484,N_1488);
and U1566 (N_1566,N_1463,N_1437);
or U1567 (N_1567,N_1427,N_1493);
nand U1568 (N_1568,N_1493,N_1468);
and U1569 (N_1569,N_1425,N_1443);
nand U1570 (N_1570,N_1492,N_1425);
nor U1571 (N_1571,N_1438,N_1496);
and U1572 (N_1572,N_1487,N_1484);
and U1573 (N_1573,N_1435,N_1461);
and U1574 (N_1574,N_1489,N_1433);
or U1575 (N_1575,N_1514,N_1546);
xor U1576 (N_1576,N_1510,N_1571);
xor U1577 (N_1577,N_1517,N_1542);
xor U1578 (N_1578,N_1563,N_1520);
nand U1579 (N_1579,N_1513,N_1531);
and U1580 (N_1580,N_1512,N_1556);
and U1581 (N_1581,N_1565,N_1501);
and U1582 (N_1582,N_1516,N_1572);
nand U1583 (N_1583,N_1507,N_1547);
nand U1584 (N_1584,N_1552,N_1558);
nor U1585 (N_1585,N_1551,N_1557);
xor U1586 (N_1586,N_1555,N_1509);
and U1587 (N_1587,N_1529,N_1535);
xnor U1588 (N_1588,N_1527,N_1569);
or U1589 (N_1589,N_1523,N_1543);
nand U1590 (N_1590,N_1504,N_1519);
and U1591 (N_1591,N_1554,N_1518);
and U1592 (N_1592,N_1540,N_1532);
nor U1593 (N_1593,N_1526,N_1505);
or U1594 (N_1594,N_1506,N_1528);
or U1595 (N_1595,N_1574,N_1570);
nand U1596 (N_1596,N_1561,N_1524);
nor U1597 (N_1597,N_1573,N_1537);
and U1598 (N_1598,N_1559,N_1544);
nand U1599 (N_1599,N_1536,N_1525);
and U1600 (N_1600,N_1503,N_1502);
or U1601 (N_1601,N_1548,N_1500);
xor U1602 (N_1602,N_1553,N_1545);
or U1603 (N_1603,N_1549,N_1550);
nor U1604 (N_1604,N_1564,N_1508);
and U1605 (N_1605,N_1515,N_1539);
nor U1606 (N_1606,N_1534,N_1533);
and U1607 (N_1607,N_1568,N_1560);
and U1608 (N_1608,N_1522,N_1521);
and U1609 (N_1609,N_1566,N_1538);
or U1610 (N_1610,N_1530,N_1567);
nand U1611 (N_1611,N_1541,N_1562);
or U1612 (N_1612,N_1511,N_1549);
or U1613 (N_1613,N_1518,N_1511);
nand U1614 (N_1614,N_1506,N_1551);
xor U1615 (N_1615,N_1504,N_1540);
nor U1616 (N_1616,N_1566,N_1567);
nand U1617 (N_1617,N_1553,N_1505);
or U1618 (N_1618,N_1522,N_1568);
or U1619 (N_1619,N_1515,N_1507);
nand U1620 (N_1620,N_1505,N_1545);
or U1621 (N_1621,N_1566,N_1500);
nand U1622 (N_1622,N_1520,N_1524);
or U1623 (N_1623,N_1530,N_1504);
or U1624 (N_1624,N_1515,N_1500);
or U1625 (N_1625,N_1525,N_1559);
xor U1626 (N_1626,N_1540,N_1552);
and U1627 (N_1627,N_1505,N_1567);
nand U1628 (N_1628,N_1525,N_1568);
xor U1629 (N_1629,N_1571,N_1534);
xor U1630 (N_1630,N_1518,N_1514);
or U1631 (N_1631,N_1511,N_1522);
nor U1632 (N_1632,N_1539,N_1531);
or U1633 (N_1633,N_1560,N_1514);
xor U1634 (N_1634,N_1519,N_1550);
nand U1635 (N_1635,N_1560,N_1557);
xor U1636 (N_1636,N_1510,N_1542);
nand U1637 (N_1637,N_1523,N_1564);
and U1638 (N_1638,N_1544,N_1529);
xnor U1639 (N_1639,N_1553,N_1541);
or U1640 (N_1640,N_1574,N_1554);
nor U1641 (N_1641,N_1543,N_1565);
nor U1642 (N_1642,N_1515,N_1560);
xnor U1643 (N_1643,N_1526,N_1568);
nor U1644 (N_1644,N_1511,N_1555);
nand U1645 (N_1645,N_1552,N_1569);
nand U1646 (N_1646,N_1540,N_1522);
or U1647 (N_1647,N_1525,N_1508);
xnor U1648 (N_1648,N_1532,N_1518);
or U1649 (N_1649,N_1552,N_1539);
xnor U1650 (N_1650,N_1589,N_1636);
xnor U1651 (N_1651,N_1594,N_1579);
nand U1652 (N_1652,N_1611,N_1614);
nand U1653 (N_1653,N_1647,N_1595);
xnor U1654 (N_1654,N_1605,N_1646);
or U1655 (N_1655,N_1616,N_1582);
and U1656 (N_1656,N_1597,N_1584);
or U1657 (N_1657,N_1604,N_1612);
nor U1658 (N_1658,N_1634,N_1613);
nand U1659 (N_1659,N_1644,N_1576);
xor U1660 (N_1660,N_1619,N_1588);
or U1661 (N_1661,N_1580,N_1607);
or U1662 (N_1662,N_1641,N_1640);
or U1663 (N_1663,N_1591,N_1601);
and U1664 (N_1664,N_1585,N_1625);
or U1665 (N_1665,N_1575,N_1583);
or U1666 (N_1666,N_1639,N_1621);
nor U1667 (N_1667,N_1578,N_1623);
and U1668 (N_1668,N_1627,N_1609);
nand U1669 (N_1669,N_1628,N_1610);
nor U1670 (N_1670,N_1596,N_1630);
or U1671 (N_1671,N_1586,N_1581);
nor U1672 (N_1672,N_1631,N_1617);
xnor U1673 (N_1673,N_1608,N_1590);
nor U1674 (N_1674,N_1632,N_1645);
xor U1675 (N_1675,N_1642,N_1577);
and U1676 (N_1676,N_1620,N_1635);
and U1677 (N_1677,N_1587,N_1629);
or U1678 (N_1678,N_1592,N_1626);
nand U1679 (N_1679,N_1643,N_1600);
xor U1680 (N_1680,N_1615,N_1622);
and U1681 (N_1681,N_1602,N_1593);
nor U1682 (N_1682,N_1598,N_1649);
nor U1683 (N_1683,N_1603,N_1618);
nand U1684 (N_1684,N_1599,N_1606);
and U1685 (N_1685,N_1637,N_1638);
and U1686 (N_1686,N_1633,N_1624);
nor U1687 (N_1687,N_1648,N_1614);
nand U1688 (N_1688,N_1626,N_1587);
nor U1689 (N_1689,N_1642,N_1620);
and U1690 (N_1690,N_1642,N_1643);
and U1691 (N_1691,N_1642,N_1582);
nand U1692 (N_1692,N_1584,N_1626);
or U1693 (N_1693,N_1642,N_1589);
xor U1694 (N_1694,N_1588,N_1575);
or U1695 (N_1695,N_1599,N_1578);
nor U1696 (N_1696,N_1575,N_1598);
nor U1697 (N_1697,N_1622,N_1610);
or U1698 (N_1698,N_1628,N_1639);
nand U1699 (N_1699,N_1607,N_1645);
xnor U1700 (N_1700,N_1632,N_1589);
xnor U1701 (N_1701,N_1597,N_1618);
nand U1702 (N_1702,N_1634,N_1592);
xor U1703 (N_1703,N_1624,N_1626);
nand U1704 (N_1704,N_1596,N_1602);
or U1705 (N_1705,N_1595,N_1619);
nor U1706 (N_1706,N_1605,N_1603);
and U1707 (N_1707,N_1585,N_1640);
nand U1708 (N_1708,N_1641,N_1580);
and U1709 (N_1709,N_1611,N_1642);
and U1710 (N_1710,N_1629,N_1642);
nand U1711 (N_1711,N_1589,N_1648);
and U1712 (N_1712,N_1595,N_1648);
or U1713 (N_1713,N_1591,N_1589);
or U1714 (N_1714,N_1631,N_1609);
xnor U1715 (N_1715,N_1633,N_1645);
or U1716 (N_1716,N_1626,N_1579);
and U1717 (N_1717,N_1602,N_1594);
nand U1718 (N_1718,N_1627,N_1596);
nand U1719 (N_1719,N_1625,N_1611);
or U1720 (N_1720,N_1641,N_1583);
nand U1721 (N_1721,N_1628,N_1577);
xnor U1722 (N_1722,N_1640,N_1575);
xnor U1723 (N_1723,N_1585,N_1617);
nand U1724 (N_1724,N_1602,N_1629);
or U1725 (N_1725,N_1671,N_1678);
and U1726 (N_1726,N_1652,N_1659);
or U1727 (N_1727,N_1670,N_1687);
nand U1728 (N_1728,N_1677,N_1718);
nor U1729 (N_1729,N_1719,N_1656);
or U1730 (N_1730,N_1667,N_1674);
or U1731 (N_1731,N_1658,N_1710);
or U1732 (N_1732,N_1686,N_1688);
xor U1733 (N_1733,N_1682,N_1693);
and U1734 (N_1734,N_1654,N_1661);
and U1735 (N_1735,N_1698,N_1657);
and U1736 (N_1736,N_1723,N_1714);
nor U1737 (N_1737,N_1692,N_1707);
nand U1738 (N_1738,N_1664,N_1653);
nor U1739 (N_1739,N_1669,N_1651);
and U1740 (N_1740,N_1720,N_1666);
xor U1741 (N_1741,N_1662,N_1706);
or U1742 (N_1742,N_1668,N_1684);
and U1743 (N_1743,N_1650,N_1694);
and U1744 (N_1744,N_1665,N_1679);
nand U1745 (N_1745,N_1655,N_1663);
nand U1746 (N_1746,N_1713,N_1675);
xor U1747 (N_1747,N_1709,N_1700);
nor U1748 (N_1748,N_1695,N_1691);
or U1749 (N_1749,N_1685,N_1673);
nor U1750 (N_1750,N_1681,N_1711);
nor U1751 (N_1751,N_1708,N_1676);
nand U1752 (N_1752,N_1712,N_1715);
xnor U1753 (N_1753,N_1672,N_1697);
xnor U1754 (N_1754,N_1716,N_1680);
or U1755 (N_1755,N_1703,N_1690);
or U1756 (N_1756,N_1724,N_1702);
or U1757 (N_1757,N_1701,N_1722);
and U1758 (N_1758,N_1683,N_1704);
or U1759 (N_1759,N_1660,N_1689);
nor U1760 (N_1760,N_1696,N_1699);
nand U1761 (N_1761,N_1717,N_1721);
or U1762 (N_1762,N_1705,N_1693);
and U1763 (N_1763,N_1691,N_1715);
nor U1764 (N_1764,N_1718,N_1708);
nand U1765 (N_1765,N_1670,N_1684);
nand U1766 (N_1766,N_1701,N_1724);
and U1767 (N_1767,N_1724,N_1689);
xnor U1768 (N_1768,N_1664,N_1716);
xor U1769 (N_1769,N_1660,N_1665);
xor U1770 (N_1770,N_1670,N_1652);
nor U1771 (N_1771,N_1670,N_1721);
and U1772 (N_1772,N_1691,N_1671);
xnor U1773 (N_1773,N_1706,N_1688);
nand U1774 (N_1774,N_1657,N_1665);
or U1775 (N_1775,N_1712,N_1658);
nor U1776 (N_1776,N_1724,N_1686);
and U1777 (N_1777,N_1710,N_1699);
nor U1778 (N_1778,N_1711,N_1669);
and U1779 (N_1779,N_1705,N_1664);
nor U1780 (N_1780,N_1715,N_1714);
xnor U1781 (N_1781,N_1711,N_1697);
xnor U1782 (N_1782,N_1720,N_1665);
xnor U1783 (N_1783,N_1679,N_1652);
xor U1784 (N_1784,N_1668,N_1687);
or U1785 (N_1785,N_1680,N_1722);
xor U1786 (N_1786,N_1692,N_1702);
or U1787 (N_1787,N_1661,N_1708);
nor U1788 (N_1788,N_1696,N_1655);
nor U1789 (N_1789,N_1693,N_1655);
nand U1790 (N_1790,N_1692,N_1665);
nor U1791 (N_1791,N_1658,N_1708);
and U1792 (N_1792,N_1701,N_1702);
and U1793 (N_1793,N_1691,N_1705);
xnor U1794 (N_1794,N_1723,N_1672);
or U1795 (N_1795,N_1653,N_1718);
xor U1796 (N_1796,N_1718,N_1687);
nor U1797 (N_1797,N_1716,N_1677);
nor U1798 (N_1798,N_1712,N_1721);
nor U1799 (N_1799,N_1702,N_1720);
nor U1800 (N_1800,N_1767,N_1782);
xnor U1801 (N_1801,N_1744,N_1752);
or U1802 (N_1802,N_1793,N_1764);
and U1803 (N_1803,N_1780,N_1751);
and U1804 (N_1804,N_1753,N_1762);
xnor U1805 (N_1805,N_1742,N_1745);
xor U1806 (N_1806,N_1772,N_1775);
and U1807 (N_1807,N_1786,N_1741);
and U1808 (N_1808,N_1787,N_1788);
xnor U1809 (N_1809,N_1795,N_1779);
xnor U1810 (N_1810,N_1784,N_1728);
nand U1811 (N_1811,N_1765,N_1774);
nand U1812 (N_1812,N_1794,N_1732);
nand U1813 (N_1813,N_1730,N_1733);
and U1814 (N_1814,N_1769,N_1799);
xnor U1815 (N_1815,N_1785,N_1760);
xnor U1816 (N_1816,N_1778,N_1796);
or U1817 (N_1817,N_1798,N_1727);
nand U1818 (N_1818,N_1743,N_1726);
nor U1819 (N_1819,N_1725,N_1759);
or U1820 (N_1820,N_1781,N_1729);
nor U1821 (N_1821,N_1761,N_1768);
nand U1822 (N_1822,N_1792,N_1746);
xnor U1823 (N_1823,N_1758,N_1749);
nand U1824 (N_1824,N_1739,N_1731);
nor U1825 (N_1825,N_1763,N_1770);
and U1826 (N_1826,N_1776,N_1735);
nor U1827 (N_1827,N_1756,N_1757);
xnor U1828 (N_1828,N_1773,N_1771);
xnor U1829 (N_1829,N_1766,N_1777);
xnor U1830 (N_1830,N_1755,N_1736);
nor U1831 (N_1831,N_1748,N_1790);
xnor U1832 (N_1832,N_1747,N_1797);
and U1833 (N_1833,N_1734,N_1750);
or U1834 (N_1834,N_1789,N_1740);
nor U1835 (N_1835,N_1738,N_1791);
nand U1836 (N_1836,N_1737,N_1754);
and U1837 (N_1837,N_1783,N_1765);
xnor U1838 (N_1838,N_1757,N_1747);
or U1839 (N_1839,N_1780,N_1745);
nor U1840 (N_1840,N_1774,N_1748);
and U1841 (N_1841,N_1759,N_1763);
xor U1842 (N_1842,N_1725,N_1765);
nor U1843 (N_1843,N_1781,N_1727);
nand U1844 (N_1844,N_1774,N_1796);
nand U1845 (N_1845,N_1734,N_1785);
or U1846 (N_1846,N_1761,N_1786);
nand U1847 (N_1847,N_1759,N_1735);
and U1848 (N_1848,N_1783,N_1788);
nor U1849 (N_1849,N_1792,N_1738);
and U1850 (N_1850,N_1742,N_1775);
nor U1851 (N_1851,N_1794,N_1738);
or U1852 (N_1852,N_1772,N_1780);
nand U1853 (N_1853,N_1798,N_1784);
nor U1854 (N_1854,N_1785,N_1755);
and U1855 (N_1855,N_1764,N_1728);
nand U1856 (N_1856,N_1753,N_1798);
nor U1857 (N_1857,N_1752,N_1730);
xor U1858 (N_1858,N_1740,N_1741);
xnor U1859 (N_1859,N_1786,N_1746);
xnor U1860 (N_1860,N_1738,N_1776);
xnor U1861 (N_1861,N_1778,N_1748);
or U1862 (N_1862,N_1785,N_1773);
and U1863 (N_1863,N_1791,N_1733);
nor U1864 (N_1864,N_1794,N_1790);
or U1865 (N_1865,N_1774,N_1781);
xnor U1866 (N_1866,N_1772,N_1735);
or U1867 (N_1867,N_1727,N_1792);
or U1868 (N_1868,N_1766,N_1748);
or U1869 (N_1869,N_1760,N_1728);
xnor U1870 (N_1870,N_1736,N_1782);
xnor U1871 (N_1871,N_1750,N_1744);
xor U1872 (N_1872,N_1799,N_1760);
or U1873 (N_1873,N_1744,N_1788);
xnor U1874 (N_1874,N_1759,N_1762);
xor U1875 (N_1875,N_1871,N_1831);
nand U1876 (N_1876,N_1813,N_1834);
nor U1877 (N_1877,N_1863,N_1818);
nand U1878 (N_1878,N_1809,N_1801);
and U1879 (N_1879,N_1859,N_1843);
and U1880 (N_1880,N_1830,N_1869);
or U1881 (N_1881,N_1815,N_1873);
or U1882 (N_1882,N_1825,N_1838);
nor U1883 (N_1883,N_1807,N_1864);
or U1884 (N_1884,N_1816,N_1829);
nand U1885 (N_1885,N_1841,N_1865);
or U1886 (N_1886,N_1861,N_1828);
and U1887 (N_1887,N_1839,N_1802);
nand U1888 (N_1888,N_1845,N_1858);
xor U1889 (N_1889,N_1857,N_1814);
and U1890 (N_1890,N_1808,N_1819);
or U1891 (N_1891,N_1862,N_1851);
nand U1892 (N_1892,N_1804,N_1817);
nor U1893 (N_1893,N_1870,N_1811);
nand U1894 (N_1894,N_1849,N_1822);
nand U1895 (N_1895,N_1847,N_1840);
or U1896 (N_1896,N_1852,N_1850);
and U1897 (N_1897,N_1835,N_1867);
nand U1898 (N_1898,N_1836,N_1827);
nor U1899 (N_1899,N_1868,N_1826);
nand U1900 (N_1900,N_1805,N_1856);
nand U1901 (N_1901,N_1832,N_1848);
xnor U1902 (N_1902,N_1833,N_1860);
nand U1903 (N_1903,N_1842,N_1806);
xnor U1904 (N_1904,N_1855,N_1821);
nor U1905 (N_1905,N_1844,N_1824);
nand U1906 (N_1906,N_1820,N_1803);
and U1907 (N_1907,N_1874,N_1837);
or U1908 (N_1908,N_1810,N_1853);
nand U1909 (N_1909,N_1800,N_1866);
or U1910 (N_1910,N_1854,N_1812);
and U1911 (N_1911,N_1846,N_1872);
xnor U1912 (N_1912,N_1823,N_1868);
and U1913 (N_1913,N_1829,N_1855);
nand U1914 (N_1914,N_1837,N_1842);
nand U1915 (N_1915,N_1809,N_1838);
nand U1916 (N_1916,N_1846,N_1854);
nand U1917 (N_1917,N_1846,N_1858);
and U1918 (N_1918,N_1873,N_1830);
or U1919 (N_1919,N_1804,N_1865);
and U1920 (N_1920,N_1841,N_1846);
or U1921 (N_1921,N_1845,N_1809);
nand U1922 (N_1922,N_1830,N_1868);
nor U1923 (N_1923,N_1812,N_1850);
nor U1924 (N_1924,N_1808,N_1854);
xnor U1925 (N_1925,N_1847,N_1802);
xnor U1926 (N_1926,N_1834,N_1843);
xor U1927 (N_1927,N_1859,N_1836);
xor U1928 (N_1928,N_1870,N_1824);
nand U1929 (N_1929,N_1821,N_1850);
and U1930 (N_1930,N_1843,N_1845);
xor U1931 (N_1931,N_1852,N_1831);
nor U1932 (N_1932,N_1863,N_1861);
or U1933 (N_1933,N_1865,N_1864);
nor U1934 (N_1934,N_1802,N_1855);
nand U1935 (N_1935,N_1801,N_1836);
nor U1936 (N_1936,N_1848,N_1854);
and U1937 (N_1937,N_1872,N_1819);
nand U1938 (N_1938,N_1838,N_1812);
and U1939 (N_1939,N_1851,N_1847);
nor U1940 (N_1940,N_1825,N_1870);
nor U1941 (N_1941,N_1805,N_1813);
or U1942 (N_1942,N_1811,N_1831);
and U1943 (N_1943,N_1831,N_1862);
nand U1944 (N_1944,N_1849,N_1862);
nor U1945 (N_1945,N_1844,N_1864);
and U1946 (N_1946,N_1827,N_1855);
or U1947 (N_1947,N_1851,N_1800);
nor U1948 (N_1948,N_1822,N_1852);
or U1949 (N_1949,N_1819,N_1839);
nor U1950 (N_1950,N_1916,N_1913);
and U1951 (N_1951,N_1879,N_1897);
nand U1952 (N_1952,N_1889,N_1906);
nand U1953 (N_1953,N_1904,N_1895);
and U1954 (N_1954,N_1898,N_1915);
and U1955 (N_1955,N_1943,N_1885);
or U1956 (N_1956,N_1890,N_1942);
xnor U1957 (N_1957,N_1903,N_1918);
and U1958 (N_1958,N_1937,N_1912);
nand U1959 (N_1959,N_1922,N_1930);
nor U1960 (N_1960,N_1934,N_1945);
or U1961 (N_1961,N_1907,N_1938);
nand U1962 (N_1962,N_1936,N_1923);
or U1963 (N_1963,N_1900,N_1917);
xnor U1964 (N_1964,N_1928,N_1944);
and U1965 (N_1965,N_1909,N_1925);
or U1966 (N_1966,N_1876,N_1947);
and U1967 (N_1967,N_1935,N_1882);
and U1968 (N_1968,N_1888,N_1941);
xnor U1969 (N_1969,N_1878,N_1931);
or U1970 (N_1970,N_1948,N_1908);
xor U1971 (N_1971,N_1881,N_1896);
and U1972 (N_1972,N_1884,N_1883);
and U1973 (N_1973,N_1927,N_1880);
nand U1974 (N_1974,N_1946,N_1919);
xnor U1975 (N_1975,N_1893,N_1902);
xnor U1976 (N_1976,N_1894,N_1887);
and U1977 (N_1977,N_1921,N_1892);
and U1978 (N_1978,N_1929,N_1932);
and U1979 (N_1979,N_1926,N_1899);
nor U1980 (N_1980,N_1933,N_1875);
nand U1981 (N_1981,N_1939,N_1901);
and U1982 (N_1982,N_1891,N_1910);
xor U1983 (N_1983,N_1886,N_1924);
nor U1984 (N_1984,N_1914,N_1920);
xor U1985 (N_1985,N_1949,N_1940);
or U1986 (N_1986,N_1911,N_1905);
and U1987 (N_1987,N_1877,N_1893);
nor U1988 (N_1988,N_1937,N_1930);
and U1989 (N_1989,N_1920,N_1912);
and U1990 (N_1990,N_1916,N_1897);
nand U1991 (N_1991,N_1912,N_1906);
xnor U1992 (N_1992,N_1933,N_1930);
or U1993 (N_1993,N_1896,N_1922);
nand U1994 (N_1994,N_1901,N_1905);
or U1995 (N_1995,N_1906,N_1895);
nand U1996 (N_1996,N_1910,N_1926);
nor U1997 (N_1997,N_1878,N_1912);
nand U1998 (N_1998,N_1908,N_1916);
xnor U1999 (N_1999,N_1879,N_1941);
nor U2000 (N_2000,N_1891,N_1939);
nor U2001 (N_2001,N_1892,N_1947);
and U2002 (N_2002,N_1942,N_1940);
nor U2003 (N_2003,N_1879,N_1906);
and U2004 (N_2004,N_1942,N_1900);
nor U2005 (N_2005,N_1878,N_1909);
or U2006 (N_2006,N_1895,N_1908);
and U2007 (N_2007,N_1905,N_1939);
or U2008 (N_2008,N_1884,N_1942);
nor U2009 (N_2009,N_1946,N_1905);
nor U2010 (N_2010,N_1890,N_1947);
nand U2011 (N_2011,N_1947,N_1904);
xnor U2012 (N_2012,N_1895,N_1935);
nor U2013 (N_2013,N_1909,N_1880);
nor U2014 (N_2014,N_1880,N_1912);
or U2015 (N_2015,N_1889,N_1938);
nand U2016 (N_2016,N_1937,N_1889);
or U2017 (N_2017,N_1949,N_1947);
xor U2018 (N_2018,N_1882,N_1891);
and U2019 (N_2019,N_1933,N_1884);
and U2020 (N_2020,N_1922,N_1935);
nand U2021 (N_2021,N_1941,N_1897);
nand U2022 (N_2022,N_1906,N_1936);
xor U2023 (N_2023,N_1942,N_1923);
and U2024 (N_2024,N_1893,N_1925);
nand U2025 (N_2025,N_1977,N_1980);
or U2026 (N_2026,N_1990,N_1955);
nor U2027 (N_2027,N_1964,N_2012);
and U2028 (N_2028,N_1981,N_1963);
nor U2029 (N_2029,N_1973,N_1966);
nor U2030 (N_2030,N_1959,N_1952);
nor U2031 (N_2031,N_1988,N_1951);
and U2032 (N_2032,N_2003,N_1953);
nand U2033 (N_2033,N_2006,N_1972);
or U2034 (N_2034,N_2021,N_2001);
and U2035 (N_2035,N_1995,N_2011);
and U2036 (N_2036,N_1956,N_2013);
and U2037 (N_2037,N_1994,N_2015);
or U2038 (N_2038,N_1984,N_1958);
or U2039 (N_2039,N_1986,N_2007);
xor U2040 (N_2040,N_1967,N_1975);
nor U2041 (N_2041,N_2023,N_1987);
xor U2042 (N_2042,N_1982,N_1971);
xor U2043 (N_2043,N_1961,N_2024);
and U2044 (N_2044,N_1965,N_2019);
and U2045 (N_2045,N_1991,N_1999);
xor U2046 (N_2046,N_1993,N_1997);
and U2047 (N_2047,N_2009,N_1962);
nor U2048 (N_2048,N_2002,N_2004);
or U2049 (N_2049,N_1969,N_2016);
xnor U2050 (N_2050,N_1985,N_2000);
nand U2051 (N_2051,N_1979,N_2014);
nor U2052 (N_2052,N_1989,N_1970);
and U2053 (N_2053,N_1954,N_1998);
nand U2054 (N_2054,N_1974,N_2020);
nand U2055 (N_2055,N_2008,N_1957);
and U2056 (N_2056,N_1960,N_2017);
or U2057 (N_2057,N_1976,N_1996);
and U2058 (N_2058,N_1950,N_1968);
and U2059 (N_2059,N_2005,N_1983);
nor U2060 (N_2060,N_1992,N_2022);
nor U2061 (N_2061,N_2010,N_2018);
or U2062 (N_2062,N_1978,N_2005);
xor U2063 (N_2063,N_2011,N_2019);
and U2064 (N_2064,N_1985,N_2019);
or U2065 (N_2065,N_1972,N_1989);
or U2066 (N_2066,N_1992,N_2021);
nor U2067 (N_2067,N_2021,N_2024);
xor U2068 (N_2068,N_1965,N_1978);
xnor U2069 (N_2069,N_2013,N_2002);
nor U2070 (N_2070,N_2019,N_1993);
nand U2071 (N_2071,N_1990,N_1999);
and U2072 (N_2072,N_1969,N_1985);
or U2073 (N_2073,N_1991,N_1981);
xnor U2074 (N_2074,N_1984,N_1954);
nor U2075 (N_2075,N_2000,N_1964);
nand U2076 (N_2076,N_1997,N_2000);
nand U2077 (N_2077,N_2022,N_2003);
or U2078 (N_2078,N_1954,N_2023);
nor U2079 (N_2079,N_2020,N_1999);
or U2080 (N_2080,N_1998,N_1961);
or U2081 (N_2081,N_2023,N_1955);
or U2082 (N_2082,N_2024,N_1990);
xor U2083 (N_2083,N_1966,N_1968);
xnor U2084 (N_2084,N_2022,N_2011);
or U2085 (N_2085,N_1988,N_2004);
and U2086 (N_2086,N_1991,N_1954);
xnor U2087 (N_2087,N_1957,N_1986);
nor U2088 (N_2088,N_1977,N_1965);
or U2089 (N_2089,N_1975,N_1953);
xnor U2090 (N_2090,N_1979,N_1956);
or U2091 (N_2091,N_1965,N_2000);
nor U2092 (N_2092,N_1952,N_2018);
nor U2093 (N_2093,N_1979,N_1993);
nor U2094 (N_2094,N_2019,N_2006);
nand U2095 (N_2095,N_2017,N_1996);
nor U2096 (N_2096,N_2003,N_1984);
and U2097 (N_2097,N_1962,N_1952);
nor U2098 (N_2098,N_1998,N_2006);
nor U2099 (N_2099,N_2012,N_1951);
nor U2100 (N_2100,N_2035,N_2075);
nor U2101 (N_2101,N_2031,N_2038);
nor U2102 (N_2102,N_2036,N_2065);
and U2103 (N_2103,N_2071,N_2048);
xnor U2104 (N_2104,N_2053,N_2044);
xor U2105 (N_2105,N_2083,N_2033);
xnor U2106 (N_2106,N_2052,N_2042);
nor U2107 (N_2107,N_2094,N_2077);
xor U2108 (N_2108,N_2080,N_2059);
or U2109 (N_2109,N_2051,N_2086);
or U2110 (N_2110,N_2078,N_2058);
and U2111 (N_2111,N_2067,N_2090);
nand U2112 (N_2112,N_2027,N_2064);
or U2113 (N_2113,N_2081,N_2054);
and U2114 (N_2114,N_2096,N_2028);
nand U2115 (N_2115,N_2062,N_2049);
or U2116 (N_2116,N_2088,N_2092);
or U2117 (N_2117,N_2050,N_2073);
and U2118 (N_2118,N_2082,N_2074);
xor U2119 (N_2119,N_2057,N_2056);
or U2120 (N_2120,N_2084,N_2060);
nor U2121 (N_2121,N_2046,N_2095);
xnor U2122 (N_2122,N_2040,N_2087);
xor U2123 (N_2123,N_2032,N_2025);
nand U2124 (N_2124,N_2070,N_2066);
nand U2125 (N_2125,N_2097,N_2037);
and U2126 (N_2126,N_2063,N_2034);
nand U2127 (N_2127,N_2093,N_2072);
and U2128 (N_2128,N_2047,N_2043);
and U2129 (N_2129,N_2061,N_2045);
and U2130 (N_2130,N_2041,N_2039);
nand U2131 (N_2131,N_2069,N_2099);
nor U2132 (N_2132,N_2085,N_2098);
or U2133 (N_2133,N_2091,N_2076);
nand U2134 (N_2134,N_2068,N_2055);
nand U2135 (N_2135,N_2026,N_2089);
nor U2136 (N_2136,N_2079,N_2030);
nor U2137 (N_2137,N_2029,N_2092);
and U2138 (N_2138,N_2057,N_2034);
and U2139 (N_2139,N_2072,N_2096);
nor U2140 (N_2140,N_2095,N_2040);
nand U2141 (N_2141,N_2074,N_2099);
or U2142 (N_2142,N_2089,N_2077);
and U2143 (N_2143,N_2037,N_2043);
nand U2144 (N_2144,N_2080,N_2097);
nand U2145 (N_2145,N_2039,N_2025);
or U2146 (N_2146,N_2032,N_2038);
nand U2147 (N_2147,N_2067,N_2060);
nor U2148 (N_2148,N_2080,N_2085);
nor U2149 (N_2149,N_2057,N_2065);
xnor U2150 (N_2150,N_2081,N_2090);
xor U2151 (N_2151,N_2053,N_2051);
nand U2152 (N_2152,N_2077,N_2099);
nand U2153 (N_2153,N_2098,N_2065);
and U2154 (N_2154,N_2063,N_2096);
and U2155 (N_2155,N_2031,N_2042);
xor U2156 (N_2156,N_2046,N_2088);
and U2157 (N_2157,N_2056,N_2034);
and U2158 (N_2158,N_2076,N_2052);
and U2159 (N_2159,N_2025,N_2076);
nand U2160 (N_2160,N_2097,N_2098);
xnor U2161 (N_2161,N_2051,N_2060);
xnor U2162 (N_2162,N_2063,N_2077);
nor U2163 (N_2163,N_2026,N_2099);
and U2164 (N_2164,N_2028,N_2064);
nor U2165 (N_2165,N_2085,N_2042);
and U2166 (N_2166,N_2070,N_2085);
nand U2167 (N_2167,N_2073,N_2062);
xnor U2168 (N_2168,N_2065,N_2064);
or U2169 (N_2169,N_2085,N_2064);
or U2170 (N_2170,N_2046,N_2045);
and U2171 (N_2171,N_2061,N_2033);
nor U2172 (N_2172,N_2070,N_2050);
and U2173 (N_2173,N_2071,N_2087);
nand U2174 (N_2174,N_2086,N_2036);
nor U2175 (N_2175,N_2173,N_2161);
xor U2176 (N_2176,N_2116,N_2110);
nand U2177 (N_2177,N_2144,N_2106);
or U2178 (N_2178,N_2101,N_2103);
xnor U2179 (N_2179,N_2167,N_2147);
nand U2180 (N_2180,N_2156,N_2138);
and U2181 (N_2181,N_2166,N_2107);
nand U2182 (N_2182,N_2109,N_2108);
or U2183 (N_2183,N_2100,N_2131);
nand U2184 (N_2184,N_2158,N_2150);
or U2185 (N_2185,N_2142,N_2117);
or U2186 (N_2186,N_2136,N_2149);
xor U2187 (N_2187,N_2134,N_2132);
xor U2188 (N_2188,N_2137,N_2130);
or U2189 (N_2189,N_2174,N_2171);
xor U2190 (N_2190,N_2160,N_2129);
nor U2191 (N_2191,N_2140,N_2157);
or U2192 (N_2192,N_2169,N_2124);
xnor U2193 (N_2193,N_2152,N_2154);
or U2194 (N_2194,N_2135,N_2120);
and U2195 (N_2195,N_2115,N_2112);
nand U2196 (N_2196,N_2126,N_2141);
or U2197 (N_2197,N_2164,N_2143);
xnor U2198 (N_2198,N_2121,N_2148);
nor U2199 (N_2199,N_2139,N_2163);
nand U2200 (N_2200,N_2127,N_2170);
nor U2201 (N_2201,N_2122,N_2172);
or U2202 (N_2202,N_2125,N_2153);
xnor U2203 (N_2203,N_2102,N_2159);
xor U2204 (N_2204,N_2119,N_2118);
nand U2205 (N_2205,N_2151,N_2146);
nor U2206 (N_2206,N_2104,N_2114);
or U2207 (N_2207,N_2105,N_2155);
nand U2208 (N_2208,N_2145,N_2165);
or U2209 (N_2209,N_2123,N_2133);
and U2210 (N_2210,N_2162,N_2168);
or U2211 (N_2211,N_2128,N_2113);
nand U2212 (N_2212,N_2111,N_2170);
xor U2213 (N_2213,N_2117,N_2140);
nand U2214 (N_2214,N_2125,N_2156);
xnor U2215 (N_2215,N_2108,N_2125);
nor U2216 (N_2216,N_2125,N_2147);
and U2217 (N_2217,N_2106,N_2140);
xnor U2218 (N_2218,N_2134,N_2136);
and U2219 (N_2219,N_2107,N_2125);
nor U2220 (N_2220,N_2156,N_2152);
nand U2221 (N_2221,N_2134,N_2115);
xnor U2222 (N_2222,N_2156,N_2163);
nor U2223 (N_2223,N_2109,N_2174);
nand U2224 (N_2224,N_2154,N_2143);
xnor U2225 (N_2225,N_2152,N_2146);
nor U2226 (N_2226,N_2116,N_2118);
or U2227 (N_2227,N_2153,N_2167);
or U2228 (N_2228,N_2172,N_2112);
xnor U2229 (N_2229,N_2100,N_2130);
nor U2230 (N_2230,N_2123,N_2168);
and U2231 (N_2231,N_2144,N_2104);
and U2232 (N_2232,N_2104,N_2161);
and U2233 (N_2233,N_2169,N_2174);
or U2234 (N_2234,N_2100,N_2136);
nand U2235 (N_2235,N_2165,N_2126);
nor U2236 (N_2236,N_2144,N_2113);
xnor U2237 (N_2237,N_2139,N_2167);
xnor U2238 (N_2238,N_2107,N_2165);
nand U2239 (N_2239,N_2120,N_2167);
nor U2240 (N_2240,N_2168,N_2151);
xnor U2241 (N_2241,N_2119,N_2107);
xor U2242 (N_2242,N_2125,N_2141);
nor U2243 (N_2243,N_2140,N_2145);
and U2244 (N_2244,N_2135,N_2129);
or U2245 (N_2245,N_2167,N_2129);
nand U2246 (N_2246,N_2124,N_2115);
nand U2247 (N_2247,N_2113,N_2104);
and U2248 (N_2248,N_2145,N_2131);
and U2249 (N_2249,N_2114,N_2131);
xnor U2250 (N_2250,N_2198,N_2176);
or U2251 (N_2251,N_2242,N_2235);
nor U2252 (N_2252,N_2229,N_2228);
or U2253 (N_2253,N_2211,N_2175);
and U2254 (N_2254,N_2191,N_2180);
xor U2255 (N_2255,N_2244,N_2192);
and U2256 (N_2256,N_2220,N_2215);
or U2257 (N_2257,N_2208,N_2184);
or U2258 (N_2258,N_2224,N_2197);
or U2259 (N_2259,N_2183,N_2195);
and U2260 (N_2260,N_2194,N_2189);
and U2261 (N_2261,N_2210,N_2193);
and U2262 (N_2262,N_2234,N_2202);
and U2263 (N_2263,N_2206,N_2177);
or U2264 (N_2264,N_2217,N_2231);
or U2265 (N_2265,N_2247,N_2240);
xnor U2266 (N_2266,N_2221,N_2209);
and U2267 (N_2267,N_2222,N_2214);
and U2268 (N_2268,N_2218,N_2225);
nor U2269 (N_2269,N_2245,N_2186);
or U2270 (N_2270,N_2216,N_2188);
or U2271 (N_2271,N_2236,N_2237);
nor U2272 (N_2272,N_2219,N_2199);
nand U2273 (N_2273,N_2185,N_2181);
and U2274 (N_2274,N_2212,N_2233);
and U2275 (N_2275,N_2227,N_2204);
or U2276 (N_2276,N_2190,N_2239);
or U2277 (N_2277,N_2201,N_2223);
nand U2278 (N_2278,N_2178,N_2243);
nand U2279 (N_2279,N_2205,N_2248);
or U2280 (N_2280,N_2249,N_2196);
xor U2281 (N_2281,N_2232,N_2182);
nor U2282 (N_2282,N_2246,N_2230);
or U2283 (N_2283,N_2213,N_2203);
xnor U2284 (N_2284,N_2207,N_2238);
nand U2285 (N_2285,N_2179,N_2187);
and U2286 (N_2286,N_2226,N_2241);
and U2287 (N_2287,N_2200,N_2208);
xnor U2288 (N_2288,N_2233,N_2206);
nand U2289 (N_2289,N_2203,N_2190);
or U2290 (N_2290,N_2198,N_2234);
nand U2291 (N_2291,N_2226,N_2207);
xor U2292 (N_2292,N_2227,N_2224);
and U2293 (N_2293,N_2237,N_2190);
xnor U2294 (N_2294,N_2211,N_2237);
xor U2295 (N_2295,N_2206,N_2244);
nand U2296 (N_2296,N_2248,N_2211);
or U2297 (N_2297,N_2223,N_2186);
and U2298 (N_2298,N_2194,N_2242);
or U2299 (N_2299,N_2210,N_2201);
nand U2300 (N_2300,N_2237,N_2198);
nor U2301 (N_2301,N_2229,N_2244);
nand U2302 (N_2302,N_2186,N_2208);
or U2303 (N_2303,N_2242,N_2179);
and U2304 (N_2304,N_2189,N_2213);
xor U2305 (N_2305,N_2247,N_2234);
nor U2306 (N_2306,N_2177,N_2207);
xor U2307 (N_2307,N_2181,N_2200);
nor U2308 (N_2308,N_2246,N_2200);
nor U2309 (N_2309,N_2229,N_2191);
or U2310 (N_2310,N_2219,N_2213);
nor U2311 (N_2311,N_2231,N_2210);
nand U2312 (N_2312,N_2217,N_2235);
xnor U2313 (N_2313,N_2183,N_2249);
xor U2314 (N_2314,N_2225,N_2248);
nor U2315 (N_2315,N_2198,N_2175);
xor U2316 (N_2316,N_2185,N_2216);
or U2317 (N_2317,N_2203,N_2223);
or U2318 (N_2318,N_2200,N_2239);
nor U2319 (N_2319,N_2248,N_2235);
nand U2320 (N_2320,N_2199,N_2216);
and U2321 (N_2321,N_2211,N_2224);
or U2322 (N_2322,N_2202,N_2224);
nor U2323 (N_2323,N_2248,N_2247);
or U2324 (N_2324,N_2205,N_2192);
nand U2325 (N_2325,N_2277,N_2323);
and U2326 (N_2326,N_2265,N_2282);
and U2327 (N_2327,N_2305,N_2251);
xnor U2328 (N_2328,N_2272,N_2319);
xnor U2329 (N_2329,N_2256,N_2263);
nor U2330 (N_2330,N_2276,N_2281);
nand U2331 (N_2331,N_2304,N_2288);
and U2332 (N_2332,N_2306,N_2274);
xnor U2333 (N_2333,N_2311,N_2250);
nand U2334 (N_2334,N_2270,N_2314);
nand U2335 (N_2335,N_2308,N_2280);
nor U2336 (N_2336,N_2262,N_2255);
xnor U2337 (N_2337,N_2278,N_2275);
nor U2338 (N_2338,N_2303,N_2254);
nor U2339 (N_2339,N_2318,N_2283);
or U2340 (N_2340,N_2320,N_2293);
nand U2341 (N_2341,N_2309,N_2313);
and U2342 (N_2342,N_2266,N_2315);
xor U2343 (N_2343,N_2324,N_2259);
or U2344 (N_2344,N_2294,N_2261);
and U2345 (N_2345,N_2287,N_2296);
or U2346 (N_2346,N_2300,N_2269);
and U2347 (N_2347,N_2301,N_2273);
xnor U2348 (N_2348,N_2286,N_2297);
nor U2349 (N_2349,N_2284,N_2267);
or U2350 (N_2350,N_2291,N_2317);
xor U2351 (N_2351,N_2292,N_2298);
xnor U2352 (N_2352,N_2316,N_2264);
xnor U2353 (N_2353,N_2295,N_2321);
and U2354 (N_2354,N_2307,N_2322);
nand U2355 (N_2355,N_2268,N_2279);
or U2356 (N_2356,N_2312,N_2285);
xnor U2357 (N_2357,N_2260,N_2258);
or U2358 (N_2358,N_2252,N_2290);
nor U2359 (N_2359,N_2289,N_2302);
xor U2360 (N_2360,N_2310,N_2253);
and U2361 (N_2361,N_2299,N_2271);
or U2362 (N_2362,N_2257,N_2306);
and U2363 (N_2363,N_2319,N_2315);
xor U2364 (N_2364,N_2254,N_2296);
xnor U2365 (N_2365,N_2293,N_2297);
and U2366 (N_2366,N_2322,N_2287);
and U2367 (N_2367,N_2255,N_2250);
and U2368 (N_2368,N_2254,N_2253);
xor U2369 (N_2369,N_2318,N_2268);
nand U2370 (N_2370,N_2324,N_2261);
and U2371 (N_2371,N_2262,N_2287);
or U2372 (N_2372,N_2276,N_2278);
or U2373 (N_2373,N_2320,N_2324);
nor U2374 (N_2374,N_2304,N_2298);
and U2375 (N_2375,N_2303,N_2301);
and U2376 (N_2376,N_2309,N_2304);
and U2377 (N_2377,N_2272,N_2258);
nor U2378 (N_2378,N_2261,N_2283);
nand U2379 (N_2379,N_2270,N_2256);
or U2380 (N_2380,N_2251,N_2259);
and U2381 (N_2381,N_2289,N_2262);
nand U2382 (N_2382,N_2267,N_2274);
nor U2383 (N_2383,N_2288,N_2270);
or U2384 (N_2384,N_2296,N_2276);
and U2385 (N_2385,N_2277,N_2320);
nor U2386 (N_2386,N_2309,N_2318);
or U2387 (N_2387,N_2272,N_2277);
nand U2388 (N_2388,N_2260,N_2259);
nor U2389 (N_2389,N_2284,N_2323);
nor U2390 (N_2390,N_2313,N_2276);
xnor U2391 (N_2391,N_2270,N_2274);
xor U2392 (N_2392,N_2261,N_2251);
xnor U2393 (N_2393,N_2263,N_2253);
and U2394 (N_2394,N_2278,N_2251);
and U2395 (N_2395,N_2284,N_2250);
nor U2396 (N_2396,N_2277,N_2306);
nor U2397 (N_2397,N_2314,N_2324);
xnor U2398 (N_2398,N_2252,N_2318);
and U2399 (N_2399,N_2267,N_2282);
xor U2400 (N_2400,N_2361,N_2399);
xnor U2401 (N_2401,N_2339,N_2356);
and U2402 (N_2402,N_2384,N_2380);
and U2403 (N_2403,N_2372,N_2341);
nand U2404 (N_2404,N_2369,N_2336);
xor U2405 (N_2405,N_2383,N_2386);
nor U2406 (N_2406,N_2374,N_2355);
and U2407 (N_2407,N_2343,N_2357);
or U2408 (N_2408,N_2368,N_2391);
and U2409 (N_2409,N_2332,N_2342);
or U2410 (N_2410,N_2364,N_2360);
and U2411 (N_2411,N_2388,N_2325);
and U2412 (N_2412,N_2340,N_2334);
and U2413 (N_2413,N_2366,N_2337);
xor U2414 (N_2414,N_2377,N_2394);
xor U2415 (N_2415,N_2375,N_2351);
and U2416 (N_2416,N_2335,N_2345);
xnor U2417 (N_2417,N_2327,N_2363);
and U2418 (N_2418,N_2385,N_2367);
nor U2419 (N_2419,N_2371,N_2397);
nand U2420 (N_2420,N_2338,N_2330);
xor U2421 (N_2421,N_2354,N_2379);
and U2422 (N_2422,N_2396,N_2331);
nor U2423 (N_2423,N_2349,N_2359);
nor U2424 (N_2424,N_2346,N_2350);
nand U2425 (N_2425,N_2387,N_2390);
nand U2426 (N_2426,N_2395,N_2382);
nand U2427 (N_2427,N_2376,N_2329);
xor U2428 (N_2428,N_2358,N_2328);
xnor U2429 (N_2429,N_2378,N_2373);
or U2430 (N_2430,N_2389,N_2347);
nor U2431 (N_2431,N_2392,N_2393);
nor U2432 (N_2432,N_2365,N_2326);
nand U2433 (N_2433,N_2353,N_2398);
xor U2434 (N_2434,N_2348,N_2352);
nor U2435 (N_2435,N_2362,N_2381);
and U2436 (N_2436,N_2333,N_2344);
nor U2437 (N_2437,N_2370,N_2381);
nor U2438 (N_2438,N_2350,N_2369);
nand U2439 (N_2439,N_2348,N_2380);
nor U2440 (N_2440,N_2377,N_2381);
nand U2441 (N_2441,N_2325,N_2362);
xor U2442 (N_2442,N_2325,N_2387);
xnor U2443 (N_2443,N_2353,N_2385);
nor U2444 (N_2444,N_2393,N_2362);
nand U2445 (N_2445,N_2377,N_2396);
xnor U2446 (N_2446,N_2369,N_2334);
xnor U2447 (N_2447,N_2340,N_2387);
xnor U2448 (N_2448,N_2392,N_2361);
nor U2449 (N_2449,N_2399,N_2398);
and U2450 (N_2450,N_2371,N_2377);
xnor U2451 (N_2451,N_2341,N_2378);
xor U2452 (N_2452,N_2346,N_2335);
and U2453 (N_2453,N_2378,N_2343);
nor U2454 (N_2454,N_2398,N_2364);
xnor U2455 (N_2455,N_2347,N_2386);
xor U2456 (N_2456,N_2364,N_2388);
or U2457 (N_2457,N_2375,N_2382);
or U2458 (N_2458,N_2353,N_2335);
nor U2459 (N_2459,N_2336,N_2349);
xor U2460 (N_2460,N_2337,N_2342);
nand U2461 (N_2461,N_2378,N_2384);
and U2462 (N_2462,N_2383,N_2326);
xor U2463 (N_2463,N_2343,N_2386);
nor U2464 (N_2464,N_2348,N_2328);
and U2465 (N_2465,N_2326,N_2362);
or U2466 (N_2466,N_2373,N_2375);
or U2467 (N_2467,N_2380,N_2340);
xor U2468 (N_2468,N_2357,N_2390);
xnor U2469 (N_2469,N_2360,N_2336);
nor U2470 (N_2470,N_2371,N_2360);
nor U2471 (N_2471,N_2392,N_2375);
xnor U2472 (N_2472,N_2385,N_2329);
or U2473 (N_2473,N_2334,N_2341);
nand U2474 (N_2474,N_2358,N_2356);
nand U2475 (N_2475,N_2426,N_2403);
or U2476 (N_2476,N_2417,N_2446);
nor U2477 (N_2477,N_2408,N_2457);
xor U2478 (N_2478,N_2405,N_2414);
xnor U2479 (N_2479,N_2466,N_2418);
nor U2480 (N_2480,N_2436,N_2404);
xor U2481 (N_2481,N_2434,N_2439);
or U2482 (N_2482,N_2419,N_2409);
nand U2483 (N_2483,N_2410,N_2471);
nor U2484 (N_2484,N_2430,N_2453);
xnor U2485 (N_2485,N_2463,N_2460);
and U2486 (N_2486,N_2447,N_2444);
nand U2487 (N_2487,N_2445,N_2448);
nor U2488 (N_2488,N_2469,N_2454);
nor U2489 (N_2489,N_2415,N_2442);
nor U2490 (N_2490,N_2411,N_2416);
xnor U2491 (N_2491,N_2423,N_2452);
xor U2492 (N_2492,N_2425,N_2441);
or U2493 (N_2493,N_2449,N_2431);
or U2494 (N_2494,N_2473,N_2458);
or U2495 (N_2495,N_2421,N_2461);
and U2496 (N_2496,N_2401,N_2438);
or U2497 (N_2497,N_2462,N_2400);
or U2498 (N_2498,N_2427,N_2459);
or U2499 (N_2499,N_2474,N_2432);
and U2500 (N_2500,N_2451,N_2422);
and U2501 (N_2501,N_2440,N_2406);
and U2502 (N_2502,N_2467,N_2464);
xor U2503 (N_2503,N_2424,N_2413);
or U2504 (N_2504,N_2472,N_2429);
nand U2505 (N_2505,N_2437,N_2470);
nor U2506 (N_2506,N_2402,N_2468);
and U2507 (N_2507,N_2465,N_2412);
nor U2508 (N_2508,N_2456,N_2433);
xnor U2509 (N_2509,N_2435,N_2443);
and U2510 (N_2510,N_2428,N_2420);
nor U2511 (N_2511,N_2407,N_2455);
nor U2512 (N_2512,N_2450,N_2430);
and U2513 (N_2513,N_2436,N_2412);
or U2514 (N_2514,N_2441,N_2433);
and U2515 (N_2515,N_2444,N_2448);
or U2516 (N_2516,N_2448,N_2433);
nor U2517 (N_2517,N_2443,N_2455);
or U2518 (N_2518,N_2428,N_2404);
nand U2519 (N_2519,N_2457,N_2429);
xnor U2520 (N_2520,N_2421,N_2457);
xor U2521 (N_2521,N_2455,N_2400);
or U2522 (N_2522,N_2419,N_2453);
nand U2523 (N_2523,N_2417,N_2414);
nor U2524 (N_2524,N_2474,N_2422);
nand U2525 (N_2525,N_2406,N_2441);
nor U2526 (N_2526,N_2403,N_2413);
nand U2527 (N_2527,N_2453,N_2470);
and U2528 (N_2528,N_2424,N_2460);
nor U2529 (N_2529,N_2422,N_2408);
nand U2530 (N_2530,N_2459,N_2405);
nor U2531 (N_2531,N_2460,N_2435);
xnor U2532 (N_2532,N_2421,N_2462);
nand U2533 (N_2533,N_2454,N_2409);
xor U2534 (N_2534,N_2457,N_2414);
or U2535 (N_2535,N_2435,N_2402);
or U2536 (N_2536,N_2427,N_2455);
and U2537 (N_2537,N_2417,N_2444);
nand U2538 (N_2538,N_2426,N_2422);
nor U2539 (N_2539,N_2457,N_2470);
or U2540 (N_2540,N_2457,N_2443);
nor U2541 (N_2541,N_2434,N_2404);
xnor U2542 (N_2542,N_2463,N_2401);
or U2543 (N_2543,N_2401,N_2430);
nor U2544 (N_2544,N_2430,N_2447);
or U2545 (N_2545,N_2442,N_2473);
xor U2546 (N_2546,N_2453,N_2425);
and U2547 (N_2547,N_2452,N_2451);
or U2548 (N_2548,N_2453,N_2456);
xnor U2549 (N_2549,N_2453,N_2422);
nor U2550 (N_2550,N_2484,N_2513);
xor U2551 (N_2551,N_2542,N_2535);
nand U2552 (N_2552,N_2525,N_2492);
xor U2553 (N_2553,N_2500,N_2501);
or U2554 (N_2554,N_2526,N_2502);
and U2555 (N_2555,N_2538,N_2507);
nor U2556 (N_2556,N_2485,N_2512);
and U2557 (N_2557,N_2546,N_2519);
nand U2558 (N_2558,N_2530,N_2534);
nand U2559 (N_2559,N_2533,N_2498);
nand U2560 (N_2560,N_2489,N_2523);
nand U2561 (N_2561,N_2475,N_2478);
and U2562 (N_2562,N_2529,N_2532);
nand U2563 (N_2563,N_2515,N_2518);
or U2564 (N_2564,N_2544,N_2545);
nor U2565 (N_2565,N_2483,N_2539);
xor U2566 (N_2566,N_2482,N_2487);
xor U2567 (N_2567,N_2508,N_2511);
xor U2568 (N_2568,N_2514,N_2520);
xor U2569 (N_2569,N_2496,N_2476);
and U2570 (N_2570,N_2488,N_2506);
and U2571 (N_2571,N_2497,N_2527);
and U2572 (N_2572,N_2549,N_2509);
and U2573 (N_2573,N_2541,N_2522);
xor U2574 (N_2574,N_2493,N_2491);
and U2575 (N_2575,N_2504,N_2543);
nor U2576 (N_2576,N_2537,N_2505);
nor U2577 (N_2577,N_2524,N_2536);
nor U2578 (N_2578,N_2517,N_2547);
xor U2579 (N_2579,N_2477,N_2516);
xnor U2580 (N_2580,N_2503,N_2494);
and U2581 (N_2581,N_2521,N_2540);
and U2582 (N_2582,N_2499,N_2479);
and U2583 (N_2583,N_2486,N_2510);
nor U2584 (N_2584,N_2480,N_2548);
nand U2585 (N_2585,N_2531,N_2481);
nand U2586 (N_2586,N_2490,N_2528);
and U2587 (N_2587,N_2495,N_2520);
nor U2588 (N_2588,N_2532,N_2478);
nand U2589 (N_2589,N_2509,N_2501);
nand U2590 (N_2590,N_2539,N_2535);
nor U2591 (N_2591,N_2542,N_2512);
and U2592 (N_2592,N_2499,N_2488);
and U2593 (N_2593,N_2496,N_2532);
nand U2594 (N_2594,N_2487,N_2479);
nand U2595 (N_2595,N_2502,N_2547);
and U2596 (N_2596,N_2522,N_2489);
nand U2597 (N_2597,N_2505,N_2535);
or U2598 (N_2598,N_2476,N_2542);
nor U2599 (N_2599,N_2534,N_2482);
and U2600 (N_2600,N_2532,N_2494);
nand U2601 (N_2601,N_2522,N_2526);
nand U2602 (N_2602,N_2538,N_2534);
xnor U2603 (N_2603,N_2477,N_2476);
xnor U2604 (N_2604,N_2515,N_2536);
nor U2605 (N_2605,N_2501,N_2525);
nor U2606 (N_2606,N_2538,N_2531);
nand U2607 (N_2607,N_2517,N_2487);
or U2608 (N_2608,N_2508,N_2493);
nor U2609 (N_2609,N_2502,N_2498);
nor U2610 (N_2610,N_2547,N_2516);
xor U2611 (N_2611,N_2519,N_2507);
and U2612 (N_2612,N_2488,N_2485);
nor U2613 (N_2613,N_2515,N_2488);
xor U2614 (N_2614,N_2481,N_2499);
nand U2615 (N_2615,N_2539,N_2498);
or U2616 (N_2616,N_2493,N_2548);
or U2617 (N_2617,N_2528,N_2480);
xor U2618 (N_2618,N_2502,N_2493);
nand U2619 (N_2619,N_2476,N_2523);
or U2620 (N_2620,N_2547,N_2514);
nor U2621 (N_2621,N_2493,N_2513);
nand U2622 (N_2622,N_2476,N_2492);
xor U2623 (N_2623,N_2534,N_2549);
xnor U2624 (N_2624,N_2509,N_2476);
nor U2625 (N_2625,N_2602,N_2590);
and U2626 (N_2626,N_2584,N_2554);
nand U2627 (N_2627,N_2593,N_2579);
or U2628 (N_2628,N_2561,N_2607);
nand U2629 (N_2629,N_2591,N_2614);
and U2630 (N_2630,N_2565,N_2577);
and U2631 (N_2631,N_2612,N_2570);
or U2632 (N_2632,N_2575,N_2599);
xor U2633 (N_2633,N_2601,N_2571);
nor U2634 (N_2634,N_2566,N_2553);
and U2635 (N_2635,N_2598,N_2617);
nand U2636 (N_2636,N_2564,N_2592);
or U2637 (N_2637,N_2594,N_2606);
nand U2638 (N_2638,N_2624,N_2619);
xor U2639 (N_2639,N_2573,N_2557);
nand U2640 (N_2640,N_2572,N_2595);
and U2641 (N_2641,N_2611,N_2618);
xnor U2642 (N_2642,N_2567,N_2589);
and U2643 (N_2643,N_2622,N_2581);
and U2644 (N_2644,N_2613,N_2615);
xor U2645 (N_2645,N_2620,N_2609);
and U2646 (N_2646,N_2562,N_2596);
xnor U2647 (N_2647,N_2556,N_2621);
and U2648 (N_2648,N_2608,N_2574);
xor U2649 (N_2649,N_2587,N_2580);
xnor U2650 (N_2650,N_2568,N_2623);
nand U2651 (N_2651,N_2569,N_2578);
or U2652 (N_2652,N_2576,N_2610);
xnor U2653 (N_2653,N_2597,N_2552);
nor U2654 (N_2654,N_2551,N_2550);
xor U2655 (N_2655,N_2600,N_2583);
xor U2656 (N_2656,N_2563,N_2585);
xor U2657 (N_2657,N_2555,N_2560);
or U2658 (N_2658,N_2586,N_2559);
nor U2659 (N_2659,N_2582,N_2603);
xnor U2660 (N_2660,N_2558,N_2604);
xor U2661 (N_2661,N_2605,N_2616);
and U2662 (N_2662,N_2588,N_2603);
and U2663 (N_2663,N_2597,N_2624);
xor U2664 (N_2664,N_2561,N_2609);
nor U2665 (N_2665,N_2566,N_2578);
or U2666 (N_2666,N_2565,N_2581);
and U2667 (N_2667,N_2620,N_2553);
xnor U2668 (N_2668,N_2619,N_2553);
nor U2669 (N_2669,N_2618,N_2612);
nor U2670 (N_2670,N_2564,N_2610);
nand U2671 (N_2671,N_2590,N_2606);
nand U2672 (N_2672,N_2552,N_2610);
or U2673 (N_2673,N_2608,N_2561);
xnor U2674 (N_2674,N_2573,N_2554);
and U2675 (N_2675,N_2568,N_2603);
and U2676 (N_2676,N_2551,N_2607);
and U2677 (N_2677,N_2583,N_2595);
or U2678 (N_2678,N_2614,N_2581);
nand U2679 (N_2679,N_2600,N_2560);
xnor U2680 (N_2680,N_2620,N_2581);
nand U2681 (N_2681,N_2597,N_2615);
xor U2682 (N_2682,N_2551,N_2558);
or U2683 (N_2683,N_2606,N_2586);
nand U2684 (N_2684,N_2599,N_2566);
or U2685 (N_2685,N_2604,N_2582);
nand U2686 (N_2686,N_2611,N_2562);
nand U2687 (N_2687,N_2604,N_2598);
nand U2688 (N_2688,N_2580,N_2553);
nor U2689 (N_2689,N_2554,N_2590);
nand U2690 (N_2690,N_2620,N_2590);
nand U2691 (N_2691,N_2563,N_2564);
and U2692 (N_2692,N_2595,N_2581);
or U2693 (N_2693,N_2558,N_2573);
or U2694 (N_2694,N_2595,N_2565);
nor U2695 (N_2695,N_2550,N_2554);
and U2696 (N_2696,N_2568,N_2590);
xor U2697 (N_2697,N_2561,N_2558);
nand U2698 (N_2698,N_2572,N_2603);
xnor U2699 (N_2699,N_2600,N_2562);
nand U2700 (N_2700,N_2678,N_2671);
and U2701 (N_2701,N_2687,N_2664);
nor U2702 (N_2702,N_2690,N_2652);
xor U2703 (N_2703,N_2627,N_2666);
nand U2704 (N_2704,N_2686,N_2634);
or U2705 (N_2705,N_2679,N_2635);
nand U2706 (N_2706,N_2684,N_2693);
nor U2707 (N_2707,N_2654,N_2682);
nor U2708 (N_2708,N_2669,N_2660);
and U2709 (N_2709,N_2656,N_2647);
nand U2710 (N_2710,N_2643,N_2645);
xor U2711 (N_2711,N_2629,N_2696);
or U2712 (N_2712,N_2641,N_2685);
nor U2713 (N_2713,N_2638,N_2665);
xnor U2714 (N_2714,N_2688,N_2655);
or U2715 (N_2715,N_2681,N_2637);
nor U2716 (N_2716,N_2698,N_2630);
and U2717 (N_2717,N_2661,N_2657);
xnor U2718 (N_2718,N_2674,N_2680);
nand U2719 (N_2719,N_2646,N_2694);
and U2720 (N_2720,N_2689,N_2672);
nor U2721 (N_2721,N_2642,N_2668);
xor U2722 (N_2722,N_2628,N_2670);
and U2723 (N_2723,N_2636,N_2691);
or U2724 (N_2724,N_2699,N_2625);
or U2725 (N_2725,N_2662,N_2640);
nor U2726 (N_2726,N_2639,N_2651);
or U2727 (N_2727,N_2697,N_2677);
or U2728 (N_2728,N_2683,N_2695);
or U2729 (N_2729,N_2658,N_2663);
or U2730 (N_2730,N_2659,N_2650);
nor U2731 (N_2731,N_2648,N_2626);
nor U2732 (N_2732,N_2644,N_2649);
nand U2733 (N_2733,N_2676,N_2667);
xnor U2734 (N_2734,N_2692,N_2631);
xnor U2735 (N_2735,N_2673,N_2653);
or U2736 (N_2736,N_2675,N_2632);
and U2737 (N_2737,N_2633,N_2656);
xnor U2738 (N_2738,N_2670,N_2633);
xnor U2739 (N_2739,N_2636,N_2676);
and U2740 (N_2740,N_2662,N_2626);
and U2741 (N_2741,N_2679,N_2645);
or U2742 (N_2742,N_2687,N_2689);
or U2743 (N_2743,N_2686,N_2644);
and U2744 (N_2744,N_2672,N_2651);
nand U2745 (N_2745,N_2627,N_2635);
nor U2746 (N_2746,N_2692,N_2649);
nand U2747 (N_2747,N_2634,N_2698);
nand U2748 (N_2748,N_2636,N_2660);
xor U2749 (N_2749,N_2665,N_2691);
and U2750 (N_2750,N_2635,N_2677);
or U2751 (N_2751,N_2648,N_2699);
nand U2752 (N_2752,N_2676,N_2671);
or U2753 (N_2753,N_2669,N_2688);
nand U2754 (N_2754,N_2682,N_2690);
nand U2755 (N_2755,N_2628,N_2652);
nand U2756 (N_2756,N_2680,N_2662);
nor U2757 (N_2757,N_2626,N_2646);
and U2758 (N_2758,N_2641,N_2687);
xnor U2759 (N_2759,N_2642,N_2635);
or U2760 (N_2760,N_2675,N_2682);
nand U2761 (N_2761,N_2646,N_2683);
or U2762 (N_2762,N_2625,N_2665);
nand U2763 (N_2763,N_2633,N_2657);
nand U2764 (N_2764,N_2648,N_2656);
xor U2765 (N_2765,N_2675,N_2679);
nor U2766 (N_2766,N_2683,N_2656);
nor U2767 (N_2767,N_2632,N_2649);
xor U2768 (N_2768,N_2682,N_2672);
nand U2769 (N_2769,N_2643,N_2674);
or U2770 (N_2770,N_2626,N_2697);
or U2771 (N_2771,N_2664,N_2632);
xor U2772 (N_2772,N_2695,N_2650);
nand U2773 (N_2773,N_2642,N_2685);
nor U2774 (N_2774,N_2644,N_2625);
or U2775 (N_2775,N_2723,N_2724);
or U2776 (N_2776,N_2774,N_2749);
nor U2777 (N_2777,N_2713,N_2735);
or U2778 (N_2778,N_2740,N_2771);
or U2779 (N_2779,N_2703,N_2748);
nor U2780 (N_2780,N_2764,N_2729);
nor U2781 (N_2781,N_2734,N_2730);
nand U2782 (N_2782,N_2707,N_2712);
xor U2783 (N_2783,N_2769,N_2747);
nand U2784 (N_2784,N_2733,N_2717);
xnor U2785 (N_2785,N_2755,N_2756);
xnor U2786 (N_2786,N_2753,N_2727);
or U2787 (N_2787,N_2742,N_2705);
and U2788 (N_2788,N_2757,N_2759);
or U2789 (N_2789,N_2765,N_2767);
nor U2790 (N_2790,N_2728,N_2743);
nand U2791 (N_2791,N_2710,N_2726);
or U2792 (N_2792,N_2773,N_2709);
or U2793 (N_2793,N_2702,N_2718);
xor U2794 (N_2794,N_2744,N_2715);
and U2795 (N_2795,N_2762,N_2766);
nand U2796 (N_2796,N_2751,N_2770);
or U2797 (N_2797,N_2741,N_2736);
or U2798 (N_2798,N_2758,N_2760);
xor U2799 (N_2799,N_2711,N_2763);
nor U2800 (N_2800,N_2739,N_2701);
nand U2801 (N_2801,N_2732,N_2704);
xor U2802 (N_2802,N_2714,N_2722);
and U2803 (N_2803,N_2768,N_2725);
xnor U2804 (N_2804,N_2752,N_2738);
nor U2805 (N_2805,N_2716,N_2720);
xnor U2806 (N_2806,N_2754,N_2745);
xor U2807 (N_2807,N_2737,N_2706);
or U2808 (N_2808,N_2708,N_2731);
nor U2809 (N_2809,N_2772,N_2721);
and U2810 (N_2810,N_2700,N_2761);
nand U2811 (N_2811,N_2750,N_2746);
or U2812 (N_2812,N_2719,N_2770);
nand U2813 (N_2813,N_2770,N_2760);
nor U2814 (N_2814,N_2749,N_2770);
xnor U2815 (N_2815,N_2728,N_2702);
nand U2816 (N_2816,N_2748,N_2767);
nand U2817 (N_2817,N_2756,N_2729);
nor U2818 (N_2818,N_2719,N_2722);
xnor U2819 (N_2819,N_2720,N_2711);
nor U2820 (N_2820,N_2758,N_2726);
and U2821 (N_2821,N_2717,N_2763);
and U2822 (N_2822,N_2769,N_2727);
xor U2823 (N_2823,N_2742,N_2761);
nand U2824 (N_2824,N_2710,N_2739);
nor U2825 (N_2825,N_2773,N_2744);
nor U2826 (N_2826,N_2711,N_2765);
and U2827 (N_2827,N_2719,N_2737);
nand U2828 (N_2828,N_2733,N_2704);
nor U2829 (N_2829,N_2720,N_2726);
or U2830 (N_2830,N_2764,N_2701);
nor U2831 (N_2831,N_2734,N_2714);
xor U2832 (N_2832,N_2747,N_2759);
xnor U2833 (N_2833,N_2740,N_2729);
or U2834 (N_2834,N_2758,N_2742);
nor U2835 (N_2835,N_2731,N_2707);
nor U2836 (N_2836,N_2716,N_2702);
nor U2837 (N_2837,N_2768,N_2757);
xnor U2838 (N_2838,N_2743,N_2709);
xor U2839 (N_2839,N_2755,N_2704);
nor U2840 (N_2840,N_2704,N_2701);
or U2841 (N_2841,N_2752,N_2705);
nand U2842 (N_2842,N_2718,N_2711);
or U2843 (N_2843,N_2769,N_2766);
or U2844 (N_2844,N_2708,N_2742);
and U2845 (N_2845,N_2731,N_2733);
and U2846 (N_2846,N_2724,N_2752);
nand U2847 (N_2847,N_2718,N_2707);
or U2848 (N_2848,N_2700,N_2719);
nand U2849 (N_2849,N_2734,N_2701);
or U2850 (N_2850,N_2834,N_2802);
nand U2851 (N_2851,N_2803,N_2826);
or U2852 (N_2852,N_2817,N_2848);
xor U2853 (N_2853,N_2830,N_2777);
and U2854 (N_2854,N_2820,N_2785);
xor U2855 (N_2855,N_2813,N_2791);
nand U2856 (N_2856,N_2779,N_2841);
xnor U2857 (N_2857,N_2784,N_2788);
nor U2858 (N_2858,N_2816,N_2805);
nor U2859 (N_2859,N_2845,N_2827);
nor U2860 (N_2860,N_2781,N_2804);
xnor U2861 (N_2861,N_2782,N_2849);
or U2862 (N_2862,N_2799,N_2831);
nand U2863 (N_2863,N_2847,N_2836);
or U2864 (N_2864,N_2833,N_2819);
nor U2865 (N_2865,N_2825,N_2795);
nand U2866 (N_2866,N_2811,N_2796);
nor U2867 (N_2867,N_2832,N_2829);
and U2868 (N_2868,N_2835,N_2823);
xor U2869 (N_2869,N_2807,N_2789);
and U2870 (N_2870,N_2775,N_2792);
xnor U2871 (N_2871,N_2839,N_2787);
or U2872 (N_2872,N_2776,N_2828);
nor U2873 (N_2873,N_2821,N_2786);
xnor U2874 (N_2874,N_2797,N_2800);
xor U2875 (N_2875,N_2794,N_2815);
nand U2876 (N_2876,N_2818,N_2808);
and U2877 (N_2877,N_2780,N_2809);
nor U2878 (N_2878,N_2838,N_2793);
and U2879 (N_2879,N_2824,N_2778);
nor U2880 (N_2880,N_2814,N_2842);
or U2881 (N_2881,N_2844,N_2806);
nand U2882 (N_2882,N_2822,N_2801);
or U2883 (N_2883,N_2812,N_2840);
or U2884 (N_2884,N_2783,N_2846);
or U2885 (N_2885,N_2798,N_2790);
nand U2886 (N_2886,N_2843,N_2810);
or U2887 (N_2887,N_2837,N_2810);
or U2888 (N_2888,N_2848,N_2778);
and U2889 (N_2889,N_2840,N_2799);
nor U2890 (N_2890,N_2837,N_2846);
and U2891 (N_2891,N_2787,N_2848);
nand U2892 (N_2892,N_2831,N_2782);
and U2893 (N_2893,N_2796,N_2806);
nor U2894 (N_2894,N_2796,N_2826);
or U2895 (N_2895,N_2830,N_2791);
or U2896 (N_2896,N_2829,N_2814);
or U2897 (N_2897,N_2785,N_2835);
and U2898 (N_2898,N_2844,N_2798);
and U2899 (N_2899,N_2778,N_2793);
nor U2900 (N_2900,N_2808,N_2792);
nor U2901 (N_2901,N_2792,N_2789);
nand U2902 (N_2902,N_2793,N_2797);
xnor U2903 (N_2903,N_2814,N_2823);
nor U2904 (N_2904,N_2775,N_2844);
or U2905 (N_2905,N_2792,N_2820);
xor U2906 (N_2906,N_2798,N_2822);
or U2907 (N_2907,N_2790,N_2779);
xor U2908 (N_2908,N_2821,N_2785);
or U2909 (N_2909,N_2794,N_2842);
nand U2910 (N_2910,N_2776,N_2805);
nor U2911 (N_2911,N_2837,N_2825);
or U2912 (N_2912,N_2779,N_2814);
or U2913 (N_2913,N_2793,N_2781);
nor U2914 (N_2914,N_2839,N_2826);
or U2915 (N_2915,N_2818,N_2829);
xnor U2916 (N_2916,N_2813,N_2778);
xnor U2917 (N_2917,N_2836,N_2844);
nand U2918 (N_2918,N_2837,N_2817);
and U2919 (N_2919,N_2818,N_2837);
and U2920 (N_2920,N_2784,N_2781);
nand U2921 (N_2921,N_2829,N_2801);
nand U2922 (N_2922,N_2788,N_2831);
xnor U2923 (N_2923,N_2846,N_2790);
and U2924 (N_2924,N_2832,N_2816);
and U2925 (N_2925,N_2891,N_2888);
or U2926 (N_2926,N_2902,N_2904);
or U2927 (N_2927,N_2897,N_2916);
and U2928 (N_2928,N_2911,N_2866);
or U2929 (N_2929,N_2869,N_2921);
nor U2930 (N_2930,N_2895,N_2913);
xnor U2931 (N_2931,N_2896,N_2868);
or U2932 (N_2932,N_2872,N_2882);
nand U2933 (N_2933,N_2892,N_2865);
xor U2934 (N_2934,N_2906,N_2910);
or U2935 (N_2935,N_2908,N_2917);
nor U2936 (N_2936,N_2899,N_2862);
nand U2937 (N_2937,N_2878,N_2890);
and U2938 (N_2938,N_2903,N_2900);
nor U2939 (N_2939,N_2885,N_2857);
or U2940 (N_2940,N_2883,N_2914);
nand U2941 (N_2941,N_2923,N_2856);
nand U2942 (N_2942,N_2877,N_2894);
or U2943 (N_2943,N_2898,N_2909);
nand U2944 (N_2944,N_2864,N_2867);
and U2945 (N_2945,N_2855,N_2915);
xnor U2946 (N_2946,N_2922,N_2873);
xor U2947 (N_2947,N_2874,N_2876);
xor U2948 (N_2948,N_2870,N_2880);
nand U2949 (N_2949,N_2881,N_2854);
nor U2950 (N_2950,N_2852,N_2920);
xnor U2951 (N_2951,N_2887,N_2850);
and U2952 (N_2952,N_2893,N_2879);
or U2953 (N_2953,N_2861,N_2858);
xnor U2954 (N_2954,N_2884,N_2875);
or U2955 (N_2955,N_2907,N_2912);
nor U2956 (N_2956,N_2919,N_2924);
or U2957 (N_2957,N_2851,N_2859);
and U2958 (N_2958,N_2863,N_2905);
xor U2959 (N_2959,N_2853,N_2901);
and U2960 (N_2960,N_2918,N_2871);
or U2961 (N_2961,N_2860,N_2886);
nor U2962 (N_2962,N_2889,N_2888);
or U2963 (N_2963,N_2867,N_2865);
nor U2964 (N_2964,N_2916,N_2857);
xor U2965 (N_2965,N_2862,N_2869);
and U2966 (N_2966,N_2913,N_2860);
and U2967 (N_2967,N_2879,N_2865);
xor U2968 (N_2968,N_2870,N_2923);
and U2969 (N_2969,N_2873,N_2897);
xnor U2970 (N_2970,N_2873,N_2858);
xnor U2971 (N_2971,N_2854,N_2924);
nand U2972 (N_2972,N_2896,N_2922);
and U2973 (N_2973,N_2856,N_2859);
and U2974 (N_2974,N_2901,N_2899);
xor U2975 (N_2975,N_2864,N_2890);
and U2976 (N_2976,N_2870,N_2855);
and U2977 (N_2977,N_2879,N_2858);
xor U2978 (N_2978,N_2880,N_2894);
xnor U2979 (N_2979,N_2898,N_2851);
nand U2980 (N_2980,N_2860,N_2882);
nor U2981 (N_2981,N_2907,N_2863);
nor U2982 (N_2982,N_2891,N_2892);
nand U2983 (N_2983,N_2914,N_2918);
nor U2984 (N_2984,N_2856,N_2885);
xor U2985 (N_2985,N_2860,N_2903);
nand U2986 (N_2986,N_2854,N_2908);
nor U2987 (N_2987,N_2892,N_2893);
xor U2988 (N_2988,N_2875,N_2899);
or U2989 (N_2989,N_2871,N_2916);
xor U2990 (N_2990,N_2892,N_2872);
nor U2991 (N_2991,N_2923,N_2917);
nand U2992 (N_2992,N_2891,N_2852);
xnor U2993 (N_2993,N_2868,N_2872);
xor U2994 (N_2994,N_2913,N_2852);
xor U2995 (N_2995,N_2891,N_2906);
nand U2996 (N_2996,N_2907,N_2895);
nor U2997 (N_2997,N_2924,N_2875);
or U2998 (N_2998,N_2895,N_2891);
or U2999 (N_2999,N_2910,N_2867);
xor UO_0 (O_0,N_2993,N_2949);
and UO_1 (O_1,N_2996,N_2999);
nor UO_2 (O_2,N_2995,N_2983);
nor UO_3 (O_3,N_2930,N_2987);
nor UO_4 (O_4,N_2951,N_2955);
and UO_5 (O_5,N_2947,N_2972);
or UO_6 (O_6,N_2977,N_2986);
and UO_7 (O_7,N_2957,N_2939);
and UO_8 (O_8,N_2981,N_2950);
and UO_9 (O_9,N_2967,N_2989);
or UO_10 (O_10,N_2997,N_2948);
and UO_11 (O_11,N_2984,N_2988);
or UO_12 (O_12,N_2991,N_2944);
xnor UO_13 (O_13,N_2942,N_2959);
xnor UO_14 (O_14,N_2956,N_2941);
xor UO_15 (O_15,N_2961,N_2998);
xor UO_16 (O_16,N_2954,N_2945);
nand UO_17 (O_17,N_2932,N_2968);
nand UO_18 (O_18,N_2934,N_2926);
or UO_19 (O_19,N_2976,N_2974);
nor UO_20 (O_20,N_2952,N_2969);
and UO_21 (O_21,N_2933,N_2940);
or UO_22 (O_22,N_2994,N_2931);
or UO_23 (O_23,N_2938,N_2965);
xor UO_24 (O_24,N_2978,N_2980);
xnor UO_25 (O_25,N_2937,N_2990);
or UO_26 (O_26,N_2946,N_2982);
xnor UO_27 (O_27,N_2929,N_2970);
nor UO_28 (O_28,N_2928,N_2962);
nor UO_29 (O_29,N_2964,N_2953);
xnor UO_30 (O_30,N_2979,N_2925);
and UO_31 (O_31,N_2943,N_2975);
nor UO_32 (O_32,N_2966,N_2960);
xor UO_33 (O_33,N_2963,N_2958);
xor UO_34 (O_34,N_2971,N_2973);
xor UO_35 (O_35,N_2935,N_2985);
nor UO_36 (O_36,N_2927,N_2936);
nand UO_37 (O_37,N_2992,N_2951);
nor UO_38 (O_38,N_2975,N_2933);
and UO_39 (O_39,N_2989,N_2963);
xnor UO_40 (O_40,N_2954,N_2949);
or UO_41 (O_41,N_2938,N_2950);
and UO_42 (O_42,N_2974,N_2925);
nor UO_43 (O_43,N_2998,N_2926);
and UO_44 (O_44,N_2984,N_2980);
or UO_45 (O_45,N_2997,N_2996);
and UO_46 (O_46,N_2969,N_2991);
nor UO_47 (O_47,N_2965,N_2950);
or UO_48 (O_48,N_2929,N_2972);
and UO_49 (O_49,N_2985,N_2956);
nor UO_50 (O_50,N_2965,N_2968);
nor UO_51 (O_51,N_2989,N_2973);
nand UO_52 (O_52,N_2993,N_2974);
and UO_53 (O_53,N_2976,N_2960);
xor UO_54 (O_54,N_2980,N_2949);
xnor UO_55 (O_55,N_2928,N_2955);
nor UO_56 (O_56,N_2940,N_2963);
xor UO_57 (O_57,N_2997,N_2942);
nor UO_58 (O_58,N_2944,N_2935);
xnor UO_59 (O_59,N_2960,N_2941);
xnor UO_60 (O_60,N_2970,N_2945);
and UO_61 (O_61,N_2937,N_2996);
and UO_62 (O_62,N_2996,N_2954);
xnor UO_63 (O_63,N_2935,N_2968);
nor UO_64 (O_64,N_2963,N_2927);
xor UO_65 (O_65,N_2952,N_2943);
nor UO_66 (O_66,N_2975,N_2927);
or UO_67 (O_67,N_2948,N_2967);
nor UO_68 (O_68,N_2958,N_2933);
nor UO_69 (O_69,N_2931,N_2967);
or UO_70 (O_70,N_2952,N_2973);
xnor UO_71 (O_71,N_2954,N_2966);
and UO_72 (O_72,N_2941,N_2972);
nor UO_73 (O_73,N_2955,N_2933);
nand UO_74 (O_74,N_2997,N_2975);
nor UO_75 (O_75,N_2929,N_2985);
and UO_76 (O_76,N_2927,N_2946);
xor UO_77 (O_77,N_2955,N_2976);
xnor UO_78 (O_78,N_2994,N_2933);
nor UO_79 (O_79,N_2973,N_2959);
nand UO_80 (O_80,N_2942,N_2961);
nor UO_81 (O_81,N_2946,N_2931);
nor UO_82 (O_82,N_2999,N_2981);
or UO_83 (O_83,N_2949,N_2934);
nor UO_84 (O_84,N_2963,N_2954);
and UO_85 (O_85,N_2951,N_2931);
xor UO_86 (O_86,N_2962,N_2983);
xnor UO_87 (O_87,N_2991,N_2951);
nor UO_88 (O_88,N_2935,N_2991);
nand UO_89 (O_89,N_2928,N_2975);
and UO_90 (O_90,N_2947,N_2998);
or UO_91 (O_91,N_2975,N_2991);
xor UO_92 (O_92,N_2960,N_2952);
nor UO_93 (O_93,N_2976,N_2983);
nor UO_94 (O_94,N_2931,N_2964);
nand UO_95 (O_95,N_2977,N_2955);
nand UO_96 (O_96,N_2926,N_2980);
nor UO_97 (O_97,N_2969,N_2978);
or UO_98 (O_98,N_2955,N_2995);
nand UO_99 (O_99,N_2968,N_2947);
or UO_100 (O_100,N_2978,N_2977);
nor UO_101 (O_101,N_2926,N_2990);
nor UO_102 (O_102,N_2983,N_2946);
xnor UO_103 (O_103,N_2996,N_2961);
nand UO_104 (O_104,N_2926,N_2939);
and UO_105 (O_105,N_2937,N_2960);
and UO_106 (O_106,N_2969,N_2976);
xor UO_107 (O_107,N_2957,N_2950);
nand UO_108 (O_108,N_2966,N_2971);
or UO_109 (O_109,N_2941,N_2955);
xnor UO_110 (O_110,N_2946,N_2935);
and UO_111 (O_111,N_2926,N_2947);
nor UO_112 (O_112,N_2928,N_2945);
nand UO_113 (O_113,N_2932,N_2982);
nor UO_114 (O_114,N_2981,N_2945);
nand UO_115 (O_115,N_2994,N_2953);
nor UO_116 (O_116,N_2946,N_2933);
nand UO_117 (O_117,N_2937,N_2992);
or UO_118 (O_118,N_2995,N_2969);
or UO_119 (O_119,N_2967,N_2993);
nand UO_120 (O_120,N_2953,N_2995);
xor UO_121 (O_121,N_2927,N_2954);
or UO_122 (O_122,N_2975,N_2952);
or UO_123 (O_123,N_2973,N_2934);
and UO_124 (O_124,N_2959,N_2930);
xnor UO_125 (O_125,N_2964,N_2935);
nor UO_126 (O_126,N_2956,N_2935);
xor UO_127 (O_127,N_2946,N_2988);
and UO_128 (O_128,N_2953,N_2925);
or UO_129 (O_129,N_2944,N_2938);
xor UO_130 (O_130,N_2991,N_2968);
nor UO_131 (O_131,N_2981,N_2951);
xnor UO_132 (O_132,N_2929,N_2971);
nor UO_133 (O_133,N_2961,N_2991);
xnor UO_134 (O_134,N_2998,N_2962);
xor UO_135 (O_135,N_2976,N_2997);
nand UO_136 (O_136,N_2957,N_2962);
xor UO_137 (O_137,N_2969,N_2928);
nand UO_138 (O_138,N_2986,N_2960);
nand UO_139 (O_139,N_2983,N_2966);
nor UO_140 (O_140,N_2953,N_2957);
nor UO_141 (O_141,N_2989,N_2969);
or UO_142 (O_142,N_2937,N_2987);
nand UO_143 (O_143,N_2958,N_2943);
or UO_144 (O_144,N_2937,N_2979);
or UO_145 (O_145,N_2961,N_2962);
xor UO_146 (O_146,N_2971,N_2964);
or UO_147 (O_147,N_2951,N_2932);
nor UO_148 (O_148,N_2967,N_2927);
xor UO_149 (O_149,N_2982,N_2958);
nand UO_150 (O_150,N_2939,N_2998);
or UO_151 (O_151,N_2944,N_2980);
nor UO_152 (O_152,N_2934,N_2935);
xnor UO_153 (O_153,N_2942,N_2957);
xor UO_154 (O_154,N_2962,N_2975);
and UO_155 (O_155,N_2927,N_2981);
and UO_156 (O_156,N_2964,N_2955);
nor UO_157 (O_157,N_2998,N_2970);
xor UO_158 (O_158,N_2944,N_2965);
or UO_159 (O_159,N_2994,N_2983);
and UO_160 (O_160,N_2926,N_2986);
xnor UO_161 (O_161,N_2961,N_2939);
nor UO_162 (O_162,N_2954,N_2998);
nand UO_163 (O_163,N_2981,N_2993);
or UO_164 (O_164,N_2973,N_2994);
xnor UO_165 (O_165,N_2933,N_2954);
or UO_166 (O_166,N_2999,N_2991);
or UO_167 (O_167,N_2940,N_2931);
or UO_168 (O_168,N_2935,N_2983);
nand UO_169 (O_169,N_2941,N_2967);
nor UO_170 (O_170,N_2952,N_2968);
nand UO_171 (O_171,N_2928,N_2947);
nor UO_172 (O_172,N_2980,N_2931);
nor UO_173 (O_173,N_2986,N_2945);
xnor UO_174 (O_174,N_2958,N_2956);
nand UO_175 (O_175,N_2997,N_2937);
nor UO_176 (O_176,N_2939,N_2992);
or UO_177 (O_177,N_2994,N_2929);
nand UO_178 (O_178,N_2995,N_2989);
xor UO_179 (O_179,N_2991,N_2946);
nor UO_180 (O_180,N_2996,N_2970);
or UO_181 (O_181,N_2967,N_2980);
xnor UO_182 (O_182,N_2996,N_2998);
xor UO_183 (O_183,N_2994,N_2980);
or UO_184 (O_184,N_2930,N_2969);
and UO_185 (O_185,N_2934,N_2930);
and UO_186 (O_186,N_2969,N_2984);
and UO_187 (O_187,N_2989,N_2966);
nor UO_188 (O_188,N_2935,N_2967);
nor UO_189 (O_189,N_2984,N_2994);
xnor UO_190 (O_190,N_2941,N_2954);
nor UO_191 (O_191,N_2978,N_2944);
and UO_192 (O_192,N_2938,N_2939);
and UO_193 (O_193,N_2957,N_2933);
xor UO_194 (O_194,N_2950,N_2932);
xnor UO_195 (O_195,N_2952,N_2996);
nor UO_196 (O_196,N_2927,N_2938);
nor UO_197 (O_197,N_2957,N_2973);
nor UO_198 (O_198,N_2991,N_2990);
xnor UO_199 (O_199,N_2939,N_2980);
nor UO_200 (O_200,N_2993,N_2979);
nand UO_201 (O_201,N_2967,N_2953);
and UO_202 (O_202,N_2964,N_2947);
nand UO_203 (O_203,N_2925,N_2956);
or UO_204 (O_204,N_2974,N_2990);
or UO_205 (O_205,N_2948,N_2977);
nand UO_206 (O_206,N_2965,N_2945);
nand UO_207 (O_207,N_2944,N_2951);
nand UO_208 (O_208,N_2934,N_2978);
or UO_209 (O_209,N_2971,N_2989);
xor UO_210 (O_210,N_2994,N_2982);
and UO_211 (O_211,N_2948,N_2970);
nor UO_212 (O_212,N_2969,N_2977);
xor UO_213 (O_213,N_2964,N_2967);
or UO_214 (O_214,N_2926,N_2984);
nand UO_215 (O_215,N_2932,N_2976);
nand UO_216 (O_216,N_2947,N_2967);
nor UO_217 (O_217,N_2951,N_2987);
or UO_218 (O_218,N_2961,N_2967);
xnor UO_219 (O_219,N_2958,N_2994);
and UO_220 (O_220,N_2932,N_2926);
and UO_221 (O_221,N_2929,N_2928);
nor UO_222 (O_222,N_2980,N_2986);
xnor UO_223 (O_223,N_2983,N_2939);
xnor UO_224 (O_224,N_2925,N_2982);
and UO_225 (O_225,N_2978,N_2998);
nand UO_226 (O_226,N_2966,N_2990);
nand UO_227 (O_227,N_2977,N_2974);
or UO_228 (O_228,N_2926,N_2979);
xnor UO_229 (O_229,N_2949,N_2995);
nor UO_230 (O_230,N_2986,N_2987);
or UO_231 (O_231,N_2932,N_2925);
nand UO_232 (O_232,N_2925,N_2993);
xor UO_233 (O_233,N_2999,N_2934);
nor UO_234 (O_234,N_2941,N_2949);
nor UO_235 (O_235,N_2966,N_2926);
or UO_236 (O_236,N_2929,N_2947);
or UO_237 (O_237,N_2982,N_2984);
nand UO_238 (O_238,N_2968,N_2974);
nand UO_239 (O_239,N_2966,N_2934);
nor UO_240 (O_240,N_2964,N_2941);
and UO_241 (O_241,N_2963,N_2961);
nor UO_242 (O_242,N_2930,N_2967);
or UO_243 (O_243,N_2954,N_2944);
nor UO_244 (O_244,N_2964,N_2929);
nand UO_245 (O_245,N_2974,N_2953);
nor UO_246 (O_246,N_2947,N_2984);
nand UO_247 (O_247,N_2957,N_2964);
and UO_248 (O_248,N_2986,N_2999);
nor UO_249 (O_249,N_2948,N_2966);
nand UO_250 (O_250,N_2943,N_2963);
or UO_251 (O_251,N_2990,N_2979);
nor UO_252 (O_252,N_2983,N_2998);
nand UO_253 (O_253,N_2979,N_2959);
xor UO_254 (O_254,N_2926,N_2965);
xor UO_255 (O_255,N_2961,N_2934);
nand UO_256 (O_256,N_2929,N_2942);
nand UO_257 (O_257,N_2936,N_2972);
and UO_258 (O_258,N_2965,N_2981);
and UO_259 (O_259,N_2947,N_2990);
or UO_260 (O_260,N_2990,N_2950);
or UO_261 (O_261,N_2988,N_2999);
nand UO_262 (O_262,N_2937,N_2972);
nand UO_263 (O_263,N_2951,N_2996);
nand UO_264 (O_264,N_2970,N_2935);
xor UO_265 (O_265,N_2957,N_2981);
and UO_266 (O_266,N_2926,N_2981);
nand UO_267 (O_267,N_2974,N_2975);
or UO_268 (O_268,N_2933,N_2948);
and UO_269 (O_269,N_2991,N_2978);
nor UO_270 (O_270,N_2931,N_2955);
or UO_271 (O_271,N_2942,N_2927);
or UO_272 (O_272,N_2956,N_2991);
or UO_273 (O_273,N_2928,N_2931);
or UO_274 (O_274,N_2967,N_2955);
nor UO_275 (O_275,N_2990,N_2980);
xnor UO_276 (O_276,N_2943,N_2927);
nand UO_277 (O_277,N_2959,N_2943);
or UO_278 (O_278,N_2936,N_2986);
xnor UO_279 (O_279,N_2932,N_2966);
or UO_280 (O_280,N_2996,N_2941);
and UO_281 (O_281,N_2999,N_2980);
nand UO_282 (O_282,N_2937,N_2925);
and UO_283 (O_283,N_2964,N_2961);
nand UO_284 (O_284,N_2965,N_2939);
xnor UO_285 (O_285,N_2930,N_2925);
nand UO_286 (O_286,N_2997,N_2986);
nor UO_287 (O_287,N_2978,N_2981);
nor UO_288 (O_288,N_2954,N_2942);
nand UO_289 (O_289,N_2954,N_2986);
and UO_290 (O_290,N_2983,N_2991);
nor UO_291 (O_291,N_2977,N_2991);
nand UO_292 (O_292,N_2936,N_2975);
nand UO_293 (O_293,N_2931,N_2959);
nor UO_294 (O_294,N_2928,N_2925);
or UO_295 (O_295,N_2958,N_2975);
nand UO_296 (O_296,N_2995,N_2960);
nor UO_297 (O_297,N_2936,N_2970);
nor UO_298 (O_298,N_2935,N_2971);
xor UO_299 (O_299,N_2987,N_2996);
nor UO_300 (O_300,N_2938,N_2966);
xnor UO_301 (O_301,N_2936,N_2931);
or UO_302 (O_302,N_2996,N_2977);
nor UO_303 (O_303,N_2928,N_2963);
xor UO_304 (O_304,N_2943,N_2999);
nor UO_305 (O_305,N_2937,N_2935);
nor UO_306 (O_306,N_2945,N_2938);
xor UO_307 (O_307,N_2963,N_2977);
or UO_308 (O_308,N_2950,N_2969);
xnor UO_309 (O_309,N_2950,N_2976);
xor UO_310 (O_310,N_2977,N_2992);
xor UO_311 (O_311,N_2976,N_2965);
xor UO_312 (O_312,N_2932,N_2996);
nand UO_313 (O_313,N_2935,N_2990);
xor UO_314 (O_314,N_2978,N_2972);
nand UO_315 (O_315,N_2940,N_2947);
and UO_316 (O_316,N_2951,N_2975);
nor UO_317 (O_317,N_2963,N_2999);
and UO_318 (O_318,N_2955,N_2961);
nor UO_319 (O_319,N_2984,N_2977);
and UO_320 (O_320,N_2960,N_2965);
and UO_321 (O_321,N_2952,N_2970);
or UO_322 (O_322,N_2948,N_2965);
nand UO_323 (O_323,N_2970,N_2994);
and UO_324 (O_324,N_2927,N_2934);
and UO_325 (O_325,N_2983,N_2965);
and UO_326 (O_326,N_2944,N_2931);
xor UO_327 (O_327,N_2938,N_2968);
xnor UO_328 (O_328,N_2945,N_2973);
nand UO_329 (O_329,N_2989,N_2953);
and UO_330 (O_330,N_2927,N_2974);
nor UO_331 (O_331,N_2948,N_2998);
nor UO_332 (O_332,N_2996,N_2982);
or UO_333 (O_333,N_2995,N_2958);
and UO_334 (O_334,N_2942,N_2953);
and UO_335 (O_335,N_2945,N_2952);
xor UO_336 (O_336,N_2965,N_2949);
and UO_337 (O_337,N_2980,N_2993);
nor UO_338 (O_338,N_2984,N_2943);
nand UO_339 (O_339,N_2940,N_2977);
xor UO_340 (O_340,N_2926,N_2983);
xor UO_341 (O_341,N_2931,N_2984);
nor UO_342 (O_342,N_2990,N_2985);
or UO_343 (O_343,N_2982,N_2999);
or UO_344 (O_344,N_2933,N_2965);
nor UO_345 (O_345,N_2981,N_2982);
and UO_346 (O_346,N_2950,N_2978);
xor UO_347 (O_347,N_2985,N_2957);
nand UO_348 (O_348,N_2978,N_2997);
xor UO_349 (O_349,N_2970,N_2966);
xor UO_350 (O_350,N_2997,N_2930);
and UO_351 (O_351,N_2988,N_2947);
or UO_352 (O_352,N_2948,N_2969);
nand UO_353 (O_353,N_2995,N_2939);
or UO_354 (O_354,N_2983,N_2950);
nor UO_355 (O_355,N_2928,N_2981);
or UO_356 (O_356,N_2952,N_2987);
xnor UO_357 (O_357,N_2978,N_2994);
and UO_358 (O_358,N_2947,N_2950);
nor UO_359 (O_359,N_2998,N_2956);
and UO_360 (O_360,N_2987,N_2926);
or UO_361 (O_361,N_2932,N_2939);
nand UO_362 (O_362,N_2982,N_2929);
and UO_363 (O_363,N_2966,N_2984);
or UO_364 (O_364,N_2965,N_2975);
and UO_365 (O_365,N_2928,N_2994);
nor UO_366 (O_366,N_2927,N_2998);
nor UO_367 (O_367,N_2970,N_2926);
and UO_368 (O_368,N_2961,N_2954);
xor UO_369 (O_369,N_2959,N_2968);
nand UO_370 (O_370,N_2951,N_2995);
and UO_371 (O_371,N_2978,N_2959);
xor UO_372 (O_372,N_2965,N_2978);
nand UO_373 (O_373,N_2959,N_2937);
xor UO_374 (O_374,N_2931,N_2957);
xnor UO_375 (O_375,N_2980,N_2972);
nand UO_376 (O_376,N_2968,N_2981);
xor UO_377 (O_377,N_2962,N_2941);
xnor UO_378 (O_378,N_2931,N_2971);
nor UO_379 (O_379,N_2930,N_2982);
nor UO_380 (O_380,N_2971,N_2933);
nor UO_381 (O_381,N_2985,N_2983);
nor UO_382 (O_382,N_2958,N_2989);
xor UO_383 (O_383,N_2940,N_2929);
nor UO_384 (O_384,N_2945,N_2976);
xnor UO_385 (O_385,N_2936,N_2983);
nand UO_386 (O_386,N_2977,N_2937);
and UO_387 (O_387,N_2985,N_2948);
xnor UO_388 (O_388,N_2960,N_2958);
nor UO_389 (O_389,N_2963,N_2957);
or UO_390 (O_390,N_2970,N_2961);
xor UO_391 (O_391,N_2980,N_2928);
nand UO_392 (O_392,N_2996,N_2980);
xor UO_393 (O_393,N_2996,N_2984);
xor UO_394 (O_394,N_2942,N_2975);
nand UO_395 (O_395,N_2948,N_2945);
or UO_396 (O_396,N_2966,N_2995);
nand UO_397 (O_397,N_2980,N_2965);
and UO_398 (O_398,N_2998,N_2942);
nand UO_399 (O_399,N_2953,N_2983);
and UO_400 (O_400,N_2955,N_2991);
and UO_401 (O_401,N_2960,N_2996);
or UO_402 (O_402,N_2949,N_2968);
or UO_403 (O_403,N_2973,N_2991);
and UO_404 (O_404,N_2930,N_2961);
or UO_405 (O_405,N_2961,N_2958);
nor UO_406 (O_406,N_2963,N_2925);
and UO_407 (O_407,N_2967,N_2995);
nand UO_408 (O_408,N_2989,N_2952);
xnor UO_409 (O_409,N_2925,N_2944);
xnor UO_410 (O_410,N_2969,N_2979);
or UO_411 (O_411,N_2967,N_2925);
and UO_412 (O_412,N_2999,N_2984);
or UO_413 (O_413,N_2985,N_2951);
nand UO_414 (O_414,N_2989,N_2961);
xor UO_415 (O_415,N_2977,N_2999);
or UO_416 (O_416,N_2948,N_2971);
and UO_417 (O_417,N_2955,N_2982);
nor UO_418 (O_418,N_2935,N_2949);
and UO_419 (O_419,N_2949,N_2999);
nor UO_420 (O_420,N_2957,N_2992);
nand UO_421 (O_421,N_2977,N_2926);
nor UO_422 (O_422,N_2984,N_2946);
or UO_423 (O_423,N_2942,N_2963);
nand UO_424 (O_424,N_2986,N_2975);
or UO_425 (O_425,N_2939,N_2967);
or UO_426 (O_426,N_2947,N_2966);
or UO_427 (O_427,N_2989,N_2983);
xor UO_428 (O_428,N_2989,N_2984);
xor UO_429 (O_429,N_2932,N_2946);
nor UO_430 (O_430,N_2971,N_2977);
nand UO_431 (O_431,N_2971,N_2961);
or UO_432 (O_432,N_2948,N_2993);
or UO_433 (O_433,N_2950,N_2977);
nor UO_434 (O_434,N_2991,N_2992);
nor UO_435 (O_435,N_2935,N_2955);
and UO_436 (O_436,N_2970,N_2940);
nor UO_437 (O_437,N_2968,N_2983);
nand UO_438 (O_438,N_2962,N_2927);
nor UO_439 (O_439,N_2969,N_2994);
xnor UO_440 (O_440,N_2985,N_2949);
nor UO_441 (O_441,N_2941,N_2936);
xnor UO_442 (O_442,N_2952,N_2955);
xor UO_443 (O_443,N_2969,N_2954);
or UO_444 (O_444,N_2956,N_2954);
xnor UO_445 (O_445,N_2954,N_2950);
or UO_446 (O_446,N_2963,N_2946);
nor UO_447 (O_447,N_2957,N_2928);
or UO_448 (O_448,N_2973,N_2962);
nand UO_449 (O_449,N_2999,N_2952);
nand UO_450 (O_450,N_2975,N_2996);
nor UO_451 (O_451,N_2953,N_2940);
or UO_452 (O_452,N_2941,N_2930);
or UO_453 (O_453,N_2970,N_2977);
xor UO_454 (O_454,N_2926,N_2959);
nor UO_455 (O_455,N_2981,N_2994);
or UO_456 (O_456,N_2994,N_2925);
nor UO_457 (O_457,N_2986,N_2970);
nor UO_458 (O_458,N_2961,N_2999);
xor UO_459 (O_459,N_2978,N_2966);
xnor UO_460 (O_460,N_2988,N_2952);
or UO_461 (O_461,N_2925,N_2950);
and UO_462 (O_462,N_2975,N_2963);
nor UO_463 (O_463,N_2935,N_2981);
and UO_464 (O_464,N_2926,N_2956);
or UO_465 (O_465,N_2950,N_2942);
or UO_466 (O_466,N_2937,N_2968);
nand UO_467 (O_467,N_2959,N_2934);
nor UO_468 (O_468,N_2937,N_2963);
and UO_469 (O_469,N_2961,N_2990);
nor UO_470 (O_470,N_2958,N_2927);
or UO_471 (O_471,N_2989,N_2972);
nand UO_472 (O_472,N_2957,N_2984);
xnor UO_473 (O_473,N_2936,N_2998);
nand UO_474 (O_474,N_2995,N_2984);
nand UO_475 (O_475,N_2936,N_2959);
or UO_476 (O_476,N_2981,N_2991);
nor UO_477 (O_477,N_2973,N_2940);
xnor UO_478 (O_478,N_2982,N_2939);
or UO_479 (O_479,N_2966,N_2943);
xnor UO_480 (O_480,N_2983,N_2932);
nor UO_481 (O_481,N_2925,N_2996);
nor UO_482 (O_482,N_2976,N_2936);
and UO_483 (O_483,N_2933,N_2987);
nor UO_484 (O_484,N_2990,N_2955);
and UO_485 (O_485,N_2944,N_2963);
nand UO_486 (O_486,N_2981,N_2936);
xor UO_487 (O_487,N_2992,N_2960);
nor UO_488 (O_488,N_2992,N_2985);
or UO_489 (O_489,N_2925,N_2940);
and UO_490 (O_490,N_2957,N_2929);
nand UO_491 (O_491,N_2983,N_2948);
and UO_492 (O_492,N_2948,N_2988);
nand UO_493 (O_493,N_2990,N_2945);
or UO_494 (O_494,N_2933,N_2964);
nor UO_495 (O_495,N_2988,N_2997);
or UO_496 (O_496,N_2925,N_2976);
xnor UO_497 (O_497,N_2997,N_2959);
nand UO_498 (O_498,N_2925,N_2995);
xor UO_499 (O_499,N_2953,N_2990);
endmodule