module basic_500_3000_500_5_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_229,In_476);
and U1 (N_1,In_109,In_387);
and U2 (N_2,In_116,In_250);
nand U3 (N_3,In_350,In_201);
and U4 (N_4,In_6,In_86);
nor U5 (N_5,In_432,In_453);
nand U6 (N_6,In_367,In_31);
and U7 (N_7,In_126,In_58);
and U8 (N_8,In_382,In_475);
or U9 (N_9,In_381,In_204);
nand U10 (N_10,In_422,In_273);
and U11 (N_11,In_154,In_437);
or U12 (N_12,In_397,In_323);
xnor U13 (N_13,In_117,In_107);
nand U14 (N_14,In_216,In_450);
nor U15 (N_15,In_416,In_182);
nor U16 (N_16,In_310,In_191);
nor U17 (N_17,In_15,In_158);
and U18 (N_18,In_365,In_359);
or U19 (N_19,In_288,In_67);
and U20 (N_20,In_334,In_366);
and U21 (N_21,In_13,In_73);
nand U22 (N_22,In_84,In_135);
xnor U23 (N_23,In_333,In_1);
nand U24 (N_24,In_51,In_344);
or U25 (N_25,In_332,In_414);
or U26 (N_26,In_452,In_42);
nand U27 (N_27,In_498,In_462);
and U28 (N_28,In_499,In_0);
nand U29 (N_29,In_9,In_436);
or U30 (N_30,In_386,In_209);
or U31 (N_31,In_120,In_411);
and U32 (N_32,In_32,In_183);
nor U33 (N_33,In_455,In_153);
or U34 (N_34,In_259,In_329);
and U35 (N_35,In_72,In_444);
or U36 (N_36,In_97,In_267);
or U37 (N_37,In_233,In_424);
or U38 (N_38,In_391,In_124);
or U39 (N_39,In_440,In_275);
nor U40 (N_40,In_426,In_188);
or U41 (N_41,In_266,In_52);
xnor U42 (N_42,In_61,In_316);
and U43 (N_43,In_203,In_459);
or U44 (N_44,In_244,In_430);
nor U45 (N_45,In_302,In_129);
or U46 (N_46,In_491,In_490);
and U47 (N_47,In_240,In_217);
nor U48 (N_48,In_243,In_138);
nor U49 (N_49,In_263,In_146);
and U50 (N_50,In_289,In_214);
and U51 (N_51,In_184,In_480);
or U52 (N_52,In_312,In_46);
or U53 (N_53,In_324,In_404);
xnor U54 (N_54,In_37,In_222);
or U55 (N_55,In_401,In_25);
nand U56 (N_56,In_252,In_136);
xnor U57 (N_57,In_26,In_375);
nor U58 (N_58,In_377,In_8);
nand U59 (N_59,In_68,In_379);
and U60 (N_60,In_82,In_446);
and U61 (N_61,In_396,In_331);
nor U62 (N_62,In_369,In_492);
and U63 (N_63,In_373,In_41);
and U64 (N_64,In_420,In_319);
and U65 (N_65,In_152,In_304);
and U66 (N_66,In_96,In_398);
and U67 (N_67,In_99,In_206);
nand U68 (N_68,In_100,In_338);
and U69 (N_69,In_296,In_322);
or U70 (N_70,In_258,In_286);
xnor U71 (N_71,In_363,In_193);
and U72 (N_72,In_24,In_56);
nor U73 (N_73,In_463,In_278);
or U74 (N_74,In_470,In_18);
nor U75 (N_75,In_134,In_468);
nand U76 (N_76,In_460,In_494);
and U77 (N_77,In_11,In_118);
nor U78 (N_78,In_208,In_142);
or U79 (N_79,In_91,In_469);
or U80 (N_80,In_357,In_106);
and U81 (N_81,In_320,In_165);
and U82 (N_82,In_147,In_140);
nand U83 (N_83,In_171,In_264);
nor U84 (N_84,In_370,In_95);
nand U85 (N_85,In_5,In_125);
and U86 (N_86,In_465,In_219);
and U87 (N_87,In_383,In_197);
or U88 (N_88,In_283,In_242);
and U89 (N_89,In_408,In_181);
or U90 (N_90,In_167,In_327);
nand U91 (N_91,In_122,In_49);
or U92 (N_92,In_128,In_248);
nand U93 (N_93,In_212,In_364);
nor U94 (N_94,In_425,In_478);
or U95 (N_95,In_23,In_335);
and U96 (N_96,In_488,In_246);
nor U97 (N_97,In_16,In_35);
xnor U98 (N_98,In_284,In_464);
or U99 (N_99,In_40,In_290);
nand U100 (N_100,In_281,In_98);
and U101 (N_101,In_340,In_336);
or U102 (N_102,In_265,In_393);
nand U103 (N_103,In_137,In_458);
nor U104 (N_104,In_345,In_38);
or U105 (N_105,In_199,In_225);
and U106 (N_106,In_55,In_441);
nor U107 (N_107,In_64,In_256);
nand U108 (N_108,In_141,In_443);
or U109 (N_109,In_287,In_211);
and U110 (N_110,In_314,In_74);
nor U111 (N_111,In_223,In_410);
and U112 (N_112,In_173,In_176);
or U113 (N_113,In_105,In_485);
nor U114 (N_114,In_348,In_221);
nor U115 (N_115,In_166,In_368);
nor U116 (N_116,In_151,In_245);
and U117 (N_117,In_90,In_268);
and U118 (N_118,In_421,In_481);
nand U119 (N_119,In_433,In_315);
and U120 (N_120,In_189,In_295);
and U121 (N_121,In_402,In_418);
nand U122 (N_122,In_356,In_92);
nor U123 (N_123,In_317,In_307);
or U124 (N_124,In_439,In_353);
and U125 (N_125,In_119,In_164);
or U126 (N_126,In_10,In_123);
nor U127 (N_127,In_54,In_360);
and U128 (N_128,In_328,In_354);
or U129 (N_129,In_133,In_351);
nand U130 (N_130,In_497,In_409);
nor U131 (N_131,In_301,In_305);
nor U132 (N_132,In_371,In_79);
nor U133 (N_133,In_130,In_113);
nand U134 (N_134,In_447,In_269);
or U135 (N_135,In_487,In_361);
nor U136 (N_136,In_438,In_484);
or U137 (N_137,In_472,In_190);
or U138 (N_138,In_80,In_419);
nor U139 (N_139,In_271,In_456);
nand U140 (N_140,In_406,In_241);
nand U141 (N_141,In_270,In_474);
and U142 (N_142,In_358,In_200);
nor U143 (N_143,In_291,In_489);
nand U144 (N_144,In_260,In_234);
nor U145 (N_145,In_347,In_461);
nor U146 (N_146,In_399,In_34);
or U147 (N_147,In_4,In_179);
and U148 (N_148,In_466,In_448);
nor U149 (N_149,In_28,In_362);
nand U150 (N_150,In_405,In_44);
nor U151 (N_151,In_19,In_88);
nor U152 (N_152,In_161,In_110);
and U153 (N_153,In_285,In_149);
nor U154 (N_154,In_477,In_14);
and U155 (N_155,In_303,In_308);
nor U156 (N_156,In_93,In_257);
nand U157 (N_157,In_435,In_277);
nor U158 (N_158,In_70,In_394);
nand U159 (N_159,In_374,In_112);
nor U160 (N_160,In_186,In_162);
or U161 (N_161,In_104,In_247);
or U162 (N_162,In_376,In_407);
nand U163 (N_163,In_218,In_321);
and U164 (N_164,In_69,In_48);
nand U165 (N_165,In_220,In_207);
nand U166 (N_166,In_372,In_157);
nor U167 (N_167,In_294,In_22);
and U168 (N_168,In_75,In_232);
nand U169 (N_169,In_213,In_103);
and U170 (N_170,In_299,In_467);
or U171 (N_171,In_325,In_71);
nor U172 (N_172,In_2,In_400);
or U173 (N_173,In_76,In_342);
nor U174 (N_174,In_449,In_7);
or U175 (N_175,In_349,In_168);
nand U176 (N_176,In_63,In_43);
nor U177 (N_177,In_27,In_471);
xnor U178 (N_178,In_427,In_50);
and U179 (N_179,In_187,In_169);
or U180 (N_180,In_280,In_493);
nor U181 (N_181,In_159,In_238);
nor U182 (N_182,In_272,In_177);
nand U183 (N_183,In_384,In_174);
nor U184 (N_184,In_235,In_318);
and U185 (N_185,In_415,In_388);
and U186 (N_186,In_196,In_160);
and U187 (N_187,In_306,In_457);
nand U188 (N_188,In_226,In_417);
nor U189 (N_189,In_343,In_194);
nand U190 (N_190,In_155,In_380);
nor U191 (N_191,In_127,In_111);
nor U192 (N_192,In_139,In_451);
or U193 (N_193,In_121,In_81);
or U194 (N_194,In_431,In_65);
and U195 (N_195,In_300,In_442);
or U196 (N_196,In_428,In_198);
nor U197 (N_197,In_389,In_101);
nand U198 (N_198,In_195,In_346);
nand U199 (N_199,In_311,In_352);
and U200 (N_200,In_131,In_224);
or U201 (N_201,In_205,In_326);
and U202 (N_202,In_403,In_77);
and U203 (N_203,In_94,In_87);
nand U204 (N_204,In_175,In_85);
nand U205 (N_205,In_172,In_282);
xnor U206 (N_206,In_3,In_279);
or U207 (N_207,In_313,In_115);
and U208 (N_208,In_292,In_255);
nand U209 (N_209,In_36,In_202);
and U210 (N_210,In_337,In_66);
nand U211 (N_211,In_108,In_385);
or U212 (N_212,In_341,In_156);
and U213 (N_213,In_145,In_413);
nor U214 (N_214,In_170,In_330);
nor U215 (N_215,In_228,In_47);
nor U216 (N_216,In_21,In_412);
nand U217 (N_217,In_339,In_274);
and U218 (N_218,In_185,In_150);
xnor U219 (N_219,In_395,In_215);
or U220 (N_220,In_293,In_180);
or U221 (N_221,In_59,In_178);
nand U222 (N_222,In_17,In_83);
or U223 (N_223,In_78,In_227);
or U224 (N_224,In_53,In_309);
and U225 (N_225,In_495,In_251);
or U226 (N_226,In_132,In_486);
nor U227 (N_227,In_392,In_445);
nand U228 (N_228,In_479,In_57);
nand U229 (N_229,In_473,In_163);
or U230 (N_230,In_231,In_355);
and U231 (N_231,In_62,In_236);
or U232 (N_232,In_262,In_482);
nand U233 (N_233,In_423,In_192);
nor U234 (N_234,In_12,In_390);
or U235 (N_235,In_148,In_210);
nand U236 (N_236,In_230,In_297);
or U237 (N_237,In_429,In_276);
nor U238 (N_238,In_45,In_39);
and U239 (N_239,In_20,In_60);
nand U240 (N_240,In_144,In_114);
or U241 (N_241,In_298,In_261);
or U242 (N_242,In_454,In_89);
nand U243 (N_243,In_254,In_29);
and U244 (N_244,In_143,In_253);
nand U245 (N_245,In_249,In_434);
nand U246 (N_246,In_496,In_483);
xor U247 (N_247,In_378,In_33);
nand U248 (N_248,In_237,In_30);
or U249 (N_249,In_239,In_102);
and U250 (N_250,In_96,In_173);
nor U251 (N_251,In_439,In_303);
nor U252 (N_252,In_434,In_8);
nand U253 (N_253,In_6,In_317);
or U254 (N_254,In_294,In_368);
and U255 (N_255,In_448,In_322);
nand U256 (N_256,In_419,In_266);
nor U257 (N_257,In_47,In_273);
nor U258 (N_258,In_210,In_484);
and U259 (N_259,In_86,In_280);
and U260 (N_260,In_91,In_377);
or U261 (N_261,In_197,In_158);
nand U262 (N_262,In_449,In_416);
nand U263 (N_263,In_318,In_10);
and U264 (N_264,In_288,In_422);
and U265 (N_265,In_225,In_129);
or U266 (N_266,In_103,In_452);
and U267 (N_267,In_279,In_380);
or U268 (N_268,In_432,In_147);
nor U269 (N_269,In_119,In_178);
nand U270 (N_270,In_428,In_179);
nand U271 (N_271,In_200,In_331);
and U272 (N_272,In_462,In_53);
or U273 (N_273,In_154,In_85);
nor U274 (N_274,In_282,In_247);
and U275 (N_275,In_462,In_230);
or U276 (N_276,In_211,In_427);
and U277 (N_277,In_70,In_244);
nor U278 (N_278,In_281,In_172);
nor U279 (N_279,In_356,In_6);
and U280 (N_280,In_303,In_13);
nor U281 (N_281,In_315,In_413);
nor U282 (N_282,In_341,In_330);
and U283 (N_283,In_13,In_200);
nor U284 (N_284,In_136,In_416);
nor U285 (N_285,In_303,In_9);
nand U286 (N_286,In_423,In_2);
nor U287 (N_287,In_340,In_91);
or U288 (N_288,In_285,In_372);
and U289 (N_289,In_198,In_436);
nor U290 (N_290,In_206,In_121);
or U291 (N_291,In_496,In_285);
nand U292 (N_292,In_336,In_393);
nand U293 (N_293,In_472,In_493);
or U294 (N_294,In_384,In_63);
nor U295 (N_295,In_145,In_81);
and U296 (N_296,In_366,In_344);
nor U297 (N_297,In_318,In_309);
or U298 (N_298,In_364,In_421);
or U299 (N_299,In_338,In_314);
nor U300 (N_300,In_444,In_231);
or U301 (N_301,In_168,In_13);
and U302 (N_302,In_498,In_401);
and U303 (N_303,In_414,In_107);
or U304 (N_304,In_282,In_467);
xor U305 (N_305,In_473,In_107);
and U306 (N_306,In_467,In_194);
or U307 (N_307,In_355,In_215);
or U308 (N_308,In_256,In_236);
nor U309 (N_309,In_176,In_373);
nor U310 (N_310,In_169,In_20);
nor U311 (N_311,In_429,In_255);
nor U312 (N_312,In_303,In_256);
or U313 (N_313,In_421,In_34);
nand U314 (N_314,In_329,In_348);
nand U315 (N_315,In_236,In_119);
and U316 (N_316,In_487,In_109);
nor U317 (N_317,In_374,In_268);
and U318 (N_318,In_69,In_415);
or U319 (N_319,In_21,In_439);
xnor U320 (N_320,In_484,In_264);
nor U321 (N_321,In_175,In_69);
and U322 (N_322,In_393,In_353);
nor U323 (N_323,In_119,In_303);
nand U324 (N_324,In_223,In_224);
and U325 (N_325,In_268,In_421);
nand U326 (N_326,In_351,In_357);
xnor U327 (N_327,In_382,In_242);
nor U328 (N_328,In_48,In_19);
nand U329 (N_329,In_252,In_105);
or U330 (N_330,In_429,In_80);
nor U331 (N_331,In_18,In_297);
and U332 (N_332,In_404,In_14);
and U333 (N_333,In_341,In_289);
or U334 (N_334,In_406,In_249);
nor U335 (N_335,In_423,In_275);
or U336 (N_336,In_320,In_364);
and U337 (N_337,In_478,In_316);
or U338 (N_338,In_463,In_112);
or U339 (N_339,In_211,In_300);
nand U340 (N_340,In_318,In_55);
xnor U341 (N_341,In_356,In_281);
nor U342 (N_342,In_70,In_457);
and U343 (N_343,In_2,In_322);
nand U344 (N_344,In_227,In_476);
and U345 (N_345,In_377,In_353);
and U346 (N_346,In_117,In_106);
nor U347 (N_347,In_288,In_433);
nor U348 (N_348,In_63,In_23);
nor U349 (N_349,In_148,In_165);
nor U350 (N_350,In_374,In_445);
or U351 (N_351,In_403,In_337);
and U352 (N_352,In_397,In_8);
and U353 (N_353,In_5,In_173);
nand U354 (N_354,In_8,In_472);
nand U355 (N_355,In_130,In_288);
and U356 (N_356,In_40,In_244);
nand U357 (N_357,In_330,In_383);
and U358 (N_358,In_8,In_205);
or U359 (N_359,In_320,In_151);
nor U360 (N_360,In_256,In_205);
nand U361 (N_361,In_190,In_269);
and U362 (N_362,In_76,In_354);
xor U363 (N_363,In_211,In_190);
or U364 (N_364,In_278,In_150);
nand U365 (N_365,In_245,In_346);
xnor U366 (N_366,In_129,In_333);
nand U367 (N_367,In_432,In_223);
and U368 (N_368,In_304,In_283);
and U369 (N_369,In_218,In_302);
nand U370 (N_370,In_277,In_40);
nand U371 (N_371,In_209,In_156);
and U372 (N_372,In_401,In_399);
nor U373 (N_373,In_256,In_484);
nand U374 (N_374,In_429,In_138);
nand U375 (N_375,In_179,In_483);
nand U376 (N_376,In_299,In_358);
and U377 (N_377,In_235,In_213);
nand U378 (N_378,In_45,In_70);
and U379 (N_379,In_398,In_344);
or U380 (N_380,In_433,In_76);
and U381 (N_381,In_189,In_110);
or U382 (N_382,In_91,In_442);
nor U383 (N_383,In_283,In_27);
nand U384 (N_384,In_352,In_409);
or U385 (N_385,In_4,In_136);
and U386 (N_386,In_128,In_409);
nand U387 (N_387,In_149,In_388);
or U388 (N_388,In_2,In_269);
nor U389 (N_389,In_382,In_484);
and U390 (N_390,In_88,In_420);
nor U391 (N_391,In_335,In_166);
nor U392 (N_392,In_375,In_435);
nor U393 (N_393,In_316,In_95);
nor U394 (N_394,In_113,In_483);
and U395 (N_395,In_405,In_102);
or U396 (N_396,In_172,In_464);
or U397 (N_397,In_70,In_429);
nand U398 (N_398,In_116,In_449);
or U399 (N_399,In_175,In_138);
nand U400 (N_400,In_306,In_125);
or U401 (N_401,In_79,In_359);
or U402 (N_402,In_350,In_72);
xor U403 (N_403,In_108,In_21);
nand U404 (N_404,In_459,In_361);
nand U405 (N_405,In_82,In_387);
or U406 (N_406,In_404,In_209);
nand U407 (N_407,In_196,In_329);
or U408 (N_408,In_106,In_409);
nor U409 (N_409,In_268,In_48);
nand U410 (N_410,In_248,In_476);
nand U411 (N_411,In_197,In_234);
and U412 (N_412,In_101,In_113);
and U413 (N_413,In_34,In_50);
nor U414 (N_414,In_262,In_309);
and U415 (N_415,In_25,In_495);
nor U416 (N_416,In_22,In_453);
and U417 (N_417,In_371,In_9);
nor U418 (N_418,In_110,In_346);
or U419 (N_419,In_295,In_110);
nand U420 (N_420,In_329,In_30);
and U421 (N_421,In_444,In_243);
or U422 (N_422,In_61,In_194);
and U423 (N_423,In_332,In_489);
nor U424 (N_424,In_391,In_157);
nand U425 (N_425,In_332,In_376);
nor U426 (N_426,In_496,In_214);
nand U427 (N_427,In_174,In_127);
nand U428 (N_428,In_333,In_11);
nor U429 (N_429,In_313,In_74);
nor U430 (N_430,In_130,In_316);
or U431 (N_431,In_65,In_496);
and U432 (N_432,In_276,In_158);
nor U433 (N_433,In_312,In_209);
nor U434 (N_434,In_163,In_73);
xor U435 (N_435,In_473,In_365);
nor U436 (N_436,In_292,In_254);
nor U437 (N_437,In_206,In_252);
nor U438 (N_438,In_455,In_55);
and U439 (N_439,In_459,In_174);
or U440 (N_440,In_164,In_196);
nor U441 (N_441,In_485,In_333);
nor U442 (N_442,In_257,In_304);
or U443 (N_443,In_273,In_140);
or U444 (N_444,In_468,In_430);
nor U445 (N_445,In_318,In_321);
or U446 (N_446,In_401,In_143);
nor U447 (N_447,In_322,In_19);
and U448 (N_448,In_491,In_165);
and U449 (N_449,In_403,In_239);
and U450 (N_450,In_51,In_186);
and U451 (N_451,In_38,In_113);
nand U452 (N_452,In_499,In_56);
xor U453 (N_453,In_168,In_417);
nor U454 (N_454,In_14,In_42);
or U455 (N_455,In_292,In_231);
or U456 (N_456,In_95,In_43);
nor U457 (N_457,In_266,In_317);
and U458 (N_458,In_318,In_366);
nor U459 (N_459,In_378,In_92);
and U460 (N_460,In_156,In_98);
or U461 (N_461,In_375,In_284);
nand U462 (N_462,In_449,In_123);
nor U463 (N_463,In_400,In_255);
and U464 (N_464,In_62,In_3);
nand U465 (N_465,In_219,In_410);
or U466 (N_466,In_197,In_376);
nand U467 (N_467,In_357,In_10);
nor U468 (N_468,In_107,In_162);
or U469 (N_469,In_271,In_255);
or U470 (N_470,In_458,In_199);
and U471 (N_471,In_457,In_148);
nor U472 (N_472,In_5,In_408);
and U473 (N_473,In_21,In_57);
nor U474 (N_474,In_332,In_369);
nor U475 (N_475,In_192,In_143);
or U476 (N_476,In_250,In_437);
xnor U477 (N_477,In_170,In_413);
nand U478 (N_478,In_241,In_343);
and U479 (N_479,In_64,In_27);
nand U480 (N_480,In_302,In_88);
nand U481 (N_481,In_230,In_83);
nor U482 (N_482,In_328,In_250);
nand U483 (N_483,In_69,In_200);
and U484 (N_484,In_345,In_56);
and U485 (N_485,In_91,In_186);
and U486 (N_486,In_43,In_199);
nor U487 (N_487,In_416,In_398);
and U488 (N_488,In_219,In_394);
and U489 (N_489,In_285,In_53);
nand U490 (N_490,In_288,In_414);
or U491 (N_491,In_98,In_254);
nand U492 (N_492,In_425,In_412);
nor U493 (N_493,In_186,In_145);
nor U494 (N_494,In_443,In_364);
nor U495 (N_495,In_261,In_114);
or U496 (N_496,In_298,In_204);
nand U497 (N_497,In_1,In_432);
nand U498 (N_498,In_407,In_351);
or U499 (N_499,In_81,In_144);
nor U500 (N_500,In_371,In_319);
nor U501 (N_501,In_59,In_330);
nand U502 (N_502,In_453,In_486);
nor U503 (N_503,In_128,In_55);
or U504 (N_504,In_316,In_401);
and U505 (N_505,In_159,In_417);
and U506 (N_506,In_441,In_424);
or U507 (N_507,In_181,In_375);
nand U508 (N_508,In_170,In_362);
and U509 (N_509,In_353,In_145);
or U510 (N_510,In_244,In_236);
xor U511 (N_511,In_63,In_95);
and U512 (N_512,In_135,In_161);
nand U513 (N_513,In_54,In_325);
nor U514 (N_514,In_127,In_248);
nand U515 (N_515,In_395,In_361);
or U516 (N_516,In_264,In_295);
or U517 (N_517,In_161,In_354);
nor U518 (N_518,In_276,In_107);
or U519 (N_519,In_156,In_23);
nor U520 (N_520,In_191,In_286);
and U521 (N_521,In_325,In_193);
or U522 (N_522,In_324,In_135);
nor U523 (N_523,In_312,In_0);
or U524 (N_524,In_196,In_226);
nor U525 (N_525,In_28,In_497);
nand U526 (N_526,In_232,In_238);
nand U527 (N_527,In_323,In_12);
nand U528 (N_528,In_80,In_16);
or U529 (N_529,In_287,In_56);
and U530 (N_530,In_474,In_102);
xor U531 (N_531,In_383,In_275);
nor U532 (N_532,In_2,In_175);
or U533 (N_533,In_339,In_356);
nor U534 (N_534,In_81,In_137);
xnor U535 (N_535,In_340,In_441);
nor U536 (N_536,In_305,In_269);
or U537 (N_537,In_80,In_131);
nand U538 (N_538,In_328,In_471);
or U539 (N_539,In_92,In_283);
and U540 (N_540,In_222,In_178);
or U541 (N_541,In_370,In_121);
or U542 (N_542,In_224,In_146);
or U543 (N_543,In_405,In_5);
nor U544 (N_544,In_48,In_235);
and U545 (N_545,In_398,In_6);
nor U546 (N_546,In_423,In_444);
and U547 (N_547,In_473,In_326);
or U548 (N_548,In_66,In_251);
and U549 (N_549,In_177,In_302);
or U550 (N_550,In_127,In_78);
nand U551 (N_551,In_416,In_409);
nand U552 (N_552,In_238,In_432);
and U553 (N_553,In_272,In_259);
or U554 (N_554,In_249,In_133);
nor U555 (N_555,In_103,In_40);
nand U556 (N_556,In_126,In_65);
or U557 (N_557,In_186,In_160);
and U558 (N_558,In_337,In_366);
nand U559 (N_559,In_321,In_232);
and U560 (N_560,In_61,In_66);
nand U561 (N_561,In_59,In_362);
nor U562 (N_562,In_314,In_115);
and U563 (N_563,In_105,In_77);
and U564 (N_564,In_302,In_176);
or U565 (N_565,In_19,In_265);
nand U566 (N_566,In_458,In_118);
or U567 (N_567,In_461,In_53);
nor U568 (N_568,In_35,In_268);
nand U569 (N_569,In_166,In_45);
xor U570 (N_570,In_216,In_468);
nand U571 (N_571,In_312,In_399);
or U572 (N_572,In_4,In_212);
or U573 (N_573,In_245,In_143);
nor U574 (N_574,In_96,In_367);
nor U575 (N_575,In_139,In_274);
xor U576 (N_576,In_336,In_20);
or U577 (N_577,In_228,In_16);
nand U578 (N_578,In_277,In_222);
nand U579 (N_579,In_229,In_370);
nand U580 (N_580,In_155,In_430);
xnor U581 (N_581,In_152,In_444);
or U582 (N_582,In_293,In_28);
or U583 (N_583,In_192,In_465);
nand U584 (N_584,In_388,In_463);
or U585 (N_585,In_262,In_221);
or U586 (N_586,In_98,In_306);
xor U587 (N_587,In_18,In_247);
nand U588 (N_588,In_197,In_360);
nand U589 (N_589,In_484,In_189);
and U590 (N_590,In_426,In_131);
or U591 (N_591,In_119,In_83);
and U592 (N_592,In_353,In_361);
or U593 (N_593,In_419,In_460);
nor U594 (N_594,In_356,In_222);
nand U595 (N_595,In_72,In_193);
nor U596 (N_596,In_170,In_92);
xnor U597 (N_597,In_210,In_132);
nor U598 (N_598,In_427,In_79);
or U599 (N_599,In_285,In_475);
or U600 (N_600,N_118,N_511);
or U601 (N_601,N_250,N_396);
nor U602 (N_602,N_484,N_388);
nand U603 (N_603,N_479,N_443);
nor U604 (N_604,N_235,N_94);
nand U605 (N_605,N_150,N_48);
and U606 (N_606,N_442,N_253);
and U607 (N_607,N_317,N_13);
nand U608 (N_608,N_402,N_41);
nand U609 (N_609,N_587,N_262);
and U610 (N_610,N_117,N_112);
or U611 (N_611,N_31,N_466);
or U612 (N_612,N_504,N_387);
or U613 (N_613,N_173,N_143);
or U614 (N_614,N_391,N_208);
nand U615 (N_615,N_97,N_25);
nor U616 (N_616,N_152,N_70);
or U617 (N_617,N_293,N_210);
nor U618 (N_618,N_80,N_404);
and U619 (N_619,N_195,N_330);
nor U620 (N_620,N_147,N_551);
and U621 (N_621,N_69,N_267);
or U622 (N_622,N_538,N_176);
nor U623 (N_623,N_216,N_483);
and U624 (N_624,N_289,N_241);
and U625 (N_625,N_40,N_542);
nand U626 (N_626,N_554,N_230);
and U627 (N_627,N_64,N_299);
and U628 (N_628,N_541,N_477);
or U629 (N_629,N_408,N_249);
or U630 (N_630,N_3,N_468);
or U631 (N_631,N_180,N_393);
or U632 (N_632,N_570,N_586);
and U633 (N_633,N_548,N_313);
nand U634 (N_634,N_578,N_157);
nand U635 (N_635,N_174,N_7);
or U636 (N_636,N_529,N_595);
nand U637 (N_637,N_426,N_342);
or U638 (N_638,N_138,N_213);
nand U639 (N_639,N_264,N_215);
or U640 (N_640,N_302,N_111);
or U641 (N_641,N_58,N_95);
nand U642 (N_642,N_236,N_370);
xnor U643 (N_643,N_107,N_364);
or U644 (N_644,N_35,N_51);
or U645 (N_645,N_355,N_188);
nand U646 (N_646,N_133,N_557);
nor U647 (N_647,N_353,N_32);
or U648 (N_648,N_247,N_261);
nand U649 (N_649,N_131,N_458);
or U650 (N_650,N_81,N_211);
and U651 (N_651,N_294,N_75);
nand U652 (N_652,N_417,N_266);
nand U653 (N_653,N_312,N_598);
and U654 (N_654,N_145,N_515);
nor U655 (N_655,N_411,N_439);
and U656 (N_656,N_183,N_192);
or U657 (N_657,N_440,N_27);
or U658 (N_658,N_462,N_190);
nand U659 (N_659,N_52,N_221);
nor U660 (N_660,N_55,N_18);
and U661 (N_661,N_49,N_418);
or U662 (N_662,N_358,N_321);
nor U663 (N_663,N_19,N_4);
or U664 (N_664,N_105,N_543);
nand U665 (N_665,N_375,N_185);
nand U666 (N_666,N_576,N_155);
nand U667 (N_667,N_121,N_296);
and U668 (N_668,N_244,N_124);
or U669 (N_669,N_327,N_405);
nand U670 (N_670,N_220,N_571);
and U671 (N_671,N_78,N_148);
or U672 (N_672,N_243,N_574);
and U673 (N_673,N_562,N_591);
or U674 (N_674,N_189,N_372);
and U675 (N_675,N_416,N_384);
nor U676 (N_676,N_360,N_378);
nor U677 (N_677,N_245,N_257);
nor U678 (N_678,N_345,N_454);
nand U679 (N_679,N_240,N_500);
or U680 (N_680,N_565,N_269);
nor U681 (N_681,N_531,N_430);
nor U682 (N_682,N_386,N_589);
nor U683 (N_683,N_274,N_219);
and U684 (N_684,N_125,N_34);
nor U685 (N_685,N_399,N_476);
nor U686 (N_686,N_456,N_184);
and U687 (N_687,N_77,N_37);
nand U688 (N_688,N_11,N_268);
and U689 (N_689,N_169,N_460);
nand U690 (N_690,N_151,N_343);
nand U691 (N_691,N_425,N_59);
nand U692 (N_692,N_301,N_170);
and U693 (N_693,N_42,N_528);
nand U694 (N_694,N_304,N_214);
nor U695 (N_695,N_222,N_305);
or U696 (N_696,N_471,N_365);
nor U697 (N_697,N_597,N_463);
nand U698 (N_698,N_316,N_287);
or U699 (N_699,N_246,N_369);
nand U700 (N_700,N_9,N_420);
or U701 (N_701,N_331,N_263);
and U702 (N_702,N_172,N_252);
nor U703 (N_703,N_68,N_567);
or U704 (N_704,N_427,N_113);
nand U705 (N_705,N_76,N_340);
nor U706 (N_706,N_14,N_102);
and U707 (N_707,N_90,N_580);
or U708 (N_708,N_315,N_10);
or U709 (N_709,N_447,N_448);
and U710 (N_710,N_564,N_127);
nor U711 (N_711,N_596,N_5);
and U712 (N_712,N_444,N_575);
or U713 (N_713,N_149,N_497);
or U714 (N_714,N_487,N_478);
and U715 (N_715,N_383,N_421);
and U716 (N_716,N_446,N_86);
and U717 (N_717,N_50,N_135);
and U718 (N_718,N_381,N_457);
or U719 (N_719,N_306,N_171);
nor U720 (N_720,N_319,N_368);
and U721 (N_721,N_482,N_218);
nand U722 (N_722,N_473,N_436);
and U723 (N_723,N_38,N_433);
nor U724 (N_724,N_311,N_196);
or U725 (N_725,N_415,N_488);
or U726 (N_726,N_126,N_165);
and U727 (N_727,N_226,N_177);
and U728 (N_728,N_322,N_517);
nand U729 (N_729,N_401,N_17);
or U730 (N_730,N_271,N_445);
or U731 (N_731,N_480,N_568);
and U732 (N_732,N_525,N_297);
or U733 (N_733,N_89,N_242);
and U734 (N_734,N_485,N_140);
nand U735 (N_735,N_361,N_83);
and U736 (N_736,N_536,N_545);
xnor U737 (N_737,N_279,N_103);
nor U738 (N_738,N_424,N_579);
or U739 (N_739,N_367,N_338);
and U740 (N_740,N_470,N_167);
and U741 (N_741,N_63,N_435);
nand U742 (N_742,N_46,N_431);
or U743 (N_743,N_339,N_258);
and U744 (N_744,N_203,N_153);
or U745 (N_745,N_337,N_530);
nor U746 (N_746,N_144,N_594);
or U747 (N_747,N_512,N_494);
nor U748 (N_748,N_204,N_374);
and U749 (N_749,N_534,N_228);
or U750 (N_750,N_231,N_397);
nand U751 (N_751,N_572,N_201);
nor U752 (N_752,N_292,N_182);
nand U753 (N_753,N_409,N_286);
and U754 (N_754,N_569,N_585);
or U755 (N_755,N_533,N_560);
and U756 (N_756,N_524,N_505);
or U757 (N_757,N_300,N_164);
and U758 (N_758,N_429,N_283);
nand U759 (N_759,N_110,N_285);
nor U760 (N_760,N_577,N_93);
or U761 (N_761,N_566,N_407);
nor U762 (N_762,N_106,N_518);
or U763 (N_763,N_581,N_362);
xor U764 (N_764,N_356,N_472);
nand U765 (N_765,N_239,N_395);
nor U766 (N_766,N_281,N_282);
or U767 (N_767,N_158,N_209);
or U768 (N_768,N_256,N_376);
and U769 (N_769,N_325,N_563);
and U770 (N_770,N_582,N_455);
nand U771 (N_771,N_16,N_537);
and U772 (N_772,N_521,N_212);
nor U773 (N_773,N_84,N_166);
nand U774 (N_774,N_277,N_71);
nand U775 (N_775,N_116,N_357);
nand U776 (N_776,N_179,N_248);
nand U777 (N_777,N_62,N_108);
or U778 (N_778,N_584,N_509);
nor U779 (N_779,N_495,N_120);
or U780 (N_780,N_298,N_66);
and U781 (N_781,N_186,N_82);
nand U782 (N_782,N_432,N_516);
nor U783 (N_783,N_168,N_520);
nor U784 (N_784,N_161,N_15);
or U785 (N_785,N_385,N_233);
nor U786 (N_786,N_474,N_229);
or U787 (N_787,N_328,N_552);
or U788 (N_788,N_22,N_26);
nand U789 (N_789,N_53,N_308);
nand U790 (N_790,N_514,N_532);
and U791 (N_791,N_503,N_160);
and U792 (N_792,N_441,N_96);
and U793 (N_793,N_414,N_100);
nand U794 (N_794,N_137,N_544);
nand U795 (N_795,N_163,N_217);
nor U796 (N_796,N_352,N_136);
or U797 (N_797,N_232,N_398);
nand U798 (N_798,N_555,N_295);
and U799 (N_799,N_141,N_593);
or U800 (N_800,N_291,N_187);
and U801 (N_801,N_47,N_67);
and U802 (N_802,N_23,N_382);
and U803 (N_803,N_104,N_335);
nor U804 (N_804,N_114,N_119);
nand U805 (N_805,N_464,N_540);
nor U806 (N_806,N_499,N_205);
or U807 (N_807,N_154,N_227);
or U808 (N_808,N_175,N_599);
and U809 (N_809,N_288,N_8);
and U810 (N_810,N_115,N_225);
nand U811 (N_811,N_486,N_556);
or U812 (N_812,N_389,N_351);
nor U813 (N_813,N_0,N_43);
or U814 (N_814,N_92,N_363);
or U815 (N_815,N_129,N_6);
nor U816 (N_816,N_465,N_583);
or U817 (N_817,N_379,N_373);
nand U818 (N_818,N_347,N_510);
nor U819 (N_819,N_539,N_492);
and U820 (N_820,N_491,N_506);
and U821 (N_821,N_501,N_392);
nor U822 (N_822,N_344,N_197);
or U823 (N_823,N_469,N_394);
and U824 (N_824,N_284,N_251);
nor U825 (N_825,N_198,N_181);
or U826 (N_826,N_24,N_526);
nor U827 (N_827,N_36,N_475);
or U828 (N_828,N_309,N_20);
nor U829 (N_829,N_65,N_21);
or U830 (N_830,N_142,N_318);
nand U831 (N_831,N_553,N_273);
nor U832 (N_832,N_265,N_303);
nand U833 (N_833,N_275,N_12);
or U834 (N_834,N_489,N_276);
or U835 (N_835,N_224,N_419);
or U836 (N_836,N_238,N_206);
nor U837 (N_837,N_332,N_450);
xnor U838 (N_838,N_324,N_422);
nand U839 (N_839,N_91,N_508);
or U840 (N_840,N_290,N_1);
nor U841 (N_841,N_326,N_354);
nand U842 (N_842,N_449,N_44);
nor U843 (N_843,N_310,N_314);
and U844 (N_844,N_333,N_380);
nand U845 (N_845,N_132,N_280);
nor U846 (N_846,N_254,N_403);
or U847 (N_847,N_202,N_346);
nor U848 (N_848,N_377,N_79);
nand U849 (N_849,N_109,N_139);
or U850 (N_850,N_359,N_87);
or U851 (N_851,N_334,N_341);
nor U852 (N_852,N_60,N_54);
or U853 (N_853,N_350,N_412);
and U854 (N_854,N_255,N_423);
nor U855 (N_855,N_260,N_307);
nand U856 (N_856,N_437,N_45);
and U857 (N_857,N_101,N_452);
or U858 (N_858,N_336,N_490);
or U859 (N_859,N_193,N_33);
nand U860 (N_860,N_191,N_592);
or U861 (N_861,N_547,N_535);
nor U862 (N_862,N_467,N_73);
nand U863 (N_863,N_371,N_406);
nor U864 (N_864,N_522,N_428);
nand U865 (N_865,N_349,N_200);
nor U866 (N_866,N_159,N_493);
or U867 (N_867,N_270,N_519);
xnor U868 (N_868,N_527,N_549);
nor U869 (N_869,N_234,N_323);
xor U870 (N_870,N_28,N_588);
and U871 (N_871,N_146,N_453);
nor U872 (N_872,N_134,N_558);
nor U873 (N_873,N_502,N_194);
or U874 (N_874,N_57,N_590);
and U875 (N_875,N_178,N_390);
nand U876 (N_876,N_413,N_85);
nand U877 (N_877,N_272,N_278);
xor U878 (N_878,N_523,N_573);
nor U879 (N_879,N_459,N_156);
nand U880 (N_880,N_259,N_400);
nand U881 (N_881,N_498,N_99);
or U882 (N_882,N_559,N_481);
or U883 (N_883,N_207,N_434);
and U884 (N_884,N_128,N_513);
and U885 (N_885,N_56,N_88);
nor U886 (N_886,N_320,N_438);
nor U887 (N_887,N_30,N_162);
nor U888 (N_888,N_561,N_74);
nand U889 (N_889,N_410,N_223);
or U890 (N_890,N_507,N_546);
nand U891 (N_891,N_237,N_550);
or U892 (N_892,N_98,N_461);
xor U893 (N_893,N_199,N_451);
or U894 (N_894,N_2,N_366);
or U895 (N_895,N_61,N_130);
nand U896 (N_896,N_348,N_72);
and U897 (N_897,N_496,N_29);
nor U898 (N_898,N_39,N_122);
or U899 (N_899,N_123,N_329);
nor U900 (N_900,N_408,N_218);
nor U901 (N_901,N_492,N_213);
nand U902 (N_902,N_239,N_33);
nand U903 (N_903,N_429,N_449);
nand U904 (N_904,N_11,N_424);
nor U905 (N_905,N_571,N_47);
and U906 (N_906,N_389,N_89);
or U907 (N_907,N_387,N_13);
or U908 (N_908,N_490,N_282);
nor U909 (N_909,N_199,N_374);
or U910 (N_910,N_187,N_398);
and U911 (N_911,N_258,N_508);
or U912 (N_912,N_21,N_400);
nand U913 (N_913,N_81,N_395);
or U914 (N_914,N_485,N_572);
nand U915 (N_915,N_543,N_589);
and U916 (N_916,N_462,N_502);
nor U917 (N_917,N_341,N_182);
and U918 (N_918,N_540,N_353);
and U919 (N_919,N_415,N_382);
or U920 (N_920,N_555,N_401);
nand U921 (N_921,N_312,N_132);
nor U922 (N_922,N_491,N_361);
and U923 (N_923,N_163,N_121);
or U924 (N_924,N_484,N_116);
and U925 (N_925,N_117,N_173);
nor U926 (N_926,N_66,N_331);
nand U927 (N_927,N_7,N_14);
or U928 (N_928,N_484,N_270);
or U929 (N_929,N_575,N_258);
and U930 (N_930,N_191,N_477);
or U931 (N_931,N_272,N_362);
nand U932 (N_932,N_433,N_471);
xor U933 (N_933,N_544,N_358);
or U934 (N_934,N_247,N_551);
nand U935 (N_935,N_143,N_589);
nand U936 (N_936,N_19,N_299);
and U937 (N_937,N_109,N_141);
and U938 (N_938,N_579,N_10);
nand U939 (N_939,N_542,N_474);
and U940 (N_940,N_525,N_32);
and U941 (N_941,N_587,N_238);
nor U942 (N_942,N_46,N_357);
nand U943 (N_943,N_397,N_193);
nand U944 (N_944,N_254,N_492);
and U945 (N_945,N_201,N_362);
nand U946 (N_946,N_155,N_385);
and U947 (N_947,N_322,N_39);
nand U948 (N_948,N_120,N_538);
nor U949 (N_949,N_166,N_497);
or U950 (N_950,N_459,N_543);
xor U951 (N_951,N_332,N_95);
or U952 (N_952,N_209,N_129);
or U953 (N_953,N_175,N_36);
nand U954 (N_954,N_488,N_135);
and U955 (N_955,N_154,N_562);
or U956 (N_956,N_456,N_399);
or U957 (N_957,N_88,N_404);
nor U958 (N_958,N_108,N_44);
or U959 (N_959,N_418,N_339);
or U960 (N_960,N_524,N_3);
nand U961 (N_961,N_99,N_487);
and U962 (N_962,N_113,N_162);
nand U963 (N_963,N_366,N_518);
or U964 (N_964,N_145,N_523);
nor U965 (N_965,N_260,N_71);
and U966 (N_966,N_396,N_184);
or U967 (N_967,N_341,N_90);
nand U968 (N_968,N_165,N_75);
nor U969 (N_969,N_587,N_250);
nor U970 (N_970,N_512,N_143);
and U971 (N_971,N_242,N_247);
nor U972 (N_972,N_163,N_226);
or U973 (N_973,N_397,N_552);
nand U974 (N_974,N_448,N_218);
nor U975 (N_975,N_431,N_92);
nand U976 (N_976,N_15,N_340);
nand U977 (N_977,N_118,N_204);
nor U978 (N_978,N_74,N_85);
nor U979 (N_979,N_520,N_433);
or U980 (N_980,N_226,N_318);
or U981 (N_981,N_239,N_278);
nor U982 (N_982,N_131,N_191);
and U983 (N_983,N_391,N_49);
or U984 (N_984,N_320,N_10);
nor U985 (N_985,N_460,N_509);
nor U986 (N_986,N_415,N_547);
nand U987 (N_987,N_226,N_512);
nor U988 (N_988,N_506,N_88);
nand U989 (N_989,N_472,N_287);
nand U990 (N_990,N_35,N_230);
or U991 (N_991,N_3,N_91);
or U992 (N_992,N_237,N_474);
nand U993 (N_993,N_50,N_372);
nand U994 (N_994,N_350,N_355);
or U995 (N_995,N_118,N_0);
nor U996 (N_996,N_353,N_370);
nand U997 (N_997,N_171,N_359);
nor U998 (N_998,N_310,N_519);
xor U999 (N_999,N_173,N_412);
nand U1000 (N_1000,N_25,N_350);
or U1001 (N_1001,N_96,N_421);
nand U1002 (N_1002,N_462,N_465);
or U1003 (N_1003,N_117,N_496);
xnor U1004 (N_1004,N_263,N_145);
nor U1005 (N_1005,N_548,N_352);
and U1006 (N_1006,N_336,N_598);
nor U1007 (N_1007,N_148,N_88);
or U1008 (N_1008,N_428,N_593);
nor U1009 (N_1009,N_594,N_459);
nor U1010 (N_1010,N_345,N_294);
or U1011 (N_1011,N_108,N_94);
and U1012 (N_1012,N_228,N_159);
nor U1013 (N_1013,N_237,N_337);
and U1014 (N_1014,N_374,N_203);
and U1015 (N_1015,N_178,N_372);
nor U1016 (N_1016,N_268,N_427);
or U1017 (N_1017,N_87,N_273);
and U1018 (N_1018,N_91,N_341);
nor U1019 (N_1019,N_580,N_284);
and U1020 (N_1020,N_325,N_476);
nand U1021 (N_1021,N_277,N_31);
or U1022 (N_1022,N_442,N_565);
nor U1023 (N_1023,N_256,N_208);
nand U1024 (N_1024,N_360,N_222);
xor U1025 (N_1025,N_157,N_236);
or U1026 (N_1026,N_140,N_341);
or U1027 (N_1027,N_184,N_73);
or U1028 (N_1028,N_148,N_313);
nor U1029 (N_1029,N_167,N_439);
and U1030 (N_1030,N_583,N_4);
nor U1031 (N_1031,N_314,N_545);
nand U1032 (N_1032,N_285,N_298);
or U1033 (N_1033,N_590,N_459);
nor U1034 (N_1034,N_238,N_339);
nor U1035 (N_1035,N_179,N_466);
or U1036 (N_1036,N_288,N_232);
and U1037 (N_1037,N_595,N_538);
nor U1038 (N_1038,N_95,N_447);
xnor U1039 (N_1039,N_468,N_595);
nor U1040 (N_1040,N_159,N_507);
or U1041 (N_1041,N_183,N_105);
and U1042 (N_1042,N_357,N_289);
nor U1043 (N_1043,N_90,N_268);
or U1044 (N_1044,N_248,N_167);
nor U1045 (N_1045,N_532,N_188);
nand U1046 (N_1046,N_107,N_199);
or U1047 (N_1047,N_333,N_472);
nor U1048 (N_1048,N_261,N_298);
and U1049 (N_1049,N_113,N_509);
and U1050 (N_1050,N_253,N_586);
nor U1051 (N_1051,N_388,N_33);
or U1052 (N_1052,N_229,N_274);
or U1053 (N_1053,N_133,N_279);
and U1054 (N_1054,N_67,N_182);
nor U1055 (N_1055,N_215,N_307);
and U1056 (N_1056,N_584,N_529);
or U1057 (N_1057,N_158,N_425);
or U1058 (N_1058,N_57,N_422);
and U1059 (N_1059,N_294,N_226);
and U1060 (N_1060,N_85,N_475);
and U1061 (N_1061,N_101,N_127);
or U1062 (N_1062,N_367,N_572);
and U1063 (N_1063,N_421,N_558);
or U1064 (N_1064,N_36,N_216);
nand U1065 (N_1065,N_191,N_454);
nand U1066 (N_1066,N_551,N_356);
and U1067 (N_1067,N_347,N_277);
or U1068 (N_1068,N_504,N_450);
nor U1069 (N_1069,N_283,N_135);
and U1070 (N_1070,N_446,N_476);
or U1071 (N_1071,N_535,N_221);
and U1072 (N_1072,N_519,N_349);
nand U1073 (N_1073,N_410,N_319);
or U1074 (N_1074,N_583,N_480);
nor U1075 (N_1075,N_510,N_401);
nand U1076 (N_1076,N_480,N_25);
nand U1077 (N_1077,N_539,N_423);
and U1078 (N_1078,N_2,N_25);
and U1079 (N_1079,N_270,N_466);
or U1080 (N_1080,N_105,N_25);
and U1081 (N_1081,N_341,N_561);
nor U1082 (N_1082,N_19,N_97);
nand U1083 (N_1083,N_17,N_83);
nor U1084 (N_1084,N_100,N_477);
nor U1085 (N_1085,N_440,N_34);
nand U1086 (N_1086,N_158,N_202);
or U1087 (N_1087,N_259,N_53);
nor U1088 (N_1088,N_295,N_471);
and U1089 (N_1089,N_589,N_276);
or U1090 (N_1090,N_115,N_479);
nor U1091 (N_1091,N_60,N_85);
or U1092 (N_1092,N_124,N_496);
nor U1093 (N_1093,N_230,N_398);
and U1094 (N_1094,N_500,N_352);
nor U1095 (N_1095,N_219,N_348);
nor U1096 (N_1096,N_574,N_595);
nor U1097 (N_1097,N_490,N_427);
nand U1098 (N_1098,N_32,N_26);
or U1099 (N_1099,N_16,N_149);
nor U1100 (N_1100,N_570,N_15);
and U1101 (N_1101,N_327,N_54);
xor U1102 (N_1102,N_441,N_145);
or U1103 (N_1103,N_553,N_494);
nand U1104 (N_1104,N_553,N_318);
nor U1105 (N_1105,N_258,N_163);
nor U1106 (N_1106,N_181,N_155);
and U1107 (N_1107,N_578,N_160);
nand U1108 (N_1108,N_60,N_258);
nor U1109 (N_1109,N_298,N_202);
nand U1110 (N_1110,N_489,N_112);
nand U1111 (N_1111,N_396,N_412);
nand U1112 (N_1112,N_78,N_469);
or U1113 (N_1113,N_132,N_387);
and U1114 (N_1114,N_463,N_552);
nor U1115 (N_1115,N_191,N_347);
nand U1116 (N_1116,N_91,N_526);
and U1117 (N_1117,N_382,N_114);
nor U1118 (N_1118,N_22,N_458);
and U1119 (N_1119,N_136,N_351);
and U1120 (N_1120,N_399,N_468);
nand U1121 (N_1121,N_92,N_263);
nor U1122 (N_1122,N_326,N_488);
or U1123 (N_1123,N_95,N_587);
nand U1124 (N_1124,N_367,N_301);
and U1125 (N_1125,N_502,N_316);
and U1126 (N_1126,N_349,N_414);
nand U1127 (N_1127,N_69,N_594);
and U1128 (N_1128,N_363,N_130);
nand U1129 (N_1129,N_268,N_483);
or U1130 (N_1130,N_539,N_363);
and U1131 (N_1131,N_174,N_562);
nor U1132 (N_1132,N_425,N_417);
nor U1133 (N_1133,N_361,N_210);
and U1134 (N_1134,N_30,N_185);
and U1135 (N_1135,N_165,N_101);
or U1136 (N_1136,N_345,N_518);
nand U1137 (N_1137,N_269,N_381);
nand U1138 (N_1138,N_208,N_118);
and U1139 (N_1139,N_535,N_162);
nor U1140 (N_1140,N_80,N_586);
and U1141 (N_1141,N_16,N_440);
nand U1142 (N_1142,N_63,N_339);
and U1143 (N_1143,N_484,N_466);
nand U1144 (N_1144,N_492,N_353);
nor U1145 (N_1145,N_468,N_243);
nor U1146 (N_1146,N_570,N_165);
and U1147 (N_1147,N_189,N_142);
nor U1148 (N_1148,N_453,N_110);
nor U1149 (N_1149,N_100,N_522);
nand U1150 (N_1150,N_82,N_156);
or U1151 (N_1151,N_581,N_138);
nor U1152 (N_1152,N_561,N_113);
nor U1153 (N_1153,N_463,N_580);
nand U1154 (N_1154,N_569,N_403);
nor U1155 (N_1155,N_403,N_490);
or U1156 (N_1156,N_479,N_221);
and U1157 (N_1157,N_239,N_465);
or U1158 (N_1158,N_376,N_366);
or U1159 (N_1159,N_283,N_516);
nor U1160 (N_1160,N_394,N_180);
nand U1161 (N_1161,N_574,N_553);
nor U1162 (N_1162,N_406,N_370);
nor U1163 (N_1163,N_69,N_437);
nor U1164 (N_1164,N_207,N_209);
nor U1165 (N_1165,N_451,N_214);
nor U1166 (N_1166,N_33,N_26);
or U1167 (N_1167,N_593,N_379);
or U1168 (N_1168,N_31,N_456);
and U1169 (N_1169,N_369,N_584);
and U1170 (N_1170,N_160,N_72);
or U1171 (N_1171,N_97,N_486);
or U1172 (N_1172,N_304,N_152);
or U1173 (N_1173,N_197,N_453);
nor U1174 (N_1174,N_479,N_259);
or U1175 (N_1175,N_350,N_578);
or U1176 (N_1176,N_394,N_343);
and U1177 (N_1177,N_203,N_396);
nand U1178 (N_1178,N_446,N_77);
nand U1179 (N_1179,N_243,N_550);
and U1180 (N_1180,N_417,N_457);
or U1181 (N_1181,N_256,N_459);
or U1182 (N_1182,N_544,N_94);
nor U1183 (N_1183,N_540,N_590);
nor U1184 (N_1184,N_244,N_532);
and U1185 (N_1185,N_186,N_256);
xnor U1186 (N_1186,N_427,N_247);
nor U1187 (N_1187,N_345,N_398);
nand U1188 (N_1188,N_587,N_220);
nand U1189 (N_1189,N_571,N_0);
nor U1190 (N_1190,N_82,N_228);
nand U1191 (N_1191,N_89,N_353);
and U1192 (N_1192,N_440,N_55);
nand U1193 (N_1193,N_295,N_364);
nand U1194 (N_1194,N_289,N_287);
or U1195 (N_1195,N_586,N_461);
nor U1196 (N_1196,N_343,N_400);
or U1197 (N_1197,N_249,N_16);
or U1198 (N_1198,N_407,N_397);
nand U1199 (N_1199,N_96,N_30);
nor U1200 (N_1200,N_639,N_660);
nor U1201 (N_1201,N_993,N_1127);
and U1202 (N_1202,N_805,N_792);
nand U1203 (N_1203,N_955,N_1064);
and U1204 (N_1204,N_623,N_657);
or U1205 (N_1205,N_1063,N_771);
and U1206 (N_1206,N_969,N_1144);
nor U1207 (N_1207,N_645,N_895);
or U1208 (N_1208,N_612,N_1056);
or U1209 (N_1209,N_829,N_712);
and U1210 (N_1210,N_1014,N_756);
nor U1211 (N_1211,N_948,N_661);
or U1212 (N_1212,N_919,N_750);
nor U1213 (N_1213,N_617,N_637);
xor U1214 (N_1214,N_619,N_605);
and U1215 (N_1215,N_974,N_733);
and U1216 (N_1216,N_673,N_706);
nand U1217 (N_1217,N_1050,N_1005);
and U1218 (N_1218,N_1112,N_1080);
nand U1219 (N_1219,N_921,N_959);
nor U1220 (N_1220,N_1052,N_1084);
nor U1221 (N_1221,N_988,N_853);
and U1222 (N_1222,N_855,N_694);
or U1223 (N_1223,N_910,N_920);
nand U1224 (N_1224,N_862,N_985);
nor U1225 (N_1225,N_1198,N_871);
and U1226 (N_1226,N_972,N_1015);
or U1227 (N_1227,N_837,N_976);
nor U1228 (N_1228,N_1114,N_834);
and U1229 (N_1229,N_1185,N_603);
nor U1230 (N_1230,N_863,N_616);
and U1231 (N_1231,N_1115,N_1013);
nand U1232 (N_1232,N_833,N_997);
nor U1233 (N_1233,N_1044,N_849);
or U1234 (N_1234,N_1136,N_752);
nor U1235 (N_1235,N_982,N_609);
nand U1236 (N_1236,N_755,N_980);
nand U1237 (N_1237,N_1116,N_1178);
nor U1238 (N_1238,N_981,N_906);
or U1239 (N_1239,N_839,N_786);
and U1240 (N_1240,N_765,N_1138);
nor U1241 (N_1241,N_634,N_717);
nor U1242 (N_1242,N_685,N_898);
nand U1243 (N_1243,N_1017,N_888);
nand U1244 (N_1244,N_736,N_1069);
or U1245 (N_1245,N_907,N_827);
nor U1246 (N_1246,N_1078,N_700);
nand U1247 (N_1247,N_817,N_1159);
or U1248 (N_1248,N_1156,N_667);
nand U1249 (N_1249,N_662,N_622);
and U1250 (N_1250,N_901,N_1197);
or U1251 (N_1251,N_949,N_613);
nand U1252 (N_1252,N_913,N_606);
nor U1253 (N_1253,N_838,N_684);
or U1254 (N_1254,N_758,N_822);
or U1255 (N_1255,N_824,N_608);
and U1256 (N_1256,N_818,N_904);
and U1257 (N_1257,N_869,N_950);
or U1258 (N_1258,N_665,N_848);
and U1259 (N_1259,N_958,N_704);
nor U1260 (N_1260,N_1167,N_820);
nor U1261 (N_1261,N_1007,N_866);
or U1262 (N_1262,N_723,N_946);
and U1263 (N_1263,N_790,N_604);
and U1264 (N_1264,N_938,N_1149);
and U1265 (N_1265,N_708,N_716);
or U1266 (N_1266,N_832,N_1032);
xor U1267 (N_1267,N_1142,N_808);
nor U1268 (N_1268,N_1026,N_851);
and U1269 (N_1269,N_923,N_928);
nor U1270 (N_1270,N_1033,N_627);
nor U1271 (N_1271,N_696,N_1035);
or U1272 (N_1272,N_914,N_726);
nand U1273 (N_1273,N_1061,N_638);
and U1274 (N_1274,N_998,N_940);
nor U1275 (N_1275,N_1164,N_648);
or U1276 (N_1276,N_1155,N_762);
xor U1277 (N_1277,N_702,N_902);
xnor U1278 (N_1278,N_654,N_669);
nor U1279 (N_1279,N_675,N_715);
nand U1280 (N_1280,N_1172,N_753);
or U1281 (N_1281,N_867,N_641);
nand U1282 (N_1282,N_737,N_1089);
or U1283 (N_1283,N_1047,N_1106);
nand U1284 (N_1284,N_957,N_1153);
nor U1285 (N_1285,N_680,N_1057);
and U1286 (N_1286,N_1092,N_990);
or U1287 (N_1287,N_699,N_1062);
nand U1288 (N_1288,N_878,N_916);
and U1289 (N_1289,N_766,N_1169);
or U1290 (N_1290,N_1188,N_1070);
nand U1291 (N_1291,N_1096,N_975);
and U1292 (N_1292,N_759,N_741);
or U1293 (N_1293,N_1000,N_924);
nand U1294 (N_1294,N_877,N_693);
nor U1295 (N_1295,N_614,N_894);
or U1296 (N_1296,N_1028,N_1125);
and U1297 (N_1297,N_814,N_740);
nor U1298 (N_1298,N_668,N_1081);
and U1299 (N_1299,N_1150,N_971);
nor U1300 (N_1300,N_1093,N_1135);
nand U1301 (N_1301,N_744,N_767);
or U1302 (N_1302,N_764,N_1141);
or U1303 (N_1303,N_688,N_1002);
and U1304 (N_1304,N_937,N_810);
and U1305 (N_1305,N_1123,N_844);
or U1306 (N_1306,N_1059,N_1184);
or U1307 (N_1307,N_621,N_807);
and U1308 (N_1308,N_886,N_772);
nor U1309 (N_1309,N_1037,N_754);
xor U1310 (N_1310,N_679,N_966);
nand U1311 (N_1311,N_881,N_670);
nand U1312 (N_1312,N_942,N_615);
nand U1313 (N_1313,N_773,N_1139);
nor U1314 (N_1314,N_655,N_811);
or U1315 (N_1315,N_1065,N_780);
nor U1316 (N_1316,N_835,N_856);
and U1317 (N_1317,N_840,N_1042);
nand U1318 (N_1318,N_678,N_801);
nand U1319 (N_1319,N_989,N_676);
or U1320 (N_1320,N_804,N_1170);
or U1321 (N_1321,N_796,N_782);
nand U1322 (N_1322,N_1071,N_1046);
and U1323 (N_1323,N_951,N_784);
or U1324 (N_1324,N_944,N_891);
or U1325 (N_1325,N_647,N_1049);
or U1326 (N_1326,N_698,N_1019);
nand U1327 (N_1327,N_987,N_903);
and U1328 (N_1328,N_1102,N_1024);
and U1329 (N_1329,N_1104,N_1072);
or U1330 (N_1330,N_1129,N_831);
and U1331 (N_1331,N_941,N_896);
nor U1332 (N_1332,N_864,N_787);
nand U1333 (N_1333,N_683,N_1189);
or U1334 (N_1334,N_802,N_611);
or U1335 (N_1335,N_632,N_1025);
nor U1336 (N_1336,N_1098,N_671);
nand U1337 (N_1337,N_1161,N_776);
or U1338 (N_1338,N_986,N_794);
and U1339 (N_1339,N_1016,N_882);
or U1340 (N_1340,N_961,N_873);
nor U1341 (N_1341,N_1103,N_663);
nor U1342 (N_1342,N_1168,N_1173);
or U1343 (N_1343,N_610,N_1105);
and U1344 (N_1344,N_964,N_666);
xor U1345 (N_1345,N_1030,N_859);
nand U1346 (N_1346,N_936,N_664);
and U1347 (N_1347,N_713,N_943);
nand U1348 (N_1348,N_727,N_629);
and U1349 (N_1349,N_636,N_1039);
or U1350 (N_1350,N_1043,N_746);
and U1351 (N_1351,N_734,N_1182);
or U1352 (N_1352,N_749,N_1094);
nor U1353 (N_1353,N_813,N_779);
nor U1354 (N_1354,N_1001,N_1154);
nand U1355 (N_1355,N_977,N_995);
nand U1356 (N_1356,N_729,N_631);
nand U1357 (N_1357,N_1036,N_659);
nand U1358 (N_1358,N_1038,N_799);
nand U1359 (N_1359,N_884,N_825);
and U1360 (N_1360,N_843,N_875);
or U1361 (N_1361,N_652,N_887);
nand U1362 (N_1362,N_893,N_651);
nand U1363 (N_1363,N_761,N_798);
nand U1364 (N_1364,N_1066,N_774);
or U1365 (N_1365,N_695,N_1137);
nor U1366 (N_1366,N_646,N_1088);
nand U1367 (N_1367,N_900,N_1012);
or U1368 (N_1368,N_751,N_994);
and U1369 (N_1369,N_653,N_1055);
nand U1370 (N_1370,N_821,N_1180);
nor U1371 (N_1371,N_1192,N_1160);
and U1372 (N_1372,N_1120,N_1126);
and U1373 (N_1373,N_640,N_747);
or U1374 (N_1374,N_710,N_601);
nor U1375 (N_1375,N_991,N_1195);
nor U1376 (N_1376,N_812,N_912);
nor U1377 (N_1377,N_1048,N_933);
or U1378 (N_1378,N_770,N_860);
nor U1379 (N_1379,N_1087,N_1091);
nand U1380 (N_1380,N_635,N_760);
and U1381 (N_1381,N_963,N_1113);
or U1382 (N_1382,N_979,N_1045);
or U1383 (N_1383,N_1109,N_777);
nand U1384 (N_1384,N_1101,N_1111);
nor U1385 (N_1385,N_939,N_890);
xnor U1386 (N_1386,N_642,N_1076);
nor U1387 (N_1387,N_999,N_1067);
xor U1388 (N_1388,N_707,N_687);
or U1389 (N_1389,N_1040,N_728);
or U1390 (N_1390,N_1027,N_1132);
nand U1391 (N_1391,N_624,N_1090);
nand U1392 (N_1392,N_677,N_865);
nand U1393 (N_1393,N_806,N_1199);
nor U1394 (N_1394,N_1128,N_845);
and U1395 (N_1395,N_1110,N_960);
or U1396 (N_1396,N_1118,N_1086);
nand U1397 (N_1397,N_952,N_690);
nor U1398 (N_1398,N_650,N_809);
or U1399 (N_1399,N_725,N_1022);
or U1400 (N_1400,N_953,N_795);
and U1401 (N_1401,N_649,N_1171);
or U1402 (N_1402,N_1006,N_1157);
nand U1403 (N_1403,N_816,N_1020);
nor U1404 (N_1404,N_1163,N_956);
nor U1405 (N_1405,N_918,N_872);
nor U1406 (N_1406,N_1133,N_1108);
nand U1407 (N_1407,N_984,N_1152);
and U1408 (N_1408,N_722,N_730);
or U1409 (N_1409,N_954,N_745);
nor U1410 (N_1410,N_1121,N_742);
or U1411 (N_1411,N_803,N_630);
and U1412 (N_1412,N_797,N_861);
or U1413 (N_1413,N_842,N_757);
nor U1414 (N_1414,N_858,N_768);
and U1415 (N_1415,N_1176,N_826);
nand U1416 (N_1416,N_1100,N_932);
and U1417 (N_1417,N_735,N_996);
nand U1418 (N_1418,N_701,N_644);
or U1419 (N_1419,N_1148,N_1179);
nand U1420 (N_1420,N_883,N_1145);
and U1421 (N_1421,N_1124,N_846);
xor U1422 (N_1422,N_970,N_1162);
nand U1423 (N_1423,N_1190,N_1021);
nand U1424 (N_1424,N_709,N_743);
nor U1425 (N_1425,N_879,N_785);
nor U1426 (N_1426,N_705,N_602);
or U1427 (N_1427,N_689,N_1165);
or U1428 (N_1428,N_1083,N_1134);
and U1429 (N_1429,N_909,N_721);
nor U1430 (N_1430,N_1095,N_800);
or U1431 (N_1431,N_1082,N_607);
or U1432 (N_1432,N_691,N_791);
nor U1433 (N_1433,N_1003,N_819);
or U1434 (N_1434,N_1077,N_1107);
or U1435 (N_1435,N_908,N_686);
nor U1436 (N_1436,N_917,N_1031);
or U1437 (N_1437,N_847,N_1151);
nor U1438 (N_1438,N_935,N_1122);
and U1439 (N_1439,N_793,N_915);
and U1440 (N_1440,N_656,N_625);
and U1441 (N_1441,N_714,N_841);
or U1442 (N_1442,N_892,N_769);
or U1443 (N_1443,N_748,N_1060);
nor U1444 (N_1444,N_718,N_965);
or U1445 (N_1445,N_719,N_967);
or U1446 (N_1446,N_732,N_1143);
or U1447 (N_1447,N_618,N_781);
xnor U1448 (N_1448,N_854,N_1079);
nor U1449 (N_1449,N_1193,N_1174);
or U1450 (N_1450,N_931,N_724);
and U1451 (N_1451,N_947,N_1004);
nand U1452 (N_1452,N_643,N_1187);
or U1453 (N_1453,N_1181,N_992);
nor U1454 (N_1454,N_899,N_905);
or U1455 (N_1455,N_885,N_731);
and U1456 (N_1456,N_1009,N_697);
nand U1457 (N_1457,N_1097,N_600);
nand U1458 (N_1458,N_850,N_1085);
or U1459 (N_1459,N_911,N_1183);
and U1460 (N_1460,N_1158,N_628);
xnor U1461 (N_1461,N_1146,N_1177);
or U1462 (N_1462,N_828,N_1099);
or U1463 (N_1463,N_620,N_763);
nor U1464 (N_1464,N_1175,N_775);
nor U1465 (N_1465,N_672,N_778);
or U1466 (N_1466,N_874,N_789);
nor U1467 (N_1467,N_1053,N_868);
xor U1468 (N_1468,N_880,N_1018);
xor U1469 (N_1469,N_1194,N_1051);
nand U1470 (N_1470,N_739,N_692);
and U1471 (N_1471,N_983,N_852);
nand U1472 (N_1472,N_1140,N_783);
and U1473 (N_1473,N_1131,N_927);
nor U1474 (N_1474,N_897,N_930);
or U1475 (N_1475,N_925,N_681);
nand U1476 (N_1476,N_711,N_836);
nand U1477 (N_1477,N_674,N_1034);
nand U1478 (N_1478,N_1075,N_658);
and U1479 (N_1479,N_870,N_1058);
nor U1480 (N_1480,N_1166,N_1029);
nor U1481 (N_1481,N_823,N_934);
and U1482 (N_1482,N_1041,N_626);
xnor U1483 (N_1483,N_720,N_876);
or U1484 (N_1484,N_1147,N_1119);
nand U1485 (N_1485,N_973,N_633);
nor U1486 (N_1486,N_978,N_889);
nor U1487 (N_1487,N_1191,N_788);
nand U1488 (N_1488,N_962,N_857);
or U1489 (N_1489,N_1073,N_1008);
nor U1490 (N_1490,N_1011,N_815);
or U1491 (N_1491,N_1130,N_1186);
and U1492 (N_1492,N_1054,N_968);
nand U1493 (N_1493,N_1074,N_1196);
nor U1494 (N_1494,N_703,N_1117);
nand U1495 (N_1495,N_738,N_926);
or U1496 (N_1496,N_1023,N_929);
nor U1497 (N_1497,N_922,N_830);
or U1498 (N_1498,N_1010,N_945);
or U1499 (N_1499,N_1068,N_682);
and U1500 (N_1500,N_613,N_1132);
nor U1501 (N_1501,N_1120,N_1129);
nor U1502 (N_1502,N_1131,N_921);
nor U1503 (N_1503,N_988,N_627);
nand U1504 (N_1504,N_777,N_996);
nor U1505 (N_1505,N_1034,N_635);
nor U1506 (N_1506,N_870,N_1005);
nand U1507 (N_1507,N_999,N_1121);
or U1508 (N_1508,N_790,N_674);
and U1509 (N_1509,N_771,N_621);
and U1510 (N_1510,N_1096,N_1014);
nor U1511 (N_1511,N_1110,N_682);
nand U1512 (N_1512,N_957,N_667);
nand U1513 (N_1513,N_944,N_1093);
nor U1514 (N_1514,N_806,N_670);
or U1515 (N_1515,N_631,N_774);
and U1516 (N_1516,N_1122,N_939);
nand U1517 (N_1517,N_852,N_904);
and U1518 (N_1518,N_713,N_1047);
nor U1519 (N_1519,N_837,N_1145);
nand U1520 (N_1520,N_710,N_662);
and U1521 (N_1521,N_1007,N_1063);
and U1522 (N_1522,N_623,N_718);
xnor U1523 (N_1523,N_826,N_749);
nand U1524 (N_1524,N_740,N_701);
nor U1525 (N_1525,N_876,N_824);
or U1526 (N_1526,N_1049,N_1176);
nand U1527 (N_1527,N_933,N_765);
nand U1528 (N_1528,N_924,N_750);
and U1529 (N_1529,N_622,N_858);
or U1530 (N_1530,N_817,N_727);
nand U1531 (N_1531,N_889,N_748);
or U1532 (N_1532,N_765,N_645);
or U1533 (N_1533,N_860,N_882);
nor U1534 (N_1534,N_1104,N_758);
nand U1535 (N_1535,N_692,N_1048);
and U1536 (N_1536,N_811,N_1058);
or U1537 (N_1537,N_1098,N_1048);
and U1538 (N_1538,N_854,N_805);
and U1539 (N_1539,N_1146,N_1080);
nand U1540 (N_1540,N_936,N_925);
and U1541 (N_1541,N_824,N_980);
or U1542 (N_1542,N_711,N_905);
or U1543 (N_1543,N_844,N_921);
nand U1544 (N_1544,N_1097,N_677);
nor U1545 (N_1545,N_1182,N_980);
or U1546 (N_1546,N_817,N_759);
or U1547 (N_1547,N_886,N_968);
or U1548 (N_1548,N_879,N_941);
and U1549 (N_1549,N_1145,N_795);
nor U1550 (N_1550,N_611,N_956);
nor U1551 (N_1551,N_972,N_789);
nand U1552 (N_1552,N_983,N_807);
nand U1553 (N_1553,N_793,N_816);
nor U1554 (N_1554,N_1193,N_1000);
or U1555 (N_1555,N_999,N_939);
or U1556 (N_1556,N_1169,N_1139);
or U1557 (N_1557,N_918,N_909);
xor U1558 (N_1558,N_990,N_901);
and U1559 (N_1559,N_1176,N_1004);
nand U1560 (N_1560,N_1128,N_1075);
nand U1561 (N_1561,N_1157,N_635);
and U1562 (N_1562,N_1168,N_602);
and U1563 (N_1563,N_1142,N_913);
and U1564 (N_1564,N_663,N_1021);
or U1565 (N_1565,N_821,N_1000);
or U1566 (N_1566,N_1138,N_878);
and U1567 (N_1567,N_728,N_1043);
nor U1568 (N_1568,N_807,N_914);
nand U1569 (N_1569,N_968,N_802);
nand U1570 (N_1570,N_888,N_1074);
and U1571 (N_1571,N_965,N_630);
nor U1572 (N_1572,N_634,N_689);
nor U1573 (N_1573,N_653,N_835);
nor U1574 (N_1574,N_764,N_1153);
nor U1575 (N_1575,N_812,N_946);
and U1576 (N_1576,N_984,N_899);
nand U1577 (N_1577,N_854,N_681);
nand U1578 (N_1578,N_1041,N_1148);
nor U1579 (N_1579,N_1001,N_876);
and U1580 (N_1580,N_750,N_926);
nor U1581 (N_1581,N_1073,N_717);
nor U1582 (N_1582,N_781,N_1045);
or U1583 (N_1583,N_951,N_707);
nand U1584 (N_1584,N_619,N_832);
nor U1585 (N_1585,N_974,N_654);
or U1586 (N_1586,N_1134,N_1064);
or U1587 (N_1587,N_756,N_687);
nor U1588 (N_1588,N_777,N_631);
and U1589 (N_1589,N_930,N_1161);
or U1590 (N_1590,N_675,N_712);
or U1591 (N_1591,N_1067,N_1005);
xnor U1592 (N_1592,N_1168,N_708);
nor U1593 (N_1593,N_605,N_886);
or U1594 (N_1594,N_1136,N_652);
or U1595 (N_1595,N_669,N_750);
and U1596 (N_1596,N_1199,N_875);
nand U1597 (N_1597,N_690,N_1135);
or U1598 (N_1598,N_1099,N_1145);
or U1599 (N_1599,N_1178,N_711);
nor U1600 (N_1600,N_733,N_998);
and U1601 (N_1601,N_1061,N_1004);
nand U1602 (N_1602,N_1140,N_749);
and U1603 (N_1603,N_648,N_1017);
nor U1604 (N_1604,N_1015,N_870);
or U1605 (N_1605,N_726,N_670);
or U1606 (N_1606,N_1135,N_1126);
or U1607 (N_1607,N_849,N_799);
and U1608 (N_1608,N_628,N_654);
nand U1609 (N_1609,N_602,N_669);
nand U1610 (N_1610,N_955,N_796);
or U1611 (N_1611,N_938,N_622);
nand U1612 (N_1612,N_678,N_611);
nand U1613 (N_1613,N_866,N_1183);
and U1614 (N_1614,N_776,N_1033);
and U1615 (N_1615,N_988,N_899);
or U1616 (N_1616,N_914,N_1130);
nand U1617 (N_1617,N_738,N_832);
nor U1618 (N_1618,N_1194,N_663);
nor U1619 (N_1619,N_985,N_1015);
and U1620 (N_1620,N_957,N_1144);
nand U1621 (N_1621,N_1053,N_877);
nor U1622 (N_1622,N_950,N_1011);
and U1623 (N_1623,N_1156,N_787);
or U1624 (N_1624,N_1077,N_855);
nor U1625 (N_1625,N_1030,N_1037);
and U1626 (N_1626,N_671,N_636);
and U1627 (N_1627,N_748,N_1098);
and U1628 (N_1628,N_1186,N_967);
nor U1629 (N_1629,N_1074,N_984);
nand U1630 (N_1630,N_790,N_744);
and U1631 (N_1631,N_1067,N_716);
or U1632 (N_1632,N_910,N_814);
nor U1633 (N_1633,N_919,N_905);
nor U1634 (N_1634,N_1110,N_749);
nor U1635 (N_1635,N_1152,N_1066);
or U1636 (N_1636,N_1184,N_721);
nand U1637 (N_1637,N_940,N_1099);
and U1638 (N_1638,N_1124,N_931);
or U1639 (N_1639,N_1105,N_685);
nand U1640 (N_1640,N_1055,N_710);
nand U1641 (N_1641,N_1154,N_963);
nand U1642 (N_1642,N_1044,N_617);
nand U1643 (N_1643,N_635,N_916);
nand U1644 (N_1644,N_1113,N_716);
and U1645 (N_1645,N_1101,N_1010);
or U1646 (N_1646,N_764,N_1180);
or U1647 (N_1647,N_978,N_1100);
xor U1648 (N_1648,N_1082,N_1174);
and U1649 (N_1649,N_882,N_1161);
nor U1650 (N_1650,N_1132,N_753);
xnor U1651 (N_1651,N_1047,N_771);
and U1652 (N_1652,N_861,N_916);
and U1653 (N_1653,N_935,N_714);
nor U1654 (N_1654,N_1101,N_1102);
nand U1655 (N_1655,N_949,N_790);
or U1656 (N_1656,N_770,N_621);
nand U1657 (N_1657,N_788,N_1131);
or U1658 (N_1658,N_735,N_630);
nor U1659 (N_1659,N_736,N_890);
or U1660 (N_1660,N_850,N_889);
nand U1661 (N_1661,N_608,N_985);
nor U1662 (N_1662,N_995,N_982);
and U1663 (N_1663,N_1059,N_1042);
or U1664 (N_1664,N_730,N_1051);
nor U1665 (N_1665,N_964,N_929);
nand U1666 (N_1666,N_972,N_852);
nand U1667 (N_1667,N_741,N_912);
nand U1668 (N_1668,N_855,N_715);
and U1669 (N_1669,N_1046,N_1074);
or U1670 (N_1670,N_977,N_632);
xnor U1671 (N_1671,N_998,N_678);
nor U1672 (N_1672,N_718,N_847);
nand U1673 (N_1673,N_659,N_754);
nand U1674 (N_1674,N_970,N_1035);
nor U1675 (N_1675,N_1142,N_911);
and U1676 (N_1676,N_840,N_893);
nor U1677 (N_1677,N_787,N_653);
nor U1678 (N_1678,N_866,N_911);
or U1679 (N_1679,N_939,N_1091);
nor U1680 (N_1680,N_1189,N_1188);
nand U1681 (N_1681,N_1034,N_807);
and U1682 (N_1682,N_700,N_807);
nand U1683 (N_1683,N_628,N_656);
or U1684 (N_1684,N_1089,N_888);
nand U1685 (N_1685,N_1027,N_671);
nand U1686 (N_1686,N_784,N_868);
or U1687 (N_1687,N_820,N_1087);
nand U1688 (N_1688,N_842,N_892);
nand U1689 (N_1689,N_1044,N_1193);
or U1690 (N_1690,N_799,N_745);
nand U1691 (N_1691,N_675,N_740);
or U1692 (N_1692,N_1019,N_818);
nand U1693 (N_1693,N_1196,N_1005);
nand U1694 (N_1694,N_714,N_860);
nand U1695 (N_1695,N_1161,N_1184);
and U1696 (N_1696,N_1129,N_1084);
nor U1697 (N_1697,N_900,N_1148);
or U1698 (N_1698,N_949,N_648);
nor U1699 (N_1699,N_1058,N_774);
nor U1700 (N_1700,N_1177,N_683);
or U1701 (N_1701,N_829,N_1192);
xnor U1702 (N_1702,N_898,N_1028);
or U1703 (N_1703,N_817,N_690);
nor U1704 (N_1704,N_615,N_676);
and U1705 (N_1705,N_707,N_791);
nand U1706 (N_1706,N_706,N_759);
nor U1707 (N_1707,N_861,N_887);
nor U1708 (N_1708,N_749,N_1154);
nor U1709 (N_1709,N_995,N_969);
nand U1710 (N_1710,N_973,N_771);
nand U1711 (N_1711,N_704,N_663);
and U1712 (N_1712,N_1169,N_691);
and U1713 (N_1713,N_877,N_870);
nand U1714 (N_1714,N_929,N_996);
nand U1715 (N_1715,N_843,N_697);
and U1716 (N_1716,N_947,N_1059);
and U1717 (N_1717,N_1005,N_839);
nor U1718 (N_1718,N_920,N_1195);
or U1719 (N_1719,N_763,N_668);
nor U1720 (N_1720,N_1009,N_782);
or U1721 (N_1721,N_658,N_961);
or U1722 (N_1722,N_1142,N_1078);
nor U1723 (N_1723,N_985,N_797);
nor U1724 (N_1724,N_1020,N_1098);
and U1725 (N_1725,N_781,N_679);
and U1726 (N_1726,N_867,N_909);
or U1727 (N_1727,N_944,N_894);
or U1728 (N_1728,N_916,N_1129);
and U1729 (N_1729,N_923,N_1066);
or U1730 (N_1730,N_716,N_718);
xor U1731 (N_1731,N_877,N_834);
nor U1732 (N_1732,N_642,N_869);
nand U1733 (N_1733,N_873,N_760);
nor U1734 (N_1734,N_743,N_1043);
and U1735 (N_1735,N_785,N_1170);
nor U1736 (N_1736,N_831,N_1198);
and U1737 (N_1737,N_693,N_794);
and U1738 (N_1738,N_1082,N_1130);
and U1739 (N_1739,N_605,N_1054);
nor U1740 (N_1740,N_999,N_1004);
and U1741 (N_1741,N_979,N_669);
and U1742 (N_1742,N_966,N_840);
nor U1743 (N_1743,N_1031,N_1012);
nand U1744 (N_1744,N_888,N_848);
nand U1745 (N_1745,N_605,N_1045);
and U1746 (N_1746,N_1104,N_799);
or U1747 (N_1747,N_880,N_646);
or U1748 (N_1748,N_1048,N_1190);
nand U1749 (N_1749,N_1114,N_866);
nor U1750 (N_1750,N_703,N_811);
nor U1751 (N_1751,N_1001,N_1037);
and U1752 (N_1752,N_622,N_627);
nor U1753 (N_1753,N_1097,N_998);
and U1754 (N_1754,N_1029,N_672);
or U1755 (N_1755,N_1009,N_634);
and U1756 (N_1756,N_1145,N_728);
and U1757 (N_1757,N_887,N_1108);
nand U1758 (N_1758,N_797,N_1017);
nor U1759 (N_1759,N_985,N_1000);
nand U1760 (N_1760,N_716,N_927);
nand U1761 (N_1761,N_928,N_1044);
or U1762 (N_1762,N_1007,N_1160);
nand U1763 (N_1763,N_955,N_695);
nand U1764 (N_1764,N_1146,N_968);
nand U1765 (N_1765,N_1146,N_1086);
or U1766 (N_1766,N_806,N_677);
nand U1767 (N_1767,N_1114,N_667);
and U1768 (N_1768,N_842,N_656);
and U1769 (N_1769,N_923,N_906);
and U1770 (N_1770,N_801,N_707);
nand U1771 (N_1771,N_808,N_1073);
nand U1772 (N_1772,N_1185,N_896);
nand U1773 (N_1773,N_847,N_933);
nand U1774 (N_1774,N_1082,N_877);
nand U1775 (N_1775,N_710,N_928);
and U1776 (N_1776,N_1168,N_687);
nand U1777 (N_1777,N_1024,N_744);
or U1778 (N_1778,N_1048,N_633);
nor U1779 (N_1779,N_910,N_978);
nand U1780 (N_1780,N_943,N_769);
or U1781 (N_1781,N_623,N_891);
and U1782 (N_1782,N_1191,N_710);
nand U1783 (N_1783,N_764,N_1124);
nand U1784 (N_1784,N_730,N_900);
nand U1785 (N_1785,N_1014,N_1192);
nand U1786 (N_1786,N_1049,N_1090);
nand U1787 (N_1787,N_1138,N_1093);
and U1788 (N_1788,N_732,N_938);
and U1789 (N_1789,N_772,N_786);
nand U1790 (N_1790,N_1155,N_643);
nor U1791 (N_1791,N_764,N_908);
and U1792 (N_1792,N_1043,N_1182);
nand U1793 (N_1793,N_815,N_901);
nand U1794 (N_1794,N_756,N_1151);
nand U1795 (N_1795,N_833,N_753);
or U1796 (N_1796,N_852,N_869);
nor U1797 (N_1797,N_1153,N_1138);
nand U1798 (N_1798,N_843,N_1156);
or U1799 (N_1799,N_1027,N_834);
nand U1800 (N_1800,N_1776,N_1380);
or U1801 (N_1801,N_1688,N_1758);
and U1802 (N_1802,N_1695,N_1791);
nor U1803 (N_1803,N_1505,N_1251);
or U1804 (N_1804,N_1790,N_1767);
nor U1805 (N_1805,N_1488,N_1554);
nor U1806 (N_1806,N_1750,N_1376);
nor U1807 (N_1807,N_1719,N_1303);
nor U1808 (N_1808,N_1589,N_1779);
and U1809 (N_1809,N_1566,N_1243);
nand U1810 (N_1810,N_1782,N_1378);
and U1811 (N_1811,N_1318,N_1305);
or U1812 (N_1812,N_1720,N_1386);
and U1813 (N_1813,N_1761,N_1619);
nor U1814 (N_1814,N_1572,N_1382);
or U1815 (N_1815,N_1694,N_1519);
nor U1816 (N_1816,N_1736,N_1207);
xnor U1817 (N_1817,N_1227,N_1266);
nand U1818 (N_1818,N_1433,N_1471);
nand U1819 (N_1819,N_1490,N_1575);
xnor U1820 (N_1820,N_1706,N_1388);
nor U1821 (N_1821,N_1289,N_1611);
and U1822 (N_1822,N_1581,N_1792);
or U1823 (N_1823,N_1390,N_1651);
nor U1824 (N_1824,N_1320,N_1285);
or U1825 (N_1825,N_1555,N_1712);
or U1826 (N_1826,N_1533,N_1258);
xnor U1827 (N_1827,N_1466,N_1665);
and U1828 (N_1828,N_1395,N_1729);
and U1829 (N_1829,N_1653,N_1584);
and U1830 (N_1830,N_1544,N_1438);
xor U1831 (N_1831,N_1236,N_1536);
or U1832 (N_1832,N_1474,N_1740);
xnor U1833 (N_1833,N_1406,N_1668);
nor U1834 (N_1834,N_1573,N_1279);
nand U1835 (N_1835,N_1673,N_1551);
and U1836 (N_1836,N_1567,N_1629);
nor U1837 (N_1837,N_1309,N_1493);
nand U1838 (N_1838,N_1260,N_1705);
nand U1839 (N_1839,N_1721,N_1447);
nor U1840 (N_1840,N_1642,N_1666);
nor U1841 (N_1841,N_1422,N_1359);
or U1842 (N_1842,N_1543,N_1787);
or U1843 (N_1843,N_1362,N_1387);
and U1844 (N_1844,N_1443,N_1714);
or U1845 (N_1845,N_1646,N_1777);
or U1846 (N_1846,N_1268,N_1654);
nand U1847 (N_1847,N_1252,N_1639);
or U1848 (N_1848,N_1702,N_1560);
nor U1849 (N_1849,N_1739,N_1707);
nor U1850 (N_1850,N_1778,N_1669);
nand U1851 (N_1851,N_1278,N_1757);
and U1852 (N_1852,N_1248,N_1297);
nand U1853 (N_1853,N_1649,N_1261);
or U1854 (N_1854,N_1331,N_1564);
and U1855 (N_1855,N_1340,N_1598);
and U1856 (N_1856,N_1615,N_1231);
nor U1857 (N_1857,N_1553,N_1256);
nand U1858 (N_1858,N_1614,N_1345);
nor U1859 (N_1859,N_1249,N_1346);
and U1860 (N_1860,N_1496,N_1738);
nand U1861 (N_1861,N_1735,N_1431);
nor U1862 (N_1862,N_1693,N_1242);
nor U1863 (N_1863,N_1394,N_1239);
nand U1864 (N_1864,N_1458,N_1637);
and U1865 (N_1865,N_1622,N_1579);
nand U1866 (N_1866,N_1218,N_1525);
nor U1867 (N_1867,N_1741,N_1770);
nor U1868 (N_1868,N_1708,N_1436);
or U1869 (N_1869,N_1607,N_1586);
and U1870 (N_1870,N_1749,N_1238);
nor U1871 (N_1871,N_1700,N_1765);
nor U1872 (N_1872,N_1437,N_1479);
nand U1873 (N_1873,N_1212,N_1407);
or U1874 (N_1874,N_1327,N_1219);
and U1875 (N_1875,N_1494,N_1364);
and U1876 (N_1876,N_1418,N_1492);
or U1877 (N_1877,N_1506,N_1764);
and U1878 (N_1878,N_1670,N_1202);
and U1879 (N_1879,N_1208,N_1635);
nor U1880 (N_1880,N_1780,N_1240);
and U1881 (N_1881,N_1703,N_1455);
nor U1882 (N_1882,N_1414,N_1457);
and U1883 (N_1883,N_1511,N_1689);
nand U1884 (N_1884,N_1491,N_1797);
nor U1885 (N_1885,N_1547,N_1569);
and U1886 (N_1886,N_1587,N_1300);
and U1887 (N_1887,N_1645,N_1323);
and U1888 (N_1888,N_1477,N_1427);
and U1889 (N_1889,N_1284,N_1424);
and U1890 (N_1890,N_1763,N_1756);
nor U1891 (N_1891,N_1214,N_1540);
nand U1892 (N_1892,N_1524,N_1223);
nand U1893 (N_1893,N_1597,N_1384);
nand U1894 (N_1894,N_1601,N_1771);
and U1895 (N_1895,N_1354,N_1552);
nand U1896 (N_1896,N_1253,N_1613);
and U1897 (N_1897,N_1401,N_1393);
nor U1898 (N_1898,N_1324,N_1576);
or U1899 (N_1899,N_1397,N_1798);
or U1900 (N_1900,N_1641,N_1617);
nor U1901 (N_1901,N_1290,N_1697);
and U1902 (N_1902,N_1472,N_1664);
or U1903 (N_1903,N_1448,N_1593);
and U1904 (N_1904,N_1785,N_1557);
and U1905 (N_1905,N_1294,N_1636);
and U1906 (N_1906,N_1531,N_1442);
nand U1907 (N_1907,N_1277,N_1726);
and U1908 (N_1908,N_1267,N_1459);
or U1909 (N_1909,N_1716,N_1475);
nor U1910 (N_1910,N_1209,N_1287);
nand U1911 (N_1911,N_1679,N_1274);
or U1912 (N_1912,N_1516,N_1262);
and U1913 (N_1913,N_1675,N_1781);
or U1914 (N_1914,N_1409,N_1396);
and U1915 (N_1915,N_1226,N_1419);
and U1916 (N_1916,N_1762,N_1451);
or U1917 (N_1917,N_1734,N_1772);
or U1918 (N_1918,N_1361,N_1621);
xor U1919 (N_1919,N_1691,N_1349);
nor U1920 (N_1920,N_1299,N_1728);
xnor U1921 (N_1921,N_1237,N_1213);
nand U1922 (N_1922,N_1201,N_1224);
or U1923 (N_1923,N_1500,N_1434);
nor U1924 (N_1924,N_1467,N_1643);
nand U1925 (N_1925,N_1353,N_1514);
nand U1926 (N_1926,N_1215,N_1273);
and U1927 (N_1927,N_1446,N_1271);
nor U1928 (N_1928,N_1216,N_1341);
or U1929 (N_1929,N_1690,N_1217);
nand U1930 (N_1930,N_1528,N_1561);
and U1931 (N_1931,N_1591,N_1504);
nor U1932 (N_1932,N_1685,N_1461);
or U1933 (N_1933,N_1704,N_1392);
or U1934 (N_1934,N_1462,N_1225);
and U1935 (N_1935,N_1545,N_1711);
nor U1936 (N_1936,N_1338,N_1468);
nand U1937 (N_1937,N_1715,N_1210);
or U1938 (N_1938,N_1339,N_1499);
and U1939 (N_1939,N_1445,N_1541);
and U1940 (N_1940,N_1610,N_1344);
and U1941 (N_1941,N_1680,N_1766);
nor U1942 (N_1942,N_1351,N_1306);
and U1943 (N_1943,N_1751,N_1565);
nor U1944 (N_1944,N_1744,N_1513);
nor U1945 (N_1945,N_1432,N_1683);
or U1946 (N_1946,N_1269,N_1507);
nor U1947 (N_1947,N_1546,N_1599);
or U1948 (N_1948,N_1754,N_1315);
nand U1949 (N_1949,N_1298,N_1530);
nor U1950 (N_1950,N_1234,N_1769);
and U1951 (N_1951,N_1737,N_1257);
xnor U1952 (N_1952,N_1747,N_1347);
or U1953 (N_1953,N_1644,N_1794);
or U1954 (N_1954,N_1568,N_1463);
xor U1955 (N_1955,N_1532,N_1502);
and U1956 (N_1956,N_1399,N_1795);
and U1957 (N_1957,N_1301,N_1510);
nor U1958 (N_1958,N_1423,N_1529);
nand U1959 (N_1959,N_1293,N_1481);
nor U1960 (N_1960,N_1348,N_1337);
nor U1961 (N_1961,N_1460,N_1247);
and U1962 (N_1962,N_1295,N_1408);
nor U1963 (N_1963,N_1632,N_1501);
or U1964 (N_1964,N_1333,N_1508);
nor U1965 (N_1965,N_1383,N_1311);
nand U1966 (N_1966,N_1275,N_1200);
or U1967 (N_1967,N_1430,N_1571);
and U1968 (N_1968,N_1667,N_1411);
nor U1969 (N_1969,N_1313,N_1381);
nor U1970 (N_1970,N_1304,N_1476);
nor U1971 (N_1971,N_1682,N_1420);
nand U1972 (N_1972,N_1701,N_1600);
nor U1973 (N_1973,N_1296,N_1580);
nand U1974 (N_1974,N_1517,N_1788);
and U1975 (N_1975,N_1444,N_1404);
xnor U1976 (N_1976,N_1487,N_1672);
and U1977 (N_1977,N_1206,N_1439);
nor U1978 (N_1978,N_1485,N_1722);
nor U1979 (N_1979,N_1281,N_1730);
nor U1980 (N_1980,N_1308,N_1241);
and U1981 (N_1981,N_1410,N_1570);
nor U1982 (N_1982,N_1698,N_1426);
nand U1983 (N_1983,N_1659,N_1283);
or U1984 (N_1984,N_1233,N_1270);
nor U1985 (N_1985,N_1656,N_1548);
nor U1986 (N_1986,N_1470,N_1374);
or U1987 (N_1987,N_1350,N_1421);
or U1988 (N_1988,N_1360,N_1332);
or U1989 (N_1989,N_1774,N_1522);
nand U1990 (N_1990,N_1366,N_1727);
nor U1991 (N_1991,N_1435,N_1687);
and U1992 (N_1992,N_1538,N_1465);
or U1993 (N_1993,N_1612,N_1692);
and U1994 (N_1994,N_1291,N_1321);
nor U1995 (N_1995,N_1441,N_1638);
or U1996 (N_1996,N_1773,N_1678);
or U1997 (N_1997,N_1539,N_1648);
nor U1998 (N_1998,N_1398,N_1742);
nand U1999 (N_1999,N_1367,N_1498);
nand U2000 (N_2000,N_1369,N_1230);
or U2001 (N_2001,N_1521,N_1732);
nand U2002 (N_2002,N_1489,N_1671);
or U2003 (N_2003,N_1609,N_1640);
and U2004 (N_2004,N_1550,N_1425);
nand U2005 (N_2005,N_1330,N_1631);
and U2006 (N_2006,N_1625,N_1783);
nand U2007 (N_2007,N_1211,N_1583);
nor U2008 (N_2008,N_1677,N_1358);
nor U2009 (N_2009,N_1265,N_1562);
or U2010 (N_2010,N_1245,N_1220);
or U2011 (N_2011,N_1577,N_1630);
nand U2012 (N_2012,N_1731,N_1662);
or U2013 (N_2013,N_1452,N_1464);
and U2014 (N_2014,N_1264,N_1413);
or U2015 (N_2015,N_1497,N_1556);
xor U2016 (N_2016,N_1317,N_1263);
and U2017 (N_2017,N_1713,N_1745);
or U2018 (N_2018,N_1755,N_1246);
and U2019 (N_2019,N_1652,N_1585);
and U2020 (N_2020,N_1542,N_1768);
nand U2021 (N_2021,N_1699,N_1753);
nor U2022 (N_2022,N_1515,N_1796);
nand U2023 (N_2023,N_1259,N_1282);
and U2024 (N_2024,N_1549,N_1307);
nand U2025 (N_2025,N_1603,N_1628);
and U2026 (N_2026,N_1595,N_1276);
nand U2027 (N_2027,N_1322,N_1391);
and U2028 (N_2028,N_1310,N_1518);
nand U2029 (N_2029,N_1608,N_1469);
nor U2030 (N_2030,N_1415,N_1400);
and U2031 (N_2031,N_1624,N_1221);
nand U2032 (N_2032,N_1663,N_1594);
nor U2033 (N_2033,N_1449,N_1328);
nor U2034 (N_2034,N_1743,N_1428);
and U2035 (N_2035,N_1709,N_1748);
and U2036 (N_2036,N_1558,N_1799);
and U2037 (N_2037,N_1696,N_1681);
and U2038 (N_2038,N_1605,N_1385);
or U2039 (N_2039,N_1775,N_1352);
or U2040 (N_2040,N_1733,N_1655);
xor U2041 (N_2041,N_1375,N_1379);
nor U2042 (N_2042,N_1658,N_1647);
or U2043 (N_2043,N_1365,N_1319);
nand U2044 (N_2044,N_1228,N_1717);
nor U2045 (N_2045,N_1389,N_1229);
nor U2046 (N_2046,N_1232,N_1793);
nor U2047 (N_2047,N_1723,N_1326);
nand U2048 (N_2048,N_1314,N_1355);
nor U2049 (N_2049,N_1292,N_1724);
nand U2050 (N_2050,N_1204,N_1483);
xnor U2051 (N_2051,N_1633,N_1784);
and U2052 (N_2052,N_1478,N_1450);
nand U2053 (N_2053,N_1454,N_1222);
or U2054 (N_2054,N_1440,N_1316);
nand U2055 (N_2055,N_1534,N_1255);
and U2056 (N_2056,N_1336,N_1616);
and U2057 (N_2057,N_1405,N_1250);
and U2058 (N_2058,N_1473,N_1520);
and U2059 (N_2059,N_1602,N_1684);
or U2060 (N_2060,N_1627,N_1371);
and U2061 (N_2061,N_1537,N_1592);
nor U2062 (N_2062,N_1760,N_1786);
or U2063 (N_2063,N_1286,N_1403);
nor U2064 (N_2064,N_1370,N_1509);
nor U2065 (N_2065,N_1280,N_1254);
nor U2066 (N_2066,N_1453,N_1789);
or U2067 (N_2067,N_1620,N_1417);
nor U2068 (N_2068,N_1634,N_1334);
nand U2069 (N_2069,N_1484,N_1752);
nor U2070 (N_2070,N_1329,N_1606);
and U2071 (N_2071,N_1660,N_1373);
nand U2072 (N_2072,N_1377,N_1590);
nor U2073 (N_2073,N_1588,N_1710);
xnor U2074 (N_2074,N_1563,N_1486);
and U2075 (N_2075,N_1235,N_1335);
nand U2076 (N_2076,N_1674,N_1456);
or U2077 (N_2077,N_1523,N_1686);
or U2078 (N_2078,N_1559,N_1512);
and U2079 (N_2079,N_1495,N_1203);
and U2080 (N_2080,N_1618,N_1342);
and U2081 (N_2081,N_1746,N_1312);
or U2082 (N_2082,N_1205,N_1503);
or U2083 (N_2083,N_1535,N_1429);
or U2084 (N_2084,N_1527,N_1357);
nand U2085 (N_2085,N_1657,N_1272);
nor U2086 (N_2086,N_1412,N_1302);
or U2087 (N_2087,N_1650,N_1578);
nor U2088 (N_2088,N_1343,N_1626);
nand U2089 (N_2089,N_1604,N_1363);
or U2090 (N_2090,N_1676,N_1582);
or U2091 (N_2091,N_1416,N_1526);
and U2092 (N_2092,N_1244,N_1623);
nand U2093 (N_2093,N_1480,N_1368);
nand U2094 (N_2094,N_1325,N_1372);
and U2095 (N_2095,N_1759,N_1356);
nand U2096 (N_2096,N_1574,N_1718);
nor U2097 (N_2097,N_1596,N_1661);
or U2098 (N_2098,N_1402,N_1725);
nand U2099 (N_2099,N_1288,N_1482);
nand U2100 (N_2100,N_1213,N_1353);
and U2101 (N_2101,N_1744,N_1313);
and U2102 (N_2102,N_1542,N_1481);
nor U2103 (N_2103,N_1631,N_1214);
nor U2104 (N_2104,N_1414,N_1332);
and U2105 (N_2105,N_1472,N_1214);
nand U2106 (N_2106,N_1758,N_1675);
or U2107 (N_2107,N_1350,N_1649);
nor U2108 (N_2108,N_1553,N_1279);
nand U2109 (N_2109,N_1660,N_1333);
nand U2110 (N_2110,N_1679,N_1704);
nand U2111 (N_2111,N_1222,N_1586);
and U2112 (N_2112,N_1588,N_1236);
and U2113 (N_2113,N_1601,N_1302);
and U2114 (N_2114,N_1790,N_1772);
nor U2115 (N_2115,N_1488,N_1453);
xnor U2116 (N_2116,N_1627,N_1286);
nor U2117 (N_2117,N_1450,N_1298);
nor U2118 (N_2118,N_1203,N_1214);
nor U2119 (N_2119,N_1704,N_1496);
nand U2120 (N_2120,N_1567,N_1700);
nand U2121 (N_2121,N_1685,N_1564);
and U2122 (N_2122,N_1201,N_1589);
nor U2123 (N_2123,N_1697,N_1361);
and U2124 (N_2124,N_1748,N_1554);
nor U2125 (N_2125,N_1334,N_1674);
and U2126 (N_2126,N_1589,N_1649);
nand U2127 (N_2127,N_1632,N_1690);
or U2128 (N_2128,N_1635,N_1279);
nand U2129 (N_2129,N_1220,N_1450);
and U2130 (N_2130,N_1573,N_1434);
or U2131 (N_2131,N_1505,N_1759);
nor U2132 (N_2132,N_1332,N_1313);
and U2133 (N_2133,N_1685,N_1613);
nor U2134 (N_2134,N_1559,N_1353);
and U2135 (N_2135,N_1475,N_1538);
nor U2136 (N_2136,N_1588,N_1573);
or U2137 (N_2137,N_1778,N_1662);
and U2138 (N_2138,N_1799,N_1724);
nor U2139 (N_2139,N_1580,N_1744);
xor U2140 (N_2140,N_1672,N_1367);
or U2141 (N_2141,N_1587,N_1257);
and U2142 (N_2142,N_1663,N_1478);
nor U2143 (N_2143,N_1477,N_1794);
and U2144 (N_2144,N_1774,N_1503);
nand U2145 (N_2145,N_1268,N_1431);
nand U2146 (N_2146,N_1379,N_1620);
and U2147 (N_2147,N_1537,N_1412);
nor U2148 (N_2148,N_1363,N_1628);
nor U2149 (N_2149,N_1525,N_1367);
nand U2150 (N_2150,N_1422,N_1660);
or U2151 (N_2151,N_1680,N_1385);
nand U2152 (N_2152,N_1706,N_1746);
nand U2153 (N_2153,N_1283,N_1475);
nor U2154 (N_2154,N_1705,N_1533);
nor U2155 (N_2155,N_1288,N_1280);
or U2156 (N_2156,N_1777,N_1657);
nor U2157 (N_2157,N_1327,N_1356);
nor U2158 (N_2158,N_1266,N_1337);
nand U2159 (N_2159,N_1312,N_1444);
or U2160 (N_2160,N_1262,N_1509);
and U2161 (N_2161,N_1703,N_1739);
nand U2162 (N_2162,N_1480,N_1340);
and U2163 (N_2163,N_1248,N_1263);
and U2164 (N_2164,N_1718,N_1572);
nand U2165 (N_2165,N_1584,N_1499);
and U2166 (N_2166,N_1771,N_1356);
and U2167 (N_2167,N_1517,N_1603);
and U2168 (N_2168,N_1749,N_1325);
or U2169 (N_2169,N_1268,N_1583);
nand U2170 (N_2170,N_1716,N_1345);
and U2171 (N_2171,N_1501,N_1753);
or U2172 (N_2172,N_1646,N_1793);
and U2173 (N_2173,N_1573,N_1689);
nor U2174 (N_2174,N_1579,N_1514);
or U2175 (N_2175,N_1213,N_1753);
nor U2176 (N_2176,N_1677,N_1753);
and U2177 (N_2177,N_1409,N_1324);
nand U2178 (N_2178,N_1430,N_1541);
or U2179 (N_2179,N_1369,N_1320);
nor U2180 (N_2180,N_1432,N_1473);
or U2181 (N_2181,N_1251,N_1246);
or U2182 (N_2182,N_1296,N_1349);
xor U2183 (N_2183,N_1554,N_1428);
and U2184 (N_2184,N_1299,N_1616);
xnor U2185 (N_2185,N_1597,N_1355);
nor U2186 (N_2186,N_1612,N_1276);
or U2187 (N_2187,N_1517,N_1771);
and U2188 (N_2188,N_1456,N_1540);
or U2189 (N_2189,N_1435,N_1732);
nor U2190 (N_2190,N_1654,N_1382);
or U2191 (N_2191,N_1230,N_1242);
or U2192 (N_2192,N_1417,N_1225);
nand U2193 (N_2193,N_1663,N_1645);
nor U2194 (N_2194,N_1730,N_1790);
nor U2195 (N_2195,N_1564,N_1614);
nand U2196 (N_2196,N_1314,N_1770);
and U2197 (N_2197,N_1227,N_1324);
nor U2198 (N_2198,N_1306,N_1622);
nand U2199 (N_2199,N_1256,N_1567);
or U2200 (N_2200,N_1350,N_1719);
nand U2201 (N_2201,N_1276,N_1480);
nand U2202 (N_2202,N_1429,N_1335);
and U2203 (N_2203,N_1254,N_1424);
xnor U2204 (N_2204,N_1766,N_1386);
nor U2205 (N_2205,N_1229,N_1768);
nor U2206 (N_2206,N_1495,N_1778);
nor U2207 (N_2207,N_1465,N_1229);
nand U2208 (N_2208,N_1407,N_1241);
and U2209 (N_2209,N_1391,N_1543);
nand U2210 (N_2210,N_1507,N_1237);
or U2211 (N_2211,N_1395,N_1284);
or U2212 (N_2212,N_1754,N_1454);
nor U2213 (N_2213,N_1771,N_1505);
nand U2214 (N_2214,N_1609,N_1400);
or U2215 (N_2215,N_1250,N_1665);
nand U2216 (N_2216,N_1738,N_1446);
and U2217 (N_2217,N_1371,N_1340);
nor U2218 (N_2218,N_1281,N_1289);
nand U2219 (N_2219,N_1285,N_1788);
nand U2220 (N_2220,N_1403,N_1695);
nor U2221 (N_2221,N_1326,N_1439);
and U2222 (N_2222,N_1316,N_1378);
and U2223 (N_2223,N_1390,N_1321);
or U2224 (N_2224,N_1768,N_1252);
nor U2225 (N_2225,N_1782,N_1775);
or U2226 (N_2226,N_1470,N_1526);
nand U2227 (N_2227,N_1384,N_1623);
and U2228 (N_2228,N_1740,N_1233);
and U2229 (N_2229,N_1331,N_1302);
nand U2230 (N_2230,N_1477,N_1250);
and U2231 (N_2231,N_1413,N_1278);
nor U2232 (N_2232,N_1276,N_1712);
nor U2233 (N_2233,N_1417,N_1697);
nor U2234 (N_2234,N_1471,N_1241);
or U2235 (N_2235,N_1760,N_1463);
nor U2236 (N_2236,N_1604,N_1513);
or U2237 (N_2237,N_1568,N_1693);
and U2238 (N_2238,N_1387,N_1551);
xor U2239 (N_2239,N_1417,N_1534);
nand U2240 (N_2240,N_1552,N_1462);
or U2241 (N_2241,N_1702,N_1464);
nor U2242 (N_2242,N_1580,N_1615);
or U2243 (N_2243,N_1591,N_1675);
xnor U2244 (N_2244,N_1270,N_1466);
nor U2245 (N_2245,N_1295,N_1744);
or U2246 (N_2246,N_1496,N_1682);
xnor U2247 (N_2247,N_1373,N_1626);
and U2248 (N_2248,N_1641,N_1720);
and U2249 (N_2249,N_1729,N_1289);
and U2250 (N_2250,N_1553,N_1236);
nor U2251 (N_2251,N_1392,N_1672);
nand U2252 (N_2252,N_1222,N_1448);
nand U2253 (N_2253,N_1608,N_1527);
nand U2254 (N_2254,N_1681,N_1538);
nand U2255 (N_2255,N_1495,N_1620);
or U2256 (N_2256,N_1703,N_1411);
xnor U2257 (N_2257,N_1555,N_1485);
or U2258 (N_2258,N_1324,N_1515);
or U2259 (N_2259,N_1554,N_1536);
nand U2260 (N_2260,N_1213,N_1462);
or U2261 (N_2261,N_1379,N_1321);
or U2262 (N_2262,N_1797,N_1668);
nor U2263 (N_2263,N_1762,N_1733);
and U2264 (N_2264,N_1455,N_1632);
and U2265 (N_2265,N_1740,N_1406);
nor U2266 (N_2266,N_1381,N_1421);
and U2267 (N_2267,N_1603,N_1481);
or U2268 (N_2268,N_1698,N_1618);
nand U2269 (N_2269,N_1265,N_1405);
xnor U2270 (N_2270,N_1475,N_1254);
nand U2271 (N_2271,N_1504,N_1323);
nand U2272 (N_2272,N_1269,N_1524);
or U2273 (N_2273,N_1786,N_1452);
nor U2274 (N_2274,N_1723,N_1414);
and U2275 (N_2275,N_1750,N_1641);
nand U2276 (N_2276,N_1781,N_1797);
and U2277 (N_2277,N_1659,N_1375);
and U2278 (N_2278,N_1598,N_1674);
or U2279 (N_2279,N_1340,N_1541);
nand U2280 (N_2280,N_1567,N_1508);
and U2281 (N_2281,N_1462,N_1497);
or U2282 (N_2282,N_1611,N_1509);
or U2283 (N_2283,N_1795,N_1255);
or U2284 (N_2284,N_1304,N_1537);
or U2285 (N_2285,N_1322,N_1310);
and U2286 (N_2286,N_1712,N_1322);
and U2287 (N_2287,N_1586,N_1647);
nor U2288 (N_2288,N_1344,N_1624);
nand U2289 (N_2289,N_1580,N_1346);
or U2290 (N_2290,N_1222,N_1211);
or U2291 (N_2291,N_1681,N_1533);
nand U2292 (N_2292,N_1447,N_1719);
nor U2293 (N_2293,N_1549,N_1566);
nand U2294 (N_2294,N_1609,N_1491);
nor U2295 (N_2295,N_1297,N_1483);
or U2296 (N_2296,N_1655,N_1303);
or U2297 (N_2297,N_1696,N_1600);
or U2298 (N_2298,N_1463,N_1443);
nand U2299 (N_2299,N_1654,N_1431);
or U2300 (N_2300,N_1240,N_1322);
and U2301 (N_2301,N_1642,N_1687);
nand U2302 (N_2302,N_1629,N_1575);
nor U2303 (N_2303,N_1790,N_1379);
nand U2304 (N_2304,N_1241,N_1388);
nor U2305 (N_2305,N_1386,N_1660);
or U2306 (N_2306,N_1218,N_1413);
or U2307 (N_2307,N_1624,N_1254);
nor U2308 (N_2308,N_1424,N_1697);
nor U2309 (N_2309,N_1633,N_1406);
or U2310 (N_2310,N_1263,N_1669);
nand U2311 (N_2311,N_1380,N_1271);
and U2312 (N_2312,N_1733,N_1511);
and U2313 (N_2313,N_1605,N_1216);
nand U2314 (N_2314,N_1630,N_1553);
nor U2315 (N_2315,N_1561,N_1610);
nand U2316 (N_2316,N_1747,N_1755);
and U2317 (N_2317,N_1696,N_1731);
nor U2318 (N_2318,N_1724,N_1712);
nor U2319 (N_2319,N_1359,N_1294);
or U2320 (N_2320,N_1572,N_1440);
nor U2321 (N_2321,N_1781,N_1615);
or U2322 (N_2322,N_1482,N_1325);
or U2323 (N_2323,N_1265,N_1436);
and U2324 (N_2324,N_1429,N_1707);
or U2325 (N_2325,N_1703,N_1444);
nand U2326 (N_2326,N_1482,N_1356);
or U2327 (N_2327,N_1689,N_1718);
nor U2328 (N_2328,N_1207,N_1705);
or U2329 (N_2329,N_1522,N_1660);
nand U2330 (N_2330,N_1699,N_1262);
nor U2331 (N_2331,N_1648,N_1605);
and U2332 (N_2332,N_1306,N_1608);
nor U2333 (N_2333,N_1471,N_1656);
or U2334 (N_2334,N_1323,N_1291);
and U2335 (N_2335,N_1617,N_1544);
or U2336 (N_2336,N_1306,N_1454);
or U2337 (N_2337,N_1770,N_1546);
nand U2338 (N_2338,N_1648,N_1510);
or U2339 (N_2339,N_1714,N_1405);
or U2340 (N_2340,N_1703,N_1612);
nand U2341 (N_2341,N_1409,N_1417);
nor U2342 (N_2342,N_1440,N_1523);
nor U2343 (N_2343,N_1503,N_1452);
or U2344 (N_2344,N_1272,N_1449);
nand U2345 (N_2345,N_1447,N_1202);
nand U2346 (N_2346,N_1799,N_1310);
or U2347 (N_2347,N_1367,N_1206);
xor U2348 (N_2348,N_1426,N_1590);
nand U2349 (N_2349,N_1585,N_1759);
or U2350 (N_2350,N_1362,N_1457);
nor U2351 (N_2351,N_1251,N_1688);
nand U2352 (N_2352,N_1758,N_1296);
nor U2353 (N_2353,N_1628,N_1549);
nor U2354 (N_2354,N_1513,N_1687);
nand U2355 (N_2355,N_1543,N_1477);
nand U2356 (N_2356,N_1206,N_1479);
nor U2357 (N_2357,N_1583,N_1697);
and U2358 (N_2358,N_1259,N_1560);
and U2359 (N_2359,N_1246,N_1636);
nor U2360 (N_2360,N_1307,N_1460);
and U2361 (N_2361,N_1300,N_1204);
nor U2362 (N_2362,N_1280,N_1690);
nor U2363 (N_2363,N_1385,N_1502);
or U2364 (N_2364,N_1634,N_1574);
nand U2365 (N_2365,N_1299,N_1469);
and U2366 (N_2366,N_1465,N_1213);
and U2367 (N_2367,N_1661,N_1494);
and U2368 (N_2368,N_1363,N_1302);
or U2369 (N_2369,N_1442,N_1755);
nor U2370 (N_2370,N_1248,N_1308);
xnor U2371 (N_2371,N_1247,N_1796);
or U2372 (N_2372,N_1559,N_1476);
nand U2373 (N_2373,N_1597,N_1567);
xnor U2374 (N_2374,N_1440,N_1329);
nor U2375 (N_2375,N_1378,N_1673);
nand U2376 (N_2376,N_1408,N_1653);
and U2377 (N_2377,N_1650,N_1381);
nand U2378 (N_2378,N_1678,N_1651);
nor U2379 (N_2379,N_1465,N_1245);
nor U2380 (N_2380,N_1670,N_1261);
or U2381 (N_2381,N_1570,N_1644);
nor U2382 (N_2382,N_1641,N_1374);
or U2383 (N_2383,N_1639,N_1735);
and U2384 (N_2384,N_1683,N_1482);
nand U2385 (N_2385,N_1342,N_1616);
nor U2386 (N_2386,N_1582,N_1408);
nand U2387 (N_2387,N_1329,N_1720);
nor U2388 (N_2388,N_1242,N_1589);
or U2389 (N_2389,N_1534,N_1595);
nand U2390 (N_2390,N_1307,N_1627);
nand U2391 (N_2391,N_1711,N_1358);
and U2392 (N_2392,N_1541,N_1496);
nor U2393 (N_2393,N_1773,N_1579);
nand U2394 (N_2394,N_1495,N_1634);
nand U2395 (N_2395,N_1651,N_1368);
and U2396 (N_2396,N_1565,N_1402);
nand U2397 (N_2397,N_1633,N_1599);
or U2398 (N_2398,N_1605,N_1288);
nor U2399 (N_2399,N_1733,N_1332);
and U2400 (N_2400,N_2280,N_2377);
and U2401 (N_2401,N_2143,N_2251);
nor U2402 (N_2402,N_1968,N_2317);
xnor U2403 (N_2403,N_2014,N_2253);
nand U2404 (N_2404,N_2157,N_2190);
nand U2405 (N_2405,N_2266,N_1920);
or U2406 (N_2406,N_1937,N_1829);
or U2407 (N_2407,N_2135,N_2325);
and U2408 (N_2408,N_2334,N_2025);
nor U2409 (N_2409,N_1967,N_2087);
or U2410 (N_2410,N_2374,N_2056);
and U2411 (N_2411,N_2298,N_2354);
nand U2412 (N_2412,N_1800,N_1921);
nor U2413 (N_2413,N_2053,N_2249);
or U2414 (N_2414,N_1962,N_2343);
nor U2415 (N_2415,N_1986,N_2282);
nor U2416 (N_2416,N_1878,N_2126);
and U2417 (N_2417,N_2389,N_1977);
nor U2418 (N_2418,N_1812,N_2122);
or U2419 (N_2419,N_2151,N_2236);
or U2420 (N_2420,N_2026,N_1973);
and U2421 (N_2421,N_1913,N_1814);
nand U2422 (N_2422,N_2082,N_2004);
or U2423 (N_2423,N_1892,N_1855);
nand U2424 (N_2424,N_2357,N_1882);
and U2425 (N_2425,N_2276,N_1999);
xnor U2426 (N_2426,N_1840,N_1988);
and U2427 (N_2427,N_1964,N_2286);
nand U2428 (N_2428,N_1843,N_2378);
or U2429 (N_2429,N_2302,N_1811);
or U2430 (N_2430,N_2081,N_2161);
or U2431 (N_2431,N_1950,N_1960);
nor U2432 (N_2432,N_1927,N_2146);
or U2433 (N_2433,N_2062,N_2133);
nand U2434 (N_2434,N_2398,N_2044);
nor U2435 (N_2435,N_1846,N_2244);
or U2436 (N_2436,N_2170,N_2273);
or U2437 (N_2437,N_2222,N_1865);
xnor U2438 (N_2438,N_2150,N_2364);
nor U2439 (N_2439,N_2338,N_1881);
and U2440 (N_2440,N_2371,N_1998);
or U2441 (N_2441,N_2326,N_2060);
and U2442 (N_2442,N_2093,N_1926);
xor U2443 (N_2443,N_2365,N_2215);
or U2444 (N_2444,N_2265,N_1871);
or U2445 (N_2445,N_2118,N_2221);
or U2446 (N_2446,N_1861,N_2305);
and U2447 (N_2447,N_2030,N_2277);
and U2448 (N_2448,N_2284,N_2156);
nor U2449 (N_2449,N_2099,N_2264);
or U2450 (N_2450,N_1987,N_1894);
and U2451 (N_2451,N_2392,N_1965);
nand U2452 (N_2452,N_2013,N_1990);
or U2453 (N_2453,N_1848,N_2106);
or U2454 (N_2454,N_2169,N_2176);
nand U2455 (N_2455,N_1922,N_2307);
or U2456 (N_2456,N_2173,N_2207);
nor U2457 (N_2457,N_2140,N_2333);
or U2458 (N_2458,N_2383,N_2361);
or U2459 (N_2459,N_1985,N_1859);
and U2460 (N_2460,N_1928,N_1895);
and U2461 (N_2461,N_2137,N_2035);
or U2462 (N_2462,N_1877,N_1948);
nor U2463 (N_2463,N_1810,N_2369);
nor U2464 (N_2464,N_2209,N_2022);
and U2465 (N_2465,N_2327,N_1803);
or U2466 (N_2466,N_2005,N_1958);
and U2467 (N_2467,N_2179,N_2310);
nor U2468 (N_2468,N_2163,N_2049);
nand U2469 (N_2469,N_1869,N_2104);
xnor U2470 (N_2470,N_2254,N_1849);
nand U2471 (N_2471,N_1902,N_2168);
and U2472 (N_2472,N_1864,N_2381);
nand U2473 (N_2473,N_1930,N_1969);
nor U2474 (N_2474,N_1815,N_2109);
nor U2475 (N_2475,N_2042,N_2091);
or U2476 (N_2476,N_2191,N_2145);
and U2477 (N_2477,N_1997,N_2233);
or U2478 (N_2478,N_1897,N_1956);
and U2479 (N_2479,N_2094,N_2351);
or U2480 (N_2480,N_1873,N_1908);
and U2481 (N_2481,N_2267,N_2029);
xor U2482 (N_2482,N_1876,N_2199);
or U2483 (N_2483,N_1917,N_2360);
nand U2484 (N_2484,N_2288,N_2153);
nand U2485 (N_2485,N_2041,N_2262);
nand U2486 (N_2486,N_2291,N_2011);
nor U2487 (N_2487,N_2188,N_2231);
or U2488 (N_2488,N_2385,N_2039);
nand U2489 (N_2489,N_2219,N_2373);
nor U2490 (N_2490,N_2223,N_2303);
nand U2491 (N_2491,N_2261,N_2217);
xor U2492 (N_2492,N_2071,N_1857);
and U2493 (N_2493,N_2050,N_2103);
xnor U2494 (N_2494,N_2387,N_2224);
nor U2495 (N_2495,N_1909,N_2319);
nand U2496 (N_2496,N_2289,N_2336);
and U2497 (N_2497,N_2388,N_1813);
or U2498 (N_2498,N_2293,N_2210);
and U2499 (N_2499,N_2355,N_2096);
and U2500 (N_2500,N_1945,N_2235);
xor U2501 (N_2501,N_2193,N_1842);
nand U2502 (N_2502,N_2154,N_1983);
or U2503 (N_2503,N_1961,N_1819);
and U2504 (N_2504,N_2084,N_1801);
nor U2505 (N_2505,N_1837,N_2362);
nand U2506 (N_2506,N_1872,N_2105);
nand U2507 (N_2507,N_2192,N_2036);
or U2508 (N_2508,N_2024,N_1888);
nand U2509 (N_2509,N_2008,N_1912);
or U2510 (N_2510,N_2088,N_1834);
and U2511 (N_2511,N_2034,N_2134);
and U2512 (N_2512,N_1805,N_1979);
or U2513 (N_2513,N_2020,N_2205);
or U2514 (N_2514,N_1978,N_1845);
or U2515 (N_2515,N_2229,N_1839);
or U2516 (N_2516,N_2363,N_1828);
nor U2517 (N_2517,N_2238,N_2358);
or U2518 (N_2518,N_2206,N_1899);
nor U2519 (N_2519,N_1953,N_2344);
or U2520 (N_2520,N_2194,N_2297);
nand U2521 (N_2521,N_2065,N_2144);
nor U2522 (N_2522,N_2306,N_2185);
nand U2523 (N_2523,N_2322,N_2195);
or U2524 (N_2524,N_2057,N_2074);
nand U2525 (N_2525,N_2021,N_1856);
or U2526 (N_2526,N_2337,N_2048);
and U2527 (N_2527,N_2038,N_2311);
and U2528 (N_2528,N_1809,N_2252);
nor U2529 (N_2529,N_1971,N_1949);
nand U2530 (N_2530,N_2308,N_1993);
nor U2531 (N_2531,N_2078,N_2067);
nor U2532 (N_2532,N_1893,N_2243);
and U2533 (N_2533,N_2032,N_2218);
and U2534 (N_2534,N_1932,N_2301);
or U2535 (N_2535,N_2001,N_2114);
and U2536 (N_2536,N_2077,N_2148);
nor U2537 (N_2537,N_2051,N_2058);
or U2538 (N_2538,N_2348,N_2250);
or U2539 (N_2539,N_1996,N_2290);
nand U2540 (N_2540,N_2023,N_2328);
or U2541 (N_2541,N_1889,N_2248);
nor U2542 (N_2542,N_2237,N_2376);
or U2543 (N_2543,N_1980,N_2059);
nor U2544 (N_2544,N_1884,N_1821);
or U2545 (N_2545,N_2108,N_1947);
or U2546 (N_2546,N_2182,N_1981);
and U2547 (N_2547,N_2230,N_2320);
and U2548 (N_2548,N_2197,N_2287);
or U2549 (N_2549,N_1954,N_2226);
and U2550 (N_2550,N_1943,N_2089);
nand U2551 (N_2551,N_2228,N_2342);
xnor U2552 (N_2552,N_2313,N_1853);
or U2553 (N_2553,N_1883,N_2040);
or U2554 (N_2554,N_1941,N_2072);
nand U2555 (N_2555,N_1989,N_1886);
xnor U2556 (N_2556,N_2012,N_1915);
nand U2557 (N_2557,N_2015,N_2183);
or U2558 (N_2558,N_2175,N_2246);
xnor U2559 (N_2559,N_2278,N_1833);
nand U2560 (N_2560,N_2214,N_2019);
nor U2561 (N_2561,N_2037,N_2349);
and U2562 (N_2562,N_1995,N_2119);
nor U2563 (N_2563,N_1804,N_2372);
nor U2564 (N_2564,N_1868,N_2227);
nor U2565 (N_2565,N_1885,N_2125);
nor U2566 (N_2566,N_1825,N_2394);
nor U2567 (N_2567,N_1816,N_2272);
nand U2568 (N_2568,N_1887,N_2115);
nand U2569 (N_2569,N_1982,N_2079);
or U2570 (N_2570,N_2332,N_2339);
nor U2571 (N_2571,N_2180,N_2159);
nor U2572 (N_2572,N_2189,N_1898);
nand U2573 (N_2573,N_1992,N_1820);
nand U2574 (N_2574,N_1931,N_2113);
nor U2575 (N_2575,N_1957,N_2356);
nand U2576 (N_2576,N_2028,N_2085);
or U2577 (N_2577,N_2080,N_1807);
nand U2578 (N_2578,N_2174,N_2257);
and U2579 (N_2579,N_1862,N_2139);
nor U2580 (N_2580,N_2341,N_1910);
or U2581 (N_2581,N_2340,N_1850);
nand U2582 (N_2582,N_1823,N_2256);
or U2583 (N_2583,N_2315,N_2110);
and U2584 (N_2584,N_1880,N_2142);
nand U2585 (N_2585,N_1827,N_2171);
nand U2586 (N_2586,N_2346,N_1901);
nand U2587 (N_2587,N_1806,N_1916);
nand U2588 (N_2588,N_1841,N_1907);
or U2589 (N_2589,N_1896,N_2211);
nand U2590 (N_2590,N_2285,N_2070);
nor U2591 (N_2591,N_2043,N_1914);
or U2592 (N_2592,N_1972,N_2352);
nand U2593 (N_2593,N_2031,N_1890);
or U2594 (N_2594,N_1852,N_1970);
and U2595 (N_2595,N_2124,N_2129);
nor U2596 (N_2596,N_1903,N_2395);
nor U2597 (N_2597,N_1938,N_1963);
nor U2598 (N_2598,N_1940,N_2164);
nor U2599 (N_2599,N_2239,N_2397);
nor U2600 (N_2600,N_2138,N_1911);
nor U2601 (N_2601,N_2380,N_2123);
or U2602 (N_2602,N_1946,N_1984);
and U2603 (N_2603,N_1994,N_1900);
nor U2604 (N_2604,N_2331,N_2064);
nand U2605 (N_2605,N_2006,N_1874);
nand U2606 (N_2606,N_1847,N_2324);
nor U2607 (N_2607,N_2158,N_1830);
nand U2608 (N_2608,N_2240,N_1860);
or U2609 (N_2609,N_2132,N_2366);
or U2610 (N_2610,N_2329,N_2271);
or U2611 (N_2611,N_2116,N_2172);
or U2612 (N_2612,N_2054,N_2283);
nand U2613 (N_2613,N_1944,N_2225);
nand U2614 (N_2614,N_2255,N_1918);
nand U2615 (N_2615,N_2263,N_2370);
nand U2616 (N_2616,N_1923,N_2202);
or U2617 (N_2617,N_2314,N_2130);
nor U2618 (N_2618,N_2242,N_2162);
and U2619 (N_2619,N_1906,N_1976);
nand U2620 (N_2620,N_2127,N_2068);
or U2621 (N_2621,N_1929,N_2399);
nor U2622 (N_2622,N_2075,N_2347);
nor U2623 (N_2623,N_2165,N_2018);
and U2624 (N_2624,N_2367,N_1951);
nand U2625 (N_2625,N_2198,N_1866);
nand U2626 (N_2626,N_2294,N_2178);
nor U2627 (N_2627,N_1808,N_2083);
nand U2628 (N_2628,N_1933,N_2033);
or U2629 (N_2629,N_1925,N_2292);
and U2630 (N_2630,N_1818,N_2121);
xnor U2631 (N_2631,N_2186,N_2149);
nor U2632 (N_2632,N_2384,N_2187);
nor U2633 (N_2633,N_2396,N_1924);
xnor U2634 (N_2634,N_2275,N_2316);
and U2635 (N_2635,N_1935,N_1858);
or U2636 (N_2636,N_2181,N_2300);
or U2637 (N_2637,N_2321,N_2312);
nor U2638 (N_2638,N_1905,N_2274);
and U2639 (N_2639,N_1952,N_2258);
and U2640 (N_2640,N_2241,N_1870);
or U2641 (N_2641,N_1939,N_1959);
and U2642 (N_2642,N_2009,N_2147);
and U2643 (N_2643,N_1838,N_2259);
and U2644 (N_2644,N_2016,N_2111);
xnor U2645 (N_2645,N_2167,N_2027);
nand U2646 (N_2646,N_2117,N_1863);
and U2647 (N_2647,N_2155,N_2391);
nand U2648 (N_2648,N_2345,N_1832);
nand U2649 (N_2649,N_2017,N_2216);
and U2650 (N_2650,N_2063,N_2152);
nor U2651 (N_2651,N_2232,N_1891);
and U2652 (N_2652,N_2112,N_2330);
nand U2653 (N_2653,N_2390,N_2386);
and U2654 (N_2654,N_2003,N_2128);
and U2655 (N_2655,N_2304,N_2069);
nor U2656 (N_2656,N_2368,N_2200);
and U2657 (N_2657,N_1879,N_2196);
and U2658 (N_2658,N_2220,N_2382);
or U2659 (N_2659,N_1974,N_1867);
or U2660 (N_2660,N_2101,N_2086);
or U2661 (N_2661,N_1904,N_2203);
and U2662 (N_2662,N_2100,N_2201);
nand U2663 (N_2663,N_2076,N_2000);
nand U2664 (N_2664,N_1822,N_2213);
or U2665 (N_2665,N_1836,N_1991);
xnor U2666 (N_2666,N_2296,N_2045);
nor U2667 (N_2667,N_2073,N_1955);
or U2668 (N_2668,N_2212,N_2007);
or U2669 (N_2669,N_2177,N_1835);
nor U2670 (N_2670,N_2097,N_1919);
nand U2671 (N_2671,N_2141,N_2204);
or U2672 (N_2672,N_2269,N_2061);
and U2673 (N_2673,N_1826,N_2107);
or U2674 (N_2674,N_2234,N_2055);
and U2675 (N_2675,N_2208,N_2047);
nand U2676 (N_2676,N_2098,N_2318);
or U2677 (N_2677,N_2095,N_1942);
and U2678 (N_2678,N_1817,N_2046);
nand U2679 (N_2679,N_2002,N_2245);
nor U2680 (N_2680,N_2010,N_1966);
or U2681 (N_2681,N_2131,N_2052);
nand U2682 (N_2682,N_2268,N_2120);
nor U2683 (N_2683,N_1824,N_2375);
and U2684 (N_2684,N_2335,N_2299);
or U2685 (N_2685,N_2166,N_1844);
nand U2686 (N_2686,N_1875,N_1936);
or U2687 (N_2687,N_2160,N_2359);
and U2688 (N_2688,N_2281,N_2393);
nor U2689 (N_2689,N_2279,N_2136);
nand U2690 (N_2690,N_2102,N_1934);
or U2691 (N_2691,N_2353,N_2066);
nand U2692 (N_2692,N_1854,N_2090);
and U2693 (N_2693,N_2309,N_2092);
and U2694 (N_2694,N_2270,N_2260);
nor U2695 (N_2695,N_1851,N_2247);
nand U2696 (N_2696,N_1831,N_1802);
nand U2697 (N_2697,N_2184,N_2379);
nand U2698 (N_2698,N_2350,N_2295);
and U2699 (N_2699,N_1975,N_2323);
and U2700 (N_2700,N_2344,N_2134);
and U2701 (N_2701,N_2394,N_2363);
or U2702 (N_2702,N_1899,N_2006);
and U2703 (N_2703,N_1910,N_2123);
and U2704 (N_2704,N_2137,N_1976);
nand U2705 (N_2705,N_2218,N_1963);
xor U2706 (N_2706,N_2328,N_2313);
nand U2707 (N_2707,N_2318,N_2036);
nand U2708 (N_2708,N_1981,N_2378);
and U2709 (N_2709,N_2128,N_1953);
nand U2710 (N_2710,N_1992,N_2106);
xnor U2711 (N_2711,N_2175,N_2085);
and U2712 (N_2712,N_2074,N_2210);
nor U2713 (N_2713,N_2024,N_2247);
nor U2714 (N_2714,N_1927,N_1832);
and U2715 (N_2715,N_1988,N_1983);
nor U2716 (N_2716,N_1950,N_2125);
nor U2717 (N_2717,N_1894,N_2221);
nand U2718 (N_2718,N_1851,N_2240);
nor U2719 (N_2719,N_2115,N_1878);
xor U2720 (N_2720,N_2254,N_2161);
and U2721 (N_2721,N_2048,N_1931);
nor U2722 (N_2722,N_2179,N_2363);
or U2723 (N_2723,N_2014,N_2047);
and U2724 (N_2724,N_1837,N_1908);
and U2725 (N_2725,N_1811,N_1915);
or U2726 (N_2726,N_2020,N_2282);
nor U2727 (N_2727,N_1827,N_2119);
nand U2728 (N_2728,N_2369,N_2172);
and U2729 (N_2729,N_1920,N_1989);
and U2730 (N_2730,N_2210,N_1845);
and U2731 (N_2731,N_2158,N_2234);
or U2732 (N_2732,N_2338,N_2093);
nor U2733 (N_2733,N_2174,N_2236);
or U2734 (N_2734,N_2010,N_2085);
nand U2735 (N_2735,N_2295,N_2119);
nor U2736 (N_2736,N_2072,N_1807);
nor U2737 (N_2737,N_2211,N_1832);
and U2738 (N_2738,N_1962,N_1869);
nor U2739 (N_2739,N_2339,N_2287);
nor U2740 (N_2740,N_2364,N_2226);
nand U2741 (N_2741,N_1986,N_2299);
nand U2742 (N_2742,N_2169,N_2390);
nor U2743 (N_2743,N_1987,N_2194);
xor U2744 (N_2744,N_2091,N_2114);
or U2745 (N_2745,N_2248,N_2363);
nor U2746 (N_2746,N_1858,N_1832);
xnor U2747 (N_2747,N_2277,N_2335);
or U2748 (N_2748,N_1882,N_2003);
or U2749 (N_2749,N_1960,N_2144);
or U2750 (N_2750,N_2190,N_1872);
nor U2751 (N_2751,N_2120,N_1892);
nand U2752 (N_2752,N_2318,N_1801);
and U2753 (N_2753,N_1906,N_2341);
nand U2754 (N_2754,N_2122,N_2130);
or U2755 (N_2755,N_2158,N_2324);
nand U2756 (N_2756,N_2381,N_2012);
nand U2757 (N_2757,N_1997,N_2310);
and U2758 (N_2758,N_1975,N_1833);
nand U2759 (N_2759,N_1876,N_2069);
or U2760 (N_2760,N_1921,N_2234);
and U2761 (N_2761,N_2047,N_1843);
xnor U2762 (N_2762,N_2128,N_2231);
nor U2763 (N_2763,N_1819,N_2103);
or U2764 (N_2764,N_1851,N_2369);
or U2765 (N_2765,N_2395,N_2150);
nor U2766 (N_2766,N_2269,N_2217);
or U2767 (N_2767,N_2131,N_2343);
or U2768 (N_2768,N_2349,N_2207);
nor U2769 (N_2769,N_2141,N_1999);
nor U2770 (N_2770,N_2139,N_2308);
or U2771 (N_2771,N_2077,N_1852);
nor U2772 (N_2772,N_1858,N_1810);
nor U2773 (N_2773,N_2314,N_2394);
and U2774 (N_2774,N_2045,N_1823);
nor U2775 (N_2775,N_1880,N_1984);
or U2776 (N_2776,N_2031,N_2123);
and U2777 (N_2777,N_2104,N_2340);
and U2778 (N_2778,N_2207,N_2329);
or U2779 (N_2779,N_2382,N_2015);
nand U2780 (N_2780,N_2266,N_1972);
nand U2781 (N_2781,N_2244,N_2181);
nor U2782 (N_2782,N_2211,N_2217);
or U2783 (N_2783,N_1847,N_1861);
or U2784 (N_2784,N_2329,N_1847);
and U2785 (N_2785,N_2309,N_2304);
nor U2786 (N_2786,N_2390,N_2322);
nor U2787 (N_2787,N_2380,N_2175);
nand U2788 (N_2788,N_2028,N_2001);
nor U2789 (N_2789,N_2030,N_2114);
xnor U2790 (N_2790,N_1950,N_2147);
nor U2791 (N_2791,N_2310,N_2134);
nand U2792 (N_2792,N_2120,N_2249);
nand U2793 (N_2793,N_2121,N_1855);
nor U2794 (N_2794,N_2217,N_2259);
nand U2795 (N_2795,N_1996,N_2011);
or U2796 (N_2796,N_1803,N_2142);
nor U2797 (N_2797,N_2176,N_1831);
or U2798 (N_2798,N_1824,N_1942);
nor U2799 (N_2799,N_1907,N_1858);
and U2800 (N_2800,N_1901,N_2348);
or U2801 (N_2801,N_2282,N_2161);
and U2802 (N_2802,N_1988,N_2119);
nor U2803 (N_2803,N_2362,N_1998);
and U2804 (N_2804,N_2238,N_2284);
nand U2805 (N_2805,N_2321,N_1976);
nor U2806 (N_2806,N_2232,N_1988);
and U2807 (N_2807,N_2174,N_1803);
or U2808 (N_2808,N_2101,N_1933);
xnor U2809 (N_2809,N_2236,N_2089);
nor U2810 (N_2810,N_2322,N_2242);
xnor U2811 (N_2811,N_2222,N_2374);
nand U2812 (N_2812,N_1822,N_2316);
nor U2813 (N_2813,N_2352,N_2106);
nand U2814 (N_2814,N_1885,N_2369);
nor U2815 (N_2815,N_1825,N_2183);
or U2816 (N_2816,N_2199,N_2275);
or U2817 (N_2817,N_2188,N_1971);
nor U2818 (N_2818,N_1895,N_1953);
xor U2819 (N_2819,N_1846,N_2229);
nor U2820 (N_2820,N_2232,N_1837);
or U2821 (N_2821,N_1973,N_2220);
and U2822 (N_2822,N_2241,N_1829);
nand U2823 (N_2823,N_1914,N_2069);
xor U2824 (N_2824,N_2363,N_1874);
nand U2825 (N_2825,N_2340,N_2152);
or U2826 (N_2826,N_2082,N_2084);
nor U2827 (N_2827,N_2299,N_1813);
or U2828 (N_2828,N_2173,N_1874);
nor U2829 (N_2829,N_1932,N_2198);
xnor U2830 (N_2830,N_2099,N_2000);
nand U2831 (N_2831,N_2354,N_1939);
nor U2832 (N_2832,N_2221,N_2094);
or U2833 (N_2833,N_1887,N_2314);
nor U2834 (N_2834,N_2092,N_2217);
or U2835 (N_2835,N_2226,N_1930);
nand U2836 (N_2836,N_2061,N_2007);
or U2837 (N_2837,N_2321,N_2005);
and U2838 (N_2838,N_2341,N_1918);
and U2839 (N_2839,N_2012,N_2086);
nand U2840 (N_2840,N_2065,N_2289);
or U2841 (N_2841,N_1860,N_1853);
nand U2842 (N_2842,N_2363,N_2393);
and U2843 (N_2843,N_2024,N_2066);
and U2844 (N_2844,N_1942,N_2068);
or U2845 (N_2845,N_1923,N_1905);
or U2846 (N_2846,N_1865,N_2087);
and U2847 (N_2847,N_2267,N_1975);
or U2848 (N_2848,N_2326,N_2168);
nand U2849 (N_2849,N_2236,N_1923);
nor U2850 (N_2850,N_2079,N_2216);
or U2851 (N_2851,N_2329,N_1823);
nand U2852 (N_2852,N_1898,N_2100);
nand U2853 (N_2853,N_1801,N_2279);
nand U2854 (N_2854,N_2297,N_1930);
nor U2855 (N_2855,N_2022,N_2056);
and U2856 (N_2856,N_1831,N_2390);
or U2857 (N_2857,N_2035,N_1848);
and U2858 (N_2858,N_2219,N_2275);
and U2859 (N_2859,N_2213,N_1865);
or U2860 (N_2860,N_2205,N_1966);
xnor U2861 (N_2861,N_2239,N_1960);
or U2862 (N_2862,N_2258,N_1978);
xor U2863 (N_2863,N_2107,N_1904);
or U2864 (N_2864,N_2017,N_1887);
nand U2865 (N_2865,N_2026,N_2281);
or U2866 (N_2866,N_2287,N_2375);
nand U2867 (N_2867,N_2385,N_1802);
and U2868 (N_2868,N_2255,N_1959);
and U2869 (N_2869,N_1800,N_2298);
nand U2870 (N_2870,N_2165,N_2145);
nand U2871 (N_2871,N_1830,N_2215);
nand U2872 (N_2872,N_2182,N_2303);
or U2873 (N_2873,N_1962,N_2349);
nor U2874 (N_2874,N_2101,N_2121);
nand U2875 (N_2875,N_2396,N_2392);
nor U2876 (N_2876,N_2004,N_2311);
nand U2877 (N_2877,N_2231,N_2332);
nand U2878 (N_2878,N_1953,N_1840);
xnor U2879 (N_2879,N_1984,N_2200);
nand U2880 (N_2880,N_2331,N_1810);
and U2881 (N_2881,N_2048,N_2037);
and U2882 (N_2882,N_2025,N_1861);
or U2883 (N_2883,N_2346,N_1871);
nor U2884 (N_2884,N_2166,N_1913);
nor U2885 (N_2885,N_2144,N_1840);
or U2886 (N_2886,N_2124,N_1947);
and U2887 (N_2887,N_2201,N_1997);
or U2888 (N_2888,N_2178,N_2112);
and U2889 (N_2889,N_2115,N_2301);
nor U2890 (N_2890,N_2141,N_2265);
nor U2891 (N_2891,N_2396,N_2379);
nand U2892 (N_2892,N_2158,N_1938);
xnor U2893 (N_2893,N_1895,N_2100);
or U2894 (N_2894,N_2233,N_2325);
nand U2895 (N_2895,N_2022,N_1835);
xnor U2896 (N_2896,N_1804,N_2244);
nand U2897 (N_2897,N_2372,N_1916);
and U2898 (N_2898,N_2042,N_1870);
nand U2899 (N_2899,N_2300,N_2014);
and U2900 (N_2900,N_2087,N_1836);
nand U2901 (N_2901,N_2394,N_1993);
nor U2902 (N_2902,N_2112,N_1893);
or U2903 (N_2903,N_1809,N_1847);
and U2904 (N_2904,N_2334,N_2203);
nand U2905 (N_2905,N_2252,N_1914);
and U2906 (N_2906,N_2142,N_1910);
nand U2907 (N_2907,N_1815,N_1861);
nand U2908 (N_2908,N_2168,N_1933);
or U2909 (N_2909,N_2376,N_1823);
nor U2910 (N_2910,N_2032,N_2049);
and U2911 (N_2911,N_1965,N_1810);
or U2912 (N_2912,N_2052,N_2097);
nor U2913 (N_2913,N_2103,N_1947);
or U2914 (N_2914,N_1946,N_2146);
nor U2915 (N_2915,N_2349,N_1802);
nand U2916 (N_2916,N_2183,N_1907);
nand U2917 (N_2917,N_2308,N_2068);
nand U2918 (N_2918,N_2228,N_2224);
xor U2919 (N_2919,N_1898,N_1811);
xor U2920 (N_2920,N_2048,N_2314);
and U2921 (N_2921,N_2033,N_2220);
or U2922 (N_2922,N_2017,N_2202);
and U2923 (N_2923,N_2003,N_2119);
nand U2924 (N_2924,N_1902,N_1946);
or U2925 (N_2925,N_1904,N_2341);
and U2926 (N_2926,N_2064,N_2133);
and U2927 (N_2927,N_2183,N_2025);
xnor U2928 (N_2928,N_2241,N_2360);
or U2929 (N_2929,N_1838,N_2087);
nand U2930 (N_2930,N_1821,N_2137);
nor U2931 (N_2931,N_2077,N_1806);
nor U2932 (N_2932,N_1913,N_1943);
and U2933 (N_2933,N_2235,N_2028);
or U2934 (N_2934,N_1868,N_2211);
or U2935 (N_2935,N_2166,N_1931);
and U2936 (N_2936,N_1915,N_1947);
or U2937 (N_2937,N_1862,N_1979);
or U2938 (N_2938,N_2270,N_2313);
xnor U2939 (N_2939,N_2290,N_2294);
or U2940 (N_2940,N_2213,N_2357);
and U2941 (N_2941,N_2109,N_1859);
nand U2942 (N_2942,N_1892,N_1802);
nor U2943 (N_2943,N_2386,N_2053);
and U2944 (N_2944,N_2399,N_1805);
or U2945 (N_2945,N_2113,N_1811);
or U2946 (N_2946,N_2066,N_1931);
nand U2947 (N_2947,N_2118,N_1847);
or U2948 (N_2948,N_1911,N_2393);
nand U2949 (N_2949,N_2189,N_2108);
or U2950 (N_2950,N_2395,N_2028);
nand U2951 (N_2951,N_2342,N_2062);
nor U2952 (N_2952,N_1850,N_2387);
nor U2953 (N_2953,N_1800,N_2367);
or U2954 (N_2954,N_1834,N_2094);
nor U2955 (N_2955,N_1997,N_2032);
and U2956 (N_2956,N_2164,N_2211);
xnor U2957 (N_2957,N_2370,N_1887);
nor U2958 (N_2958,N_1994,N_1943);
and U2959 (N_2959,N_2372,N_1899);
nor U2960 (N_2960,N_2282,N_2332);
or U2961 (N_2961,N_2216,N_2241);
nor U2962 (N_2962,N_1811,N_2005);
nor U2963 (N_2963,N_1821,N_2206);
nand U2964 (N_2964,N_1986,N_1858);
or U2965 (N_2965,N_2323,N_2349);
and U2966 (N_2966,N_2211,N_1880);
nor U2967 (N_2967,N_2082,N_1967);
nand U2968 (N_2968,N_2204,N_2182);
nor U2969 (N_2969,N_1956,N_1870);
or U2970 (N_2970,N_1928,N_2077);
nand U2971 (N_2971,N_1936,N_2394);
and U2972 (N_2972,N_2029,N_1819);
nand U2973 (N_2973,N_1840,N_1836);
or U2974 (N_2974,N_1849,N_1944);
and U2975 (N_2975,N_2294,N_2237);
or U2976 (N_2976,N_1993,N_2389);
nand U2977 (N_2977,N_1975,N_2110);
and U2978 (N_2978,N_2011,N_2083);
and U2979 (N_2979,N_1891,N_2017);
nor U2980 (N_2980,N_2178,N_2130);
nor U2981 (N_2981,N_2208,N_2071);
nor U2982 (N_2982,N_1866,N_1913);
and U2983 (N_2983,N_2206,N_2155);
and U2984 (N_2984,N_1880,N_1978);
and U2985 (N_2985,N_1963,N_2078);
nor U2986 (N_2986,N_2282,N_1853);
nor U2987 (N_2987,N_2389,N_2014);
and U2988 (N_2988,N_2177,N_2285);
nand U2989 (N_2989,N_1896,N_2348);
nand U2990 (N_2990,N_2221,N_1800);
and U2991 (N_2991,N_2162,N_1809);
or U2992 (N_2992,N_1823,N_2129);
and U2993 (N_2993,N_2322,N_2087);
nand U2994 (N_2994,N_2324,N_2350);
nor U2995 (N_2995,N_2097,N_2383);
nor U2996 (N_2996,N_1818,N_1904);
and U2997 (N_2997,N_1935,N_2345);
nor U2998 (N_2998,N_2376,N_2022);
nand U2999 (N_2999,N_2393,N_2369);
nor UO_0 (O_0,N_2578,N_2459);
and UO_1 (O_1,N_2886,N_2999);
or UO_2 (O_2,N_2761,N_2877);
and UO_3 (O_3,N_2815,N_2585);
and UO_4 (O_4,N_2705,N_2837);
nor UO_5 (O_5,N_2954,N_2703);
and UO_6 (O_6,N_2612,N_2456);
nand UO_7 (O_7,N_2532,N_2723);
nor UO_8 (O_8,N_2697,N_2783);
or UO_9 (O_9,N_2590,N_2662);
nor UO_10 (O_10,N_2484,N_2831);
and UO_11 (O_11,N_2643,N_2843);
nand UO_12 (O_12,N_2556,N_2919);
nor UO_13 (O_13,N_2911,N_2602);
nor UO_14 (O_14,N_2838,N_2944);
and UO_15 (O_15,N_2908,N_2460);
nand UO_16 (O_16,N_2547,N_2902);
nor UO_17 (O_17,N_2782,N_2762);
nor UO_18 (O_18,N_2490,N_2404);
nand UO_19 (O_19,N_2409,N_2882);
nand UO_20 (O_20,N_2511,N_2934);
nand UO_21 (O_21,N_2966,N_2881);
nand UO_22 (O_22,N_2770,N_2870);
and UO_23 (O_23,N_2403,N_2763);
or UO_24 (O_24,N_2415,N_2480);
nand UO_25 (O_25,N_2854,N_2827);
or UO_26 (O_26,N_2833,N_2978);
nand UO_27 (O_27,N_2533,N_2803);
nand UO_28 (O_28,N_2988,N_2563);
nand UO_29 (O_29,N_2936,N_2917);
and UO_30 (O_30,N_2967,N_2401);
or UO_31 (O_31,N_2990,N_2771);
xor UO_32 (O_32,N_2669,N_2892);
and UO_33 (O_33,N_2501,N_2435);
or UO_34 (O_34,N_2644,N_2949);
and UO_35 (O_35,N_2981,N_2737);
nor UO_36 (O_36,N_2494,N_2743);
and UO_37 (O_37,N_2959,N_2577);
and UO_38 (O_38,N_2795,N_2668);
nor UO_39 (O_39,N_2557,N_2876);
nand UO_40 (O_40,N_2451,N_2727);
or UO_41 (O_41,N_2961,N_2735);
nand UO_42 (O_42,N_2586,N_2527);
or UO_43 (O_43,N_2745,N_2521);
nor UO_44 (O_44,N_2498,N_2613);
nor UO_45 (O_45,N_2823,N_2879);
or UO_46 (O_46,N_2710,N_2913);
or UO_47 (O_47,N_2589,N_2901);
or UO_48 (O_48,N_2410,N_2458);
nor UO_49 (O_49,N_2638,N_2564);
and UO_50 (O_50,N_2692,N_2926);
nor UO_51 (O_51,N_2765,N_2839);
and UO_52 (O_52,N_2847,N_2660);
nand UO_53 (O_53,N_2529,N_2817);
xnor UO_54 (O_54,N_2989,N_2943);
and UO_55 (O_55,N_2719,N_2848);
nor UO_56 (O_56,N_2894,N_2706);
or UO_57 (O_57,N_2522,N_2849);
and UO_58 (O_58,N_2555,N_2691);
and UO_59 (O_59,N_2536,N_2704);
nand UO_60 (O_60,N_2641,N_2813);
or UO_61 (O_61,N_2429,N_2627);
and UO_62 (O_62,N_2587,N_2463);
xor UO_63 (O_63,N_2957,N_2654);
nand UO_64 (O_64,N_2543,N_2445);
nand UO_65 (O_65,N_2758,N_2678);
or UO_66 (O_66,N_2581,N_2407);
or UO_67 (O_67,N_2768,N_2434);
or UO_68 (O_68,N_2576,N_2506);
nand UO_69 (O_69,N_2729,N_2732);
nand UO_70 (O_70,N_2424,N_2816);
nand UO_71 (O_71,N_2888,N_2568);
nand UO_72 (O_72,N_2979,N_2673);
and UO_73 (O_73,N_2773,N_2923);
and UO_74 (O_74,N_2826,N_2998);
nor UO_75 (O_75,N_2916,N_2753);
nor UO_76 (O_76,N_2977,N_2452);
or UO_77 (O_77,N_2534,N_2559);
or UO_78 (O_78,N_2714,N_2797);
or UO_79 (O_79,N_2575,N_2971);
nand UO_80 (O_80,N_2596,N_2930);
or UO_81 (O_81,N_2465,N_2679);
or UO_82 (O_82,N_2814,N_2818);
nand UO_83 (O_83,N_2799,N_2804);
nand UO_84 (O_84,N_2860,N_2756);
xnor UO_85 (O_85,N_2976,N_2423);
or UO_86 (O_86,N_2698,N_2927);
nor UO_87 (O_87,N_2680,N_2426);
nand UO_88 (O_88,N_2552,N_2523);
nor UO_89 (O_89,N_2507,N_2965);
nor UO_90 (O_90,N_2752,N_2497);
or UO_91 (O_91,N_2566,N_2608);
nand UO_92 (O_92,N_2525,N_2953);
or UO_93 (O_93,N_2938,N_2801);
nor UO_94 (O_94,N_2531,N_2647);
nor UO_95 (O_95,N_2755,N_2866);
and UO_96 (O_96,N_2477,N_2614);
and UO_97 (O_97,N_2569,N_2677);
and UO_98 (O_98,N_2747,N_2515);
nor UO_99 (O_99,N_2562,N_2832);
and UO_100 (O_100,N_2650,N_2964);
xnor UO_101 (O_101,N_2702,N_2545);
nand UO_102 (O_102,N_2489,N_2715);
nand UO_103 (O_103,N_2995,N_2819);
nor UO_104 (O_104,N_2800,N_2991);
nor UO_105 (O_105,N_2872,N_2798);
nor UO_106 (O_106,N_2645,N_2775);
nor UO_107 (O_107,N_2655,N_2418);
or UO_108 (O_108,N_2925,N_2609);
or UO_109 (O_109,N_2924,N_2402);
xnor UO_110 (O_110,N_2840,N_2659);
and UO_111 (O_111,N_2666,N_2920);
nor UO_112 (O_112,N_2736,N_2883);
nor UO_113 (O_113,N_2946,N_2457);
nand UO_114 (O_114,N_2658,N_2950);
nand UO_115 (O_115,N_2885,N_2663);
and UO_116 (O_116,N_2520,N_2621);
nand UO_117 (O_117,N_2859,N_2631);
nor UO_118 (O_118,N_2963,N_2975);
nand UO_119 (O_119,N_2896,N_2842);
nand UO_120 (O_120,N_2425,N_2772);
and UO_121 (O_121,N_2906,N_2852);
xor UO_122 (O_122,N_2665,N_2582);
or UO_123 (O_123,N_2437,N_2649);
nand UO_124 (O_124,N_2508,N_2416);
nor UO_125 (O_125,N_2895,N_2897);
nand UO_126 (O_126,N_2873,N_2808);
or UO_127 (O_127,N_2462,N_2629);
and UO_128 (O_128,N_2742,N_2603);
or UO_129 (O_129,N_2535,N_2574);
nand UO_130 (O_130,N_2730,N_2793);
nand UO_131 (O_131,N_2413,N_2802);
nor UO_132 (O_132,N_2540,N_2855);
nand UO_133 (O_133,N_2811,N_2444);
nor UO_134 (O_134,N_2648,N_2996);
nand UO_135 (O_135,N_2661,N_2900);
nor UO_136 (O_136,N_2769,N_2514);
and UO_137 (O_137,N_2518,N_2734);
nor UO_138 (O_138,N_2790,N_2664);
nand UO_139 (O_139,N_2986,N_2420);
nor UO_140 (O_140,N_2604,N_2711);
or UO_141 (O_141,N_2640,N_2476);
nand UO_142 (O_142,N_2740,N_2720);
or UO_143 (O_143,N_2421,N_2724);
nor UO_144 (O_144,N_2709,N_2549);
or UO_145 (O_145,N_2594,N_2526);
and UO_146 (O_146,N_2903,N_2683);
nand UO_147 (O_147,N_2670,N_2467);
nand UO_148 (O_148,N_2905,N_2980);
or UO_149 (O_149,N_2937,N_2622);
nor UO_150 (O_150,N_2942,N_2405);
or UO_151 (O_151,N_2750,N_2513);
and UO_152 (O_152,N_2955,N_2721);
nand UO_153 (O_153,N_2824,N_2992);
nor UO_154 (O_154,N_2759,N_2579);
and UO_155 (O_155,N_2417,N_2940);
nor UO_156 (O_156,N_2931,N_2438);
nor UO_157 (O_157,N_2646,N_2561);
or UO_158 (O_158,N_2779,N_2496);
nand UO_159 (O_159,N_2858,N_2466);
nand UO_160 (O_160,N_2400,N_2810);
and UO_161 (O_161,N_2947,N_2909);
or UO_162 (O_162,N_2812,N_2478);
nand UO_163 (O_163,N_2760,N_2567);
or UO_164 (O_164,N_2442,N_2542);
nor UO_165 (O_165,N_2461,N_2516);
and UO_166 (O_166,N_2408,N_2470);
and UO_167 (O_167,N_2972,N_2548);
or UO_168 (O_168,N_2541,N_2699);
nand UO_169 (O_169,N_2597,N_2583);
or UO_170 (O_170,N_2898,N_2486);
nand UO_171 (O_171,N_2777,N_2483);
and UO_172 (O_172,N_2822,N_2432);
nand UO_173 (O_173,N_2841,N_2871);
xnor UO_174 (O_174,N_2412,N_2993);
or UO_175 (O_175,N_2615,N_2616);
and UO_176 (O_176,N_2607,N_2899);
or UO_177 (O_177,N_2878,N_2571);
nor UO_178 (O_178,N_2792,N_2922);
nor UO_179 (O_179,N_2475,N_2411);
nand UO_180 (O_180,N_2455,N_2974);
nor UO_181 (O_181,N_2544,N_2716);
nand UO_182 (O_182,N_2845,N_2731);
or UO_183 (O_183,N_2956,N_2726);
or UO_184 (O_184,N_2688,N_2969);
and UO_185 (O_185,N_2474,N_2887);
nor UO_186 (O_186,N_2471,N_2524);
nand UO_187 (O_187,N_2443,N_2794);
or UO_188 (O_188,N_2836,N_2558);
or UO_189 (O_189,N_2505,N_2406);
nor UO_190 (O_190,N_2748,N_2865);
nand UO_191 (O_191,N_2606,N_2553);
nor UO_192 (O_192,N_2844,N_2932);
or UO_193 (O_193,N_2912,N_2893);
or UO_194 (O_194,N_2502,N_2652);
or UO_195 (O_195,N_2890,N_2933);
nand UO_196 (O_196,N_2994,N_2611);
or UO_197 (O_197,N_2910,N_2733);
and UO_198 (O_198,N_2781,N_2573);
xor UO_199 (O_199,N_2874,N_2626);
or UO_200 (O_200,N_2828,N_2690);
and UO_201 (O_201,N_2970,N_2637);
nor UO_202 (O_202,N_2767,N_2469);
or UO_203 (O_203,N_2528,N_2450);
nand UO_204 (O_204,N_2725,N_2809);
nand UO_205 (O_205,N_2778,N_2473);
nor UO_206 (O_206,N_2864,N_2774);
and UO_207 (O_207,N_2952,N_2973);
nand UO_208 (O_208,N_2517,N_2674);
nand UO_209 (O_209,N_2595,N_2684);
or UO_210 (O_210,N_2538,N_2928);
nor UO_211 (O_211,N_2789,N_2962);
and UO_212 (O_212,N_2997,N_2675);
and UO_213 (O_213,N_2509,N_2914);
nor UO_214 (O_214,N_2875,N_2983);
or UO_215 (O_215,N_2982,N_2918);
nor UO_216 (O_216,N_2757,N_2984);
nor UO_217 (O_217,N_2512,N_2601);
nor UO_218 (O_218,N_2672,N_2805);
or UO_219 (O_219,N_2554,N_2958);
or UO_220 (O_220,N_2550,N_2633);
nor UO_221 (O_221,N_2570,N_2850);
nand UO_222 (O_222,N_2620,N_2481);
or UO_223 (O_223,N_2929,N_2530);
nand UO_224 (O_224,N_2754,N_2537);
nand UO_225 (O_225,N_2436,N_2468);
nor UO_226 (O_226,N_2776,N_2565);
nor UO_227 (O_227,N_2867,N_2851);
nor UO_228 (O_228,N_2695,N_2796);
and UO_229 (O_229,N_2600,N_2766);
nor UO_230 (O_230,N_2653,N_2863);
or UO_231 (O_231,N_2588,N_2440);
or UO_232 (O_232,N_2807,N_2951);
or UO_233 (O_233,N_2488,N_2712);
or UO_234 (O_234,N_2449,N_2676);
xor UO_235 (O_235,N_2492,N_2493);
and UO_236 (O_236,N_2430,N_2806);
and UO_237 (O_237,N_2427,N_2788);
nor UO_238 (O_238,N_2717,N_2464);
or UO_239 (O_239,N_2539,N_2584);
nor UO_240 (O_240,N_2551,N_2694);
or UO_241 (O_241,N_2656,N_2935);
nand UO_242 (O_242,N_2985,N_2428);
and UO_243 (O_243,N_2884,N_2619);
nand UO_244 (O_244,N_2713,N_2746);
nand UO_245 (O_245,N_2657,N_2700);
nand UO_246 (O_246,N_2667,N_2829);
and UO_247 (O_247,N_2447,N_2605);
or UO_248 (O_248,N_2945,N_2907);
or UO_249 (O_249,N_2433,N_2960);
and UO_250 (O_250,N_2718,N_2610);
nand UO_251 (O_251,N_2439,N_2749);
or UO_252 (O_252,N_2728,N_2682);
or UO_253 (O_253,N_2708,N_2921);
or UO_254 (O_254,N_2448,N_2889);
and UO_255 (O_255,N_2510,N_2503);
and UO_256 (O_256,N_2623,N_2830);
or UO_257 (O_257,N_2987,N_2495);
nand UO_258 (O_258,N_2636,N_2642);
and UO_259 (O_259,N_2500,N_2580);
nand UO_260 (O_260,N_2880,N_2634);
nor UO_261 (O_261,N_2707,N_2422);
nor UO_262 (O_262,N_2791,N_2780);
and UO_263 (O_263,N_2485,N_2693);
and UO_264 (O_264,N_2862,N_2628);
nor UO_265 (O_265,N_2834,N_2915);
nor UO_266 (O_266,N_2482,N_2948);
nand UO_267 (O_267,N_2431,N_2491);
nand UO_268 (O_268,N_2592,N_2868);
nand UO_269 (O_269,N_2968,N_2617);
nand UO_270 (O_270,N_2741,N_2546);
and UO_271 (O_271,N_2519,N_2651);
or UO_272 (O_272,N_2499,N_2696);
or UO_273 (O_273,N_2681,N_2591);
and UO_274 (O_274,N_2472,N_2738);
nand UO_275 (O_275,N_2414,N_2441);
and UO_276 (O_276,N_2487,N_2689);
and UO_277 (O_277,N_2904,N_2504);
nand UO_278 (O_278,N_2856,N_2625);
or UO_279 (O_279,N_2479,N_2572);
xnor UO_280 (O_280,N_2939,N_2419);
or UO_281 (O_281,N_2869,N_2632);
and UO_282 (O_282,N_2446,N_2787);
and UO_283 (O_283,N_2635,N_2701);
or UO_284 (O_284,N_2857,N_2599);
and UO_285 (O_285,N_2560,N_2593);
nor UO_286 (O_286,N_2825,N_2685);
nor UO_287 (O_287,N_2835,N_2821);
nor UO_288 (O_288,N_2687,N_2744);
and UO_289 (O_289,N_2618,N_2846);
nor UO_290 (O_290,N_2739,N_2891);
or UO_291 (O_291,N_2722,N_2454);
or UO_292 (O_292,N_2751,N_2820);
or UO_293 (O_293,N_2630,N_2941);
and UO_294 (O_294,N_2624,N_2784);
and UO_295 (O_295,N_2786,N_2785);
nor UO_296 (O_296,N_2764,N_2686);
and UO_297 (O_297,N_2861,N_2671);
or UO_298 (O_298,N_2598,N_2853);
nand UO_299 (O_299,N_2453,N_2639);
nand UO_300 (O_300,N_2764,N_2729);
nand UO_301 (O_301,N_2757,N_2500);
nand UO_302 (O_302,N_2776,N_2536);
and UO_303 (O_303,N_2625,N_2712);
or UO_304 (O_304,N_2911,N_2681);
nand UO_305 (O_305,N_2608,N_2895);
and UO_306 (O_306,N_2978,N_2599);
nand UO_307 (O_307,N_2676,N_2471);
and UO_308 (O_308,N_2821,N_2415);
and UO_309 (O_309,N_2627,N_2553);
xnor UO_310 (O_310,N_2502,N_2981);
or UO_311 (O_311,N_2615,N_2516);
nand UO_312 (O_312,N_2708,N_2986);
nand UO_313 (O_313,N_2921,N_2794);
nand UO_314 (O_314,N_2707,N_2725);
nand UO_315 (O_315,N_2772,N_2505);
nor UO_316 (O_316,N_2755,N_2430);
and UO_317 (O_317,N_2824,N_2792);
or UO_318 (O_318,N_2494,N_2710);
or UO_319 (O_319,N_2854,N_2736);
or UO_320 (O_320,N_2934,N_2491);
xnor UO_321 (O_321,N_2845,N_2641);
nand UO_322 (O_322,N_2442,N_2703);
or UO_323 (O_323,N_2964,N_2834);
nand UO_324 (O_324,N_2497,N_2549);
nor UO_325 (O_325,N_2429,N_2860);
nand UO_326 (O_326,N_2899,N_2455);
and UO_327 (O_327,N_2416,N_2699);
and UO_328 (O_328,N_2401,N_2907);
or UO_329 (O_329,N_2703,N_2892);
or UO_330 (O_330,N_2934,N_2940);
nor UO_331 (O_331,N_2978,N_2696);
or UO_332 (O_332,N_2529,N_2744);
and UO_333 (O_333,N_2492,N_2424);
nor UO_334 (O_334,N_2827,N_2777);
or UO_335 (O_335,N_2605,N_2755);
or UO_336 (O_336,N_2978,N_2937);
or UO_337 (O_337,N_2547,N_2891);
and UO_338 (O_338,N_2621,N_2885);
or UO_339 (O_339,N_2690,N_2952);
or UO_340 (O_340,N_2789,N_2409);
or UO_341 (O_341,N_2687,N_2435);
or UO_342 (O_342,N_2435,N_2624);
or UO_343 (O_343,N_2771,N_2582);
and UO_344 (O_344,N_2672,N_2437);
or UO_345 (O_345,N_2513,N_2967);
and UO_346 (O_346,N_2837,N_2970);
nand UO_347 (O_347,N_2547,N_2477);
nor UO_348 (O_348,N_2786,N_2550);
xor UO_349 (O_349,N_2640,N_2769);
or UO_350 (O_350,N_2548,N_2630);
nand UO_351 (O_351,N_2455,N_2496);
and UO_352 (O_352,N_2981,N_2988);
nor UO_353 (O_353,N_2717,N_2546);
or UO_354 (O_354,N_2979,N_2885);
and UO_355 (O_355,N_2494,N_2580);
or UO_356 (O_356,N_2574,N_2726);
nor UO_357 (O_357,N_2768,N_2469);
nor UO_358 (O_358,N_2668,N_2437);
or UO_359 (O_359,N_2881,N_2562);
nand UO_360 (O_360,N_2681,N_2461);
and UO_361 (O_361,N_2939,N_2523);
nand UO_362 (O_362,N_2562,N_2768);
nand UO_363 (O_363,N_2923,N_2765);
and UO_364 (O_364,N_2611,N_2519);
nor UO_365 (O_365,N_2931,N_2725);
and UO_366 (O_366,N_2805,N_2744);
and UO_367 (O_367,N_2631,N_2860);
or UO_368 (O_368,N_2580,N_2810);
nand UO_369 (O_369,N_2896,N_2499);
nor UO_370 (O_370,N_2968,N_2425);
and UO_371 (O_371,N_2787,N_2504);
or UO_372 (O_372,N_2720,N_2601);
xor UO_373 (O_373,N_2712,N_2978);
and UO_374 (O_374,N_2771,N_2918);
nor UO_375 (O_375,N_2460,N_2836);
or UO_376 (O_376,N_2514,N_2527);
xor UO_377 (O_377,N_2827,N_2813);
or UO_378 (O_378,N_2686,N_2909);
and UO_379 (O_379,N_2825,N_2523);
nand UO_380 (O_380,N_2755,N_2760);
or UO_381 (O_381,N_2876,N_2555);
and UO_382 (O_382,N_2745,N_2686);
nor UO_383 (O_383,N_2454,N_2904);
and UO_384 (O_384,N_2431,N_2585);
nand UO_385 (O_385,N_2573,N_2673);
and UO_386 (O_386,N_2478,N_2869);
and UO_387 (O_387,N_2647,N_2493);
xnor UO_388 (O_388,N_2924,N_2742);
nand UO_389 (O_389,N_2772,N_2986);
xor UO_390 (O_390,N_2507,N_2718);
nand UO_391 (O_391,N_2513,N_2789);
or UO_392 (O_392,N_2487,N_2905);
nand UO_393 (O_393,N_2518,N_2593);
and UO_394 (O_394,N_2898,N_2587);
nand UO_395 (O_395,N_2580,N_2410);
xnor UO_396 (O_396,N_2938,N_2934);
or UO_397 (O_397,N_2497,N_2474);
nand UO_398 (O_398,N_2646,N_2471);
or UO_399 (O_399,N_2876,N_2917);
and UO_400 (O_400,N_2671,N_2631);
xnor UO_401 (O_401,N_2876,N_2872);
nand UO_402 (O_402,N_2404,N_2569);
nand UO_403 (O_403,N_2528,N_2492);
nand UO_404 (O_404,N_2644,N_2753);
and UO_405 (O_405,N_2610,N_2489);
nor UO_406 (O_406,N_2686,N_2814);
and UO_407 (O_407,N_2634,N_2871);
nand UO_408 (O_408,N_2864,N_2824);
nand UO_409 (O_409,N_2456,N_2540);
and UO_410 (O_410,N_2981,N_2825);
nor UO_411 (O_411,N_2857,N_2487);
nor UO_412 (O_412,N_2902,N_2607);
nor UO_413 (O_413,N_2620,N_2909);
nor UO_414 (O_414,N_2965,N_2938);
nand UO_415 (O_415,N_2717,N_2515);
or UO_416 (O_416,N_2781,N_2512);
nor UO_417 (O_417,N_2782,N_2927);
or UO_418 (O_418,N_2809,N_2426);
or UO_419 (O_419,N_2896,N_2844);
nand UO_420 (O_420,N_2671,N_2879);
nand UO_421 (O_421,N_2703,N_2478);
or UO_422 (O_422,N_2475,N_2482);
nor UO_423 (O_423,N_2968,N_2421);
and UO_424 (O_424,N_2826,N_2691);
and UO_425 (O_425,N_2660,N_2575);
nor UO_426 (O_426,N_2562,N_2567);
nor UO_427 (O_427,N_2971,N_2986);
and UO_428 (O_428,N_2625,N_2722);
and UO_429 (O_429,N_2850,N_2965);
nor UO_430 (O_430,N_2485,N_2890);
or UO_431 (O_431,N_2957,N_2808);
or UO_432 (O_432,N_2464,N_2813);
and UO_433 (O_433,N_2424,N_2822);
and UO_434 (O_434,N_2547,N_2966);
nor UO_435 (O_435,N_2990,N_2609);
or UO_436 (O_436,N_2880,N_2878);
xnor UO_437 (O_437,N_2501,N_2980);
nor UO_438 (O_438,N_2604,N_2446);
or UO_439 (O_439,N_2565,N_2591);
nor UO_440 (O_440,N_2463,N_2783);
or UO_441 (O_441,N_2953,N_2924);
nand UO_442 (O_442,N_2907,N_2792);
xor UO_443 (O_443,N_2898,N_2737);
or UO_444 (O_444,N_2815,N_2698);
nand UO_445 (O_445,N_2607,N_2889);
and UO_446 (O_446,N_2615,N_2506);
and UO_447 (O_447,N_2437,N_2495);
nand UO_448 (O_448,N_2770,N_2848);
nand UO_449 (O_449,N_2410,N_2431);
xor UO_450 (O_450,N_2503,N_2682);
nand UO_451 (O_451,N_2487,N_2555);
nand UO_452 (O_452,N_2820,N_2721);
nand UO_453 (O_453,N_2421,N_2919);
nor UO_454 (O_454,N_2554,N_2486);
nor UO_455 (O_455,N_2628,N_2969);
nand UO_456 (O_456,N_2967,N_2533);
or UO_457 (O_457,N_2775,N_2492);
nand UO_458 (O_458,N_2425,N_2473);
and UO_459 (O_459,N_2954,N_2738);
xor UO_460 (O_460,N_2535,N_2710);
and UO_461 (O_461,N_2653,N_2766);
nand UO_462 (O_462,N_2918,N_2934);
and UO_463 (O_463,N_2730,N_2757);
nand UO_464 (O_464,N_2839,N_2999);
or UO_465 (O_465,N_2599,N_2432);
or UO_466 (O_466,N_2743,N_2994);
or UO_467 (O_467,N_2648,N_2945);
and UO_468 (O_468,N_2595,N_2900);
nand UO_469 (O_469,N_2829,N_2411);
nor UO_470 (O_470,N_2950,N_2918);
xor UO_471 (O_471,N_2805,N_2742);
nand UO_472 (O_472,N_2943,N_2825);
or UO_473 (O_473,N_2599,N_2819);
or UO_474 (O_474,N_2684,N_2982);
nor UO_475 (O_475,N_2810,N_2591);
nor UO_476 (O_476,N_2460,N_2617);
or UO_477 (O_477,N_2479,N_2443);
nand UO_478 (O_478,N_2938,N_2788);
and UO_479 (O_479,N_2724,N_2843);
and UO_480 (O_480,N_2510,N_2463);
nor UO_481 (O_481,N_2597,N_2935);
nor UO_482 (O_482,N_2766,N_2590);
and UO_483 (O_483,N_2494,N_2446);
and UO_484 (O_484,N_2559,N_2810);
and UO_485 (O_485,N_2687,N_2639);
and UO_486 (O_486,N_2526,N_2619);
and UO_487 (O_487,N_2436,N_2719);
nor UO_488 (O_488,N_2568,N_2670);
nand UO_489 (O_489,N_2407,N_2759);
nor UO_490 (O_490,N_2809,N_2646);
and UO_491 (O_491,N_2731,N_2485);
or UO_492 (O_492,N_2487,N_2740);
or UO_493 (O_493,N_2639,N_2540);
nor UO_494 (O_494,N_2543,N_2683);
nand UO_495 (O_495,N_2492,N_2649);
and UO_496 (O_496,N_2422,N_2959);
or UO_497 (O_497,N_2436,N_2737);
nand UO_498 (O_498,N_2694,N_2727);
or UO_499 (O_499,N_2700,N_2640);
endmodule