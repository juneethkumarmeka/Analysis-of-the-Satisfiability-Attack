module basic_3000_30000_3500_5_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_2412,In_2962);
or U1 (N_1,In_1584,In_747);
nand U2 (N_2,In_1270,In_1137);
nand U3 (N_3,In_1365,In_1854);
and U4 (N_4,In_298,In_150);
xnor U5 (N_5,In_1367,In_2475);
nor U6 (N_6,In_62,In_2782);
nand U7 (N_7,In_642,In_997);
and U8 (N_8,In_2035,In_2342);
xnor U9 (N_9,In_1423,In_1363);
xor U10 (N_10,In_2836,In_1296);
xnor U11 (N_11,In_163,In_2586);
xnor U12 (N_12,In_2866,In_1269);
nor U13 (N_13,In_654,In_409);
and U14 (N_14,In_264,In_289);
and U15 (N_15,In_630,In_1736);
xnor U16 (N_16,In_219,In_1657);
nor U17 (N_17,In_2409,In_2476);
nor U18 (N_18,In_937,In_17);
nor U19 (N_19,In_1393,In_1526);
or U20 (N_20,In_435,In_959);
or U21 (N_21,In_1543,In_1847);
or U22 (N_22,In_2200,In_1963);
and U23 (N_23,In_2307,In_2148);
nor U24 (N_24,In_1904,In_1728);
nor U25 (N_25,In_746,In_2313);
nand U26 (N_26,In_2713,In_229);
nand U27 (N_27,In_16,In_2974);
or U28 (N_28,In_479,In_1790);
and U29 (N_29,In_1630,In_2523);
and U30 (N_30,In_2769,In_784);
nor U31 (N_31,In_2583,In_1710);
xnor U32 (N_32,In_240,In_831);
or U33 (N_33,In_1848,In_2244);
nor U34 (N_34,In_1595,In_582);
xor U35 (N_35,In_100,In_556);
xnor U36 (N_36,In_1714,In_2139);
or U37 (N_37,In_2529,In_1748);
or U38 (N_38,In_1538,In_879);
and U39 (N_39,In_1061,In_647);
or U40 (N_40,In_2908,In_2504);
or U41 (N_41,In_2846,In_1077);
nor U42 (N_42,In_2755,In_2210);
nand U43 (N_43,In_1693,In_2125);
and U44 (N_44,In_34,In_680);
nor U45 (N_45,In_611,In_2262);
and U46 (N_46,In_2803,In_2317);
nand U47 (N_47,In_759,In_659);
nand U48 (N_48,In_1274,In_797);
xnor U49 (N_49,In_893,In_1784);
nand U50 (N_50,In_819,In_2135);
or U51 (N_51,In_201,In_512);
and U52 (N_52,In_550,In_2001);
or U53 (N_53,In_2033,In_449);
or U54 (N_54,In_473,In_2233);
nand U55 (N_55,In_2043,In_1919);
nand U56 (N_56,In_1913,In_664);
xor U57 (N_57,In_314,In_522);
nor U58 (N_58,In_2059,In_596);
xor U59 (N_59,In_1647,In_554);
nand U60 (N_60,In_1525,In_2902);
or U61 (N_61,In_2424,In_606);
nor U62 (N_62,In_2518,In_941);
nand U63 (N_63,In_1263,In_2889);
nand U64 (N_64,In_1221,In_1444);
or U65 (N_65,In_603,In_1148);
nor U66 (N_66,In_711,In_2253);
or U67 (N_67,In_2270,In_2015);
and U68 (N_68,In_2153,In_1315);
nor U69 (N_69,In_1495,In_2410);
or U70 (N_70,In_368,In_251);
and U71 (N_71,In_2344,In_350);
nor U72 (N_72,In_2876,In_1976);
nand U73 (N_73,In_1473,In_1516);
nor U74 (N_74,In_2407,In_1433);
or U75 (N_75,In_48,In_978);
nor U76 (N_76,In_622,In_261);
nor U77 (N_77,In_962,In_826);
nor U78 (N_78,In_1889,In_425);
nand U79 (N_79,In_1011,In_2380);
and U80 (N_80,In_1399,In_2141);
and U81 (N_81,In_2415,In_297);
xnor U82 (N_82,In_249,In_1929);
nor U83 (N_83,In_1534,In_1503);
xnor U84 (N_84,In_2184,In_2347);
or U85 (N_85,In_468,In_1129);
and U86 (N_86,In_2396,In_45);
or U87 (N_87,In_1414,In_644);
and U88 (N_88,In_2392,In_2705);
xor U89 (N_89,In_1028,In_2609);
or U90 (N_90,In_5,In_2459);
nand U91 (N_91,In_1350,In_246);
nand U92 (N_92,In_1022,In_77);
and U93 (N_93,In_1089,In_2165);
xor U94 (N_94,In_2708,In_87);
nand U95 (N_95,In_2134,In_2500);
nand U96 (N_96,In_520,In_818);
nand U97 (N_97,In_95,In_2677);
or U98 (N_98,In_28,In_528);
and U99 (N_99,In_840,In_1793);
nor U100 (N_100,In_1067,In_1469);
xnor U101 (N_101,In_263,In_1877);
nor U102 (N_102,In_1537,In_2478);
nor U103 (N_103,In_151,In_2463);
nand U104 (N_104,In_2764,In_652);
and U105 (N_105,In_2095,In_1771);
or U106 (N_106,In_599,In_33);
or U107 (N_107,In_996,In_2056);
nand U108 (N_108,In_2002,In_2867);
nor U109 (N_109,In_1260,In_1500);
nand U110 (N_110,In_417,In_2368);
xnor U111 (N_111,In_2601,In_2023);
and U112 (N_112,In_1696,In_2800);
nor U113 (N_113,In_2497,In_1573);
and U114 (N_114,In_542,In_1004);
or U115 (N_115,In_1236,In_106);
nor U116 (N_116,In_552,In_1582);
nand U117 (N_117,In_1151,In_1716);
nor U118 (N_118,In_2144,In_2488);
or U119 (N_119,In_1039,In_2711);
or U120 (N_120,In_2413,In_1391);
nor U121 (N_121,In_1862,In_2492);
nand U122 (N_122,In_593,In_531);
or U123 (N_123,In_1897,In_1914);
nand U124 (N_124,In_523,In_299);
nand U125 (N_125,In_1967,In_2498);
nor U126 (N_126,In_1997,In_2838);
and U127 (N_127,In_916,In_156);
and U128 (N_128,In_1762,In_1344);
nor U129 (N_129,In_846,In_85);
and U130 (N_130,In_1819,In_384);
nand U131 (N_131,In_159,In_1141);
and U132 (N_132,In_252,In_811);
nor U133 (N_133,In_269,In_2272);
or U134 (N_134,In_2738,In_353);
and U135 (N_135,In_82,In_336);
nand U136 (N_136,In_2528,In_2024);
or U137 (N_137,In_568,In_1596);
nor U138 (N_138,In_2054,In_1353);
nor U139 (N_139,In_2473,In_2771);
or U140 (N_140,In_1203,In_2398);
nand U141 (N_141,In_963,In_2108);
and U142 (N_142,In_2248,In_381);
nor U143 (N_143,In_2110,In_1464);
or U144 (N_144,In_2919,In_2978);
or U145 (N_145,In_2823,In_1139);
nand U146 (N_146,In_2762,In_2801);
and U147 (N_147,In_2798,In_2460);
xnor U148 (N_148,In_2188,In_2997);
xor U149 (N_149,In_1899,In_2532);
nor U150 (N_150,In_1551,In_2615);
xor U151 (N_151,In_567,In_312);
or U152 (N_152,In_2552,In_2625);
nor U153 (N_153,In_1686,In_2802);
nand U154 (N_154,In_2915,In_1618);
nand U155 (N_155,In_1978,In_406);
nand U156 (N_156,In_1799,In_1825);
nor U157 (N_157,In_2282,In_1163);
nand U158 (N_158,In_1428,In_977);
or U159 (N_159,In_1901,In_2290);
nor U160 (N_160,In_2495,In_905);
and U161 (N_161,In_2223,In_86);
nand U162 (N_162,In_1189,In_1430);
or U163 (N_163,In_2589,In_2926);
nor U164 (N_164,In_632,In_259);
xnor U165 (N_165,In_634,In_827);
nor U166 (N_166,In_355,In_1776);
xor U167 (N_167,In_2855,In_1304);
or U168 (N_168,In_2303,In_1785);
or U169 (N_169,In_2780,In_152);
nor U170 (N_170,In_1333,In_370);
nand U171 (N_171,In_1542,In_1337);
and U172 (N_172,In_2701,In_2694);
and U173 (N_173,In_660,In_1082);
xnor U174 (N_174,In_56,In_2390);
and U175 (N_175,In_2297,In_1772);
and U176 (N_176,In_641,In_1222);
nand U177 (N_177,In_576,In_1217);
xor U178 (N_178,In_2903,In_843);
xnor U179 (N_179,In_1727,In_391);
and U180 (N_180,In_105,In_1896);
nor U181 (N_181,In_421,In_608);
nor U182 (N_182,In_2496,In_1589);
nor U183 (N_183,In_170,In_825);
nand U184 (N_184,In_1588,In_272);
nand U185 (N_185,In_591,In_663);
or U186 (N_186,In_1427,In_1070);
nand U187 (N_187,In_1317,In_572);
or U188 (N_188,In_123,In_1741);
and U189 (N_189,In_2740,In_1559);
or U190 (N_190,In_999,In_2287);
nor U191 (N_191,In_2316,In_2101);
and U192 (N_192,In_1988,In_861);
xnor U193 (N_193,In_967,In_2227);
nor U194 (N_194,In_196,In_2852);
and U195 (N_195,In_1770,In_292);
xor U196 (N_196,In_1611,In_975);
and U197 (N_197,In_53,In_1462);
and U198 (N_198,In_906,In_1900);
and U199 (N_199,In_2382,In_2880);
xor U200 (N_200,In_752,In_2587);
or U201 (N_201,In_2292,In_964);
nand U202 (N_202,In_2952,In_378);
and U203 (N_203,In_2183,In_847);
or U204 (N_204,In_1628,In_571);
nand U205 (N_205,In_2222,In_2482);
nand U206 (N_206,In_1112,In_548);
and U207 (N_207,In_2779,In_1868);
nand U208 (N_208,In_1321,In_2097);
and U209 (N_209,In_2543,In_2123);
or U210 (N_210,In_2825,In_2517);
or U211 (N_211,In_1658,In_358);
or U212 (N_212,In_867,In_1697);
nor U213 (N_213,In_1049,In_808);
nand U214 (N_214,In_2197,In_1147);
or U215 (N_215,In_2696,In_2616);
xor U216 (N_216,In_2774,In_2891);
and U217 (N_217,In_404,In_1612);
nand U218 (N_218,In_594,In_1016);
nor U219 (N_219,In_1177,In_1577);
nor U220 (N_220,In_2428,In_1403);
nand U221 (N_221,In_1051,In_1198);
nand U222 (N_222,In_688,In_237);
or U223 (N_223,In_2387,In_2850);
and U224 (N_224,In_1272,In_1104);
nand U225 (N_225,In_2343,In_2076);
nand U226 (N_226,In_2987,In_411);
and U227 (N_227,In_2449,In_738);
nor U228 (N_228,In_1838,In_1472);
or U229 (N_229,In_1431,In_1152);
nand U230 (N_230,In_1835,In_318);
and U231 (N_231,In_2323,In_2910);
or U232 (N_232,In_1911,In_1401);
and U233 (N_233,In_841,In_2220);
or U234 (N_234,In_2806,In_2191);
xnor U235 (N_235,In_1328,In_418);
nor U236 (N_236,In_1247,In_770);
or U237 (N_237,In_439,In_1283);
or U238 (N_238,In_1927,In_181);
or U239 (N_239,In_1458,In_2685);
and U240 (N_240,In_852,In_1338);
nand U241 (N_241,In_557,In_2775);
or U242 (N_242,In_2074,In_521);
nor U243 (N_243,In_646,In_2457);
nor U244 (N_244,In_1801,In_2048);
nand U245 (N_245,In_1873,In_2558);
nor U246 (N_246,In_1759,In_1088);
nand U247 (N_247,In_986,In_2005);
nand U248 (N_248,In_1368,In_869);
xor U249 (N_249,In_1757,In_1340);
xor U250 (N_250,In_444,In_416);
or U251 (N_251,In_1223,In_842);
or U252 (N_252,In_1621,In_1497);
and U253 (N_253,In_2758,In_2374);
and U254 (N_254,In_1306,In_904);
nand U255 (N_255,In_293,In_1432);
nand U256 (N_256,In_1634,In_796);
xor U257 (N_257,In_2028,In_442);
nor U258 (N_258,In_683,In_2393);
nor U259 (N_259,In_1673,In_2541);
or U260 (N_260,In_720,In_1753);
and U261 (N_261,In_2691,In_1782);
nor U262 (N_262,In_29,In_2301);
nor U263 (N_263,In_1761,In_483);
nand U264 (N_264,In_2397,In_2888);
or U265 (N_265,In_58,In_114);
nand U266 (N_266,In_2814,In_195);
or U267 (N_267,In_2358,In_1360);
xor U268 (N_268,In_450,In_2238);
nand U269 (N_269,In_2958,In_2405);
and U270 (N_270,In_2075,In_1097);
and U271 (N_271,In_2673,In_2267);
xnor U272 (N_272,In_2314,In_509);
nor U273 (N_273,In_1982,In_1859);
nor U274 (N_274,In_2717,In_2266);
nor U275 (N_275,In_98,In_1406);
nand U276 (N_276,In_1098,In_1455);
or U277 (N_277,In_2026,In_2534);
nand U278 (N_278,In_262,In_1265);
nand U279 (N_279,In_1064,In_1898);
nand U280 (N_280,In_2688,In_1685);
or U281 (N_281,In_1320,In_2168);
or U282 (N_282,In_426,In_280);
and U283 (N_283,In_396,In_2752);
or U284 (N_284,In_2635,In_1912);
nand U285 (N_285,In_737,In_1530);
nand U286 (N_286,In_2111,In_706);
xor U287 (N_287,In_1169,In_1470);
nand U288 (N_288,In_2471,In_1950);
and U289 (N_289,In_1522,In_2280);
nand U290 (N_290,In_1324,In_1438);
or U291 (N_291,In_2166,In_1851);
and U292 (N_292,In_2564,In_1974);
or U293 (N_293,In_1124,In_2723);
nand U294 (N_294,In_2832,In_535);
or U295 (N_295,In_726,In_1521);
or U296 (N_296,In_1035,In_1593);
nor U297 (N_297,In_2115,In_727);
xor U298 (N_298,In_1273,In_97);
nand U299 (N_299,In_146,In_193);
or U300 (N_300,In_856,In_2324);
and U301 (N_301,In_2450,In_431);
nand U302 (N_302,In_2025,In_1499);
nand U303 (N_303,In_2960,In_1200);
nor U304 (N_304,In_171,In_376);
nand U305 (N_305,In_1303,In_2536);
or U306 (N_306,In_2647,In_241);
and U307 (N_307,In_2418,In_2605);
nand U308 (N_308,In_774,In_2379);
nand U309 (N_309,In_1763,In_2785);
nor U310 (N_310,In_2560,In_741);
nand U311 (N_311,In_2931,In_1695);
nor U312 (N_312,In_661,In_2051);
and U313 (N_313,In_682,In_886);
or U314 (N_314,In_1990,In_1535);
and U315 (N_315,In_2864,In_2268);
xor U316 (N_316,In_2240,In_2044);
or U317 (N_317,In_2922,In_1740);
and U318 (N_318,In_1606,In_1711);
nor U319 (N_319,In_2310,In_2467);
and U320 (N_320,In_2009,In_1533);
nand U321 (N_321,In_71,In_2817);
and U322 (N_322,In_2863,In_666);
nand U323 (N_323,In_143,In_2660);
xnor U324 (N_324,In_1466,In_2055);
nor U325 (N_325,In_2665,In_1562);
nand U326 (N_326,In_390,In_681);
xor U327 (N_327,In_438,In_69);
nor U328 (N_328,In_2008,In_573);
nor U329 (N_329,In_422,In_1188);
or U330 (N_330,In_1867,In_2841);
and U331 (N_331,In_2563,In_402);
or U332 (N_332,In_1185,In_223);
and U333 (N_333,In_2377,In_534);
nor U334 (N_334,In_352,In_2225);
and U335 (N_335,In_2699,In_1511);
nor U336 (N_336,In_1482,In_1150);
nor U337 (N_337,In_853,In_133);
or U338 (N_338,In_2352,In_408);
and U339 (N_339,In_2736,In_1342);
or U340 (N_340,In_625,In_742);
nand U341 (N_341,In_2527,In_2716);
nor U342 (N_342,In_1923,In_2146);
or U343 (N_343,In_1308,In_779);
nand U344 (N_344,In_1992,In_2204);
nor U345 (N_345,In_109,In_1758);
nand U346 (N_346,In_1479,In_1378);
nand U347 (N_347,In_1037,In_961);
nand U348 (N_348,In_1441,In_2251);
xnor U349 (N_349,In_533,In_810);
nor U350 (N_350,In_1021,In_1837);
nor U351 (N_351,In_751,In_2901);
xor U352 (N_352,In_2162,In_2524);
and U353 (N_353,In_1578,In_216);
or U354 (N_354,In_1703,In_1166);
nand U355 (N_355,In_1831,In_1845);
and U356 (N_356,In_864,In_1883);
xnor U357 (N_357,In_530,In_870);
nor U358 (N_358,In_2972,In_2670);
and U359 (N_359,In_1517,In_1347);
or U360 (N_360,In_1048,In_1820);
or U361 (N_361,In_2087,In_2444);
and U362 (N_362,In_2892,In_2422);
or U363 (N_363,In_627,In_1465);
and U364 (N_364,In_61,In_1172);
nor U365 (N_365,In_1631,In_2417);
nor U366 (N_366,In_1174,In_1531);
and U367 (N_367,In_2603,In_2751);
nand U368 (N_368,In_1952,In_1078);
nor U369 (N_369,In_1398,In_954);
nand U370 (N_370,In_2329,In_1069);
nor U371 (N_371,In_2917,In_1407);
and U372 (N_372,In_457,In_2084);
nor U373 (N_373,In_175,In_1953);
or U374 (N_374,In_1386,In_1092);
or U375 (N_375,In_1192,In_2215);
or U376 (N_376,In_1824,In_2425);
or U377 (N_377,In_281,In_1817);
and U378 (N_378,In_1213,In_942);
or U379 (N_379,In_2363,In_822);
or U380 (N_380,In_344,In_1767);
and U381 (N_381,In_1181,In_1038);
xnor U382 (N_382,In_993,In_119);
nand U383 (N_383,In_2870,In_2928);
or U384 (N_384,In_605,In_2137);
nor U385 (N_385,In_2787,In_1481);
nand U386 (N_386,In_2038,In_515);
or U387 (N_387,In_423,In_2720);
and U388 (N_388,In_885,In_1445);
nor U389 (N_389,In_1519,In_2799);
nand U390 (N_390,In_2693,In_2429);
nand U391 (N_391,In_2192,In_2650);
nand U392 (N_392,In_2907,In_2333);
and U393 (N_393,In_2474,In_331);
and U394 (N_394,In_2066,In_676);
and U395 (N_395,In_1865,In_712);
and U396 (N_396,In_2707,In_324);
nor U397 (N_397,In_1044,In_2201);
or U398 (N_398,In_320,In_1170);
or U399 (N_399,In_1332,In_2017);
or U400 (N_400,In_969,In_341);
xnor U401 (N_401,In_2768,In_2298);
and U402 (N_402,In_2871,In_1384);
or U403 (N_403,In_1193,In_1677);
nor U404 (N_404,In_769,In_474);
nand U405 (N_405,In_1640,In_1604);
nand U406 (N_406,In_990,In_2419);
nor U407 (N_407,In_1327,In_1938);
or U408 (N_408,In_43,In_1626);
and U409 (N_409,In_428,In_1843);
or U410 (N_410,In_1764,In_2989);
or U411 (N_411,In_165,In_2172);
or U412 (N_412,In_600,In_2856);
nor U413 (N_413,In_2721,In_707);
xnor U414 (N_414,In_813,In_311);
nor U415 (N_415,In_140,In_366);
nand U416 (N_416,In_913,In_2875);
and U417 (N_417,In_2218,In_1449);
nand U418 (N_418,In_173,In_874);
and U419 (N_419,In_2232,In_1587);
nand U420 (N_420,In_1777,In_777);
and U421 (N_421,In_2209,In_499);
nor U422 (N_422,In_2672,In_1295);
and U423 (N_423,In_1749,In_2283);
nor U424 (N_424,In_2975,In_2834);
nand U425 (N_425,In_1943,In_372);
nor U426 (N_426,In_2029,In_2991);
nor U427 (N_427,In_168,In_1760);
or U428 (N_428,In_854,In_2837);
or U429 (N_429,In_651,In_1940);
nand U430 (N_430,In_2535,In_1167);
nand U431 (N_431,In_2509,In_1581);
nand U432 (N_432,In_549,In_807);
nand U433 (N_433,In_1625,In_136);
nor U434 (N_434,In_2439,In_945);
and U435 (N_435,In_1539,In_92);
xor U436 (N_436,In_2895,In_2468);
and U437 (N_437,In_351,In_2749);
nand U438 (N_438,In_598,In_21);
nor U439 (N_439,In_2100,In_2948);
nor U440 (N_440,In_898,In_1488);
and U441 (N_441,In_273,In_2120);
nor U442 (N_442,In_805,In_958);
nand U443 (N_443,In_1597,In_2851);
and U444 (N_444,In_2264,In_7);
nand U445 (N_445,In_1318,In_461);
and U446 (N_446,In_2531,In_1258);
nand U447 (N_447,In_1833,In_13);
or U448 (N_448,In_1370,In_2753);
or U449 (N_449,In_702,In_487);
nand U450 (N_450,In_364,In_1394);
xnor U451 (N_451,In_1291,In_2942);
nor U452 (N_452,In_1352,In_2639);
nor U453 (N_453,In_1507,In_2568);
xor U454 (N_454,In_257,In_51);
nand U455 (N_455,In_2763,In_1564);
xor U456 (N_456,In_1805,In_83);
nand U457 (N_457,In_1781,In_296);
nor U458 (N_458,In_675,In_2150);
or U459 (N_459,In_1373,In_112);
or U460 (N_460,In_2132,In_2858);
nor U461 (N_461,In_1955,In_2039);
and U462 (N_462,In_1168,In_317);
and U463 (N_463,In_2127,In_212);
nor U464 (N_464,In_2430,In_427);
or U465 (N_465,In_1683,In_239);
nand U466 (N_466,In_2149,In_2530);
and U467 (N_467,In_1815,In_2058);
and U468 (N_468,In_2164,In_1461);
or U469 (N_469,In_2260,In_546);
or U470 (N_470,In_1074,In_2619);
nand U471 (N_471,In_1251,In_668);
or U472 (N_472,In_2868,In_1880);
nand U473 (N_473,In_346,In_430);
nand U474 (N_474,In_519,In_1655);
and U475 (N_475,In_302,In_1920);
nor U476 (N_476,In_2163,In_2304);
and U477 (N_477,In_2448,In_1572);
and U478 (N_478,In_1860,In_1857);
nand U479 (N_479,In_2747,In_1766);
or U480 (N_480,In_1671,In_699);
xor U481 (N_481,In_1842,In_2542);
xnor U482 (N_482,In_649,In_23);
or U483 (N_483,In_2041,In_1257);
nor U484 (N_484,In_2052,In_127);
xnor U485 (N_485,In_2250,In_1108);
xnor U486 (N_486,In_2385,In_708);
and U487 (N_487,In_2746,In_2886);
or U488 (N_488,In_776,In_2353);
and U489 (N_489,In_2367,In_1812);
xor U490 (N_490,In_1161,In_2982);
nor U491 (N_491,In_529,In_1754);
xor U492 (N_492,In_2581,In_859);
and U493 (N_493,In_743,In_876);
nand U494 (N_494,In_700,In_1422);
and U495 (N_495,In_984,In_79);
xnor U496 (N_496,In_1629,In_1238);
and U497 (N_497,In_2435,In_2899);
nor U498 (N_498,In_1882,In_1909);
and U499 (N_499,In_980,In_2570);
or U500 (N_500,In_66,In_1709);
and U501 (N_501,In_817,In_1620);
and U502 (N_502,In_2442,In_2477);
nor U503 (N_503,In_1520,In_2641);
or U504 (N_504,In_1649,In_2666);
and U505 (N_505,In_543,In_2273);
nor U506 (N_506,In_745,In_1316);
and U507 (N_507,In_2933,In_2332);
nor U508 (N_508,In_1447,In_1334);
and U509 (N_509,In_721,In_2649);
and U510 (N_510,In_1680,In_2849);
or U511 (N_511,In_1459,In_373);
nor U512 (N_512,In_1404,In_2845);
nand U513 (N_513,In_2890,In_2219);
xnor U514 (N_514,In_1734,In_1576);
nor U515 (N_515,In_1856,In_74);
or U516 (N_516,In_517,In_2582);
nor U517 (N_517,In_1411,In_2019);
or U518 (N_518,In_210,In_857);
and U519 (N_519,In_1925,In_1025);
nor U520 (N_520,In_1326,In_478);
or U521 (N_521,In_2462,In_1349);
or U522 (N_522,In_2626,In_386);
or U523 (N_523,In_1580,In_2395);
or U524 (N_524,In_383,In_360);
nor U525 (N_525,In_2932,In_773);
xnor U526 (N_526,In_1162,In_764);
or U527 (N_527,In_918,In_2548);
or U528 (N_528,In_653,In_881);
and U529 (N_529,In_2617,In_2546);
nor U530 (N_530,In_2810,In_678);
and U531 (N_531,In_224,In_903);
or U532 (N_532,In_1288,In_2556);
nor U533 (N_533,In_710,In_1385);
nor U534 (N_534,In_382,In_1259);
or U535 (N_535,In_672,In_2179);
or U536 (N_536,In_2735,In_198);
nand U537 (N_537,In_1550,In_1371);
and U538 (N_538,In_875,In_326);
and U539 (N_539,In_1730,In_1962);
and U540 (N_540,In_2512,In_388);
and U541 (N_541,In_1096,In_399);
and U542 (N_542,In_1972,In_279);
nand U543 (N_543,In_658,In_141);
and U544 (N_544,In_1586,In_126);
nor U545 (N_545,In_1656,In_832);
or U546 (N_546,In_1298,In_1547);
nor U547 (N_547,In_1669,In_2373);
nor U548 (N_548,In_2391,In_956);
or U549 (N_549,In_9,In_1600);
or U550 (N_550,In_1506,In_514);
and U551 (N_551,In_491,In_6);
and U552 (N_552,In_2585,In_380);
nor U553 (N_553,In_778,In_1229);
nor U554 (N_554,In_2483,In_120);
nand U555 (N_555,In_436,In_1592);
xor U556 (N_556,In_2571,In_2403);
and U557 (N_557,In_332,In_90);
or U558 (N_558,In_2760,In_2965);
nor U559 (N_559,In_2037,In_690);
nor U560 (N_560,In_1540,In_621);
xnor U561 (N_561,In_816,In_1609);
xnor U562 (N_562,In_2678,In_951);
nand U563 (N_563,In_2383,In_182);
or U564 (N_564,In_361,In_466);
nand U565 (N_565,In_617,In_750);
and U566 (N_566,In_1248,In_489);
or U567 (N_567,In_2129,In_72);
or U568 (N_568,In_2401,In_403);
nand U569 (N_569,In_2697,In_54);
and U570 (N_570,In_2784,In_2274);
or U571 (N_571,In_1878,In_1807);
and U572 (N_572,In_1692,In_2594);
and U573 (N_573,In_441,In_1816);
and U574 (N_574,In_192,In_493);
and U575 (N_575,In_2466,In_938);
or U576 (N_576,In_736,In_2487);
nor U577 (N_577,In_2645,In_1250);
nor U578 (N_578,In_145,In_1999);
or U579 (N_579,In_1099,In_2362);
and U580 (N_580,In_793,In_695);
and U581 (N_581,In_2447,In_844);
or U582 (N_582,In_1871,In_2388);
nor U583 (N_583,In_2211,In_1388);
xnor U584 (N_584,In_1651,In_991);
nand U585 (N_585,In_2724,In_1814);
nor U586 (N_586,In_2511,In_1);
and U587 (N_587,In_767,In_481);
xor U588 (N_588,In_1959,In_2319);
and U589 (N_589,In_367,In_2376);
nand U590 (N_590,In_1494,In_2657);
and U591 (N_591,In_130,In_1619);
nor U592 (N_592,In_1164,In_2472);
and U593 (N_593,In_2205,In_1267);
nand U594 (N_594,In_2239,In_2652);
nor U595 (N_595,In_1617,In_1951);
or U596 (N_596,In_587,In_1063);
or U597 (N_597,In_2078,In_2203);
nand U598 (N_598,In_2016,In_2731);
nor U599 (N_599,In_1268,In_410);
nor U600 (N_600,In_979,In_2207);
and U601 (N_601,In_983,In_2992);
nor U602 (N_602,In_2370,In_134);
or U603 (N_603,In_2638,In_282);
and U604 (N_604,In_2453,In_218);
or U605 (N_605,In_2194,In_615);
and U606 (N_606,In_1788,In_1235);
or U607 (N_607,In_508,In_290);
nand U608 (N_608,In_375,In_1452);
or U609 (N_609,In_2860,In_2328);
and U610 (N_610,In_2426,In_1888);
or U611 (N_611,In_2829,In_1977);
and U612 (N_612,In_1661,In_30);
or U613 (N_613,In_677,In_1961);
nor U614 (N_614,In_1713,In_2633);
nand U615 (N_615,In_1093,In_1712);
xnor U616 (N_616,In_771,In_1701);
xor U617 (N_617,In_319,In_1195);
and U618 (N_618,In_1775,In_2826);
or U619 (N_619,In_460,In_1058);
nand U620 (N_620,In_2706,In_694);
xor U621 (N_621,In_944,In_1515);
and U622 (N_622,In_872,In_1145);
nand U623 (N_623,In_1726,In_496);
or U624 (N_624,In_884,In_801);
nor U625 (N_625,In_2254,In_2230);
nor U626 (N_626,In_1644,In_227);
and U627 (N_627,In_1241,In_1389);
nor U628 (N_628,In_1830,In_305);
nand U629 (N_629,In_1751,In_949);
and U630 (N_630,In_862,In_982);
or U631 (N_631,In_2947,In_2011);
or U632 (N_632,In_2072,In_965);
nand U633 (N_633,In_2874,In_640);
and U634 (N_634,In_202,In_2335);
xnor U635 (N_635,In_2510,In_64);
nor U636 (N_636,In_19,In_1369);
and U637 (N_637,In_1153,In_1623);
or U638 (N_638,In_1107,In_8);
nor U639 (N_639,In_1142,In_52);
nor U640 (N_640,In_463,In_1355);
nor U641 (N_641,In_2683,In_2339);
and U642 (N_642,In_1983,In_586);
nor U643 (N_643,In_2815,In_327);
xor U644 (N_644,In_716,In_936);
nor U645 (N_645,In_2446,In_2984);
xnor U646 (N_646,In_1264,In_1379);
nor U647 (N_647,In_2246,In_2461);
nand U648 (N_648,In_2357,In_2940);
nand U649 (N_649,In_1690,In_2351);
xnor U650 (N_650,In_972,In_2632);
or U651 (N_651,In_149,In_2853);
nor U652 (N_652,In_2573,In_824);
xor U653 (N_653,In_111,In_1942);
or U654 (N_654,In_1906,In_1555);
or U655 (N_655,In_1638,In_2664);
xnor U656 (N_656,In_729,In_1056);
nand U657 (N_657,In_2526,In_1822);
and U658 (N_658,In_2096,In_2004);
nor U659 (N_659,In_2356,In_337);
or U660 (N_660,In_768,In_2255);
or U661 (N_661,In_1382,In_245);
nor U662 (N_662,In_635,In_1239);
nand U663 (N_663,In_2956,In_1616);
and U664 (N_664,In_1993,In_693);
xor U665 (N_665,In_1756,In_1182);
and U666 (N_666,In_135,In_907);
nand U667 (N_667,In_2783,In_446);
or U668 (N_668,In_766,In_1276);
nand U669 (N_669,In_1202,In_2896);
nand U670 (N_670,In_1682,In_1297);
and U671 (N_671,In_2767,In_2325);
or U672 (N_672,In_933,In_1738);
or U673 (N_673,In_704,In_2174);
or U674 (N_674,In_2451,In_1558);
and U675 (N_675,In_1797,In_1841);
nor U676 (N_676,In_2702,In_1737);
or U677 (N_677,In_2226,In_2082);
or U678 (N_678,In_1226,In_99);
or U679 (N_679,In_714,In_756);
nor U680 (N_680,In_486,In_155);
nand U681 (N_681,In_2176,In_1287);
and U682 (N_682,In_1986,In_2216);
nand U683 (N_683,In_1874,In_2369);
nor U684 (N_684,In_50,In_2263);
and U685 (N_685,In_2117,In_2659);
nor U686 (N_686,In_2464,In_2883);
and U687 (N_687,In_1636,In_2602);
xor U688 (N_688,In_1157,In_1305);
nor U689 (N_689,In_1158,In_1855);
or U690 (N_690,In_2480,In_1918);
nand U691 (N_691,In_1413,In_2923);
nor U692 (N_692,In_2946,In_2680);
or U693 (N_693,In_1454,In_2077);
nand U694 (N_694,In_323,In_1599);
or U695 (N_695,In_1210,In_2490);
nand U696 (N_696,In_2465,In_792);
and U697 (N_697,In_220,In_1448);
or U698 (N_698,In_2913,In_2550);
or U699 (N_699,In_2709,In_2621);
or U700 (N_700,In_798,In_1523);
nor U701 (N_701,In_1633,In_1007);
and U702 (N_702,In_2350,In_2190);
nor U703 (N_703,In_2271,In_2805);
xnor U704 (N_704,In_1122,In_762);
nand U705 (N_705,In_1010,In_2545);
and U706 (N_706,In_1341,In_1645);
nor U707 (N_707,In_2961,In_84);
or U708 (N_708,In_1040,In_901);
nor U709 (N_709,In_2224,In_1417);
nor U710 (N_710,In_2142,In_189);
and U711 (N_711,In_1800,In_2692);
nor U712 (N_712,In_283,In_1780);
or U713 (N_713,In_2790,In_131);
nor U714 (N_714,In_2712,In_2627);
nor U715 (N_715,In_559,In_2791);
or U716 (N_716,In_345,In_2613);
and U717 (N_717,In_734,In_1425);
xor U718 (N_718,In_1498,In_765);
or U719 (N_719,In_829,In_1421);
nor U720 (N_720,In_2734,In_234);
nand U721 (N_721,In_2489,In_1729);
or U722 (N_722,In_288,In_1944);
or U723 (N_723,In_2640,In_1585);
xnor U724 (N_724,In_484,In_863);
nand U725 (N_725,In_2818,In_2929);
and U726 (N_726,In_2154,In_920);
and U727 (N_727,In_37,In_948);
nor U728 (N_728,In_705,In_685);
and U729 (N_729,In_1310,In_1556);
or U730 (N_730,In_2909,In_2765);
and U731 (N_731,In_1262,In_40);
nor U732 (N_732,In_2656,In_185);
and U733 (N_733,In_1934,In_2985);
or U734 (N_734,In_2018,In_1665);
nor U735 (N_735,In_1255,In_462);
nand U736 (N_736,In_2807,In_2745);
nor U737 (N_737,In_2136,In_2327);
or U738 (N_738,In_2642,In_1424);
nand U739 (N_739,In_1654,In_2916);
nand U740 (N_740,In_2995,In_2265);
nor U741 (N_741,In_1408,In_725);
and U742 (N_742,In_1380,In_2399);
nor U743 (N_743,In_1437,In_1663);
and U744 (N_744,In_834,In_2359);
and U745 (N_745,In_233,In_2859);
nor U746 (N_746,In_2857,In_41);
nor U747 (N_747,In_1362,In_2436);
nand U748 (N_748,In_1397,In_723);
nand U749 (N_749,In_2557,In_2228);
nor U750 (N_750,In_1375,In_618);
or U751 (N_751,In_349,In_1325);
and U752 (N_752,In_2334,In_851);
nand U753 (N_753,In_1121,In_2572);
or U754 (N_754,In_1916,In_719);
xnor U755 (N_755,In_614,In_174);
nand U756 (N_756,In_1227,In_1935);
xor U757 (N_757,In_256,In_1561);
and U758 (N_758,In_2067,In_1571);
nor U759 (N_759,In_1966,In_2257);
nor U760 (N_760,In_637,In_57);
and U761 (N_761,In_482,In_2979);
or U762 (N_762,In_786,In_1662);
nand U763 (N_763,In_1605,In_1109);
or U764 (N_764,In_2157,In_1949);
nor U765 (N_765,In_2578,In_1314);
or U766 (N_766,In_1405,In_501);
and U767 (N_767,In_648,In_1778);
and U768 (N_768,In_1354,In_1718);
and U769 (N_769,In_799,In_2539);
or U770 (N_770,In_923,In_1917);
nor U771 (N_771,In_2715,In_2113);
nand U772 (N_772,In_1343,In_362);
nand U773 (N_773,In_347,In_1228);
and U774 (N_774,In_1708,In_2469);
or U775 (N_775,In_67,In_242);
or U776 (N_776,In_2414,In_643);
nand U777 (N_777,In_1960,In_122);
and U778 (N_778,In_1244,In_2293);
or U779 (N_779,In_2241,In_492);
and U780 (N_780,In_2634,In_740);
nand U781 (N_781,In_2516,In_2898);
or U782 (N_782,In_294,In_267);
nand U783 (N_783,In_1957,In_2728);
and U784 (N_784,In_2894,In_2973);
or U785 (N_785,In_379,In_1019);
and U786 (N_786,In_1672,In_1691);
nor U787 (N_787,In_2371,In_2456);
nand U788 (N_788,In_129,In_899);
nor U789 (N_789,In_1936,In_1256);
or U790 (N_790,In_39,In_2365);
and U791 (N_791,In_541,In_2943);
nor U792 (N_792,In_101,In_164);
or U793 (N_793,In_454,In_2623);
and U794 (N_794,In_148,In_1643);
and U795 (N_795,In_1496,In_987);
and U796 (N_796,In_1209,In_2458);
or U797 (N_797,In_340,In_2420);
nand U798 (N_798,In_180,In_276);
or U799 (N_799,In_1339,In_194);
or U800 (N_800,In_601,In_208);
xor U801 (N_801,In_2732,In_1694);
nor U802 (N_802,In_316,In_2930);
nand U803 (N_803,In_665,In_2862);
and U804 (N_804,In_1279,In_138);
xnor U805 (N_805,In_124,In_260);
and U806 (N_806,In_1613,In_1047);
xor U807 (N_807,In_2700,In_2584);
or U808 (N_808,In_2651,In_2950);
nor U809 (N_809,In_1062,In_655);
and U810 (N_810,In_2126,In_2554);
nand U811 (N_811,In_2180,In_574);
or U812 (N_812,In_1285,In_1984);
or U813 (N_813,In_139,In_357);
or U814 (N_814,In_2045,In_2593);
nor U815 (N_815,In_2404,In_1552);
nand U816 (N_816,In_2668,In_1869);
or U817 (N_817,In_1073,In_214);
nor U818 (N_818,In_1066,In_562);
or U819 (N_819,In_1744,In_313);
or U820 (N_820,In_2882,In_547);
nor U821 (N_821,In_1474,In_1434);
nand U822 (N_822,In_2839,In_2155);
and U823 (N_823,In_763,In_2121);
nor U824 (N_824,In_1915,In_2681);
xnor U825 (N_825,In_1958,In_2437);
nor U826 (N_826,In_1372,In_2949);
nor U827 (N_827,In_1115,In_616);
nand U828 (N_828,In_1975,In_2522);
nand U829 (N_829,In_1302,In_1249);
nor U830 (N_830,In_815,In_566);
nor U831 (N_831,In_2105,In_1652);
nand U832 (N_832,In_1307,In_308);
or U833 (N_833,In_2648,In_1946);
or U834 (N_834,In_1480,In_873);
nor U835 (N_835,In_172,In_957);
and U836 (N_836,In_31,In_917);
nand U837 (N_837,In_278,In_1087);
or U838 (N_838,In_415,In_14);
nand U839 (N_839,In_2007,In_929);
nand U840 (N_840,In_1207,In_70);
or U841 (N_841,In_2820,In_1668);
xnor U842 (N_842,In_2349,In_2499);
nand U843 (N_843,In_1075,In_2118);
xnor U844 (N_844,In_1903,In_2969);
nor U845 (N_845,In_467,In_1995);
or U846 (N_846,In_1116,In_1964);
xor U847 (N_847,In_2555,In_2773);
or U848 (N_848,In_2629,In_589);
nor U849 (N_849,In_1133,In_2877);
and U850 (N_850,In_2331,In_2010);
nor U851 (N_851,In_1560,In_2833);
nor U852 (N_852,In_2690,In_1548);
and U853 (N_853,In_761,In_2221);
nor U854 (N_854,In_1123,In_1970);
and U855 (N_855,In_2599,In_2674);
xnor U856 (N_856,In_2079,In_497);
or U857 (N_857,In_2727,In_253);
or U858 (N_858,In_1313,In_748);
nor U859 (N_859,In_1528,In_1013);
nand U860 (N_860,In_1136,In_633);
and U861 (N_861,In_1704,In_2361);
nor U862 (N_862,In_505,In_749);
and U863 (N_863,In_270,In_2286);
nand U864 (N_864,In_671,In_1091);
nand U865 (N_865,In_631,In_268);
nand U866 (N_866,In_2507,In_1731);
nand U867 (N_867,In_2348,In_1381);
or U868 (N_868,In_563,In_1796);
nand U869 (N_869,In_1792,In_338);
nand U870 (N_870,In_2198,In_670);
and U871 (N_871,In_231,In_577);
xnor U872 (N_872,In_2576,In_115);
and U873 (N_873,In_2322,In_2741);
nor U874 (N_874,In_2187,In_414);
and U875 (N_875,In_780,In_511);
nand U876 (N_876,In_1743,In_2091);
and U877 (N_877,In_1853,In_1410);
or U878 (N_878,In_2772,In_926);
xnor U879 (N_879,In_532,In_579);
and U880 (N_880,In_887,In_1366);
nand U881 (N_881,In_2156,In_398);
nand U882 (N_882,In_2575,In_1721);
or U883 (N_883,In_539,In_2515);
or U884 (N_884,In_1907,In_739);
nand U885 (N_885,In_513,In_2217);
nand U886 (N_886,In_2759,In_500);
nor U887 (N_887,In_2937,In_2296);
nand U888 (N_888,In_221,In_1689);
nor U889 (N_889,In_1284,In_1610);
xor U890 (N_890,In_2595,In_335);
nand U891 (N_891,In_2671,In_882);
nor U892 (N_892,In_2354,In_1941);
xnor U893 (N_893,In_1246,In_758);
or U894 (N_894,In_1557,In_2481);
or U895 (N_895,In_1688,In_284);
nand U896 (N_896,In_1965,In_2143);
or U897 (N_897,In_561,In_1197);
nand U898 (N_898,In_2704,In_1872);
and U899 (N_899,In_2631,In_2062);
and U900 (N_900,In_697,In_1852);
nor U901 (N_901,In_1985,In_2088);
and U902 (N_902,In_2245,In_1130);
or U903 (N_903,In_2493,In_1215);
nor U904 (N_904,In_1106,In_1429);
xnor U905 (N_905,In_1110,In_1277);
or U906 (N_906,In_858,In_540);
and U907 (N_907,In_1681,In_1052);
nand U908 (N_908,In_733,In_1803);
xor U909 (N_909,In_1234,In_2063);
and U910 (N_910,In_1622,In_2795);
and U911 (N_911,In_2021,In_2655);
xnor U912 (N_912,In_569,In_2533);
or U913 (N_913,In_2996,In_310);
and U914 (N_914,In_1336,In_2147);
and U915 (N_915,In_789,In_407);
and U916 (N_916,In_2042,In_1839);
or U917 (N_917,In_2378,In_2089);
xnor U918 (N_918,In_2686,In_2102);
nand U919 (N_919,In_1233,In_2822);
nand U920 (N_920,In_1135,In_2030);
nand U921 (N_921,In_2093,In_1083);
or U922 (N_922,In_1601,In_1675);
nand U923 (N_923,In_1850,In_2596);
nand U924 (N_924,In_1165,In_1146);
nand U925 (N_925,In_609,In_1419);
xor U926 (N_926,In_2336,In_1442);
xnor U927 (N_927,In_1720,In_503);
or U928 (N_928,In_472,In_2830);
and U929 (N_929,In_1330,In_2071);
nand U930 (N_930,In_91,In_144);
nor U931 (N_931,In_1436,In_1527);
and U932 (N_932,In_2905,In_2070);
and U933 (N_933,In_2193,In_1705);
or U934 (N_934,In_485,In_2366);
and U935 (N_935,In_1159,In_526);
and U936 (N_936,In_1245,In_1742);
and U937 (N_937,In_1514,In_2491);
nor U938 (N_938,In_2938,In_1504);
or U939 (N_939,In_760,In_2630);
nand U940 (N_940,In_78,In_1309);
xor U941 (N_941,In_1849,In_2718);
nor U942 (N_942,In_437,In_1509);
or U943 (N_943,In_2326,In_465);
xor U944 (N_944,In_1881,In_911);
or U945 (N_945,In_2235,In_2981);
xnor U946 (N_946,In_2520,In_2000);
nand U947 (N_947,In_96,In_788);
or U948 (N_948,In_359,In_1676);
nor U949 (N_949,In_902,In_333);
and U950 (N_950,In_728,In_2119);
and U951 (N_951,In_2116,In_420);
nor U952 (N_952,In_2506,In_2689);
nor U953 (N_953,In_225,In_2486);
and U954 (N_954,In_717,In_555);
or U955 (N_955,In_393,In_2879);
and U956 (N_956,In_1026,In_2797);
and U957 (N_957,In_1012,In_2861);
or U958 (N_958,In_525,In_925);
nand U959 (N_959,In_1905,In_2604);
and U960 (N_960,In_304,In_1351);
nand U961 (N_961,In_713,In_2687);
xor U962 (N_962,In_447,In_1117);
nand U963 (N_963,In_2847,In_2725);
and U964 (N_964,In_2729,In_2152);
xor U965 (N_965,In_1861,In_2169);
xor U966 (N_966,In_1512,In_186);
and U967 (N_967,In_1746,In_480);
nand U968 (N_968,In_1921,In_2934);
nand U969 (N_969,In_325,In_679);
nand U970 (N_970,In_998,In_775);
or U971 (N_971,In_1664,In_2844);
xor U972 (N_972,In_1971,In_1420);
nand U973 (N_973,In_1568,In_1180);
nand U974 (N_974,In_102,In_1443);
nor U975 (N_975,In_2811,In_2050);
nand U976 (N_976,In_1773,In_2214);
and U977 (N_977,In_1524,In_2980);
nor U978 (N_978,In_1364,In_2733);
nor U979 (N_979,In_2804,In_1300);
and U980 (N_980,In_2047,In_1478);
or U981 (N_981,In_915,In_167);
nor U982 (N_982,In_153,In_2355);
or U983 (N_983,In_828,In_1928);
or U984 (N_984,In_2330,In_2027);
and U985 (N_985,In_2967,In_306);
and U986 (N_986,In_1191,In_451);
xor U987 (N_987,In_800,In_354);
or U988 (N_988,In_1666,In_2750);
and U989 (N_989,In_1968,In_2537);
nand U990 (N_990,In_2781,In_2389);
or U991 (N_991,In_924,In_2646);
or U992 (N_992,In_2375,In_871);
or U993 (N_993,In_1508,In_537);
nor U994 (N_994,In_2703,In_2598);
or U995 (N_995,In_1536,In_371);
or U996 (N_996,In_2964,In_785);
or U997 (N_997,In_459,In_698);
nand U998 (N_998,In_565,In_2140);
and U999 (N_999,In_2675,In_2754);
nand U1000 (N_1000,In_2189,In_2454);
nor U1001 (N_1001,In_2580,In_2320);
and U1002 (N_1002,In_1821,In_620);
nor U1003 (N_1003,In_1409,In_2566);
or U1004 (N_1004,In_1910,In_588);
nor U1005 (N_1005,In_1131,In_1870);
xor U1006 (N_1006,In_2513,In_2085);
or U1007 (N_1007,In_2663,In_2036);
nand U1008 (N_1008,In_2252,In_1707);
nor U1009 (N_1009,In_866,In_1598);
nor U1010 (N_1010,In_2243,In_1029);
or U1011 (N_1011,In_55,In_2824);
nor U1012 (N_1012,In_453,In_2970);
nand U1013 (N_1013,In_1128,In_636);
nor U1014 (N_1014,In_1783,In_2080);
or U1015 (N_1015,In_1723,In_2452);
nand U1016 (N_1016,In_2614,In_889);
nand U1017 (N_1017,In_2927,In_12);
xnor U1018 (N_1018,In_1144,In_830);
nand U1019 (N_1019,In_2726,In_1045);
nor U1020 (N_1020,In_440,In_2269);
nor U1021 (N_1021,In_1006,In_1005);
and U1022 (N_1022,In_2561,In_395);
xor U1023 (N_1023,In_1237,In_1127);
and U1024 (N_1024,In_2835,In_1266);
nand U1025 (N_1025,In_183,In_424);
or U1026 (N_1026,In_804,In_343);
nor U1027 (N_1027,In_137,In_1700);
nor U1028 (N_1028,In_2503,In_1034);
xnor U1029 (N_1029,In_2341,In_914);
and U1030 (N_1030,In_860,In_2840);
nand U1031 (N_1031,In_2730,In_271);
xnor U1032 (N_1032,In_2073,In_1293);
nor U1033 (N_1033,In_1608,In_365);
nand U1034 (N_1034,In_1699,In_2284);
xnor U1035 (N_1035,In_2766,In_328);
nand U1036 (N_1036,In_1426,In_476);
nor U1037 (N_1037,In_2549,In_657);
or U1038 (N_1038,In_2494,In_1892);
nand U1039 (N_1039,In_334,In_80);
nand U1040 (N_1040,In_394,In_1545);
nor U1041 (N_1041,In_602,In_1294);
or U1042 (N_1042,In_2569,In_772);
nor U1043 (N_1043,In_65,In_94);
nand U1044 (N_1044,In_1954,In_1811);
and U1045 (N_1045,In_2551,In_2669);
and U1046 (N_1046,In_2258,In_204);
or U1047 (N_1047,In_1674,In_1050);
or U1048 (N_1048,In_744,In_1932);
nand U1049 (N_1049,In_277,In_2103);
or U1050 (N_1050,In_1902,In_692);
nand U1051 (N_1051,In_2289,In_2789);
nor U1052 (N_1052,In_63,In_2976);
nor U1053 (N_1053,In_2049,In_199);
nand U1054 (N_1054,In_1126,In_2770);
nor U1055 (N_1055,In_639,In_1224);
and U1056 (N_1056,In_932,In_1173);
and U1057 (N_1057,In_348,In_142);
or U1058 (N_1058,In_1908,In_1160);
nand U1059 (N_1059,In_2161,In_922);
or U1060 (N_1060,In_1702,In_1632);
or U1061 (N_1061,In_833,In_2406);
and U1062 (N_1062,In_1491,In_2778);
or U1063 (N_1063,In_1184,In_2786);
or U1064 (N_1064,In_1739,In_1715);
nand U1065 (N_1065,In_2206,In_934);
or U1066 (N_1066,In_2090,In_650);
nand U1067 (N_1067,In_2951,In_2285);
or U1068 (N_1068,In_125,In_908);
xor U1069 (N_1069,In_1023,In_1068);
nor U1070 (N_1070,In_1724,In_1301);
and U1071 (N_1071,In_1768,In_1891);
xor U1072 (N_1072,In_2276,In_1893);
xnor U1073 (N_1073,In_2591,In_837);
or U1074 (N_1074,In_1487,In_232);
or U1075 (N_1075,In_178,In_1745);
or U1076 (N_1076,In_868,In_2993);
and U1077 (N_1077,In_1637,In_518);
nor U1078 (N_1078,In_1876,In_2869);
or U1079 (N_1079,In_2173,In_2918);
and U1080 (N_1080,In_2776,In_1826);
nor U1081 (N_1081,In_2434,In_2094);
and U1082 (N_1082,In_689,In_2411);
xor U1083 (N_1083,In_1566,In_1980);
or U1084 (N_1084,In_433,In_387);
nor U1085 (N_1085,In_1059,In_11);
nand U1086 (N_1086,In_939,In_878);
or U1087 (N_1087,In_1991,In_940);
and U1088 (N_1088,In_1086,In_1100);
and U1089 (N_1089,In_1290,In_1377);
nand U1090 (N_1090,In_1510,In_1046);
or U1091 (N_1091,In_1947,In_1468);
and U1092 (N_1092,In_1884,In_1402);
or U1093 (N_1093,In_1219,In_507);
or U1094 (N_1094,In_2821,In_1143);
or U1095 (N_1095,In_1392,In_179);
and U1096 (N_1096,In_2231,In_1886);
or U1097 (N_1097,In_116,In_110);
nand U1098 (N_1098,In_892,In_2281);
and U1099 (N_1099,In_988,In_211);
nor U1100 (N_1100,In_2171,In_1646);
or U1101 (N_1101,In_44,In_2057);
nor U1102 (N_1102,In_1583,In_2878);
or U1103 (N_1103,In_1798,In_1667);
nand U1104 (N_1104,In_1356,In_176);
nor U1105 (N_1105,In_2935,In_2983);
xor U1106 (N_1106,In_1008,In_1453);
and U1107 (N_1107,In_1017,In_2945);
and U1108 (N_1108,In_2302,In_724);
nand U1109 (N_1109,In_1374,In_1501);
nand U1110 (N_1110,In_2046,In_896);
xnor U1111 (N_1111,In_2470,In_1806);
nand U1112 (N_1112,In_1994,In_1036);
nor U1113 (N_1113,In_303,In_1866);
nand U1114 (N_1114,In_2308,In_1684);
or U1115 (N_1115,In_1650,In_1615);
or U1116 (N_1116,In_985,In_2809);
or U1117 (N_1117,In_1639,In_107);
or U1118 (N_1118,In_1001,In_1080);
nor U1119 (N_1119,In_894,In_981);
and U1120 (N_1120,In_2914,In_578);
or U1121 (N_1121,In_2954,In_2695);
or U1122 (N_1122,In_1890,In_2872);
nand U1123 (N_1123,In_1020,In_2756);
or U1124 (N_1124,In_2212,In_464);
and U1125 (N_1125,In_287,In_2291);
or U1126 (N_1126,In_412,In_469);
or U1127 (N_1127,In_498,In_0);
or U1128 (N_1128,In_502,In_989);
and U1129 (N_1129,In_191,In_731);
and U1130 (N_1130,In_177,In_1030);
and U1131 (N_1131,In_2612,In_2624);
nand U1132 (N_1132,In_26,In_2012);
or U1133 (N_1133,In_2433,In_397);
nand U1134 (N_1134,In_1687,In_1120);
or U1135 (N_1135,In_1218,In_754);
xnor U1136 (N_1136,In_931,In_88);
xor U1137 (N_1137,In_1641,In_2618);
or U1138 (N_1138,In_2953,In_2151);
or U1139 (N_1139,In_1642,In_974);
nor U1140 (N_1140,In_960,In_1489);
and U1141 (N_1141,In_1024,In_2345);
nand U1142 (N_1142,In_1002,In_2968);
and U1143 (N_1143,In_1031,In_2337);
or U1144 (N_1144,In_2567,In_1053);
or U1145 (N_1145,In_2653,In_1483);
or U1146 (N_1146,In_2900,In_803);
and U1147 (N_1147,In_2299,In_595);
and U1148 (N_1148,In_2540,In_1670);
and U1149 (N_1149,In_2525,In_1042);
nor U1150 (N_1150,In_104,In_166);
nand U1151 (N_1151,In_2608,In_1015);
nand U1152 (N_1152,In_2181,In_2416);
nor U1153 (N_1153,In_2032,In_2195);
nand U1154 (N_1154,In_161,In_2966);
xor U1155 (N_1155,In_1948,In_108);
nor U1156 (N_1156,In_2338,In_1933);
nor U1157 (N_1157,In_2106,In_2060);
and U1158 (N_1158,In_2607,In_322);
or U1159 (N_1159,In_2547,In_2743);
or U1160 (N_1160,In_169,In_2441);
and U1161 (N_1161,In_2921,In_1698);
nand U1162 (N_1162,In_1653,In_209);
nand U1163 (N_1163,In_68,In_888);
xor U1164 (N_1164,In_1348,In_1450);
nor U1165 (N_1165,In_2064,In_2259);
nor U1166 (N_1166,In_1183,In_2131);
and U1167 (N_1167,In_2022,In_2792);
or U1168 (N_1168,In_330,In_1114);
nand U1169 (N_1169,In_2114,In_2234);
nand U1170 (N_1170,In_2484,In_81);
nor U1171 (N_1171,In_1225,In_1635);
or U1172 (N_1172,In_1505,In_2924);
and U1173 (N_1173,In_516,In_2553);
nor U1174 (N_1174,In_258,In_787);
and U1175 (N_1175,In_1931,In_2138);
and U1176 (N_1176,In_880,In_1201);
nand U1177 (N_1177,In_1286,In_2177);
or U1178 (N_1178,In_1813,In_1476);
or U1179 (N_1179,In_203,In_2592);
and U1180 (N_1180,In_952,In_623);
nor U1181 (N_1181,In_475,In_2565);
nand U1182 (N_1182,In_2208,In_1231);
and U1183 (N_1183,In_2944,In_2013);
and U1184 (N_1184,In_2588,In_782);
nand U1185 (N_1185,In_1111,In_849);
and U1186 (N_1186,In_2300,In_35);
nand U1187 (N_1187,In_553,In_2508);
and U1188 (N_1188,In_1828,In_1574);
nor U1189 (N_1189,In_2794,In_1084);
and U1190 (N_1190,In_1105,In_1125);
or U1191 (N_1191,In_2662,In_968);
nand U1192 (N_1192,In_2986,In_2848);
or U1193 (N_1193,In_36,In_1810);
and U1194 (N_1194,In_2247,In_1361);
nand U1195 (N_1195,In_188,In_47);
and U1196 (N_1196,In_2812,In_558);
nand U1197 (N_1197,In_1484,In_1575);
and U1198 (N_1198,In_592,In_2577);
nand U1199 (N_1199,In_1922,In_1832);
or U1200 (N_1200,In_564,In_995);
or U1201 (N_1201,In_1275,In_1887);
and U1202 (N_1202,In_2994,In_1054);
nand U1203 (N_1203,In_1000,In_1864);
and U1204 (N_1204,In_1118,In_2904);
or U1205 (N_1205,In_1199,In_919);
nor U1206 (N_1206,In_89,In_2679);
and U1207 (N_1207,In_2479,In_673);
and U1208 (N_1208,In_2443,In_1750);
nand U1209 (N_1209,In_2574,In_584);
and U1210 (N_1210,In_2408,In_2098);
and U1211 (N_1211,In_946,In_2501);
and U1212 (N_1212,In_970,In_2003);
or U1213 (N_1213,In_275,In_1989);
nor U1214 (N_1214,In_2977,In_2684);
nand U1215 (N_1215,In_2971,In_1930);
xor U1216 (N_1216,In_59,In_2843);
nor U1217 (N_1217,In_494,In_1331);
and U1218 (N_1218,In_1553,In_1055);
and U1219 (N_1219,In_1998,In_1945);
nor U1220 (N_1220,In_1591,In_2340);
and U1221 (N_1221,In_1240,In_883);
nor U1222 (N_1222,In_506,In_2242);
and U1223 (N_1223,In_265,In_992);
xnor U1224 (N_1224,In_638,In_158);
or U1225 (N_1225,In_669,In_2606);
and U1226 (N_1226,In_1014,In_2261);
nand U1227 (N_1227,In_1119,In_2676);
or U1228 (N_1228,In_2394,In_1156);
nand U1229 (N_1229,In_321,In_1033);
xnor U1230 (N_1230,In_1594,In_890);
xnor U1231 (N_1231,In_1095,In_2505);
and U1232 (N_1232,In_2175,In_1791);
and U1233 (N_1233,In_1311,In_2213);
and U1234 (N_1234,In_128,In_691);
nand U1235 (N_1235,In_2236,In_1230);
nor U1236 (N_1236,In_1563,In_667);
or U1237 (N_1237,In_783,In_2170);
and U1238 (N_1238,In_2610,In_1076);
nor U1239 (N_1239,In_1376,In_400);
nand U1240 (N_1240,In_560,In_757);
nand U1241 (N_1241,In_2107,In_1541);
nor U1242 (N_1242,In_2963,In_2485);
or U1243 (N_1243,In_1493,In_2777);
and U1244 (N_1244,In_2714,In_2122);
nor U1245 (N_1245,In_1057,In_1926);
nor U1246 (N_1246,In_495,In_1787);
or U1247 (N_1247,In_2590,In_662);
xor U1248 (N_1248,In_1786,In_1802);
nor U1249 (N_1249,In_117,In_1463);
xor U1250 (N_1250,In_2400,In_1138);
nand U1251 (N_1251,In_538,In_1292);
or U1252 (N_1252,In_835,In_950);
nand U1253 (N_1253,In_2636,In_2288);
nor U1254 (N_1254,In_1885,In_2318);
nor U1255 (N_1255,In_1544,In_580);
or U1256 (N_1256,In_994,In_291);
or U1257 (N_1257,In_1973,In_2514);
nor U1258 (N_1258,In_604,In_206);
nor U1259 (N_1259,In_1179,In_1312);
nor U1260 (N_1260,In_2682,In_2423);
or U1261 (N_1261,In_1969,In_802);
or U1262 (N_1262,In_2719,In_1567);
nor U1263 (N_1263,In_1678,In_2842);
xnor U1264 (N_1264,In_1937,In_973);
nand U1265 (N_1265,In_1502,In_1323);
nand U1266 (N_1266,In_2311,In_213);
nor U1267 (N_1267,In_1149,In_118);
nor U1268 (N_1268,In_2321,In_452);
nor U1269 (N_1269,In_619,In_1722);
and U1270 (N_1270,In_1132,In_1041);
and U1271 (N_1271,In_2906,In_490);
or U1272 (N_1272,In_551,In_389);
xnor U1273 (N_1273,In_1603,In_2158);
and U1274 (N_1274,In_686,In_2294);
or U1275 (N_1275,In_1242,In_315);
and U1276 (N_1276,In_488,In_1844);
nand U1277 (N_1277,In_2999,In_2068);
nor U1278 (N_1278,In_1418,In_1735);
or U1279 (N_1279,In_301,In_2865);
or U1280 (N_1280,In_401,In_307);
nand U1281 (N_1281,In_1281,In_2034);
nor U1282 (N_1282,In_2959,In_1204);
nand U1283 (N_1283,In_1467,In_1490);
and U1284 (N_1284,In_2742,In_1032);
nand U1285 (N_1285,In_510,In_405);
and U1286 (N_1286,In_60,In_266);
and U1287 (N_1287,In_1840,In_1299);
nor U1288 (N_1288,In_455,In_2519);
xor U1289 (N_1289,In_814,In_2196);
and U1290 (N_1290,In_1446,In_385);
and U1291 (N_1291,In_197,In_2);
nand U1292 (N_1292,In_2386,In_1003);
nor U1293 (N_1293,In_2104,In_2813);
nand U1294 (N_1294,In_1846,In_1134);
nor U1295 (N_1295,In_2109,In_1607);
nor U1296 (N_1296,In_20,In_1319);
or U1297 (N_1297,In_162,In_236);
or U1298 (N_1298,In_2167,In_1719);
xor U1299 (N_1299,In_2427,In_1602);
nand U1300 (N_1300,In_2381,In_715);
nor U1301 (N_1301,In_2099,In_687);
and U1302 (N_1302,In_850,In_228);
and U1303 (N_1303,In_1569,In_456);
nand U1304 (N_1304,In_470,In_1475);
or U1305 (N_1305,In_1194,In_1090);
and U1306 (N_1306,In_1624,In_248);
and U1307 (N_1307,In_2160,In_2061);
nor U1308 (N_1308,In_1570,In_855);
xnor U1309 (N_1309,In_342,In_722);
or U1310 (N_1310,In_2315,In_1072);
or U1311 (N_1311,In_200,In_943);
and U1312 (N_1312,In_2438,In_2372);
nor U1313 (N_1313,In_2628,In_2306);
or U1314 (N_1314,In_1390,In_2455);
and U1315 (N_1315,In_25,In_1085);
or U1316 (N_1316,In_1187,In_2643);
xnor U1317 (N_1317,In_217,In_2816);
or U1318 (N_1318,In_701,In_392);
nand U1319 (N_1319,In_2178,In_76);
or U1320 (N_1320,In_1809,In_585);
or U1321 (N_1321,In_339,In_1113);
nor U1322 (N_1322,In_429,In_1829);
nand U1323 (N_1323,In_2722,In_2939);
and U1324 (N_1324,In_2562,In_2893);
nand U1325 (N_1325,In_2364,In_674);
nand U1326 (N_1326,In_2911,In_132);
or U1327 (N_1327,In_75,In_329);
nand U1328 (N_1328,In_718,In_2092);
and U1329 (N_1329,In_877,In_2831);
and U1330 (N_1330,In_2502,In_2854);
nor U1331 (N_1331,In_38,In_1823);
or U1332 (N_1332,In_2887,In_1322);
xor U1333 (N_1333,In_1774,In_42);
nand U1334 (N_1334,In_1439,In_1679);
or U1335 (N_1335,In_795,In_2897);
and U1336 (N_1336,In_1765,In_222);
and U1337 (N_1337,In_1357,In_536);
nor U1338 (N_1338,In_1094,In_544);
or U1339 (N_1339,In_2538,In_732);
nor U1340 (N_1340,In_1492,In_1206);
or U1341 (N_1341,In_2185,In_1252);
and U1342 (N_1342,In_821,In_2069);
xnor U1343 (N_1343,In_477,In_820);
or U1344 (N_1344,In_2279,In_1747);
xor U1345 (N_1345,In_1101,In_2521);
nor U1346 (N_1346,In_1289,In_1789);
or U1347 (N_1347,In_545,In_154);
nand U1348 (N_1348,In_927,In_953);
or U1349 (N_1349,In_910,In_24);
and U1350 (N_1350,In_1043,In_794);
nand U1351 (N_1351,In_1996,In_1794);
nor U1352 (N_1352,In_703,In_2256);
nor U1353 (N_1353,In_1808,In_2312);
nor U1354 (N_1354,In_838,In_1627);
or U1355 (N_1355,In_1186,In_3);
nand U1356 (N_1356,In_147,In_1103);
and U1357 (N_1357,In_1987,In_2432);
or U1358 (N_1358,In_1211,In_1271);
and U1359 (N_1359,In_1416,In_2957);
or U1360 (N_1360,In_2295,In_971);
or U1361 (N_1361,In_684,In_2249);
xnor U1362 (N_1362,In_2920,In_1529);
and U1363 (N_1363,In_1939,In_865);
nand U1364 (N_1364,In_839,In_1400);
nor U1365 (N_1365,In_2873,In_2654);
and U1366 (N_1366,In_255,In_1154);
and U1367 (N_1367,In_300,In_215);
or U1368 (N_1368,In_1779,In_2611);
nand U1369 (N_1369,In_1732,In_1214);
xor U1370 (N_1370,In_190,In_1769);
or U1371 (N_1371,In_1383,In_356);
or U1372 (N_1372,In_1208,In_730);
or U1373 (N_1373,In_1212,In_2199);
nand U1374 (N_1374,In_2182,In_1278);
xor U1375 (N_1375,In_15,In_250);
and U1376 (N_1376,In_1532,In_1346);
nand U1377 (N_1377,In_2421,In_2936);
nand U1378 (N_1378,In_1518,In_2644);
xnor U1379 (N_1379,In_1979,In_2881);
or U1380 (N_1380,In_935,In_226);
nor U1381 (N_1381,In_1079,In_2579);
or U1382 (N_1382,In_295,In_2739);
nand U1383 (N_1383,In_2040,In_581);
nand U1384 (N_1384,In_2130,In_1485);
nor U1385 (N_1385,In_1579,In_4);
nor U1386 (N_1386,In_1956,In_445);
and U1387 (N_1387,In_1477,In_755);
or U1388 (N_1388,In_2661,In_2360);
nand U1389 (N_1389,In_254,In_443);
nand U1390 (N_1390,In_895,In_806);
nor U1391 (N_1391,In_1280,In_1457);
or U1392 (N_1392,In_2237,In_1243);
nor U1393 (N_1393,In_2081,In_709);
and U1394 (N_1394,In_32,In_2808);
or U1395 (N_1395,In_836,In_1549);
nor U1396 (N_1396,In_10,In_575);
nand U1397 (N_1397,In_1733,In_1834);
nand U1398 (N_1398,In_2658,In_458);
or U1399 (N_1399,In_1190,In_103);
nor U1400 (N_1400,In_2202,In_781);
or U1401 (N_1401,In_157,In_909);
nand U1402 (N_1402,In_2402,In_2128);
nand U1403 (N_1403,In_1706,In_22);
nand U1404 (N_1404,In_2020,In_2384);
or U1405 (N_1405,In_947,In_1027);
nand U1406 (N_1406,In_610,In_1282);
and U1407 (N_1407,In_1795,In_18);
and U1408 (N_1408,In_2006,In_2305);
nor U1409 (N_1409,In_230,In_2819);
nor U1410 (N_1410,In_1009,In_27);
xnor U1411 (N_1411,In_1894,In_369);
nor U1412 (N_1412,In_1513,In_238);
nor U1413 (N_1413,In_1412,In_656);
and U1414 (N_1414,In_49,In_1065);
and U1415 (N_1415,In_2925,In_2827);
or U1416 (N_1416,In_791,In_1081);
or U1417 (N_1417,In_1725,In_753);
and U1418 (N_1418,In_891,In_1395);
and U1419 (N_1419,In_955,In_93);
or U1420 (N_1420,In_2744,In_2988);
nand U1421 (N_1421,In_583,In_2065);
and U1422 (N_1422,In_1755,In_1818);
nand U1423 (N_1423,In_1648,In_2159);
or U1424 (N_1424,In_1018,In_1924);
nand U1425 (N_1425,In_823,In_1981);
or U1426 (N_1426,In_243,In_1345);
nor U1427 (N_1427,In_1471,In_2544);
nor U1428 (N_1428,In_612,In_2884);
nor U1429 (N_1429,In_607,In_2710);
nand U1430 (N_1430,In_419,In_976);
and U1431 (N_1431,In_2600,In_2309);
or U1432 (N_1432,In_2955,In_2793);
nand U1433 (N_1433,In_1875,In_1836);
nand U1434 (N_1434,In_2031,In_735);
nor U1435 (N_1435,In_900,In_309);
nand U1436 (N_1436,In_160,In_2737);
and U1437 (N_1437,In_2229,In_1590);
or U1438 (N_1438,In_1614,In_2748);
and U1439 (N_1439,In_645,In_1335);
or U1440 (N_1440,In_848,In_1329);
or U1441 (N_1441,In_928,In_1827);
and U1442 (N_1442,In_285,In_1060);
and U1443 (N_1443,In_1220,In_1140);
and U1444 (N_1444,In_2014,In_244);
nand U1445 (N_1445,In_1565,In_845);
and U1446 (N_1446,In_235,In_2620);
and U1447 (N_1447,In_2186,In_1486);
nand U1448 (N_1448,In_1804,In_2912);
nand U1449 (N_1449,In_613,In_2941);
or U1450 (N_1450,In_2597,In_2667);
nor U1451 (N_1451,In_1717,In_2796);
nor U1452 (N_1452,In_286,In_897);
nand U1453 (N_1453,In_2145,In_1071);
nand U1454 (N_1454,In_966,In_2440);
and U1455 (N_1455,In_1253,In_930);
or U1456 (N_1456,In_1232,In_629);
xnor U1457 (N_1457,In_184,In_809);
or U1458 (N_1458,In_247,In_1175);
nand U1459 (N_1459,In_1205,In_413);
nand U1460 (N_1460,In_2761,In_2431);
nand U1461 (N_1461,In_1415,In_2637);
nor U1462 (N_1462,In_696,In_434);
nand U1463 (N_1463,In_527,In_1171);
xnor U1464 (N_1464,In_1176,In_2998);
nand U1465 (N_1465,In_1387,In_2278);
or U1466 (N_1466,In_1196,In_1858);
or U1467 (N_1467,In_1359,In_363);
nor U1468 (N_1468,In_187,In_73);
xor U1469 (N_1469,In_1102,In_205);
xor U1470 (N_1470,In_2346,In_1863);
nand U1471 (N_1471,In_1216,In_1178);
nor U1472 (N_1472,In_2885,In_121);
and U1473 (N_1473,In_1261,In_1554);
and U1474 (N_1474,In_2277,In_1254);
nand U1475 (N_1475,In_377,In_790);
nand U1476 (N_1476,In_912,In_2757);
xnor U1477 (N_1477,In_590,In_1460);
nand U1478 (N_1478,In_570,In_432);
or U1479 (N_1479,In_2828,In_812);
nor U1480 (N_1480,In_1435,In_2275);
and U1481 (N_1481,In_46,In_1752);
nand U1482 (N_1482,In_2445,In_1660);
and U1483 (N_1483,In_921,In_2053);
nand U1484 (N_1484,In_2990,In_504);
and U1485 (N_1485,In_2112,In_2698);
nand U1486 (N_1486,In_2124,In_1451);
nor U1487 (N_1487,In_1895,In_374);
and U1488 (N_1488,In_1659,In_1358);
or U1489 (N_1489,In_2086,In_2788);
nand U1490 (N_1490,In_1456,In_113);
nand U1491 (N_1491,In_1440,In_2559);
and U1492 (N_1492,In_628,In_471);
xor U1493 (N_1493,In_624,In_524);
and U1494 (N_1494,In_1155,In_597);
nor U1495 (N_1495,In_274,In_626);
and U1496 (N_1496,In_1546,In_448);
or U1497 (N_1497,In_1879,In_2083);
nand U1498 (N_1498,In_207,In_1396);
nor U1499 (N_1499,In_2622,In_2133);
nand U1500 (N_1500,In_205,In_2936);
or U1501 (N_1501,In_1600,In_2332);
nand U1502 (N_1502,In_369,In_756);
nor U1503 (N_1503,In_1159,In_1154);
nor U1504 (N_1504,In_2236,In_165);
and U1505 (N_1505,In_1368,In_1502);
and U1506 (N_1506,In_428,In_2571);
and U1507 (N_1507,In_141,In_1640);
nand U1508 (N_1508,In_2073,In_773);
xnor U1509 (N_1509,In_114,In_2030);
nand U1510 (N_1510,In_120,In_1450);
xor U1511 (N_1511,In_1504,In_2913);
or U1512 (N_1512,In_785,In_2279);
and U1513 (N_1513,In_1308,In_184);
xor U1514 (N_1514,In_2810,In_897);
or U1515 (N_1515,In_672,In_1894);
xnor U1516 (N_1516,In_2158,In_1022);
nor U1517 (N_1517,In_2172,In_923);
and U1518 (N_1518,In_1196,In_910);
nand U1519 (N_1519,In_646,In_1450);
nand U1520 (N_1520,In_2475,In_1696);
nor U1521 (N_1521,In_413,In_1251);
nor U1522 (N_1522,In_1517,In_1026);
nor U1523 (N_1523,In_1358,In_1637);
or U1524 (N_1524,In_577,In_2078);
xor U1525 (N_1525,In_349,In_1478);
or U1526 (N_1526,In_1170,In_1593);
and U1527 (N_1527,In_2030,In_1047);
or U1528 (N_1528,In_2986,In_1294);
and U1529 (N_1529,In_1638,In_2401);
nor U1530 (N_1530,In_688,In_472);
or U1531 (N_1531,In_230,In_2438);
nor U1532 (N_1532,In_2490,In_1294);
or U1533 (N_1533,In_2876,In_610);
nor U1534 (N_1534,In_2677,In_2569);
nor U1535 (N_1535,In_606,In_1237);
and U1536 (N_1536,In_1131,In_1952);
nor U1537 (N_1537,In_1667,In_2536);
nand U1538 (N_1538,In_1224,In_2376);
or U1539 (N_1539,In_1071,In_2546);
and U1540 (N_1540,In_564,In_163);
or U1541 (N_1541,In_2908,In_868);
or U1542 (N_1542,In_2290,In_112);
and U1543 (N_1543,In_2203,In_383);
and U1544 (N_1544,In_148,In_889);
or U1545 (N_1545,In_2923,In_498);
and U1546 (N_1546,In_397,In_372);
or U1547 (N_1547,In_2008,In_1736);
xor U1548 (N_1548,In_1977,In_1159);
and U1549 (N_1549,In_1237,In_2058);
or U1550 (N_1550,In_1659,In_2235);
nor U1551 (N_1551,In_1979,In_671);
or U1552 (N_1552,In_2170,In_2163);
nor U1553 (N_1553,In_816,In_1546);
and U1554 (N_1554,In_0,In_1685);
xnor U1555 (N_1555,In_2208,In_1214);
nand U1556 (N_1556,In_76,In_530);
and U1557 (N_1557,In_1645,In_874);
nand U1558 (N_1558,In_691,In_1488);
nand U1559 (N_1559,In_1898,In_384);
nor U1560 (N_1560,In_2367,In_2427);
or U1561 (N_1561,In_1236,In_1560);
or U1562 (N_1562,In_1494,In_1003);
or U1563 (N_1563,In_1254,In_666);
nor U1564 (N_1564,In_2365,In_1852);
nand U1565 (N_1565,In_1572,In_1107);
xnor U1566 (N_1566,In_1475,In_301);
or U1567 (N_1567,In_240,In_936);
nand U1568 (N_1568,In_2930,In_2751);
or U1569 (N_1569,In_2772,In_2347);
or U1570 (N_1570,In_2367,In_143);
and U1571 (N_1571,In_979,In_2811);
and U1572 (N_1572,In_2332,In_2307);
nor U1573 (N_1573,In_1568,In_2284);
nor U1574 (N_1574,In_2078,In_418);
nor U1575 (N_1575,In_2477,In_1335);
or U1576 (N_1576,In_1414,In_505);
nand U1577 (N_1577,In_214,In_1627);
and U1578 (N_1578,In_592,In_322);
or U1579 (N_1579,In_1630,In_387);
nor U1580 (N_1580,In_1023,In_1236);
and U1581 (N_1581,In_1546,In_1910);
nor U1582 (N_1582,In_1381,In_2966);
nor U1583 (N_1583,In_36,In_720);
nand U1584 (N_1584,In_1129,In_182);
nand U1585 (N_1585,In_778,In_1);
nand U1586 (N_1586,In_2360,In_2408);
xor U1587 (N_1587,In_2486,In_1796);
and U1588 (N_1588,In_556,In_45);
or U1589 (N_1589,In_2776,In_2237);
nor U1590 (N_1590,In_1200,In_727);
or U1591 (N_1591,In_1847,In_1551);
nand U1592 (N_1592,In_832,In_1201);
and U1593 (N_1593,In_275,In_357);
nor U1594 (N_1594,In_769,In_2732);
and U1595 (N_1595,In_2833,In_2829);
and U1596 (N_1596,In_1405,In_1683);
or U1597 (N_1597,In_192,In_2988);
nand U1598 (N_1598,In_656,In_1712);
nor U1599 (N_1599,In_1797,In_1557);
xor U1600 (N_1600,In_2519,In_2188);
nand U1601 (N_1601,In_2061,In_507);
or U1602 (N_1602,In_897,In_610);
nand U1603 (N_1603,In_2764,In_789);
nand U1604 (N_1604,In_2154,In_1856);
nor U1605 (N_1605,In_2930,In_39);
xnor U1606 (N_1606,In_1616,In_1514);
nand U1607 (N_1607,In_663,In_462);
or U1608 (N_1608,In_2765,In_2880);
nand U1609 (N_1609,In_14,In_1606);
or U1610 (N_1610,In_2000,In_2328);
and U1611 (N_1611,In_873,In_2816);
nand U1612 (N_1612,In_2761,In_1577);
nand U1613 (N_1613,In_2468,In_2921);
or U1614 (N_1614,In_1356,In_856);
nand U1615 (N_1615,In_2769,In_699);
nand U1616 (N_1616,In_1438,In_2797);
nand U1617 (N_1617,In_1693,In_1035);
nand U1618 (N_1618,In_1827,In_1298);
nand U1619 (N_1619,In_1133,In_287);
nor U1620 (N_1620,In_2178,In_2839);
and U1621 (N_1621,In_1565,In_822);
xnor U1622 (N_1622,In_8,In_1828);
nand U1623 (N_1623,In_1230,In_43);
or U1624 (N_1624,In_2162,In_1938);
xor U1625 (N_1625,In_749,In_520);
and U1626 (N_1626,In_2591,In_2637);
or U1627 (N_1627,In_999,In_1576);
and U1628 (N_1628,In_218,In_1694);
and U1629 (N_1629,In_291,In_738);
and U1630 (N_1630,In_1953,In_76);
nor U1631 (N_1631,In_2413,In_2232);
or U1632 (N_1632,In_2330,In_409);
or U1633 (N_1633,In_735,In_1048);
nor U1634 (N_1634,In_2942,In_983);
or U1635 (N_1635,In_2561,In_2618);
or U1636 (N_1636,In_2126,In_298);
and U1637 (N_1637,In_2035,In_1546);
nor U1638 (N_1638,In_42,In_2459);
nor U1639 (N_1639,In_941,In_1304);
xnor U1640 (N_1640,In_10,In_2367);
nor U1641 (N_1641,In_2672,In_665);
and U1642 (N_1642,In_670,In_806);
nand U1643 (N_1643,In_280,In_2265);
nor U1644 (N_1644,In_2752,In_1501);
or U1645 (N_1645,In_2224,In_825);
xor U1646 (N_1646,In_1240,In_632);
or U1647 (N_1647,In_1315,In_1062);
or U1648 (N_1648,In_1938,In_2370);
nand U1649 (N_1649,In_2611,In_1483);
or U1650 (N_1650,In_715,In_215);
nor U1651 (N_1651,In_878,In_1592);
and U1652 (N_1652,In_1513,In_125);
xnor U1653 (N_1653,In_1037,In_1271);
nand U1654 (N_1654,In_2281,In_1081);
or U1655 (N_1655,In_2067,In_833);
nand U1656 (N_1656,In_2822,In_2225);
and U1657 (N_1657,In_1238,In_2161);
or U1658 (N_1658,In_2623,In_2544);
nand U1659 (N_1659,In_506,In_128);
and U1660 (N_1660,In_1091,In_1590);
nor U1661 (N_1661,In_1754,In_2857);
nor U1662 (N_1662,In_713,In_2538);
and U1663 (N_1663,In_2350,In_1724);
and U1664 (N_1664,In_407,In_799);
or U1665 (N_1665,In_2296,In_141);
nand U1666 (N_1666,In_1798,In_570);
nand U1667 (N_1667,In_459,In_32);
and U1668 (N_1668,In_2659,In_2990);
and U1669 (N_1669,In_253,In_2840);
nor U1670 (N_1670,In_2500,In_1816);
nor U1671 (N_1671,In_565,In_2873);
nand U1672 (N_1672,In_1901,In_263);
and U1673 (N_1673,In_269,In_2553);
nor U1674 (N_1674,In_170,In_1472);
or U1675 (N_1675,In_1622,In_2152);
nand U1676 (N_1676,In_1300,In_2064);
or U1677 (N_1677,In_2914,In_1487);
or U1678 (N_1678,In_633,In_402);
or U1679 (N_1679,In_1287,In_2217);
nand U1680 (N_1680,In_620,In_2345);
nor U1681 (N_1681,In_1062,In_1285);
or U1682 (N_1682,In_1933,In_2129);
xnor U1683 (N_1683,In_1779,In_1777);
and U1684 (N_1684,In_1402,In_2127);
and U1685 (N_1685,In_18,In_352);
nor U1686 (N_1686,In_2898,In_507);
nor U1687 (N_1687,In_2610,In_2557);
nand U1688 (N_1688,In_2388,In_2030);
or U1689 (N_1689,In_354,In_1169);
nand U1690 (N_1690,In_508,In_781);
nor U1691 (N_1691,In_2440,In_767);
and U1692 (N_1692,In_2472,In_256);
or U1693 (N_1693,In_738,In_1681);
xor U1694 (N_1694,In_1574,In_2185);
xnor U1695 (N_1695,In_211,In_2606);
nor U1696 (N_1696,In_2766,In_2394);
or U1697 (N_1697,In_2696,In_72);
nor U1698 (N_1698,In_939,In_2790);
xor U1699 (N_1699,In_2103,In_724);
or U1700 (N_1700,In_1718,In_111);
nand U1701 (N_1701,In_1211,In_2342);
nand U1702 (N_1702,In_164,In_121);
nand U1703 (N_1703,In_2449,In_1180);
xnor U1704 (N_1704,In_1924,In_1994);
or U1705 (N_1705,In_2340,In_1812);
nand U1706 (N_1706,In_1441,In_2423);
or U1707 (N_1707,In_1163,In_1559);
xnor U1708 (N_1708,In_1269,In_1748);
or U1709 (N_1709,In_2747,In_519);
xnor U1710 (N_1710,In_2336,In_684);
nand U1711 (N_1711,In_1590,In_103);
or U1712 (N_1712,In_1697,In_516);
xor U1713 (N_1713,In_2017,In_227);
or U1714 (N_1714,In_1615,In_2366);
or U1715 (N_1715,In_1646,In_1736);
and U1716 (N_1716,In_690,In_853);
nor U1717 (N_1717,In_724,In_416);
nor U1718 (N_1718,In_879,In_790);
xnor U1719 (N_1719,In_839,In_179);
nor U1720 (N_1720,In_894,In_1970);
xnor U1721 (N_1721,In_2084,In_258);
nand U1722 (N_1722,In_1561,In_839);
nor U1723 (N_1723,In_172,In_2172);
or U1724 (N_1724,In_162,In_428);
and U1725 (N_1725,In_118,In_2512);
or U1726 (N_1726,In_212,In_2795);
and U1727 (N_1727,In_2144,In_1166);
nand U1728 (N_1728,In_1096,In_2087);
or U1729 (N_1729,In_1788,In_453);
and U1730 (N_1730,In_1059,In_2107);
or U1731 (N_1731,In_2313,In_1090);
and U1732 (N_1732,In_940,In_1550);
nand U1733 (N_1733,In_2819,In_813);
and U1734 (N_1734,In_1707,In_1328);
and U1735 (N_1735,In_2277,In_2033);
nand U1736 (N_1736,In_2243,In_2527);
nand U1737 (N_1737,In_2087,In_708);
nand U1738 (N_1738,In_146,In_173);
or U1739 (N_1739,In_2336,In_1920);
nor U1740 (N_1740,In_2471,In_2695);
nor U1741 (N_1741,In_1812,In_617);
nand U1742 (N_1742,In_2356,In_345);
xnor U1743 (N_1743,In_2392,In_2608);
and U1744 (N_1744,In_2532,In_1254);
or U1745 (N_1745,In_1109,In_577);
and U1746 (N_1746,In_1706,In_2659);
and U1747 (N_1747,In_2178,In_798);
nor U1748 (N_1748,In_53,In_1761);
nand U1749 (N_1749,In_2806,In_2450);
and U1750 (N_1750,In_1901,In_2789);
and U1751 (N_1751,In_1573,In_1760);
nand U1752 (N_1752,In_996,In_2699);
and U1753 (N_1753,In_2873,In_255);
and U1754 (N_1754,In_992,In_1941);
nor U1755 (N_1755,In_1087,In_435);
and U1756 (N_1756,In_1737,In_489);
nand U1757 (N_1757,In_1861,In_2747);
or U1758 (N_1758,In_2395,In_249);
and U1759 (N_1759,In_1471,In_2723);
nand U1760 (N_1760,In_2287,In_2198);
nand U1761 (N_1761,In_1922,In_445);
and U1762 (N_1762,In_1467,In_2611);
nor U1763 (N_1763,In_1539,In_1342);
nor U1764 (N_1764,In_138,In_175);
nand U1765 (N_1765,In_2089,In_1265);
or U1766 (N_1766,In_2982,In_2608);
nor U1767 (N_1767,In_1904,In_185);
nor U1768 (N_1768,In_1184,In_85);
nand U1769 (N_1769,In_221,In_1764);
and U1770 (N_1770,In_1025,In_2906);
nand U1771 (N_1771,In_2972,In_1212);
nor U1772 (N_1772,In_1948,In_2213);
xnor U1773 (N_1773,In_2683,In_2450);
or U1774 (N_1774,In_1090,In_2312);
nand U1775 (N_1775,In_561,In_1910);
or U1776 (N_1776,In_1881,In_1058);
or U1777 (N_1777,In_2314,In_645);
and U1778 (N_1778,In_1867,In_5);
nand U1779 (N_1779,In_2155,In_902);
nor U1780 (N_1780,In_2741,In_518);
and U1781 (N_1781,In_2223,In_1621);
nor U1782 (N_1782,In_329,In_1902);
nand U1783 (N_1783,In_1163,In_1408);
or U1784 (N_1784,In_2100,In_2331);
or U1785 (N_1785,In_1670,In_1943);
nor U1786 (N_1786,In_2553,In_1118);
xnor U1787 (N_1787,In_18,In_1782);
or U1788 (N_1788,In_767,In_1542);
or U1789 (N_1789,In_339,In_1570);
nor U1790 (N_1790,In_1833,In_2723);
and U1791 (N_1791,In_2121,In_2842);
xor U1792 (N_1792,In_1259,In_2984);
nor U1793 (N_1793,In_2641,In_709);
or U1794 (N_1794,In_2688,In_2600);
nand U1795 (N_1795,In_885,In_2261);
nor U1796 (N_1796,In_1020,In_143);
nand U1797 (N_1797,In_553,In_1722);
nor U1798 (N_1798,In_95,In_2244);
xor U1799 (N_1799,In_1813,In_1400);
nor U1800 (N_1800,In_222,In_1356);
or U1801 (N_1801,In_241,In_2256);
or U1802 (N_1802,In_2533,In_56);
and U1803 (N_1803,In_1649,In_2420);
nand U1804 (N_1804,In_917,In_1378);
xor U1805 (N_1805,In_2354,In_552);
nor U1806 (N_1806,In_1128,In_78);
nand U1807 (N_1807,In_2429,In_1143);
or U1808 (N_1808,In_1363,In_533);
nor U1809 (N_1809,In_686,In_1605);
nor U1810 (N_1810,In_1780,In_7);
nand U1811 (N_1811,In_2305,In_2383);
and U1812 (N_1812,In_1287,In_317);
and U1813 (N_1813,In_285,In_2872);
nor U1814 (N_1814,In_755,In_2741);
or U1815 (N_1815,In_1878,In_1941);
nor U1816 (N_1816,In_2504,In_1349);
nor U1817 (N_1817,In_2147,In_1366);
nand U1818 (N_1818,In_1295,In_984);
nor U1819 (N_1819,In_507,In_2483);
and U1820 (N_1820,In_1643,In_1676);
nor U1821 (N_1821,In_248,In_2268);
and U1822 (N_1822,In_537,In_402);
or U1823 (N_1823,In_70,In_574);
xnor U1824 (N_1824,In_2483,In_2044);
nand U1825 (N_1825,In_2999,In_484);
nor U1826 (N_1826,In_2815,In_1792);
and U1827 (N_1827,In_2088,In_342);
and U1828 (N_1828,In_1445,In_1596);
nor U1829 (N_1829,In_518,In_4);
nor U1830 (N_1830,In_2985,In_911);
or U1831 (N_1831,In_806,In_110);
nor U1832 (N_1832,In_1821,In_1744);
nand U1833 (N_1833,In_1966,In_1473);
nor U1834 (N_1834,In_465,In_2520);
nor U1835 (N_1835,In_2833,In_249);
and U1836 (N_1836,In_1822,In_699);
or U1837 (N_1837,In_26,In_2103);
and U1838 (N_1838,In_1519,In_213);
nor U1839 (N_1839,In_1025,In_2935);
nand U1840 (N_1840,In_829,In_1186);
or U1841 (N_1841,In_1158,In_2253);
nand U1842 (N_1842,In_326,In_1177);
or U1843 (N_1843,In_2320,In_2406);
and U1844 (N_1844,In_2152,In_1612);
nand U1845 (N_1845,In_1638,In_146);
nor U1846 (N_1846,In_1707,In_1853);
nor U1847 (N_1847,In_1161,In_2533);
nor U1848 (N_1848,In_644,In_2291);
xnor U1849 (N_1849,In_414,In_448);
nand U1850 (N_1850,In_649,In_2100);
and U1851 (N_1851,In_2096,In_576);
nor U1852 (N_1852,In_2592,In_2026);
nor U1853 (N_1853,In_2542,In_1279);
and U1854 (N_1854,In_1108,In_1797);
nor U1855 (N_1855,In_921,In_2494);
xnor U1856 (N_1856,In_2049,In_2486);
nand U1857 (N_1857,In_2593,In_2299);
and U1858 (N_1858,In_1507,In_2153);
and U1859 (N_1859,In_113,In_581);
nor U1860 (N_1860,In_649,In_1553);
nor U1861 (N_1861,In_2648,In_1703);
or U1862 (N_1862,In_1985,In_1981);
or U1863 (N_1863,In_2337,In_2445);
nand U1864 (N_1864,In_444,In_1571);
nor U1865 (N_1865,In_2249,In_2466);
and U1866 (N_1866,In_2840,In_1287);
nor U1867 (N_1867,In_1709,In_827);
and U1868 (N_1868,In_1192,In_2196);
nor U1869 (N_1869,In_2866,In_1758);
nor U1870 (N_1870,In_1009,In_854);
nand U1871 (N_1871,In_879,In_1493);
or U1872 (N_1872,In_375,In_1928);
nand U1873 (N_1873,In_361,In_1131);
nor U1874 (N_1874,In_2152,In_2915);
and U1875 (N_1875,In_166,In_2310);
nand U1876 (N_1876,In_1302,In_2499);
and U1877 (N_1877,In_1274,In_1304);
and U1878 (N_1878,In_2111,In_1341);
and U1879 (N_1879,In_765,In_2151);
or U1880 (N_1880,In_2206,In_1668);
xnor U1881 (N_1881,In_1290,In_2422);
and U1882 (N_1882,In_2417,In_1032);
and U1883 (N_1883,In_545,In_1078);
and U1884 (N_1884,In_784,In_2183);
xor U1885 (N_1885,In_1439,In_1403);
nor U1886 (N_1886,In_1975,In_719);
nand U1887 (N_1887,In_2569,In_863);
nand U1888 (N_1888,In_2001,In_1694);
nor U1889 (N_1889,In_1803,In_765);
or U1890 (N_1890,In_687,In_2316);
and U1891 (N_1891,In_940,In_2082);
nor U1892 (N_1892,In_1679,In_2226);
xnor U1893 (N_1893,In_1884,In_1430);
or U1894 (N_1894,In_1040,In_2212);
nand U1895 (N_1895,In_1450,In_2757);
and U1896 (N_1896,In_2395,In_2142);
or U1897 (N_1897,In_2001,In_1552);
or U1898 (N_1898,In_860,In_1345);
and U1899 (N_1899,In_1556,In_1572);
and U1900 (N_1900,In_1806,In_2352);
nand U1901 (N_1901,In_1524,In_166);
nand U1902 (N_1902,In_2732,In_839);
nor U1903 (N_1903,In_695,In_995);
or U1904 (N_1904,In_540,In_2559);
nor U1905 (N_1905,In_480,In_489);
nor U1906 (N_1906,In_2212,In_977);
and U1907 (N_1907,In_105,In_968);
nand U1908 (N_1908,In_1710,In_893);
nor U1909 (N_1909,In_141,In_1670);
nor U1910 (N_1910,In_2486,In_1574);
nand U1911 (N_1911,In_1041,In_2002);
or U1912 (N_1912,In_859,In_159);
nor U1913 (N_1913,In_2689,In_1671);
and U1914 (N_1914,In_1679,In_2128);
nand U1915 (N_1915,In_945,In_689);
nand U1916 (N_1916,In_991,In_2620);
xnor U1917 (N_1917,In_2996,In_639);
xor U1918 (N_1918,In_2310,In_663);
nand U1919 (N_1919,In_494,In_829);
nand U1920 (N_1920,In_1887,In_2003);
or U1921 (N_1921,In_2701,In_1491);
or U1922 (N_1922,In_174,In_2180);
and U1923 (N_1923,In_2844,In_303);
nand U1924 (N_1924,In_908,In_1056);
nand U1925 (N_1925,In_2392,In_486);
or U1926 (N_1926,In_1245,In_2934);
nand U1927 (N_1927,In_2694,In_2175);
nor U1928 (N_1928,In_2124,In_797);
nand U1929 (N_1929,In_495,In_2609);
or U1930 (N_1930,In_1003,In_2967);
or U1931 (N_1931,In_2640,In_2838);
nor U1932 (N_1932,In_1489,In_721);
nand U1933 (N_1933,In_89,In_1726);
nand U1934 (N_1934,In_628,In_2688);
or U1935 (N_1935,In_2818,In_2756);
nand U1936 (N_1936,In_377,In_2621);
nand U1937 (N_1937,In_866,In_1174);
nand U1938 (N_1938,In_698,In_373);
nor U1939 (N_1939,In_2202,In_2697);
and U1940 (N_1940,In_2407,In_344);
and U1941 (N_1941,In_638,In_1238);
or U1942 (N_1942,In_2501,In_1986);
and U1943 (N_1943,In_2679,In_794);
and U1944 (N_1944,In_2328,In_1428);
nand U1945 (N_1945,In_199,In_721);
or U1946 (N_1946,In_627,In_1528);
nor U1947 (N_1947,In_910,In_2954);
nand U1948 (N_1948,In_1731,In_1271);
and U1949 (N_1949,In_1795,In_919);
and U1950 (N_1950,In_2717,In_1230);
nor U1951 (N_1951,In_2941,In_1936);
and U1952 (N_1952,In_1491,In_790);
and U1953 (N_1953,In_1577,In_778);
nand U1954 (N_1954,In_2419,In_421);
or U1955 (N_1955,In_402,In_1506);
nand U1956 (N_1956,In_2920,In_930);
or U1957 (N_1957,In_669,In_2678);
or U1958 (N_1958,In_1784,In_744);
nor U1959 (N_1959,In_1708,In_2583);
or U1960 (N_1960,In_1840,In_408);
xnor U1961 (N_1961,In_1608,In_2323);
and U1962 (N_1962,In_1176,In_815);
or U1963 (N_1963,In_2442,In_652);
nand U1964 (N_1964,In_1958,In_2018);
nand U1965 (N_1965,In_207,In_2388);
nor U1966 (N_1966,In_748,In_2474);
or U1967 (N_1967,In_503,In_1214);
or U1968 (N_1968,In_2955,In_2883);
nand U1969 (N_1969,In_2278,In_1688);
or U1970 (N_1970,In_133,In_223);
or U1971 (N_1971,In_1034,In_2349);
nand U1972 (N_1972,In_112,In_1421);
nand U1973 (N_1973,In_491,In_1273);
or U1974 (N_1974,In_526,In_2731);
nor U1975 (N_1975,In_2798,In_2162);
or U1976 (N_1976,In_942,In_1589);
xnor U1977 (N_1977,In_2521,In_2339);
nand U1978 (N_1978,In_1552,In_1875);
xnor U1979 (N_1979,In_2247,In_743);
and U1980 (N_1980,In_1362,In_2306);
nand U1981 (N_1981,In_483,In_1691);
nand U1982 (N_1982,In_887,In_1552);
or U1983 (N_1983,In_193,In_1541);
nand U1984 (N_1984,In_1618,In_2380);
xnor U1985 (N_1985,In_1643,In_333);
xor U1986 (N_1986,In_2553,In_2934);
nor U1987 (N_1987,In_844,In_19);
nor U1988 (N_1988,In_2911,In_216);
or U1989 (N_1989,In_1127,In_234);
and U1990 (N_1990,In_1542,In_2676);
nand U1991 (N_1991,In_78,In_1329);
and U1992 (N_1992,In_2782,In_1738);
and U1993 (N_1993,In_1839,In_611);
nand U1994 (N_1994,In_1135,In_1485);
or U1995 (N_1995,In_2493,In_2004);
and U1996 (N_1996,In_362,In_650);
nor U1997 (N_1997,In_982,In_1664);
xor U1998 (N_1998,In_561,In_483);
nand U1999 (N_1999,In_2416,In_2005);
nor U2000 (N_2000,In_1468,In_165);
nor U2001 (N_2001,In_2343,In_851);
nor U2002 (N_2002,In_427,In_955);
nand U2003 (N_2003,In_230,In_538);
or U2004 (N_2004,In_906,In_602);
nand U2005 (N_2005,In_818,In_1837);
nor U2006 (N_2006,In_351,In_2067);
nand U2007 (N_2007,In_122,In_332);
nand U2008 (N_2008,In_208,In_1784);
nand U2009 (N_2009,In_2752,In_2875);
nor U2010 (N_2010,In_2380,In_1702);
and U2011 (N_2011,In_2878,In_1130);
or U2012 (N_2012,In_46,In_2920);
nor U2013 (N_2013,In_2548,In_615);
nand U2014 (N_2014,In_2217,In_1362);
and U2015 (N_2015,In_85,In_1015);
nor U2016 (N_2016,In_1728,In_655);
and U2017 (N_2017,In_1159,In_1646);
or U2018 (N_2018,In_186,In_394);
and U2019 (N_2019,In_651,In_2549);
nor U2020 (N_2020,In_1624,In_1196);
or U2021 (N_2021,In_2293,In_1492);
xnor U2022 (N_2022,In_1428,In_784);
or U2023 (N_2023,In_1820,In_1651);
nor U2024 (N_2024,In_1536,In_2897);
nor U2025 (N_2025,In_2482,In_1908);
xnor U2026 (N_2026,In_1890,In_2493);
nor U2027 (N_2027,In_2689,In_1674);
nor U2028 (N_2028,In_189,In_1174);
and U2029 (N_2029,In_2144,In_734);
nor U2030 (N_2030,In_2747,In_1375);
nand U2031 (N_2031,In_2787,In_1112);
or U2032 (N_2032,In_1034,In_1243);
nand U2033 (N_2033,In_708,In_926);
or U2034 (N_2034,In_1610,In_2156);
or U2035 (N_2035,In_2293,In_1730);
and U2036 (N_2036,In_2336,In_2824);
nor U2037 (N_2037,In_1527,In_1976);
and U2038 (N_2038,In_1708,In_1695);
or U2039 (N_2039,In_2079,In_1730);
nor U2040 (N_2040,In_2140,In_1405);
nor U2041 (N_2041,In_809,In_1791);
and U2042 (N_2042,In_1143,In_1037);
xor U2043 (N_2043,In_1749,In_1645);
and U2044 (N_2044,In_1521,In_2455);
and U2045 (N_2045,In_1459,In_2397);
xnor U2046 (N_2046,In_2753,In_258);
or U2047 (N_2047,In_1247,In_386);
or U2048 (N_2048,In_661,In_2803);
nand U2049 (N_2049,In_793,In_292);
nor U2050 (N_2050,In_545,In_1794);
or U2051 (N_2051,In_2714,In_91);
or U2052 (N_2052,In_756,In_2628);
nor U2053 (N_2053,In_2952,In_2298);
or U2054 (N_2054,In_258,In_1399);
nand U2055 (N_2055,In_1056,In_1735);
nor U2056 (N_2056,In_628,In_1421);
or U2057 (N_2057,In_2997,In_1385);
xor U2058 (N_2058,In_2146,In_2963);
or U2059 (N_2059,In_2241,In_2978);
nor U2060 (N_2060,In_1598,In_86);
nand U2061 (N_2061,In_2050,In_2130);
nor U2062 (N_2062,In_2797,In_1460);
or U2063 (N_2063,In_1807,In_1521);
or U2064 (N_2064,In_2127,In_2465);
nor U2065 (N_2065,In_2266,In_864);
nand U2066 (N_2066,In_1641,In_29);
nand U2067 (N_2067,In_839,In_1522);
or U2068 (N_2068,In_771,In_5);
nor U2069 (N_2069,In_2783,In_1785);
nor U2070 (N_2070,In_2506,In_1636);
and U2071 (N_2071,In_434,In_1382);
nand U2072 (N_2072,In_1229,In_2901);
nand U2073 (N_2073,In_2698,In_235);
or U2074 (N_2074,In_319,In_2927);
nand U2075 (N_2075,In_2132,In_1505);
xor U2076 (N_2076,In_2014,In_1649);
and U2077 (N_2077,In_2888,In_2457);
or U2078 (N_2078,In_2133,In_1067);
nor U2079 (N_2079,In_2111,In_1473);
nor U2080 (N_2080,In_2491,In_1455);
nor U2081 (N_2081,In_2467,In_654);
nor U2082 (N_2082,In_200,In_1084);
nor U2083 (N_2083,In_1730,In_509);
nor U2084 (N_2084,In_1800,In_1310);
nor U2085 (N_2085,In_1647,In_597);
and U2086 (N_2086,In_2080,In_74);
nand U2087 (N_2087,In_1786,In_2430);
nor U2088 (N_2088,In_1399,In_303);
xor U2089 (N_2089,In_921,In_1899);
or U2090 (N_2090,In_54,In_1391);
and U2091 (N_2091,In_2799,In_1861);
or U2092 (N_2092,In_1610,In_1141);
nor U2093 (N_2093,In_557,In_2712);
nand U2094 (N_2094,In_1112,In_1760);
xnor U2095 (N_2095,In_1533,In_2397);
and U2096 (N_2096,In_2836,In_2097);
and U2097 (N_2097,In_844,In_2082);
and U2098 (N_2098,In_1776,In_1936);
xor U2099 (N_2099,In_1323,In_2198);
nand U2100 (N_2100,In_1632,In_1965);
and U2101 (N_2101,In_2980,In_2837);
and U2102 (N_2102,In_1059,In_1695);
xnor U2103 (N_2103,In_668,In_756);
or U2104 (N_2104,In_1564,In_1518);
nor U2105 (N_2105,In_2881,In_1058);
or U2106 (N_2106,In_2225,In_185);
and U2107 (N_2107,In_896,In_118);
nand U2108 (N_2108,In_2317,In_1073);
nand U2109 (N_2109,In_2176,In_1284);
or U2110 (N_2110,In_2438,In_1757);
nand U2111 (N_2111,In_859,In_889);
or U2112 (N_2112,In_2153,In_2555);
nor U2113 (N_2113,In_463,In_2826);
xor U2114 (N_2114,In_1503,In_21);
or U2115 (N_2115,In_1857,In_2364);
xnor U2116 (N_2116,In_2725,In_2917);
or U2117 (N_2117,In_126,In_2937);
and U2118 (N_2118,In_2234,In_11);
nor U2119 (N_2119,In_2414,In_2956);
or U2120 (N_2120,In_2236,In_1342);
nor U2121 (N_2121,In_367,In_2122);
nor U2122 (N_2122,In_1646,In_482);
and U2123 (N_2123,In_17,In_2023);
nand U2124 (N_2124,In_783,In_2740);
or U2125 (N_2125,In_1143,In_2991);
or U2126 (N_2126,In_93,In_1050);
nand U2127 (N_2127,In_204,In_1385);
or U2128 (N_2128,In_887,In_980);
nor U2129 (N_2129,In_2482,In_2586);
xor U2130 (N_2130,In_528,In_2214);
nor U2131 (N_2131,In_2261,In_1909);
nand U2132 (N_2132,In_484,In_258);
nand U2133 (N_2133,In_2445,In_440);
or U2134 (N_2134,In_2607,In_1898);
nor U2135 (N_2135,In_1813,In_1427);
nand U2136 (N_2136,In_1632,In_584);
nor U2137 (N_2137,In_2963,In_1256);
and U2138 (N_2138,In_801,In_2013);
and U2139 (N_2139,In_700,In_1963);
nand U2140 (N_2140,In_2672,In_1551);
or U2141 (N_2141,In_1413,In_580);
nand U2142 (N_2142,In_297,In_1236);
or U2143 (N_2143,In_492,In_518);
nand U2144 (N_2144,In_345,In_768);
xnor U2145 (N_2145,In_531,In_2711);
and U2146 (N_2146,In_2,In_58);
or U2147 (N_2147,In_1738,In_2235);
nor U2148 (N_2148,In_999,In_2411);
or U2149 (N_2149,In_2025,In_2983);
or U2150 (N_2150,In_198,In_2801);
and U2151 (N_2151,In_206,In_1565);
nor U2152 (N_2152,In_1170,In_1127);
or U2153 (N_2153,In_1017,In_1495);
nor U2154 (N_2154,In_1800,In_1544);
or U2155 (N_2155,In_857,In_493);
xnor U2156 (N_2156,In_548,In_1635);
nand U2157 (N_2157,In_1234,In_1715);
xnor U2158 (N_2158,In_696,In_1705);
nor U2159 (N_2159,In_1630,In_731);
nor U2160 (N_2160,In_1827,In_2976);
or U2161 (N_2161,In_853,In_1639);
nor U2162 (N_2162,In_709,In_1537);
and U2163 (N_2163,In_2526,In_571);
nand U2164 (N_2164,In_1848,In_1757);
nand U2165 (N_2165,In_1803,In_364);
nor U2166 (N_2166,In_2571,In_960);
nor U2167 (N_2167,In_2745,In_974);
or U2168 (N_2168,In_1675,In_322);
nor U2169 (N_2169,In_898,In_2829);
nor U2170 (N_2170,In_2143,In_1196);
or U2171 (N_2171,In_251,In_863);
nand U2172 (N_2172,In_590,In_1959);
xnor U2173 (N_2173,In_1273,In_1603);
xnor U2174 (N_2174,In_1779,In_2475);
nor U2175 (N_2175,In_700,In_2355);
and U2176 (N_2176,In_599,In_771);
and U2177 (N_2177,In_951,In_198);
and U2178 (N_2178,In_2987,In_967);
nand U2179 (N_2179,In_1196,In_1011);
and U2180 (N_2180,In_1166,In_50);
and U2181 (N_2181,In_267,In_2426);
and U2182 (N_2182,In_962,In_2055);
or U2183 (N_2183,In_2045,In_605);
and U2184 (N_2184,In_491,In_1566);
or U2185 (N_2185,In_2586,In_1793);
nand U2186 (N_2186,In_1528,In_1861);
nand U2187 (N_2187,In_2386,In_310);
and U2188 (N_2188,In_2444,In_274);
and U2189 (N_2189,In_2391,In_347);
and U2190 (N_2190,In_2553,In_658);
or U2191 (N_2191,In_869,In_2974);
nor U2192 (N_2192,In_2470,In_2871);
xor U2193 (N_2193,In_2184,In_283);
nand U2194 (N_2194,In_2499,In_2828);
nand U2195 (N_2195,In_1591,In_2511);
nand U2196 (N_2196,In_564,In_2815);
nor U2197 (N_2197,In_399,In_301);
nand U2198 (N_2198,In_1752,In_2805);
and U2199 (N_2199,In_2734,In_1127);
nor U2200 (N_2200,In_1735,In_1894);
and U2201 (N_2201,In_578,In_1654);
and U2202 (N_2202,In_2737,In_2034);
nor U2203 (N_2203,In_1447,In_2146);
and U2204 (N_2204,In_1897,In_81);
and U2205 (N_2205,In_403,In_2284);
xor U2206 (N_2206,In_2317,In_202);
or U2207 (N_2207,In_2215,In_2860);
nand U2208 (N_2208,In_1365,In_2418);
nand U2209 (N_2209,In_1892,In_375);
nor U2210 (N_2210,In_539,In_1448);
nor U2211 (N_2211,In_256,In_1314);
nor U2212 (N_2212,In_1867,In_1264);
and U2213 (N_2213,In_1012,In_2821);
or U2214 (N_2214,In_1763,In_513);
nor U2215 (N_2215,In_2627,In_2323);
nand U2216 (N_2216,In_1474,In_1538);
nand U2217 (N_2217,In_1008,In_520);
or U2218 (N_2218,In_1790,In_2903);
nand U2219 (N_2219,In_44,In_2266);
nand U2220 (N_2220,In_222,In_432);
nor U2221 (N_2221,In_515,In_651);
nand U2222 (N_2222,In_1569,In_777);
nor U2223 (N_2223,In_1903,In_73);
or U2224 (N_2224,In_1382,In_716);
nand U2225 (N_2225,In_2067,In_524);
nand U2226 (N_2226,In_2147,In_1296);
and U2227 (N_2227,In_1601,In_1449);
xor U2228 (N_2228,In_968,In_2207);
xnor U2229 (N_2229,In_891,In_2931);
and U2230 (N_2230,In_551,In_352);
or U2231 (N_2231,In_843,In_2127);
nand U2232 (N_2232,In_1618,In_832);
nand U2233 (N_2233,In_452,In_24);
and U2234 (N_2234,In_1839,In_1751);
or U2235 (N_2235,In_2038,In_1870);
nor U2236 (N_2236,In_2722,In_1041);
or U2237 (N_2237,In_130,In_941);
nand U2238 (N_2238,In_2485,In_2153);
nor U2239 (N_2239,In_1311,In_1262);
or U2240 (N_2240,In_294,In_2973);
nor U2241 (N_2241,In_2746,In_1906);
or U2242 (N_2242,In_2832,In_2551);
nor U2243 (N_2243,In_1586,In_2845);
xnor U2244 (N_2244,In_2078,In_1311);
xnor U2245 (N_2245,In_2623,In_2538);
and U2246 (N_2246,In_734,In_923);
xnor U2247 (N_2247,In_2188,In_1177);
and U2248 (N_2248,In_1511,In_769);
nor U2249 (N_2249,In_1164,In_835);
nor U2250 (N_2250,In_1313,In_1276);
or U2251 (N_2251,In_1829,In_2292);
or U2252 (N_2252,In_2703,In_2359);
nand U2253 (N_2253,In_2554,In_2040);
or U2254 (N_2254,In_2064,In_1729);
nand U2255 (N_2255,In_1793,In_1967);
nand U2256 (N_2256,In_1184,In_1232);
nor U2257 (N_2257,In_386,In_1157);
and U2258 (N_2258,In_270,In_2549);
or U2259 (N_2259,In_880,In_1744);
nor U2260 (N_2260,In_1255,In_1821);
and U2261 (N_2261,In_2609,In_537);
and U2262 (N_2262,In_708,In_2553);
or U2263 (N_2263,In_2876,In_456);
nor U2264 (N_2264,In_456,In_1849);
nand U2265 (N_2265,In_1089,In_387);
or U2266 (N_2266,In_2232,In_379);
nand U2267 (N_2267,In_410,In_2988);
and U2268 (N_2268,In_1255,In_48);
and U2269 (N_2269,In_2726,In_2554);
nor U2270 (N_2270,In_604,In_1787);
or U2271 (N_2271,In_1740,In_133);
or U2272 (N_2272,In_1390,In_2123);
nand U2273 (N_2273,In_1212,In_601);
nand U2274 (N_2274,In_597,In_1972);
nand U2275 (N_2275,In_644,In_1693);
nor U2276 (N_2276,In_2037,In_2241);
nand U2277 (N_2277,In_49,In_72);
and U2278 (N_2278,In_999,In_114);
or U2279 (N_2279,In_1635,In_2028);
nand U2280 (N_2280,In_2099,In_311);
xor U2281 (N_2281,In_1592,In_1538);
or U2282 (N_2282,In_232,In_2930);
and U2283 (N_2283,In_2390,In_1951);
nor U2284 (N_2284,In_2314,In_1164);
xor U2285 (N_2285,In_411,In_605);
and U2286 (N_2286,In_1683,In_454);
and U2287 (N_2287,In_939,In_2281);
nor U2288 (N_2288,In_160,In_1693);
nand U2289 (N_2289,In_1130,In_462);
and U2290 (N_2290,In_1723,In_912);
xnor U2291 (N_2291,In_2111,In_828);
nor U2292 (N_2292,In_1685,In_1294);
or U2293 (N_2293,In_77,In_980);
and U2294 (N_2294,In_1808,In_625);
and U2295 (N_2295,In_1693,In_2578);
nor U2296 (N_2296,In_1644,In_211);
nor U2297 (N_2297,In_794,In_111);
and U2298 (N_2298,In_2462,In_2830);
xor U2299 (N_2299,In_1601,In_1605);
nand U2300 (N_2300,In_1337,In_1095);
and U2301 (N_2301,In_649,In_1238);
nor U2302 (N_2302,In_2323,In_1263);
xnor U2303 (N_2303,In_2289,In_1257);
nor U2304 (N_2304,In_669,In_746);
nand U2305 (N_2305,In_595,In_2854);
and U2306 (N_2306,In_299,In_639);
nand U2307 (N_2307,In_1435,In_67);
and U2308 (N_2308,In_476,In_393);
nor U2309 (N_2309,In_1132,In_693);
or U2310 (N_2310,In_948,In_1017);
and U2311 (N_2311,In_1967,In_2946);
or U2312 (N_2312,In_1705,In_1664);
nand U2313 (N_2313,In_1059,In_2972);
or U2314 (N_2314,In_802,In_454);
xnor U2315 (N_2315,In_346,In_987);
nand U2316 (N_2316,In_2790,In_287);
or U2317 (N_2317,In_336,In_980);
xnor U2318 (N_2318,In_974,In_2460);
nand U2319 (N_2319,In_578,In_89);
and U2320 (N_2320,In_116,In_2471);
and U2321 (N_2321,In_1971,In_2214);
nand U2322 (N_2322,In_2014,In_2686);
or U2323 (N_2323,In_613,In_2932);
xnor U2324 (N_2324,In_1452,In_1934);
nand U2325 (N_2325,In_1968,In_2228);
and U2326 (N_2326,In_2148,In_1738);
or U2327 (N_2327,In_2012,In_2563);
nand U2328 (N_2328,In_1994,In_1078);
nand U2329 (N_2329,In_1113,In_2833);
and U2330 (N_2330,In_1111,In_1931);
nand U2331 (N_2331,In_1623,In_744);
nand U2332 (N_2332,In_2218,In_1438);
and U2333 (N_2333,In_2604,In_2858);
or U2334 (N_2334,In_1981,In_1784);
xor U2335 (N_2335,In_1304,In_1649);
or U2336 (N_2336,In_984,In_2026);
or U2337 (N_2337,In_2874,In_1032);
and U2338 (N_2338,In_279,In_1012);
nand U2339 (N_2339,In_1426,In_1956);
or U2340 (N_2340,In_1531,In_1760);
and U2341 (N_2341,In_1521,In_2757);
nor U2342 (N_2342,In_2377,In_661);
nor U2343 (N_2343,In_2974,In_204);
and U2344 (N_2344,In_472,In_2613);
nand U2345 (N_2345,In_304,In_2143);
nor U2346 (N_2346,In_2128,In_1566);
nand U2347 (N_2347,In_2017,In_492);
and U2348 (N_2348,In_578,In_514);
nand U2349 (N_2349,In_865,In_1909);
nand U2350 (N_2350,In_2235,In_1106);
nor U2351 (N_2351,In_2677,In_1554);
nand U2352 (N_2352,In_340,In_2300);
nor U2353 (N_2353,In_1604,In_1626);
nand U2354 (N_2354,In_111,In_2541);
nor U2355 (N_2355,In_1380,In_720);
and U2356 (N_2356,In_401,In_2211);
nand U2357 (N_2357,In_2664,In_2494);
nand U2358 (N_2358,In_2934,In_2686);
nor U2359 (N_2359,In_1668,In_571);
and U2360 (N_2360,In_2402,In_1268);
nand U2361 (N_2361,In_1473,In_2632);
or U2362 (N_2362,In_1829,In_711);
nand U2363 (N_2363,In_2272,In_1471);
nand U2364 (N_2364,In_2143,In_1869);
nand U2365 (N_2365,In_44,In_25);
nor U2366 (N_2366,In_2863,In_1149);
nand U2367 (N_2367,In_1138,In_2678);
and U2368 (N_2368,In_1161,In_2465);
nand U2369 (N_2369,In_2181,In_1909);
xnor U2370 (N_2370,In_313,In_1108);
nand U2371 (N_2371,In_954,In_1552);
nor U2372 (N_2372,In_126,In_2890);
nand U2373 (N_2373,In_1715,In_2395);
and U2374 (N_2374,In_1842,In_1860);
or U2375 (N_2375,In_1617,In_2746);
or U2376 (N_2376,In_258,In_1311);
or U2377 (N_2377,In_2281,In_2339);
nor U2378 (N_2378,In_2803,In_2069);
nand U2379 (N_2379,In_2822,In_2037);
or U2380 (N_2380,In_47,In_1789);
nor U2381 (N_2381,In_2112,In_127);
or U2382 (N_2382,In_1861,In_2871);
nor U2383 (N_2383,In_2660,In_1385);
or U2384 (N_2384,In_731,In_1812);
or U2385 (N_2385,In_2506,In_1180);
or U2386 (N_2386,In_2286,In_2873);
nand U2387 (N_2387,In_2488,In_493);
or U2388 (N_2388,In_2834,In_380);
nand U2389 (N_2389,In_1363,In_2315);
or U2390 (N_2390,In_462,In_1299);
nor U2391 (N_2391,In_53,In_2404);
xor U2392 (N_2392,In_2477,In_957);
and U2393 (N_2393,In_1536,In_1129);
or U2394 (N_2394,In_2091,In_2611);
xnor U2395 (N_2395,In_1908,In_2420);
nor U2396 (N_2396,In_2632,In_2427);
nand U2397 (N_2397,In_630,In_390);
xor U2398 (N_2398,In_888,In_1940);
nand U2399 (N_2399,In_2009,In_451);
or U2400 (N_2400,In_2446,In_501);
nor U2401 (N_2401,In_2216,In_2409);
and U2402 (N_2402,In_1541,In_1774);
or U2403 (N_2403,In_1769,In_276);
or U2404 (N_2404,In_256,In_238);
nor U2405 (N_2405,In_1694,In_2636);
xnor U2406 (N_2406,In_650,In_276);
xnor U2407 (N_2407,In_44,In_928);
or U2408 (N_2408,In_1175,In_1699);
nor U2409 (N_2409,In_2090,In_2543);
and U2410 (N_2410,In_928,In_1205);
nand U2411 (N_2411,In_1052,In_1698);
or U2412 (N_2412,In_651,In_2852);
or U2413 (N_2413,In_137,In_1969);
and U2414 (N_2414,In_2763,In_2925);
nand U2415 (N_2415,In_1122,In_816);
nand U2416 (N_2416,In_1753,In_599);
xor U2417 (N_2417,In_2182,In_1612);
and U2418 (N_2418,In_2989,In_1487);
and U2419 (N_2419,In_2082,In_2539);
or U2420 (N_2420,In_133,In_1849);
and U2421 (N_2421,In_2020,In_2172);
xor U2422 (N_2422,In_2921,In_1034);
xnor U2423 (N_2423,In_665,In_871);
and U2424 (N_2424,In_2341,In_296);
nor U2425 (N_2425,In_1267,In_2641);
or U2426 (N_2426,In_499,In_15);
nor U2427 (N_2427,In_1312,In_35);
nand U2428 (N_2428,In_2263,In_1277);
and U2429 (N_2429,In_632,In_91);
nor U2430 (N_2430,In_1322,In_2064);
nor U2431 (N_2431,In_1930,In_966);
nor U2432 (N_2432,In_2489,In_456);
and U2433 (N_2433,In_1501,In_2893);
and U2434 (N_2434,In_685,In_2997);
or U2435 (N_2435,In_20,In_197);
xnor U2436 (N_2436,In_2750,In_2181);
and U2437 (N_2437,In_2549,In_2390);
xor U2438 (N_2438,In_2160,In_1564);
and U2439 (N_2439,In_847,In_2968);
and U2440 (N_2440,In_1836,In_978);
or U2441 (N_2441,In_1181,In_1223);
nand U2442 (N_2442,In_1071,In_1027);
xnor U2443 (N_2443,In_2479,In_1490);
nand U2444 (N_2444,In_2712,In_741);
nor U2445 (N_2445,In_1063,In_2165);
xnor U2446 (N_2446,In_2645,In_2851);
or U2447 (N_2447,In_124,In_70);
nand U2448 (N_2448,In_295,In_970);
nor U2449 (N_2449,In_1200,In_2358);
xor U2450 (N_2450,In_19,In_498);
xor U2451 (N_2451,In_1466,In_1339);
nand U2452 (N_2452,In_2616,In_1556);
nand U2453 (N_2453,In_775,In_1664);
nand U2454 (N_2454,In_505,In_541);
xor U2455 (N_2455,In_1403,In_244);
xor U2456 (N_2456,In_1956,In_1626);
xnor U2457 (N_2457,In_1590,In_1812);
or U2458 (N_2458,In_2734,In_931);
nor U2459 (N_2459,In_1912,In_2168);
and U2460 (N_2460,In_2287,In_292);
nand U2461 (N_2461,In_1305,In_2912);
or U2462 (N_2462,In_875,In_1886);
xnor U2463 (N_2463,In_1340,In_2557);
and U2464 (N_2464,In_323,In_2774);
and U2465 (N_2465,In_498,In_2830);
nand U2466 (N_2466,In_835,In_829);
or U2467 (N_2467,In_2477,In_2439);
or U2468 (N_2468,In_2062,In_2281);
or U2469 (N_2469,In_1152,In_1757);
nor U2470 (N_2470,In_987,In_563);
or U2471 (N_2471,In_160,In_598);
and U2472 (N_2472,In_1289,In_2244);
and U2473 (N_2473,In_768,In_2484);
xor U2474 (N_2474,In_7,In_2488);
nand U2475 (N_2475,In_1368,In_2363);
or U2476 (N_2476,In_1872,In_2295);
xor U2477 (N_2477,In_1626,In_298);
nor U2478 (N_2478,In_945,In_2482);
and U2479 (N_2479,In_2626,In_2345);
and U2480 (N_2480,In_995,In_2695);
nor U2481 (N_2481,In_2895,In_197);
nand U2482 (N_2482,In_1559,In_1219);
and U2483 (N_2483,In_2828,In_1979);
nand U2484 (N_2484,In_1384,In_2665);
xor U2485 (N_2485,In_2480,In_795);
and U2486 (N_2486,In_233,In_1740);
nand U2487 (N_2487,In_2350,In_1316);
and U2488 (N_2488,In_394,In_1667);
nand U2489 (N_2489,In_1942,In_1342);
or U2490 (N_2490,In_2555,In_1140);
xor U2491 (N_2491,In_1787,In_857);
nor U2492 (N_2492,In_1451,In_831);
and U2493 (N_2493,In_2551,In_2899);
nand U2494 (N_2494,In_1819,In_1710);
and U2495 (N_2495,In_751,In_97);
or U2496 (N_2496,In_26,In_1890);
or U2497 (N_2497,In_2754,In_1018);
nor U2498 (N_2498,In_2866,In_1809);
or U2499 (N_2499,In_8,In_1829);
or U2500 (N_2500,In_329,In_2318);
nor U2501 (N_2501,In_961,In_615);
or U2502 (N_2502,In_1122,In_1333);
or U2503 (N_2503,In_420,In_1150);
or U2504 (N_2504,In_1965,In_1737);
and U2505 (N_2505,In_2740,In_503);
xnor U2506 (N_2506,In_2127,In_614);
nand U2507 (N_2507,In_1238,In_740);
nor U2508 (N_2508,In_2414,In_673);
nor U2509 (N_2509,In_1128,In_80);
nand U2510 (N_2510,In_61,In_2960);
and U2511 (N_2511,In_1400,In_2563);
or U2512 (N_2512,In_2761,In_1745);
or U2513 (N_2513,In_2236,In_2749);
nand U2514 (N_2514,In_1699,In_2039);
nand U2515 (N_2515,In_180,In_2298);
and U2516 (N_2516,In_888,In_2483);
xor U2517 (N_2517,In_2673,In_637);
and U2518 (N_2518,In_604,In_2047);
and U2519 (N_2519,In_2222,In_2052);
nand U2520 (N_2520,In_1914,In_465);
and U2521 (N_2521,In_1142,In_591);
nand U2522 (N_2522,In_2019,In_1139);
nor U2523 (N_2523,In_90,In_1695);
or U2524 (N_2524,In_384,In_2156);
and U2525 (N_2525,In_1383,In_683);
xnor U2526 (N_2526,In_1846,In_458);
xnor U2527 (N_2527,In_1072,In_561);
and U2528 (N_2528,In_1398,In_499);
nand U2529 (N_2529,In_1141,In_333);
and U2530 (N_2530,In_1955,In_1870);
nand U2531 (N_2531,In_2973,In_1083);
nand U2532 (N_2532,In_1829,In_2318);
nor U2533 (N_2533,In_1888,In_1452);
nand U2534 (N_2534,In_576,In_1095);
nand U2535 (N_2535,In_2019,In_1345);
and U2536 (N_2536,In_2586,In_2679);
and U2537 (N_2537,In_727,In_119);
and U2538 (N_2538,In_824,In_483);
or U2539 (N_2539,In_2500,In_1966);
nor U2540 (N_2540,In_2972,In_1435);
or U2541 (N_2541,In_2085,In_1226);
nand U2542 (N_2542,In_804,In_655);
nor U2543 (N_2543,In_73,In_2708);
nor U2544 (N_2544,In_5,In_1164);
or U2545 (N_2545,In_1358,In_829);
nand U2546 (N_2546,In_242,In_763);
and U2547 (N_2547,In_2731,In_2765);
or U2548 (N_2548,In_918,In_716);
xor U2549 (N_2549,In_2674,In_972);
xor U2550 (N_2550,In_1806,In_395);
or U2551 (N_2551,In_2035,In_768);
or U2552 (N_2552,In_1178,In_167);
and U2553 (N_2553,In_2577,In_2444);
nor U2554 (N_2554,In_2375,In_2758);
nand U2555 (N_2555,In_2202,In_43);
or U2556 (N_2556,In_725,In_1675);
and U2557 (N_2557,In_1930,In_2099);
nand U2558 (N_2558,In_568,In_1427);
nor U2559 (N_2559,In_2035,In_710);
and U2560 (N_2560,In_836,In_2751);
or U2561 (N_2561,In_2976,In_469);
or U2562 (N_2562,In_2274,In_1779);
xnor U2563 (N_2563,In_1812,In_1947);
nand U2564 (N_2564,In_2039,In_2544);
nor U2565 (N_2565,In_1678,In_2825);
and U2566 (N_2566,In_2232,In_1028);
nand U2567 (N_2567,In_2820,In_1865);
or U2568 (N_2568,In_194,In_624);
nand U2569 (N_2569,In_1531,In_470);
nor U2570 (N_2570,In_2366,In_194);
or U2571 (N_2571,In_1539,In_2513);
nand U2572 (N_2572,In_1907,In_1321);
nand U2573 (N_2573,In_2933,In_1249);
and U2574 (N_2574,In_1248,In_1092);
xor U2575 (N_2575,In_2720,In_1246);
and U2576 (N_2576,In_2438,In_1386);
and U2577 (N_2577,In_119,In_2814);
or U2578 (N_2578,In_1699,In_1866);
nor U2579 (N_2579,In_2460,In_2976);
nand U2580 (N_2580,In_1676,In_752);
and U2581 (N_2581,In_1301,In_1495);
or U2582 (N_2582,In_1278,In_719);
nand U2583 (N_2583,In_2898,In_2073);
and U2584 (N_2584,In_202,In_2186);
and U2585 (N_2585,In_2536,In_2563);
nor U2586 (N_2586,In_2907,In_1735);
and U2587 (N_2587,In_591,In_632);
or U2588 (N_2588,In_2540,In_2408);
nor U2589 (N_2589,In_215,In_2755);
xor U2590 (N_2590,In_1288,In_2520);
and U2591 (N_2591,In_2797,In_1495);
nand U2592 (N_2592,In_1118,In_2031);
nand U2593 (N_2593,In_2799,In_1406);
or U2594 (N_2594,In_738,In_2227);
nand U2595 (N_2595,In_1303,In_129);
nand U2596 (N_2596,In_2403,In_1716);
nand U2597 (N_2597,In_2382,In_1571);
or U2598 (N_2598,In_87,In_1030);
nor U2599 (N_2599,In_1221,In_490);
nor U2600 (N_2600,In_2094,In_764);
nor U2601 (N_2601,In_2618,In_2043);
or U2602 (N_2602,In_1430,In_2753);
nor U2603 (N_2603,In_1384,In_2300);
and U2604 (N_2604,In_1583,In_2937);
and U2605 (N_2605,In_1350,In_1795);
or U2606 (N_2606,In_2028,In_1916);
and U2607 (N_2607,In_2979,In_1371);
nor U2608 (N_2608,In_668,In_1715);
or U2609 (N_2609,In_1216,In_1834);
nand U2610 (N_2610,In_2139,In_2453);
or U2611 (N_2611,In_1940,In_2918);
and U2612 (N_2612,In_1414,In_615);
nor U2613 (N_2613,In_1382,In_1365);
xnor U2614 (N_2614,In_794,In_1897);
or U2615 (N_2615,In_1990,In_1732);
xor U2616 (N_2616,In_1634,In_2345);
and U2617 (N_2617,In_922,In_382);
or U2618 (N_2618,In_1303,In_1540);
xor U2619 (N_2619,In_401,In_1719);
and U2620 (N_2620,In_558,In_1500);
and U2621 (N_2621,In_1799,In_2567);
and U2622 (N_2622,In_1426,In_1138);
or U2623 (N_2623,In_1419,In_2264);
or U2624 (N_2624,In_1929,In_23);
nand U2625 (N_2625,In_319,In_2190);
or U2626 (N_2626,In_2663,In_887);
or U2627 (N_2627,In_2155,In_296);
xnor U2628 (N_2628,In_284,In_2030);
nand U2629 (N_2629,In_867,In_2081);
nor U2630 (N_2630,In_377,In_1601);
xnor U2631 (N_2631,In_2710,In_2046);
and U2632 (N_2632,In_443,In_271);
xor U2633 (N_2633,In_2533,In_1051);
nand U2634 (N_2634,In_1120,In_2365);
nand U2635 (N_2635,In_2563,In_2108);
xor U2636 (N_2636,In_2364,In_2820);
and U2637 (N_2637,In_2998,In_2412);
nor U2638 (N_2638,In_2154,In_1287);
xor U2639 (N_2639,In_1726,In_750);
nand U2640 (N_2640,In_1037,In_1033);
xor U2641 (N_2641,In_1973,In_1340);
nor U2642 (N_2642,In_1514,In_2977);
or U2643 (N_2643,In_2924,In_1897);
nor U2644 (N_2644,In_2741,In_1830);
xnor U2645 (N_2645,In_1160,In_2338);
xor U2646 (N_2646,In_2525,In_1116);
or U2647 (N_2647,In_2193,In_324);
xor U2648 (N_2648,In_2479,In_2316);
or U2649 (N_2649,In_55,In_1288);
and U2650 (N_2650,In_704,In_1717);
and U2651 (N_2651,In_484,In_478);
xor U2652 (N_2652,In_1763,In_2169);
and U2653 (N_2653,In_2132,In_452);
nand U2654 (N_2654,In_1794,In_920);
nor U2655 (N_2655,In_1334,In_2551);
and U2656 (N_2656,In_2516,In_1706);
or U2657 (N_2657,In_304,In_2596);
and U2658 (N_2658,In_2514,In_2848);
or U2659 (N_2659,In_246,In_1246);
and U2660 (N_2660,In_1333,In_253);
or U2661 (N_2661,In_2715,In_1035);
nor U2662 (N_2662,In_1378,In_1673);
nand U2663 (N_2663,In_23,In_2570);
xnor U2664 (N_2664,In_2066,In_1886);
and U2665 (N_2665,In_2294,In_47);
xnor U2666 (N_2666,In_1631,In_2559);
and U2667 (N_2667,In_1505,In_111);
or U2668 (N_2668,In_1735,In_2447);
nand U2669 (N_2669,In_2087,In_1158);
or U2670 (N_2670,In_2800,In_1258);
xnor U2671 (N_2671,In_1545,In_1888);
or U2672 (N_2672,In_1689,In_1647);
nand U2673 (N_2673,In_2964,In_581);
nor U2674 (N_2674,In_597,In_2368);
and U2675 (N_2675,In_502,In_1796);
and U2676 (N_2676,In_2284,In_332);
nand U2677 (N_2677,In_571,In_25);
and U2678 (N_2678,In_1494,In_1456);
and U2679 (N_2679,In_41,In_2789);
or U2680 (N_2680,In_2910,In_1979);
nor U2681 (N_2681,In_1588,In_1142);
or U2682 (N_2682,In_2232,In_791);
and U2683 (N_2683,In_2643,In_256);
nand U2684 (N_2684,In_2440,In_1677);
and U2685 (N_2685,In_896,In_1535);
and U2686 (N_2686,In_768,In_323);
and U2687 (N_2687,In_1036,In_2041);
and U2688 (N_2688,In_471,In_2771);
or U2689 (N_2689,In_874,In_2394);
or U2690 (N_2690,In_1516,In_2130);
xnor U2691 (N_2691,In_2458,In_2056);
and U2692 (N_2692,In_2795,In_1484);
nand U2693 (N_2693,In_1780,In_1553);
xnor U2694 (N_2694,In_2666,In_1812);
nand U2695 (N_2695,In_778,In_6);
and U2696 (N_2696,In_713,In_2618);
nor U2697 (N_2697,In_1410,In_1291);
nand U2698 (N_2698,In_2122,In_2833);
nand U2699 (N_2699,In_1224,In_1738);
and U2700 (N_2700,In_1861,In_448);
and U2701 (N_2701,In_79,In_2552);
nor U2702 (N_2702,In_1832,In_1833);
nor U2703 (N_2703,In_315,In_950);
or U2704 (N_2704,In_2911,In_2025);
xor U2705 (N_2705,In_1800,In_1333);
xnor U2706 (N_2706,In_190,In_1552);
nor U2707 (N_2707,In_2349,In_1147);
nor U2708 (N_2708,In_1771,In_1487);
nor U2709 (N_2709,In_1858,In_1237);
nor U2710 (N_2710,In_250,In_614);
or U2711 (N_2711,In_426,In_370);
or U2712 (N_2712,In_1129,In_2761);
nand U2713 (N_2713,In_1182,In_579);
nor U2714 (N_2714,In_1646,In_1532);
nand U2715 (N_2715,In_2644,In_1508);
or U2716 (N_2716,In_866,In_2290);
nor U2717 (N_2717,In_502,In_1139);
or U2718 (N_2718,In_1856,In_563);
nor U2719 (N_2719,In_1984,In_1646);
nand U2720 (N_2720,In_475,In_2131);
nand U2721 (N_2721,In_2400,In_557);
nor U2722 (N_2722,In_88,In_1183);
and U2723 (N_2723,In_375,In_1956);
nand U2724 (N_2724,In_2473,In_1207);
and U2725 (N_2725,In_2200,In_1835);
xor U2726 (N_2726,In_235,In_1635);
and U2727 (N_2727,In_497,In_1437);
or U2728 (N_2728,In_2898,In_2214);
xor U2729 (N_2729,In_2470,In_1585);
nor U2730 (N_2730,In_2964,In_2970);
nor U2731 (N_2731,In_2322,In_1135);
and U2732 (N_2732,In_817,In_1139);
nand U2733 (N_2733,In_2004,In_2810);
and U2734 (N_2734,In_1945,In_985);
nor U2735 (N_2735,In_2909,In_316);
nand U2736 (N_2736,In_2236,In_2768);
or U2737 (N_2737,In_512,In_2671);
nor U2738 (N_2738,In_644,In_2999);
or U2739 (N_2739,In_2943,In_2167);
nor U2740 (N_2740,In_553,In_2053);
nand U2741 (N_2741,In_763,In_2047);
xor U2742 (N_2742,In_2285,In_329);
nor U2743 (N_2743,In_782,In_2470);
and U2744 (N_2744,In_789,In_2927);
nand U2745 (N_2745,In_1730,In_368);
nor U2746 (N_2746,In_1112,In_2688);
and U2747 (N_2747,In_2848,In_1140);
xnor U2748 (N_2748,In_953,In_239);
or U2749 (N_2749,In_2439,In_1127);
nand U2750 (N_2750,In_2286,In_2718);
nor U2751 (N_2751,In_211,In_2705);
and U2752 (N_2752,In_2089,In_382);
xnor U2753 (N_2753,In_1193,In_2022);
nor U2754 (N_2754,In_1312,In_1882);
nand U2755 (N_2755,In_2681,In_2302);
and U2756 (N_2756,In_2296,In_680);
nor U2757 (N_2757,In_753,In_2114);
nand U2758 (N_2758,In_1611,In_2429);
and U2759 (N_2759,In_24,In_2174);
nand U2760 (N_2760,In_817,In_479);
nor U2761 (N_2761,In_1700,In_2933);
nand U2762 (N_2762,In_2551,In_2780);
nand U2763 (N_2763,In_1016,In_2711);
nand U2764 (N_2764,In_2981,In_319);
xor U2765 (N_2765,In_2256,In_130);
xnor U2766 (N_2766,In_1969,In_2119);
nor U2767 (N_2767,In_215,In_2416);
and U2768 (N_2768,In_2905,In_307);
or U2769 (N_2769,In_2774,In_231);
nor U2770 (N_2770,In_1284,In_2839);
nand U2771 (N_2771,In_1335,In_1764);
and U2772 (N_2772,In_653,In_249);
nor U2773 (N_2773,In_1632,In_467);
nor U2774 (N_2774,In_837,In_1097);
xor U2775 (N_2775,In_2154,In_216);
and U2776 (N_2776,In_279,In_121);
nand U2777 (N_2777,In_1489,In_997);
nor U2778 (N_2778,In_2989,In_2543);
or U2779 (N_2779,In_1436,In_2215);
or U2780 (N_2780,In_912,In_1863);
and U2781 (N_2781,In_2267,In_1729);
nor U2782 (N_2782,In_2112,In_95);
and U2783 (N_2783,In_2359,In_287);
nand U2784 (N_2784,In_267,In_2611);
nand U2785 (N_2785,In_1414,In_2913);
nand U2786 (N_2786,In_1786,In_2835);
xnor U2787 (N_2787,In_204,In_2765);
nand U2788 (N_2788,In_478,In_1235);
nor U2789 (N_2789,In_225,In_2893);
and U2790 (N_2790,In_52,In_1855);
xor U2791 (N_2791,In_2022,In_65);
or U2792 (N_2792,In_545,In_1363);
nand U2793 (N_2793,In_2056,In_3);
or U2794 (N_2794,In_2301,In_127);
nor U2795 (N_2795,In_348,In_58);
and U2796 (N_2796,In_2004,In_1045);
or U2797 (N_2797,In_2218,In_2071);
nand U2798 (N_2798,In_2315,In_1008);
nor U2799 (N_2799,In_1136,In_2637);
nor U2800 (N_2800,In_731,In_987);
nand U2801 (N_2801,In_1008,In_2424);
nand U2802 (N_2802,In_1935,In_1706);
nor U2803 (N_2803,In_438,In_1873);
nand U2804 (N_2804,In_1366,In_2887);
xor U2805 (N_2805,In_2938,In_170);
nand U2806 (N_2806,In_997,In_589);
or U2807 (N_2807,In_1654,In_2989);
nand U2808 (N_2808,In_463,In_1882);
xor U2809 (N_2809,In_638,In_957);
or U2810 (N_2810,In_332,In_1398);
or U2811 (N_2811,In_2525,In_2212);
and U2812 (N_2812,In_1754,In_2211);
nor U2813 (N_2813,In_58,In_2970);
nor U2814 (N_2814,In_1577,In_1263);
nor U2815 (N_2815,In_2567,In_2852);
or U2816 (N_2816,In_1593,In_2259);
nor U2817 (N_2817,In_883,In_284);
xor U2818 (N_2818,In_772,In_2019);
and U2819 (N_2819,In_2944,In_361);
nand U2820 (N_2820,In_1402,In_1927);
nand U2821 (N_2821,In_956,In_226);
nor U2822 (N_2822,In_231,In_2227);
nand U2823 (N_2823,In_1864,In_2015);
nor U2824 (N_2824,In_2814,In_2766);
nand U2825 (N_2825,In_1046,In_1023);
or U2826 (N_2826,In_1336,In_2714);
nor U2827 (N_2827,In_1927,In_2153);
and U2828 (N_2828,In_321,In_2839);
and U2829 (N_2829,In_2130,In_2172);
and U2830 (N_2830,In_1973,In_2583);
nand U2831 (N_2831,In_2074,In_1956);
or U2832 (N_2832,In_2013,In_1197);
nor U2833 (N_2833,In_1304,In_1573);
or U2834 (N_2834,In_566,In_1661);
and U2835 (N_2835,In_1151,In_2093);
or U2836 (N_2836,In_822,In_2387);
or U2837 (N_2837,In_2579,In_293);
and U2838 (N_2838,In_921,In_366);
nand U2839 (N_2839,In_841,In_428);
nand U2840 (N_2840,In_2193,In_1045);
and U2841 (N_2841,In_165,In_1712);
nand U2842 (N_2842,In_967,In_451);
nand U2843 (N_2843,In_232,In_1484);
or U2844 (N_2844,In_1833,In_2134);
nor U2845 (N_2845,In_2436,In_2554);
and U2846 (N_2846,In_69,In_2461);
nand U2847 (N_2847,In_1407,In_753);
or U2848 (N_2848,In_1866,In_937);
nand U2849 (N_2849,In_470,In_2024);
or U2850 (N_2850,In_2180,In_2021);
nand U2851 (N_2851,In_1750,In_1396);
and U2852 (N_2852,In_894,In_356);
nand U2853 (N_2853,In_2229,In_137);
nor U2854 (N_2854,In_1885,In_97);
and U2855 (N_2855,In_2259,In_1673);
nand U2856 (N_2856,In_1529,In_2793);
or U2857 (N_2857,In_1768,In_1492);
or U2858 (N_2858,In_2989,In_1931);
nor U2859 (N_2859,In_2227,In_425);
xor U2860 (N_2860,In_93,In_349);
and U2861 (N_2861,In_2455,In_960);
or U2862 (N_2862,In_1196,In_939);
xor U2863 (N_2863,In_1750,In_636);
xnor U2864 (N_2864,In_521,In_1425);
and U2865 (N_2865,In_693,In_2903);
nand U2866 (N_2866,In_403,In_1353);
nor U2867 (N_2867,In_1455,In_623);
nand U2868 (N_2868,In_2768,In_984);
or U2869 (N_2869,In_2278,In_2493);
nor U2870 (N_2870,In_942,In_2241);
nand U2871 (N_2871,In_961,In_1620);
nor U2872 (N_2872,In_809,In_2256);
nor U2873 (N_2873,In_2719,In_1335);
and U2874 (N_2874,In_925,In_2481);
or U2875 (N_2875,In_466,In_2418);
xor U2876 (N_2876,In_1274,In_11);
and U2877 (N_2877,In_2944,In_2930);
xnor U2878 (N_2878,In_272,In_677);
nand U2879 (N_2879,In_1839,In_373);
or U2880 (N_2880,In_2046,In_2562);
or U2881 (N_2881,In_1046,In_174);
nor U2882 (N_2882,In_2765,In_631);
nor U2883 (N_2883,In_1438,In_2550);
and U2884 (N_2884,In_2371,In_1876);
or U2885 (N_2885,In_520,In_2589);
nor U2886 (N_2886,In_1653,In_981);
nor U2887 (N_2887,In_2374,In_2602);
nor U2888 (N_2888,In_2058,In_2121);
xor U2889 (N_2889,In_75,In_2887);
nor U2890 (N_2890,In_1816,In_1132);
nand U2891 (N_2891,In_258,In_231);
or U2892 (N_2892,In_2797,In_2485);
nand U2893 (N_2893,In_2415,In_635);
nor U2894 (N_2894,In_1915,In_140);
and U2895 (N_2895,In_2769,In_1355);
nor U2896 (N_2896,In_1869,In_2130);
nor U2897 (N_2897,In_227,In_2136);
xnor U2898 (N_2898,In_1470,In_2406);
nor U2899 (N_2899,In_442,In_2691);
and U2900 (N_2900,In_1599,In_2706);
nand U2901 (N_2901,In_2122,In_2476);
or U2902 (N_2902,In_2095,In_2636);
nor U2903 (N_2903,In_499,In_2244);
xnor U2904 (N_2904,In_176,In_2584);
nand U2905 (N_2905,In_1580,In_1721);
and U2906 (N_2906,In_1512,In_435);
and U2907 (N_2907,In_2378,In_1712);
nand U2908 (N_2908,In_1048,In_2261);
nor U2909 (N_2909,In_2864,In_2353);
nand U2910 (N_2910,In_2158,In_2528);
xor U2911 (N_2911,In_337,In_472);
xor U2912 (N_2912,In_2357,In_1871);
or U2913 (N_2913,In_1683,In_2999);
nand U2914 (N_2914,In_1953,In_1608);
nor U2915 (N_2915,In_1441,In_2031);
and U2916 (N_2916,In_743,In_1840);
nor U2917 (N_2917,In_2567,In_141);
nor U2918 (N_2918,In_843,In_2065);
or U2919 (N_2919,In_2283,In_944);
nand U2920 (N_2920,In_355,In_1668);
xnor U2921 (N_2921,In_2565,In_1841);
nand U2922 (N_2922,In_2907,In_1054);
and U2923 (N_2923,In_779,In_2953);
nand U2924 (N_2924,In_878,In_1394);
xnor U2925 (N_2925,In_1149,In_493);
and U2926 (N_2926,In_673,In_2228);
or U2927 (N_2927,In_1131,In_577);
nand U2928 (N_2928,In_2292,In_47);
nor U2929 (N_2929,In_2139,In_1186);
and U2930 (N_2930,In_2762,In_2645);
nand U2931 (N_2931,In_2438,In_315);
and U2932 (N_2932,In_1135,In_2661);
nand U2933 (N_2933,In_1863,In_2628);
nand U2934 (N_2934,In_173,In_515);
and U2935 (N_2935,In_2354,In_2729);
and U2936 (N_2936,In_2881,In_384);
and U2937 (N_2937,In_1478,In_1074);
and U2938 (N_2938,In_1240,In_811);
and U2939 (N_2939,In_852,In_1860);
or U2940 (N_2940,In_1037,In_405);
and U2941 (N_2941,In_762,In_998);
or U2942 (N_2942,In_640,In_64);
or U2943 (N_2943,In_74,In_612);
and U2944 (N_2944,In_2167,In_413);
and U2945 (N_2945,In_2488,In_2549);
nand U2946 (N_2946,In_757,In_2709);
nor U2947 (N_2947,In_1930,In_2190);
or U2948 (N_2948,In_0,In_1515);
xor U2949 (N_2949,In_270,In_1784);
or U2950 (N_2950,In_1967,In_992);
nand U2951 (N_2951,In_87,In_2643);
nor U2952 (N_2952,In_1478,In_323);
and U2953 (N_2953,In_2743,In_1716);
nor U2954 (N_2954,In_2069,In_752);
xor U2955 (N_2955,In_1006,In_1944);
xnor U2956 (N_2956,In_2382,In_2901);
or U2957 (N_2957,In_1673,In_2614);
nor U2958 (N_2958,In_1702,In_2082);
and U2959 (N_2959,In_2062,In_1123);
xnor U2960 (N_2960,In_2960,In_107);
nor U2961 (N_2961,In_615,In_213);
or U2962 (N_2962,In_1749,In_2438);
nor U2963 (N_2963,In_761,In_1502);
or U2964 (N_2964,In_2968,In_852);
nand U2965 (N_2965,In_2153,In_2852);
or U2966 (N_2966,In_1291,In_1723);
nor U2967 (N_2967,In_879,In_2732);
and U2968 (N_2968,In_445,In_1927);
and U2969 (N_2969,In_2284,In_1095);
and U2970 (N_2970,In_2366,In_379);
and U2971 (N_2971,In_2703,In_1309);
and U2972 (N_2972,In_1052,In_614);
and U2973 (N_2973,In_2919,In_2673);
nand U2974 (N_2974,In_523,In_1559);
nand U2975 (N_2975,In_1927,In_1327);
xor U2976 (N_2976,In_1488,In_8);
nand U2977 (N_2977,In_2625,In_789);
and U2978 (N_2978,In_2313,In_1790);
nor U2979 (N_2979,In_2306,In_2961);
or U2980 (N_2980,In_2062,In_1273);
or U2981 (N_2981,In_2069,In_1244);
nor U2982 (N_2982,In_1979,In_1420);
and U2983 (N_2983,In_2233,In_1243);
xnor U2984 (N_2984,In_1138,In_919);
or U2985 (N_2985,In_2178,In_1337);
and U2986 (N_2986,In_1962,In_2741);
xnor U2987 (N_2987,In_1978,In_2689);
or U2988 (N_2988,In_2905,In_2283);
nand U2989 (N_2989,In_1943,In_1426);
nor U2990 (N_2990,In_788,In_2351);
and U2991 (N_2991,In_643,In_1725);
or U2992 (N_2992,In_2168,In_1101);
xnor U2993 (N_2993,In_2568,In_1680);
and U2994 (N_2994,In_1659,In_1183);
or U2995 (N_2995,In_2609,In_1805);
nor U2996 (N_2996,In_2944,In_530);
nor U2997 (N_2997,In_2039,In_27);
or U2998 (N_2998,In_394,In_2627);
nand U2999 (N_2999,In_93,In_2839);
and U3000 (N_3000,In_1377,In_297);
xor U3001 (N_3001,In_270,In_198);
nor U3002 (N_3002,In_2430,In_747);
and U3003 (N_3003,In_830,In_847);
or U3004 (N_3004,In_2210,In_1566);
nand U3005 (N_3005,In_2181,In_1334);
nor U3006 (N_3006,In_479,In_172);
and U3007 (N_3007,In_2355,In_59);
or U3008 (N_3008,In_2074,In_2901);
nor U3009 (N_3009,In_1821,In_2402);
nor U3010 (N_3010,In_2431,In_2951);
nand U3011 (N_3011,In_450,In_2399);
or U3012 (N_3012,In_2523,In_1600);
nor U3013 (N_3013,In_243,In_2201);
nand U3014 (N_3014,In_59,In_2787);
nand U3015 (N_3015,In_991,In_824);
and U3016 (N_3016,In_1006,In_211);
and U3017 (N_3017,In_806,In_1482);
and U3018 (N_3018,In_1243,In_2564);
nand U3019 (N_3019,In_193,In_341);
or U3020 (N_3020,In_1099,In_2805);
nand U3021 (N_3021,In_1331,In_1601);
nor U3022 (N_3022,In_194,In_2);
and U3023 (N_3023,In_914,In_1249);
nand U3024 (N_3024,In_2968,In_855);
xnor U3025 (N_3025,In_2033,In_797);
xor U3026 (N_3026,In_1299,In_2033);
nor U3027 (N_3027,In_772,In_488);
nand U3028 (N_3028,In_2817,In_494);
and U3029 (N_3029,In_652,In_2028);
or U3030 (N_3030,In_864,In_2755);
nand U3031 (N_3031,In_146,In_281);
or U3032 (N_3032,In_1426,In_1126);
nand U3033 (N_3033,In_774,In_2207);
or U3034 (N_3034,In_414,In_1683);
nand U3035 (N_3035,In_509,In_1276);
and U3036 (N_3036,In_2372,In_1496);
nand U3037 (N_3037,In_1661,In_1233);
or U3038 (N_3038,In_312,In_2128);
nor U3039 (N_3039,In_2606,In_1836);
xnor U3040 (N_3040,In_2212,In_2727);
and U3041 (N_3041,In_10,In_405);
or U3042 (N_3042,In_2291,In_1904);
xnor U3043 (N_3043,In_1082,In_223);
nand U3044 (N_3044,In_2899,In_1912);
or U3045 (N_3045,In_240,In_2614);
xnor U3046 (N_3046,In_819,In_913);
nand U3047 (N_3047,In_227,In_2497);
and U3048 (N_3048,In_232,In_1257);
and U3049 (N_3049,In_603,In_2203);
xnor U3050 (N_3050,In_331,In_615);
nand U3051 (N_3051,In_2015,In_546);
nor U3052 (N_3052,In_1419,In_1363);
or U3053 (N_3053,In_1823,In_2035);
nor U3054 (N_3054,In_2514,In_2982);
nor U3055 (N_3055,In_577,In_2827);
and U3056 (N_3056,In_2608,In_753);
and U3057 (N_3057,In_2690,In_1115);
or U3058 (N_3058,In_46,In_2126);
nand U3059 (N_3059,In_1476,In_131);
nand U3060 (N_3060,In_1146,In_433);
nand U3061 (N_3061,In_651,In_2535);
nor U3062 (N_3062,In_2737,In_1871);
nand U3063 (N_3063,In_1274,In_2607);
or U3064 (N_3064,In_413,In_696);
and U3065 (N_3065,In_2734,In_2481);
xor U3066 (N_3066,In_2342,In_2239);
or U3067 (N_3067,In_2845,In_1341);
nor U3068 (N_3068,In_1451,In_894);
and U3069 (N_3069,In_2081,In_2945);
and U3070 (N_3070,In_1430,In_2600);
nand U3071 (N_3071,In_665,In_2205);
nor U3072 (N_3072,In_2732,In_2826);
nor U3073 (N_3073,In_166,In_1623);
nor U3074 (N_3074,In_2455,In_386);
nor U3075 (N_3075,In_1122,In_620);
and U3076 (N_3076,In_1142,In_2337);
nor U3077 (N_3077,In_1288,In_2553);
or U3078 (N_3078,In_368,In_1561);
nand U3079 (N_3079,In_718,In_2494);
and U3080 (N_3080,In_2067,In_1535);
nand U3081 (N_3081,In_2527,In_819);
or U3082 (N_3082,In_2497,In_2196);
or U3083 (N_3083,In_1508,In_1846);
nor U3084 (N_3084,In_1455,In_2398);
nand U3085 (N_3085,In_991,In_55);
or U3086 (N_3086,In_2487,In_2469);
nor U3087 (N_3087,In_625,In_2521);
or U3088 (N_3088,In_542,In_159);
xnor U3089 (N_3089,In_2305,In_1047);
nor U3090 (N_3090,In_2894,In_784);
nor U3091 (N_3091,In_1404,In_2070);
nor U3092 (N_3092,In_2755,In_2441);
or U3093 (N_3093,In_20,In_1569);
nor U3094 (N_3094,In_2882,In_2539);
and U3095 (N_3095,In_1526,In_1216);
nor U3096 (N_3096,In_1661,In_2348);
and U3097 (N_3097,In_1114,In_1846);
xnor U3098 (N_3098,In_775,In_874);
xor U3099 (N_3099,In_1026,In_2325);
and U3100 (N_3100,In_1710,In_482);
and U3101 (N_3101,In_2344,In_1763);
or U3102 (N_3102,In_1965,In_493);
nand U3103 (N_3103,In_1631,In_2692);
nor U3104 (N_3104,In_1312,In_2098);
xor U3105 (N_3105,In_2753,In_1462);
or U3106 (N_3106,In_2187,In_1983);
or U3107 (N_3107,In_718,In_1478);
nand U3108 (N_3108,In_475,In_1605);
nor U3109 (N_3109,In_1709,In_716);
or U3110 (N_3110,In_1791,In_2760);
xor U3111 (N_3111,In_2933,In_2370);
nand U3112 (N_3112,In_2793,In_1223);
nand U3113 (N_3113,In_133,In_1189);
nand U3114 (N_3114,In_1065,In_1646);
or U3115 (N_3115,In_1528,In_2700);
and U3116 (N_3116,In_27,In_1097);
nand U3117 (N_3117,In_2549,In_1055);
nor U3118 (N_3118,In_2900,In_710);
nor U3119 (N_3119,In_898,In_1625);
nor U3120 (N_3120,In_1009,In_1593);
and U3121 (N_3121,In_2814,In_502);
or U3122 (N_3122,In_570,In_2568);
nor U3123 (N_3123,In_292,In_2463);
nand U3124 (N_3124,In_46,In_860);
xor U3125 (N_3125,In_1233,In_501);
nand U3126 (N_3126,In_1317,In_1069);
nor U3127 (N_3127,In_2568,In_914);
nor U3128 (N_3128,In_2177,In_1870);
and U3129 (N_3129,In_827,In_2977);
and U3130 (N_3130,In_372,In_786);
nand U3131 (N_3131,In_354,In_2871);
or U3132 (N_3132,In_1497,In_1644);
or U3133 (N_3133,In_2137,In_891);
and U3134 (N_3134,In_840,In_2884);
or U3135 (N_3135,In_2780,In_1016);
nand U3136 (N_3136,In_809,In_19);
or U3137 (N_3137,In_1877,In_805);
or U3138 (N_3138,In_2935,In_1724);
and U3139 (N_3139,In_363,In_2308);
and U3140 (N_3140,In_1986,In_267);
nor U3141 (N_3141,In_2218,In_2533);
nor U3142 (N_3142,In_2561,In_1837);
or U3143 (N_3143,In_1211,In_920);
nand U3144 (N_3144,In_2629,In_2429);
and U3145 (N_3145,In_1454,In_191);
nor U3146 (N_3146,In_2166,In_2248);
or U3147 (N_3147,In_2824,In_1331);
nand U3148 (N_3148,In_685,In_403);
nor U3149 (N_3149,In_987,In_218);
nor U3150 (N_3150,In_1269,In_1567);
and U3151 (N_3151,In_2995,In_2217);
xor U3152 (N_3152,In_918,In_1110);
or U3153 (N_3153,In_2933,In_2653);
nand U3154 (N_3154,In_2865,In_1544);
nor U3155 (N_3155,In_1108,In_2548);
and U3156 (N_3156,In_1550,In_2203);
xor U3157 (N_3157,In_247,In_2248);
or U3158 (N_3158,In_2832,In_1768);
nor U3159 (N_3159,In_2052,In_1257);
and U3160 (N_3160,In_704,In_618);
and U3161 (N_3161,In_1263,In_124);
nor U3162 (N_3162,In_1171,In_2628);
or U3163 (N_3163,In_2111,In_604);
and U3164 (N_3164,In_495,In_1226);
nor U3165 (N_3165,In_2512,In_943);
or U3166 (N_3166,In_1883,In_542);
xor U3167 (N_3167,In_417,In_932);
nor U3168 (N_3168,In_826,In_1625);
nor U3169 (N_3169,In_736,In_777);
nand U3170 (N_3170,In_190,In_2580);
nor U3171 (N_3171,In_506,In_1226);
xnor U3172 (N_3172,In_1883,In_2968);
nor U3173 (N_3173,In_2258,In_2701);
or U3174 (N_3174,In_2206,In_725);
and U3175 (N_3175,In_2531,In_2790);
or U3176 (N_3176,In_323,In_2250);
and U3177 (N_3177,In_930,In_1176);
or U3178 (N_3178,In_2414,In_2785);
xor U3179 (N_3179,In_729,In_1227);
and U3180 (N_3180,In_1456,In_1306);
or U3181 (N_3181,In_303,In_1498);
or U3182 (N_3182,In_1894,In_2876);
and U3183 (N_3183,In_2938,In_132);
nor U3184 (N_3184,In_492,In_2320);
and U3185 (N_3185,In_2120,In_2002);
and U3186 (N_3186,In_2186,In_2218);
nand U3187 (N_3187,In_1638,In_396);
and U3188 (N_3188,In_299,In_1390);
nand U3189 (N_3189,In_2941,In_183);
or U3190 (N_3190,In_690,In_863);
and U3191 (N_3191,In_1150,In_2435);
nand U3192 (N_3192,In_2819,In_1525);
nand U3193 (N_3193,In_103,In_1033);
and U3194 (N_3194,In_1514,In_2002);
and U3195 (N_3195,In_2925,In_929);
nand U3196 (N_3196,In_640,In_1768);
xor U3197 (N_3197,In_1243,In_1749);
xor U3198 (N_3198,In_2531,In_1643);
and U3199 (N_3199,In_2994,In_902);
and U3200 (N_3200,In_1071,In_1879);
nor U3201 (N_3201,In_1298,In_1858);
nand U3202 (N_3202,In_1597,In_32);
nand U3203 (N_3203,In_2020,In_1369);
xor U3204 (N_3204,In_1835,In_2399);
and U3205 (N_3205,In_134,In_1971);
nor U3206 (N_3206,In_2700,In_2348);
nor U3207 (N_3207,In_1165,In_2453);
and U3208 (N_3208,In_541,In_1461);
and U3209 (N_3209,In_2384,In_888);
or U3210 (N_3210,In_1294,In_2848);
and U3211 (N_3211,In_1373,In_2791);
nor U3212 (N_3212,In_1319,In_2737);
nand U3213 (N_3213,In_1065,In_2070);
nor U3214 (N_3214,In_2861,In_1340);
and U3215 (N_3215,In_1390,In_1117);
nand U3216 (N_3216,In_2745,In_2350);
and U3217 (N_3217,In_1485,In_2409);
nor U3218 (N_3218,In_1073,In_2028);
nor U3219 (N_3219,In_847,In_525);
or U3220 (N_3220,In_1126,In_328);
nand U3221 (N_3221,In_1699,In_2850);
xor U3222 (N_3222,In_1868,In_1460);
or U3223 (N_3223,In_2983,In_1876);
or U3224 (N_3224,In_1591,In_590);
and U3225 (N_3225,In_446,In_533);
and U3226 (N_3226,In_1961,In_1275);
nand U3227 (N_3227,In_168,In_324);
xor U3228 (N_3228,In_1515,In_1083);
nor U3229 (N_3229,In_1330,In_1497);
and U3230 (N_3230,In_2482,In_1198);
nor U3231 (N_3231,In_2326,In_2327);
xor U3232 (N_3232,In_1068,In_220);
and U3233 (N_3233,In_729,In_1773);
or U3234 (N_3234,In_204,In_39);
or U3235 (N_3235,In_1374,In_2201);
nor U3236 (N_3236,In_2443,In_2256);
and U3237 (N_3237,In_209,In_2197);
xnor U3238 (N_3238,In_1766,In_421);
nor U3239 (N_3239,In_825,In_236);
nand U3240 (N_3240,In_2996,In_2093);
xnor U3241 (N_3241,In_2558,In_1882);
nor U3242 (N_3242,In_2918,In_2220);
and U3243 (N_3243,In_2342,In_1164);
or U3244 (N_3244,In_1876,In_1133);
or U3245 (N_3245,In_2731,In_1362);
nand U3246 (N_3246,In_1799,In_422);
nor U3247 (N_3247,In_2233,In_2454);
nand U3248 (N_3248,In_2446,In_2527);
and U3249 (N_3249,In_2119,In_1721);
or U3250 (N_3250,In_488,In_1999);
nand U3251 (N_3251,In_897,In_1687);
nand U3252 (N_3252,In_1409,In_2053);
and U3253 (N_3253,In_1007,In_2120);
and U3254 (N_3254,In_2283,In_449);
nand U3255 (N_3255,In_416,In_127);
nor U3256 (N_3256,In_1731,In_1703);
nor U3257 (N_3257,In_900,In_621);
and U3258 (N_3258,In_674,In_583);
nor U3259 (N_3259,In_1922,In_2767);
or U3260 (N_3260,In_1972,In_714);
and U3261 (N_3261,In_2639,In_146);
or U3262 (N_3262,In_1043,In_2230);
nor U3263 (N_3263,In_749,In_323);
nor U3264 (N_3264,In_554,In_1226);
and U3265 (N_3265,In_323,In_390);
nor U3266 (N_3266,In_421,In_2385);
nor U3267 (N_3267,In_1926,In_1658);
xnor U3268 (N_3268,In_2023,In_1299);
nand U3269 (N_3269,In_1221,In_566);
or U3270 (N_3270,In_2846,In_2276);
xnor U3271 (N_3271,In_2420,In_222);
nor U3272 (N_3272,In_2341,In_1410);
and U3273 (N_3273,In_264,In_1699);
nand U3274 (N_3274,In_1351,In_1177);
nand U3275 (N_3275,In_190,In_680);
nand U3276 (N_3276,In_2509,In_2442);
and U3277 (N_3277,In_2807,In_489);
nor U3278 (N_3278,In_584,In_2718);
and U3279 (N_3279,In_1377,In_2577);
nand U3280 (N_3280,In_1825,In_1970);
or U3281 (N_3281,In_2303,In_1717);
xor U3282 (N_3282,In_984,In_208);
nor U3283 (N_3283,In_2768,In_1096);
or U3284 (N_3284,In_11,In_1779);
and U3285 (N_3285,In_18,In_1188);
nand U3286 (N_3286,In_2729,In_1);
nand U3287 (N_3287,In_1790,In_2488);
nand U3288 (N_3288,In_1857,In_2919);
and U3289 (N_3289,In_848,In_567);
or U3290 (N_3290,In_2712,In_2341);
or U3291 (N_3291,In_225,In_1616);
and U3292 (N_3292,In_533,In_97);
nor U3293 (N_3293,In_1036,In_2228);
nor U3294 (N_3294,In_1265,In_1179);
nand U3295 (N_3295,In_2946,In_2510);
or U3296 (N_3296,In_1555,In_1101);
and U3297 (N_3297,In_1232,In_205);
xor U3298 (N_3298,In_1031,In_1908);
and U3299 (N_3299,In_1877,In_2799);
xnor U3300 (N_3300,In_418,In_1278);
nand U3301 (N_3301,In_1656,In_2180);
xor U3302 (N_3302,In_1346,In_2837);
nand U3303 (N_3303,In_2359,In_1159);
nor U3304 (N_3304,In_108,In_487);
or U3305 (N_3305,In_498,In_2491);
xnor U3306 (N_3306,In_1147,In_2321);
or U3307 (N_3307,In_1247,In_1169);
nor U3308 (N_3308,In_1729,In_2758);
and U3309 (N_3309,In_1183,In_354);
and U3310 (N_3310,In_2655,In_2048);
nor U3311 (N_3311,In_2396,In_1932);
and U3312 (N_3312,In_2153,In_2938);
or U3313 (N_3313,In_358,In_1326);
and U3314 (N_3314,In_1967,In_599);
or U3315 (N_3315,In_2664,In_37);
or U3316 (N_3316,In_1195,In_1643);
nand U3317 (N_3317,In_2611,In_886);
nor U3318 (N_3318,In_1851,In_2643);
nand U3319 (N_3319,In_2326,In_1312);
or U3320 (N_3320,In_608,In_2840);
nand U3321 (N_3321,In_1248,In_91);
or U3322 (N_3322,In_265,In_913);
nand U3323 (N_3323,In_2036,In_1576);
and U3324 (N_3324,In_2690,In_322);
xnor U3325 (N_3325,In_1800,In_1657);
or U3326 (N_3326,In_2882,In_2286);
nand U3327 (N_3327,In_742,In_355);
nor U3328 (N_3328,In_1295,In_342);
or U3329 (N_3329,In_2754,In_2359);
and U3330 (N_3330,In_439,In_2699);
xnor U3331 (N_3331,In_1541,In_383);
or U3332 (N_3332,In_941,In_767);
and U3333 (N_3333,In_2810,In_2777);
nor U3334 (N_3334,In_1691,In_2989);
nor U3335 (N_3335,In_343,In_2410);
xor U3336 (N_3336,In_396,In_1170);
or U3337 (N_3337,In_944,In_2656);
and U3338 (N_3338,In_2817,In_1416);
and U3339 (N_3339,In_878,In_986);
nand U3340 (N_3340,In_2639,In_2245);
and U3341 (N_3341,In_2944,In_1787);
and U3342 (N_3342,In_1279,In_985);
nor U3343 (N_3343,In_1048,In_2598);
xor U3344 (N_3344,In_1876,In_2342);
and U3345 (N_3345,In_2502,In_2263);
and U3346 (N_3346,In_233,In_1040);
and U3347 (N_3347,In_2253,In_2401);
or U3348 (N_3348,In_812,In_2654);
or U3349 (N_3349,In_2373,In_436);
xnor U3350 (N_3350,In_1466,In_1800);
nor U3351 (N_3351,In_1186,In_321);
xor U3352 (N_3352,In_956,In_300);
xnor U3353 (N_3353,In_1085,In_942);
nor U3354 (N_3354,In_1476,In_2910);
or U3355 (N_3355,In_353,In_1442);
xnor U3356 (N_3356,In_1313,In_1765);
or U3357 (N_3357,In_85,In_1567);
or U3358 (N_3358,In_2167,In_1256);
or U3359 (N_3359,In_1475,In_2520);
or U3360 (N_3360,In_1589,In_699);
and U3361 (N_3361,In_2395,In_1014);
or U3362 (N_3362,In_115,In_1828);
nand U3363 (N_3363,In_2704,In_1234);
and U3364 (N_3364,In_2092,In_2938);
xnor U3365 (N_3365,In_2948,In_2465);
nor U3366 (N_3366,In_1847,In_794);
nand U3367 (N_3367,In_1212,In_1348);
nor U3368 (N_3368,In_2168,In_384);
xnor U3369 (N_3369,In_1487,In_1355);
nand U3370 (N_3370,In_2568,In_1283);
nand U3371 (N_3371,In_2603,In_1874);
or U3372 (N_3372,In_2377,In_2835);
nand U3373 (N_3373,In_142,In_143);
nand U3374 (N_3374,In_229,In_1493);
and U3375 (N_3375,In_894,In_143);
nand U3376 (N_3376,In_2847,In_2678);
and U3377 (N_3377,In_1052,In_810);
and U3378 (N_3378,In_17,In_276);
nand U3379 (N_3379,In_2919,In_602);
nand U3380 (N_3380,In_2469,In_1538);
or U3381 (N_3381,In_1735,In_1462);
or U3382 (N_3382,In_1198,In_1298);
and U3383 (N_3383,In_2815,In_1691);
or U3384 (N_3384,In_879,In_372);
or U3385 (N_3385,In_2148,In_2172);
and U3386 (N_3386,In_1941,In_414);
or U3387 (N_3387,In_1981,In_2265);
or U3388 (N_3388,In_735,In_2703);
xnor U3389 (N_3389,In_2946,In_2068);
nor U3390 (N_3390,In_2262,In_404);
nand U3391 (N_3391,In_1967,In_2947);
xor U3392 (N_3392,In_134,In_1004);
and U3393 (N_3393,In_634,In_1128);
and U3394 (N_3394,In_1414,In_887);
and U3395 (N_3395,In_125,In_337);
or U3396 (N_3396,In_1845,In_1615);
nand U3397 (N_3397,In_1285,In_362);
nor U3398 (N_3398,In_1751,In_1042);
xor U3399 (N_3399,In_233,In_2169);
nor U3400 (N_3400,In_1643,In_349);
nor U3401 (N_3401,In_1432,In_1364);
nand U3402 (N_3402,In_1870,In_2634);
xor U3403 (N_3403,In_42,In_1808);
nor U3404 (N_3404,In_755,In_963);
or U3405 (N_3405,In_237,In_109);
nor U3406 (N_3406,In_2820,In_2208);
or U3407 (N_3407,In_701,In_2037);
or U3408 (N_3408,In_137,In_2500);
nand U3409 (N_3409,In_1408,In_1765);
xnor U3410 (N_3410,In_1333,In_1931);
nor U3411 (N_3411,In_755,In_2164);
and U3412 (N_3412,In_2203,In_2456);
nand U3413 (N_3413,In_2823,In_418);
nor U3414 (N_3414,In_1224,In_2611);
or U3415 (N_3415,In_2197,In_1353);
nand U3416 (N_3416,In_874,In_2389);
nand U3417 (N_3417,In_110,In_2535);
xnor U3418 (N_3418,In_2241,In_828);
and U3419 (N_3419,In_1948,In_1038);
nand U3420 (N_3420,In_2612,In_657);
and U3421 (N_3421,In_281,In_2202);
and U3422 (N_3422,In_1116,In_256);
nor U3423 (N_3423,In_148,In_1320);
and U3424 (N_3424,In_2253,In_2841);
nor U3425 (N_3425,In_800,In_586);
or U3426 (N_3426,In_1055,In_534);
nand U3427 (N_3427,In_2857,In_515);
and U3428 (N_3428,In_2299,In_843);
nand U3429 (N_3429,In_2890,In_1807);
or U3430 (N_3430,In_776,In_184);
xnor U3431 (N_3431,In_542,In_1245);
or U3432 (N_3432,In_165,In_2209);
nor U3433 (N_3433,In_1255,In_863);
nor U3434 (N_3434,In_2321,In_840);
nand U3435 (N_3435,In_2155,In_1965);
nand U3436 (N_3436,In_2729,In_493);
nand U3437 (N_3437,In_1580,In_2880);
nand U3438 (N_3438,In_1072,In_518);
nand U3439 (N_3439,In_337,In_2490);
nor U3440 (N_3440,In_104,In_378);
or U3441 (N_3441,In_2167,In_1185);
and U3442 (N_3442,In_490,In_388);
or U3443 (N_3443,In_1363,In_2519);
or U3444 (N_3444,In_473,In_873);
nand U3445 (N_3445,In_664,In_725);
and U3446 (N_3446,In_21,In_2196);
or U3447 (N_3447,In_801,In_1644);
and U3448 (N_3448,In_1058,In_1045);
and U3449 (N_3449,In_110,In_1927);
nand U3450 (N_3450,In_1056,In_1158);
nand U3451 (N_3451,In_1246,In_2288);
nor U3452 (N_3452,In_58,In_1439);
nand U3453 (N_3453,In_807,In_1460);
xor U3454 (N_3454,In_995,In_699);
nor U3455 (N_3455,In_1501,In_2887);
xnor U3456 (N_3456,In_2500,In_1795);
xor U3457 (N_3457,In_749,In_1753);
or U3458 (N_3458,In_2855,In_2482);
and U3459 (N_3459,In_2505,In_2414);
nand U3460 (N_3460,In_2971,In_258);
nor U3461 (N_3461,In_1806,In_1274);
or U3462 (N_3462,In_2974,In_2559);
nand U3463 (N_3463,In_2795,In_1898);
or U3464 (N_3464,In_1770,In_1196);
nor U3465 (N_3465,In_2357,In_1799);
nand U3466 (N_3466,In_1681,In_2011);
nor U3467 (N_3467,In_1920,In_671);
or U3468 (N_3468,In_2805,In_2277);
or U3469 (N_3469,In_1688,In_1938);
nand U3470 (N_3470,In_909,In_213);
nand U3471 (N_3471,In_1131,In_1907);
or U3472 (N_3472,In_2967,In_2946);
nand U3473 (N_3473,In_634,In_2111);
and U3474 (N_3474,In_954,In_1290);
xnor U3475 (N_3475,In_2831,In_409);
or U3476 (N_3476,In_553,In_2367);
nand U3477 (N_3477,In_2849,In_940);
nand U3478 (N_3478,In_296,In_187);
and U3479 (N_3479,In_1187,In_1617);
nand U3480 (N_3480,In_2849,In_587);
nor U3481 (N_3481,In_1769,In_593);
and U3482 (N_3482,In_2153,In_2382);
and U3483 (N_3483,In_241,In_61);
and U3484 (N_3484,In_1591,In_1682);
nand U3485 (N_3485,In_2422,In_2350);
nand U3486 (N_3486,In_1826,In_1455);
nor U3487 (N_3487,In_725,In_2737);
and U3488 (N_3488,In_2094,In_1330);
or U3489 (N_3489,In_1118,In_2160);
or U3490 (N_3490,In_2648,In_1262);
and U3491 (N_3491,In_399,In_1068);
or U3492 (N_3492,In_1791,In_2436);
xor U3493 (N_3493,In_1047,In_1125);
nand U3494 (N_3494,In_1470,In_147);
and U3495 (N_3495,In_2954,In_1789);
and U3496 (N_3496,In_1632,In_613);
nor U3497 (N_3497,In_915,In_1817);
nand U3498 (N_3498,In_2168,In_1779);
nor U3499 (N_3499,In_1274,In_1118);
or U3500 (N_3500,In_844,In_817);
or U3501 (N_3501,In_2731,In_689);
xor U3502 (N_3502,In_2925,In_1271);
and U3503 (N_3503,In_2281,In_1063);
and U3504 (N_3504,In_2085,In_2083);
nand U3505 (N_3505,In_2318,In_900);
and U3506 (N_3506,In_1174,In_656);
and U3507 (N_3507,In_653,In_1660);
and U3508 (N_3508,In_2777,In_2318);
or U3509 (N_3509,In_858,In_312);
and U3510 (N_3510,In_1460,In_1936);
and U3511 (N_3511,In_1424,In_997);
or U3512 (N_3512,In_57,In_1851);
nand U3513 (N_3513,In_395,In_405);
nor U3514 (N_3514,In_1770,In_1943);
nor U3515 (N_3515,In_2351,In_2095);
and U3516 (N_3516,In_2239,In_339);
and U3517 (N_3517,In_1357,In_2845);
and U3518 (N_3518,In_2864,In_1884);
and U3519 (N_3519,In_1857,In_2731);
nand U3520 (N_3520,In_468,In_1580);
or U3521 (N_3521,In_1599,In_91);
nand U3522 (N_3522,In_1282,In_275);
nand U3523 (N_3523,In_1495,In_1562);
or U3524 (N_3524,In_360,In_653);
nor U3525 (N_3525,In_911,In_2775);
nand U3526 (N_3526,In_603,In_2843);
nor U3527 (N_3527,In_2085,In_1358);
and U3528 (N_3528,In_854,In_1033);
and U3529 (N_3529,In_2569,In_149);
nand U3530 (N_3530,In_293,In_2447);
nand U3531 (N_3531,In_2033,In_692);
and U3532 (N_3532,In_907,In_380);
nor U3533 (N_3533,In_2856,In_2064);
or U3534 (N_3534,In_1790,In_2970);
or U3535 (N_3535,In_2996,In_2023);
or U3536 (N_3536,In_1272,In_1067);
or U3537 (N_3537,In_2407,In_114);
and U3538 (N_3538,In_2186,In_1133);
nand U3539 (N_3539,In_2878,In_869);
nand U3540 (N_3540,In_1816,In_1365);
and U3541 (N_3541,In_252,In_2620);
and U3542 (N_3542,In_515,In_1799);
and U3543 (N_3543,In_630,In_819);
and U3544 (N_3544,In_110,In_285);
or U3545 (N_3545,In_2355,In_2694);
nor U3546 (N_3546,In_1837,In_1342);
nand U3547 (N_3547,In_1689,In_1900);
and U3548 (N_3548,In_1508,In_2732);
nor U3549 (N_3549,In_1494,In_305);
nand U3550 (N_3550,In_398,In_2247);
and U3551 (N_3551,In_394,In_2951);
nand U3552 (N_3552,In_934,In_884);
and U3553 (N_3553,In_2717,In_612);
or U3554 (N_3554,In_2376,In_1986);
and U3555 (N_3555,In_984,In_607);
and U3556 (N_3556,In_216,In_549);
nand U3557 (N_3557,In_949,In_1334);
nor U3558 (N_3558,In_113,In_1083);
nor U3559 (N_3559,In_929,In_2817);
nand U3560 (N_3560,In_1174,In_2958);
or U3561 (N_3561,In_1556,In_2568);
and U3562 (N_3562,In_1510,In_2400);
and U3563 (N_3563,In_351,In_2400);
and U3564 (N_3564,In_2865,In_2878);
or U3565 (N_3565,In_969,In_1660);
xor U3566 (N_3566,In_1050,In_1412);
and U3567 (N_3567,In_335,In_1544);
nor U3568 (N_3568,In_2128,In_2850);
or U3569 (N_3569,In_982,In_1696);
nor U3570 (N_3570,In_343,In_2244);
nand U3571 (N_3571,In_447,In_1836);
or U3572 (N_3572,In_1860,In_2859);
nor U3573 (N_3573,In_2317,In_2102);
nand U3574 (N_3574,In_1901,In_2739);
nor U3575 (N_3575,In_2402,In_203);
nand U3576 (N_3576,In_1697,In_2645);
nor U3577 (N_3577,In_2308,In_344);
or U3578 (N_3578,In_2432,In_704);
and U3579 (N_3579,In_2703,In_1400);
nand U3580 (N_3580,In_2829,In_1327);
or U3581 (N_3581,In_643,In_2612);
nand U3582 (N_3582,In_652,In_1684);
or U3583 (N_3583,In_379,In_1);
nand U3584 (N_3584,In_2884,In_1483);
nand U3585 (N_3585,In_1842,In_272);
nand U3586 (N_3586,In_14,In_2145);
nand U3587 (N_3587,In_2597,In_1925);
or U3588 (N_3588,In_2229,In_361);
nor U3589 (N_3589,In_102,In_2977);
nor U3590 (N_3590,In_1909,In_1747);
nor U3591 (N_3591,In_320,In_2142);
or U3592 (N_3592,In_431,In_1622);
nand U3593 (N_3593,In_2829,In_1274);
nor U3594 (N_3594,In_1060,In_1613);
xor U3595 (N_3595,In_1062,In_1341);
or U3596 (N_3596,In_310,In_2412);
or U3597 (N_3597,In_1312,In_691);
nor U3598 (N_3598,In_1146,In_458);
and U3599 (N_3599,In_2394,In_2158);
or U3600 (N_3600,In_591,In_2109);
and U3601 (N_3601,In_1517,In_2403);
or U3602 (N_3602,In_1352,In_41);
nand U3603 (N_3603,In_2761,In_2566);
nor U3604 (N_3604,In_1696,In_1772);
or U3605 (N_3605,In_2452,In_733);
nand U3606 (N_3606,In_573,In_2525);
and U3607 (N_3607,In_1328,In_2359);
and U3608 (N_3608,In_2442,In_1977);
or U3609 (N_3609,In_100,In_1793);
and U3610 (N_3610,In_2273,In_1479);
nand U3611 (N_3611,In_705,In_1140);
nand U3612 (N_3612,In_367,In_2511);
nor U3613 (N_3613,In_1253,In_783);
and U3614 (N_3614,In_2238,In_931);
nand U3615 (N_3615,In_2591,In_2181);
nand U3616 (N_3616,In_1721,In_1262);
nand U3617 (N_3617,In_1484,In_1407);
xnor U3618 (N_3618,In_229,In_2069);
nor U3619 (N_3619,In_1308,In_1418);
xnor U3620 (N_3620,In_2625,In_2880);
and U3621 (N_3621,In_2706,In_593);
and U3622 (N_3622,In_2595,In_2016);
and U3623 (N_3623,In_615,In_430);
and U3624 (N_3624,In_1582,In_1921);
xor U3625 (N_3625,In_540,In_1620);
and U3626 (N_3626,In_869,In_2846);
or U3627 (N_3627,In_2745,In_136);
nor U3628 (N_3628,In_1922,In_502);
or U3629 (N_3629,In_1871,In_654);
and U3630 (N_3630,In_779,In_221);
nand U3631 (N_3631,In_1378,In_1745);
and U3632 (N_3632,In_1490,In_1892);
and U3633 (N_3633,In_1412,In_2270);
nor U3634 (N_3634,In_1872,In_2566);
nand U3635 (N_3635,In_2969,In_2912);
nor U3636 (N_3636,In_508,In_855);
nand U3637 (N_3637,In_976,In_2723);
or U3638 (N_3638,In_751,In_2531);
nor U3639 (N_3639,In_2821,In_1965);
nor U3640 (N_3640,In_2482,In_1457);
nand U3641 (N_3641,In_2889,In_1692);
or U3642 (N_3642,In_2425,In_2272);
and U3643 (N_3643,In_2050,In_1188);
or U3644 (N_3644,In_491,In_384);
nor U3645 (N_3645,In_1185,In_625);
nand U3646 (N_3646,In_45,In_523);
and U3647 (N_3647,In_2244,In_457);
and U3648 (N_3648,In_1426,In_2208);
nor U3649 (N_3649,In_1578,In_2066);
nand U3650 (N_3650,In_2256,In_452);
or U3651 (N_3651,In_2274,In_1296);
or U3652 (N_3652,In_1335,In_1482);
or U3653 (N_3653,In_417,In_769);
and U3654 (N_3654,In_2747,In_771);
or U3655 (N_3655,In_1075,In_1040);
nor U3656 (N_3656,In_1680,In_2457);
and U3657 (N_3657,In_2916,In_2040);
nand U3658 (N_3658,In_2973,In_848);
nand U3659 (N_3659,In_445,In_755);
xor U3660 (N_3660,In_1944,In_1686);
and U3661 (N_3661,In_1515,In_2781);
nand U3662 (N_3662,In_1728,In_1609);
and U3663 (N_3663,In_1561,In_1300);
or U3664 (N_3664,In_2594,In_1746);
nor U3665 (N_3665,In_321,In_2052);
xnor U3666 (N_3666,In_2462,In_653);
nor U3667 (N_3667,In_2094,In_1448);
nor U3668 (N_3668,In_715,In_2339);
nor U3669 (N_3669,In_2780,In_2871);
or U3670 (N_3670,In_2129,In_2380);
nor U3671 (N_3671,In_2895,In_2642);
or U3672 (N_3672,In_296,In_1073);
nor U3673 (N_3673,In_2321,In_1156);
nor U3674 (N_3674,In_2791,In_712);
and U3675 (N_3675,In_2986,In_560);
nor U3676 (N_3676,In_2181,In_1425);
xor U3677 (N_3677,In_313,In_117);
and U3678 (N_3678,In_2702,In_804);
xnor U3679 (N_3679,In_1917,In_311);
nor U3680 (N_3680,In_2250,In_646);
or U3681 (N_3681,In_549,In_1700);
nor U3682 (N_3682,In_410,In_737);
and U3683 (N_3683,In_780,In_2567);
xnor U3684 (N_3684,In_2356,In_1769);
xor U3685 (N_3685,In_2301,In_128);
and U3686 (N_3686,In_2021,In_2209);
nor U3687 (N_3687,In_657,In_2638);
nor U3688 (N_3688,In_466,In_1775);
or U3689 (N_3689,In_2067,In_197);
and U3690 (N_3690,In_742,In_32);
nor U3691 (N_3691,In_220,In_208);
nor U3692 (N_3692,In_2999,In_1136);
nand U3693 (N_3693,In_2747,In_2839);
and U3694 (N_3694,In_428,In_1013);
nor U3695 (N_3695,In_1420,In_1622);
or U3696 (N_3696,In_1666,In_2303);
xnor U3697 (N_3697,In_2942,In_296);
nand U3698 (N_3698,In_1023,In_286);
xnor U3699 (N_3699,In_151,In_1816);
nor U3700 (N_3700,In_1083,In_1348);
or U3701 (N_3701,In_2229,In_2894);
and U3702 (N_3702,In_1261,In_1858);
or U3703 (N_3703,In_950,In_1225);
or U3704 (N_3704,In_207,In_1725);
and U3705 (N_3705,In_47,In_2330);
nor U3706 (N_3706,In_2436,In_2995);
and U3707 (N_3707,In_1937,In_348);
and U3708 (N_3708,In_400,In_2089);
nor U3709 (N_3709,In_2420,In_37);
nor U3710 (N_3710,In_2100,In_320);
and U3711 (N_3711,In_1737,In_236);
nor U3712 (N_3712,In_2984,In_1018);
xor U3713 (N_3713,In_2175,In_1442);
and U3714 (N_3714,In_1284,In_866);
xor U3715 (N_3715,In_1166,In_2761);
or U3716 (N_3716,In_2249,In_1093);
or U3717 (N_3717,In_1372,In_1416);
nor U3718 (N_3718,In_79,In_2471);
and U3719 (N_3719,In_2353,In_913);
nor U3720 (N_3720,In_2875,In_125);
nor U3721 (N_3721,In_2832,In_732);
and U3722 (N_3722,In_1165,In_2810);
nor U3723 (N_3723,In_2884,In_2269);
or U3724 (N_3724,In_1662,In_826);
nor U3725 (N_3725,In_1403,In_198);
nor U3726 (N_3726,In_1690,In_489);
or U3727 (N_3727,In_1022,In_145);
or U3728 (N_3728,In_2163,In_471);
nor U3729 (N_3729,In_1069,In_1187);
or U3730 (N_3730,In_3,In_209);
nand U3731 (N_3731,In_2227,In_2523);
nor U3732 (N_3732,In_1390,In_320);
nand U3733 (N_3733,In_1547,In_650);
and U3734 (N_3734,In_1940,In_2153);
and U3735 (N_3735,In_2981,In_1642);
nor U3736 (N_3736,In_765,In_1906);
nor U3737 (N_3737,In_1967,In_886);
or U3738 (N_3738,In_2076,In_74);
nor U3739 (N_3739,In_2577,In_2539);
and U3740 (N_3740,In_1327,In_2738);
nand U3741 (N_3741,In_1755,In_2571);
and U3742 (N_3742,In_1873,In_1110);
or U3743 (N_3743,In_864,In_1583);
nor U3744 (N_3744,In_2661,In_889);
xor U3745 (N_3745,In_1782,In_1351);
and U3746 (N_3746,In_195,In_2903);
or U3747 (N_3747,In_881,In_878);
nor U3748 (N_3748,In_2200,In_154);
nor U3749 (N_3749,In_406,In_1455);
or U3750 (N_3750,In_253,In_1419);
or U3751 (N_3751,In_1232,In_2150);
or U3752 (N_3752,In_2512,In_1745);
nor U3753 (N_3753,In_1426,In_2290);
and U3754 (N_3754,In_547,In_1894);
and U3755 (N_3755,In_2031,In_1412);
nand U3756 (N_3756,In_2481,In_430);
xor U3757 (N_3757,In_917,In_2031);
nor U3758 (N_3758,In_2744,In_55);
or U3759 (N_3759,In_1760,In_37);
nor U3760 (N_3760,In_2078,In_1859);
or U3761 (N_3761,In_470,In_2095);
nor U3762 (N_3762,In_1253,In_1918);
nor U3763 (N_3763,In_1878,In_1434);
or U3764 (N_3764,In_2377,In_1877);
nor U3765 (N_3765,In_2109,In_43);
and U3766 (N_3766,In_741,In_1751);
and U3767 (N_3767,In_54,In_2792);
and U3768 (N_3768,In_1800,In_2130);
nor U3769 (N_3769,In_555,In_867);
nand U3770 (N_3770,In_1162,In_1767);
xnor U3771 (N_3771,In_2095,In_1902);
nand U3772 (N_3772,In_1585,In_2585);
xor U3773 (N_3773,In_1150,In_2929);
or U3774 (N_3774,In_429,In_2751);
nor U3775 (N_3775,In_944,In_1378);
or U3776 (N_3776,In_1293,In_1634);
nor U3777 (N_3777,In_1908,In_646);
or U3778 (N_3778,In_2058,In_412);
nor U3779 (N_3779,In_1240,In_2763);
nand U3780 (N_3780,In_1530,In_2552);
or U3781 (N_3781,In_1229,In_1819);
nand U3782 (N_3782,In_858,In_1432);
nor U3783 (N_3783,In_1099,In_2939);
or U3784 (N_3784,In_1545,In_44);
nand U3785 (N_3785,In_594,In_2636);
nor U3786 (N_3786,In_1081,In_1426);
and U3787 (N_3787,In_1337,In_787);
nor U3788 (N_3788,In_2580,In_2209);
xnor U3789 (N_3789,In_2646,In_1109);
or U3790 (N_3790,In_238,In_2080);
or U3791 (N_3791,In_1224,In_2827);
and U3792 (N_3792,In_1812,In_955);
nand U3793 (N_3793,In_1325,In_2958);
nand U3794 (N_3794,In_1394,In_244);
xor U3795 (N_3795,In_1105,In_2907);
nor U3796 (N_3796,In_78,In_1474);
nor U3797 (N_3797,In_1709,In_1071);
nand U3798 (N_3798,In_2458,In_2306);
nor U3799 (N_3799,In_2045,In_304);
or U3800 (N_3800,In_1281,In_2810);
and U3801 (N_3801,In_651,In_2197);
nor U3802 (N_3802,In_776,In_326);
and U3803 (N_3803,In_1260,In_613);
nor U3804 (N_3804,In_2491,In_1880);
nand U3805 (N_3805,In_966,In_568);
nor U3806 (N_3806,In_712,In_2035);
or U3807 (N_3807,In_1476,In_304);
xnor U3808 (N_3808,In_1464,In_794);
nor U3809 (N_3809,In_2867,In_753);
nand U3810 (N_3810,In_1822,In_1768);
and U3811 (N_3811,In_2248,In_155);
nand U3812 (N_3812,In_2527,In_2925);
nand U3813 (N_3813,In_501,In_2773);
nand U3814 (N_3814,In_1649,In_991);
and U3815 (N_3815,In_2785,In_1436);
or U3816 (N_3816,In_2362,In_2313);
nor U3817 (N_3817,In_1733,In_952);
and U3818 (N_3818,In_655,In_71);
nand U3819 (N_3819,In_2221,In_1396);
or U3820 (N_3820,In_1578,In_522);
or U3821 (N_3821,In_1090,In_1883);
and U3822 (N_3822,In_2447,In_2441);
nand U3823 (N_3823,In_1004,In_2584);
or U3824 (N_3824,In_742,In_2120);
or U3825 (N_3825,In_1508,In_214);
nand U3826 (N_3826,In_2368,In_856);
or U3827 (N_3827,In_1859,In_2047);
nor U3828 (N_3828,In_1338,In_2523);
nand U3829 (N_3829,In_697,In_657);
nand U3830 (N_3830,In_1115,In_2784);
and U3831 (N_3831,In_764,In_1047);
or U3832 (N_3832,In_129,In_1174);
nor U3833 (N_3833,In_2812,In_1301);
nor U3834 (N_3834,In_2487,In_960);
and U3835 (N_3835,In_2660,In_2275);
nand U3836 (N_3836,In_651,In_1610);
and U3837 (N_3837,In_2517,In_1392);
or U3838 (N_3838,In_335,In_530);
xor U3839 (N_3839,In_61,In_2169);
nand U3840 (N_3840,In_1708,In_333);
xnor U3841 (N_3841,In_1026,In_2401);
and U3842 (N_3842,In_946,In_1683);
nand U3843 (N_3843,In_2057,In_1644);
or U3844 (N_3844,In_2687,In_1385);
and U3845 (N_3845,In_2037,In_1894);
and U3846 (N_3846,In_1534,In_2706);
and U3847 (N_3847,In_219,In_1596);
nand U3848 (N_3848,In_524,In_1083);
or U3849 (N_3849,In_1813,In_1158);
nand U3850 (N_3850,In_2697,In_1222);
nor U3851 (N_3851,In_154,In_274);
nor U3852 (N_3852,In_1761,In_1984);
or U3853 (N_3853,In_2946,In_420);
nor U3854 (N_3854,In_978,In_1844);
nand U3855 (N_3855,In_860,In_2676);
and U3856 (N_3856,In_857,In_1456);
xor U3857 (N_3857,In_949,In_2855);
and U3858 (N_3858,In_1737,In_1483);
and U3859 (N_3859,In_1258,In_355);
or U3860 (N_3860,In_2725,In_2247);
nand U3861 (N_3861,In_1856,In_2785);
or U3862 (N_3862,In_967,In_1170);
nand U3863 (N_3863,In_1928,In_18);
nand U3864 (N_3864,In_546,In_1277);
and U3865 (N_3865,In_2278,In_301);
and U3866 (N_3866,In_1564,In_2410);
and U3867 (N_3867,In_2149,In_1876);
nor U3868 (N_3868,In_1833,In_2495);
nor U3869 (N_3869,In_1732,In_959);
nor U3870 (N_3870,In_1173,In_1942);
nand U3871 (N_3871,In_1735,In_245);
nand U3872 (N_3872,In_728,In_2649);
and U3873 (N_3873,In_2289,In_2319);
nand U3874 (N_3874,In_2808,In_1484);
nand U3875 (N_3875,In_1461,In_1676);
or U3876 (N_3876,In_909,In_1158);
nand U3877 (N_3877,In_2874,In_1030);
nand U3878 (N_3878,In_132,In_1213);
nand U3879 (N_3879,In_1019,In_1985);
nand U3880 (N_3880,In_9,In_1289);
or U3881 (N_3881,In_2304,In_236);
and U3882 (N_3882,In_2622,In_2707);
or U3883 (N_3883,In_838,In_2402);
and U3884 (N_3884,In_940,In_850);
nand U3885 (N_3885,In_1788,In_2821);
xor U3886 (N_3886,In_78,In_2588);
nand U3887 (N_3887,In_712,In_1337);
nor U3888 (N_3888,In_2617,In_1561);
or U3889 (N_3889,In_2501,In_2841);
nand U3890 (N_3890,In_1215,In_53);
or U3891 (N_3891,In_1173,In_739);
nor U3892 (N_3892,In_1506,In_1636);
nand U3893 (N_3893,In_233,In_2342);
and U3894 (N_3894,In_2571,In_233);
or U3895 (N_3895,In_2906,In_211);
xor U3896 (N_3896,In_1498,In_204);
or U3897 (N_3897,In_650,In_1455);
or U3898 (N_3898,In_1623,In_675);
and U3899 (N_3899,In_924,In_1725);
and U3900 (N_3900,In_2917,In_60);
or U3901 (N_3901,In_234,In_537);
nor U3902 (N_3902,In_1375,In_338);
nand U3903 (N_3903,In_1516,In_2278);
or U3904 (N_3904,In_2119,In_1515);
and U3905 (N_3905,In_2015,In_566);
and U3906 (N_3906,In_2164,In_1272);
or U3907 (N_3907,In_2319,In_2539);
or U3908 (N_3908,In_2819,In_705);
and U3909 (N_3909,In_2930,In_1947);
nor U3910 (N_3910,In_720,In_1235);
xor U3911 (N_3911,In_1750,In_1141);
or U3912 (N_3912,In_1083,In_501);
nor U3913 (N_3913,In_705,In_2895);
and U3914 (N_3914,In_1635,In_1529);
nand U3915 (N_3915,In_1483,In_1697);
nand U3916 (N_3916,In_469,In_408);
and U3917 (N_3917,In_2881,In_663);
and U3918 (N_3918,In_701,In_2888);
xor U3919 (N_3919,In_2149,In_2291);
or U3920 (N_3920,In_1126,In_1698);
and U3921 (N_3921,In_1253,In_2838);
nor U3922 (N_3922,In_2433,In_1284);
and U3923 (N_3923,In_2826,In_600);
or U3924 (N_3924,In_386,In_2038);
nand U3925 (N_3925,In_1505,In_262);
xor U3926 (N_3926,In_2092,In_1480);
nand U3927 (N_3927,In_1070,In_1518);
or U3928 (N_3928,In_2503,In_2395);
or U3929 (N_3929,In_1508,In_2286);
or U3930 (N_3930,In_629,In_2430);
and U3931 (N_3931,In_219,In_715);
nor U3932 (N_3932,In_990,In_2460);
and U3933 (N_3933,In_1800,In_482);
or U3934 (N_3934,In_2372,In_677);
nand U3935 (N_3935,In_1933,In_1226);
and U3936 (N_3936,In_10,In_2107);
nor U3937 (N_3937,In_1575,In_1252);
or U3938 (N_3938,In_2021,In_1688);
nand U3939 (N_3939,In_1957,In_273);
and U3940 (N_3940,In_298,In_310);
or U3941 (N_3941,In_92,In_1568);
or U3942 (N_3942,In_1078,In_2724);
or U3943 (N_3943,In_1126,In_1268);
or U3944 (N_3944,In_2098,In_2858);
or U3945 (N_3945,In_1115,In_2646);
or U3946 (N_3946,In_2668,In_402);
or U3947 (N_3947,In_2175,In_2658);
and U3948 (N_3948,In_2365,In_2589);
and U3949 (N_3949,In_447,In_2900);
nor U3950 (N_3950,In_2451,In_2547);
nand U3951 (N_3951,In_2420,In_55);
or U3952 (N_3952,In_2165,In_2543);
nor U3953 (N_3953,In_1481,In_1415);
xnor U3954 (N_3954,In_2154,In_1088);
and U3955 (N_3955,In_908,In_1249);
nor U3956 (N_3956,In_1736,In_159);
and U3957 (N_3957,In_1313,In_1847);
nor U3958 (N_3958,In_385,In_117);
nand U3959 (N_3959,In_2065,In_1513);
nor U3960 (N_3960,In_1500,In_1264);
nor U3961 (N_3961,In_1850,In_1194);
and U3962 (N_3962,In_1572,In_395);
and U3963 (N_3963,In_2395,In_1816);
nor U3964 (N_3964,In_2235,In_2757);
nor U3965 (N_3965,In_2244,In_1525);
nand U3966 (N_3966,In_2203,In_2777);
xor U3967 (N_3967,In_2955,In_2561);
and U3968 (N_3968,In_2028,In_1767);
nand U3969 (N_3969,In_304,In_2640);
and U3970 (N_3970,In_525,In_2677);
xor U3971 (N_3971,In_2586,In_223);
nand U3972 (N_3972,In_2907,In_677);
nor U3973 (N_3973,In_2305,In_1001);
nor U3974 (N_3974,In_1864,In_2366);
and U3975 (N_3975,In_887,In_1837);
nor U3976 (N_3976,In_502,In_617);
nor U3977 (N_3977,In_2141,In_2610);
xor U3978 (N_3978,In_2771,In_211);
or U3979 (N_3979,In_2371,In_355);
and U3980 (N_3980,In_1202,In_1095);
nand U3981 (N_3981,In_1830,In_2644);
nor U3982 (N_3982,In_1239,In_255);
nand U3983 (N_3983,In_799,In_784);
and U3984 (N_3984,In_2823,In_58);
and U3985 (N_3985,In_1097,In_1918);
nor U3986 (N_3986,In_1842,In_2444);
or U3987 (N_3987,In_2379,In_438);
xnor U3988 (N_3988,In_2586,In_1638);
and U3989 (N_3989,In_696,In_566);
nand U3990 (N_3990,In_1522,In_6);
xnor U3991 (N_3991,In_2234,In_1402);
or U3992 (N_3992,In_468,In_794);
nand U3993 (N_3993,In_1008,In_883);
and U3994 (N_3994,In_1141,In_133);
or U3995 (N_3995,In_2865,In_2706);
or U3996 (N_3996,In_2160,In_523);
nor U3997 (N_3997,In_1275,In_2722);
or U3998 (N_3998,In_2811,In_604);
and U3999 (N_3999,In_1880,In_613);
nand U4000 (N_4000,In_252,In_2510);
nor U4001 (N_4001,In_1314,In_486);
nand U4002 (N_4002,In_2672,In_2315);
or U4003 (N_4003,In_1649,In_1530);
xnor U4004 (N_4004,In_392,In_530);
nand U4005 (N_4005,In_2916,In_1375);
or U4006 (N_4006,In_1417,In_2856);
or U4007 (N_4007,In_375,In_201);
nand U4008 (N_4008,In_1077,In_2916);
nand U4009 (N_4009,In_1758,In_731);
nand U4010 (N_4010,In_524,In_2787);
or U4011 (N_4011,In_454,In_575);
or U4012 (N_4012,In_2026,In_2844);
nand U4013 (N_4013,In_445,In_143);
or U4014 (N_4014,In_2648,In_295);
nand U4015 (N_4015,In_467,In_482);
xnor U4016 (N_4016,In_2042,In_2197);
nand U4017 (N_4017,In_85,In_300);
and U4018 (N_4018,In_2608,In_716);
nand U4019 (N_4019,In_861,In_1902);
nor U4020 (N_4020,In_845,In_436);
nand U4021 (N_4021,In_1656,In_1304);
and U4022 (N_4022,In_38,In_1832);
xor U4023 (N_4023,In_29,In_323);
and U4024 (N_4024,In_988,In_1867);
or U4025 (N_4025,In_1650,In_1496);
nor U4026 (N_4026,In_164,In_606);
nand U4027 (N_4027,In_397,In_1473);
nand U4028 (N_4028,In_1839,In_2151);
nand U4029 (N_4029,In_410,In_2334);
or U4030 (N_4030,In_1013,In_2555);
and U4031 (N_4031,In_559,In_183);
nand U4032 (N_4032,In_1675,In_954);
or U4033 (N_4033,In_823,In_336);
nor U4034 (N_4034,In_2223,In_1745);
nand U4035 (N_4035,In_846,In_2556);
nor U4036 (N_4036,In_2650,In_1185);
or U4037 (N_4037,In_2465,In_1772);
and U4038 (N_4038,In_1819,In_2319);
xnor U4039 (N_4039,In_2096,In_1423);
and U4040 (N_4040,In_1898,In_2087);
or U4041 (N_4041,In_23,In_945);
nand U4042 (N_4042,In_1170,In_1685);
nand U4043 (N_4043,In_2674,In_987);
xor U4044 (N_4044,In_1598,In_953);
and U4045 (N_4045,In_2961,In_1727);
nor U4046 (N_4046,In_2924,In_1802);
or U4047 (N_4047,In_1378,In_1847);
and U4048 (N_4048,In_84,In_2573);
nand U4049 (N_4049,In_1491,In_575);
nand U4050 (N_4050,In_2633,In_2882);
nand U4051 (N_4051,In_2533,In_896);
or U4052 (N_4052,In_2204,In_1437);
and U4053 (N_4053,In_1491,In_2449);
and U4054 (N_4054,In_1149,In_2390);
nor U4055 (N_4055,In_306,In_119);
nor U4056 (N_4056,In_1038,In_2153);
nand U4057 (N_4057,In_1476,In_2129);
xnor U4058 (N_4058,In_1988,In_1160);
nand U4059 (N_4059,In_431,In_1322);
or U4060 (N_4060,In_1325,In_1510);
and U4061 (N_4061,In_2217,In_1173);
or U4062 (N_4062,In_2760,In_815);
xor U4063 (N_4063,In_2872,In_2637);
and U4064 (N_4064,In_1629,In_910);
and U4065 (N_4065,In_124,In_102);
or U4066 (N_4066,In_799,In_865);
nor U4067 (N_4067,In_651,In_2605);
and U4068 (N_4068,In_2940,In_2813);
and U4069 (N_4069,In_1758,In_1984);
and U4070 (N_4070,In_1672,In_2162);
nand U4071 (N_4071,In_2786,In_585);
and U4072 (N_4072,In_2030,In_787);
nand U4073 (N_4073,In_1989,In_2540);
nand U4074 (N_4074,In_1743,In_1974);
xor U4075 (N_4075,In_2322,In_2201);
nand U4076 (N_4076,In_2360,In_2874);
nand U4077 (N_4077,In_449,In_1366);
and U4078 (N_4078,In_300,In_1730);
nand U4079 (N_4079,In_2150,In_2210);
nor U4080 (N_4080,In_254,In_1868);
nor U4081 (N_4081,In_426,In_2250);
nor U4082 (N_4082,In_1346,In_389);
or U4083 (N_4083,In_1564,In_103);
nor U4084 (N_4084,In_89,In_783);
xor U4085 (N_4085,In_2344,In_156);
xor U4086 (N_4086,In_1460,In_2245);
nand U4087 (N_4087,In_1429,In_2441);
or U4088 (N_4088,In_1839,In_943);
and U4089 (N_4089,In_1773,In_1275);
nor U4090 (N_4090,In_1865,In_839);
and U4091 (N_4091,In_1740,In_1022);
and U4092 (N_4092,In_1740,In_1765);
xor U4093 (N_4093,In_722,In_354);
or U4094 (N_4094,In_53,In_1700);
or U4095 (N_4095,In_1810,In_2962);
nand U4096 (N_4096,In_2252,In_2283);
and U4097 (N_4097,In_1888,In_1241);
or U4098 (N_4098,In_215,In_61);
or U4099 (N_4099,In_666,In_583);
or U4100 (N_4100,In_127,In_1858);
nor U4101 (N_4101,In_342,In_1882);
xnor U4102 (N_4102,In_1782,In_1944);
nand U4103 (N_4103,In_982,In_1669);
xor U4104 (N_4104,In_2490,In_471);
xor U4105 (N_4105,In_2235,In_2443);
xnor U4106 (N_4106,In_2540,In_1898);
nand U4107 (N_4107,In_1555,In_2456);
and U4108 (N_4108,In_634,In_2008);
xor U4109 (N_4109,In_1066,In_1433);
nor U4110 (N_4110,In_1973,In_1591);
or U4111 (N_4111,In_1536,In_2522);
nor U4112 (N_4112,In_339,In_2307);
nor U4113 (N_4113,In_1858,In_2019);
nor U4114 (N_4114,In_2739,In_1472);
xor U4115 (N_4115,In_2114,In_1873);
and U4116 (N_4116,In_225,In_1071);
and U4117 (N_4117,In_1451,In_1979);
and U4118 (N_4118,In_2486,In_2077);
nor U4119 (N_4119,In_133,In_348);
or U4120 (N_4120,In_1434,In_638);
nand U4121 (N_4121,In_2023,In_2948);
and U4122 (N_4122,In_2725,In_356);
nor U4123 (N_4123,In_1795,In_2573);
nor U4124 (N_4124,In_1286,In_2392);
or U4125 (N_4125,In_2108,In_211);
or U4126 (N_4126,In_2163,In_1828);
and U4127 (N_4127,In_699,In_2134);
nand U4128 (N_4128,In_1235,In_1222);
nor U4129 (N_4129,In_1658,In_1885);
nand U4130 (N_4130,In_2984,In_2615);
xnor U4131 (N_4131,In_2781,In_1495);
nand U4132 (N_4132,In_2534,In_2253);
nand U4133 (N_4133,In_1,In_2855);
nor U4134 (N_4134,In_2796,In_454);
and U4135 (N_4135,In_2034,In_2477);
nand U4136 (N_4136,In_13,In_1689);
nand U4137 (N_4137,In_324,In_1175);
nor U4138 (N_4138,In_933,In_2619);
nor U4139 (N_4139,In_353,In_943);
and U4140 (N_4140,In_639,In_2421);
or U4141 (N_4141,In_1436,In_1102);
or U4142 (N_4142,In_888,In_246);
nor U4143 (N_4143,In_586,In_1743);
nand U4144 (N_4144,In_2445,In_2950);
or U4145 (N_4145,In_2548,In_2537);
nor U4146 (N_4146,In_1261,In_1539);
and U4147 (N_4147,In_767,In_2148);
or U4148 (N_4148,In_1320,In_1186);
nor U4149 (N_4149,In_245,In_944);
or U4150 (N_4150,In_1658,In_2031);
nor U4151 (N_4151,In_2801,In_316);
or U4152 (N_4152,In_2396,In_670);
or U4153 (N_4153,In_740,In_707);
and U4154 (N_4154,In_2339,In_1347);
nor U4155 (N_4155,In_1443,In_2106);
xnor U4156 (N_4156,In_1368,In_1815);
xnor U4157 (N_4157,In_1419,In_291);
xor U4158 (N_4158,In_1439,In_850);
nor U4159 (N_4159,In_2184,In_2597);
nand U4160 (N_4160,In_1615,In_2104);
or U4161 (N_4161,In_160,In_1641);
and U4162 (N_4162,In_481,In_1014);
nand U4163 (N_4163,In_2931,In_2932);
xor U4164 (N_4164,In_163,In_2890);
and U4165 (N_4165,In_163,In_1848);
nand U4166 (N_4166,In_389,In_128);
nand U4167 (N_4167,In_2058,In_124);
or U4168 (N_4168,In_2147,In_2633);
xnor U4169 (N_4169,In_817,In_2538);
nand U4170 (N_4170,In_1012,In_2467);
nor U4171 (N_4171,In_2059,In_118);
nor U4172 (N_4172,In_1807,In_1374);
and U4173 (N_4173,In_921,In_525);
nor U4174 (N_4174,In_2414,In_2023);
nor U4175 (N_4175,In_1243,In_1010);
and U4176 (N_4176,In_66,In_2452);
nand U4177 (N_4177,In_1788,In_483);
or U4178 (N_4178,In_0,In_778);
nor U4179 (N_4179,In_504,In_337);
and U4180 (N_4180,In_2477,In_2995);
and U4181 (N_4181,In_1972,In_1671);
nor U4182 (N_4182,In_404,In_291);
and U4183 (N_4183,In_1520,In_766);
and U4184 (N_4184,In_819,In_615);
or U4185 (N_4185,In_2734,In_2003);
nand U4186 (N_4186,In_2426,In_826);
or U4187 (N_4187,In_1418,In_1448);
xor U4188 (N_4188,In_876,In_2068);
nor U4189 (N_4189,In_2410,In_424);
and U4190 (N_4190,In_954,In_2206);
nand U4191 (N_4191,In_195,In_1087);
nor U4192 (N_4192,In_1816,In_2607);
nor U4193 (N_4193,In_2066,In_1871);
and U4194 (N_4194,In_1829,In_932);
nor U4195 (N_4195,In_2315,In_618);
nand U4196 (N_4196,In_951,In_2234);
nand U4197 (N_4197,In_2644,In_2103);
nor U4198 (N_4198,In_723,In_522);
or U4199 (N_4199,In_2343,In_1473);
nand U4200 (N_4200,In_40,In_1656);
nor U4201 (N_4201,In_537,In_1576);
and U4202 (N_4202,In_1199,In_2812);
nand U4203 (N_4203,In_1963,In_1207);
and U4204 (N_4204,In_2283,In_2272);
nor U4205 (N_4205,In_237,In_128);
or U4206 (N_4206,In_915,In_2503);
nand U4207 (N_4207,In_2016,In_1943);
nand U4208 (N_4208,In_852,In_177);
and U4209 (N_4209,In_1125,In_2522);
and U4210 (N_4210,In_1560,In_33);
xnor U4211 (N_4211,In_1266,In_482);
and U4212 (N_4212,In_1527,In_1713);
nor U4213 (N_4213,In_2497,In_1984);
and U4214 (N_4214,In_2993,In_1104);
or U4215 (N_4215,In_2321,In_1537);
nor U4216 (N_4216,In_2199,In_1373);
nand U4217 (N_4217,In_544,In_403);
and U4218 (N_4218,In_1923,In_1156);
nand U4219 (N_4219,In_926,In_354);
xor U4220 (N_4220,In_2332,In_2166);
nand U4221 (N_4221,In_1710,In_1724);
and U4222 (N_4222,In_1727,In_114);
nor U4223 (N_4223,In_1006,In_2027);
and U4224 (N_4224,In_1441,In_517);
or U4225 (N_4225,In_9,In_1146);
nand U4226 (N_4226,In_1817,In_2206);
nor U4227 (N_4227,In_2059,In_854);
xnor U4228 (N_4228,In_2180,In_2332);
nand U4229 (N_4229,In_503,In_1808);
nor U4230 (N_4230,In_1201,In_1021);
and U4231 (N_4231,In_2693,In_229);
nor U4232 (N_4232,In_523,In_2194);
or U4233 (N_4233,In_2385,In_2913);
nand U4234 (N_4234,In_2689,In_1170);
nor U4235 (N_4235,In_2286,In_2870);
and U4236 (N_4236,In_2804,In_1143);
or U4237 (N_4237,In_1492,In_2388);
nand U4238 (N_4238,In_2567,In_1987);
nand U4239 (N_4239,In_2069,In_627);
nand U4240 (N_4240,In_2953,In_1102);
nand U4241 (N_4241,In_1771,In_2168);
and U4242 (N_4242,In_782,In_93);
or U4243 (N_4243,In_1636,In_1380);
and U4244 (N_4244,In_2543,In_2884);
nand U4245 (N_4245,In_1098,In_2597);
nand U4246 (N_4246,In_1065,In_886);
or U4247 (N_4247,In_2094,In_976);
nand U4248 (N_4248,In_1500,In_1520);
and U4249 (N_4249,In_1483,In_145);
nor U4250 (N_4250,In_2731,In_1754);
nand U4251 (N_4251,In_2702,In_274);
nand U4252 (N_4252,In_321,In_1755);
or U4253 (N_4253,In_525,In_2795);
and U4254 (N_4254,In_1625,In_2188);
and U4255 (N_4255,In_1659,In_2594);
and U4256 (N_4256,In_2625,In_2023);
or U4257 (N_4257,In_1125,In_2887);
and U4258 (N_4258,In_1407,In_2066);
or U4259 (N_4259,In_655,In_2658);
and U4260 (N_4260,In_1391,In_2279);
xnor U4261 (N_4261,In_314,In_2785);
nand U4262 (N_4262,In_2365,In_224);
nand U4263 (N_4263,In_412,In_2566);
nor U4264 (N_4264,In_2007,In_2067);
nor U4265 (N_4265,In_387,In_2797);
and U4266 (N_4266,In_42,In_762);
xnor U4267 (N_4267,In_1052,In_195);
nand U4268 (N_4268,In_330,In_1569);
xnor U4269 (N_4269,In_680,In_1538);
xnor U4270 (N_4270,In_231,In_886);
nor U4271 (N_4271,In_2046,In_2583);
and U4272 (N_4272,In_2165,In_2701);
and U4273 (N_4273,In_2765,In_2582);
nor U4274 (N_4274,In_1479,In_739);
nor U4275 (N_4275,In_595,In_1408);
and U4276 (N_4276,In_701,In_227);
or U4277 (N_4277,In_203,In_2803);
xor U4278 (N_4278,In_1490,In_1018);
nand U4279 (N_4279,In_1514,In_516);
and U4280 (N_4280,In_1052,In_958);
and U4281 (N_4281,In_140,In_1493);
or U4282 (N_4282,In_2449,In_2564);
or U4283 (N_4283,In_955,In_1223);
and U4284 (N_4284,In_2105,In_1326);
or U4285 (N_4285,In_414,In_1496);
or U4286 (N_4286,In_1766,In_61);
nand U4287 (N_4287,In_908,In_356);
nand U4288 (N_4288,In_2658,In_43);
or U4289 (N_4289,In_2244,In_1834);
and U4290 (N_4290,In_1407,In_1211);
xnor U4291 (N_4291,In_1665,In_1630);
xnor U4292 (N_4292,In_2368,In_587);
and U4293 (N_4293,In_1841,In_681);
nand U4294 (N_4294,In_398,In_417);
nand U4295 (N_4295,In_2322,In_2174);
nor U4296 (N_4296,In_1688,In_2608);
and U4297 (N_4297,In_2500,In_1894);
or U4298 (N_4298,In_24,In_2582);
xor U4299 (N_4299,In_2479,In_2428);
nor U4300 (N_4300,In_1284,In_439);
xor U4301 (N_4301,In_260,In_1992);
or U4302 (N_4302,In_1806,In_1882);
and U4303 (N_4303,In_538,In_1452);
nor U4304 (N_4304,In_1493,In_1061);
nand U4305 (N_4305,In_68,In_2880);
and U4306 (N_4306,In_1389,In_2749);
and U4307 (N_4307,In_1145,In_945);
nand U4308 (N_4308,In_2752,In_2809);
or U4309 (N_4309,In_659,In_2131);
nor U4310 (N_4310,In_2092,In_1054);
and U4311 (N_4311,In_219,In_1262);
or U4312 (N_4312,In_2097,In_2808);
nor U4313 (N_4313,In_2575,In_2985);
and U4314 (N_4314,In_2006,In_2815);
or U4315 (N_4315,In_2364,In_897);
and U4316 (N_4316,In_423,In_2429);
xor U4317 (N_4317,In_1381,In_1400);
or U4318 (N_4318,In_2778,In_2434);
or U4319 (N_4319,In_615,In_112);
nor U4320 (N_4320,In_864,In_2076);
nand U4321 (N_4321,In_278,In_1960);
xnor U4322 (N_4322,In_1408,In_2984);
or U4323 (N_4323,In_149,In_953);
nor U4324 (N_4324,In_85,In_803);
or U4325 (N_4325,In_2987,In_640);
nand U4326 (N_4326,In_1936,In_1352);
or U4327 (N_4327,In_268,In_2681);
and U4328 (N_4328,In_182,In_590);
and U4329 (N_4329,In_2598,In_922);
xor U4330 (N_4330,In_175,In_2856);
nand U4331 (N_4331,In_2487,In_1866);
nor U4332 (N_4332,In_2528,In_1927);
or U4333 (N_4333,In_1526,In_1981);
nand U4334 (N_4334,In_2025,In_2279);
and U4335 (N_4335,In_2398,In_2506);
and U4336 (N_4336,In_1924,In_2418);
and U4337 (N_4337,In_1262,In_152);
nor U4338 (N_4338,In_2718,In_466);
xnor U4339 (N_4339,In_383,In_1587);
nand U4340 (N_4340,In_2688,In_1851);
nor U4341 (N_4341,In_2067,In_209);
nor U4342 (N_4342,In_753,In_1695);
or U4343 (N_4343,In_850,In_2956);
nand U4344 (N_4344,In_325,In_2133);
nand U4345 (N_4345,In_2123,In_541);
nor U4346 (N_4346,In_2128,In_2188);
nand U4347 (N_4347,In_1884,In_1023);
or U4348 (N_4348,In_1428,In_1603);
or U4349 (N_4349,In_1892,In_765);
nand U4350 (N_4350,In_639,In_1803);
nand U4351 (N_4351,In_2625,In_1133);
nor U4352 (N_4352,In_1669,In_2022);
nor U4353 (N_4353,In_497,In_279);
nor U4354 (N_4354,In_1527,In_1529);
nor U4355 (N_4355,In_732,In_580);
nand U4356 (N_4356,In_1856,In_1676);
or U4357 (N_4357,In_1098,In_330);
nor U4358 (N_4358,In_928,In_2153);
and U4359 (N_4359,In_2435,In_2818);
nand U4360 (N_4360,In_697,In_2593);
nor U4361 (N_4361,In_2368,In_2739);
or U4362 (N_4362,In_567,In_1266);
nor U4363 (N_4363,In_211,In_2295);
nor U4364 (N_4364,In_986,In_1816);
nand U4365 (N_4365,In_2746,In_2786);
or U4366 (N_4366,In_243,In_2037);
or U4367 (N_4367,In_448,In_2086);
or U4368 (N_4368,In_321,In_895);
xor U4369 (N_4369,In_1533,In_1297);
nor U4370 (N_4370,In_2854,In_1664);
or U4371 (N_4371,In_220,In_2276);
nand U4372 (N_4372,In_956,In_448);
or U4373 (N_4373,In_1641,In_2245);
xor U4374 (N_4374,In_983,In_470);
nor U4375 (N_4375,In_2071,In_2368);
nand U4376 (N_4376,In_2944,In_2355);
or U4377 (N_4377,In_2402,In_373);
nor U4378 (N_4378,In_756,In_815);
nor U4379 (N_4379,In_398,In_1019);
nor U4380 (N_4380,In_2149,In_1440);
or U4381 (N_4381,In_1854,In_621);
nand U4382 (N_4382,In_2366,In_2715);
xor U4383 (N_4383,In_402,In_304);
nor U4384 (N_4384,In_2689,In_1160);
and U4385 (N_4385,In_2158,In_856);
nor U4386 (N_4386,In_55,In_854);
or U4387 (N_4387,In_2052,In_322);
xor U4388 (N_4388,In_800,In_1566);
nor U4389 (N_4389,In_1361,In_1253);
nor U4390 (N_4390,In_855,In_1810);
nor U4391 (N_4391,In_1042,In_1702);
nor U4392 (N_4392,In_2472,In_449);
or U4393 (N_4393,In_1038,In_2102);
nand U4394 (N_4394,In_1503,In_1443);
nand U4395 (N_4395,In_1931,In_1312);
nand U4396 (N_4396,In_927,In_677);
xor U4397 (N_4397,In_1689,In_553);
nand U4398 (N_4398,In_18,In_2591);
nand U4399 (N_4399,In_1331,In_1419);
nand U4400 (N_4400,In_1169,In_1355);
nor U4401 (N_4401,In_1864,In_1507);
nor U4402 (N_4402,In_1427,In_1440);
nor U4403 (N_4403,In_2216,In_2269);
xnor U4404 (N_4404,In_2149,In_1377);
nand U4405 (N_4405,In_1044,In_2400);
nand U4406 (N_4406,In_537,In_224);
and U4407 (N_4407,In_2378,In_414);
nor U4408 (N_4408,In_1033,In_27);
nand U4409 (N_4409,In_606,In_402);
or U4410 (N_4410,In_163,In_2484);
or U4411 (N_4411,In_2656,In_1100);
or U4412 (N_4412,In_1485,In_924);
or U4413 (N_4413,In_171,In_1661);
nand U4414 (N_4414,In_1008,In_1329);
nor U4415 (N_4415,In_49,In_244);
and U4416 (N_4416,In_320,In_710);
nor U4417 (N_4417,In_118,In_2065);
nand U4418 (N_4418,In_2881,In_1648);
and U4419 (N_4419,In_2421,In_1272);
and U4420 (N_4420,In_913,In_2307);
or U4421 (N_4421,In_2218,In_2876);
nor U4422 (N_4422,In_1897,In_2767);
nor U4423 (N_4423,In_2516,In_1663);
and U4424 (N_4424,In_2715,In_1612);
or U4425 (N_4425,In_111,In_1999);
nand U4426 (N_4426,In_668,In_1075);
nor U4427 (N_4427,In_278,In_248);
and U4428 (N_4428,In_1761,In_2404);
or U4429 (N_4429,In_2441,In_1452);
nor U4430 (N_4430,In_2813,In_341);
or U4431 (N_4431,In_1014,In_1102);
nor U4432 (N_4432,In_902,In_2339);
nand U4433 (N_4433,In_1074,In_135);
nand U4434 (N_4434,In_2762,In_6);
and U4435 (N_4435,In_2780,In_1167);
or U4436 (N_4436,In_1652,In_496);
and U4437 (N_4437,In_391,In_451);
and U4438 (N_4438,In_1986,In_2489);
nand U4439 (N_4439,In_640,In_2274);
or U4440 (N_4440,In_2914,In_1633);
or U4441 (N_4441,In_2618,In_2044);
nor U4442 (N_4442,In_2572,In_1915);
or U4443 (N_4443,In_1781,In_2032);
or U4444 (N_4444,In_105,In_1908);
nor U4445 (N_4445,In_2444,In_971);
nor U4446 (N_4446,In_2799,In_498);
or U4447 (N_4447,In_1168,In_376);
nor U4448 (N_4448,In_2001,In_1082);
xnor U4449 (N_4449,In_1072,In_897);
nor U4450 (N_4450,In_2992,In_946);
or U4451 (N_4451,In_2096,In_1410);
nor U4452 (N_4452,In_1932,In_1436);
or U4453 (N_4453,In_913,In_1976);
nor U4454 (N_4454,In_1682,In_2596);
or U4455 (N_4455,In_993,In_1368);
nor U4456 (N_4456,In_1758,In_2050);
nand U4457 (N_4457,In_1282,In_2799);
nand U4458 (N_4458,In_643,In_2940);
or U4459 (N_4459,In_2439,In_2299);
and U4460 (N_4460,In_1725,In_1386);
nand U4461 (N_4461,In_2606,In_2936);
and U4462 (N_4462,In_233,In_1049);
nor U4463 (N_4463,In_2247,In_2143);
nor U4464 (N_4464,In_1005,In_444);
or U4465 (N_4465,In_1805,In_2856);
and U4466 (N_4466,In_2809,In_655);
and U4467 (N_4467,In_706,In_103);
or U4468 (N_4468,In_117,In_907);
nand U4469 (N_4469,In_2717,In_1335);
and U4470 (N_4470,In_1974,In_1776);
xnor U4471 (N_4471,In_1559,In_1280);
and U4472 (N_4472,In_1966,In_886);
and U4473 (N_4473,In_1157,In_2371);
nand U4474 (N_4474,In_400,In_1474);
nand U4475 (N_4475,In_896,In_2837);
nand U4476 (N_4476,In_910,In_183);
nand U4477 (N_4477,In_534,In_16);
or U4478 (N_4478,In_565,In_2254);
and U4479 (N_4479,In_1424,In_2683);
or U4480 (N_4480,In_119,In_327);
and U4481 (N_4481,In_2558,In_1207);
and U4482 (N_4482,In_2214,In_328);
or U4483 (N_4483,In_1468,In_2922);
nand U4484 (N_4484,In_1000,In_805);
or U4485 (N_4485,In_2837,In_1625);
or U4486 (N_4486,In_2682,In_1347);
nand U4487 (N_4487,In_1804,In_1329);
nand U4488 (N_4488,In_2162,In_496);
xor U4489 (N_4489,In_2880,In_933);
nor U4490 (N_4490,In_1633,In_686);
nand U4491 (N_4491,In_2350,In_2160);
xnor U4492 (N_4492,In_1728,In_688);
nor U4493 (N_4493,In_2222,In_1803);
nand U4494 (N_4494,In_2539,In_1679);
nor U4495 (N_4495,In_1714,In_1475);
nor U4496 (N_4496,In_2303,In_2827);
and U4497 (N_4497,In_99,In_1322);
or U4498 (N_4498,In_1759,In_332);
and U4499 (N_4499,In_334,In_2620);
or U4500 (N_4500,In_2001,In_2832);
or U4501 (N_4501,In_2555,In_152);
or U4502 (N_4502,In_89,In_1576);
and U4503 (N_4503,In_1283,In_2435);
and U4504 (N_4504,In_654,In_380);
or U4505 (N_4505,In_2954,In_2073);
or U4506 (N_4506,In_1481,In_2062);
nor U4507 (N_4507,In_132,In_1094);
nand U4508 (N_4508,In_159,In_2478);
or U4509 (N_4509,In_2700,In_620);
or U4510 (N_4510,In_2517,In_330);
and U4511 (N_4511,In_667,In_2219);
xnor U4512 (N_4512,In_344,In_592);
nor U4513 (N_4513,In_724,In_2627);
or U4514 (N_4514,In_492,In_140);
and U4515 (N_4515,In_2517,In_1796);
nand U4516 (N_4516,In_2420,In_890);
and U4517 (N_4517,In_1558,In_1958);
and U4518 (N_4518,In_163,In_2214);
or U4519 (N_4519,In_2089,In_2091);
nor U4520 (N_4520,In_676,In_560);
and U4521 (N_4521,In_1772,In_2321);
nor U4522 (N_4522,In_2214,In_2317);
nand U4523 (N_4523,In_2937,In_227);
and U4524 (N_4524,In_2844,In_2935);
nand U4525 (N_4525,In_474,In_2322);
and U4526 (N_4526,In_1451,In_1603);
and U4527 (N_4527,In_1912,In_1890);
or U4528 (N_4528,In_7,In_1406);
and U4529 (N_4529,In_1084,In_2793);
and U4530 (N_4530,In_1856,In_1270);
and U4531 (N_4531,In_823,In_2896);
xor U4532 (N_4532,In_1206,In_1285);
nor U4533 (N_4533,In_1761,In_900);
or U4534 (N_4534,In_145,In_1646);
xnor U4535 (N_4535,In_2729,In_2647);
nand U4536 (N_4536,In_1334,In_828);
nand U4537 (N_4537,In_843,In_501);
nor U4538 (N_4538,In_2236,In_1413);
or U4539 (N_4539,In_1148,In_1408);
nand U4540 (N_4540,In_1974,In_120);
nand U4541 (N_4541,In_632,In_1104);
nand U4542 (N_4542,In_2882,In_2810);
nand U4543 (N_4543,In_51,In_1584);
xor U4544 (N_4544,In_1910,In_2731);
nor U4545 (N_4545,In_2872,In_1170);
or U4546 (N_4546,In_863,In_271);
or U4547 (N_4547,In_2688,In_2636);
or U4548 (N_4548,In_2527,In_1893);
nand U4549 (N_4549,In_1987,In_730);
or U4550 (N_4550,In_79,In_211);
nand U4551 (N_4551,In_2701,In_1138);
nand U4552 (N_4552,In_2838,In_2203);
nand U4553 (N_4553,In_268,In_2420);
and U4554 (N_4554,In_946,In_565);
nand U4555 (N_4555,In_1754,In_1998);
nor U4556 (N_4556,In_721,In_2680);
nor U4557 (N_4557,In_1338,In_2607);
or U4558 (N_4558,In_1444,In_2895);
nor U4559 (N_4559,In_169,In_495);
nor U4560 (N_4560,In_612,In_1734);
nor U4561 (N_4561,In_1195,In_1960);
nor U4562 (N_4562,In_165,In_575);
nand U4563 (N_4563,In_650,In_305);
or U4564 (N_4564,In_1520,In_1373);
and U4565 (N_4565,In_1912,In_2917);
and U4566 (N_4566,In_272,In_1637);
or U4567 (N_4567,In_311,In_1390);
nor U4568 (N_4568,In_1435,In_2636);
xnor U4569 (N_4569,In_1065,In_1384);
or U4570 (N_4570,In_2562,In_1033);
and U4571 (N_4571,In_1446,In_2815);
nand U4572 (N_4572,In_2862,In_2215);
nand U4573 (N_4573,In_2180,In_1974);
nand U4574 (N_4574,In_1848,In_883);
or U4575 (N_4575,In_1727,In_572);
nor U4576 (N_4576,In_1221,In_636);
nor U4577 (N_4577,In_286,In_2028);
xnor U4578 (N_4578,In_2559,In_59);
nor U4579 (N_4579,In_2660,In_1440);
nand U4580 (N_4580,In_889,In_2501);
nand U4581 (N_4581,In_1663,In_226);
and U4582 (N_4582,In_2622,In_1734);
nor U4583 (N_4583,In_2186,In_359);
and U4584 (N_4584,In_39,In_743);
or U4585 (N_4585,In_2458,In_2514);
nor U4586 (N_4586,In_2389,In_959);
or U4587 (N_4587,In_837,In_74);
and U4588 (N_4588,In_2986,In_1149);
or U4589 (N_4589,In_1342,In_2630);
or U4590 (N_4590,In_752,In_1645);
nor U4591 (N_4591,In_11,In_2406);
nand U4592 (N_4592,In_2409,In_1716);
nand U4593 (N_4593,In_2573,In_15);
nand U4594 (N_4594,In_120,In_2698);
and U4595 (N_4595,In_1621,In_2009);
nor U4596 (N_4596,In_369,In_2613);
or U4597 (N_4597,In_2492,In_899);
nand U4598 (N_4598,In_2727,In_869);
nand U4599 (N_4599,In_2061,In_1335);
nand U4600 (N_4600,In_1215,In_1461);
nor U4601 (N_4601,In_1674,In_360);
or U4602 (N_4602,In_1166,In_2108);
and U4603 (N_4603,In_894,In_2827);
nand U4604 (N_4604,In_2064,In_2290);
nor U4605 (N_4605,In_1049,In_1828);
nand U4606 (N_4606,In_2187,In_1463);
nand U4607 (N_4607,In_694,In_709);
nand U4608 (N_4608,In_1603,In_531);
and U4609 (N_4609,In_228,In_585);
and U4610 (N_4610,In_2757,In_604);
and U4611 (N_4611,In_793,In_1420);
nand U4612 (N_4612,In_2932,In_2383);
nand U4613 (N_4613,In_1921,In_2401);
and U4614 (N_4614,In_1450,In_2821);
nor U4615 (N_4615,In_1728,In_453);
or U4616 (N_4616,In_2135,In_2636);
nor U4617 (N_4617,In_2809,In_2330);
xnor U4618 (N_4618,In_1502,In_991);
nor U4619 (N_4619,In_352,In_1945);
nor U4620 (N_4620,In_2107,In_2033);
xor U4621 (N_4621,In_1196,In_199);
or U4622 (N_4622,In_2142,In_2775);
and U4623 (N_4623,In_1728,In_1782);
or U4624 (N_4624,In_2779,In_1781);
or U4625 (N_4625,In_1295,In_288);
nor U4626 (N_4626,In_921,In_834);
and U4627 (N_4627,In_1273,In_1397);
and U4628 (N_4628,In_245,In_1327);
nand U4629 (N_4629,In_2627,In_826);
xor U4630 (N_4630,In_1728,In_1513);
nor U4631 (N_4631,In_945,In_1998);
nor U4632 (N_4632,In_2771,In_1701);
nor U4633 (N_4633,In_1522,In_1944);
xor U4634 (N_4634,In_2848,In_697);
nand U4635 (N_4635,In_1309,In_2626);
xor U4636 (N_4636,In_777,In_2876);
nand U4637 (N_4637,In_2046,In_2749);
nand U4638 (N_4638,In_162,In_2498);
nor U4639 (N_4639,In_1259,In_2275);
or U4640 (N_4640,In_2663,In_2118);
xnor U4641 (N_4641,In_216,In_388);
nor U4642 (N_4642,In_707,In_2448);
and U4643 (N_4643,In_954,In_2751);
nor U4644 (N_4644,In_2759,In_632);
nand U4645 (N_4645,In_1064,In_2454);
and U4646 (N_4646,In_1525,In_2984);
and U4647 (N_4647,In_2959,In_1262);
xnor U4648 (N_4648,In_1417,In_1496);
and U4649 (N_4649,In_1441,In_692);
xnor U4650 (N_4650,In_2120,In_2762);
nand U4651 (N_4651,In_1948,In_1048);
nand U4652 (N_4652,In_2833,In_738);
nor U4653 (N_4653,In_2086,In_2390);
nor U4654 (N_4654,In_688,In_576);
and U4655 (N_4655,In_1455,In_2681);
xnor U4656 (N_4656,In_1065,In_159);
xnor U4657 (N_4657,In_2927,In_1956);
xnor U4658 (N_4658,In_1343,In_218);
or U4659 (N_4659,In_360,In_308);
nand U4660 (N_4660,In_1105,In_1033);
xnor U4661 (N_4661,In_2857,In_682);
nand U4662 (N_4662,In_298,In_2706);
or U4663 (N_4663,In_635,In_167);
and U4664 (N_4664,In_2965,In_1416);
nand U4665 (N_4665,In_1629,In_1964);
nor U4666 (N_4666,In_2198,In_363);
and U4667 (N_4667,In_2989,In_1919);
nor U4668 (N_4668,In_1742,In_1240);
or U4669 (N_4669,In_360,In_86);
nor U4670 (N_4670,In_1538,In_2418);
or U4671 (N_4671,In_950,In_2933);
nor U4672 (N_4672,In_991,In_925);
nor U4673 (N_4673,In_2490,In_418);
nor U4674 (N_4674,In_2532,In_2778);
xor U4675 (N_4675,In_1464,In_1758);
nand U4676 (N_4676,In_1651,In_162);
or U4677 (N_4677,In_2267,In_2992);
nor U4678 (N_4678,In_1143,In_2550);
nor U4679 (N_4679,In_2330,In_1278);
xor U4680 (N_4680,In_2109,In_1870);
or U4681 (N_4681,In_2092,In_2006);
or U4682 (N_4682,In_120,In_151);
or U4683 (N_4683,In_2661,In_1661);
xor U4684 (N_4684,In_482,In_468);
nand U4685 (N_4685,In_317,In_1146);
and U4686 (N_4686,In_2920,In_2714);
nand U4687 (N_4687,In_55,In_405);
nand U4688 (N_4688,In_876,In_1087);
nand U4689 (N_4689,In_2840,In_2312);
nand U4690 (N_4690,In_2178,In_1531);
nor U4691 (N_4691,In_1495,In_1665);
nor U4692 (N_4692,In_1675,In_883);
xnor U4693 (N_4693,In_856,In_288);
nor U4694 (N_4694,In_444,In_1833);
and U4695 (N_4695,In_2334,In_720);
and U4696 (N_4696,In_2141,In_1030);
nand U4697 (N_4697,In_1014,In_2689);
and U4698 (N_4698,In_2816,In_2275);
xor U4699 (N_4699,In_2714,In_233);
and U4700 (N_4700,In_1929,In_1557);
nand U4701 (N_4701,In_2798,In_1011);
and U4702 (N_4702,In_379,In_1832);
nor U4703 (N_4703,In_1504,In_2887);
or U4704 (N_4704,In_1571,In_2504);
nand U4705 (N_4705,In_247,In_1490);
and U4706 (N_4706,In_2366,In_45);
or U4707 (N_4707,In_405,In_2591);
or U4708 (N_4708,In_2783,In_1993);
and U4709 (N_4709,In_741,In_63);
or U4710 (N_4710,In_1961,In_1568);
nand U4711 (N_4711,In_689,In_1877);
nor U4712 (N_4712,In_293,In_2223);
or U4713 (N_4713,In_1353,In_2610);
nor U4714 (N_4714,In_543,In_975);
nor U4715 (N_4715,In_804,In_2611);
nor U4716 (N_4716,In_2496,In_1788);
nand U4717 (N_4717,In_2495,In_2684);
nor U4718 (N_4718,In_1751,In_1382);
or U4719 (N_4719,In_853,In_603);
or U4720 (N_4720,In_1691,In_2978);
nand U4721 (N_4721,In_850,In_811);
and U4722 (N_4722,In_583,In_581);
xnor U4723 (N_4723,In_523,In_942);
nand U4724 (N_4724,In_2027,In_365);
nor U4725 (N_4725,In_2663,In_2283);
and U4726 (N_4726,In_834,In_852);
nand U4727 (N_4727,In_836,In_144);
nor U4728 (N_4728,In_1771,In_2588);
and U4729 (N_4729,In_1777,In_707);
nor U4730 (N_4730,In_2034,In_2778);
xor U4731 (N_4731,In_2578,In_84);
or U4732 (N_4732,In_1335,In_2264);
nand U4733 (N_4733,In_478,In_173);
and U4734 (N_4734,In_432,In_2931);
nor U4735 (N_4735,In_545,In_1066);
and U4736 (N_4736,In_2533,In_214);
nand U4737 (N_4737,In_1616,In_945);
nand U4738 (N_4738,In_2528,In_860);
and U4739 (N_4739,In_2180,In_1425);
nor U4740 (N_4740,In_2114,In_1720);
xnor U4741 (N_4741,In_1587,In_2716);
or U4742 (N_4742,In_982,In_2081);
nor U4743 (N_4743,In_1282,In_2288);
nor U4744 (N_4744,In_2406,In_2807);
and U4745 (N_4745,In_103,In_1192);
xor U4746 (N_4746,In_593,In_1679);
nand U4747 (N_4747,In_2825,In_2281);
xnor U4748 (N_4748,In_1212,In_1852);
nand U4749 (N_4749,In_2167,In_2492);
nor U4750 (N_4750,In_43,In_2663);
or U4751 (N_4751,In_2304,In_1321);
and U4752 (N_4752,In_831,In_1116);
nand U4753 (N_4753,In_2912,In_2002);
or U4754 (N_4754,In_1706,In_325);
xor U4755 (N_4755,In_1617,In_1001);
and U4756 (N_4756,In_749,In_2506);
and U4757 (N_4757,In_975,In_342);
or U4758 (N_4758,In_1118,In_1042);
xnor U4759 (N_4759,In_349,In_2925);
and U4760 (N_4760,In_542,In_844);
nor U4761 (N_4761,In_784,In_1912);
or U4762 (N_4762,In_741,In_801);
or U4763 (N_4763,In_458,In_397);
or U4764 (N_4764,In_2950,In_2958);
and U4765 (N_4765,In_991,In_1363);
or U4766 (N_4766,In_335,In_50);
nand U4767 (N_4767,In_1466,In_1947);
nand U4768 (N_4768,In_365,In_1421);
and U4769 (N_4769,In_2764,In_181);
and U4770 (N_4770,In_971,In_1985);
nor U4771 (N_4771,In_2043,In_2285);
nand U4772 (N_4772,In_1157,In_1944);
and U4773 (N_4773,In_690,In_1194);
and U4774 (N_4774,In_454,In_492);
nand U4775 (N_4775,In_1334,In_378);
xnor U4776 (N_4776,In_2991,In_58);
nor U4777 (N_4777,In_1077,In_1892);
xnor U4778 (N_4778,In_1414,In_638);
xor U4779 (N_4779,In_1289,In_765);
or U4780 (N_4780,In_1882,In_1511);
and U4781 (N_4781,In_2570,In_2584);
or U4782 (N_4782,In_579,In_19);
xor U4783 (N_4783,In_27,In_1096);
nand U4784 (N_4784,In_1553,In_1692);
or U4785 (N_4785,In_1544,In_752);
nand U4786 (N_4786,In_1724,In_103);
nor U4787 (N_4787,In_2728,In_195);
or U4788 (N_4788,In_1229,In_939);
nor U4789 (N_4789,In_2747,In_149);
or U4790 (N_4790,In_82,In_1498);
and U4791 (N_4791,In_2709,In_2030);
and U4792 (N_4792,In_2156,In_1559);
and U4793 (N_4793,In_2075,In_823);
or U4794 (N_4794,In_146,In_1252);
or U4795 (N_4795,In_1696,In_1955);
nor U4796 (N_4796,In_2617,In_2695);
and U4797 (N_4797,In_626,In_485);
and U4798 (N_4798,In_530,In_544);
or U4799 (N_4799,In_2849,In_377);
or U4800 (N_4800,In_2717,In_1215);
or U4801 (N_4801,In_1708,In_1469);
and U4802 (N_4802,In_2041,In_2658);
xor U4803 (N_4803,In_1462,In_2529);
xor U4804 (N_4804,In_378,In_26);
and U4805 (N_4805,In_1238,In_2779);
xor U4806 (N_4806,In_791,In_1556);
nand U4807 (N_4807,In_1829,In_1132);
and U4808 (N_4808,In_364,In_2067);
or U4809 (N_4809,In_29,In_796);
nand U4810 (N_4810,In_1616,In_983);
nor U4811 (N_4811,In_302,In_1581);
nor U4812 (N_4812,In_33,In_81);
nor U4813 (N_4813,In_2622,In_2519);
nor U4814 (N_4814,In_954,In_2058);
or U4815 (N_4815,In_559,In_350);
and U4816 (N_4816,In_2730,In_1199);
nor U4817 (N_4817,In_2135,In_2230);
xnor U4818 (N_4818,In_2887,In_1849);
or U4819 (N_4819,In_2045,In_112);
and U4820 (N_4820,In_1575,In_646);
nand U4821 (N_4821,In_1455,In_2329);
and U4822 (N_4822,In_2127,In_1129);
nor U4823 (N_4823,In_2088,In_861);
nor U4824 (N_4824,In_1497,In_407);
xnor U4825 (N_4825,In_2188,In_2214);
and U4826 (N_4826,In_2734,In_2778);
nor U4827 (N_4827,In_1564,In_739);
or U4828 (N_4828,In_2771,In_425);
nand U4829 (N_4829,In_932,In_73);
and U4830 (N_4830,In_1316,In_920);
and U4831 (N_4831,In_1621,In_2755);
nand U4832 (N_4832,In_1955,In_2685);
or U4833 (N_4833,In_1314,In_1753);
or U4834 (N_4834,In_2606,In_1795);
and U4835 (N_4835,In_85,In_2609);
nor U4836 (N_4836,In_1804,In_2288);
or U4837 (N_4837,In_1519,In_2352);
and U4838 (N_4838,In_2071,In_1998);
or U4839 (N_4839,In_422,In_2197);
and U4840 (N_4840,In_1280,In_26);
and U4841 (N_4841,In_126,In_1282);
xor U4842 (N_4842,In_1011,In_2284);
nor U4843 (N_4843,In_875,In_1166);
and U4844 (N_4844,In_2398,In_1947);
nor U4845 (N_4845,In_1586,In_2461);
nor U4846 (N_4846,In_1476,In_502);
or U4847 (N_4847,In_2919,In_1256);
nor U4848 (N_4848,In_1904,In_443);
nor U4849 (N_4849,In_2725,In_1942);
nor U4850 (N_4850,In_108,In_2880);
or U4851 (N_4851,In_2327,In_2562);
and U4852 (N_4852,In_1956,In_1746);
and U4853 (N_4853,In_2191,In_1073);
or U4854 (N_4854,In_2579,In_2322);
nand U4855 (N_4855,In_1851,In_901);
xor U4856 (N_4856,In_2183,In_679);
nand U4857 (N_4857,In_112,In_2475);
nor U4858 (N_4858,In_2066,In_1431);
nand U4859 (N_4859,In_359,In_2724);
nand U4860 (N_4860,In_2176,In_70);
or U4861 (N_4861,In_816,In_2478);
xnor U4862 (N_4862,In_586,In_1887);
xor U4863 (N_4863,In_2407,In_1405);
nand U4864 (N_4864,In_631,In_1993);
nand U4865 (N_4865,In_1843,In_1758);
nand U4866 (N_4866,In_1804,In_413);
or U4867 (N_4867,In_158,In_2011);
nor U4868 (N_4868,In_459,In_131);
nor U4869 (N_4869,In_625,In_539);
and U4870 (N_4870,In_2846,In_1056);
or U4871 (N_4871,In_2868,In_2290);
nand U4872 (N_4872,In_986,In_1875);
nor U4873 (N_4873,In_470,In_1052);
and U4874 (N_4874,In_2088,In_2252);
and U4875 (N_4875,In_1801,In_546);
or U4876 (N_4876,In_2116,In_932);
nand U4877 (N_4877,In_514,In_2290);
nor U4878 (N_4878,In_279,In_2573);
or U4879 (N_4879,In_1456,In_2452);
or U4880 (N_4880,In_296,In_1621);
nor U4881 (N_4881,In_2031,In_1792);
xor U4882 (N_4882,In_2739,In_562);
or U4883 (N_4883,In_581,In_2312);
nor U4884 (N_4884,In_77,In_2577);
and U4885 (N_4885,In_1752,In_1259);
and U4886 (N_4886,In_2449,In_1218);
xor U4887 (N_4887,In_2601,In_440);
or U4888 (N_4888,In_1382,In_2502);
or U4889 (N_4889,In_962,In_2017);
nor U4890 (N_4890,In_1142,In_1926);
nand U4891 (N_4891,In_2581,In_395);
or U4892 (N_4892,In_1947,In_2162);
or U4893 (N_4893,In_1881,In_2623);
xnor U4894 (N_4894,In_1807,In_2260);
xor U4895 (N_4895,In_1296,In_360);
or U4896 (N_4896,In_66,In_2001);
nor U4897 (N_4897,In_533,In_1309);
nand U4898 (N_4898,In_100,In_2053);
or U4899 (N_4899,In_580,In_2412);
nor U4900 (N_4900,In_1273,In_1511);
xor U4901 (N_4901,In_536,In_143);
or U4902 (N_4902,In_1763,In_2843);
nand U4903 (N_4903,In_1453,In_2218);
or U4904 (N_4904,In_1669,In_2521);
xnor U4905 (N_4905,In_415,In_2770);
nand U4906 (N_4906,In_1558,In_2479);
nand U4907 (N_4907,In_2609,In_787);
or U4908 (N_4908,In_2499,In_719);
or U4909 (N_4909,In_1773,In_266);
nor U4910 (N_4910,In_1801,In_1741);
and U4911 (N_4911,In_1415,In_1590);
and U4912 (N_4912,In_1266,In_1687);
or U4913 (N_4913,In_2408,In_745);
or U4914 (N_4914,In_224,In_2126);
or U4915 (N_4915,In_990,In_709);
nand U4916 (N_4916,In_1007,In_1544);
or U4917 (N_4917,In_1196,In_838);
nor U4918 (N_4918,In_12,In_2966);
nand U4919 (N_4919,In_1900,In_484);
or U4920 (N_4920,In_2197,In_2347);
nand U4921 (N_4921,In_355,In_701);
and U4922 (N_4922,In_1731,In_36);
and U4923 (N_4923,In_2119,In_341);
nor U4924 (N_4924,In_1906,In_2836);
nor U4925 (N_4925,In_1526,In_1691);
and U4926 (N_4926,In_1609,In_757);
nor U4927 (N_4927,In_737,In_2912);
and U4928 (N_4928,In_2008,In_488);
nand U4929 (N_4929,In_2341,In_1794);
or U4930 (N_4930,In_628,In_479);
nand U4931 (N_4931,In_1793,In_950);
or U4932 (N_4932,In_435,In_2704);
nor U4933 (N_4933,In_2383,In_318);
nand U4934 (N_4934,In_1062,In_2250);
xnor U4935 (N_4935,In_2525,In_1203);
or U4936 (N_4936,In_2573,In_1152);
or U4937 (N_4937,In_328,In_514);
xnor U4938 (N_4938,In_1300,In_298);
and U4939 (N_4939,In_1254,In_2558);
nand U4940 (N_4940,In_2021,In_703);
nor U4941 (N_4941,In_1491,In_2292);
nor U4942 (N_4942,In_355,In_2424);
and U4943 (N_4943,In_1571,In_2289);
xor U4944 (N_4944,In_280,In_445);
nor U4945 (N_4945,In_1737,In_2567);
xnor U4946 (N_4946,In_1345,In_38);
nand U4947 (N_4947,In_1745,In_249);
or U4948 (N_4948,In_1614,In_1766);
nor U4949 (N_4949,In_2326,In_2726);
and U4950 (N_4950,In_818,In_346);
and U4951 (N_4951,In_2335,In_2331);
xor U4952 (N_4952,In_2265,In_1321);
nor U4953 (N_4953,In_1441,In_609);
or U4954 (N_4954,In_711,In_1051);
xnor U4955 (N_4955,In_651,In_2564);
nand U4956 (N_4956,In_1857,In_187);
xnor U4957 (N_4957,In_2758,In_2589);
nor U4958 (N_4958,In_913,In_1624);
xnor U4959 (N_4959,In_312,In_2488);
or U4960 (N_4960,In_1124,In_551);
nor U4961 (N_4961,In_2370,In_872);
or U4962 (N_4962,In_1417,In_2419);
nor U4963 (N_4963,In_1677,In_2182);
and U4964 (N_4964,In_1082,In_1250);
nand U4965 (N_4965,In_1537,In_1172);
or U4966 (N_4966,In_2142,In_1528);
and U4967 (N_4967,In_1184,In_236);
nand U4968 (N_4968,In_789,In_2336);
nand U4969 (N_4969,In_1055,In_1341);
and U4970 (N_4970,In_1332,In_2768);
nor U4971 (N_4971,In_2297,In_2049);
nor U4972 (N_4972,In_1293,In_2703);
or U4973 (N_4973,In_1092,In_1486);
nand U4974 (N_4974,In_478,In_500);
and U4975 (N_4975,In_346,In_2568);
or U4976 (N_4976,In_484,In_2606);
xor U4977 (N_4977,In_2480,In_1539);
nor U4978 (N_4978,In_721,In_659);
nand U4979 (N_4979,In_786,In_77);
or U4980 (N_4980,In_282,In_552);
or U4981 (N_4981,In_79,In_2769);
and U4982 (N_4982,In_314,In_2);
nor U4983 (N_4983,In_146,In_1390);
nor U4984 (N_4984,In_2773,In_358);
nor U4985 (N_4985,In_1638,In_1289);
nor U4986 (N_4986,In_877,In_622);
nand U4987 (N_4987,In_1648,In_2542);
xnor U4988 (N_4988,In_2315,In_1813);
or U4989 (N_4989,In_367,In_2150);
nor U4990 (N_4990,In_1969,In_1751);
and U4991 (N_4991,In_2086,In_1779);
or U4992 (N_4992,In_1926,In_1550);
and U4993 (N_4993,In_1062,In_610);
xor U4994 (N_4994,In_1804,In_2081);
nor U4995 (N_4995,In_1874,In_1908);
nand U4996 (N_4996,In_204,In_2802);
nor U4997 (N_4997,In_1717,In_1669);
nand U4998 (N_4998,In_2783,In_2265);
and U4999 (N_4999,In_1132,In_1732);
nor U5000 (N_5000,In_2826,In_2051);
nand U5001 (N_5001,In_347,In_163);
and U5002 (N_5002,In_1686,In_380);
nor U5003 (N_5003,In_197,In_2469);
and U5004 (N_5004,In_2791,In_1507);
or U5005 (N_5005,In_755,In_652);
and U5006 (N_5006,In_865,In_642);
nor U5007 (N_5007,In_2830,In_2693);
nor U5008 (N_5008,In_1531,In_22);
or U5009 (N_5009,In_2146,In_2034);
nor U5010 (N_5010,In_282,In_407);
or U5011 (N_5011,In_1915,In_1027);
nand U5012 (N_5012,In_533,In_104);
xor U5013 (N_5013,In_2699,In_1919);
nor U5014 (N_5014,In_304,In_2505);
nand U5015 (N_5015,In_5,In_1558);
nand U5016 (N_5016,In_2563,In_2715);
nand U5017 (N_5017,In_837,In_1557);
nor U5018 (N_5018,In_1320,In_807);
nand U5019 (N_5019,In_910,In_1889);
and U5020 (N_5020,In_1047,In_2054);
and U5021 (N_5021,In_2149,In_905);
or U5022 (N_5022,In_1190,In_2190);
nor U5023 (N_5023,In_2957,In_286);
nor U5024 (N_5024,In_155,In_1790);
or U5025 (N_5025,In_1529,In_2581);
and U5026 (N_5026,In_2843,In_1764);
nor U5027 (N_5027,In_2689,In_1596);
or U5028 (N_5028,In_314,In_1284);
or U5029 (N_5029,In_2727,In_175);
nor U5030 (N_5030,In_622,In_90);
nor U5031 (N_5031,In_446,In_1209);
nor U5032 (N_5032,In_1709,In_479);
nor U5033 (N_5033,In_2230,In_2860);
nor U5034 (N_5034,In_2874,In_1874);
or U5035 (N_5035,In_1825,In_2303);
and U5036 (N_5036,In_1868,In_427);
nand U5037 (N_5037,In_1187,In_1562);
and U5038 (N_5038,In_1214,In_1577);
nand U5039 (N_5039,In_2019,In_1188);
nand U5040 (N_5040,In_1429,In_2746);
or U5041 (N_5041,In_1281,In_348);
nand U5042 (N_5042,In_2103,In_2786);
nand U5043 (N_5043,In_2722,In_1393);
or U5044 (N_5044,In_5,In_1025);
nand U5045 (N_5045,In_2578,In_431);
and U5046 (N_5046,In_451,In_982);
or U5047 (N_5047,In_73,In_1699);
nand U5048 (N_5048,In_1447,In_1939);
nor U5049 (N_5049,In_2360,In_1492);
or U5050 (N_5050,In_2556,In_1390);
nand U5051 (N_5051,In_432,In_1450);
and U5052 (N_5052,In_2907,In_222);
nor U5053 (N_5053,In_2362,In_790);
nand U5054 (N_5054,In_2101,In_381);
xnor U5055 (N_5055,In_2512,In_1272);
and U5056 (N_5056,In_1086,In_1166);
or U5057 (N_5057,In_1142,In_2451);
nand U5058 (N_5058,In_2980,In_2887);
or U5059 (N_5059,In_441,In_2816);
or U5060 (N_5060,In_174,In_1872);
and U5061 (N_5061,In_1120,In_2132);
or U5062 (N_5062,In_2063,In_418);
or U5063 (N_5063,In_1364,In_2910);
and U5064 (N_5064,In_137,In_1490);
or U5065 (N_5065,In_1788,In_216);
xor U5066 (N_5066,In_1557,In_2935);
nor U5067 (N_5067,In_2689,In_1970);
or U5068 (N_5068,In_1132,In_2452);
and U5069 (N_5069,In_589,In_762);
nand U5070 (N_5070,In_705,In_2556);
or U5071 (N_5071,In_289,In_732);
nand U5072 (N_5072,In_1405,In_2867);
and U5073 (N_5073,In_1118,In_1443);
xor U5074 (N_5074,In_1966,In_2102);
nand U5075 (N_5075,In_1692,In_921);
xnor U5076 (N_5076,In_1444,In_2597);
xor U5077 (N_5077,In_968,In_56);
xor U5078 (N_5078,In_2513,In_2154);
nand U5079 (N_5079,In_2066,In_2886);
nand U5080 (N_5080,In_1683,In_630);
xor U5081 (N_5081,In_2022,In_2709);
and U5082 (N_5082,In_1516,In_299);
nand U5083 (N_5083,In_748,In_960);
and U5084 (N_5084,In_2314,In_198);
nand U5085 (N_5085,In_2009,In_1246);
nand U5086 (N_5086,In_2792,In_384);
nand U5087 (N_5087,In_732,In_307);
nor U5088 (N_5088,In_411,In_72);
and U5089 (N_5089,In_1661,In_387);
nor U5090 (N_5090,In_422,In_2127);
xnor U5091 (N_5091,In_1469,In_1031);
and U5092 (N_5092,In_539,In_1600);
and U5093 (N_5093,In_715,In_1849);
nand U5094 (N_5094,In_645,In_2951);
nand U5095 (N_5095,In_385,In_242);
or U5096 (N_5096,In_137,In_398);
nand U5097 (N_5097,In_2925,In_1693);
nor U5098 (N_5098,In_2935,In_1769);
nor U5099 (N_5099,In_177,In_769);
nor U5100 (N_5100,In_327,In_224);
or U5101 (N_5101,In_2558,In_2857);
nor U5102 (N_5102,In_1808,In_1553);
or U5103 (N_5103,In_1873,In_2744);
nor U5104 (N_5104,In_1593,In_1011);
nand U5105 (N_5105,In_1915,In_922);
xnor U5106 (N_5106,In_2981,In_2756);
nand U5107 (N_5107,In_1498,In_1395);
and U5108 (N_5108,In_2524,In_197);
nand U5109 (N_5109,In_2640,In_2657);
or U5110 (N_5110,In_2381,In_1668);
nor U5111 (N_5111,In_144,In_1974);
or U5112 (N_5112,In_2350,In_2982);
and U5113 (N_5113,In_766,In_2969);
nor U5114 (N_5114,In_2783,In_945);
xnor U5115 (N_5115,In_850,In_2773);
nor U5116 (N_5116,In_2401,In_1160);
or U5117 (N_5117,In_400,In_1673);
nand U5118 (N_5118,In_2624,In_1121);
nand U5119 (N_5119,In_1169,In_969);
nand U5120 (N_5120,In_79,In_949);
nor U5121 (N_5121,In_1943,In_2567);
nand U5122 (N_5122,In_2404,In_891);
nor U5123 (N_5123,In_1451,In_1149);
nor U5124 (N_5124,In_2150,In_2991);
and U5125 (N_5125,In_2749,In_1841);
and U5126 (N_5126,In_1917,In_2975);
nor U5127 (N_5127,In_745,In_56);
xnor U5128 (N_5128,In_2778,In_617);
nor U5129 (N_5129,In_2322,In_2642);
xor U5130 (N_5130,In_2331,In_1837);
and U5131 (N_5131,In_835,In_2059);
nand U5132 (N_5132,In_1343,In_1892);
and U5133 (N_5133,In_2771,In_2182);
nor U5134 (N_5134,In_2164,In_587);
or U5135 (N_5135,In_786,In_2471);
nor U5136 (N_5136,In_1270,In_660);
nand U5137 (N_5137,In_93,In_1769);
xnor U5138 (N_5138,In_1238,In_2384);
nand U5139 (N_5139,In_2743,In_2163);
nand U5140 (N_5140,In_896,In_1721);
or U5141 (N_5141,In_483,In_2961);
or U5142 (N_5142,In_2207,In_510);
or U5143 (N_5143,In_1931,In_832);
or U5144 (N_5144,In_1743,In_2855);
and U5145 (N_5145,In_979,In_492);
nand U5146 (N_5146,In_2902,In_1982);
and U5147 (N_5147,In_2525,In_2019);
nand U5148 (N_5148,In_2450,In_1369);
and U5149 (N_5149,In_1005,In_1441);
nand U5150 (N_5150,In_1025,In_374);
or U5151 (N_5151,In_869,In_2025);
nand U5152 (N_5152,In_1601,In_998);
and U5153 (N_5153,In_921,In_1500);
and U5154 (N_5154,In_865,In_2073);
nand U5155 (N_5155,In_1145,In_1688);
xnor U5156 (N_5156,In_2870,In_497);
nand U5157 (N_5157,In_2559,In_814);
and U5158 (N_5158,In_95,In_1964);
nand U5159 (N_5159,In_2440,In_1435);
or U5160 (N_5160,In_1209,In_776);
nand U5161 (N_5161,In_742,In_2653);
nor U5162 (N_5162,In_2925,In_2580);
or U5163 (N_5163,In_1210,In_1369);
and U5164 (N_5164,In_1019,In_1907);
nor U5165 (N_5165,In_1008,In_436);
or U5166 (N_5166,In_662,In_1242);
nand U5167 (N_5167,In_2588,In_501);
and U5168 (N_5168,In_1089,In_568);
or U5169 (N_5169,In_1275,In_1020);
nand U5170 (N_5170,In_1061,In_2778);
xnor U5171 (N_5171,In_2202,In_896);
and U5172 (N_5172,In_303,In_2051);
or U5173 (N_5173,In_469,In_764);
nand U5174 (N_5174,In_1801,In_2693);
nand U5175 (N_5175,In_2561,In_2634);
and U5176 (N_5176,In_2466,In_2612);
nor U5177 (N_5177,In_65,In_1959);
or U5178 (N_5178,In_2930,In_2332);
and U5179 (N_5179,In_1262,In_793);
or U5180 (N_5180,In_16,In_947);
xor U5181 (N_5181,In_878,In_2211);
and U5182 (N_5182,In_2535,In_1314);
or U5183 (N_5183,In_1341,In_1631);
or U5184 (N_5184,In_2267,In_2665);
nand U5185 (N_5185,In_1703,In_247);
and U5186 (N_5186,In_161,In_2874);
nor U5187 (N_5187,In_2095,In_775);
nand U5188 (N_5188,In_1512,In_527);
or U5189 (N_5189,In_1212,In_2209);
xor U5190 (N_5190,In_2056,In_2323);
nor U5191 (N_5191,In_2958,In_1104);
and U5192 (N_5192,In_1177,In_1185);
nand U5193 (N_5193,In_2140,In_1529);
nor U5194 (N_5194,In_1988,In_2889);
nand U5195 (N_5195,In_2582,In_109);
and U5196 (N_5196,In_2879,In_2919);
nand U5197 (N_5197,In_259,In_1124);
xnor U5198 (N_5198,In_770,In_661);
nor U5199 (N_5199,In_2114,In_1640);
or U5200 (N_5200,In_130,In_561);
or U5201 (N_5201,In_1177,In_394);
xor U5202 (N_5202,In_306,In_1304);
nand U5203 (N_5203,In_2393,In_1382);
and U5204 (N_5204,In_848,In_2923);
nand U5205 (N_5205,In_2413,In_43);
or U5206 (N_5206,In_2509,In_471);
nand U5207 (N_5207,In_1529,In_2613);
nor U5208 (N_5208,In_2879,In_1822);
nor U5209 (N_5209,In_88,In_2073);
nor U5210 (N_5210,In_2602,In_2238);
nand U5211 (N_5211,In_2912,In_56);
and U5212 (N_5212,In_337,In_2269);
nor U5213 (N_5213,In_289,In_2524);
xor U5214 (N_5214,In_1566,In_1607);
or U5215 (N_5215,In_1020,In_646);
and U5216 (N_5216,In_1610,In_1325);
nand U5217 (N_5217,In_119,In_1549);
or U5218 (N_5218,In_2512,In_2733);
or U5219 (N_5219,In_213,In_1325);
and U5220 (N_5220,In_2610,In_1895);
nand U5221 (N_5221,In_231,In_2757);
and U5222 (N_5222,In_2897,In_233);
or U5223 (N_5223,In_348,In_2790);
nand U5224 (N_5224,In_1354,In_2983);
nor U5225 (N_5225,In_458,In_1095);
and U5226 (N_5226,In_2599,In_2757);
and U5227 (N_5227,In_863,In_2689);
nor U5228 (N_5228,In_1124,In_1367);
or U5229 (N_5229,In_2387,In_1811);
and U5230 (N_5230,In_2879,In_2500);
nand U5231 (N_5231,In_498,In_1654);
and U5232 (N_5232,In_1329,In_39);
or U5233 (N_5233,In_231,In_2689);
nor U5234 (N_5234,In_154,In_2342);
nor U5235 (N_5235,In_2129,In_2167);
nor U5236 (N_5236,In_291,In_2958);
nor U5237 (N_5237,In_1516,In_614);
or U5238 (N_5238,In_2825,In_1113);
and U5239 (N_5239,In_580,In_2571);
nor U5240 (N_5240,In_1716,In_2049);
or U5241 (N_5241,In_701,In_1165);
or U5242 (N_5242,In_1968,In_1429);
and U5243 (N_5243,In_2566,In_1150);
and U5244 (N_5244,In_1881,In_2354);
or U5245 (N_5245,In_2197,In_1643);
or U5246 (N_5246,In_2043,In_551);
and U5247 (N_5247,In_1541,In_474);
or U5248 (N_5248,In_2761,In_1834);
xor U5249 (N_5249,In_2495,In_2415);
xnor U5250 (N_5250,In_978,In_1438);
or U5251 (N_5251,In_2737,In_404);
and U5252 (N_5252,In_2066,In_1691);
nor U5253 (N_5253,In_1967,In_514);
and U5254 (N_5254,In_1156,In_887);
nand U5255 (N_5255,In_1012,In_221);
and U5256 (N_5256,In_616,In_2249);
nor U5257 (N_5257,In_859,In_1957);
nor U5258 (N_5258,In_2306,In_792);
nor U5259 (N_5259,In_1319,In_1359);
nand U5260 (N_5260,In_441,In_1472);
or U5261 (N_5261,In_2087,In_177);
and U5262 (N_5262,In_2280,In_2527);
and U5263 (N_5263,In_1700,In_2464);
and U5264 (N_5264,In_155,In_2821);
and U5265 (N_5265,In_2076,In_2794);
nand U5266 (N_5266,In_475,In_1814);
xnor U5267 (N_5267,In_2631,In_14);
or U5268 (N_5268,In_2162,In_487);
nand U5269 (N_5269,In_2965,In_1977);
xnor U5270 (N_5270,In_260,In_2199);
nor U5271 (N_5271,In_1743,In_996);
nor U5272 (N_5272,In_2389,In_1061);
or U5273 (N_5273,In_1258,In_1498);
nand U5274 (N_5274,In_278,In_2609);
or U5275 (N_5275,In_2907,In_186);
nor U5276 (N_5276,In_458,In_217);
nand U5277 (N_5277,In_649,In_537);
nand U5278 (N_5278,In_1862,In_2814);
nor U5279 (N_5279,In_857,In_263);
nand U5280 (N_5280,In_1777,In_1292);
nor U5281 (N_5281,In_502,In_1863);
or U5282 (N_5282,In_984,In_1452);
nor U5283 (N_5283,In_56,In_1011);
xor U5284 (N_5284,In_1907,In_2214);
or U5285 (N_5285,In_1644,In_1493);
and U5286 (N_5286,In_1656,In_1071);
or U5287 (N_5287,In_608,In_1625);
nand U5288 (N_5288,In_2302,In_2490);
nand U5289 (N_5289,In_2494,In_1670);
or U5290 (N_5290,In_1164,In_1639);
nand U5291 (N_5291,In_685,In_2672);
and U5292 (N_5292,In_2108,In_903);
nand U5293 (N_5293,In_633,In_2044);
nor U5294 (N_5294,In_1016,In_400);
nor U5295 (N_5295,In_1217,In_1113);
nor U5296 (N_5296,In_2817,In_1136);
and U5297 (N_5297,In_1657,In_1928);
nand U5298 (N_5298,In_2484,In_2405);
xnor U5299 (N_5299,In_575,In_1380);
or U5300 (N_5300,In_1607,In_675);
or U5301 (N_5301,In_1801,In_1850);
nand U5302 (N_5302,In_1683,In_1550);
nand U5303 (N_5303,In_263,In_2814);
nor U5304 (N_5304,In_112,In_2460);
nor U5305 (N_5305,In_360,In_133);
nor U5306 (N_5306,In_2011,In_487);
or U5307 (N_5307,In_313,In_1215);
nand U5308 (N_5308,In_518,In_831);
nand U5309 (N_5309,In_1114,In_2849);
nor U5310 (N_5310,In_142,In_1438);
nand U5311 (N_5311,In_723,In_808);
and U5312 (N_5312,In_272,In_2332);
nor U5313 (N_5313,In_1832,In_355);
nand U5314 (N_5314,In_2546,In_666);
nor U5315 (N_5315,In_1517,In_467);
nand U5316 (N_5316,In_2941,In_1412);
nand U5317 (N_5317,In_565,In_2005);
or U5318 (N_5318,In_112,In_326);
and U5319 (N_5319,In_2472,In_1394);
nand U5320 (N_5320,In_1289,In_1960);
nor U5321 (N_5321,In_728,In_2082);
and U5322 (N_5322,In_1365,In_2237);
nor U5323 (N_5323,In_1636,In_2711);
nand U5324 (N_5324,In_2459,In_1954);
or U5325 (N_5325,In_1826,In_2484);
or U5326 (N_5326,In_1988,In_1229);
nand U5327 (N_5327,In_1342,In_2659);
xor U5328 (N_5328,In_2335,In_1186);
or U5329 (N_5329,In_1014,In_429);
nand U5330 (N_5330,In_332,In_562);
or U5331 (N_5331,In_2793,In_2646);
nand U5332 (N_5332,In_822,In_402);
nor U5333 (N_5333,In_2717,In_109);
and U5334 (N_5334,In_1973,In_1101);
and U5335 (N_5335,In_606,In_1000);
nor U5336 (N_5336,In_962,In_885);
nor U5337 (N_5337,In_2610,In_48);
nor U5338 (N_5338,In_132,In_2529);
and U5339 (N_5339,In_15,In_1792);
nand U5340 (N_5340,In_677,In_2072);
nand U5341 (N_5341,In_2047,In_1809);
or U5342 (N_5342,In_1440,In_26);
xnor U5343 (N_5343,In_492,In_670);
and U5344 (N_5344,In_2992,In_546);
xnor U5345 (N_5345,In_1764,In_198);
xnor U5346 (N_5346,In_570,In_1020);
nor U5347 (N_5347,In_2649,In_410);
nand U5348 (N_5348,In_1912,In_651);
xnor U5349 (N_5349,In_2667,In_2701);
and U5350 (N_5350,In_1738,In_2266);
or U5351 (N_5351,In_2719,In_513);
xnor U5352 (N_5352,In_580,In_148);
or U5353 (N_5353,In_2592,In_636);
and U5354 (N_5354,In_363,In_2958);
or U5355 (N_5355,In_319,In_2343);
or U5356 (N_5356,In_1836,In_1892);
nor U5357 (N_5357,In_1793,In_933);
nor U5358 (N_5358,In_750,In_688);
nor U5359 (N_5359,In_1055,In_1065);
nand U5360 (N_5360,In_1847,In_1829);
xor U5361 (N_5361,In_941,In_1475);
and U5362 (N_5362,In_450,In_2496);
xor U5363 (N_5363,In_2885,In_2406);
nor U5364 (N_5364,In_2225,In_159);
nand U5365 (N_5365,In_1820,In_2755);
nor U5366 (N_5366,In_1049,In_1349);
nor U5367 (N_5367,In_243,In_1002);
nor U5368 (N_5368,In_1287,In_2789);
nand U5369 (N_5369,In_2599,In_392);
and U5370 (N_5370,In_217,In_1103);
or U5371 (N_5371,In_600,In_226);
xnor U5372 (N_5372,In_1521,In_1447);
and U5373 (N_5373,In_1802,In_1664);
nand U5374 (N_5374,In_441,In_433);
nor U5375 (N_5375,In_1801,In_2824);
nand U5376 (N_5376,In_864,In_83);
or U5377 (N_5377,In_2313,In_2448);
or U5378 (N_5378,In_2203,In_2613);
nand U5379 (N_5379,In_498,In_104);
or U5380 (N_5380,In_771,In_2460);
nand U5381 (N_5381,In_2297,In_434);
xor U5382 (N_5382,In_883,In_779);
and U5383 (N_5383,In_2730,In_1839);
or U5384 (N_5384,In_2739,In_1220);
and U5385 (N_5385,In_2121,In_2320);
nor U5386 (N_5386,In_277,In_2995);
nor U5387 (N_5387,In_1187,In_2116);
and U5388 (N_5388,In_2654,In_1366);
nand U5389 (N_5389,In_892,In_2527);
xnor U5390 (N_5390,In_1092,In_857);
and U5391 (N_5391,In_1079,In_2752);
or U5392 (N_5392,In_1641,In_2390);
or U5393 (N_5393,In_974,In_1917);
nand U5394 (N_5394,In_1050,In_2503);
nor U5395 (N_5395,In_1384,In_360);
xor U5396 (N_5396,In_1519,In_480);
and U5397 (N_5397,In_2960,In_1408);
nand U5398 (N_5398,In_1391,In_1408);
or U5399 (N_5399,In_2602,In_2944);
or U5400 (N_5400,In_1248,In_1581);
nand U5401 (N_5401,In_650,In_2062);
and U5402 (N_5402,In_2314,In_2911);
and U5403 (N_5403,In_850,In_555);
xor U5404 (N_5404,In_2407,In_2517);
and U5405 (N_5405,In_1148,In_553);
and U5406 (N_5406,In_2572,In_2723);
nand U5407 (N_5407,In_1779,In_1636);
xnor U5408 (N_5408,In_2774,In_1933);
nand U5409 (N_5409,In_988,In_2538);
or U5410 (N_5410,In_2354,In_1412);
and U5411 (N_5411,In_1211,In_2778);
or U5412 (N_5412,In_1470,In_345);
and U5413 (N_5413,In_338,In_1861);
nor U5414 (N_5414,In_1536,In_2550);
xnor U5415 (N_5415,In_2810,In_2405);
and U5416 (N_5416,In_1527,In_2112);
and U5417 (N_5417,In_199,In_619);
nor U5418 (N_5418,In_2819,In_2970);
or U5419 (N_5419,In_1097,In_2271);
or U5420 (N_5420,In_1610,In_39);
or U5421 (N_5421,In_2338,In_109);
nand U5422 (N_5422,In_2137,In_379);
and U5423 (N_5423,In_2186,In_2493);
and U5424 (N_5424,In_2233,In_2250);
nand U5425 (N_5425,In_1282,In_1179);
nor U5426 (N_5426,In_472,In_89);
nand U5427 (N_5427,In_934,In_1848);
and U5428 (N_5428,In_2673,In_1720);
nand U5429 (N_5429,In_1803,In_424);
and U5430 (N_5430,In_827,In_2145);
or U5431 (N_5431,In_1348,In_2787);
and U5432 (N_5432,In_2439,In_274);
or U5433 (N_5433,In_1536,In_2365);
and U5434 (N_5434,In_1105,In_2411);
or U5435 (N_5435,In_2906,In_361);
xor U5436 (N_5436,In_2151,In_298);
or U5437 (N_5437,In_1114,In_1140);
and U5438 (N_5438,In_834,In_620);
nand U5439 (N_5439,In_1449,In_1096);
and U5440 (N_5440,In_2887,In_329);
nand U5441 (N_5441,In_826,In_2410);
or U5442 (N_5442,In_2731,In_1927);
xor U5443 (N_5443,In_1741,In_1037);
and U5444 (N_5444,In_1037,In_1980);
or U5445 (N_5445,In_602,In_1004);
or U5446 (N_5446,In_2921,In_1338);
xnor U5447 (N_5447,In_132,In_1547);
nand U5448 (N_5448,In_353,In_2333);
or U5449 (N_5449,In_1217,In_1408);
and U5450 (N_5450,In_598,In_108);
and U5451 (N_5451,In_1782,In_2408);
nor U5452 (N_5452,In_2771,In_476);
or U5453 (N_5453,In_649,In_1155);
nor U5454 (N_5454,In_1637,In_2047);
or U5455 (N_5455,In_1541,In_1376);
nand U5456 (N_5456,In_663,In_1389);
nor U5457 (N_5457,In_1428,In_2402);
nor U5458 (N_5458,In_2304,In_2038);
nand U5459 (N_5459,In_701,In_2082);
nand U5460 (N_5460,In_2240,In_1132);
nor U5461 (N_5461,In_2492,In_669);
and U5462 (N_5462,In_2872,In_1503);
nor U5463 (N_5463,In_2188,In_1160);
and U5464 (N_5464,In_2053,In_2722);
or U5465 (N_5465,In_2512,In_1623);
nor U5466 (N_5466,In_178,In_1004);
or U5467 (N_5467,In_1239,In_1967);
nand U5468 (N_5468,In_1031,In_2310);
nor U5469 (N_5469,In_2218,In_1668);
and U5470 (N_5470,In_1220,In_297);
and U5471 (N_5471,In_1671,In_28);
and U5472 (N_5472,In_1958,In_231);
nor U5473 (N_5473,In_2588,In_956);
and U5474 (N_5474,In_1352,In_1026);
xnor U5475 (N_5475,In_2237,In_2279);
and U5476 (N_5476,In_1285,In_1694);
or U5477 (N_5477,In_2520,In_1941);
and U5478 (N_5478,In_594,In_314);
and U5479 (N_5479,In_1583,In_1672);
or U5480 (N_5480,In_1573,In_700);
nor U5481 (N_5481,In_834,In_1057);
or U5482 (N_5482,In_4,In_2600);
nand U5483 (N_5483,In_2253,In_1394);
nor U5484 (N_5484,In_1959,In_2894);
or U5485 (N_5485,In_648,In_2692);
nor U5486 (N_5486,In_660,In_2970);
and U5487 (N_5487,In_955,In_132);
and U5488 (N_5488,In_788,In_2691);
nor U5489 (N_5489,In_1966,In_641);
or U5490 (N_5490,In_577,In_2450);
nor U5491 (N_5491,In_2485,In_284);
nand U5492 (N_5492,In_1269,In_1080);
or U5493 (N_5493,In_2537,In_2397);
nand U5494 (N_5494,In_510,In_2884);
or U5495 (N_5495,In_1085,In_1487);
nor U5496 (N_5496,In_1996,In_1642);
nor U5497 (N_5497,In_1998,In_2626);
and U5498 (N_5498,In_1115,In_2416);
nor U5499 (N_5499,In_1354,In_451);
and U5500 (N_5500,In_2077,In_2144);
or U5501 (N_5501,In_235,In_1334);
or U5502 (N_5502,In_1476,In_1484);
nand U5503 (N_5503,In_353,In_1929);
and U5504 (N_5504,In_2926,In_1455);
xor U5505 (N_5505,In_1556,In_1728);
nand U5506 (N_5506,In_1249,In_1598);
or U5507 (N_5507,In_2236,In_1736);
nand U5508 (N_5508,In_1552,In_1014);
nor U5509 (N_5509,In_866,In_1006);
or U5510 (N_5510,In_4,In_1954);
nand U5511 (N_5511,In_605,In_1092);
and U5512 (N_5512,In_1902,In_1812);
xor U5513 (N_5513,In_2290,In_424);
nor U5514 (N_5514,In_313,In_483);
nand U5515 (N_5515,In_2034,In_959);
nor U5516 (N_5516,In_2254,In_1277);
and U5517 (N_5517,In_822,In_2358);
and U5518 (N_5518,In_1793,In_453);
or U5519 (N_5519,In_1747,In_165);
nor U5520 (N_5520,In_2896,In_1487);
or U5521 (N_5521,In_2919,In_479);
and U5522 (N_5522,In_491,In_2370);
and U5523 (N_5523,In_1090,In_83);
and U5524 (N_5524,In_311,In_2539);
and U5525 (N_5525,In_1995,In_2028);
or U5526 (N_5526,In_1621,In_749);
or U5527 (N_5527,In_2304,In_1842);
nor U5528 (N_5528,In_1061,In_435);
xor U5529 (N_5529,In_2280,In_2648);
or U5530 (N_5530,In_1471,In_1961);
nand U5531 (N_5531,In_116,In_1260);
and U5532 (N_5532,In_2003,In_413);
xnor U5533 (N_5533,In_657,In_345);
nor U5534 (N_5534,In_2028,In_2071);
xor U5535 (N_5535,In_129,In_1180);
or U5536 (N_5536,In_1424,In_2671);
nor U5537 (N_5537,In_2479,In_290);
nor U5538 (N_5538,In_855,In_2173);
nor U5539 (N_5539,In_561,In_2126);
nor U5540 (N_5540,In_967,In_384);
or U5541 (N_5541,In_1468,In_213);
or U5542 (N_5542,In_909,In_2841);
xnor U5543 (N_5543,In_2021,In_253);
or U5544 (N_5544,In_846,In_572);
or U5545 (N_5545,In_136,In_2188);
and U5546 (N_5546,In_2153,In_2987);
nand U5547 (N_5547,In_2775,In_2356);
nor U5548 (N_5548,In_581,In_641);
and U5549 (N_5549,In_1710,In_2601);
xor U5550 (N_5550,In_2460,In_2154);
xor U5551 (N_5551,In_1121,In_1551);
nand U5552 (N_5552,In_2651,In_2083);
and U5553 (N_5553,In_1832,In_534);
nor U5554 (N_5554,In_2871,In_932);
and U5555 (N_5555,In_1911,In_1);
or U5556 (N_5556,In_2626,In_2329);
or U5557 (N_5557,In_2155,In_2853);
nor U5558 (N_5558,In_1236,In_2659);
or U5559 (N_5559,In_659,In_2023);
and U5560 (N_5560,In_97,In_2097);
nand U5561 (N_5561,In_1342,In_1512);
nor U5562 (N_5562,In_977,In_1960);
nand U5563 (N_5563,In_935,In_695);
and U5564 (N_5564,In_704,In_2205);
or U5565 (N_5565,In_396,In_1551);
nand U5566 (N_5566,In_650,In_755);
nor U5567 (N_5567,In_1246,In_499);
nand U5568 (N_5568,In_2631,In_1975);
xor U5569 (N_5569,In_1660,In_2866);
nor U5570 (N_5570,In_2179,In_418);
nor U5571 (N_5571,In_972,In_2887);
and U5572 (N_5572,In_1060,In_1625);
nor U5573 (N_5573,In_50,In_2148);
and U5574 (N_5574,In_2529,In_505);
nand U5575 (N_5575,In_1421,In_568);
or U5576 (N_5576,In_1969,In_2764);
nor U5577 (N_5577,In_1472,In_735);
nand U5578 (N_5578,In_2527,In_550);
or U5579 (N_5579,In_1003,In_2238);
nor U5580 (N_5580,In_105,In_2411);
nand U5581 (N_5581,In_1450,In_923);
and U5582 (N_5582,In_1736,In_529);
nand U5583 (N_5583,In_1933,In_1210);
nor U5584 (N_5584,In_2731,In_1872);
or U5585 (N_5585,In_2204,In_2324);
nand U5586 (N_5586,In_1589,In_786);
nor U5587 (N_5587,In_413,In_2364);
xnor U5588 (N_5588,In_1654,In_2127);
nor U5589 (N_5589,In_2697,In_1558);
or U5590 (N_5590,In_1173,In_1107);
nor U5591 (N_5591,In_2570,In_1772);
or U5592 (N_5592,In_2831,In_1342);
and U5593 (N_5593,In_745,In_2056);
nand U5594 (N_5594,In_1071,In_173);
nor U5595 (N_5595,In_2354,In_426);
or U5596 (N_5596,In_6,In_2428);
nand U5597 (N_5597,In_2859,In_971);
nor U5598 (N_5598,In_476,In_963);
nand U5599 (N_5599,In_1974,In_2716);
and U5600 (N_5600,In_525,In_2340);
and U5601 (N_5601,In_1168,In_158);
and U5602 (N_5602,In_1665,In_53);
and U5603 (N_5603,In_1724,In_2939);
or U5604 (N_5604,In_2236,In_662);
nand U5605 (N_5605,In_612,In_64);
or U5606 (N_5606,In_2506,In_2021);
or U5607 (N_5607,In_2977,In_874);
nor U5608 (N_5608,In_1366,In_1167);
nand U5609 (N_5609,In_2686,In_1500);
nand U5610 (N_5610,In_1089,In_979);
and U5611 (N_5611,In_2983,In_1892);
nor U5612 (N_5612,In_2146,In_1970);
or U5613 (N_5613,In_1847,In_2139);
nor U5614 (N_5614,In_2714,In_1023);
or U5615 (N_5615,In_1784,In_295);
or U5616 (N_5616,In_2176,In_99);
or U5617 (N_5617,In_1147,In_346);
nand U5618 (N_5618,In_723,In_795);
and U5619 (N_5619,In_382,In_1855);
nor U5620 (N_5620,In_1751,In_686);
or U5621 (N_5621,In_686,In_918);
and U5622 (N_5622,In_2791,In_2714);
nor U5623 (N_5623,In_1809,In_1293);
nand U5624 (N_5624,In_2436,In_1600);
nor U5625 (N_5625,In_1839,In_1789);
nor U5626 (N_5626,In_2246,In_778);
or U5627 (N_5627,In_1322,In_1314);
nand U5628 (N_5628,In_289,In_2879);
nand U5629 (N_5629,In_1006,In_1143);
or U5630 (N_5630,In_734,In_450);
nor U5631 (N_5631,In_2364,In_1979);
nor U5632 (N_5632,In_2873,In_1075);
nor U5633 (N_5633,In_323,In_1725);
and U5634 (N_5634,In_1500,In_990);
and U5635 (N_5635,In_857,In_896);
or U5636 (N_5636,In_1037,In_2346);
and U5637 (N_5637,In_2530,In_109);
nand U5638 (N_5638,In_482,In_1134);
nand U5639 (N_5639,In_1494,In_980);
and U5640 (N_5640,In_1616,In_987);
or U5641 (N_5641,In_2491,In_2076);
xnor U5642 (N_5642,In_2036,In_869);
nand U5643 (N_5643,In_517,In_1190);
nand U5644 (N_5644,In_1957,In_1740);
xnor U5645 (N_5645,In_1044,In_2311);
nor U5646 (N_5646,In_58,In_1131);
xor U5647 (N_5647,In_1578,In_344);
and U5648 (N_5648,In_725,In_1892);
and U5649 (N_5649,In_2083,In_2758);
xnor U5650 (N_5650,In_2899,In_2532);
or U5651 (N_5651,In_261,In_92);
and U5652 (N_5652,In_680,In_831);
and U5653 (N_5653,In_2348,In_1344);
or U5654 (N_5654,In_2644,In_919);
or U5655 (N_5655,In_2057,In_1681);
nor U5656 (N_5656,In_210,In_2675);
nand U5657 (N_5657,In_101,In_2189);
and U5658 (N_5658,In_1943,In_2149);
nand U5659 (N_5659,In_766,In_1736);
and U5660 (N_5660,In_603,In_1855);
or U5661 (N_5661,In_1641,In_1341);
nand U5662 (N_5662,In_1562,In_1248);
xnor U5663 (N_5663,In_523,In_1996);
nand U5664 (N_5664,In_801,In_2849);
nor U5665 (N_5665,In_1518,In_249);
nor U5666 (N_5666,In_967,In_2349);
or U5667 (N_5667,In_2261,In_2793);
nand U5668 (N_5668,In_1641,In_2416);
xnor U5669 (N_5669,In_2975,In_2706);
nand U5670 (N_5670,In_618,In_528);
or U5671 (N_5671,In_1997,In_2820);
nor U5672 (N_5672,In_217,In_2140);
xnor U5673 (N_5673,In_1718,In_2980);
or U5674 (N_5674,In_1745,In_292);
or U5675 (N_5675,In_1274,In_1798);
nor U5676 (N_5676,In_519,In_125);
nand U5677 (N_5677,In_1162,In_263);
and U5678 (N_5678,In_558,In_553);
or U5679 (N_5679,In_2073,In_495);
nor U5680 (N_5680,In_2216,In_268);
nand U5681 (N_5681,In_1904,In_2617);
and U5682 (N_5682,In_715,In_2828);
nor U5683 (N_5683,In_601,In_676);
xnor U5684 (N_5684,In_65,In_2973);
nor U5685 (N_5685,In_493,In_1747);
and U5686 (N_5686,In_1409,In_1899);
and U5687 (N_5687,In_274,In_2414);
nand U5688 (N_5688,In_2387,In_2802);
nand U5689 (N_5689,In_996,In_666);
nand U5690 (N_5690,In_2331,In_810);
and U5691 (N_5691,In_80,In_445);
xnor U5692 (N_5692,In_686,In_2496);
nand U5693 (N_5693,In_2290,In_299);
nand U5694 (N_5694,In_2085,In_1486);
nor U5695 (N_5695,In_2233,In_2343);
or U5696 (N_5696,In_186,In_579);
nand U5697 (N_5697,In_2331,In_2172);
nor U5698 (N_5698,In_1848,In_2054);
and U5699 (N_5699,In_2345,In_20);
xor U5700 (N_5700,In_315,In_2613);
xnor U5701 (N_5701,In_2117,In_1654);
and U5702 (N_5702,In_1234,In_2055);
nand U5703 (N_5703,In_1422,In_2860);
nand U5704 (N_5704,In_1797,In_1589);
xor U5705 (N_5705,In_1625,In_1366);
or U5706 (N_5706,In_542,In_1882);
nand U5707 (N_5707,In_611,In_965);
nand U5708 (N_5708,In_2264,In_585);
nand U5709 (N_5709,In_1511,In_374);
or U5710 (N_5710,In_2921,In_828);
nand U5711 (N_5711,In_1333,In_124);
or U5712 (N_5712,In_1501,In_2663);
nand U5713 (N_5713,In_606,In_1333);
nor U5714 (N_5714,In_2926,In_352);
nor U5715 (N_5715,In_2256,In_1885);
nand U5716 (N_5716,In_1797,In_350);
and U5717 (N_5717,In_1137,In_563);
or U5718 (N_5718,In_422,In_1805);
or U5719 (N_5719,In_1876,In_2443);
and U5720 (N_5720,In_1623,In_1091);
nand U5721 (N_5721,In_2939,In_2708);
nor U5722 (N_5722,In_989,In_1828);
nor U5723 (N_5723,In_1039,In_1312);
and U5724 (N_5724,In_1895,In_903);
nand U5725 (N_5725,In_2246,In_494);
nand U5726 (N_5726,In_2578,In_2716);
nand U5727 (N_5727,In_531,In_1118);
nor U5728 (N_5728,In_2558,In_569);
nor U5729 (N_5729,In_1125,In_1641);
and U5730 (N_5730,In_869,In_643);
and U5731 (N_5731,In_2765,In_2882);
nor U5732 (N_5732,In_275,In_2363);
and U5733 (N_5733,In_1387,In_2827);
or U5734 (N_5734,In_1525,In_2383);
nor U5735 (N_5735,In_1416,In_1412);
and U5736 (N_5736,In_1360,In_2841);
nor U5737 (N_5737,In_903,In_582);
xnor U5738 (N_5738,In_1358,In_1676);
nand U5739 (N_5739,In_2107,In_164);
nor U5740 (N_5740,In_1553,In_1611);
and U5741 (N_5741,In_1968,In_2571);
and U5742 (N_5742,In_2701,In_141);
or U5743 (N_5743,In_2876,In_2455);
nand U5744 (N_5744,In_2384,In_2265);
or U5745 (N_5745,In_877,In_2905);
and U5746 (N_5746,In_502,In_562);
or U5747 (N_5747,In_1096,In_992);
nor U5748 (N_5748,In_809,In_926);
or U5749 (N_5749,In_1318,In_2110);
and U5750 (N_5750,In_1107,In_174);
and U5751 (N_5751,In_1456,In_2490);
and U5752 (N_5752,In_2636,In_1710);
and U5753 (N_5753,In_1985,In_2267);
and U5754 (N_5754,In_2734,In_2518);
or U5755 (N_5755,In_1623,In_12);
nor U5756 (N_5756,In_112,In_2580);
and U5757 (N_5757,In_2124,In_2239);
xnor U5758 (N_5758,In_687,In_2556);
or U5759 (N_5759,In_774,In_1407);
nand U5760 (N_5760,In_104,In_597);
nor U5761 (N_5761,In_29,In_1961);
xor U5762 (N_5762,In_1635,In_85);
nand U5763 (N_5763,In_2244,In_916);
xnor U5764 (N_5764,In_297,In_1247);
and U5765 (N_5765,In_731,In_2487);
nor U5766 (N_5766,In_2373,In_899);
nand U5767 (N_5767,In_417,In_2483);
nor U5768 (N_5768,In_544,In_1155);
and U5769 (N_5769,In_1673,In_1539);
nor U5770 (N_5770,In_1425,In_171);
nand U5771 (N_5771,In_902,In_284);
or U5772 (N_5772,In_1556,In_804);
nand U5773 (N_5773,In_2780,In_2018);
or U5774 (N_5774,In_1628,In_1547);
or U5775 (N_5775,In_1648,In_2051);
nand U5776 (N_5776,In_1955,In_760);
or U5777 (N_5777,In_2315,In_2059);
nand U5778 (N_5778,In_2332,In_1071);
nand U5779 (N_5779,In_2933,In_516);
or U5780 (N_5780,In_1881,In_490);
nand U5781 (N_5781,In_1828,In_2942);
nor U5782 (N_5782,In_862,In_860);
and U5783 (N_5783,In_2948,In_2962);
or U5784 (N_5784,In_2298,In_2105);
nor U5785 (N_5785,In_2557,In_2633);
nand U5786 (N_5786,In_2774,In_678);
and U5787 (N_5787,In_2992,In_906);
nand U5788 (N_5788,In_2939,In_162);
or U5789 (N_5789,In_2354,In_1742);
nand U5790 (N_5790,In_1080,In_2846);
or U5791 (N_5791,In_2959,In_2010);
nand U5792 (N_5792,In_1068,In_1372);
and U5793 (N_5793,In_1377,In_75);
nand U5794 (N_5794,In_1190,In_731);
xnor U5795 (N_5795,In_2842,In_1642);
xor U5796 (N_5796,In_2452,In_1668);
and U5797 (N_5797,In_303,In_1572);
and U5798 (N_5798,In_1566,In_992);
xor U5799 (N_5799,In_949,In_2791);
nand U5800 (N_5800,In_2812,In_2700);
nand U5801 (N_5801,In_212,In_2422);
nand U5802 (N_5802,In_2313,In_2945);
nor U5803 (N_5803,In_2880,In_2160);
nand U5804 (N_5804,In_1287,In_498);
nor U5805 (N_5805,In_461,In_1636);
or U5806 (N_5806,In_1267,In_2014);
nor U5807 (N_5807,In_1731,In_1187);
nor U5808 (N_5808,In_1244,In_1081);
or U5809 (N_5809,In_386,In_2730);
and U5810 (N_5810,In_479,In_2683);
and U5811 (N_5811,In_1551,In_1024);
or U5812 (N_5812,In_129,In_1814);
nand U5813 (N_5813,In_554,In_2551);
nor U5814 (N_5814,In_333,In_1362);
and U5815 (N_5815,In_1247,In_765);
and U5816 (N_5816,In_2683,In_2427);
or U5817 (N_5817,In_1590,In_1979);
nor U5818 (N_5818,In_682,In_390);
nand U5819 (N_5819,In_2508,In_1698);
nand U5820 (N_5820,In_2792,In_1146);
nor U5821 (N_5821,In_2106,In_2355);
nand U5822 (N_5822,In_2923,In_75);
nor U5823 (N_5823,In_928,In_1484);
and U5824 (N_5824,In_2115,In_1819);
nor U5825 (N_5825,In_209,In_2401);
nand U5826 (N_5826,In_2201,In_2678);
and U5827 (N_5827,In_1267,In_1210);
or U5828 (N_5828,In_2944,In_1471);
nand U5829 (N_5829,In_739,In_742);
nand U5830 (N_5830,In_835,In_1423);
nor U5831 (N_5831,In_8,In_1594);
nor U5832 (N_5832,In_2851,In_2543);
nor U5833 (N_5833,In_2241,In_1314);
nand U5834 (N_5834,In_1152,In_234);
xnor U5835 (N_5835,In_844,In_1337);
nand U5836 (N_5836,In_1484,In_132);
nor U5837 (N_5837,In_2346,In_1338);
and U5838 (N_5838,In_205,In_1963);
nor U5839 (N_5839,In_2510,In_2911);
nor U5840 (N_5840,In_2277,In_1201);
nand U5841 (N_5841,In_2754,In_2187);
xor U5842 (N_5842,In_601,In_834);
nor U5843 (N_5843,In_1569,In_545);
nand U5844 (N_5844,In_242,In_1703);
nor U5845 (N_5845,In_2053,In_1289);
or U5846 (N_5846,In_2107,In_1270);
nand U5847 (N_5847,In_1101,In_2086);
and U5848 (N_5848,In_1214,In_1936);
nand U5849 (N_5849,In_604,In_2304);
or U5850 (N_5850,In_2736,In_2017);
nand U5851 (N_5851,In_30,In_1884);
or U5852 (N_5852,In_1464,In_631);
and U5853 (N_5853,In_269,In_368);
nor U5854 (N_5854,In_103,In_1941);
xor U5855 (N_5855,In_595,In_1756);
and U5856 (N_5856,In_1795,In_754);
nor U5857 (N_5857,In_2686,In_2613);
or U5858 (N_5858,In_2503,In_137);
xnor U5859 (N_5859,In_2057,In_1457);
nand U5860 (N_5860,In_1181,In_207);
nor U5861 (N_5861,In_2525,In_114);
nand U5862 (N_5862,In_1298,In_1936);
and U5863 (N_5863,In_2762,In_2954);
nor U5864 (N_5864,In_2430,In_2348);
or U5865 (N_5865,In_2812,In_2366);
nand U5866 (N_5866,In_216,In_385);
or U5867 (N_5867,In_946,In_2449);
or U5868 (N_5868,In_2587,In_1120);
and U5869 (N_5869,In_318,In_400);
or U5870 (N_5870,In_727,In_273);
or U5871 (N_5871,In_1151,In_2104);
nor U5872 (N_5872,In_2280,In_959);
nor U5873 (N_5873,In_1298,In_900);
nor U5874 (N_5874,In_2586,In_657);
nor U5875 (N_5875,In_1114,In_1159);
nand U5876 (N_5876,In_109,In_1943);
or U5877 (N_5877,In_649,In_2425);
xnor U5878 (N_5878,In_793,In_2326);
nor U5879 (N_5879,In_2043,In_2818);
or U5880 (N_5880,In_1200,In_621);
nor U5881 (N_5881,In_1673,In_1706);
and U5882 (N_5882,In_311,In_1993);
or U5883 (N_5883,In_1612,In_799);
and U5884 (N_5884,In_2527,In_2935);
xnor U5885 (N_5885,In_2540,In_292);
and U5886 (N_5886,In_529,In_565);
nor U5887 (N_5887,In_1216,In_1765);
nor U5888 (N_5888,In_2227,In_2323);
xnor U5889 (N_5889,In_737,In_97);
xnor U5890 (N_5890,In_1630,In_609);
or U5891 (N_5891,In_2069,In_515);
or U5892 (N_5892,In_2390,In_2651);
nor U5893 (N_5893,In_1564,In_43);
nand U5894 (N_5894,In_570,In_1577);
nor U5895 (N_5895,In_2845,In_1068);
xnor U5896 (N_5896,In_1866,In_1787);
or U5897 (N_5897,In_1126,In_2301);
nor U5898 (N_5898,In_1306,In_1806);
nor U5899 (N_5899,In_1424,In_2085);
xnor U5900 (N_5900,In_128,In_1677);
nor U5901 (N_5901,In_1848,In_1402);
xnor U5902 (N_5902,In_1075,In_915);
and U5903 (N_5903,In_635,In_1707);
nand U5904 (N_5904,In_17,In_1945);
and U5905 (N_5905,In_2333,In_1447);
nand U5906 (N_5906,In_2865,In_652);
nand U5907 (N_5907,In_187,In_1634);
and U5908 (N_5908,In_2091,In_519);
or U5909 (N_5909,In_251,In_877);
nor U5910 (N_5910,In_2097,In_2007);
nand U5911 (N_5911,In_1498,In_2801);
and U5912 (N_5912,In_1868,In_2241);
nand U5913 (N_5913,In_2129,In_919);
or U5914 (N_5914,In_987,In_852);
nand U5915 (N_5915,In_2846,In_2869);
or U5916 (N_5916,In_598,In_1117);
nand U5917 (N_5917,In_2008,In_1471);
xor U5918 (N_5918,In_2919,In_2596);
nor U5919 (N_5919,In_1814,In_1141);
and U5920 (N_5920,In_2963,In_2278);
nand U5921 (N_5921,In_726,In_2388);
nand U5922 (N_5922,In_1870,In_2965);
nor U5923 (N_5923,In_613,In_395);
or U5924 (N_5924,In_864,In_2446);
nand U5925 (N_5925,In_2740,In_623);
and U5926 (N_5926,In_1496,In_357);
or U5927 (N_5927,In_771,In_464);
and U5928 (N_5928,In_2523,In_492);
nand U5929 (N_5929,In_1173,In_2440);
xnor U5930 (N_5930,In_210,In_2839);
nor U5931 (N_5931,In_1846,In_744);
nor U5932 (N_5932,In_1795,In_1188);
and U5933 (N_5933,In_945,In_1702);
or U5934 (N_5934,In_807,In_1547);
or U5935 (N_5935,In_2985,In_2230);
nor U5936 (N_5936,In_2246,In_936);
nor U5937 (N_5937,In_2770,In_967);
nand U5938 (N_5938,In_550,In_2938);
or U5939 (N_5939,In_1157,In_1260);
or U5940 (N_5940,In_869,In_2124);
nand U5941 (N_5941,In_2553,In_2124);
xor U5942 (N_5942,In_289,In_1374);
or U5943 (N_5943,In_1637,In_1301);
nor U5944 (N_5944,In_614,In_98);
nand U5945 (N_5945,In_1281,In_1038);
xor U5946 (N_5946,In_1350,In_1671);
nand U5947 (N_5947,In_2930,In_2843);
xor U5948 (N_5948,In_1626,In_1932);
nand U5949 (N_5949,In_844,In_2623);
or U5950 (N_5950,In_2339,In_1419);
nand U5951 (N_5951,In_84,In_1500);
nor U5952 (N_5952,In_1003,In_809);
nor U5953 (N_5953,In_1235,In_2532);
or U5954 (N_5954,In_1922,In_1594);
nor U5955 (N_5955,In_1715,In_901);
or U5956 (N_5956,In_61,In_1936);
or U5957 (N_5957,In_2545,In_1350);
and U5958 (N_5958,In_1245,In_2237);
and U5959 (N_5959,In_1434,In_2808);
nand U5960 (N_5960,In_2643,In_327);
and U5961 (N_5961,In_2926,In_470);
and U5962 (N_5962,In_1910,In_316);
or U5963 (N_5963,In_2207,In_1441);
nand U5964 (N_5964,In_752,In_295);
nor U5965 (N_5965,In_914,In_2988);
nand U5966 (N_5966,In_1169,In_2318);
nand U5967 (N_5967,In_2343,In_1500);
and U5968 (N_5968,In_1046,In_378);
and U5969 (N_5969,In_1017,In_2373);
and U5970 (N_5970,In_1098,In_1921);
nand U5971 (N_5971,In_635,In_565);
or U5972 (N_5972,In_194,In_2195);
and U5973 (N_5973,In_1449,In_2162);
nand U5974 (N_5974,In_1323,In_2259);
and U5975 (N_5975,In_3,In_1181);
or U5976 (N_5976,In_1324,In_2203);
nand U5977 (N_5977,In_2744,In_1706);
nor U5978 (N_5978,In_896,In_481);
and U5979 (N_5979,In_2426,In_2299);
and U5980 (N_5980,In_2606,In_744);
nor U5981 (N_5981,In_785,In_2195);
nand U5982 (N_5982,In_699,In_526);
and U5983 (N_5983,In_1101,In_1552);
and U5984 (N_5984,In_1127,In_732);
nor U5985 (N_5985,In_428,In_2232);
nor U5986 (N_5986,In_309,In_2261);
and U5987 (N_5987,In_1879,In_1248);
and U5988 (N_5988,In_1160,In_1580);
nor U5989 (N_5989,In_413,In_1181);
or U5990 (N_5990,In_2820,In_289);
nor U5991 (N_5991,In_2115,In_780);
and U5992 (N_5992,In_1374,In_1155);
and U5993 (N_5993,In_2394,In_819);
or U5994 (N_5994,In_2684,In_523);
or U5995 (N_5995,In_2960,In_1811);
or U5996 (N_5996,In_1908,In_1351);
nor U5997 (N_5997,In_1025,In_748);
nor U5998 (N_5998,In_1450,In_1429);
and U5999 (N_5999,In_1229,In_951);
nand U6000 (N_6000,N_797,N_578);
nor U6001 (N_6001,N_2859,N_2200);
nand U6002 (N_6002,N_1623,N_5041);
nand U6003 (N_6003,N_4682,N_5845);
nand U6004 (N_6004,N_5807,N_5259);
nor U6005 (N_6005,N_822,N_41);
or U6006 (N_6006,N_661,N_548);
nor U6007 (N_6007,N_4467,N_3929);
and U6008 (N_6008,N_3404,N_1497);
and U6009 (N_6009,N_2375,N_994);
or U6010 (N_6010,N_3633,N_4591);
xor U6011 (N_6011,N_537,N_4617);
nand U6012 (N_6012,N_4182,N_2794);
nand U6013 (N_6013,N_3989,N_188);
xnor U6014 (N_6014,N_5420,N_4075);
xor U6015 (N_6015,N_5040,N_1501);
nor U6016 (N_6016,N_4600,N_31);
and U6017 (N_6017,N_2997,N_5818);
and U6018 (N_6018,N_1710,N_2669);
nor U6019 (N_6019,N_5799,N_5646);
nand U6020 (N_6020,N_3525,N_2345);
and U6021 (N_6021,N_4933,N_5050);
nor U6022 (N_6022,N_1894,N_2426);
and U6023 (N_6023,N_5132,N_1771);
or U6024 (N_6024,N_4681,N_4662);
and U6025 (N_6025,N_3017,N_1945);
and U6026 (N_6026,N_3492,N_5944);
and U6027 (N_6027,N_4572,N_5523);
and U6028 (N_6028,N_3379,N_5430);
nand U6029 (N_6029,N_5087,N_4639);
nand U6030 (N_6030,N_5366,N_3490);
nand U6031 (N_6031,N_1616,N_1764);
nand U6032 (N_6032,N_1031,N_4926);
nand U6033 (N_6033,N_3669,N_605);
and U6034 (N_6034,N_3002,N_734);
nand U6035 (N_6035,N_1073,N_1293);
nand U6036 (N_6036,N_5679,N_3988);
nor U6037 (N_6037,N_51,N_3352);
xnor U6038 (N_6038,N_5276,N_3541);
nand U6039 (N_6039,N_3118,N_3408);
nor U6040 (N_6040,N_2240,N_4376);
nand U6041 (N_6041,N_4373,N_5334);
or U6042 (N_6042,N_1388,N_582);
or U6043 (N_6043,N_5978,N_2770);
or U6044 (N_6044,N_4430,N_3454);
and U6045 (N_6045,N_3417,N_5566);
nor U6046 (N_6046,N_556,N_4858);
nand U6047 (N_6047,N_695,N_5491);
and U6048 (N_6048,N_2142,N_2901);
nand U6049 (N_6049,N_550,N_2875);
nand U6050 (N_6050,N_1376,N_918);
and U6051 (N_6051,N_3188,N_5494);
or U6052 (N_6052,N_4936,N_1163);
xnor U6053 (N_6053,N_4200,N_3363);
nor U6054 (N_6054,N_1586,N_4406);
nor U6055 (N_6055,N_513,N_3259);
and U6056 (N_6056,N_2366,N_588);
or U6057 (N_6057,N_2391,N_5480);
nor U6058 (N_6058,N_4538,N_2125);
nand U6059 (N_6059,N_3519,N_323);
nand U6060 (N_6060,N_1199,N_1047);
nor U6061 (N_6061,N_1347,N_496);
nor U6062 (N_6062,N_5591,N_877);
and U6063 (N_6063,N_1495,N_4924);
or U6064 (N_6064,N_5587,N_563);
nor U6065 (N_6065,N_2439,N_5383);
xnor U6066 (N_6066,N_4768,N_1526);
and U6067 (N_6067,N_203,N_2441);
and U6068 (N_6068,N_1825,N_2981);
or U6069 (N_6069,N_5840,N_4152);
nand U6070 (N_6070,N_1723,N_1342);
nor U6071 (N_6071,N_2839,N_1652);
or U6072 (N_6072,N_5801,N_4257);
and U6073 (N_6073,N_1631,N_375);
or U6074 (N_6074,N_5335,N_1731);
nand U6075 (N_6075,N_4421,N_1570);
and U6076 (N_6076,N_5036,N_229);
nor U6077 (N_6077,N_5286,N_2098);
and U6078 (N_6078,N_5526,N_5316);
and U6079 (N_6079,N_5340,N_3652);
nor U6080 (N_6080,N_343,N_5529);
and U6081 (N_6081,N_3504,N_5950);
nand U6082 (N_6082,N_2648,N_5594);
nand U6083 (N_6083,N_2510,N_3673);
and U6084 (N_6084,N_4105,N_5022);
nor U6085 (N_6085,N_445,N_5290);
nand U6086 (N_6086,N_3770,N_2908);
and U6087 (N_6087,N_1533,N_2049);
nor U6088 (N_6088,N_1386,N_1837);
nor U6089 (N_6089,N_1310,N_220);
nand U6090 (N_6090,N_1970,N_596);
and U6091 (N_6091,N_4855,N_1254);
or U6092 (N_6092,N_1987,N_1428);
or U6093 (N_6093,N_5226,N_3640);
and U6094 (N_6094,N_4577,N_740);
nor U6095 (N_6095,N_3883,N_5681);
and U6096 (N_6096,N_3040,N_2363);
nor U6097 (N_6097,N_4811,N_3376);
or U6098 (N_6098,N_924,N_2507);
or U6099 (N_6099,N_2016,N_2842);
and U6100 (N_6100,N_2036,N_115);
or U6101 (N_6101,N_3748,N_3555);
or U6102 (N_6102,N_4663,N_1530);
and U6103 (N_6103,N_665,N_1795);
nand U6104 (N_6104,N_3416,N_795);
nand U6105 (N_6105,N_1080,N_1517);
or U6106 (N_6106,N_330,N_86);
nand U6107 (N_6107,N_4080,N_2879);
or U6108 (N_6108,N_4063,N_3201);
nand U6109 (N_6109,N_182,N_2050);
nor U6110 (N_6110,N_2547,N_2357);
and U6111 (N_6111,N_4747,N_2198);
or U6112 (N_6112,N_4206,N_1767);
nor U6113 (N_6113,N_1929,N_3372);
nand U6114 (N_6114,N_5304,N_3647);
and U6115 (N_6115,N_2671,N_5856);
nor U6116 (N_6116,N_5999,N_744);
nand U6117 (N_6117,N_42,N_2038);
and U6118 (N_6118,N_1176,N_4215);
nand U6119 (N_6119,N_836,N_448);
nor U6120 (N_6120,N_3406,N_2664);
nor U6121 (N_6121,N_5005,N_3998);
xor U6122 (N_6122,N_2867,N_3203);
and U6123 (N_6123,N_4575,N_5541);
xor U6124 (N_6124,N_1593,N_4966);
or U6125 (N_6125,N_1012,N_1704);
nand U6126 (N_6126,N_692,N_469);
or U6127 (N_6127,N_3461,N_1819);
nand U6128 (N_6128,N_3339,N_5583);
or U6129 (N_6129,N_3445,N_2673);
nand U6130 (N_6130,N_3191,N_2549);
nor U6131 (N_6131,N_2392,N_699);
xnor U6132 (N_6132,N_4311,N_2067);
or U6133 (N_6133,N_3233,N_1991);
xor U6134 (N_6134,N_1249,N_4438);
nand U6135 (N_6135,N_5149,N_5424);
xor U6136 (N_6136,N_5016,N_3288);
or U6137 (N_6137,N_5957,N_4930);
nand U6138 (N_6138,N_1452,N_319);
nor U6139 (N_6139,N_3333,N_3122);
and U6140 (N_6140,N_4998,N_3790);
nor U6141 (N_6141,N_219,N_1202);
nand U6142 (N_6142,N_3892,N_1128);
nand U6143 (N_6143,N_2451,N_4491);
nor U6144 (N_6144,N_5795,N_3522);
nand U6145 (N_6145,N_1626,N_4156);
xnor U6146 (N_6146,N_1367,N_5339);
xnor U6147 (N_6147,N_1658,N_3390);
nand U6148 (N_6148,N_4917,N_2741);
and U6149 (N_6149,N_128,N_1093);
nand U6150 (N_6150,N_1446,N_4274);
or U6151 (N_6151,N_93,N_3389);
nand U6152 (N_6152,N_5524,N_5625);
nor U6153 (N_6153,N_4873,N_2256);
nand U6154 (N_6154,N_4767,N_2204);
and U6155 (N_6155,N_2083,N_893);
nand U6156 (N_6156,N_3769,N_2935);
nand U6157 (N_6157,N_5805,N_1307);
nand U6158 (N_6158,N_5467,N_3733);
or U6159 (N_6159,N_2783,N_5387);
or U6160 (N_6160,N_4095,N_1886);
and U6161 (N_6161,N_5300,N_3211);
or U6162 (N_6162,N_4729,N_3049);
nand U6163 (N_6163,N_4451,N_304);
nand U6164 (N_6164,N_4932,N_4440);
nand U6165 (N_6165,N_5013,N_3126);
and U6166 (N_6166,N_1865,N_2045);
xor U6167 (N_6167,N_4359,N_5636);
nor U6168 (N_6168,N_3,N_865);
nor U6169 (N_6169,N_5251,N_3586);
nand U6170 (N_6170,N_2534,N_718);
nand U6171 (N_6171,N_5696,N_5633);
nor U6172 (N_6172,N_1655,N_2925);
nor U6173 (N_6173,N_447,N_1339);
or U6174 (N_6174,N_3195,N_2866);
nand U6175 (N_6175,N_3248,N_930);
nor U6176 (N_6176,N_2290,N_811);
and U6177 (N_6177,N_4089,N_4646);
xnor U6178 (N_6178,N_2405,N_3134);
and U6179 (N_6179,N_5662,N_1605);
xor U6180 (N_6180,N_5240,N_4615);
and U6181 (N_6181,N_5153,N_4425);
nand U6182 (N_6182,N_5769,N_5262);
xor U6183 (N_6183,N_3974,N_4412);
and U6184 (N_6184,N_3907,N_4341);
nor U6185 (N_6185,N_5266,N_4202);
nand U6186 (N_6186,N_4053,N_4893);
nand U6187 (N_6187,N_1360,N_4526);
nor U6188 (N_6188,N_2499,N_2550);
xnor U6189 (N_6189,N_2597,N_1089);
or U6190 (N_6190,N_4717,N_2927);
and U6191 (N_6191,N_4715,N_3571);
or U6192 (N_6192,N_1736,N_470);
nor U6193 (N_6193,N_2327,N_1488);
or U6194 (N_6194,N_2896,N_5894);
and U6195 (N_6195,N_5138,N_4846);
xor U6196 (N_6196,N_2931,N_4249);
nor U6197 (N_6197,N_4817,N_1131);
or U6198 (N_6198,N_952,N_3059);
nor U6199 (N_6199,N_2462,N_3047);
or U6200 (N_6200,N_406,N_3478);
nand U6201 (N_6201,N_4276,N_2591);
or U6202 (N_6202,N_4698,N_2789);
or U6203 (N_6203,N_1294,N_1644);
or U6204 (N_6204,N_5349,N_5927);
or U6205 (N_6205,N_2257,N_46);
nand U6206 (N_6206,N_449,N_3030);
or U6207 (N_6207,N_3976,N_5450);
and U6208 (N_6208,N_1839,N_3133);
nand U6209 (N_6209,N_3598,N_3582);
and U6210 (N_6210,N_2460,N_3308);
nor U6211 (N_6211,N_3192,N_23);
or U6212 (N_6212,N_807,N_1926);
or U6213 (N_6213,N_5298,N_4340);
and U6214 (N_6214,N_3833,N_1461);
nand U6215 (N_6215,N_3986,N_4083);
or U6216 (N_6216,N_4132,N_3480);
nand U6217 (N_6217,N_957,N_1086);
and U6218 (N_6218,N_5687,N_3128);
or U6219 (N_6219,N_3491,N_987);
and U6220 (N_6220,N_613,N_1684);
and U6221 (N_6221,N_5510,N_4568);
nor U6222 (N_6222,N_3275,N_5949);
nor U6223 (N_6223,N_4149,N_813);
nand U6224 (N_6224,N_326,N_2918);
xnor U6225 (N_6225,N_3013,N_202);
and U6226 (N_6226,N_5873,N_3531);
nor U6227 (N_6227,N_2580,N_5830);
or U6228 (N_6228,N_3577,N_2370);
and U6229 (N_6229,N_3025,N_878);
nand U6230 (N_6230,N_5284,N_1538);
nor U6231 (N_6231,N_5230,N_5060);
nand U6232 (N_6232,N_1755,N_2078);
and U6233 (N_6233,N_2403,N_1782);
or U6234 (N_6234,N_4522,N_3570);
or U6235 (N_6235,N_3696,N_30);
xnor U6236 (N_6236,N_4207,N_3872);
nor U6237 (N_6237,N_2563,N_114);
or U6238 (N_6238,N_4939,N_4432);
or U6239 (N_6239,N_761,N_4145);
nand U6240 (N_6240,N_2063,N_4454);
nor U6241 (N_6241,N_2118,N_3709);
nor U6242 (N_6242,N_1918,N_2685);
or U6243 (N_6243,N_3289,N_4822);
nand U6244 (N_6244,N_3991,N_2238);
xor U6245 (N_6245,N_5393,N_2620);
and U6246 (N_6246,N_1236,N_5425);
nor U6247 (N_6247,N_2593,N_1171);
nand U6248 (N_6248,N_5462,N_5075);
and U6249 (N_6249,N_566,N_4942);
nand U6250 (N_6250,N_494,N_5874);
and U6251 (N_6251,N_1705,N_3517);
and U6252 (N_6252,N_5175,N_1326);
and U6253 (N_6253,N_5731,N_3039);
nor U6254 (N_6254,N_712,N_532);
nand U6255 (N_6255,N_1017,N_526);
or U6256 (N_6256,N_2590,N_299);
and U6257 (N_6257,N_1726,N_887);
or U6258 (N_6258,N_4177,N_2860);
or U6259 (N_6259,N_2598,N_735);
nand U6260 (N_6260,N_941,N_1035);
nor U6261 (N_6261,N_4316,N_2724);
and U6262 (N_6262,N_4929,N_4306);
nand U6263 (N_6263,N_3380,N_5697);
nor U6264 (N_6264,N_4716,N_2231);
nand U6265 (N_6265,N_1550,N_1242);
nor U6266 (N_6266,N_5573,N_56);
and U6267 (N_6267,N_4755,N_4141);
and U6268 (N_6268,N_1132,N_1735);
or U6269 (N_6269,N_639,N_270);
nand U6270 (N_6270,N_2605,N_3237);
and U6271 (N_6271,N_1406,N_2400);
and U6272 (N_6272,N_5373,N_4040);
nor U6273 (N_6273,N_910,N_1474);
nor U6274 (N_6274,N_1272,N_272);
nand U6275 (N_6275,N_1481,N_3583);
and U6276 (N_6276,N_2746,N_454);
and U6277 (N_6277,N_5753,N_5444);
and U6278 (N_6278,N_3723,N_3905);
nand U6279 (N_6279,N_4898,N_2861);
or U6280 (N_6280,N_5260,N_2585);
nand U6281 (N_6281,N_458,N_4530);
nor U6282 (N_6282,N_4308,N_5505);
and U6283 (N_6283,N_4876,N_4632);
xnor U6284 (N_6284,N_105,N_2153);
or U6285 (N_6285,N_4070,N_2304);
or U6286 (N_6286,N_4258,N_2682);
or U6287 (N_6287,N_685,N_1935);
nand U6288 (N_6288,N_2989,N_4000);
nand U6289 (N_6289,N_5553,N_2934);
and U6290 (N_6290,N_2279,N_5980);
and U6291 (N_6291,N_4622,N_748);
nand U6292 (N_6292,N_4518,N_5421);
and U6293 (N_6293,N_5466,N_3698);
and U6294 (N_6294,N_4500,N_5747);
xor U6295 (N_6295,N_5324,N_2141);
or U6296 (N_6296,N_3928,N_87);
or U6297 (N_6297,N_2830,N_4244);
and U6298 (N_6298,N_5461,N_3407);
nand U6299 (N_6299,N_348,N_5991);
nand U6300 (N_6300,N_3184,N_4969);
xor U6301 (N_6301,N_5185,N_5144);
nor U6302 (N_6302,N_2571,N_2005);
nor U6303 (N_6303,N_1599,N_1983);
nand U6304 (N_6304,N_5415,N_881);
or U6305 (N_6305,N_2980,N_3801);
or U6306 (N_6306,N_3925,N_248);
and U6307 (N_6307,N_450,N_4041);
nor U6308 (N_6308,N_4205,N_2898);
or U6309 (N_6309,N_336,N_3557);
nor U6310 (N_6310,N_1629,N_269);
or U6311 (N_6311,N_4766,N_4475);
nor U6312 (N_6312,N_3452,N_3750);
and U6313 (N_6313,N_2071,N_5066);
or U6314 (N_6314,N_5200,N_2251);
and U6315 (N_6315,N_5618,N_1742);
nand U6316 (N_6316,N_5150,N_1756);
and U6317 (N_6317,N_4489,N_4543);
and U6318 (N_6318,N_3336,N_5055);
or U6319 (N_6319,N_2709,N_2288);
or U6320 (N_6320,N_391,N_3533);
or U6321 (N_6321,N_1919,N_5151);
or U6322 (N_6322,N_2225,N_5294);
and U6323 (N_6323,N_2275,N_2641);
or U6324 (N_6324,N_570,N_3662);
nand U6325 (N_6325,N_2386,N_2693);
nand U6326 (N_6326,N_4702,N_776);
or U6327 (N_6327,N_606,N_390);
and U6328 (N_6328,N_1632,N_1589);
nor U6329 (N_6329,N_1722,N_1947);
nor U6330 (N_6330,N_5832,N_2611);
nor U6331 (N_6331,N_497,N_4913);
nand U6332 (N_6332,N_2321,N_620);
nor U6333 (N_6333,N_1602,N_830);
nor U6334 (N_6334,N_5976,N_1953);
and U6335 (N_6335,N_5893,N_5813);
xor U6336 (N_6336,N_5416,N_5402);
and U6337 (N_6337,N_4051,N_4428);
nor U6338 (N_6338,N_4624,N_790);
nand U6339 (N_6339,N_2052,N_3057);
or U6340 (N_6340,N_542,N_5848);
or U6341 (N_6341,N_2721,N_1603);
and U6342 (N_6342,N_736,N_1915);
nor U6343 (N_6343,N_4955,N_2120);
or U6344 (N_6344,N_4305,N_5126);
and U6345 (N_6345,N_1387,N_898);
nand U6346 (N_6346,N_1170,N_412);
nor U6347 (N_6347,N_1287,N_1668);
nor U6348 (N_6348,N_5164,N_2466);
and U6349 (N_6349,N_5725,N_841);
nor U6350 (N_6350,N_4834,N_1963);
and U6351 (N_6351,N_867,N_1799);
and U6352 (N_6352,N_633,N_2668);
or U6353 (N_6353,N_3561,N_875);
or U6354 (N_6354,N_4787,N_2284);
xnor U6355 (N_6355,N_2947,N_2502);
nor U6356 (N_6356,N_2396,N_2469);
nor U6357 (N_6357,N_2185,N_4180);
or U6358 (N_6358,N_3546,N_1288);
or U6359 (N_6359,N_752,N_5855);
nor U6360 (N_6360,N_5490,N_561);
or U6361 (N_6361,N_5699,N_831);
or U6362 (N_6362,N_3756,N_3311);
nor U6363 (N_6363,N_5033,N_4928);
or U6364 (N_6364,N_3614,N_1322);
or U6365 (N_6365,N_2139,N_3123);
nor U6366 (N_6366,N_4970,N_3719);
nor U6367 (N_6367,N_1590,N_1037);
or U6368 (N_6368,N_5321,N_672);
nor U6369 (N_6369,N_3219,N_2862);
and U6370 (N_6370,N_522,N_2608);
or U6371 (N_6371,N_2224,N_16);
xor U6372 (N_6372,N_3368,N_482);
nor U6373 (N_6373,N_1627,N_3979);
and U6374 (N_6374,N_4107,N_492);
and U6375 (N_6375,N_5837,N_5802);
nand U6376 (N_6376,N_3834,N_4414);
or U6377 (N_6377,N_5015,N_3117);
nor U6378 (N_6378,N_2882,N_395);
nor U6379 (N_6379,N_1305,N_3479);
or U6380 (N_6380,N_5501,N_5977);
or U6381 (N_6381,N_3643,N_2915);
nor U6382 (N_6382,N_4488,N_2751);
nand U6383 (N_6383,N_2303,N_432);
or U6384 (N_6384,N_1761,N_2798);
and U6385 (N_6385,N_1715,N_5849);
nand U6386 (N_6386,N_1924,N_2412);
xnor U6387 (N_6387,N_4806,N_546);
or U6388 (N_6388,N_2184,N_4974);
and U6389 (N_6389,N_3388,N_1464);
nand U6390 (N_6390,N_451,N_5095);
and U6391 (N_6391,N_2261,N_5826);
or U6392 (N_6392,N_552,N_2891);
nor U6393 (N_6393,N_2034,N_1480);
or U6394 (N_6394,N_3249,N_1359);
or U6395 (N_6395,N_1773,N_1544);
nor U6396 (N_6396,N_5859,N_2979);
and U6397 (N_6397,N_3537,N_4794);
or U6398 (N_6398,N_4762,N_4757);
nor U6399 (N_6399,N_1707,N_3220);
and U6400 (N_6400,N_5273,N_747);
or U6401 (N_6401,N_4162,N_5863);
nand U6402 (N_6402,N_2335,N_280);
nand U6403 (N_6403,N_1453,N_5224);
xnor U6404 (N_6404,N_3244,N_1341);
xor U6405 (N_6405,N_758,N_1058);
nor U6406 (N_6406,N_3864,N_5852);
or U6407 (N_6407,N_3215,N_510);
and U6408 (N_6408,N_3212,N_3163);
and U6409 (N_6409,N_2632,N_4761);
nand U6410 (N_6410,N_947,N_4687);
or U6411 (N_6411,N_5209,N_1636);
nor U6412 (N_6412,N_1133,N_1628);
nand U6413 (N_6413,N_4976,N_3593);
nor U6414 (N_6414,N_1262,N_464);
or U6415 (N_6415,N_4706,N_3205);
nand U6416 (N_6416,N_1548,N_5632);
nand U6417 (N_6417,N_2320,N_2186);
or U6418 (N_6418,N_1139,N_4602);
and U6419 (N_6419,N_667,N_2110);
nand U6420 (N_6420,N_111,N_3657);
nand U6421 (N_6421,N_1233,N_3292);
and U6422 (N_6422,N_2066,N_3682);
or U6423 (N_6423,N_284,N_4732);
xor U6424 (N_6424,N_622,N_4736);
or U6425 (N_6425,N_4980,N_5248);
nor U6426 (N_6426,N_5857,N_2904);
and U6427 (N_6427,N_4288,N_3736);
nor U6428 (N_6428,N_1787,N_3966);
xor U6429 (N_6429,N_5436,N_213);
or U6430 (N_6430,N_5481,N_5596);
nor U6431 (N_6431,N_2094,N_4650);
nand U6432 (N_6432,N_3015,N_4704);
nor U6433 (N_6433,N_2670,N_4461);
and U6434 (N_6434,N_5154,N_4374);
nand U6435 (N_6435,N_5943,N_1247);
or U6436 (N_6436,N_4866,N_3022);
and U6437 (N_6437,N_3793,N_4754);
xnor U6438 (N_6438,N_4388,N_5888);
nand U6439 (N_6439,N_3313,N_5323);
or U6440 (N_6440,N_1664,N_1881);
and U6441 (N_6441,N_4569,N_4712);
xor U6442 (N_6442,N_3291,N_5942);
nand U6443 (N_6443,N_715,N_2802);
nor U6444 (N_6444,N_2222,N_3664);
nor U6445 (N_6445,N_3660,N_1984);
nand U6446 (N_6446,N_3939,N_1990);
nor U6447 (N_6447,N_17,N_5918);
and U6448 (N_6448,N_3584,N_315);
nand U6449 (N_6449,N_1346,N_7);
nand U6450 (N_6450,N_5563,N_4441);
nor U6451 (N_6451,N_245,N_3766);
and U6452 (N_6452,N_1621,N_1185);
and U6453 (N_6453,N_5287,N_1059);
nand U6454 (N_6454,N_936,N_1317);
nor U6455 (N_6455,N_5508,N_5655);
or U6456 (N_6456,N_1999,N_3937);
and U6457 (N_6457,N_69,N_5434);
nand U6458 (N_6458,N_1229,N_638);
or U6459 (N_6459,N_2277,N_356);
and U6460 (N_6460,N_1181,N_3306);
or U6461 (N_6461,N_1124,N_2265);
nand U6462 (N_6462,N_559,N_2458);
xor U6463 (N_6463,N_4369,N_2509);
or U6464 (N_6464,N_3323,N_5348);
nand U6465 (N_6465,N_5449,N_3509);
or U6466 (N_6466,N_4985,N_2992);
and U6467 (N_6467,N_5345,N_4036);
or U6468 (N_6468,N_1023,N_2607);
or U6469 (N_6469,N_886,N_3846);
nor U6470 (N_6470,N_5891,N_2413);
nor U6471 (N_6471,N_1808,N_2619);
or U6472 (N_6472,N_226,N_2354);
or U6473 (N_6473,N_2427,N_760);
nand U6474 (N_6474,N_2229,N_5228);
xor U6475 (N_6475,N_5790,N_3398);
nor U6476 (N_6476,N_3969,N_4212);
and U6477 (N_6477,N_4556,N_4077);
or U6478 (N_6478,N_3970,N_2630);
or U6479 (N_6479,N_2291,N_2171);
or U6480 (N_6480,N_5382,N_4192);
nand U6481 (N_6481,N_619,N_1175);
nor U6482 (N_6482,N_2324,N_1209);
and U6483 (N_6483,N_2621,N_4143);
and U6484 (N_6484,N_3109,N_2476);
nor U6485 (N_6485,N_864,N_3505);
xor U6486 (N_6486,N_2180,N_4870);
nand U6487 (N_6487,N_3838,N_960);
and U6488 (N_6488,N_3495,N_907);
nand U6489 (N_6489,N_1729,N_2022);
nor U6490 (N_6490,N_1425,N_895);
and U6491 (N_6491,N_1671,N_707);
and U6492 (N_6492,N_2459,N_325);
or U6493 (N_6493,N_5191,N_4015);
nor U6494 (N_6494,N_3520,N_525);
nor U6495 (N_6495,N_119,N_4171);
nand U6496 (N_6496,N_1643,N_3646);
and U6497 (N_6497,N_473,N_5301);
nor U6498 (N_6498,N_2592,N_1724);
and U6499 (N_6499,N_1980,N_1496);
and U6500 (N_6500,N_34,N_3107);
and U6501 (N_6501,N_855,N_5320);
and U6502 (N_6502,N_5322,N_3863);
and U6503 (N_6503,N_2811,N_1955);
nor U6504 (N_6504,N_4493,N_5307);
nand U6505 (N_6505,N_5838,N_5280);
nand U6506 (N_6506,N_5463,N_1315);
and U6507 (N_6507,N_4387,N_2076);
or U6508 (N_6508,N_1469,N_5559);
nand U6509 (N_6509,N_3337,N_4719);
and U6510 (N_6510,N_4914,N_300);
nand U6511 (N_6511,N_3786,N_5333);
nor U6512 (N_6512,N_279,N_2361);
nand U6513 (N_6513,N_3011,N_3960);
and U6514 (N_6514,N_3052,N_902);
and U6515 (N_6515,N_5247,N_2216);
or U6516 (N_6516,N_757,N_2126);
or U6517 (N_6517,N_9,N_650);
nand U6518 (N_6518,N_2624,N_5923);
and U6519 (N_6519,N_600,N_5546);
or U6520 (N_6520,N_5053,N_2813);
nand U6521 (N_6521,N_2021,N_1845);
nor U6522 (N_6522,N_558,N_4273);
and U6523 (N_6523,N_2878,N_3512);
and U6524 (N_6524,N_4385,N_5118);
and U6525 (N_6525,N_1774,N_2649);
nor U6526 (N_6526,N_401,N_5285);
nor U6527 (N_6527,N_4660,N_3508);
or U6528 (N_6528,N_2637,N_845);
and U6529 (N_6529,N_2040,N_2828);
or U6530 (N_6530,N_901,N_1149);
xor U6531 (N_6531,N_55,N_1228);
and U6532 (N_6532,N_4750,N_1781);
and U6533 (N_6533,N_549,N_5303);
nand U6534 (N_6534,N_5825,N_749);
nor U6535 (N_6535,N_1213,N_1261);
nor U6536 (N_6536,N_5428,N_2834);
or U6537 (N_6537,N_2892,N_1524);
or U6538 (N_6538,N_44,N_3060);
and U6539 (N_6539,N_1665,N_4919);
nor U6540 (N_6540,N_3327,N_5647);
or U6541 (N_6541,N_2310,N_2388);
or U6542 (N_6542,N_428,N_5581);
xnor U6543 (N_6543,N_4034,N_5884);
or U6544 (N_6544,N_1607,N_1519);
or U6545 (N_6545,N_4726,N_2161);
nor U6546 (N_6546,N_1145,N_2779);
and U6547 (N_6547,N_5751,N_5935);
nand U6548 (N_6548,N_2764,N_4620);
or U6549 (N_6549,N_5374,N_4799);
or U6550 (N_6550,N_1079,N_4973);
or U6551 (N_6551,N_4098,N_5770);
or U6552 (N_6552,N_5445,N_5232);
nor U6553 (N_6553,N_3361,N_3744);
or U6554 (N_6554,N_2395,N_5565);
xor U6555 (N_6555,N_2656,N_2951);
xor U6556 (N_6556,N_2958,N_4112);
nor U6557 (N_6557,N_2876,N_1415);
and U6558 (N_6558,N_4424,N_3050);
xnor U6559 (N_6559,N_5292,N_67);
or U6560 (N_6560,N_3365,N_5879);
nand U6561 (N_6561,N_3995,N_5610);
nor U6562 (N_6562,N_140,N_2870);
and U6563 (N_6563,N_3626,N_2823);
xor U6564 (N_6564,N_4847,N_1297);
or U6565 (N_6565,N_4635,N_5584);
nand U6566 (N_6566,N_1884,N_1741);
and U6567 (N_6567,N_1189,N_92);
nor U6568 (N_6568,N_5722,N_4218);
and U6569 (N_6569,N_4471,N_4150);
nand U6570 (N_6570,N_676,N_3155);
nor U6571 (N_6571,N_1558,N_4029);
or U6572 (N_6572,N_409,N_113);
and U6573 (N_6573,N_2368,N_2533);
nor U6574 (N_6574,N_4032,N_4618);
or U6575 (N_6575,N_2129,N_1269);
or U6576 (N_6576,N_5034,N_531);
nor U6577 (N_6577,N_5869,N_3279);
or U6578 (N_6578,N_2385,N_2695);
or U6579 (N_6579,N_274,N_4355);
nand U6580 (N_6580,N_3874,N_3559);
nand U6581 (N_6581,N_3261,N_1115);
or U6582 (N_6582,N_4850,N_4158);
nand U6583 (N_6583,N_3532,N_205);
nor U6584 (N_6584,N_5982,N_419);
nand U6585 (N_6585,N_3899,N_4184);
or U6586 (N_6586,N_4469,N_355);
nand U6587 (N_6587,N_2893,N_3886);
and U6588 (N_6588,N_1908,N_3482);
xnor U6589 (N_6589,N_172,N_859);
or U6590 (N_6590,N_5672,N_2138);
nor U6591 (N_6591,N_4444,N_809);
or U6592 (N_6592,N_4364,N_95);
nor U6593 (N_6593,N_2750,N_4948);
or U6594 (N_6594,N_5086,N_4514);
nand U6595 (N_6595,N_3674,N_5734);
and U6596 (N_6596,N_3785,N_788);
or U6597 (N_6597,N_1559,N_2775);
nor U6598 (N_6598,N_815,N_1780);
and U6599 (N_6599,N_350,N_2192);
nand U6600 (N_6600,N_335,N_1419);
and U6601 (N_6601,N_3572,N_81);
and U6602 (N_6602,N_2188,N_14);
and U6603 (N_6603,N_3827,N_3415);
and U6604 (N_6604,N_168,N_5692);
and U6605 (N_6605,N_2610,N_5651);
or U6606 (N_6606,N_5535,N_671);
or U6607 (N_6607,N_3513,N_5302);
nor U6608 (N_6608,N_4110,N_623);
xor U6609 (N_6609,N_152,N_365);
nor U6610 (N_6610,N_4951,N_1728);
nand U6611 (N_6611,N_3999,N_3705);
and U6612 (N_6612,N_2097,N_5203);
and U6613 (N_6613,N_5970,N_1564);
and U6614 (N_6614,N_1725,N_2259);
xor U6615 (N_6615,N_2372,N_2864);
nor U6616 (N_6616,N_4140,N_688);
and U6617 (N_6617,N_2230,N_4419);
or U6618 (N_6618,N_4278,N_5527);
and U6619 (N_6619,N_493,N_3198);
or U6620 (N_6620,N_3320,N_4291);
and U6621 (N_6621,N_5483,N_1477);
or U6622 (N_6622,N_1087,N_360);
or U6623 (N_6623,N_1932,N_177);
xor U6624 (N_6624,N_2272,N_3617);
xor U6625 (N_6625,N_3083,N_2752);
or U6626 (N_6626,N_1662,N_3239);
and U6627 (N_6627,N_5435,N_914);
and U6628 (N_6628,N_3878,N_2220);
nor U6629 (N_6629,N_2053,N_985);
xnor U6630 (N_6630,N_3762,N_2011);
nor U6631 (N_6631,N_5782,N_5243);
and U6632 (N_6632,N_799,N_4565);
or U6633 (N_6633,N_677,N_1043);
or U6634 (N_6634,N_3282,N_631);
nand U6635 (N_6635,N_427,N_1216);
or U6636 (N_6636,N_2821,N_5028);
nand U6637 (N_6637,N_1878,N_4803);
and U6638 (N_6638,N_3018,N_1549);
nor U6639 (N_6639,N_1299,N_5069);
and U6640 (N_6640,N_4246,N_3189);
or U6641 (N_6641,N_3689,N_2705);
nand U6642 (N_6642,N_1577,N_3916);
xnor U6643 (N_6643,N_5715,N_1323);
and U6644 (N_6644,N_1235,N_2243);
nand U6645 (N_6645,N_819,N_2936);
nor U6646 (N_6646,N_1498,N_2850);
nor U6647 (N_6647,N_2900,N_2984);
or U6648 (N_6648,N_3355,N_3611);
nor U6649 (N_6649,N_1896,N_5966);
or U6650 (N_6650,N_2603,N_5989);
xnor U6651 (N_6651,N_1336,N_3395);
nor U6652 (N_6652,N_1484,N_3277);
xnor U6653 (N_6653,N_1557,N_175);
nand U6654 (N_6654,N_2493,N_2048);
and U6655 (N_6655,N_5534,N_2541);
nor U6656 (N_6656,N_5457,N_4299);
nand U6657 (N_6657,N_5834,N_1536);
nand U6658 (N_6658,N_5992,N_3920);
or U6659 (N_6659,N_3114,N_2480);
nor U6660 (N_6660,N_2877,N_2636);
or U6661 (N_6661,N_2924,N_256);
xnor U6662 (N_6662,N_938,N_2218);
nor U6663 (N_6663,N_2848,N_1904);
or U6664 (N_6664,N_820,N_3104);
or U6665 (N_6665,N_738,N_3470);
xor U6666 (N_6666,N_3314,N_2851);
nand U6667 (N_6667,N_517,N_1523);
nand U6668 (N_6668,N_4473,N_4154);
or U6669 (N_6669,N_2456,N_1195);
xnor U6670 (N_6670,N_2911,N_1745);
xnor U6671 (N_6671,N_850,N_3160);
or U6672 (N_6672,N_3247,N_1231);
and U6673 (N_6673,N_4453,N_2377);
and U6674 (N_6674,N_3803,N_3199);
nor U6675 (N_6675,N_3156,N_911);
nor U6676 (N_6676,N_2626,N_5084);
or U6677 (N_6677,N_5575,N_4413);
nand U6678 (N_6678,N_709,N_0);
xor U6679 (N_6679,N_5114,N_1022);
or U6680 (N_6680,N_2683,N_3934);
nor U6681 (N_6681,N_842,N_4781);
and U6682 (N_6682,N_5960,N_303);
and U6683 (N_6683,N_2857,N_4882);
or U6684 (N_6684,N_5338,N_4512);
nor U6685 (N_6685,N_644,N_2568);
or U6686 (N_6686,N_3858,N_103);
nand U6687 (N_6687,N_680,N_2638);
or U6688 (N_6688,N_431,N_2351);
and U6689 (N_6689,N_988,N_4818);
nand U6690 (N_6690,N_2573,N_3540);
or U6691 (N_6691,N_5227,N_837);
nor U6692 (N_6692,N_2614,N_5652);
or U6693 (N_6693,N_5735,N_2824);
and U6694 (N_6694,N_3168,N_870);
nand U6695 (N_6695,N_5570,N_1610);
and U6696 (N_6696,N_1330,N_1950);
and U6697 (N_6697,N_5048,N_1936);
nor U6698 (N_6698,N_2564,N_1522);
nand U6699 (N_6699,N_5475,N_3831);
nor U6700 (N_6700,N_2754,N_2807);
nor U6701 (N_6701,N_1817,N_3453);
and U6702 (N_6702,N_424,N_1210);
or U6703 (N_6703,N_4656,N_1978);
xnor U6704 (N_6704,N_1830,N_4668);
nor U6705 (N_6705,N_4742,N_3464);
or U6706 (N_6706,N_3550,N_4231);
or U6707 (N_6707,N_1925,N_5308);
nand U6708 (N_6708,N_4446,N_4232);
or U6709 (N_6709,N_530,N_1098);
nand U6710 (N_6710,N_5775,N_885);
nand U6711 (N_6711,N_3940,N_5979);
or U6712 (N_6712,N_3130,N_3216);
nand U6713 (N_6713,N_5554,N_5160);
nor U6714 (N_6714,N_4261,N_2755);
xnor U6715 (N_6715,N_1815,N_3909);
and U6716 (N_6716,N_3366,N_5641);
and U6717 (N_6717,N_4820,N_2657);
xnor U6718 (N_6718,N_1828,N_5907);
nand U6719 (N_6719,N_5101,N_2690);
xor U6720 (N_6720,N_2030,N_2943);
and U6721 (N_6721,N_239,N_2863);
nand U6722 (N_6722,N_5352,N_4476);
or U6723 (N_6723,N_2089,N_5104);
and U6724 (N_6724,N_1591,N_5601);
xnor U6725 (N_6725,N_4398,N_4555);
or U6726 (N_6726,N_2162,N_1848);
nand U6727 (N_6727,N_4330,N_4988);
or U6728 (N_6728,N_341,N_555);
nand U6729 (N_6729,N_2954,N_651);
nand U6730 (N_6730,N_3171,N_196);
nor U6731 (N_6731,N_3426,N_3845);
xor U6732 (N_6732,N_3321,N_1889);
or U6733 (N_6733,N_1001,N_4760);
nand U6734 (N_6734,N_3627,N_169);
nor U6735 (N_6735,N_4020,N_800);
or U6736 (N_6736,N_2601,N_1020);
nand U6737 (N_6737,N_2430,N_5119);
nand U6738 (N_6738,N_2276,N_689);
or U6739 (N_6739,N_3399,N_277);
or U6740 (N_6740,N_2181,N_3996);
xnor U6741 (N_6741,N_380,N_1416);
or U6742 (N_6742,N_3258,N_5314);
nor U6743 (N_6743,N_288,N_3356);
or U6744 (N_6744,N_3042,N_1958);
nand U6745 (N_6745,N_3903,N_1097);
xor U6746 (N_6746,N_3534,N_4049);
and U6747 (N_6747,N_1617,N_3401);
or U6748 (N_6748,N_3433,N_2604);
nor U6749 (N_6749,N_4745,N_2930);
nand U6750 (N_6750,N_2301,N_1650);
and U6751 (N_6751,N_3746,N_216);
nand U6752 (N_6752,N_4133,N_5497);
or U6753 (N_6753,N_1314,N_4164);
and U6754 (N_6754,N_2114,N_5630);
xor U6755 (N_6755,N_3706,N_2562);
nand U6756 (N_6756,N_349,N_1806);
nand U6757 (N_6757,N_71,N_832);
and U6758 (N_6758,N_4483,N_4956);
nor U6759 (N_6759,N_2064,N_455);
xnor U6760 (N_6760,N_5555,N_3590);
nor U6761 (N_6761,N_1747,N_5781);
and U6762 (N_6762,N_583,N_3494);
nand U6763 (N_6763,N_306,N_4744);
nor U6764 (N_6764,N_4515,N_1788);
and U6765 (N_6765,N_3307,N_945);
or U6766 (N_6766,N_2616,N_358);
or U6767 (N_6767,N_5403,N_3094);
or U6768 (N_6768,N_1528,N_4418);
and U6769 (N_6769,N_110,N_834);
nor U6770 (N_6770,N_1700,N_2596);
nor U6771 (N_6771,N_3560,N_1850);
and U6772 (N_6772,N_5768,N_4612);
nand U6773 (N_6773,N_2497,N_313);
nand U6774 (N_6774,N_5702,N_4225);
or U6775 (N_6775,N_1504,N_1666);
nor U6776 (N_6776,N_3129,N_1686);
nor U6777 (N_6777,N_2727,N_3100);
and U6778 (N_6778,N_408,N_4400);
nand U6779 (N_6779,N_4775,N_4361);
nand U6780 (N_6780,N_2163,N_388);
nand U6781 (N_6781,N_4124,N_1499);
or U6782 (N_6782,N_1466,N_2437);
nor U6783 (N_6783,N_4353,N_3449);
nand U6784 (N_6784,N_4375,N_3080);
nand U6785 (N_6785,N_3090,N_5720);
nand U6786 (N_6786,N_38,N_2843);
and U6787 (N_6787,N_208,N_2704);
or U6788 (N_6788,N_3392,N_1823);
nand U6789 (N_6789,N_528,N_3102);
or U6790 (N_6790,N_3477,N_149);
xor U6791 (N_6791,N_3562,N_3502);
or U6792 (N_6792,N_3469,N_351);
or U6793 (N_6793,N_2529,N_4081);
nor U6794 (N_6794,N_3856,N_53);
nor U6795 (N_6795,N_533,N_3581);
and U6796 (N_6796,N_4864,N_4125);
or U6797 (N_6797,N_146,N_2806);
or U6798 (N_6798,N_3567,N_4513);
or U6799 (N_6799,N_2482,N_3255);
nor U6800 (N_6800,N_1997,N_5707);
and U6801 (N_6801,N_5597,N_4896);
nor U6802 (N_6802,N_240,N_5311);
or U6803 (N_6803,N_2618,N_3424);
nor U6804 (N_6804,N_2663,N_1361);
or U6805 (N_6805,N_4025,N_4384);
or U6806 (N_6806,N_1214,N_4269);
nand U6807 (N_6807,N_1188,N_711);
xnor U6808 (N_6808,N_4393,N_562);
nor U6809 (N_6809,N_3257,N_3843);
nand U6810 (N_6810,N_3947,N_3839);
nand U6811 (N_6811,N_5344,N_503);
or U6812 (N_6812,N_1816,N_4601);
or U6813 (N_6813,N_2341,N_777);
xor U6814 (N_6814,N_965,N_5117);
and U6815 (N_6815,N_871,N_995);
nor U6816 (N_6816,N_3463,N_892);
nor U6817 (N_6817,N_3993,N_2105);
nand U6818 (N_6818,N_5532,N_529);
or U6819 (N_6819,N_1455,N_295);
nor U6820 (N_6820,N_5068,N_4693);
nor U6821 (N_6821,N_1612,N_2854);
nor U6822 (N_6822,N_2825,N_2101);
nand U6823 (N_6823,N_2814,N_2401);
and U6824 (N_6824,N_385,N_456);
nor U6825 (N_6825,N_4027,N_2945);
or U6826 (N_6826,N_2974,N_2205);
or U6827 (N_6827,N_5381,N_414);
nand U6828 (N_6828,N_384,N_3644);
xor U6829 (N_6829,N_4343,N_5924);
and U6830 (N_6830,N_362,N_1454);
xor U6831 (N_6831,N_4753,N_5789);
xor U6832 (N_6832,N_2332,N_1021);
nand U6833 (N_6833,N_2500,N_154);
or U6834 (N_6834,N_5614,N_1754);
and U6835 (N_6835,N_211,N_768);
or U6836 (N_6836,N_2719,N_2890);
xor U6837 (N_6837,N_5111,N_4644);
and U6838 (N_6838,N_5097,N_163);
nand U6839 (N_6839,N_2278,N_3943);
or U6840 (N_6840,N_40,N_33);
or U6841 (N_6841,N_1338,N_5188);
nor U6842 (N_6842,N_5872,N_5961);
nor U6843 (N_6843,N_2556,N_4735);
or U6844 (N_6844,N_2577,N_4405);
nand U6845 (N_6845,N_2211,N_377);
nor U6846 (N_6846,N_3904,N_2913);
nor U6847 (N_6847,N_2058,N_5724);
nand U6848 (N_6848,N_4860,N_5020);
xnor U6849 (N_6849,N_716,N_3527);
xnor U6850 (N_6850,N_478,N_4155);
and U6851 (N_6851,N_2521,N_5275);
and U6852 (N_6852,N_2699,N_5002);
and U6853 (N_6853,N_1951,N_4763);
nand U6854 (N_6854,N_4194,N_3295);
nand U6855 (N_6855,N_4123,N_1717);
or U6856 (N_6856,N_4074,N_624);
nand U6857 (N_6857,N_3891,N_29);
or U6858 (N_6858,N_2506,N_1398);
or U6859 (N_6859,N_2991,N_4902);
and U6860 (N_6860,N_2096,N_3262);
nand U6861 (N_6861,N_4751,N_969);
nor U6862 (N_6862,N_4292,N_135);
or U6863 (N_6863,N_5673,N_2152);
nor U6864 (N_6864,N_900,N_4664);
and U6865 (N_6865,N_3737,N_3132);
nor U6866 (N_6866,N_805,N_4114);
nor U6867 (N_6867,N_4727,N_2492);
nand U6868 (N_6868,N_499,N_1027);
or U6869 (N_6869,N_5103,N_2144);
xor U6870 (N_6870,N_4911,N_4665);
xor U6871 (N_6871,N_5184,N_773);
and U6872 (N_6872,N_1653,N_4429);
and U6873 (N_6873,N_3860,N_4907);
nand U6874 (N_6874,N_5492,N_1220);
nor U6875 (N_6875,N_1660,N_4496);
or U6876 (N_6876,N_2902,N_4067);
nand U6877 (N_6877,N_1719,N_1067);
nand U6878 (N_6878,N_5774,N_5426);
nand U6879 (N_6879,N_955,N_4759);
or U6880 (N_6880,N_45,N_889);
or U6881 (N_6881,N_3910,N_4637);
nor U6882 (N_6882,N_2213,N_4268);
and U6883 (N_6883,N_501,N_339);
nor U6884 (N_6884,N_5824,N_2044);
or U6885 (N_6885,N_5983,N_2517);
nor U6886 (N_6886,N_849,N_5410);
nor U6887 (N_6887,N_5777,N_4528);
nand U6888 (N_6888,N_1385,N_4694);
and U6889 (N_6889,N_3972,N_1797);
or U6890 (N_6890,N_4950,N_5507);
nor U6891 (N_6891,N_59,N_1566);
or U6892 (N_6892,N_2369,N_1578);
nor U6893 (N_6893,N_1794,N_5897);
xnor U6894 (N_6894,N_5379,N_5684);
and U6895 (N_6895,N_4718,N_252);
nand U6896 (N_6896,N_1870,N_1205);
or U6897 (N_6897,N_803,N_2306);
xnor U6898 (N_6898,N_5589,N_2099);
nor U6899 (N_6899,N_1648,N_5540);
or U6900 (N_6900,N_4654,N_4509);
nor U6901 (N_6901,N_1121,N_2552);
and U6902 (N_6902,N_4519,N_1692);
and U6903 (N_6903,N_5582,N_982);
or U6904 (N_6904,N_2317,N_439);
or U6905 (N_6905,N_1165,N_5956);
and U6906 (N_6906,N_1887,N_1108);
nor U6907 (N_6907,N_5617,N_5009);
nand U6908 (N_6908,N_5560,N_4151);
xnor U6909 (N_6909,N_3773,N_5000);
nor U6910 (N_6910,N_3936,N_872);
and U6911 (N_6911,N_13,N_2095);
nand U6912 (N_6912,N_2708,N_3190);
and U6913 (N_6913,N_2849,N_2343);
or U6914 (N_6914,N_5800,N_3641);
nand U6915 (N_6915,N_1669,N_5422);
nor U6916 (N_6916,N_433,N_268);
and U6917 (N_6917,N_2987,N_4078);
nand U6918 (N_6918,N_3553,N_998);
or U6919 (N_6919,N_2025,N_770);
nand U6920 (N_6920,N_4671,N_5237);
and U6921 (N_6921,N_5914,N_3120);
and U6922 (N_6922,N_5268,N_2068);
nor U6923 (N_6923,N_4462,N_3420);
and U6924 (N_6924,N_4506,N_1107);
or U6925 (N_6925,N_2778,N_4284);
nand U6926 (N_6926,N_944,N_4999);
nor U6927 (N_6927,N_4836,N_5796);
nand U6928 (N_6928,N_4166,N_5128);
and U6929 (N_6929,N_3254,N_2772);
xnor U6930 (N_6930,N_1274,N_2287);
or U6931 (N_6931,N_926,N_4138);
and U6932 (N_6932,N_5190,N_1917);
nor U6933 (N_6933,N_4723,N_5252);
xor U6934 (N_6934,N_1066,N_3384);
nor U6935 (N_6935,N_5804,N_4022);
and U6936 (N_6936,N_3428,N_3791);
nor U6937 (N_6937,N_2241,N_899);
nand U6938 (N_6938,N_230,N_964);
or U6939 (N_6939,N_3418,N_3784);
and U6940 (N_6940,N_1417,N_1995);
and U6941 (N_6941,N_2575,N_5089);
xor U6942 (N_6942,N_5356,N_193);
and U6943 (N_6943,N_2446,N_4172);
xor U6944 (N_6944,N_255,N_1289);
xnor U6945 (N_6945,N_3543,N_1620);
and U6946 (N_6946,N_3442,N_5061);
nor U6947 (N_6947,N_18,N_5210);
or U6948 (N_6948,N_3318,N_764);
or U6949 (N_6949,N_3604,N_2143);
and U6950 (N_6950,N_1706,N_4833);
nand U6951 (N_6951,N_4339,N_3077);
nand U6952 (N_6952,N_1458,N_4399);
nor U6953 (N_6953,N_1721,N_2841);
or U6954 (N_6954,N_2838,N_4352);
and U6955 (N_6955,N_1948,N_5667);
and U6956 (N_6956,N_3659,N_4944);
and U6957 (N_6957,N_3183,N_5578);
nand U6958 (N_6958,N_5690,N_5574);
nand U6959 (N_6959,N_3594,N_802);
and U6960 (N_6960,N_3981,N_5744);
or U6961 (N_6961,N_950,N_5370);
nor U6962 (N_6962,N_975,N_4527);
nor U6963 (N_6963,N_3004,N_4146);
or U6964 (N_6964,N_3064,N_4821);
nor U6965 (N_6965,N_5336,N_2907);
or U6966 (N_6966,N_3739,N_915);
nand U6967 (N_6967,N_170,N_4434);
or U6968 (N_6968,N_3780,N_4128);
and U6969 (N_6969,N_4659,N_144);
and U6970 (N_6970,N_5847,N_5386);
and U6971 (N_6971,N_5905,N_5442);
and U6972 (N_6972,N_3754,N_4317);
nor U6973 (N_6973,N_3564,N_5313);
and U6974 (N_6974,N_4195,N_2572);
or U6975 (N_6975,N_5728,N_438);
nand U6976 (N_6976,N_4465,N_5661);
or U6977 (N_6977,N_3334,N_5605);
or U6978 (N_6978,N_5109,N_1587);
or U6979 (N_6979,N_1117,N_4566);
and U6980 (N_6980,N_5295,N_2639);
nand U6981 (N_6981,N_1718,N_1321);
nand U6982 (N_6982,N_756,N_1749);
nor U6983 (N_6983,N_1711,N_4903);
or U6984 (N_6984,N_4802,N_1252);
xnor U6985 (N_6985,N_4275,N_64);
nand U6986 (N_6986,N_96,N_713);
nor U6987 (N_6987,N_771,N_4925);
nor U6988 (N_6988,N_3115,N_4266);
and U6989 (N_6989,N_244,N_282);
and U6990 (N_6990,N_714,N_2054);
nand U6991 (N_6991,N_4370,N_590);
nand U6992 (N_6992,N_3458,N_4962);
or U6993 (N_6993,N_2504,N_4119);
and U6994 (N_6994,N_3524,N_4532);
and U6995 (N_6995,N_4720,N_5207);
or U6996 (N_6996,N_2075,N_5900);
nor U6997 (N_6997,N_4542,N_5972);
nand U6998 (N_6998,N_466,N_467);
nand U6999 (N_6999,N_2817,N_2157);
xor U7000 (N_7000,N_4627,N_5470);
or U7001 (N_7001,N_4658,N_167);
and U7002 (N_7002,N_5443,N_5951);
and U7003 (N_7003,N_567,N_1155);
nor U7004 (N_7004,N_371,N_74);
xor U7005 (N_7005,N_407,N_4529);
and U7006 (N_7006,N_1281,N_1637);
nand U7007 (N_7007,N_4807,N_4511);
nor U7008 (N_7008,N_787,N_4841);
nor U7009 (N_7009,N_4014,N_5482);
nor U7010 (N_7010,N_1152,N_260);
nand U7011 (N_7011,N_5689,N_3642);
nor U7012 (N_7012,N_3747,N_1467);
and U7013 (N_7013,N_3093,N_3542);
and U7014 (N_7014,N_2475,N_422);
and U7015 (N_7015,N_3810,N_3783);
nor U7016 (N_7016,N_3310,N_4472);
nand U7017 (N_7017,N_241,N_2961);
xnor U7018 (N_7018,N_2519,N_2923);
nor U7019 (N_7019,N_129,N_2666);
or U7020 (N_7020,N_3949,N_3862);
nor U7021 (N_7021,N_1099,N_4810);
and U7022 (N_7022,N_5081,N_2262);
xor U7023 (N_7023,N_39,N_2199);
or U7024 (N_7024,N_1245,N_861);
xor U7025 (N_7025,N_5439,N_5572);
nand U7026 (N_7026,N_1260,N_3743);
nand U7027 (N_7027,N_4892,N_1801);
or U7028 (N_7028,N_1443,N_3854);
nand U7029 (N_7029,N_5793,N_2037);
and U7030 (N_7030,N_5199,N_4243);
nor U7031 (N_7031,N_2674,N_1026);
and U7032 (N_7032,N_5599,N_5831);
and U7033 (N_7033,N_1449,N_3214);
nand U7034 (N_7034,N_27,N_1019);
or U7035 (N_7035,N_696,N_703);
xnor U7036 (N_7036,N_1681,N_3752);
and U7037 (N_7037,N_242,N_3732);
nor U7038 (N_7038,N_1308,N_4691);
or U7039 (N_7039,N_374,N_3613);
or U7040 (N_7040,N_3054,N_979);
xor U7041 (N_7041,N_4436,N_4307);
and U7042 (N_7042,N_5530,N_1275);
nand U7043 (N_7043,N_3419,N_989);
nor U7044 (N_7044,N_1611,N_5562);
or U7045 (N_7045,N_4563,N_762);
and U7046 (N_7046,N_2855,N_4788);
and U7047 (N_7047,N_3136,N_5472);
nor U7048 (N_7048,N_264,N_5265);
nand U7049 (N_7049,N_686,N_251);
nand U7050 (N_7050,N_3599,N_271);
and U7051 (N_7051,N_3097,N_2004);
nor U7052 (N_7052,N_1010,N_3632);
nor U7053 (N_7053,N_5254,N_3888);
or U7054 (N_7054,N_243,N_2132);
and U7055 (N_7055,N_2508,N_5712);
nand U7056 (N_7056,N_4394,N_5908);
nand U7057 (N_7057,N_186,N_908);
or U7058 (N_7058,N_3089,N_28);
and U7059 (N_7059,N_430,N_3978);
nand U7060 (N_7060,N_3683,N_5045);
nor U7061 (N_7061,N_3354,N_4252);
nor U7062 (N_7062,N_5821,N_1270);
and U7063 (N_7063,N_483,N_2921);
nor U7064 (N_7064,N_5544,N_922);
nand U7065 (N_7065,N_4746,N_3252);
nand U7066 (N_7066,N_4501,N_3713);
nand U7067 (N_7067,N_127,N_2172);
and U7068 (N_7068,N_164,N_2374);
nor U7069 (N_7069,N_2996,N_2769);
and U7070 (N_7070,N_511,N_5108);
or U7071 (N_7071,N_3950,N_4830);
nand U7072 (N_7072,N_3885,N_2454);
nor U7073 (N_7073,N_1542,N_1651);
and U7074 (N_7074,N_1224,N_2090);
nor U7075 (N_7075,N_2108,N_4816);
nor U7076 (N_7076,N_162,N_4439);
xor U7077 (N_7077,N_3088,N_5078);
xor U7078 (N_7078,N_4101,N_212);
nand U7079 (N_7079,N_4069,N_2014);
nand U7080 (N_7080,N_5052,N_6);
nand U7081 (N_7081,N_5904,N_1873);
and U7082 (N_7082,N_2461,N_2886);
nor U7083 (N_7083,N_393,N_1834);
xnor U7084 (N_7084,N_1829,N_276);
xor U7085 (N_7085,N_191,N_8);
and U7086 (N_7086,N_2352,N_1541);
nor U7087 (N_7087,N_1957,N_453);
nor U7088 (N_7088,N_1070,N_3068);
xnor U7089 (N_7089,N_3804,N_2111);
nand U7090 (N_7090,N_4785,N_823);
and U7091 (N_7091,N_321,N_1221);
or U7092 (N_7092,N_1268,N_3069);
and U7093 (N_7093,N_3772,N_3958);
xor U7094 (N_7094,N_925,N_2874);
nand U7095 (N_7095,N_1772,N_3959);
nand U7096 (N_7096,N_1778,N_5543);
and U7097 (N_7097,N_357,N_98);
and U7098 (N_7098,N_1364,N_2026);
nor U7099 (N_7099,N_2191,N_4437);
or U7100 (N_7100,N_5091,N_920);
and U7101 (N_7101,N_5035,N_1048);
nor U7102 (N_7102,N_2350,N_2318);
nand U7103 (N_7103,N_781,N_3848);
and U7104 (N_7104,N_4641,N_1191);
or U7105 (N_7105,N_5072,N_967);
and U7106 (N_7106,N_1110,N_2905);
and U7107 (N_7107,N_857,N_3953);
and U7108 (N_7108,N_1861,N_3085);
or U7109 (N_7109,N_1583,N_4738);
or U7110 (N_7110,N_5718,N_5644);
nand U7111 (N_7111,N_5385,N_3394);
nand U7112 (N_7112,N_2540,N_192);
nand U7113 (N_7113,N_3151,N_4277);
nand U7114 (N_7114,N_5244,N_3340);
nor U7115 (N_7115,N_1956,N_2367);
nand U7116 (N_7116,N_2425,N_5354);
and U7117 (N_7117,N_1426,N_3667);
and U7118 (N_7118,N_5658,N_2822);
and U7119 (N_7119,N_2136,N_3521);
nor U7120 (N_7120,N_3460,N_3253);
or U7121 (N_7121,N_4259,N_2757);
nor U7122 (N_7122,N_5453,N_704);
or U7123 (N_7123,N_1877,N_5743);
and U7124 (N_7124,N_1327,N_5169);
nor U7125 (N_7125,N_4910,N_4570);
nand U7126 (N_7126,N_223,N_1403);
xnor U7127 (N_7127,N_2156,N_3410);
and U7128 (N_7128,N_3154,N_3402);
and U7129 (N_7129,N_2498,N_1401);
nand U7130 (N_7130,N_3493,N_1479);
or U7131 (N_7131,N_5620,N_3434);
nand U7132 (N_7132,N_3797,N_3137);
and U7133 (N_7133,N_3894,N_1846);
nor U7134 (N_7134,N_2576,N_1197);
nand U7135 (N_7135,N_2561,N_2043);
nand U7136 (N_7136,N_3703,N_5936);
or U7137 (N_7137,N_545,N_1374);
nand U7138 (N_7138,N_4852,N_1300);
nand U7139 (N_7139,N_2414,N_5930);
or U7140 (N_7140,N_5922,N_4332);
or U7141 (N_7141,N_2716,N_4201);
nor U7142 (N_7142,N_1639,N_1363);
nand U7143 (N_7143,N_5217,N_5129);
or U7144 (N_7144,N_5854,N_1263);
nand U7145 (N_7145,N_4581,N_5342);
or U7146 (N_7146,N_3853,N_1377);
and U7147 (N_7147,N_2336,N_1259);
and U7148 (N_7148,N_3507,N_3471);
and U7149 (N_7149,N_626,N_5858);
nor U7150 (N_7150,N_292,N_602);
xor U7151 (N_7151,N_933,N_2226);
nand U7152 (N_7152,N_4079,N_5738);
nand U7153 (N_7153,N_1414,N_4169);
nor U7154 (N_7154,N_3427,N_1109);
xor U7155 (N_7155,N_3921,N_153);
nand U7156 (N_7156,N_194,N_1039);
and U7157 (N_7157,N_19,N_3961);
nor U7158 (N_7158,N_3300,N_5080);
and U7159 (N_7159,N_1770,N_553);
and U7160 (N_7160,N_4228,N_4521);
nand U7161 (N_7161,N_519,N_3964);
or U7162 (N_7162,N_1814,N_4862);
nand U7163 (N_7163,N_3725,N_1015);
or U7164 (N_7164,N_3051,N_1378);
nor U7165 (N_7165,N_91,N_1531);
nor U7166 (N_7166,N_3496,N_4984);
nand U7167 (N_7167,N_4586,N_2124);
and U7168 (N_7168,N_3923,N_2645);
xor U7169 (N_7169,N_4590,N_2387);
and U7170 (N_7170,N_509,N_2298);
and U7171 (N_7171,N_4844,N_1333);
xnor U7172 (N_7172,N_798,N_4118);
and U7173 (N_7173,N_1193,N_2675);
or U7174 (N_7174,N_3957,N_4675);
nor U7175 (N_7175,N_2155,N_4296);
nor U7176 (N_7176,N_5264,N_4122);
or U7177 (N_7177,N_1,N_5783);
nand U7178 (N_7178,N_2474,N_4008);
or U7179 (N_7179,N_731,N_5642);
nand U7180 (N_7180,N_5341,N_5042);
and U7181 (N_7181,N_421,N_1399);
nand U7182 (N_7182,N_974,N_4731);
or U7183 (N_7183,N_5668,N_3185);
nand U7184 (N_7184,N_3649,N_3113);
and U7185 (N_7185,N_235,N_3962);
or U7186 (N_7186,N_2617,N_4889);
and U7187 (N_7187,N_1291,N_301);
and U7188 (N_7188,N_1485,N_3963);
nand U7189 (N_7189,N_4829,N_2232);
and U7190 (N_7190,N_2625,N_2844);
or U7191 (N_7191,N_3071,N_2409);
nor U7192 (N_7192,N_2164,N_4245);
xor U7193 (N_7193,N_2788,N_5616);
nor U7194 (N_7194,N_5551,N_1324);
or U7195 (N_7195,N_2732,N_3378);
or U7196 (N_7196,N_209,N_5746);
and U7197 (N_7197,N_1920,N_3835);
and U7198 (N_7198,N_396,N_664);
and U7199 (N_7199,N_2922,N_3242);
nand U7200 (N_7200,N_4853,N_5065);
nand U7201 (N_7201,N_953,N_2416);
nor U7202 (N_7202,N_1407,N_2883);
xnor U7203 (N_7203,N_2187,N_3634);
and U7204 (N_7204,N_3143,N_3767);
or U7205 (N_7205,N_5958,N_2219);
nand U7206 (N_7206,N_4573,N_2445);
nand U7207 (N_7207,N_2895,N_3707);
nand U7208 (N_7208,N_2121,N_4211);
and U7209 (N_7209,N_2473,N_1104);
nor U7210 (N_7210,N_2555,N_3987);
nand U7211 (N_7211,N_2281,N_4549);
xnor U7212 (N_7212,N_333,N_3152);
xnor U7213 (N_7213,N_1624,N_3879);
and U7214 (N_7214,N_4173,N_1311);
and U7215 (N_7215,N_5012,N_3021);
nand U7216 (N_7216,N_4442,N_2856);
nand U7217 (N_7217,N_2978,N_1529);
or U7218 (N_7218,N_5198,N_4545);
and U7219 (N_7219,N_2937,N_4728);
nor U7220 (N_7220,N_3729,N_2995);
and U7221 (N_7221,N_1052,N_1081);
nor U7222 (N_7222,N_3035,N_4724);
nand U7223 (N_7223,N_5788,N_5902);
nor U7224 (N_7224,N_5648,N_890);
nor U7225 (N_7225,N_4740,N_12);
or U7226 (N_7226,N_4048,N_4603);
nor U7227 (N_7227,N_3578,N_309);
or U7228 (N_7228,N_576,N_4979);
or U7229 (N_7229,N_5170,N_5705);
and U7230 (N_7230,N_2800,N_2681);
xnor U7231 (N_7231,N_5851,N_5389);
nand U7232 (N_7232,N_5148,N_2920);
nand U7233 (N_7233,N_5468,N_1304);
or U7234 (N_7234,N_2744,N_2560);
nand U7235 (N_7235,N_94,N_565);
or U7236 (N_7236,N_5974,N_5656);
nand U7237 (N_7237,N_3941,N_5853);
or U7238 (N_7238,N_5182,N_3202);
and U7239 (N_7239,N_1156,N_706);
nand U7240 (N_7240,N_263,N_1352);
nand U7241 (N_7241,N_2296,N_1740);
nand U7242 (N_7242,N_968,N_3997);
xnor U7243 (N_7243,N_3377,N_50);
xnor U7244 (N_7244,N_293,N_2820);
and U7245 (N_7245,N_1635,N_3605);
nand U7246 (N_7246,N_5634,N_3251);
nor U7247 (N_7247,N_1283,N_5073);
nand U7248 (N_7248,N_3514,N_5708);
and U7249 (N_7249,N_2260,N_4992);
nand U7250 (N_7250,N_4176,N_4780);
or U7251 (N_7251,N_3672,N_846);
nor U7252 (N_7252,N_5283,N_5351);
nand U7253 (N_7253,N_2970,N_4989);
nand U7254 (N_7254,N_2150,N_992);
or U7255 (N_7255,N_3761,N_3396);
xor U7256 (N_7256,N_1146,N_2364);
or U7257 (N_7257,N_4697,N_4946);
nand U7258 (N_7258,N_1137,N_3096);
nor U7259 (N_7259,N_4504,N_2165);
and U7260 (N_7260,N_1885,N_5455);
nand U7261 (N_7261,N_3547,N_2131);
nand U7262 (N_7262,N_2210,N_3164);
nand U7263 (N_7263,N_4019,N_3842);
nor U7264 (N_7264,N_4126,N_4606);
nand U7265 (N_7265,N_2189,N_3441);
and U7266 (N_7266,N_2847,N_1222);
nor U7267 (N_7267,N_5919,N_2178);
or U7268 (N_7268,N_5815,N_2270);
nor U7269 (N_7269,N_4289,N_595);
nand U7270 (N_7270,N_1371,N_5400);
or U7271 (N_7271,N_1095,N_397);
nor U7272 (N_7272,N_2274,N_3087);
xor U7273 (N_7273,N_2376,N_4062);
and U7274 (N_7274,N_3119,N_5984);
xnor U7275 (N_7275,N_4854,N_4782);
nor U7276 (N_7276,N_1656,N_5056);
or U7277 (N_7277,N_5357,N_4010);
nand U7278 (N_7278,N_1677,N_1543);
or U7279 (N_7279,N_662,N_515);
or U7280 (N_7280,N_3023,N_3938);
or U7281 (N_7281,N_5558,N_5369);
nor U7282 (N_7282,N_2609,N_3348);
nor U7283 (N_7283,N_1579,N_535);
or U7284 (N_7284,N_472,N_2333);
or U7285 (N_7285,N_2348,N_2223);
nor U7286 (N_7286,N_1227,N_1638);
nor U7287 (N_7287,N_327,N_2986);
or U7288 (N_7288,N_1113,N_990);
nand U7289 (N_7289,N_1854,N_457);
and U7290 (N_7290,N_4574,N_5538);
nand U7291 (N_7291,N_1094,N_4337);
nand U7292 (N_7292,N_769,N_126);
or U7293 (N_7293,N_5135,N_3722);
or U7294 (N_7294,N_3236,N_1906);
or U7295 (N_7295,N_4262,N_2023);
and U7296 (N_7296,N_4487,N_3715);
and U7297 (N_7297,N_946,N_4065);
or U7298 (N_7298,N_560,N_3326);
or U7299 (N_7299,N_4085,N_3029);
or U7300 (N_7300,N_5607,N_5660);
nand U7301 (N_7301,N_2382,N_2623);
nor U7302 (N_7302,N_3075,N_1096);
xnor U7303 (N_7303,N_4342,N_1910);
nor U7304 (N_7304,N_1064,N_364);
or U7305 (N_7305,N_5216,N_3545);
nor U7306 (N_7306,N_3230,N_5939);
or U7307 (N_7307,N_1051,N_4960);
and U7308 (N_7308,N_1641,N_2481);
nor U7309 (N_7309,N_2006,N_5528);
and U7310 (N_7310,N_827,N_3070);
and U7311 (N_7311,N_2526,N_1046);
nand U7312 (N_7312,N_125,N_3447);
or U7313 (N_7313,N_2906,N_418);
xor U7314 (N_7314,N_5604,N_2267);
nor U7315 (N_7315,N_4804,N_3086);
nor U7316 (N_7316,N_863,N_3924);
and U7317 (N_7317,N_3385,N_4016);
or U7318 (N_7318,N_4377,N_4251);
or U7319 (N_7319,N_923,N_564);
nand U7320 (N_7320,N_1647,N_3591);
nor U7321 (N_7321,N_3932,N_5046);
xor U7322 (N_7322,N_3965,N_1649);
nand U7323 (N_7323,N_2133,N_403);
xnor U7324 (N_7324,N_508,N_1595);
and U7325 (N_7325,N_5367,N_2444);
or U7326 (N_7326,N_1490,N_5967);
or U7327 (N_7327,N_4607,N_3286);
nand U7328 (N_7328,N_2994,N_5099);
and U7329 (N_7329,N_4204,N_4420);
nand U7330 (N_7330,N_3774,N_2092);
or U7331 (N_7331,N_3721,N_4510);
and U7332 (N_7332,N_3821,N_879);
and U7333 (N_7333,N_5044,N_97);
nor U7334 (N_7334,N_3685,N_4097);
nand U7335 (N_7335,N_5864,N_2438);
nor U7336 (N_7336,N_1243,N_3072);
and U7337 (N_7337,N_416,N_1029);
and U7338 (N_7338,N_4033,N_5399);
or U7339 (N_7339,N_4879,N_3009);
nand U7340 (N_7340,N_1092,N_2538);
nand U7341 (N_7341,N_5568,N_2762);
or U7342 (N_7342,N_1439,N_60);
or U7343 (N_7343,N_3587,N_1030);
xnor U7344 (N_7344,N_3990,N_1836);
nand U7345 (N_7345,N_1518,N_5533);
and U7346 (N_7346,N_4734,N_507);
or U7347 (N_7347,N_5197,N_5628);
and U7348 (N_7348,N_4046,N_4092);
and U7349 (N_7349,N_3444,N_1302);
nand U7350 (N_7350,N_5306,N_15);
xnor U7351 (N_7351,N_4843,N_4401);
nor U7352 (N_7352,N_3898,N_3283);
nand U7353 (N_7353,N_5571,N_5677);
nor U7354 (N_7354,N_5158,N_2201);
nand U7355 (N_7355,N_1056,N_1005);
nand U7356 (N_7356,N_5639,N_1619);
nand U7357 (N_7357,N_4497,N_3374);
or U7358 (N_7358,N_3697,N_2292);
nor U7359 (N_7359,N_4459,N_5585);
xor U7360 (N_7360,N_5401,N_4240);
nand U7361 (N_7361,N_2973,N_4028);
nor U7362 (N_7362,N_2872,N_5229);
and U7363 (N_7363,N_2447,N_3329);
or U7364 (N_7364,N_4611,N_1508);
xor U7365 (N_7365,N_5116,N_928);
or U7366 (N_7366,N_1429,N_1685);
or U7367 (N_7367,N_1279,N_1996);
xor U7368 (N_7368,N_3148,N_4579);
or U7369 (N_7369,N_2881,N_2565);
or U7370 (N_7370,N_4174,N_634);
or U7371 (N_7371,N_1285,N_866);
nand U7372 (N_7372,N_1698,N_4378);
nand U7373 (N_7373,N_2214,N_5809);
nand U7374 (N_7374,N_2109,N_3179);
nor U7375 (N_7375,N_1255,N_1525);
or U7376 (N_7376,N_2271,N_2212);
nor U7377 (N_7377,N_5931,N_4900);
nand U7378 (N_7378,N_3280,N_3276);
xnor U7379 (N_7379,N_3173,N_5365);
and U7380 (N_7380,N_479,N_68);
nor U7381 (N_7381,N_543,N_1369);
and U7382 (N_7382,N_2464,N_5518);
nor U7383 (N_7383,N_3579,N_3062);
or U7384 (N_7384,N_2147,N_5567);
and U7385 (N_7385,N_2467,N_2263);
nand U7386 (N_7386,N_801,N_4170);
or U7387 (N_7387,N_2939,N_3443);
xnor U7388 (N_7388,N_2631,N_2587);
or U7389 (N_7389,N_2252,N_32);
nor U7390 (N_7390,N_940,N_5844);
or U7391 (N_7391,N_5018,N_1927);
nand U7392 (N_7392,N_3802,N_4815);
nand U7393 (N_7393,N_796,N_682);
xnor U7394 (N_7394,N_1246,N_2266);
nand U7395 (N_7395,N_2865,N_1412);
nor U7396 (N_7396,N_4039,N_1792);
nor U7397 (N_7397,N_5142,N_882);
nor U7398 (N_7398,N_1103,N_4769);
and U7399 (N_7399,N_116,N_2799);
nor U7400 (N_7400,N_2999,N_3243);
nor U7401 (N_7401,N_257,N_1512);
and U7402 (N_7402,N_4448,N_3226);
nor U7403 (N_7403,N_3663,N_5007);
nor U7404 (N_7404,N_2146,N_2039);
nor U7405 (N_7405,N_1601,N_4707);
or U7406 (N_7406,N_917,N_4776);
nor U7407 (N_7407,N_1286,N_1858);
nand U7408 (N_7408,N_5638,N_1125);
nor U7409 (N_7409,N_2766,N_4825);
nor U7410 (N_7410,N_1120,N_3933);
or U7411 (N_7411,N_1042,N_5417);
nor U7412 (N_7412,N_137,N_1489);
and U7413 (N_7413,N_1786,N_4422);
nor U7414 (N_7414,N_725,N_1460);
and U7415 (N_7415,N_539,N_3944);
nor U7416 (N_7416,N_3437,N_1041);
nand U7417 (N_7417,N_2602,N_4877);
nor U7418 (N_7418,N_5868,N_3548);
nand U7419 (N_7419,N_904,N_5773);
nand U7420 (N_7420,N_4621,N_592);
or U7421 (N_7421,N_2104,N_4703);
and U7422 (N_7422,N_83,N_4625);
xor U7423 (N_7423,N_2300,N_4626);
or U7424 (N_7424,N_117,N_72);
xor U7425 (N_7425,N_5926,N_1897);
nand U7426 (N_7426,N_5159,N_463);
or U7427 (N_7427,N_10,N_1690);
xnor U7428 (N_7428,N_1940,N_4883);
nand U7429 (N_7429,N_3225,N_184);
xor U7430 (N_7430,N_2106,N_1232);
nor U7431 (N_7431,N_4905,N_2853);
nor U7432 (N_7432,N_76,N_698);
and U7433 (N_7433,N_3840,N_3956);
nand U7434 (N_7434,N_35,N_5742);
nor U7435 (N_7435,N_2432,N_1083);
and U7436 (N_7436,N_4562,N_4443);
nand U7437 (N_7437,N_4772,N_5234);
xor U7438 (N_7438,N_963,N_21);
nor U7439 (N_7439,N_4520,N_5934);
and U7440 (N_7440,N_308,N_4279);
nand U7441 (N_7441,N_4188,N_2805);
nand U7442 (N_7442,N_3044,N_3485);
nand U7443 (N_7443,N_1798,N_883);
nand U7444 (N_7444,N_1157,N_3628);
nor U7445 (N_7445,N_5098,N_1129);
or U7446 (N_7446,N_4131,N_1588);
or U7447 (N_7447,N_426,N_1922);
nand U7448 (N_7448,N_5709,N_2868);
nand U7449 (N_7449,N_954,N_224);
nand U7450 (N_7450,N_5877,N_314);
nand U7451 (N_7451,N_3297,N_4994);
nand U7452 (N_7452,N_225,N_5635);
nand U7453 (N_7453,N_2888,N_3193);
and U7454 (N_7454,N_4957,N_5219);
or U7455 (N_7455,N_547,N_5833);
or U7456 (N_7456,N_3565,N_3176);
nor U7457 (N_7457,N_1383,N_5969);
xor U7458 (N_7458,N_1992,N_5688);
and U7459 (N_7459,N_5238,N_1891);
xnor U7460 (N_7460,N_4031,N_2019);
nand U7461 (N_7461,N_2326,N_5947);
nor U7462 (N_7462,N_2491,N_1921);
or U7463 (N_7463,N_1573,N_959);
nor U7464 (N_7464,N_4923,N_381);
or U7465 (N_7465,N_724,N_1391);
or U7466 (N_7466,N_2389,N_1796);
and U7467 (N_7467,N_3603,N_5817);
xnor U7468 (N_7468,N_1765,N_4312);
nor U7469 (N_7469,N_774,N_387);
nor U7470 (N_7470,N_4379,N_3877);
nand U7471 (N_7471,N_1392,N_5107);
or U7472 (N_7472,N_2919,N_5090);
nand U7473 (N_7473,N_4552,N_5772);
nor U7474 (N_7474,N_5603,N_1200);
and U7475 (N_7475,N_4619,N_3635);
nor U7476 (N_7476,N_5112,N_5172);
and U7477 (N_7477,N_3116,N_792);
xnor U7478 (N_7478,N_1832,N_5194);
nor U7479 (N_7479,N_5319,N_635);
and U7480 (N_7480,N_5171,N_338);
nor U7481 (N_7481,N_2010,N_1841);
nand U7482 (N_7482,N_2559,N_5816);
nand U7483 (N_7483,N_2100,N_5432);
nand U7484 (N_7484,N_2170,N_2644);
or U7485 (N_7485,N_1971,N_5876);
nor U7486 (N_7486,N_5350,N_4498);
or U7487 (N_7487,N_3615,N_1257);
nand U7488 (N_7488,N_2686,N_1142);
or U7489 (N_7489,N_2969,N_5183);
nor U7490 (N_7490,N_3665,N_4390);
xor U7491 (N_7491,N_5423,N_5014);
or U7492 (N_7492,N_862,N_2522);
nor U7493 (N_7493,N_4784,N_1077);
and U7494 (N_7494,N_4314,N_3716);
or U7495 (N_7495,N_1944,N_22);
nor U7496 (N_7496,N_3296,N_5727);
nor U7497 (N_7497,N_206,N_2554);
nor U7498 (N_7498,N_465,N_3081);
nor U7499 (N_7499,N_259,N_3631);
and U7500 (N_7500,N_70,N_4190);
and U7501 (N_7501,N_4953,N_4001);
nor U7502 (N_7502,N_2293,N_1790);
nor U7503 (N_7503,N_4921,N_359);
nand U7504 (N_7504,N_5411,N_2889);
nor U7505 (N_7505,N_3166,N_812);
or U7506 (N_7506,N_3450,N_3229);
nand U7507 (N_7507,N_5364,N_4456);
or U7508 (N_7508,N_1818,N_2938);
and U7509 (N_7509,N_180,N_5839);
and U7510 (N_7510,N_2653,N_5819);
and U7511 (N_7511,N_2314,N_1733);
nand U7512 (N_7512,N_231,N_3830);
or U7513 (N_7513,N_2676,N_3001);
nand U7514 (N_7514,N_147,N_3552);
nor U7515 (N_7515,N_5177,N_506);
and U7516 (N_7516,N_1126,N_4544);
or U7517 (N_7517,N_5975,N_4294);
or U7518 (N_7518,N_1344,N_498);
nand U7519 (N_7519,N_462,N_4918);
nand U7520 (N_7520,N_2313,N_1592);
or U7521 (N_7521,N_5096,N_2127);
or U7522 (N_7522,N_1143,N_3638);
or U7523 (N_7523,N_5459,N_5139);
nand U7524 (N_7524,N_5010,N_367);
or U7525 (N_7525,N_5315,N_5397);
or U7526 (N_7526,N_4977,N_3636);
or U7527 (N_7527,N_1276,N_3816);
nor U7528 (N_7528,N_1154,N_2135);
or U7529 (N_7529,N_1618,N_3610);
and U7530 (N_7530,N_5161,N_1208);
or U7531 (N_7531,N_973,N_5998);
and U7532 (N_7532,N_382,N_2247);
and U7533 (N_7533,N_4683,N_5384);
nand U7534 (N_7534,N_1006,N_2176);
nand U7535 (N_7535,N_2707,N_637);
and U7536 (N_7536,N_5408,N_3589);
nand U7537 (N_7537,N_2511,N_3720);
or U7538 (N_7538,N_3175,N_5913);
nand U7539 (N_7539,N_4407,N_3955);
and U7540 (N_7540,N_2342,N_5756);
nor U7541 (N_7541,N_5309,N_3850);
nand U7542 (N_7542,N_1675,N_5269);
xor U7543 (N_7543,N_1493,N_3922);
nor U7544 (N_7544,N_4991,N_1679);
or U7545 (N_7545,N_1568,N_2539);
nor U7546 (N_7546,N_3061,N_1551);
nor U7547 (N_7547,N_3692,N_3078);
or U7548 (N_7548,N_2711,N_124);
and U7549 (N_7549,N_4692,N_791);
nand U7550 (N_7550,N_4630,N_3745);
or U7551 (N_7551,N_4233,N_1844);
and U7552 (N_7552,N_5437,N_2254);
nand U7553 (N_7553,N_913,N_3935);
nand U7554 (N_7554,N_2735,N_104);
or U7555 (N_7555,N_5760,N_3855);
nor U7556 (N_7556,N_109,N_5332);
nand U7557 (N_7557,N_5971,N_4199);
and U7558 (N_7558,N_4826,N_1337);
xor U7559 (N_7559,N_5448,N_5469);
nand U7560 (N_7560,N_5627,N_2680);
and U7561 (N_7561,N_189,N_2134);
nand U7562 (N_7562,N_4674,N_3806);
or U7563 (N_7563,N_4690,N_2899);
nand U7564 (N_7564,N_577,N_5829);
nand U7565 (N_7565,N_5762,N_3967);
and U7566 (N_7566,N_1803,N_5737);
nor U7567 (N_7567,N_1166,N_4002);
nand U7568 (N_7568,N_5059,N_3127);
or U7569 (N_7569,N_201,N_4012);
xnor U7570 (N_7570,N_943,N_4517);
or U7571 (N_7571,N_2353,N_3034);
or U7572 (N_7572,N_1827,N_5649);
xor U7573 (N_7573,N_666,N_1111);
nor U7574 (N_7574,N_62,N_5626);
and U7575 (N_7575,N_3694,N_2785);
or U7576 (N_7576,N_5741,N_1779);
and U7577 (N_7577,N_5703,N_1513);
and U7578 (N_7578,N_853,N_2684);
and U7579 (N_7579,N_4408,N_2208);
and U7580 (N_7580,N_4832,N_261);
and U7581 (N_7581,N_2760,N_1775);
nand U7582 (N_7582,N_5140,N_2736);
xor U7583 (N_7583,N_2655,N_5331);
nand U7584 (N_7584,N_217,N_4224);
or U7585 (N_7585,N_1250,N_3782);
xor U7586 (N_7586,N_4881,N_2007);
nor U7587 (N_7587,N_3499,N_3817);
or U7588 (N_7588,N_3914,N_37);
xnor U7589 (N_7589,N_3079,N_2059);
and U7590 (N_7590,N_2852,N_5032);
nor U7591 (N_7591,N_1468,N_2928);
xnor U7592 (N_7592,N_4302,N_5822);
nand U7593 (N_7593,N_5606,N_3919);
nor U7594 (N_7594,N_24,N_3501);
nand U7595 (N_7595,N_118,N_523);
nor U7596 (N_7596,N_3218,N_311);
nor U7597 (N_7597,N_4964,N_755);
or U7598 (N_7598,N_1943,N_3411);
or U7599 (N_7599,N_2722,N_4891);
nor U7600 (N_7600,N_5669,N_1356);
or U7601 (N_7601,N_1172,N_1860);
nor U7602 (N_7602,N_690,N_939);
nor U7603 (N_7603,N_4163,N_1203);
and U7604 (N_7604,N_1994,N_4774);
and U7605 (N_7605,N_2237,N_2728);
nand U7606 (N_7606,N_1630,N_4450);
nand U7607 (N_7607,N_1678,N_554);
and U7608 (N_7608,N_5409,N_919);
xor U7609 (N_7609,N_4867,N_621);
nor U7610 (N_7610,N_2202,N_2269);
or U7611 (N_7611,N_4589,N_1633);
nand U7612 (N_7612,N_4179,N_2532);
xor U7613 (N_7613,N_5985,N_471);
and U7614 (N_7614,N_1362,N_5814);
nor U7615 (N_7615,N_4792,N_3048);
nor U7616 (N_7616,N_4739,N_2768);
or U7617 (N_7617,N_4965,N_3149);
nand U7618 (N_7618,N_3409,N_1301);
or U7619 (N_7619,N_4219,N_2167);
or U7620 (N_7620,N_1448,N_4303);
or U7621 (N_7621,N_648,N_2379);
nand U7622 (N_7622,N_4267,N_2091);
nand U7623 (N_7623,N_297,N_4196);
nor U7624 (N_7624,N_5719,N_929);
or U7625 (N_7625,N_4106,N_1251);
xor U7626 (N_7626,N_1527,N_3432);
nor U7627 (N_7627,N_5803,N_3108);
and U7628 (N_7628,N_3825,N_281);
nor U7629 (N_7629,N_4906,N_123);
and U7630 (N_7630,N_2221,N_5965);
nand U7631 (N_7631,N_3781,N_1440);
nor U7632 (N_7632,N_1938,N_4885);
or U7633 (N_7633,N_4695,N_4916);
nand U7634 (N_7634,N_4861,N_179);
xnor U7635 (N_7635,N_3332,N_615);
xor U7636 (N_7636,N_5070,N_2513);
nand U7637 (N_7637,N_2407,N_4354);
and U7638 (N_7638,N_2518,N_5479);
and U7639 (N_7639,N_1600,N_3359);
and U7640 (N_7640,N_285,N_2215);
nor U7641 (N_7641,N_1486,N_5557);
nor U7642 (N_7642,N_1893,N_2836);
and U7643 (N_7643,N_5921,N_5181);
nand U7644 (N_7644,N_5214,N_90);
nand U7645 (N_7645,N_5130,N_1682);
nor U7646 (N_7646,N_1694,N_888);
xnor U7647 (N_7647,N_373,N_5502);
nand U7648 (N_7648,N_2041,N_4845);
nor U7649 (N_7649,N_3483,N_1680);
nand U7650 (N_7650,N_1088,N_2331);
nor U7651 (N_7651,N_2137,N_3558);
xnor U7652 (N_7652,N_4937,N_1395);
nand U7653 (N_7653,N_618,N_2008);
nand U7654 (N_7654,N_3755,N_5245);
nor U7655 (N_7655,N_1753,N_411);
nand U7656 (N_7656,N_4856,N_79);
nand U7657 (N_7657,N_3592,N_2960);
nand U7658 (N_7658,N_4696,N_2887);
nor U7659 (N_7659,N_1420,N_66);
and U7660 (N_7660,N_4347,N_1007);
nor U7661 (N_7661,N_1404,N_783);
xor U7662 (N_7662,N_5823,N_5860);
nand U7663 (N_7663,N_2584,N_2957);
xnor U7664 (N_7664,N_4952,N_5500);
or U7665 (N_7665,N_3260,N_891);
nand U7666 (N_7666,N_4191,N_3893);
nor U7667 (N_7667,N_1437,N_2660);
xnor U7668 (N_7668,N_670,N_1500);
nor U7669 (N_7669,N_4915,N_2737);
nor U7670 (N_7670,N_3265,N_2753);
xnor U7671 (N_7671,N_2819,N_2177);
xor U7672 (N_7672,N_4007,N_1150);
nand U7673 (N_7673,N_2740,N_2373);
and U7674 (N_7674,N_4793,N_3303);
or U7675 (N_7675,N_2282,N_2588);
and U7676 (N_7676,N_5460,N_2952);
and U7677 (N_7677,N_3691,N_2929);
nor U7678 (N_7678,N_4593,N_2194);
nor U7679 (N_7679,N_5771,N_5011);
xor U7680 (N_7680,N_2417,N_4786);
and U7681 (N_7681,N_5710,N_4208);
nor U7682 (N_7682,N_3322,N_5064);
nand U7683 (N_7683,N_5539,N_1138);
nand U7684 (N_7684,N_1375,N_2544);
and U7685 (N_7685,N_2193,N_2420);
xor U7686 (N_7686,N_3135,N_4592);
nand U7687 (N_7687,N_4814,N_3881);
or U7688 (N_7688,N_4087,N_2536);
xor U7689 (N_7689,N_5911,N_3690);
nor U7690 (N_7690,N_4356,N_4661);
and U7691 (N_7691,N_77,N_3063);
and U7692 (N_7692,N_5836,N_5909);
and U7693 (N_7693,N_1147,N_876);
or U7694 (N_7694,N_5004,N_3677);
and U7695 (N_7695,N_347,N_5106);
nor U7696 (N_7696,N_3373,N_3169);
nor U7697 (N_7697,N_1712,N_3873);
nor U7698 (N_7698,N_782,N_4835);
nor U7699 (N_7699,N_4402,N_4653);
or U7700 (N_7700,N_4888,N_3556);
and U7701 (N_7701,N_145,N_1751);
nand U7702 (N_7702,N_4368,N_1565);
or U7703 (N_7703,N_3319,N_2956);
xnor U7704 (N_7704,N_3041,N_5916);
or U7705 (N_7705,N_839,N_1563);
nor U7706 (N_7706,N_1390,N_2634);
nor U7707 (N_7707,N_4426,N_3758);
and U7708 (N_7708,N_4954,N_3267);
and U7709 (N_7709,N_1396,N_2390);
and U7710 (N_7710,N_5550,N_1646);
nand U7711 (N_7711,N_829,N_5179);
xor U7712 (N_7712,N_601,N_2065);
nor U7713 (N_7713,N_2659,N_1849);
nor U7714 (N_7714,N_2880,N_4458);
nand U7715 (N_7715,N_199,N_3740);
xor U7716 (N_7716,N_5682,N_5024);
nor U7717 (N_7717,N_3222,N_468);
xor U7718 (N_7718,N_121,N_2912);
xor U7719 (N_7719,N_2322,N_2816);
nand U7720 (N_7720,N_4213,N_2203);
xnor U7721 (N_7721,N_2916,N_150);
or U7722 (N_7722,N_1713,N_2028);
or U7723 (N_7723,N_4819,N_4403);
nor U7724 (N_7724,N_156,N_833);
nor U7725 (N_7725,N_4238,N_4733);
or U7726 (N_7726,N_3868,N_2479);
nor U7727 (N_7727,N_3948,N_1985);
xnor U7728 (N_7728,N_2440,N_1084);
and U7729 (N_7729,N_1575,N_3622);
and U7730 (N_7730,N_1883,N_2182);
nor U7731 (N_7731,N_3607,N_3272);
and U7732 (N_7732,N_4455,N_2346);
nor U7733 (N_7733,N_3382,N_1040);
and U7734 (N_7734,N_2712,N_5100);
nor U7735 (N_7735,N_2558,N_410);
nand U7736 (N_7736,N_2073,N_1852);
nand U7737 (N_7737,N_3984,N_4395);
nand U7738 (N_7738,N_5946,N_784);
nor U7739 (N_7739,N_794,N_1672);
nor U7740 (N_7740,N_4711,N_5440);
or U7741 (N_7741,N_3896,N_2312);
nor U7742 (N_7742,N_5088,N_2528);
nand U7743 (N_7743,N_1340,N_5429);
or U7744 (N_7744,N_2470,N_4584);
or U7745 (N_7745,N_1013,N_3569);
and U7746 (N_7746,N_4326,N_5643);
nor U7747 (N_7747,N_5353,N_1183);
nand U7748 (N_7748,N_1492,N_1914);
or U7749 (N_7749,N_1148,N_657);
nand U7750 (N_7750,N_3876,N_1898);
xor U7751 (N_7751,N_4209,N_1476);
nand U7752 (N_7752,N_4485,N_1427);
nand U7753 (N_7753,N_5493,N_4613);
nand U7754 (N_7754,N_873,N_2228);
and U7755 (N_7755,N_4349,N_4021);
or U7756 (N_7756,N_3224,N_1141);
and U7757 (N_7757,N_1511,N_2581);
or U7758 (N_7758,N_4700,N_4790);
nand U7759 (N_7759,N_2897,N_5929);
nand U7760 (N_7760,N_3112,N_1874);
nor U7761 (N_7761,N_3456,N_5092);
and U7762 (N_7762,N_1487,N_5763);
and U7763 (N_7763,N_2672,N_3731);
nand U7764 (N_7764,N_3335,N_3317);
and U7765 (N_7765,N_4773,N_1596);
and U7766 (N_7766,N_5,N_4324);
nand U7767 (N_7767,N_5657,N_642);
or U7768 (N_7768,N_1789,N_1567);
nand U7769 (N_7769,N_5133,N_1561);
nand U7770 (N_7770,N_4038,N_5812);
and U7771 (N_7771,N_4055,N_25);
xnor U7772 (N_7772,N_1604,N_1237);
nand U7773 (N_7773,N_2449,N_935);
or U7774 (N_7774,N_2743,N_3601);
nor U7775 (N_7775,N_702,N_1218);
nor U7776 (N_7776,N_4344,N_3367);
nand U7777 (N_7777,N_630,N_4839);
or U7778 (N_7778,N_1697,N_2035);
nand U7779 (N_7779,N_3585,N_678);
and U7780 (N_7780,N_3270,N_1011);
nor U7781 (N_7781,N_1226,N_3309);
nor U7782 (N_7782,N_1319,N_2885);
and U7783 (N_7783,N_4217,N_2738);
and U7784 (N_7784,N_2484,N_4534);
and U7785 (N_7785,N_2309,N_2826);
nand U7786 (N_7786,N_4863,N_610);
nand U7787 (N_7787,N_3430,N_3866);
or U7788 (N_7788,N_3165,N_4059);
and U7789 (N_7789,N_3468,N_5318);
and U7790 (N_7790,N_1032,N_2725);
nand U7791 (N_7791,N_442,N_1292);
nand U7792 (N_7792,N_1034,N_4972);
nor U7793 (N_7793,N_4967,N_5293);
nand U7794 (N_7794,N_5706,N_173);
xnor U7795 (N_7795,N_1024,N_4466);
and U7796 (N_7796,N_1609,N_4842);
xor U7797 (N_7797,N_3500,N_5147);
or U7798 (N_7798,N_4875,N_5754);
and U7799 (N_7799,N_2250,N_5282);
nand U7800 (N_7800,N_5156,N_3157);
and U7801 (N_7801,N_5006,N_1835);
xnor U7802 (N_7802,N_1169,N_4023);
nand U7803 (N_7803,N_4397,N_2316);
nand U7804 (N_7804,N_2145,N_693);
or U7805 (N_7805,N_4897,N_5025);
xor U7806 (N_7806,N_3462,N_5941);
nor U7807 (N_7807,N_1762,N_1805);
or U7808 (N_7808,N_2024,N_962);
nor U7809 (N_7809,N_3139,N_679);
or U7810 (N_7810,N_4857,N_5038);
or U7811 (N_7811,N_986,N_1597);
or U7812 (N_7812,N_436,N_884);
nand U7813 (N_7813,N_675,N_580);
nand U7814 (N_7814,N_663,N_2966);
nand U7815 (N_7815,N_4824,N_3871);
nand U7816 (N_7816,N_654,N_4285);
and U7817 (N_7817,N_3484,N_3397);
nor U7818 (N_7818,N_5920,N_4508);
or U7819 (N_7819,N_5376,N_3597);
xnor U7820 (N_7820,N_2399,N_1954);
or U7821 (N_7821,N_1663,N_5784);
and U7822 (N_7822,N_5359,N_956);
or U7823 (N_7823,N_4295,N_2691);
or U7824 (N_7824,N_4651,N_1182);
or U7825 (N_7825,N_4323,N_157);
nor U7826 (N_7826,N_3828,N_332);
nand U7827 (N_7827,N_2158,N_329);
and U7828 (N_7828,N_3315,N_2640);
nand U7829 (N_7829,N_4721,N_1959);
and U7830 (N_7830,N_2701,N_4134);
nand U7831 (N_7831,N_2365,N_3353);
or U7832 (N_7832,N_5906,N_3832);
nand U7833 (N_7833,N_4121,N_730);
nor U7834 (N_7834,N_1355,N_1683);
nor U7835 (N_7835,N_4474,N_2017);
and U7836 (N_7836,N_2702,N_2207);
and U7837 (N_7837,N_3459,N_544);
nand U7838 (N_7838,N_5094,N_3796);
nand U7839 (N_7839,N_2285,N_4934);
or U7840 (N_7840,N_3679,N_722);
or U7841 (N_7841,N_2359,N_3019);
or U7842 (N_7842,N_2173,N_4433);
and U7843 (N_7843,N_2085,N_5997);
or U7844 (N_7844,N_283,N_3431);
and U7845 (N_7845,N_3954,N_141);
nor U7846 (N_7846,N_1645,N_3110);
nor U7847 (N_7847,N_5786,N_4524);
or U7848 (N_7848,N_3653,N_3875);
xor U7849 (N_7849,N_3264,N_1540);
nor U7850 (N_7850,N_2168,N_2815);
or U7851 (N_7851,N_912,N_4350);
nand U7852 (N_7852,N_1053,N_4610);
and U7853 (N_7853,N_810,N_2362);
and U7854 (N_7854,N_5875,N_434);
xnor U7855 (N_7855,N_5779,N_3625);
and U7856 (N_7856,N_207,N_4082);
or U7857 (N_7857,N_130,N_443);
or U7858 (N_7858,N_4457,N_1993);
nor U7859 (N_7859,N_134,N_1280);
nor U7860 (N_7860,N_3852,N_2371);
nand U7861 (N_7861,N_1296,N_1760);
or U7862 (N_7862,N_298,N_1923);
and U7863 (N_7863,N_3596,N_2567);
or U7864 (N_7864,N_3414,N_3344);
nand U7865 (N_7865,N_2308,N_5141);
xor U7866 (N_7866,N_3695,N_1785);
nor U7867 (N_7867,N_3971,N_2903);
nor U7868 (N_7868,N_3554,N_4778);
and U7869 (N_7869,N_1061,N_534);
nand U7870 (N_7870,N_2397,N_3618);
nand U7871 (N_7871,N_5933,N_2174);
xnor U7872 (N_7872,N_2112,N_5412);
or U7873 (N_7873,N_3290,N_487);
nor U7874 (N_7874,N_5152,N_691);
and U7875 (N_7875,N_4628,N_2000);
or U7876 (N_7876,N_1888,N_3765);
nand U7877 (N_7877,N_2589,N_2998);
or U7878 (N_7878,N_132,N_2027);
nor U7879 (N_7879,N_629,N_61);
xnor U7880 (N_7880,N_5187,N_3764);
and U7881 (N_7881,N_4890,N_3056);
and U7882 (N_7882,N_5001,N_2206);
and U7883 (N_7883,N_3798,N_1343);
and U7884 (N_7884,N_4940,N_3457);
or U7885 (N_7885,N_1539,N_5267);
or U7886 (N_7886,N_1556,N_49);
and U7887 (N_7887,N_4011,N_2151);
and U7888 (N_7888,N_3338,N_2394);
nand U7889 (N_7889,N_2579,N_858);
and U7890 (N_7890,N_3038,N_5464);
or U7891 (N_7891,N_2537,N_1207);
nand U7892 (N_7892,N_2964,N_2747);
or U7893 (N_7893,N_1661,N_3241);
and U7894 (N_7894,N_1598,N_1465);
or U7895 (N_7895,N_3476,N_4234);
nor U7896 (N_7896,N_1123,N_5665);
or U7897 (N_7897,N_1879,N_3053);
and U7898 (N_7898,N_3913,N_927);
and U7899 (N_7899,N_4777,N_5988);
nor U7900 (N_7900,N_536,N_1777);
and U7901 (N_7901,N_5166,N_1423);
nand U7902 (N_7902,N_3421,N_4073);
nor U7903 (N_7903,N_402,N_3400);
and U7904 (N_7904,N_312,N_5405);
or U7905 (N_7905,N_1634,N_4480);
nand U7906 (N_7906,N_5895,N_4629);
xnor U7907 (N_7907,N_1800,N_2514);
xor U7908 (N_7908,N_3324,N_2643);
or U7909 (N_7909,N_3003,N_2628);
or U7910 (N_7910,N_848,N_331);
or U7911 (N_7911,N_4239,N_1018);
nor U7912 (N_7912,N_2688,N_334);
nand U7913 (N_7913,N_2983,N_2967);
nand U7914 (N_7914,N_3274,N_5372);
nor U7915 (N_7915,N_3412,N_1072);
nand U7916 (N_7916,N_2599,N_3815);
and U7917 (N_7917,N_4657,N_1422);
nand U7918 (N_7918,N_4554,N_3498);
nand U7919 (N_7919,N_3043,N_214);
nand U7920 (N_7920,N_2694,N_5305);
and U7921 (N_7921,N_3775,N_178);
xnor U7922 (N_7922,N_5750,N_4178);
nand U7923 (N_7923,N_4237,N_3381);
or U7924 (N_7924,N_4071,N_5766);
or U7925 (N_7925,N_2246,N_337);
nor U7926 (N_7926,N_5937,N_1379);
nor U7927 (N_7927,N_2234,N_151);
or U7928 (N_7928,N_267,N_5987);
nand U7929 (N_7929,N_1560,N_5878);
and U7930 (N_7930,N_5683,N_5167);
nand U7931 (N_7931,N_1112,N_2471);
xnor U7932 (N_7932,N_3238,N_1977);
or U7933 (N_7933,N_423,N_3302);
or U7934 (N_7934,N_2337,N_3440);
or U7935 (N_7935,N_2299,N_2344);
or U7936 (N_7936,N_4971,N_2305);
nand U7937 (N_7937,N_2255,N_1160);
and U7938 (N_7938,N_1981,N_2494);
and U7939 (N_7939,N_1998,N_575);
nand U7940 (N_7940,N_3701,N_165);
nand U7941 (N_7941,N_4214,N_4331);
and U7942 (N_7942,N_745,N_318);
nand U7943 (N_7943,N_825,N_1078);
and U7944 (N_7944,N_5615,N_717);
nand U7945 (N_7945,N_4535,N_3724);
and U7946 (N_7946,N_2360,N_2490);
xor U7947 (N_7947,N_4319,N_2831);
and U7948 (N_7948,N_1127,N_3422);
xnor U7949 (N_7949,N_3688,N_3726);
and U7950 (N_7950,N_653,N_3234);
nor U7951 (N_7951,N_4427,N_3349);
nand U7952 (N_7952,N_1546,N_572);
and U7953 (N_7953,N_4139,N_1657);
and U7954 (N_7954,N_5739,N_459);
nor U7955 (N_7955,N_5892,N_5261);
and U7956 (N_7956,N_701,N_5548);
and U7957 (N_7957,N_4996,N_2975);
and U7958 (N_7958,N_1357,N_5810);
nand U7959 (N_7959,N_3684,N_108);
and U7960 (N_7960,N_636,N_4688);
nand U7961 (N_7961,N_2548,N_1044);
nand U7962 (N_7962,N_937,N_2253);
or U7963 (N_7963,N_3675,N_1313);
nor U7964 (N_7964,N_4005,N_4959);
or U7965 (N_7965,N_4334,N_3612);
or U7966 (N_7966,N_2002,N_3516);
xor U7967 (N_7967,N_1472,N_949);
nand U7968 (N_7968,N_1937,N_869);
xnor U7969 (N_7969,N_2787,N_324);
or U7970 (N_7970,N_2758,N_1397);
nor U7971 (N_7971,N_2113,N_1768);
nor U7972 (N_7972,N_4300,N_1654);
or U7973 (N_7973,N_1353,N_5621);
xnor U7974 (N_7974,N_5513,N_2988);
and U7975 (N_7975,N_249,N_643);
and U7976 (N_7976,N_4338,N_5310);
or U7977 (N_7977,N_2453,N_4254);
xor U7978 (N_7978,N_5253,N_3357);
or U7979 (N_7979,N_5043,N_3915);
and U7980 (N_7980,N_2651,N_5134);
or U7981 (N_7981,N_2505,N_4539);
nand U7982 (N_7982,N_1271,N_5127);
or U7983 (N_7983,N_1091,N_4546);
and U7984 (N_7984,N_1931,N_4636);
xor U7985 (N_7985,N_1613,N_75);
nand U7986 (N_7986,N_1892,N_5394);
and U7987 (N_7987,N_4868,N_5058);
or U7988 (N_7988,N_1393,N_5730);
and U7989 (N_7989,N_2797,N_669);
nor U7990 (N_7990,N_5165,N_1444);
nor U7991 (N_7991,N_5640,N_5700);
and U7992 (N_7992,N_4391,N_4494);
xor U7993 (N_7993,N_1709,N_4756);
or U7994 (N_7994,N_3968,N_5202);
nand U7995 (N_7995,N_2566,N_3822);
nand U7996 (N_7996,N_5312,N_3686);
or U7997 (N_7997,N_1973,N_1405);
xor U7998 (N_7998,N_4222,N_4525);
or U7999 (N_7999,N_2942,N_183);
and U8000 (N_8000,N_3325,N_4795);
or U8001 (N_8001,N_847,N_3749);
and U8002 (N_8002,N_500,N_1875);
nor U8003 (N_8003,N_2463,N_2742);
nand U8004 (N_8004,N_3014,N_273);
nor U8005 (N_8005,N_5263,N_991);
or U8006 (N_8006,N_2197,N_2606);
or U8007 (N_8007,N_1776,N_5609);
or U8008 (N_8008,N_826,N_3727);
or U8009 (N_8009,N_1670,N_5717);
or U8010 (N_8010,N_3836,N_5071);
and U8011 (N_8011,N_4297,N_4576);
and U8012 (N_8012,N_4328,N_3687);
and U8013 (N_8013,N_3751,N_4363);
and U8014 (N_8014,N_5427,N_1503);
or U8015 (N_8015,N_4808,N_5137);
nand U8016 (N_8016,N_2723,N_1194);
or U8017 (N_8017,N_4280,N_2434);
and U8018 (N_8018,N_5588,N_5579);
and U8019 (N_8019,N_1876,N_1491);
or U8020 (N_8020,N_3101,N_557);
and U8021 (N_8021,N_3341,N_5414);
nand U8022 (N_8022,N_3370,N_2248);
xor U8023 (N_8023,N_4616,N_4144);
or U8024 (N_8024,N_2329,N_2489);
nand U8025 (N_8025,N_793,N_5564);
or U8026 (N_8026,N_5477,N_1161);
or U8027 (N_8027,N_983,N_5915);
and U8028 (N_8028,N_4030,N_821);
or U8029 (N_8029,N_3177,N_4061);
nor U8030 (N_8030,N_4313,N_4499);
or U8031 (N_8031,N_681,N_4409);
nand U8032 (N_8032,N_4052,N_616);
or U8033 (N_8033,N_1435,N_1843);
or U8034 (N_8034,N_4859,N_1187);
nor U8035 (N_8035,N_505,N_2808);
nor U8036 (N_8036,N_1961,N_1584);
nor U8037 (N_8037,N_5886,N_2264);
nand U8038 (N_8038,N_52,N_708);
nand U8039 (N_8039,N_4287,N_5023);
xnor U8040 (N_8040,N_1320,N_4113);
nand U8041 (N_8041,N_4221,N_1345);
nor U8042 (N_8042,N_5030,N_3221);
and U8043 (N_8043,N_694,N_368);
nor U8044 (N_8044,N_2286,N_4248);
xor U8045 (N_8045,N_2330,N_5740);
and U8046 (N_8046,N_452,N_1100);
nor U8047 (N_8047,N_250,N_389);
and U8048 (N_8048,N_4241,N_3194);
or U8049 (N_8049,N_2169,N_1689);
and U8050 (N_8050,N_5155,N_1691);
nand U8051 (N_8051,N_4161,N_571);
and U8052 (N_8052,N_3945,N_775);
or U8053 (N_8053,N_980,N_3800);
or U8054 (N_8054,N_2486,N_1370);
or U8055 (N_8055,N_4958,N_3639);
nand U8056 (N_8056,N_4153,N_3472);
and U8057 (N_8057,N_5885,N_2717);
or U8058 (N_8058,N_2183,N_5288);
nor U8059 (N_8059,N_4410,N_5515);
nand U8060 (N_8060,N_2615,N_2227);
or U8061 (N_8061,N_3768,N_1857);
nand U8062 (N_8062,N_4531,N_4282);
xor U8063 (N_8063,N_2062,N_3268);
or U8064 (N_8064,N_3240,N_4779);
and U8065 (N_8065,N_5180,N_1867);
nor U8066 (N_8066,N_3481,N_3884);
and U8067 (N_8067,N_3145,N_604);
xor U8068 (N_8068,N_5079,N_1038);
or U8069 (N_8069,N_5246,N_112);
or U8070 (N_8070,N_1553,N_2349);
nand U8071 (N_8071,N_1180,N_647);
nand U8072 (N_8072,N_4054,N_3809);
xnor U8073 (N_8073,N_1763,N_1895);
or U8074 (N_8074,N_1028,N_2117);
and U8075 (N_8075,N_1673,N_3813);
nand U8076 (N_8076,N_4770,N_3150);
and U8077 (N_8077,N_4634,N_2759);
nor U8078 (N_8078,N_1580,N_4136);
or U8079 (N_8079,N_1102,N_475);
nor U8080 (N_8080,N_1329,N_1520);
nor U8081 (N_8081,N_5917,N_3391);
or U8082 (N_8082,N_687,N_5438);
or U8083 (N_8083,N_187,N_446);
or U8084 (N_8084,N_3413,N_1625);
nand U8085 (N_8085,N_3232,N_3036);
and U8086 (N_8086,N_2530,N_131);
or U8087 (N_8087,N_2380,N_4798);
and U8088 (N_8088,N_5206,N_739);
and U8089 (N_8089,N_5645,N_1582);
nor U8090 (N_8090,N_2457,N_597);
nor U8091 (N_8091,N_2796,N_2428);
and U8092 (N_8092,N_2015,N_1909);
and U8093 (N_8093,N_4789,N_1933);
nor U8094 (N_8094,N_1219,N_4599);
nor U8095 (N_8095,N_4801,N_4056);
nor U8096 (N_8096,N_5631,N_2411);
nor U8097 (N_8097,N_2718,N_4272);
or U8098 (N_8098,N_1510,N_860);
nand U8099 (N_8099,N_4941,N_4823);
and U8100 (N_8100,N_2756,N_1471);
and U8101 (N_8101,N_3814,N_2393);
xnor U8102 (N_8102,N_1859,N_4111);
and U8103 (N_8103,N_4633,N_5704);
nand U8104 (N_8104,N_366,N_136);
nand U8105 (N_8105,N_5487,N_4878);
nor U8106 (N_8106,N_2020,N_1284);
nor U8107 (N_8107,N_3007,N_1076);
xor U8108 (N_8108,N_4148,N_4447);
xor U8109 (N_8109,N_262,N_1368);
nor U8110 (N_8110,N_2543,N_1273);
and U8111 (N_8111,N_1332,N_684);
or U8112 (N_8112,N_5157,N_197);
or U8113 (N_8113,N_1810,N_5329);
nor U8114 (N_8114,N_386,N_5948);
and U8115 (N_8115,N_5576,N_1968);
and U8116 (N_8116,N_2244,N_710);
nand U8117 (N_8117,N_2496,N_4383);
nand U8118 (N_8118,N_5767,N_3805);
or U8119 (N_8119,N_1769,N_275);
and U8120 (N_8120,N_2650,N_3714);
or U8121 (N_8121,N_3210,N_2696);
and U8122 (N_8122,N_1872,N_2001);
nand U8123 (N_8123,N_476,N_461);
nor U8124 (N_8124,N_166,N_4949);
xor U8125 (N_8125,N_1941,N_3734);
or U8126 (N_8126,N_3371,N_1118);
and U8127 (N_8127,N_1838,N_3882);
or U8128 (N_8128,N_3231,N_2398);
and U8129 (N_8129,N_5828,N_1475);
nor U8130 (N_8130,N_5208,N_1433);
xnor U8131 (N_8131,N_2450,N_2812);
nor U8132 (N_8132,N_4578,N_4304);
and U8133 (N_8133,N_316,N_2774);
nand U8134 (N_8134,N_5274,N_1622);
xor U8135 (N_8135,N_683,N_2600);
or U8136 (N_8136,N_5146,N_3037);
nand U8137 (N_8137,N_3347,N_3350);
nor U8138 (N_8138,N_2790,N_673);
or U8139 (N_8139,N_1173,N_2869);
nor U8140 (N_8140,N_1750,N_3167);
xor U8141 (N_8141,N_5694,N_5029);
nor U8142 (N_8142,N_3263,N_4100);
or U8143 (N_8143,N_1212,N_1306);
nand U8144 (N_8144,N_3712,N_524);
nor U8145 (N_8145,N_291,N_4470);
and U8146 (N_8146,N_3575,N_921);
nor U8147 (N_8147,N_460,N_3890);
and U8148 (N_8148,N_4679,N_435);
or U8149 (N_8149,N_1256,N_107);
nand U8150 (N_8150,N_5368,N_4094);
nand U8151 (N_8151,N_4849,N_4223);
and U8152 (N_8152,N_2646,N_2733);
or U8153 (N_8153,N_5953,N_5664);
and U8154 (N_8154,N_3209,N_1025);
nor U8155 (N_8155,N_4673,N_5008);
and U8156 (N_8156,N_2542,N_3671);
nor U8157 (N_8157,N_3506,N_4652);
or U8158 (N_8158,N_3473,N_5835);
nor U8159 (N_8159,N_4104,N_5121);
and U8160 (N_8160,N_1009,N_5898);
xnor U8161 (N_8161,N_440,N_3759);
and U8162 (N_8162,N_185,N_1899);
or U8163 (N_8163,N_1516,N_4995);
xnor U8164 (N_8164,N_1702,N_5624);
and U8165 (N_8165,N_2033,N_3859);
nor U8166 (N_8166,N_733,N_2933);
and U8167 (N_8167,N_3131,N_4741);
or U8168 (N_8168,N_1802,N_1976);
and U8169 (N_8169,N_521,N_3792);
and U8170 (N_8170,N_4993,N_5549);
nor U8171 (N_8171,N_3095,N_3566);
nor U8172 (N_8172,N_2667,N_2478);
and U8173 (N_8173,N_1693,N_3076);
or U8174 (N_8174,N_4392,N_4336);
and U8175 (N_8175,N_1069,N_221);
nand U8176 (N_8176,N_2894,N_3668);
nor U8177 (N_8177,N_4686,N_1949);
nor U8178 (N_8178,N_3906,N_5778);
nand U8179 (N_8179,N_1905,N_2442);
or U8180 (N_8180,N_4899,N_3902);
or U8181 (N_8181,N_737,N_4066);
or U8182 (N_8182,N_4874,N_3144);
and U8183 (N_8183,N_2745,N_569);
nand U8184 (N_8184,N_4235,N_984);
or U8185 (N_8185,N_4096,N_1277);
or U8186 (N_8186,N_3870,N_1413);
nor U8187 (N_8187,N_415,N_4689);
or U8188 (N_8188,N_1809,N_1509);
nand U8189 (N_8189,N_5654,N_5595);
nand U8190 (N_8190,N_2909,N_971);
or U8191 (N_8191,N_2273,N_587);
or U8192 (N_8192,N_5806,N_2149);
or U8193 (N_8193,N_3026,N_3387);
xnor U8194 (N_8194,N_4024,N_585);
or U8195 (N_8195,N_1701,N_5995);
and U8196 (N_8196,N_4035,N_480);
and U8197 (N_8197,N_5577,N_133);
and U8198 (N_8198,N_5765,N_4604);
and U8199 (N_8199,N_3204,N_2697);
or U8200 (N_8200,N_3757,N_3467);
and U8201 (N_8201,N_139,N_4886);
nand U8202 (N_8202,N_5912,N_835);
and U8203 (N_8203,N_4006,N_1380);
nor U8204 (N_8204,N_1045,N_1381);
xor U8205 (N_8205,N_1552,N_1303);
xor U8206 (N_8206,N_5213,N_2654);
and U8207 (N_8207,N_3197,N_2431);
xor U8208 (N_8208,N_3187,N_1136);
nand U8209 (N_8209,N_3351,N_5398);
or U8210 (N_8210,N_3946,N_4167);
or U8211 (N_8211,N_5593,N_3146);
or U8212 (N_8212,N_5123,N_3271);
nand U8213 (N_8213,N_5143,N_2726);
nor U8214 (N_8214,N_3358,N_4791);
and U8215 (N_8215,N_579,N_481);
and U8216 (N_8216,N_195,N_1869);
nand U8217 (N_8217,N_1164,N_1594);
and U8218 (N_8218,N_628,N_5105);
nand U8219 (N_8219,N_4463,N_5431);
nor U8220 (N_8220,N_425,N_4255);
xnor U8221 (N_8221,N_2069,N_3010);
xor U8222 (N_8222,N_4445,N_2289);
or U8223 (N_8223,N_5698,N_2148);
nand U8224 (N_8224,N_2582,N_404);
and U8225 (N_8225,N_4242,N_2803);
nor U8226 (N_8226,N_594,N_1206);
xnor U8227 (N_8227,N_4583,N_3369);
nand U8228 (N_8228,N_5986,N_3819);
nor U8229 (N_8229,N_1351,N_2315);
nor U8230 (N_8230,N_4362,N_3648);
and U8231 (N_8231,N_3982,N_4931);
and U8232 (N_8232,N_3887,N_2871);
xor U8233 (N_8233,N_3269,N_4523);
nor U8234 (N_8234,N_2072,N_5650);
nand U8235 (N_8235,N_3027,N_3977);
nand U8236 (N_8236,N_753,N_2107);
and U8237 (N_8237,N_3435,N_1807);
or U8238 (N_8238,N_5973,N_5729);
nor U8239 (N_8239,N_1198,N_668);
or U8240 (N_8240,N_1217,N_1000);
and U8241 (N_8241,N_1853,N_516);
and U8242 (N_8242,N_5396,N_489);
and U8243 (N_8243,N_444,N_3304);
and U8244 (N_8244,N_5392,N_328);
nand U8245 (N_8245,N_2944,N_4655);
or U8246 (N_8246,N_58,N_4649);
or U8247 (N_8247,N_538,N_2115);
nor U8248 (N_8248,N_3158,N_4076);
nand U8249 (N_8249,N_3779,N_5317);
and U8250 (N_8250,N_5685,N_705);
or U8251 (N_8251,N_5195,N_3008);
nand U8252 (N_8252,N_1864,N_5785);
or U8253 (N_8253,N_4321,N_2715);
nand U8254 (N_8254,N_1979,N_3293);
nor U8255 (N_8255,N_1695,N_2423);
and U8256 (N_8256,N_763,N_1532);
nand U8257 (N_8257,N_3217,N_4137);
nand U8258 (N_8258,N_607,N_844);
nor U8259 (N_8259,N_3438,N_2443);
nor U8260 (N_8260,N_4320,N_5063);
nand U8261 (N_8261,N_4978,N_5120);
nor U8262 (N_8262,N_1267,N_1162);
nand U8263 (N_8263,N_5233,N_2829);
or U8264 (N_8264,N_2531,N_353);
nand U8265 (N_8265,N_3926,N_3600);
xor U8266 (N_8266,N_970,N_751);
nor U8267 (N_8267,N_2982,N_2629);
nor U8268 (N_8268,N_5556,N_4502);
nor U8269 (N_8269,N_5938,N_1196);
nor U8270 (N_8270,N_5255,N_3595);
nor U8271 (N_8271,N_3841,N_3656);
or U8272 (N_8272,N_2809,N_3602);
xor U8273 (N_8273,N_5377,N_3763);
xor U8274 (N_8274,N_227,N_106);
xor U8275 (N_8275,N_581,N_3178);
nand U8276 (N_8276,N_3487,N_4551);
and U8277 (N_8277,N_3510,N_1116);
nand U8278 (N_8278,N_2780,N_5278);
or U8279 (N_8279,N_2503,N_1515);
or U8280 (N_8280,N_1211,N_5204);
or U8281 (N_8281,N_2977,N_2953);
nand U8282 (N_8282,N_996,N_3159);
and U8283 (N_8283,N_352,N_2963);
and U8284 (N_8284,N_54,N_1821);
and U8285 (N_8285,N_4168,N_3563);
and U8286 (N_8286,N_1382,N_3930);
xnor U8287 (N_8287,N_3180,N_1348);
or U8288 (N_8288,N_4884,N_4709);
nor U8289 (N_8289,N_4666,N_3655);
nand U8290 (N_8290,N_1988,N_2515);
or U8291 (N_8291,N_3897,N_5945);
nand U8292 (N_8292,N_237,N_5145);
nor U8293 (N_8293,N_5811,N_4713);
nor U8294 (N_8294,N_2154,N_5903);
or U8295 (N_8295,N_5456,N_3735);
and U8296 (N_8296,N_2159,N_1004);
nand U8297 (N_8297,N_3580,N_3141);
nor U8298 (N_8298,N_4165,N_2791);
or U8299 (N_8299,N_700,N_1642);
or U8300 (N_8300,N_3466,N_1409);
and U8301 (N_8301,N_138,N_1930);
nor U8302 (N_8302,N_2116,N_3074);
nor U8303 (N_8303,N_3788,N_5346);
nor U8304 (N_8304,N_3918,N_2003);
or U8305 (N_8305,N_344,N_5347);
xor U8306 (N_8306,N_1547,N_5325);
or U8307 (N_8307,N_4560,N_4220);
and U8308 (N_8308,N_977,N_1952);
and U8309 (N_8309,N_4187,N_1074);
nand U8310 (N_8310,N_4372,N_2661);
and U8311 (N_8311,N_5622,N_3718);
nor U8312 (N_8312,N_3654,N_3865);
or U8313 (N_8313,N_1855,N_78);
nor U8314 (N_8314,N_1240,N_5882);
nor U8315 (N_8315,N_3681,N_2081);
and U8316 (N_8316,N_2884,N_4699);
and U8317 (N_8317,N_1014,N_4758);
or U8318 (N_8318,N_2122,N_3032);
nand U8319 (N_8319,N_5990,N_3826);
nand U8320 (N_8320,N_3704,N_3511);
and U8321 (N_8321,N_2832,N_4813);
and U8322 (N_8322,N_3911,N_3005);
nor U8323 (N_8323,N_3711,N_5296);
nand U8324 (N_8324,N_2665,N_307);
nand U8325 (N_8325,N_1418,N_5910);
nand U8326 (N_8326,N_1177,N_1554);
nor U8327 (N_8327,N_4389,N_5051);
or U8328 (N_8328,N_3994,N_5963);
and U8329 (N_8329,N_2972,N_3000);
nand U8330 (N_8330,N_1298,N_2422);
xnor U8331 (N_8331,N_5764,N_4283);
nor U8332 (N_8332,N_4838,N_1975);
nand U8333 (N_8333,N_2917,N_2258);
xnor U8334 (N_8334,N_3028,N_302);
nand U8335 (N_8335,N_3098,N_286);
xnor U8336 (N_8336,N_5162,N_1290);
nand U8337 (N_8337,N_765,N_2677);
nand U8338 (N_8338,N_614,N_1856);
xnor U8339 (N_8339,N_4548,N_568);
nand U8340 (N_8340,N_1811,N_593);
nor U8341 (N_8341,N_4348,N_4093);
nor U8342 (N_8342,N_1457,N_3912);
nand U8343 (N_8343,N_2703,N_2527);
and U8344 (N_8344,N_1606,N_1349);
xnor U8345 (N_8345,N_4920,N_1608);
xor U8346 (N_8346,N_640,N_2652);
nand U8347 (N_8347,N_5192,N_1325);
nor U8348 (N_8348,N_785,N_73);
xnor U8349 (N_8349,N_4764,N_101);
nor U8350 (N_8350,N_2408,N_4335);
or U8351 (N_8351,N_5827,N_5039);
xor U8352 (N_8352,N_372,N_4908);
nor U8353 (N_8353,N_2079,N_3621);
nand U8354 (N_8354,N_4226,N_3847);
or U8355 (N_8355,N_766,N_1033);
nand U8356 (N_8356,N_3544,N_2057);
nor U8357 (N_8357,N_4186,N_3055);
and U8358 (N_8358,N_2084,N_399);
or U8359 (N_8359,N_4997,N_3539);
or U8360 (N_8360,N_4026,N_490);
nand U8361 (N_8361,N_1438,N_234);
nor U8362 (N_8362,N_4765,N_1640);
nor U8363 (N_8363,N_1535,N_2858);
nor U8364 (N_8364,N_1822,N_4160);
nand U8365 (N_8365,N_3142,N_3951);
nand U8366 (N_8366,N_4058,N_4536);
and U8367 (N_8367,N_1851,N_2595);
and U8368 (N_8368,N_3616,N_2710);
xor U8369 (N_8369,N_1965,N_5637);
nor U8370 (N_8370,N_5752,N_843);
or U8371 (N_8371,N_5486,N_4198);
and U8372 (N_8372,N_2501,N_3103);
nor U8373 (N_8373,N_310,N_5205);
nor U8374 (N_8374,N_2406,N_1463);
and U8375 (N_8375,N_198,N_4710);
and U8376 (N_8376,N_1366,N_4380);
xnor U8377 (N_8377,N_5451,N_2586);
or U8378 (N_8378,N_5390,N_1434);
and U8379 (N_8379,N_4345,N_2700);
nor U8380 (N_8380,N_4325,N_3741);
xnor U8381 (N_8381,N_3016,N_4927);
nand U8382 (N_8382,N_1036,N_655);
or U8383 (N_8383,N_2339,N_3375);
or U8384 (N_8384,N_981,N_4559);
or U8385 (N_8385,N_161,N_4827);
nor U8386 (N_8386,N_342,N_441);
nor U8387 (N_8387,N_1408,N_5713);
and U8388 (N_8388,N_4871,N_2570);
nand U8389 (N_8389,N_1295,N_2845);
nand U8390 (N_8390,N_2801,N_5174);
and U8391 (N_8391,N_3006,N_3033);
or U8392 (N_8392,N_1421,N_5031);
and U8393 (N_8393,N_4017,N_5476);
nand U8394 (N_8394,N_4645,N_656);
or U8395 (N_8395,N_4367,N_2140);
or U8396 (N_8396,N_1696,N_1813);
xor U8397 (N_8397,N_5361,N_3386);
or U8398 (N_8398,N_1082,N_3362);
nor U8399 (N_8399,N_5471,N_2338);
xnor U8400 (N_8400,N_3807,N_645);
nor U8401 (N_8401,N_1253,N_5675);
nand U8402 (N_8402,N_3760,N_1140);
and U8403 (N_8403,N_174,N_5733);
xor U8404 (N_8404,N_2553,N_5522);
nor U8405 (N_8405,N_4415,N_4227);
nand U8406 (N_8406,N_1225,N_3693);
nand U8407 (N_8407,N_5732,N_5019);
nor U8408 (N_8408,N_4561,N_2765);
nand U8409 (N_8409,N_804,N_398);
and U8410 (N_8410,N_5489,N_3235);
or U8411 (N_8411,N_2483,N_3503);
and U8412 (N_8412,N_3676,N_143);
or U8413 (N_8413,N_5054,N_617);
and U8414 (N_8414,N_2993,N_4935);
nand U8415 (N_8415,N_719,N_1328);
nand U8416 (N_8416,N_5561,N_3889);
nor U8417 (N_8417,N_5062,N_3799);
or U8418 (N_8418,N_632,N_4203);
or U8419 (N_8419,N_5236,N_4250);
or U8420 (N_8420,N_1431,N_1201);
nand U8421 (N_8421,N_5691,N_4678);
and U8422 (N_8422,N_1424,N_3106);
nor U8423 (N_8423,N_2914,N_1144);
nand U8424 (N_8424,N_5083,N_759);
and U8425 (N_8425,N_2175,N_3084);
and U8426 (N_8426,N_3670,N_3857);
xnor U8427 (N_8427,N_1791,N_2249);
and U8428 (N_8428,N_4945,N_2804);
nand U8429 (N_8429,N_4812,N_1372);
nand U8430 (N_8430,N_317,N_26);
xor U8431 (N_8431,N_2383,N_2123);
nor U8432 (N_8432,N_4894,N_4449);
nor U8433 (N_8433,N_2334,N_3012);
xor U8434 (N_8434,N_1964,N_1130);
and U8435 (N_8435,N_3661,N_3298);
xor U8436 (N_8436,N_2687,N_2013);
or U8437 (N_8437,N_3851,N_5256);
nand U8438 (N_8438,N_504,N_3488);
and U8439 (N_8439,N_1699,N_934);
nor U8440 (N_8440,N_5964,N_5748);
xor U8441 (N_8441,N_2436,N_4828);
nand U8442 (N_8442,N_43,N_4503);
xor U8443 (N_8443,N_2435,N_1688);
and U8444 (N_8444,N_1049,N_2662);
xnor U8445 (N_8445,N_3082,N_4263);
nand U8446 (N_8446,N_4327,N_814);
nor U8447 (N_8447,N_5592,N_5473);
nand U8448 (N_8448,N_1441,N_4064);
or U8449 (N_8449,N_4018,N_1230);
xnor U8450 (N_8450,N_204,N_400);
nor U8451 (N_8451,N_4982,N_5498);
and U8452 (N_8452,N_3172,N_1085);
or U8453 (N_8453,N_1114,N_2209);
nor U8454 (N_8454,N_2465,N_3629);
nand U8455 (N_8455,N_5289,N_159);
nor U8456 (N_8456,N_2196,N_5862);
nor U8457 (N_8457,N_4672,N_4103);
and U8458 (N_8458,N_2574,N_868);
nand U8459 (N_8459,N_2940,N_1571);
xnor U8460 (N_8460,N_4983,N_1134);
xor U8461 (N_8461,N_4647,N_4068);
nor U8462 (N_8462,N_3228,N_2976);
or U8463 (N_8463,N_1442,N_5297);
and U8464 (N_8464,N_1350,N_840);
and U8465 (N_8465,N_4090,N_5968);
and U8466 (N_8466,N_2325,N_2402);
and U8467 (N_8467,N_2070,N_4680);
nand U8468 (N_8468,N_99,N_3281);
nand U8469 (N_8469,N_1282,N_697);
or U8470 (N_8470,N_5761,N_296);
nand U8471 (N_8471,N_3829,N_1659);
and U8472 (N_8472,N_429,N_5093);
nor U8473 (N_8473,N_1783,N_817);
and U8474 (N_8474,N_1687,N_1868);
or U8475 (N_8475,N_5776,N_1916);
nand U8476 (N_8476,N_1708,N_4486);
and U8477 (N_8477,N_3429,N_5545);
and U8478 (N_8478,N_1410,N_148);
and U8479 (N_8479,N_2731,N_3301);
xnor U8480 (N_8480,N_2633,N_247);
or U8481 (N_8481,N_1537,N_2594);
and U8482 (N_8482,N_5270,N_1871);
or U8483 (N_8483,N_584,N_659);
xnor U8484 (N_8484,N_3530,N_4648);
nor U8485 (N_8485,N_305,N_2734);
and U8486 (N_8486,N_4631,N_1939);
nor U8487 (N_8487,N_89,N_2949);
and U8488 (N_8488,N_906,N_2713);
nor U8489 (N_8489,N_1581,N_4482);
nor U8490 (N_8490,N_5082,N_1054);
and U8491 (N_8491,N_5512,N_160);
xnor U8492 (N_8492,N_2415,N_1730);
and U8493 (N_8493,N_2985,N_828);
nor U8494 (N_8494,N_5701,N_4623);
nor U8495 (N_8495,N_1459,N_4460);
xnor U8496 (N_8496,N_3342,N_4464);
nand U8497 (N_8497,N_5619,N_5478);
nand U8498 (N_8498,N_880,N_2749);
or U8499 (N_8499,N_1521,N_1065);
or U8500 (N_8500,N_5074,N_2545);
nor U8501 (N_8501,N_997,N_5186);
nand U8502 (N_8502,N_1473,N_5867);
or U8503 (N_8503,N_3730,N_1737);
xor U8504 (N_8504,N_290,N_5360);
nand U8505 (N_8505,N_2307,N_586);
nand U8506 (N_8506,N_4730,N_370);
xor U8507 (N_8507,N_4417,N_5598);
nand U8508 (N_8508,N_2195,N_2404);
nor U8509 (N_8509,N_4404,N_5870);
nor U8510 (N_8510,N_3058,N_1309);
and U8511 (N_8511,N_4484,N_1003);
and U8512 (N_8512,N_4507,N_611);
nand U8513 (N_8513,N_5343,N_2130);
nand U8514 (N_8514,N_2488,N_4045);
or U8515 (N_8515,N_1192,N_1451);
nor U8516 (N_8516,N_2233,N_340);
and U8517 (N_8517,N_1101,N_2730);
and U8518 (N_8518,N_951,N_413);
and U8519 (N_8519,N_852,N_3343);
and U8520 (N_8520,N_3608,N_1966);
or U8521 (N_8521,N_1748,N_4887);
nand U8522 (N_8522,N_5932,N_236);
nor U8523 (N_8523,N_5113,N_5250);
xor U8524 (N_8524,N_5608,N_3624);
and U8525 (N_8525,N_246,N_894);
nor U8526 (N_8526,N_1758,N_4749);
and U8527 (N_8527,N_3574,N_999);
or U8528 (N_8528,N_3147,N_574);
and U8529 (N_8529,N_5797,N_2495);
or U8530 (N_8530,N_1862,N_1840);
or U8531 (N_8531,N_2990,N_931);
or U8532 (N_8532,N_2910,N_743);
nor U8533 (N_8533,N_2578,N_2047);
and U8534 (N_8534,N_2077,N_4701);
or U8535 (N_8535,N_599,N_3811);
nor U8536 (N_8536,N_896,N_3917);
nor U8537 (N_8537,N_5418,N_4614);
nand U8538 (N_8538,N_5355,N_2523);
nand U8539 (N_8539,N_4193,N_1820);
or U8540 (N_8540,N_1482,N_4580);
or U8541 (N_8541,N_4057,N_2295);
nor U8542 (N_8542,N_728,N_5225);
and U8543 (N_8543,N_3446,N_5509);
or U8544 (N_8544,N_3383,N_5196);
nand U8545 (N_8545,N_2302,N_1373);
or U8546 (N_8546,N_3207,N_2433);
nand U8547 (N_8547,N_254,N_383);
or U8548 (N_8548,N_1757,N_5600);
xnor U8549 (N_8549,N_3992,N_4981);
and U8550 (N_8550,N_1050,N_5110);
xnor U8551 (N_8551,N_1960,N_2358);
or U8552 (N_8552,N_1804,N_3031);
nor U8553 (N_8553,N_3294,N_4912);
nand U8554 (N_8554,N_1057,N_1831);
and U8555 (N_8555,N_5085,N_3523);
and U8556 (N_8556,N_3403,N_3900);
nor U8557 (N_8557,N_5842,N_3549);
and U8558 (N_8558,N_966,N_5890);
nor U8559 (N_8559,N_5666,N_612);
and U8560 (N_8560,N_2512,N_4904);
and U8561 (N_8561,N_3650,N_2635);
and U8562 (N_8562,N_3908,N_3535);
or U8563 (N_8563,N_1882,N_1506);
and U8564 (N_8564,N_4564,N_3105);
nand U8565 (N_8565,N_598,N_5590);
nor U8566 (N_8566,N_2612,N_5281);
or U8567 (N_8567,N_1866,N_5511);
nand U8568 (N_8568,N_4797,N_2642);
or U8569 (N_8569,N_20,N_2056);
nor U8570 (N_8570,N_2051,N_3091);
and U8571 (N_8571,N_1265,N_1055);
or U8572 (N_8572,N_786,N_4004);
or U8573 (N_8573,N_5337,N_5794);
or U8574 (N_8574,N_1436,N_1316);
nor U8575 (N_8575,N_3497,N_603);
nand U8576 (N_8576,N_1793,N_4265);
or U8577 (N_8577,N_1153,N_741);
and U8578 (N_8578,N_1842,N_3206);
or U8579 (N_8579,N_2082,N_1732);
and U8580 (N_8580,N_3538,N_5328);
nand U8581 (N_8581,N_1248,N_4909);
and U8582 (N_8582,N_5850,N_1278);
nand U8583 (N_8583,N_3250,N_2932);
and U8584 (N_8584,N_3666,N_2627);
or U8585 (N_8585,N_3678,N_2835);
or U8586 (N_8586,N_5454,N_4748);
or U8587 (N_8587,N_5887,N_2452);
nand U8588 (N_8588,N_2840,N_874);
or U8589 (N_8589,N_1982,N_346);
xnor U8590 (N_8590,N_4301,N_4286);
and U8591 (N_8591,N_215,N_5067);
or U8592 (N_8592,N_5272,N_5506);
nor U8593 (N_8593,N_1119,N_1928);
or U8594 (N_8594,N_3065,N_4135);
nor U8595 (N_8595,N_5378,N_2516);
nor U8596 (N_8596,N_5586,N_4371);
nand U8597 (N_8597,N_4260,N_3256);
or U8598 (N_8598,N_354,N_176);
or U8599 (N_8599,N_2319,N_2242);
xnor U8600 (N_8600,N_3869,N_4479);
or U8601 (N_8601,N_3024,N_4264);
nand U8602 (N_8602,N_2948,N_1494);
or U8603 (N_8603,N_1833,N_2421);
nand U8604 (N_8604,N_3186,N_158);
nand U8605 (N_8605,N_3623,N_726);
xor U8606 (N_8606,N_5242,N_485);
or U8607 (N_8607,N_5258,N_3448);
nand U8608 (N_8608,N_1716,N_2525);
nand U8609 (N_8609,N_2093,N_5504);
xor U8610 (N_8610,N_5122,N_1902);
nand U8611 (N_8611,N_4553,N_1241);
and U8612 (N_8612,N_2692,N_3927);
and U8613 (N_8613,N_2217,N_1912);
or U8614 (N_8614,N_1720,N_1727);
and U8615 (N_8615,N_720,N_1986);
nor U8616 (N_8616,N_4533,N_2833);
xor U8617 (N_8617,N_5629,N_2179);
nor U8618 (N_8618,N_1890,N_1934);
nand U8619 (N_8619,N_5520,N_5952);
or U8620 (N_8620,N_3808,N_1106);
or U8621 (N_8621,N_3973,N_5027);
nand U8622 (N_8622,N_5755,N_4183);
nor U8623 (N_8623,N_3518,N_2311);
and U8624 (N_8624,N_2622,N_2647);
and U8625 (N_8625,N_2166,N_4142);
and U8626 (N_8626,N_320,N_905);
and U8627 (N_8627,N_3227,N_4129);
and U8628 (N_8628,N_1674,N_4880);
or U8629 (N_8629,N_1062,N_4947);
nand U8630 (N_8630,N_3536,N_2487);
xor U8631 (N_8631,N_5496,N_5678);
nand U8632 (N_8632,N_1903,N_1562);
or U8633 (N_8633,N_1766,N_4315);
or U8634 (N_8634,N_5076,N_1090);
xor U8635 (N_8635,N_1151,N_5220);
and U8636 (N_8636,N_5484,N_2950);
and U8637 (N_8637,N_2160,N_363);
or U8638 (N_8638,N_1312,N_948);
or U8639 (N_8639,N_514,N_5277);
nand U8640 (N_8640,N_780,N_3700);
xor U8641 (N_8641,N_2771,N_2551);
and U8642 (N_8642,N_5465,N_5714);
xnor U8643 (N_8643,N_518,N_5201);
or U8644 (N_8644,N_3045,N_2032);
xnor U8645 (N_8645,N_4197,N_4084);
and U8646 (N_8646,N_3208,N_1505);
nor U8647 (N_8647,N_1572,N_746);
nor U8648 (N_8648,N_1900,N_4181);
nor U8649 (N_8649,N_4478,N_3680);
xor U8650 (N_8650,N_361,N_2468);
or U8651 (N_8651,N_5168,N_3515);
and U8652 (N_8652,N_4115,N_2773);
nor U8653 (N_8653,N_5889,N_1462);
and U8654 (N_8654,N_4540,N_5380);
nand U8655 (N_8655,N_527,N_2965);
xnor U8656 (N_8656,N_11,N_5925);
nor U8657 (N_8657,N_5017,N_916);
nand U8658 (N_8658,N_5580,N_3360);
nand U8659 (N_8659,N_4185,N_3778);
nor U8660 (N_8660,N_3330,N_3170);
xnor U8661 (N_8661,N_4642,N_4230);
or U8662 (N_8662,N_3423,N_2782);
or U8663 (N_8663,N_5215,N_2781);
and U8664 (N_8664,N_5671,N_2678);
or U8665 (N_8665,N_3742,N_36);
and U8666 (N_8666,N_3273,N_238);
nand U8667 (N_8667,N_4943,N_4541);
or U8668 (N_8668,N_2583,N_5047);
xor U8669 (N_8669,N_3328,N_5680);
or U8670 (N_8670,N_5131,N_5861);
nor U8671 (N_8671,N_181,N_2941);
nor U8672 (N_8672,N_1478,N_3861);
nor U8673 (N_8673,N_1008,N_4571);
xor U8674 (N_8674,N_4477,N_4381);
and U8675 (N_8675,N_1734,N_2786);
xor U8676 (N_8676,N_1174,N_641);
and U8677 (N_8677,N_3609,N_3489);
nand U8678 (N_8678,N_2472,N_5446);
and U8679 (N_8679,N_5612,N_2381);
nor U8680 (N_8680,N_5485,N_3551);
or U8681 (N_8681,N_5447,N_5758);
nor U8682 (N_8682,N_5676,N_5955);
nand U8683 (N_8683,N_3651,N_4537);
nand U8684 (N_8684,N_2784,N_4091);
or U8685 (N_8685,N_233,N_5326);
and U8686 (N_8686,N_4783,N_1962);
and U8687 (N_8687,N_3436,N_4598);
nor U8688 (N_8688,N_376,N_824);
xor U8689 (N_8689,N_5711,N_4492);
nand U8690 (N_8690,N_222,N_2236);
nand U8691 (N_8691,N_589,N_2235);
nor U8692 (N_8692,N_345,N_287);
and U8693 (N_8693,N_5519,N_5846);
or U8694 (N_8694,N_4216,N_1244);
nor U8695 (N_8695,N_1974,N_1178);
nand U8696 (N_8696,N_4159,N_1969);
xor U8697 (N_8697,N_660,N_3880);
or U8698 (N_8698,N_2088,N_2419);
nand U8699 (N_8699,N_3020,N_909);
or U8700 (N_8700,N_4557,N_2810);
nor U8701 (N_8701,N_4281,N_658);
or U8702 (N_8702,N_3121,N_1075);
nor U8703 (N_8703,N_4037,N_2239);
or U8704 (N_8704,N_2046,N_47);
nand U8705 (N_8705,N_4596,N_417);
nor U8706 (N_8706,N_5115,N_4901);
nor U8707 (N_8707,N_5954,N_993);
or U8708 (N_8708,N_3364,N_4771);
and U8709 (N_8709,N_4669,N_4550);
nor U8710 (N_8710,N_2873,N_4365);
nor U8711 (N_8711,N_502,N_4594);
or U8712 (N_8712,N_1258,N_2793);
xor U8713 (N_8713,N_3067,N_5488);
nor U8714 (N_8714,N_5049,N_3266);
and U8715 (N_8715,N_1135,N_4396);
nor U8716 (N_8716,N_4086,N_4490);
nor U8717 (N_8717,N_1179,N_5395);
nand U8718 (N_8718,N_155,N_5021);
nand U8719 (N_8719,N_5218,N_5723);
and U8720 (N_8720,N_5003,N_405);
and U8721 (N_8721,N_484,N_3345);
nand U8722 (N_8722,N_2569,N_5745);
nand U8723 (N_8723,N_4938,N_3312);
and U8724 (N_8724,N_3213,N_512);
or U8725 (N_8725,N_5940,N_2268);
xnor U8726 (N_8726,N_3753,N_5212);
nor U8727 (N_8727,N_2546,N_818);
nand U8728 (N_8728,N_3331,N_5883);
xnor U8729 (N_8729,N_5757,N_477);
nor U8730 (N_8730,N_1060,N_3299);
nand U8731 (N_8731,N_4975,N_3161);
and U8732 (N_8732,N_3702,N_3066);
xnor U8733 (N_8733,N_2720,N_1190);
nand U8734 (N_8734,N_3576,N_4271);
xor U8735 (N_8735,N_1913,N_392);
nand U8736 (N_8736,N_5371,N_1739);
nand U8737 (N_8737,N_721,N_1746);
nor U8738 (N_8738,N_2706,N_4587);
nor U8739 (N_8739,N_1470,N_2714);
nand U8740 (N_8740,N_1514,N_4667);
nor U8741 (N_8741,N_3316,N_4175);
or U8742 (N_8742,N_2042,N_5452);
nor U8743 (N_8743,N_5611,N_2328);
xor U8744 (N_8744,N_437,N_85);
nor U8745 (N_8745,N_4567,N_5026);
and U8746 (N_8746,N_1266,N_4102);
nor U8747 (N_8747,N_4872,N_4840);
nand U8748 (N_8748,N_2777,N_1743);
and U8749 (N_8749,N_5791,N_2340);
xor U8750 (N_8750,N_4358,N_2846);
or U8751 (N_8751,N_4481,N_3287);
or U8752 (N_8752,N_2190,N_732);
xnor U8753 (N_8753,N_491,N_723);
or U8754 (N_8754,N_2763,N_3789);
or U8755 (N_8755,N_4608,N_3474);
nand U8756 (N_8756,N_4189,N_2103);
nand U8757 (N_8757,N_5602,N_1204);
nand U8758 (N_8758,N_5077,N_4318);
or U8759 (N_8759,N_84,N_190);
nor U8760 (N_8760,N_2297,N_5542);
nor U8761 (N_8761,N_2060,N_5257);
nand U8762 (N_8762,N_1615,N_520);
xor U8763 (N_8763,N_1389,N_609);
and U8764 (N_8764,N_2795,N_3174);
and U8765 (N_8765,N_3728,N_57);
nand U8766 (N_8766,N_2485,N_1071);
and U8767 (N_8767,N_5173,N_5327);
and U8768 (N_8768,N_2012,N_3245);
xnor U8769 (N_8769,N_5759,N_2955);
nand U8770 (N_8770,N_4322,N_4547);
xnor U8771 (N_8771,N_4147,N_5866);
nor U8772 (N_8772,N_1738,N_3823);
or U8773 (N_8773,N_1354,N_65);
nand U8774 (N_8774,N_4597,N_2962);
and U8775 (N_8775,N_3588,N_4708);
nor U8776 (N_8776,N_3901,N_5241);
and U8777 (N_8777,N_4752,N_3820);
nand U8778 (N_8778,N_1016,N_4088);
nand U8779 (N_8779,N_5716,N_903);
and U8780 (N_8780,N_200,N_2524);
nor U8781 (N_8781,N_5125,N_3818);
nor U8782 (N_8782,N_727,N_4360);
nand U8783 (N_8783,N_5531,N_4116);
nor U8784 (N_8784,N_4676,N_4060);
xnor U8785 (N_8785,N_379,N_4831);
nand U8786 (N_8786,N_2429,N_2792);
xnor U8787 (N_8787,N_2946,N_5358);
nand U8788 (N_8788,N_294,N_5780);
and U8789 (N_8789,N_5896,N_742);
or U8790 (N_8790,N_5792,N_1847);
or U8791 (N_8791,N_4108,N_4737);
or U8792 (N_8792,N_5670,N_1234);
and U8793 (N_8793,N_958,N_218);
and U8794 (N_8794,N_5291,N_4044);
xor U8795 (N_8795,N_3849,N_5391);
and U8796 (N_8796,N_4585,N_5330);
nand U8797 (N_8797,N_4714,N_1784);
and U8798 (N_8798,N_4120,N_4677);
and U8799 (N_8799,N_3393,N_63);
nor U8800 (N_8800,N_5525,N_1400);
nor U8801 (N_8801,N_3284,N_1411);
xnor U8802 (N_8802,N_2968,N_3975);
nand U8803 (N_8803,N_2119,N_3465);
and U8804 (N_8804,N_3196,N_3223);
nor U8805 (N_8805,N_5552,N_3425);
nor U8806 (N_8806,N_5880,N_5178);
or U8807 (N_8807,N_142,N_4452);
nand U8808 (N_8808,N_2477,N_2384);
and U8809 (N_8809,N_369,N_5057);
and U8810 (N_8810,N_289,N_5407);
and U8811 (N_8811,N_976,N_591);
nand U8812 (N_8812,N_2535,N_5962);
or U8813 (N_8813,N_5433,N_1168);
or U8814 (N_8814,N_3980,N_4050);
nor U8815 (N_8815,N_2557,N_4987);
and U8816 (N_8816,N_4640,N_3985);
or U8817 (N_8817,N_228,N_3710);
nand U8818 (N_8818,N_2029,N_5623);
or U8819 (N_8819,N_4411,N_2698);
and U8820 (N_8820,N_3529,N_3606);
nand U8821 (N_8821,N_5787,N_378);
or U8822 (N_8822,N_4609,N_3405);
and U8823 (N_8823,N_3812,N_4670);
xnor U8824 (N_8824,N_646,N_627);
nand U8825 (N_8825,N_3046,N_4298);
and U8826 (N_8826,N_754,N_1159);
or U8827 (N_8827,N_5441,N_1358);
nand U8828 (N_8828,N_5749,N_80);
and U8829 (N_8829,N_102,N_1574);
or U8830 (N_8830,N_5136,N_2294);
nand U8831 (N_8831,N_2086,N_1972);
nand U8832 (N_8832,N_3092,N_5843);
or U8833 (N_8833,N_3200,N_4684);
or U8834 (N_8834,N_838,N_122);
or U8835 (N_8835,N_3099,N_3451);
and U8836 (N_8836,N_420,N_2347);
or U8837 (N_8837,N_5959,N_972);
nor U8838 (N_8838,N_4588,N_4329);
xnor U8839 (N_8839,N_2245,N_4743);
or U8840 (N_8840,N_394,N_4837);
or U8841 (N_8841,N_5547,N_1667);
or U8842 (N_8842,N_2767,N_278);
and U8843 (N_8843,N_1063,N_5865);
nand U8844 (N_8844,N_4253,N_1824);
or U8845 (N_8845,N_5404,N_4416);
or U8846 (N_8846,N_488,N_1759);
nor U8847 (N_8847,N_2520,N_4003);
xor U8848 (N_8848,N_1585,N_1167);
xor U8849 (N_8849,N_540,N_5299);
and U8850 (N_8850,N_4963,N_5928);
nor U8851 (N_8851,N_3931,N_5211);
and U8852 (N_8852,N_1752,N_4968);
nor U8853 (N_8853,N_3125,N_322);
or U8854 (N_8854,N_5569,N_1812);
nand U8855 (N_8855,N_4229,N_2926);
nor U8856 (N_8856,N_4351,N_2061);
or U8857 (N_8857,N_2679,N_5516);
xnor U8858 (N_8858,N_2455,N_5537);
nor U8859 (N_8859,N_2355,N_808);
and U8860 (N_8860,N_729,N_5419);
and U8861 (N_8861,N_1967,N_1184);
or U8862 (N_8862,N_4685,N_5221);
nor U8863 (N_8863,N_932,N_3140);
and U8864 (N_8864,N_1907,N_5993);
and U8865 (N_8865,N_4382,N_4423);
nor U8866 (N_8866,N_5388,N_3952);
and U8867 (N_8867,N_5102,N_1215);
nor U8868 (N_8868,N_2689,N_3455);
xnor U8869 (N_8869,N_2102,N_5981);
or U8870 (N_8870,N_4013,N_2018);
and U8871 (N_8871,N_2,N_806);
and U8872 (N_8872,N_2729,N_3162);
nand U8873 (N_8873,N_3777,N_1676);
or U8874 (N_8874,N_5536,N_2424);
or U8875 (N_8875,N_772,N_4582);
nand U8876 (N_8876,N_1394,N_779);
xor U8877 (N_8877,N_4,N_5521);
nor U8878 (N_8878,N_1483,N_1880);
or U8879 (N_8879,N_816,N_4366);
xor U8880 (N_8880,N_82,N_608);
nor U8881 (N_8881,N_541,N_171);
or U8882 (N_8882,N_5375,N_1576);
and U8883 (N_8883,N_4505,N_4961);
nor U8884 (N_8884,N_5413,N_5899);
nand U8885 (N_8885,N_5663,N_3837);
or U8886 (N_8886,N_3708,N_4210);
nand U8887 (N_8887,N_3568,N_5517);
and U8888 (N_8888,N_5239,N_100);
xor U8889 (N_8889,N_5222,N_3246);
nand U8890 (N_8890,N_3867,N_1703);
and U8891 (N_8891,N_1456,N_1714);
nor U8892 (N_8892,N_3787,N_4431);
or U8893 (N_8893,N_1569,N_1507);
nand U8894 (N_8894,N_232,N_3138);
nor U8895 (N_8895,N_4109,N_3824);
nand U8896 (N_8896,N_4516,N_5176);
nor U8897 (N_8897,N_649,N_3528);
or U8898 (N_8898,N_652,N_4386);
and U8899 (N_8899,N_3699,N_3526);
nand U8900 (N_8900,N_4722,N_3073);
nor U8901 (N_8901,N_961,N_2748);
nor U8902 (N_8902,N_4468,N_5499);
or U8903 (N_8903,N_674,N_210);
nor U8904 (N_8904,N_1432,N_3305);
nor U8905 (N_8905,N_3795,N_2739);
nand U8906 (N_8906,N_625,N_1744);
or U8907 (N_8907,N_1555,N_4986);
nand U8908 (N_8908,N_4042,N_2074);
xor U8909 (N_8909,N_897,N_1445);
or U8910 (N_8910,N_1430,N_767);
and U8911 (N_8911,N_3573,N_4130);
nand U8912 (N_8912,N_4256,N_1989);
and U8913 (N_8913,N_5503,N_1447);
nor U8914 (N_8914,N_3717,N_2323);
nand U8915 (N_8915,N_5514,N_3181);
or U8916 (N_8916,N_3486,N_978);
nor U8917 (N_8917,N_750,N_5495);
nor U8918 (N_8918,N_5841,N_942);
and U8919 (N_8919,N_2280,N_1331);
or U8920 (N_8920,N_1614,N_3942);
nand U8921 (N_8921,N_4895,N_4346);
xnor U8922 (N_8922,N_5721,N_5124);
nor U8923 (N_8923,N_5363,N_3794);
xor U8924 (N_8924,N_3278,N_5223);
nor U8925 (N_8925,N_1186,N_856);
xnor U8926 (N_8926,N_1122,N_2128);
nand U8927 (N_8927,N_3637,N_486);
nor U8928 (N_8928,N_4236,N_495);
or U8929 (N_8929,N_1911,N_3738);
nand U8930 (N_8930,N_5996,N_5235);
nand U8931 (N_8931,N_5808,N_4157);
and U8932 (N_8932,N_4595,N_4869);
nand U8933 (N_8933,N_1264,N_2837);
or U8934 (N_8934,N_1942,N_4805);
nand U8935 (N_8935,N_2055,N_3111);
or U8936 (N_8936,N_5686,N_5871);
and U8937 (N_8937,N_1105,N_4290);
xnor U8938 (N_8938,N_2613,N_1826);
nand U8939 (N_8939,N_5458,N_4796);
nor U8940 (N_8940,N_5231,N_3346);
or U8941 (N_8941,N_778,N_4127);
nand U8942 (N_8942,N_1002,N_4865);
and U8943 (N_8943,N_5279,N_258);
or U8944 (N_8944,N_3645,N_2959);
and U8945 (N_8945,N_4725,N_854);
or U8946 (N_8946,N_1545,N_5901);
nor U8947 (N_8947,N_5163,N_2971);
nor U8948 (N_8948,N_1946,N_2009);
xnor U8949 (N_8949,N_789,N_48);
nand U8950 (N_8950,N_5726,N_5362);
and U8951 (N_8951,N_2410,N_4009);
nand U8952 (N_8952,N_5474,N_4333);
or U8953 (N_8953,N_5820,N_3983);
or U8954 (N_8954,N_1158,N_3182);
nor U8955 (N_8955,N_1334,N_4293);
xnor U8956 (N_8956,N_3620,N_2418);
or U8957 (N_8957,N_2448,N_4435);
and U8958 (N_8958,N_2356,N_4309);
and U8959 (N_8959,N_4848,N_253);
nand U8960 (N_8960,N_3895,N_4809);
nand U8961 (N_8961,N_4357,N_4043);
or U8962 (N_8962,N_5674,N_2283);
or U8963 (N_8963,N_3124,N_5193);
nor U8964 (N_8964,N_1335,N_5037);
nand U8965 (N_8965,N_5695,N_1384);
nand U8966 (N_8966,N_851,N_2827);
xor U8967 (N_8967,N_4495,N_5881);
or U8968 (N_8968,N_4922,N_4605);
or U8969 (N_8969,N_1238,N_5798);
and U8970 (N_8970,N_3475,N_5736);
nand U8971 (N_8971,N_1402,N_4800);
nor U8972 (N_8972,N_1068,N_4705);
or U8973 (N_8973,N_1223,N_4558);
and U8974 (N_8974,N_551,N_5613);
or U8975 (N_8975,N_5189,N_4117);
or U8976 (N_8976,N_3844,N_3630);
nand U8977 (N_8977,N_1450,N_5693);
nand U8978 (N_8978,N_2087,N_5653);
nor U8979 (N_8979,N_3776,N_4047);
and U8980 (N_8980,N_3619,N_2031);
nand U8981 (N_8981,N_5994,N_1502);
and U8982 (N_8982,N_3439,N_265);
nand U8983 (N_8983,N_5659,N_4851);
nand U8984 (N_8984,N_1318,N_573);
and U8985 (N_8985,N_4072,N_1365);
and U8986 (N_8986,N_3153,N_1534);
nor U8987 (N_8987,N_3658,N_2761);
nor U8988 (N_8988,N_474,N_5271);
nor U8989 (N_8989,N_4310,N_2378);
nand U8990 (N_8990,N_2080,N_1901);
nor U8991 (N_8991,N_3285,N_4643);
or U8992 (N_8992,N_4270,N_1239);
or U8993 (N_8993,N_1863,N_4247);
nor U8994 (N_8994,N_5406,N_120);
and U8995 (N_8995,N_2818,N_88);
nor U8996 (N_8996,N_4099,N_266);
nor U8997 (N_8997,N_3771,N_4638);
or U8998 (N_8998,N_4990,N_2658);
nor U8999 (N_8999,N_5249,N_2776);
nand U9000 (N_9000,N_2882,N_755);
or U9001 (N_9001,N_2849,N_3308);
or U9002 (N_9002,N_4596,N_5271);
nand U9003 (N_9003,N_3593,N_1479);
or U9004 (N_9004,N_1871,N_452);
and U9005 (N_9005,N_2959,N_1809);
and U9006 (N_9006,N_3721,N_3328);
xnor U9007 (N_9007,N_235,N_3943);
nor U9008 (N_9008,N_190,N_3346);
nor U9009 (N_9009,N_5587,N_3374);
or U9010 (N_9010,N_5871,N_1317);
nand U9011 (N_9011,N_1412,N_799);
nor U9012 (N_9012,N_2146,N_2050);
xnor U9013 (N_9013,N_3451,N_4403);
nand U9014 (N_9014,N_218,N_2812);
or U9015 (N_9015,N_675,N_3067);
or U9016 (N_9016,N_2285,N_2311);
nor U9017 (N_9017,N_735,N_2403);
or U9018 (N_9018,N_3875,N_636);
and U9019 (N_9019,N_4665,N_2685);
and U9020 (N_9020,N_2892,N_296);
and U9021 (N_9021,N_2429,N_4197);
and U9022 (N_9022,N_4569,N_5532);
and U9023 (N_9023,N_5350,N_201);
nor U9024 (N_9024,N_1004,N_2567);
and U9025 (N_9025,N_3179,N_2244);
and U9026 (N_9026,N_2731,N_5136);
and U9027 (N_9027,N_4794,N_550);
and U9028 (N_9028,N_492,N_1014);
xnor U9029 (N_9029,N_5646,N_2425);
and U9030 (N_9030,N_1895,N_5196);
and U9031 (N_9031,N_17,N_5347);
nand U9032 (N_9032,N_4818,N_1283);
or U9033 (N_9033,N_4396,N_5804);
or U9034 (N_9034,N_2084,N_1313);
nor U9035 (N_9035,N_4240,N_879);
and U9036 (N_9036,N_5739,N_2921);
nand U9037 (N_9037,N_1472,N_4528);
or U9038 (N_9038,N_1833,N_388);
nand U9039 (N_9039,N_1275,N_1291);
nor U9040 (N_9040,N_1795,N_3205);
nor U9041 (N_9041,N_3235,N_5388);
and U9042 (N_9042,N_3515,N_496);
nand U9043 (N_9043,N_1432,N_4125);
nand U9044 (N_9044,N_5262,N_4864);
nor U9045 (N_9045,N_2496,N_3486);
nand U9046 (N_9046,N_1579,N_1587);
or U9047 (N_9047,N_4344,N_2352);
nand U9048 (N_9048,N_4245,N_2563);
and U9049 (N_9049,N_2065,N_3105);
nand U9050 (N_9050,N_381,N_3219);
and U9051 (N_9051,N_4344,N_2052);
or U9052 (N_9052,N_4203,N_2176);
xor U9053 (N_9053,N_4798,N_5045);
and U9054 (N_9054,N_5315,N_2482);
and U9055 (N_9055,N_5095,N_4182);
and U9056 (N_9056,N_4562,N_4627);
xor U9057 (N_9057,N_5570,N_1360);
xor U9058 (N_9058,N_4164,N_4265);
xnor U9059 (N_9059,N_1062,N_3198);
nand U9060 (N_9060,N_0,N_2486);
nor U9061 (N_9061,N_3647,N_2143);
or U9062 (N_9062,N_2403,N_5135);
nand U9063 (N_9063,N_2203,N_5374);
nand U9064 (N_9064,N_1501,N_779);
xor U9065 (N_9065,N_3462,N_4052);
or U9066 (N_9066,N_1556,N_5810);
and U9067 (N_9067,N_2479,N_4026);
or U9068 (N_9068,N_5871,N_4550);
or U9069 (N_9069,N_3225,N_3494);
nor U9070 (N_9070,N_4985,N_2694);
nand U9071 (N_9071,N_5668,N_2776);
or U9072 (N_9072,N_4165,N_1578);
or U9073 (N_9073,N_2351,N_4079);
nor U9074 (N_9074,N_1177,N_606);
nand U9075 (N_9075,N_3657,N_1730);
or U9076 (N_9076,N_239,N_4769);
nand U9077 (N_9077,N_3891,N_358);
and U9078 (N_9078,N_5945,N_505);
nand U9079 (N_9079,N_5690,N_3724);
nor U9080 (N_9080,N_5127,N_3503);
nand U9081 (N_9081,N_5897,N_1400);
or U9082 (N_9082,N_5868,N_921);
or U9083 (N_9083,N_3175,N_1482);
nor U9084 (N_9084,N_5804,N_854);
and U9085 (N_9085,N_5563,N_1341);
xor U9086 (N_9086,N_535,N_3914);
and U9087 (N_9087,N_2039,N_1150);
or U9088 (N_9088,N_5719,N_2995);
xnor U9089 (N_9089,N_1876,N_2229);
nand U9090 (N_9090,N_4842,N_3349);
xor U9091 (N_9091,N_751,N_628);
or U9092 (N_9092,N_4144,N_5967);
or U9093 (N_9093,N_3156,N_69);
or U9094 (N_9094,N_1277,N_852);
or U9095 (N_9095,N_3091,N_3697);
xnor U9096 (N_9096,N_3329,N_2509);
or U9097 (N_9097,N_4387,N_500);
and U9098 (N_9098,N_1135,N_1450);
or U9099 (N_9099,N_3164,N_3200);
or U9100 (N_9100,N_2545,N_4778);
and U9101 (N_9101,N_505,N_138);
or U9102 (N_9102,N_3511,N_4454);
nor U9103 (N_9103,N_5887,N_2937);
nor U9104 (N_9104,N_4615,N_727);
and U9105 (N_9105,N_940,N_5918);
xor U9106 (N_9106,N_3946,N_4173);
or U9107 (N_9107,N_3972,N_1487);
nand U9108 (N_9108,N_1023,N_4600);
nand U9109 (N_9109,N_505,N_4445);
and U9110 (N_9110,N_1647,N_1348);
nand U9111 (N_9111,N_3650,N_879);
or U9112 (N_9112,N_1711,N_2610);
and U9113 (N_9113,N_3144,N_2918);
xor U9114 (N_9114,N_3171,N_1397);
nand U9115 (N_9115,N_807,N_3089);
xor U9116 (N_9116,N_344,N_156);
nor U9117 (N_9117,N_4247,N_4232);
and U9118 (N_9118,N_4328,N_1005);
nand U9119 (N_9119,N_4348,N_59);
nand U9120 (N_9120,N_2643,N_3644);
or U9121 (N_9121,N_3041,N_3236);
nor U9122 (N_9122,N_2435,N_2497);
xnor U9123 (N_9123,N_4769,N_4375);
and U9124 (N_9124,N_4189,N_2948);
nand U9125 (N_9125,N_3563,N_1580);
xnor U9126 (N_9126,N_535,N_3704);
nor U9127 (N_9127,N_2126,N_2216);
xnor U9128 (N_9128,N_681,N_4221);
or U9129 (N_9129,N_127,N_339);
nand U9130 (N_9130,N_4795,N_5280);
nor U9131 (N_9131,N_5055,N_2229);
nand U9132 (N_9132,N_5137,N_2049);
nor U9133 (N_9133,N_2585,N_2403);
nand U9134 (N_9134,N_3374,N_2389);
nand U9135 (N_9135,N_5247,N_4162);
nand U9136 (N_9136,N_3824,N_4783);
nand U9137 (N_9137,N_2850,N_3474);
nor U9138 (N_9138,N_1565,N_4355);
or U9139 (N_9139,N_183,N_4311);
or U9140 (N_9140,N_2027,N_4162);
or U9141 (N_9141,N_1062,N_2119);
and U9142 (N_9142,N_2542,N_1887);
nor U9143 (N_9143,N_3620,N_960);
and U9144 (N_9144,N_405,N_1905);
nor U9145 (N_9145,N_2635,N_4984);
nand U9146 (N_9146,N_5578,N_455);
nor U9147 (N_9147,N_2118,N_673);
nor U9148 (N_9148,N_5251,N_4183);
and U9149 (N_9149,N_2752,N_2686);
or U9150 (N_9150,N_3553,N_2286);
and U9151 (N_9151,N_588,N_3508);
nor U9152 (N_9152,N_1655,N_1529);
and U9153 (N_9153,N_2481,N_2042);
and U9154 (N_9154,N_4833,N_5334);
nor U9155 (N_9155,N_2812,N_112);
nor U9156 (N_9156,N_4107,N_2191);
or U9157 (N_9157,N_879,N_5331);
nor U9158 (N_9158,N_3367,N_5992);
xor U9159 (N_9159,N_2866,N_3113);
nand U9160 (N_9160,N_4514,N_178);
or U9161 (N_9161,N_898,N_5116);
and U9162 (N_9162,N_3798,N_1406);
xnor U9163 (N_9163,N_5781,N_2669);
or U9164 (N_9164,N_2650,N_5015);
and U9165 (N_9165,N_2695,N_2227);
xnor U9166 (N_9166,N_5422,N_3060);
or U9167 (N_9167,N_572,N_1959);
nor U9168 (N_9168,N_232,N_1598);
nand U9169 (N_9169,N_2363,N_4265);
and U9170 (N_9170,N_5040,N_1852);
or U9171 (N_9171,N_3016,N_2449);
nor U9172 (N_9172,N_1453,N_4403);
xor U9173 (N_9173,N_2555,N_1532);
and U9174 (N_9174,N_2330,N_1893);
nor U9175 (N_9175,N_4280,N_702);
xor U9176 (N_9176,N_2012,N_452);
nor U9177 (N_9177,N_3895,N_836);
nand U9178 (N_9178,N_3274,N_5475);
and U9179 (N_9179,N_2567,N_905);
nand U9180 (N_9180,N_2648,N_2919);
and U9181 (N_9181,N_837,N_5408);
nand U9182 (N_9182,N_2547,N_1799);
nor U9183 (N_9183,N_4510,N_2017);
and U9184 (N_9184,N_1511,N_2483);
or U9185 (N_9185,N_3979,N_4627);
or U9186 (N_9186,N_5563,N_1958);
nor U9187 (N_9187,N_2307,N_4932);
or U9188 (N_9188,N_2340,N_5302);
nor U9189 (N_9189,N_3071,N_678);
or U9190 (N_9190,N_1207,N_1021);
and U9191 (N_9191,N_1955,N_1282);
xor U9192 (N_9192,N_2769,N_2779);
and U9193 (N_9193,N_1883,N_4155);
xor U9194 (N_9194,N_1984,N_4820);
nand U9195 (N_9195,N_816,N_2770);
nand U9196 (N_9196,N_1369,N_2526);
and U9197 (N_9197,N_2297,N_1075);
nor U9198 (N_9198,N_3855,N_4644);
and U9199 (N_9199,N_2823,N_4327);
nor U9200 (N_9200,N_4858,N_1485);
nand U9201 (N_9201,N_4060,N_4482);
nand U9202 (N_9202,N_2150,N_3976);
or U9203 (N_9203,N_5130,N_4758);
or U9204 (N_9204,N_1358,N_4926);
nand U9205 (N_9205,N_1565,N_156);
nor U9206 (N_9206,N_2948,N_3817);
or U9207 (N_9207,N_2871,N_2151);
or U9208 (N_9208,N_5786,N_690);
nor U9209 (N_9209,N_5938,N_5907);
nand U9210 (N_9210,N_4872,N_3425);
and U9211 (N_9211,N_1777,N_1413);
and U9212 (N_9212,N_5703,N_3706);
or U9213 (N_9213,N_678,N_739);
nor U9214 (N_9214,N_59,N_4791);
or U9215 (N_9215,N_218,N_2438);
nand U9216 (N_9216,N_5957,N_2009);
nand U9217 (N_9217,N_733,N_2643);
nor U9218 (N_9218,N_2463,N_1399);
xor U9219 (N_9219,N_4769,N_3468);
nand U9220 (N_9220,N_5488,N_3962);
nor U9221 (N_9221,N_968,N_5716);
and U9222 (N_9222,N_2667,N_5565);
nand U9223 (N_9223,N_5034,N_4575);
nand U9224 (N_9224,N_1086,N_4201);
nor U9225 (N_9225,N_3939,N_764);
nor U9226 (N_9226,N_4411,N_1930);
and U9227 (N_9227,N_5568,N_1153);
or U9228 (N_9228,N_4563,N_761);
nand U9229 (N_9229,N_2661,N_1530);
nor U9230 (N_9230,N_2675,N_93);
nand U9231 (N_9231,N_1184,N_1874);
nor U9232 (N_9232,N_4416,N_2438);
nand U9233 (N_9233,N_4694,N_1207);
nor U9234 (N_9234,N_4660,N_5536);
or U9235 (N_9235,N_2763,N_3305);
xnor U9236 (N_9236,N_2814,N_1816);
nor U9237 (N_9237,N_3946,N_5662);
nand U9238 (N_9238,N_2971,N_3239);
xnor U9239 (N_9239,N_4119,N_1353);
xor U9240 (N_9240,N_2110,N_4946);
and U9241 (N_9241,N_2106,N_5157);
or U9242 (N_9242,N_2193,N_2423);
or U9243 (N_9243,N_4053,N_1350);
or U9244 (N_9244,N_1834,N_1525);
nand U9245 (N_9245,N_845,N_1066);
nor U9246 (N_9246,N_1446,N_5868);
nand U9247 (N_9247,N_3571,N_1140);
and U9248 (N_9248,N_3190,N_1719);
nor U9249 (N_9249,N_3077,N_2103);
or U9250 (N_9250,N_5980,N_583);
or U9251 (N_9251,N_5305,N_2138);
xor U9252 (N_9252,N_5083,N_4321);
nand U9253 (N_9253,N_3125,N_2268);
nor U9254 (N_9254,N_2915,N_5751);
nor U9255 (N_9255,N_4488,N_3847);
nand U9256 (N_9256,N_1286,N_3467);
nand U9257 (N_9257,N_5739,N_5688);
nand U9258 (N_9258,N_2842,N_3400);
or U9259 (N_9259,N_2568,N_3268);
nor U9260 (N_9260,N_780,N_1552);
and U9261 (N_9261,N_4259,N_3397);
and U9262 (N_9262,N_248,N_4930);
and U9263 (N_9263,N_4265,N_5498);
or U9264 (N_9264,N_861,N_1950);
or U9265 (N_9265,N_2190,N_670);
nand U9266 (N_9266,N_4084,N_549);
nand U9267 (N_9267,N_2056,N_4591);
nand U9268 (N_9268,N_5918,N_3188);
or U9269 (N_9269,N_1712,N_5987);
nand U9270 (N_9270,N_1820,N_234);
nand U9271 (N_9271,N_4008,N_4193);
nand U9272 (N_9272,N_5906,N_4463);
nor U9273 (N_9273,N_5292,N_4101);
nand U9274 (N_9274,N_2072,N_2370);
or U9275 (N_9275,N_2667,N_5590);
xor U9276 (N_9276,N_167,N_4508);
nor U9277 (N_9277,N_2357,N_2293);
and U9278 (N_9278,N_1330,N_1432);
and U9279 (N_9279,N_427,N_2440);
nor U9280 (N_9280,N_321,N_4543);
nor U9281 (N_9281,N_416,N_1363);
nor U9282 (N_9282,N_3476,N_2546);
or U9283 (N_9283,N_2737,N_3498);
and U9284 (N_9284,N_5010,N_1554);
and U9285 (N_9285,N_380,N_729);
or U9286 (N_9286,N_4915,N_2799);
or U9287 (N_9287,N_234,N_596);
or U9288 (N_9288,N_2021,N_4968);
nor U9289 (N_9289,N_389,N_3985);
nor U9290 (N_9290,N_1715,N_1497);
nor U9291 (N_9291,N_3380,N_3144);
or U9292 (N_9292,N_2930,N_5723);
nor U9293 (N_9293,N_3828,N_3968);
or U9294 (N_9294,N_503,N_301);
nand U9295 (N_9295,N_3303,N_661);
nand U9296 (N_9296,N_3049,N_479);
and U9297 (N_9297,N_3674,N_49);
nand U9298 (N_9298,N_2558,N_2968);
or U9299 (N_9299,N_5683,N_994);
nand U9300 (N_9300,N_1845,N_1756);
or U9301 (N_9301,N_1999,N_3593);
nor U9302 (N_9302,N_1565,N_1452);
xnor U9303 (N_9303,N_1468,N_4248);
or U9304 (N_9304,N_3648,N_4010);
nor U9305 (N_9305,N_5928,N_3738);
or U9306 (N_9306,N_514,N_2336);
nand U9307 (N_9307,N_470,N_2945);
or U9308 (N_9308,N_2728,N_1872);
and U9309 (N_9309,N_3659,N_4713);
or U9310 (N_9310,N_5527,N_5243);
or U9311 (N_9311,N_611,N_5677);
nor U9312 (N_9312,N_4270,N_261);
and U9313 (N_9313,N_4708,N_1624);
or U9314 (N_9314,N_2648,N_46);
or U9315 (N_9315,N_139,N_284);
nor U9316 (N_9316,N_1799,N_2678);
and U9317 (N_9317,N_758,N_2170);
or U9318 (N_9318,N_592,N_3020);
or U9319 (N_9319,N_5456,N_19);
and U9320 (N_9320,N_3178,N_3753);
and U9321 (N_9321,N_3362,N_4571);
nor U9322 (N_9322,N_3890,N_5407);
or U9323 (N_9323,N_2621,N_2991);
nor U9324 (N_9324,N_2879,N_1529);
or U9325 (N_9325,N_2864,N_733);
or U9326 (N_9326,N_5678,N_2032);
or U9327 (N_9327,N_4385,N_3273);
or U9328 (N_9328,N_1811,N_3169);
nand U9329 (N_9329,N_4878,N_2248);
nor U9330 (N_9330,N_1593,N_5262);
or U9331 (N_9331,N_5083,N_267);
or U9332 (N_9332,N_2668,N_1057);
nand U9333 (N_9333,N_4805,N_4750);
nor U9334 (N_9334,N_5093,N_2127);
and U9335 (N_9335,N_4449,N_5610);
nor U9336 (N_9336,N_2278,N_1818);
nand U9337 (N_9337,N_104,N_1151);
xnor U9338 (N_9338,N_1248,N_989);
nor U9339 (N_9339,N_964,N_3508);
or U9340 (N_9340,N_602,N_209);
and U9341 (N_9341,N_1521,N_5464);
nand U9342 (N_9342,N_5503,N_3881);
or U9343 (N_9343,N_818,N_1824);
nor U9344 (N_9344,N_3036,N_63);
and U9345 (N_9345,N_4613,N_1061);
nand U9346 (N_9346,N_4234,N_3300);
and U9347 (N_9347,N_148,N_5477);
nand U9348 (N_9348,N_5024,N_4485);
and U9349 (N_9349,N_3391,N_3758);
and U9350 (N_9350,N_3727,N_5456);
xnor U9351 (N_9351,N_5890,N_4601);
or U9352 (N_9352,N_5749,N_630);
or U9353 (N_9353,N_1739,N_4170);
nand U9354 (N_9354,N_5640,N_4341);
and U9355 (N_9355,N_3248,N_3642);
nand U9356 (N_9356,N_5510,N_2581);
and U9357 (N_9357,N_395,N_4646);
nand U9358 (N_9358,N_525,N_4454);
nor U9359 (N_9359,N_4452,N_5505);
and U9360 (N_9360,N_2574,N_3097);
nor U9361 (N_9361,N_1219,N_1624);
and U9362 (N_9362,N_710,N_5430);
nand U9363 (N_9363,N_1768,N_2528);
or U9364 (N_9364,N_4250,N_1025);
and U9365 (N_9365,N_5420,N_443);
and U9366 (N_9366,N_2732,N_4270);
nor U9367 (N_9367,N_4846,N_1699);
or U9368 (N_9368,N_3387,N_2711);
xor U9369 (N_9369,N_1578,N_3063);
and U9370 (N_9370,N_273,N_3831);
nor U9371 (N_9371,N_4520,N_482);
xnor U9372 (N_9372,N_687,N_4269);
nand U9373 (N_9373,N_3410,N_4452);
nor U9374 (N_9374,N_4189,N_1761);
nand U9375 (N_9375,N_2999,N_1653);
xnor U9376 (N_9376,N_5719,N_5177);
and U9377 (N_9377,N_572,N_4128);
nand U9378 (N_9378,N_5586,N_2115);
xnor U9379 (N_9379,N_4107,N_2583);
or U9380 (N_9380,N_3096,N_5555);
nand U9381 (N_9381,N_2001,N_5985);
nand U9382 (N_9382,N_4606,N_5920);
or U9383 (N_9383,N_1494,N_1656);
nor U9384 (N_9384,N_619,N_2216);
and U9385 (N_9385,N_4041,N_1030);
nand U9386 (N_9386,N_2377,N_4486);
nand U9387 (N_9387,N_3800,N_1739);
nand U9388 (N_9388,N_3685,N_1452);
nand U9389 (N_9389,N_3244,N_3663);
and U9390 (N_9390,N_5407,N_1166);
nand U9391 (N_9391,N_4900,N_1898);
nor U9392 (N_9392,N_635,N_5850);
and U9393 (N_9393,N_5498,N_2191);
nor U9394 (N_9394,N_1775,N_5946);
nor U9395 (N_9395,N_1706,N_4423);
or U9396 (N_9396,N_5887,N_1726);
xor U9397 (N_9397,N_3632,N_5708);
nor U9398 (N_9398,N_2393,N_5381);
nor U9399 (N_9399,N_5536,N_5001);
nor U9400 (N_9400,N_655,N_1892);
or U9401 (N_9401,N_5214,N_394);
nor U9402 (N_9402,N_1938,N_3788);
nor U9403 (N_9403,N_1953,N_110);
nand U9404 (N_9404,N_2777,N_1760);
or U9405 (N_9405,N_4609,N_3111);
nand U9406 (N_9406,N_445,N_5661);
or U9407 (N_9407,N_1399,N_4241);
nand U9408 (N_9408,N_5693,N_1010);
nand U9409 (N_9409,N_237,N_1216);
and U9410 (N_9410,N_5240,N_4778);
or U9411 (N_9411,N_297,N_3543);
xnor U9412 (N_9412,N_5333,N_2706);
xnor U9413 (N_9413,N_729,N_2970);
and U9414 (N_9414,N_2503,N_1170);
or U9415 (N_9415,N_4121,N_4910);
and U9416 (N_9416,N_779,N_3876);
or U9417 (N_9417,N_5729,N_4187);
nand U9418 (N_9418,N_2850,N_5570);
or U9419 (N_9419,N_941,N_1539);
or U9420 (N_9420,N_59,N_1751);
nand U9421 (N_9421,N_2887,N_4940);
nor U9422 (N_9422,N_3620,N_1971);
and U9423 (N_9423,N_4123,N_3189);
nand U9424 (N_9424,N_5348,N_4307);
nor U9425 (N_9425,N_2769,N_3659);
and U9426 (N_9426,N_667,N_687);
or U9427 (N_9427,N_3834,N_3818);
and U9428 (N_9428,N_4877,N_4899);
nand U9429 (N_9429,N_1437,N_5615);
nand U9430 (N_9430,N_999,N_4709);
xnor U9431 (N_9431,N_1907,N_2786);
xnor U9432 (N_9432,N_5790,N_1391);
xor U9433 (N_9433,N_3296,N_3911);
and U9434 (N_9434,N_5724,N_4372);
or U9435 (N_9435,N_752,N_4388);
and U9436 (N_9436,N_463,N_3981);
nor U9437 (N_9437,N_5831,N_792);
nand U9438 (N_9438,N_2530,N_4594);
and U9439 (N_9439,N_1392,N_4704);
or U9440 (N_9440,N_5001,N_5207);
xor U9441 (N_9441,N_2916,N_3328);
nand U9442 (N_9442,N_2818,N_4960);
nand U9443 (N_9443,N_4875,N_3814);
nor U9444 (N_9444,N_2539,N_5696);
nand U9445 (N_9445,N_1521,N_729);
nor U9446 (N_9446,N_1207,N_4014);
and U9447 (N_9447,N_1307,N_600);
nand U9448 (N_9448,N_3991,N_3615);
and U9449 (N_9449,N_5523,N_5425);
xor U9450 (N_9450,N_279,N_574);
nand U9451 (N_9451,N_574,N_971);
or U9452 (N_9452,N_1084,N_4667);
nand U9453 (N_9453,N_3845,N_317);
nand U9454 (N_9454,N_4433,N_1848);
and U9455 (N_9455,N_4980,N_580);
and U9456 (N_9456,N_4465,N_3117);
and U9457 (N_9457,N_1106,N_2588);
and U9458 (N_9458,N_4508,N_5859);
nand U9459 (N_9459,N_831,N_1023);
or U9460 (N_9460,N_4383,N_2022);
nand U9461 (N_9461,N_2169,N_2700);
nand U9462 (N_9462,N_4473,N_3955);
xor U9463 (N_9463,N_3390,N_733);
xor U9464 (N_9464,N_2712,N_4164);
nor U9465 (N_9465,N_467,N_3614);
or U9466 (N_9466,N_5677,N_4401);
xnor U9467 (N_9467,N_1288,N_3267);
xnor U9468 (N_9468,N_947,N_3045);
or U9469 (N_9469,N_3673,N_1955);
and U9470 (N_9470,N_924,N_1152);
and U9471 (N_9471,N_3323,N_3904);
or U9472 (N_9472,N_2749,N_1842);
and U9473 (N_9473,N_4031,N_266);
or U9474 (N_9474,N_517,N_3727);
or U9475 (N_9475,N_217,N_1161);
nor U9476 (N_9476,N_2960,N_5553);
nor U9477 (N_9477,N_1192,N_3024);
and U9478 (N_9478,N_3192,N_616);
xnor U9479 (N_9479,N_954,N_3842);
nor U9480 (N_9480,N_695,N_4112);
or U9481 (N_9481,N_3499,N_3821);
nor U9482 (N_9482,N_5991,N_3535);
or U9483 (N_9483,N_3634,N_3239);
nand U9484 (N_9484,N_2853,N_2595);
or U9485 (N_9485,N_2203,N_5194);
nor U9486 (N_9486,N_1641,N_5912);
nand U9487 (N_9487,N_1812,N_3064);
or U9488 (N_9488,N_325,N_3593);
and U9489 (N_9489,N_5706,N_3457);
xor U9490 (N_9490,N_2916,N_5981);
nor U9491 (N_9491,N_2525,N_1221);
nand U9492 (N_9492,N_4552,N_2934);
nand U9493 (N_9493,N_5479,N_2016);
nor U9494 (N_9494,N_3134,N_1701);
and U9495 (N_9495,N_5362,N_804);
and U9496 (N_9496,N_4797,N_5149);
nand U9497 (N_9497,N_3461,N_749);
and U9498 (N_9498,N_5200,N_750);
and U9499 (N_9499,N_2619,N_2125);
and U9500 (N_9500,N_1875,N_114);
or U9501 (N_9501,N_2966,N_3121);
xor U9502 (N_9502,N_4078,N_3946);
nand U9503 (N_9503,N_2141,N_5330);
nor U9504 (N_9504,N_255,N_5453);
xor U9505 (N_9505,N_2350,N_4909);
xnor U9506 (N_9506,N_2892,N_2828);
or U9507 (N_9507,N_2681,N_3672);
or U9508 (N_9508,N_5072,N_5537);
and U9509 (N_9509,N_5627,N_1790);
nor U9510 (N_9510,N_5875,N_67);
nor U9511 (N_9511,N_3134,N_1426);
and U9512 (N_9512,N_4765,N_3561);
or U9513 (N_9513,N_1997,N_4350);
nand U9514 (N_9514,N_5135,N_1254);
nand U9515 (N_9515,N_5569,N_1504);
xor U9516 (N_9516,N_1080,N_1365);
or U9517 (N_9517,N_376,N_5467);
or U9518 (N_9518,N_254,N_5709);
nor U9519 (N_9519,N_1506,N_3761);
nand U9520 (N_9520,N_1637,N_2328);
nand U9521 (N_9521,N_1385,N_913);
nand U9522 (N_9522,N_5754,N_746);
nand U9523 (N_9523,N_2021,N_5381);
nand U9524 (N_9524,N_200,N_4564);
and U9525 (N_9525,N_1457,N_3450);
or U9526 (N_9526,N_1230,N_978);
or U9527 (N_9527,N_3008,N_4470);
nor U9528 (N_9528,N_2977,N_1103);
or U9529 (N_9529,N_5263,N_3985);
nand U9530 (N_9530,N_474,N_441);
nand U9531 (N_9531,N_4107,N_5099);
xor U9532 (N_9532,N_3059,N_1907);
and U9533 (N_9533,N_2818,N_2121);
nand U9534 (N_9534,N_3869,N_3533);
nor U9535 (N_9535,N_339,N_5659);
nor U9536 (N_9536,N_2559,N_5056);
nor U9537 (N_9537,N_3500,N_5067);
nor U9538 (N_9538,N_336,N_2069);
and U9539 (N_9539,N_4999,N_5875);
xor U9540 (N_9540,N_962,N_1707);
and U9541 (N_9541,N_565,N_2140);
and U9542 (N_9542,N_2445,N_5582);
and U9543 (N_9543,N_2818,N_1332);
nor U9544 (N_9544,N_459,N_1299);
nor U9545 (N_9545,N_4847,N_5795);
and U9546 (N_9546,N_4017,N_2462);
nor U9547 (N_9547,N_374,N_3144);
nand U9548 (N_9548,N_2640,N_2363);
xnor U9549 (N_9549,N_5293,N_4819);
nand U9550 (N_9550,N_5870,N_1775);
or U9551 (N_9551,N_357,N_4335);
nand U9552 (N_9552,N_5051,N_5588);
nand U9553 (N_9553,N_4198,N_329);
nor U9554 (N_9554,N_1241,N_858);
or U9555 (N_9555,N_1301,N_3118);
nor U9556 (N_9556,N_5099,N_5647);
nor U9557 (N_9557,N_3343,N_1218);
xnor U9558 (N_9558,N_1154,N_336);
or U9559 (N_9559,N_5626,N_5415);
xnor U9560 (N_9560,N_2587,N_4269);
or U9561 (N_9561,N_448,N_4470);
nand U9562 (N_9562,N_1360,N_5159);
or U9563 (N_9563,N_5779,N_3677);
nor U9564 (N_9564,N_2446,N_1283);
nand U9565 (N_9565,N_2806,N_5279);
or U9566 (N_9566,N_2566,N_5304);
nand U9567 (N_9567,N_3449,N_2415);
or U9568 (N_9568,N_4449,N_2833);
or U9569 (N_9569,N_649,N_5403);
and U9570 (N_9570,N_1378,N_1790);
nor U9571 (N_9571,N_52,N_487);
xor U9572 (N_9572,N_944,N_1496);
nand U9573 (N_9573,N_2494,N_3580);
and U9574 (N_9574,N_785,N_2651);
nand U9575 (N_9575,N_4853,N_3994);
and U9576 (N_9576,N_2221,N_1798);
and U9577 (N_9577,N_5032,N_4459);
nand U9578 (N_9578,N_5254,N_2471);
or U9579 (N_9579,N_4496,N_4726);
xnor U9580 (N_9580,N_3991,N_2216);
and U9581 (N_9581,N_1051,N_5374);
nor U9582 (N_9582,N_3054,N_5209);
and U9583 (N_9583,N_5278,N_3288);
xor U9584 (N_9584,N_4423,N_1022);
nor U9585 (N_9585,N_4769,N_2397);
nand U9586 (N_9586,N_5258,N_3551);
nor U9587 (N_9587,N_2448,N_863);
and U9588 (N_9588,N_2523,N_2589);
nand U9589 (N_9589,N_3021,N_3159);
and U9590 (N_9590,N_112,N_2695);
xor U9591 (N_9591,N_5254,N_3044);
nor U9592 (N_9592,N_5120,N_5277);
nand U9593 (N_9593,N_867,N_3892);
xnor U9594 (N_9594,N_5721,N_349);
and U9595 (N_9595,N_1748,N_3943);
nand U9596 (N_9596,N_3890,N_2893);
or U9597 (N_9597,N_1934,N_5119);
or U9598 (N_9598,N_1769,N_1864);
or U9599 (N_9599,N_4569,N_4562);
nor U9600 (N_9600,N_4023,N_728);
nor U9601 (N_9601,N_769,N_3284);
nand U9602 (N_9602,N_1074,N_4574);
or U9603 (N_9603,N_4463,N_1315);
nand U9604 (N_9604,N_92,N_684);
xnor U9605 (N_9605,N_5571,N_3366);
xor U9606 (N_9606,N_3527,N_2227);
xnor U9607 (N_9607,N_173,N_544);
nand U9608 (N_9608,N_2742,N_5168);
nor U9609 (N_9609,N_5777,N_4396);
xor U9610 (N_9610,N_3406,N_4854);
or U9611 (N_9611,N_5095,N_1606);
or U9612 (N_9612,N_3603,N_2125);
nand U9613 (N_9613,N_5513,N_4739);
or U9614 (N_9614,N_616,N_2522);
or U9615 (N_9615,N_1331,N_514);
and U9616 (N_9616,N_4895,N_131);
nand U9617 (N_9617,N_373,N_343);
and U9618 (N_9618,N_760,N_3475);
nand U9619 (N_9619,N_5890,N_527);
or U9620 (N_9620,N_3991,N_2253);
or U9621 (N_9621,N_4119,N_350);
and U9622 (N_9622,N_222,N_415);
and U9623 (N_9623,N_2887,N_3233);
nand U9624 (N_9624,N_3257,N_4552);
nand U9625 (N_9625,N_749,N_2563);
or U9626 (N_9626,N_1432,N_1014);
and U9627 (N_9627,N_2240,N_4107);
or U9628 (N_9628,N_4938,N_3387);
or U9629 (N_9629,N_5831,N_1588);
nor U9630 (N_9630,N_5130,N_1844);
nor U9631 (N_9631,N_669,N_5332);
and U9632 (N_9632,N_3824,N_4062);
nand U9633 (N_9633,N_2650,N_2308);
or U9634 (N_9634,N_4698,N_2765);
nand U9635 (N_9635,N_4039,N_5877);
or U9636 (N_9636,N_4266,N_2376);
and U9637 (N_9637,N_5055,N_80);
nand U9638 (N_9638,N_831,N_1084);
nor U9639 (N_9639,N_5962,N_940);
nor U9640 (N_9640,N_5316,N_2066);
nor U9641 (N_9641,N_1679,N_2177);
or U9642 (N_9642,N_2653,N_1070);
and U9643 (N_9643,N_4964,N_2017);
or U9644 (N_9644,N_1518,N_268);
nand U9645 (N_9645,N_808,N_4809);
or U9646 (N_9646,N_4440,N_3277);
and U9647 (N_9647,N_3091,N_2282);
xor U9648 (N_9648,N_2374,N_1696);
and U9649 (N_9649,N_5545,N_145);
or U9650 (N_9650,N_300,N_3808);
nor U9651 (N_9651,N_5197,N_3381);
and U9652 (N_9652,N_2151,N_4553);
nand U9653 (N_9653,N_941,N_3168);
or U9654 (N_9654,N_3598,N_3509);
xnor U9655 (N_9655,N_5784,N_559);
or U9656 (N_9656,N_2304,N_455);
or U9657 (N_9657,N_4268,N_4118);
nand U9658 (N_9658,N_3662,N_4063);
xor U9659 (N_9659,N_5726,N_2371);
nor U9660 (N_9660,N_1687,N_5606);
nand U9661 (N_9661,N_479,N_4668);
xor U9662 (N_9662,N_1155,N_2876);
nor U9663 (N_9663,N_3715,N_3828);
nor U9664 (N_9664,N_1485,N_5331);
nand U9665 (N_9665,N_2383,N_2895);
nand U9666 (N_9666,N_1759,N_109);
nor U9667 (N_9667,N_2681,N_2937);
nand U9668 (N_9668,N_5055,N_1487);
nand U9669 (N_9669,N_3486,N_384);
nand U9670 (N_9670,N_5087,N_5948);
nand U9671 (N_9671,N_4225,N_3181);
and U9672 (N_9672,N_1747,N_3765);
and U9673 (N_9673,N_4199,N_3529);
nor U9674 (N_9674,N_520,N_1979);
nor U9675 (N_9675,N_322,N_1765);
and U9676 (N_9676,N_3255,N_3137);
nand U9677 (N_9677,N_3839,N_5157);
nor U9678 (N_9678,N_5080,N_89);
and U9679 (N_9679,N_2498,N_1127);
or U9680 (N_9680,N_3578,N_141);
or U9681 (N_9681,N_5314,N_1038);
and U9682 (N_9682,N_5658,N_5274);
nand U9683 (N_9683,N_5585,N_5849);
and U9684 (N_9684,N_1871,N_4180);
nor U9685 (N_9685,N_4445,N_2161);
or U9686 (N_9686,N_1166,N_1931);
xor U9687 (N_9687,N_2133,N_2267);
nand U9688 (N_9688,N_4928,N_4685);
or U9689 (N_9689,N_710,N_138);
xnor U9690 (N_9690,N_2214,N_2108);
nand U9691 (N_9691,N_5967,N_5537);
and U9692 (N_9692,N_786,N_2562);
nor U9693 (N_9693,N_5353,N_4093);
nor U9694 (N_9694,N_1980,N_188);
nor U9695 (N_9695,N_3322,N_5398);
and U9696 (N_9696,N_4020,N_5350);
nor U9697 (N_9697,N_935,N_5206);
or U9698 (N_9698,N_5266,N_5077);
or U9699 (N_9699,N_3114,N_3495);
nand U9700 (N_9700,N_4357,N_2658);
nor U9701 (N_9701,N_4360,N_5728);
nor U9702 (N_9702,N_3502,N_1874);
or U9703 (N_9703,N_1585,N_1057);
nor U9704 (N_9704,N_1366,N_5958);
or U9705 (N_9705,N_423,N_4577);
nand U9706 (N_9706,N_2305,N_4446);
nor U9707 (N_9707,N_4448,N_4148);
nor U9708 (N_9708,N_3305,N_564);
nor U9709 (N_9709,N_3930,N_123);
nand U9710 (N_9710,N_3444,N_172);
or U9711 (N_9711,N_138,N_4744);
or U9712 (N_9712,N_930,N_3781);
or U9713 (N_9713,N_3845,N_4094);
nand U9714 (N_9714,N_937,N_2629);
nand U9715 (N_9715,N_4997,N_2770);
or U9716 (N_9716,N_3007,N_3779);
or U9717 (N_9717,N_202,N_2485);
nand U9718 (N_9718,N_5372,N_2083);
and U9719 (N_9719,N_151,N_5671);
nor U9720 (N_9720,N_4981,N_5727);
or U9721 (N_9721,N_2631,N_3575);
or U9722 (N_9722,N_5238,N_5534);
or U9723 (N_9723,N_2429,N_5208);
or U9724 (N_9724,N_1494,N_3672);
xor U9725 (N_9725,N_1336,N_3718);
or U9726 (N_9726,N_5916,N_21);
and U9727 (N_9727,N_5327,N_2054);
nor U9728 (N_9728,N_2103,N_1706);
and U9729 (N_9729,N_3123,N_798);
and U9730 (N_9730,N_1585,N_1345);
nand U9731 (N_9731,N_2104,N_5231);
nor U9732 (N_9732,N_5639,N_2982);
nand U9733 (N_9733,N_5518,N_2143);
and U9734 (N_9734,N_4053,N_2004);
xor U9735 (N_9735,N_393,N_85);
nand U9736 (N_9736,N_3070,N_1404);
and U9737 (N_9737,N_159,N_3396);
and U9738 (N_9738,N_1708,N_2168);
and U9739 (N_9739,N_4765,N_1669);
nor U9740 (N_9740,N_1099,N_5700);
nor U9741 (N_9741,N_1049,N_5649);
nand U9742 (N_9742,N_5984,N_4388);
nor U9743 (N_9743,N_146,N_5800);
nor U9744 (N_9744,N_2244,N_4032);
xor U9745 (N_9745,N_3586,N_4863);
nor U9746 (N_9746,N_5386,N_751);
and U9747 (N_9747,N_5351,N_5382);
or U9748 (N_9748,N_969,N_2128);
or U9749 (N_9749,N_1470,N_329);
or U9750 (N_9750,N_4201,N_1101);
or U9751 (N_9751,N_1006,N_2714);
and U9752 (N_9752,N_4578,N_3756);
or U9753 (N_9753,N_149,N_4594);
nor U9754 (N_9754,N_1017,N_3335);
or U9755 (N_9755,N_4539,N_4759);
xnor U9756 (N_9756,N_3510,N_4705);
or U9757 (N_9757,N_3969,N_636);
nor U9758 (N_9758,N_1926,N_5793);
xor U9759 (N_9759,N_1407,N_5041);
and U9760 (N_9760,N_748,N_1696);
and U9761 (N_9761,N_3602,N_5542);
nand U9762 (N_9762,N_1933,N_269);
nand U9763 (N_9763,N_3451,N_1838);
or U9764 (N_9764,N_1656,N_4311);
or U9765 (N_9765,N_5202,N_2846);
and U9766 (N_9766,N_2954,N_5266);
and U9767 (N_9767,N_466,N_3793);
and U9768 (N_9768,N_4,N_5410);
nor U9769 (N_9769,N_5581,N_2856);
and U9770 (N_9770,N_3736,N_1207);
nor U9771 (N_9771,N_3474,N_2921);
nor U9772 (N_9772,N_4929,N_5808);
nand U9773 (N_9773,N_838,N_3129);
xnor U9774 (N_9774,N_4270,N_2797);
xnor U9775 (N_9775,N_3576,N_4516);
nor U9776 (N_9776,N_2812,N_3090);
nand U9777 (N_9777,N_2148,N_3081);
and U9778 (N_9778,N_1882,N_3410);
and U9779 (N_9779,N_1316,N_3976);
and U9780 (N_9780,N_2666,N_1210);
or U9781 (N_9781,N_3935,N_4307);
or U9782 (N_9782,N_3137,N_1957);
and U9783 (N_9783,N_3439,N_1758);
nand U9784 (N_9784,N_4358,N_473);
or U9785 (N_9785,N_2806,N_2484);
or U9786 (N_9786,N_2418,N_342);
nand U9787 (N_9787,N_4579,N_3926);
nor U9788 (N_9788,N_4725,N_5100);
nor U9789 (N_9789,N_1134,N_4435);
nor U9790 (N_9790,N_1319,N_4396);
and U9791 (N_9791,N_3100,N_5311);
and U9792 (N_9792,N_679,N_5162);
and U9793 (N_9793,N_4652,N_4791);
nand U9794 (N_9794,N_3057,N_1812);
nand U9795 (N_9795,N_5132,N_2916);
nand U9796 (N_9796,N_2355,N_3597);
or U9797 (N_9797,N_3836,N_330);
and U9798 (N_9798,N_2928,N_3022);
or U9799 (N_9799,N_3006,N_4242);
nand U9800 (N_9800,N_4670,N_5361);
nor U9801 (N_9801,N_2833,N_2878);
and U9802 (N_9802,N_4441,N_1769);
nand U9803 (N_9803,N_4165,N_2704);
nand U9804 (N_9804,N_4872,N_2921);
nand U9805 (N_9805,N_3462,N_1047);
or U9806 (N_9806,N_5826,N_2458);
nand U9807 (N_9807,N_2246,N_945);
nand U9808 (N_9808,N_1200,N_3434);
nor U9809 (N_9809,N_2006,N_2433);
xnor U9810 (N_9810,N_3180,N_3441);
or U9811 (N_9811,N_4105,N_394);
or U9812 (N_9812,N_1779,N_5118);
nand U9813 (N_9813,N_3873,N_4275);
and U9814 (N_9814,N_479,N_568);
nand U9815 (N_9815,N_4256,N_5796);
nor U9816 (N_9816,N_4917,N_269);
and U9817 (N_9817,N_4352,N_2439);
or U9818 (N_9818,N_621,N_2845);
nand U9819 (N_9819,N_501,N_2537);
nand U9820 (N_9820,N_1048,N_281);
and U9821 (N_9821,N_5164,N_2051);
xnor U9822 (N_9822,N_371,N_749);
nand U9823 (N_9823,N_2247,N_5575);
or U9824 (N_9824,N_2939,N_1249);
nand U9825 (N_9825,N_3137,N_1583);
xnor U9826 (N_9826,N_5426,N_2543);
xnor U9827 (N_9827,N_2552,N_3507);
and U9828 (N_9828,N_3251,N_389);
or U9829 (N_9829,N_966,N_1876);
and U9830 (N_9830,N_354,N_3075);
or U9831 (N_9831,N_321,N_3987);
and U9832 (N_9832,N_2759,N_1361);
nand U9833 (N_9833,N_2934,N_4678);
or U9834 (N_9834,N_3820,N_5548);
nand U9835 (N_9835,N_4767,N_4245);
and U9836 (N_9836,N_5397,N_3406);
nand U9837 (N_9837,N_1745,N_2356);
or U9838 (N_9838,N_2087,N_485);
nand U9839 (N_9839,N_600,N_5998);
and U9840 (N_9840,N_3260,N_382);
nand U9841 (N_9841,N_5584,N_158);
nor U9842 (N_9842,N_31,N_2758);
nand U9843 (N_9843,N_645,N_2486);
or U9844 (N_9844,N_273,N_2088);
nand U9845 (N_9845,N_2343,N_1932);
and U9846 (N_9846,N_2065,N_4771);
and U9847 (N_9847,N_5151,N_3213);
nor U9848 (N_9848,N_4335,N_374);
and U9849 (N_9849,N_882,N_767);
or U9850 (N_9850,N_1061,N_2990);
nand U9851 (N_9851,N_1206,N_5030);
nor U9852 (N_9852,N_5473,N_3684);
and U9853 (N_9853,N_202,N_3941);
nand U9854 (N_9854,N_2695,N_4143);
nand U9855 (N_9855,N_2842,N_4927);
or U9856 (N_9856,N_3659,N_1637);
xor U9857 (N_9857,N_78,N_3021);
nand U9858 (N_9858,N_1378,N_4772);
and U9859 (N_9859,N_4522,N_527);
and U9860 (N_9860,N_1002,N_5943);
nand U9861 (N_9861,N_3948,N_3741);
and U9862 (N_9862,N_46,N_3536);
xnor U9863 (N_9863,N_3251,N_4617);
nor U9864 (N_9864,N_3575,N_4235);
or U9865 (N_9865,N_2424,N_1399);
or U9866 (N_9866,N_959,N_3814);
or U9867 (N_9867,N_460,N_583);
or U9868 (N_9868,N_5869,N_5903);
nand U9869 (N_9869,N_5413,N_978);
or U9870 (N_9870,N_2613,N_3188);
and U9871 (N_9871,N_2220,N_2743);
xnor U9872 (N_9872,N_4473,N_4969);
and U9873 (N_9873,N_4202,N_925);
nor U9874 (N_9874,N_5630,N_3021);
and U9875 (N_9875,N_2746,N_441);
nor U9876 (N_9876,N_3520,N_1869);
nand U9877 (N_9877,N_1203,N_2037);
nor U9878 (N_9878,N_4161,N_1656);
or U9879 (N_9879,N_5153,N_2944);
and U9880 (N_9880,N_664,N_2643);
or U9881 (N_9881,N_4711,N_5586);
nor U9882 (N_9882,N_822,N_4055);
xor U9883 (N_9883,N_5043,N_4574);
nand U9884 (N_9884,N_1958,N_2253);
or U9885 (N_9885,N_4150,N_5390);
nand U9886 (N_9886,N_5506,N_5329);
or U9887 (N_9887,N_1303,N_4694);
nand U9888 (N_9888,N_1395,N_416);
and U9889 (N_9889,N_2385,N_3103);
or U9890 (N_9890,N_3003,N_336);
or U9891 (N_9891,N_1145,N_3761);
nor U9892 (N_9892,N_117,N_963);
nor U9893 (N_9893,N_3926,N_4403);
nor U9894 (N_9894,N_4623,N_1191);
and U9895 (N_9895,N_527,N_5547);
nor U9896 (N_9896,N_4129,N_3019);
xor U9897 (N_9897,N_3234,N_1778);
or U9898 (N_9898,N_3563,N_4913);
or U9899 (N_9899,N_319,N_2185);
or U9900 (N_9900,N_5617,N_1077);
or U9901 (N_9901,N_3992,N_417);
nor U9902 (N_9902,N_3953,N_4356);
or U9903 (N_9903,N_1410,N_5007);
nand U9904 (N_9904,N_1067,N_2506);
nand U9905 (N_9905,N_2536,N_1694);
nor U9906 (N_9906,N_1051,N_1429);
and U9907 (N_9907,N_3649,N_5331);
and U9908 (N_9908,N_5685,N_1192);
xnor U9909 (N_9909,N_5680,N_4840);
and U9910 (N_9910,N_490,N_3533);
nor U9911 (N_9911,N_239,N_688);
and U9912 (N_9912,N_5458,N_1120);
xor U9913 (N_9913,N_1263,N_695);
or U9914 (N_9914,N_5595,N_1169);
or U9915 (N_9915,N_3972,N_5788);
or U9916 (N_9916,N_5665,N_4670);
nand U9917 (N_9917,N_3173,N_2824);
xnor U9918 (N_9918,N_2192,N_2841);
or U9919 (N_9919,N_274,N_5909);
nand U9920 (N_9920,N_3654,N_5839);
and U9921 (N_9921,N_178,N_1581);
or U9922 (N_9922,N_673,N_665);
or U9923 (N_9923,N_1070,N_4483);
or U9924 (N_9924,N_4203,N_1499);
nor U9925 (N_9925,N_1581,N_2994);
xnor U9926 (N_9926,N_3454,N_3322);
nor U9927 (N_9927,N_4410,N_1061);
or U9928 (N_9928,N_409,N_3142);
and U9929 (N_9929,N_290,N_5472);
nand U9930 (N_9930,N_609,N_349);
nand U9931 (N_9931,N_4606,N_1337);
and U9932 (N_9932,N_2256,N_1570);
and U9933 (N_9933,N_1584,N_3862);
nand U9934 (N_9934,N_5125,N_744);
xnor U9935 (N_9935,N_788,N_3820);
or U9936 (N_9936,N_5309,N_5839);
or U9937 (N_9937,N_1089,N_4213);
or U9938 (N_9938,N_52,N_1832);
and U9939 (N_9939,N_1092,N_3800);
or U9940 (N_9940,N_3266,N_951);
nor U9941 (N_9941,N_3914,N_4637);
and U9942 (N_9942,N_1162,N_578);
xnor U9943 (N_9943,N_2225,N_5138);
and U9944 (N_9944,N_4785,N_5421);
nor U9945 (N_9945,N_3095,N_4098);
and U9946 (N_9946,N_3916,N_3127);
nand U9947 (N_9947,N_915,N_3272);
xor U9948 (N_9948,N_3967,N_872);
nand U9949 (N_9949,N_1104,N_4464);
or U9950 (N_9950,N_1885,N_3851);
xnor U9951 (N_9951,N_1486,N_160);
or U9952 (N_9952,N_5709,N_2188);
nor U9953 (N_9953,N_94,N_4829);
and U9954 (N_9954,N_862,N_5352);
nand U9955 (N_9955,N_4083,N_1530);
nand U9956 (N_9956,N_5636,N_5976);
nand U9957 (N_9957,N_4344,N_4664);
nand U9958 (N_9958,N_505,N_1447);
or U9959 (N_9959,N_5176,N_3312);
nor U9960 (N_9960,N_97,N_511);
and U9961 (N_9961,N_397,N_1724);
nor U9962 (N_9962,N_1938,N_714);
nor U9963 (N_9963,N_2518,N_3391);
or U9964 (N_9964,N_2187,N_3664);
and U9965 (N_9965,N_1931,N_89);
or U9966 (N_9966,N_1369,N_545);
xnor U9967 (N_9967,N_1181,N_4988);
nand U9968 (N_9968,N_4713,N_5934);
or U9969 (N_9969,N_3860,N_2983);
and U9970 (N_9970,N_1706,N_3327);
nor U9971 (N_9971,N_4654,N_1715);
xnor U9972 (N_9972,N_3791,N_1215);
nand U9973 (N_9973,N_3248,N_2604);
or U9974 (N_9974,N_2125,N_1131);
nor U9975 (N_9975,N_1617,N_332);
and U9976 (N_9976,N_4150,N_5183);
xnor U9977 (N_9977,N_5948,N_763);
nand U9978 (N_9978,N_5080,N_1582);
nand U9979 (N_9979,N_3985,N_5986);
nor U9980 (N_9980,N_3345,N_3737);
nor U9981 (N_9981,N_3380,N_180);
nor U9982 (N_9982,N_4460,N_68);
xnor U9983 (N_9983,N_2183,N_3988);
and U9984 (N_9984,N_3585,N_494);
xnor U9985 (N_9985,N_2993,N_4744);
or U9986 (N_9986,N_4487,N_2248);
or U9987 (N_9987,N_3424,N_4619);
nor U9988 (N_9988,N_1925,N_3453);
nor U9989 (N_9989,N_145,N_2068);
nor U9990 (N_9990,N_706,N_2049);
nor U9991 (N_9991,N_780,N_5768);
nand U9992 (N_9992,N_1124,N_714);
and U9993 (N_9993,N_3109,N_2357);
nor U9994 (N_9994,N_747,N_201);
nor U9995 (N_9995,N_5319,N_5069);
or U9996 (N_9996,N_2477,N_4871);
xnor U9997 (N_9997,N_5266,N_3141);
and U9998 (N_9998,N_184,N_1694);
nand U9999 (N_9999,N_3979,N_5719);
and U10000 (N_10000,N_5849,N_5272);
nor U10001 (N_10001,N_3148,N_558);
or U10002 (N_10002,N_2149,N_5119);
or U10003 (N_10003,N_3941,N_2325);
and U10004 (N_10004,N_4604,N_4995);
nand U10005 (N_10005,N_2981,N_4346);
or U10006 (N_10006,N_1222,N_4594);
and U10007 (N_10007,N_4387,N_3016);
and U10008 (N_10008,N_2007,N_4259);
nor U10009 (N_10009,N_4833,N_5969);
or U10010 (N_10010,N_2800,N_4712);
nor U10011 (N_10011,N_5056,N_2798);
or U10012 (N_10012,N_237,N_3422);
and U10013 (N_10013,N_699,N_2699);
or U10014 (N_10014,N_2631,N_1112);
xnor U10015 (N_10015,N_3168,N_3359);
nand U10016 (N_10016,N_631,N_4450);
and U10017 (N_10017,N_4689,N_3994);
and U10018 (N_10018,N_4907,N_529);
and U10019 (N_10019,N_1441,N_3324);
or U10020 (N_10020,N_286,N_1604);
and U10021 (N_10021,N_2115,N_4797);
nor U10022 (N_10022,N_463,N_1947);
and U10023 (N_10023,N_3733,N_125);
and U10024 (N_10024,N_1885,N_314);
xor U10025 (N_10025,N_3971,N_313);
nand U10026 (N_10026,N_5067,N_3073);
or U10027 (N_10027,N_512,N_4685);
or U10028 (N_10028,N_828,N_153);
and U10029 (N_10029,N_3981,N_3842);
and U10030 (N_10030,N_882,N_4329);
and U10031 (N_10031,N_1931,N_397);
nand U10032 (N_10032,N_4237,N_1132);
and U10033 (N_10033,N_4401,N_3788);
or U10034 (N_10034,N_4647,N_3374);
or U10035 (N_10035,N_5314,N_4113);
nand U10036 (N_10036,N_5767,N_5778);
nand U10037 (N_10037,N_1534,N_2828);
nand U10038 (N_10038,N_3446,N_3147);
nor U10039 (N_10039,N_2153,N_1892);
or U10040 (N_10040,N_5221,N_1978);
or U10041 (N_10041,N_4600,N_5168);
or U10042 (N_10042,N_3198,N_310);
or U10043 (N_10043,N_1411,N_2364);
or U10044 (N_10044,N_3861,N_5729);
or U10045 (N_10045,N_1154,N_4081);
and U10046 (N_10046,N_4577,N_435);
and U10047 (N_10047,N_4589,N_1861);
nand U10048 (N_10048,N_5515,N_1009);
xnor U10049 (N_10049,N_903,N_336);
or U10050 (N_10050,N_4631,N_2027);
nand U10051 (N_10051,N_3096,N_5613);
nand U10052 (N_10052,N_4497,N_5941);
xor U10053 (N_10053,N_4365,N_1435);
or U10054 (N_10054,N_1047,N_4701);
nor U10055 (N_10055,N_4918,N_3653);
nand U10056 (N_10056,N_4212,N_1431);
nand U10057 (N_10057,N_1963,N_4233);
and U10058 (N_10058,N_5487,N_34);
or U10059 (N_10059,N_2319,N_3943);
nand U10060 (N_10060,N_4636,N_633);
xnor U10061 (N_10061,N_4114,N_4268);
nor U10062 (N_10062,N_888,N_2598);
xor U10063 (N_10063,N_5975,N_411);
nand U10064 (N_10064,N_5268,N_1690);
nand U10065 (N_10065,N_1734,N_2890);
and U10066 (N_10066,N_4248,N_864);
and U10067 (N_10067,N_2317,N_259);
and U10068 (N_10068,N_1502,N_3672);
or U10069 (N_10069,N_2610,N_3865);
nor U10070 (N_10070,N_2126,N_2494);
or U10071 (N_10071,N_2671,N_2075);
nand U10072 (N_10072,N_4847,N_5330);
and U10073 (N_10073,N_128,N_3387);
nor U10074 (N_10074,N_1557,N_2299);
or U10075 (N_10075,N_4674,N_5921);
and U10076 (N_10076,N_3727,N_5987);
nor U10077 (N_10077,N_1815,N_5630);
or U10078 (N_10078,N_2077,N_5057);
and U10079 (N_10079,N_554,N_5870);
nor U10080 (N_10080,N_4274,N_1920);
nand U10081 (N_10081,N_5246,N_3436);
and U10082 (N_10082,N_3131,N_1671);
nor U10083 (N_10083,N_3852,N_4789);
nand U10084 (N_10084,N_4046,N_4010);
nor U10085 (N_10085,N_115,N_4522);
nor U10086 (N_10086,N_3477,N_5036);
nand U10087 (N_10087,N_5696,N_5807);
nor U10088 (N_10088,N_4207,N_4662);
xor U10089 (N_10089,N_1208,N_2980);
nand U10090 (N_10090,N_4802,N_5984);
or U10091 (N_10091,N_611,N_879);
nor U10092 (N_10092,N_5183,N_4550);
or U10093 (N_10093,N_3773,N_3823);
and U10094 (N_10094,N_5184,N_1841);
nand U10095 (N_10095,N_3497,N_4101);
nand U10096 (N_10096,N_5059,N_4473);
nand U10097 (N_10097,N_4504,N_546);
and U10098 (N_10098,N_2113,N_4024);
and U10099 (N_10099,N_4028,N_4833);
nand U10100 (N_10100,N_5586,N_5167);
and U10101 (N_10101,N_2695,N_5374);
nand U10102 (N_10102,N_3694,N_4282);
and U10103 (N_10103,N_1772,N_5761);
nand U10104 (N_10104,N_4820,N_2879);
nand U10105 (N_10105,N_5654,N_5640);
and U10106 (N_10106,N_3117,N_3297);
nor U10107 (N_10107,N_2861,N_3616);
nor U10108 (N_10108,N_498,N_1748);
and U10109 (N_10109,N_1628,N_3508);
nor U10110 (N_10110,N_1775,N_5819);
or U10111 (N_10111,N_5014,N_3065);
nor U10112 (N_10112,N_873,N_3222);
and U10113 (N_10113,N_686,N_2753);
xor U10114 (N_10114,N_4651,N_5772);
nand U10115 (N_10115,N_88,N_4562);
nand U10116 (N_10116,N_5958,N_1202);
and U10117 (N_10117,N_888,N_4169);
nor U10118 (N_10118,N_343,N_4086);
or U10119 (N_10119,N_5976,N_2339);
or U10120 (N_10120,N_128,N_169);
or U10121 (N_10121,N_292,N_4332);
and U10122 (N_10122,N_2812,N_1284);
or U10123 (N_10123,N_5108,N_3580);
nand U10124 (N_10124,N_5429,N_2349);
and U10125 (N_10125,N_5081,N_469);
and U10126 (N_10126,N_5379,N_4433);
nand U10127 (N_10127,N_1529,N_3395);
nand U10128 (N_10128,N_3212,N_5975);
and U10129 (N_10129,N_4345,N_5701);
xnor U10130 (N_10130,N_2251,N_1550);
and U10131 (N_10131,N_1840,N_3078);
or U10132 (N_10132,N_3754,N_1441);
nor U10133 (N_10133,N_5273,N_5566);
or U10134 (N_10134,N_1436,N_2518);
or U10135 (N_10135,N_1204,N_5378);
and U10136 (N_10136,N_2740,N_4980);
xor U10137 (N_10137,N_2888,N_557);
nand U10138 (N_10138,N_4981,N_3031);
and U10139 (N_10139,N_2937,N_567);
nor U10140 (N_10140,N_2817,N_2833);
and U10141 (N_10141,N_475,N_810);
nor U10142 (N_10142,N_310,N_1135);
or U10143 (N_10143,N_846,N_5233);
nor U10144 (N_10144,N_1391,N_383);
xor U10145 (N_10145,N_196,N_3822);
or U10146 (N_10146,N_533,N_5467);
nand U10147 (N_10147,N_573,N_3438);
nand U10148 (N_10148,N_2009,N_679);
and U10149 (N_10149,N_3374,N_674);
nand U10150 (N_10150,N_3664,N_3407);
nand U10151 (N_10151,N_1055,N_1585);
nor U10152 (N_10152,N_4010,N_805);
or U10153 (N_10153,N_3626,N_2662);
nand U10154 (N_10154,N_2910,N_2585);
xor U10155 (N_10155,N_4969,N_2102);
nand U10156 (N_10156,N_444,N_790);
nand U10157 (N_10157,N_3120,N_24);
or U10158 (N_10158,N_1804,N_5722);
or U10159 (N_10159,N_4903,N_2858);
xnor U10160 (N_10160,N_5086,N_5789);
xor U10161 (N_10161,N_2193,N_4823);
or U10162 (N_10162,N_5317,N_86);
nor U10163 (N_10163,N_3449,N_1381);
or U10164 (N_10164,N_5598,N_838);
nand U10165 (N_10165,N_1206,N_2208);
or U10166 (N_10166,N_1038,N_4018);
nor U10167 (N_10167,N_682,N_261);
or U10168 (N_10168,N_4629,N_2787);
nor U10169 (N_10169,N_409,N_3815);
or U10170 (N_10170,N_1027,N_4509);
and U10171 (N_10171,N_426,N_3842);
nor U10172 (N_10172,N_5506,N_5536);
or U10173 (N_10173,N_4120,N_5656);
nand U10174 (N_10174,N_1906,N_2502);
or U10175 (N_10175,N_3664,N_664);
nor U10176 (N_10176,N_3220,N_2192);
nand U10177 (N_10177,N_2906,N_5383);
or U10178 (N_10178,N_852,N_5252);
nand U10179 (N_10179,N_3431,N_1180);
and U10180 (N_10180,N_5715,N_2345);
or U10181 (N_10181,N_2997,N_79);
and U10182 (N_10182,N_4462,N_5059);
and U10183 (N_10183,N_2568,N_388);
or U10184 (N_10184,N_5052,N_4610);
and U10185 (N_10185,N_2014,N_2098);
nand U10186 (N_10186,N_1224,N_1896);
or U10187 (N_10187,N_3749,N_5691);
nor U10188 (N_10188,N_695,N_2325);
nand U10189 (N_10189,N_5396,N_5628);
nor U10190 (N_10190,N_74,N_4521);
nand U10191 (N_10191,N_4785,N_4088);
and U10192 (N_10192,N_1076,N_5445);
xor U10193 (N_10193,N_1581,N_1142);
nand U10194 (N_10194,N_1931,N_4638);
nor U10195 (N_10195,N_4091,N_2555);
and U10196 (N_10196,N_4626,N_943);
nand U10197 (N_10197,N_2159,N_1346);
or U10198 (N_10198,N_1342,N_3680);
and U10199 (N_10199,N_3854,N_4453);
or U10200 (N_10200,N_1969,N_3778);
or U10201 (N_10201,N_5588,N_4594);
nand U10202 (N_10202,N_1278,N_5868);
nor U10203 (N_10203,N_2391,N_1087);
and U10204 (N_10204,N_1066,N_3716);
nor U10205 (N_10205,N_4694,N_3925);
nor U10206 (N_10206,N_1100,N_1945);
nand U10207 (N_10207,N_1266,N_810);
nor U10208 (N_10208,N_3494,N_113);
nor U10209 (N_10209,N_5279,N_1633);
nand U10210 (N_10210,N_3537,N_2067);
and U10211 (N_10211,N_1174,N_1611);
or U10212 (N_10212,N_5884,N_2951);
and U10213 (N_10213,N_2080,N_2947);
nor U10214 (N_10214,N_3592,N_1900);
nor U10215 (N_10215,N_87,N_4006);
and U10216 (N_10216,N_3330,N_1218);
or U10217 (N_10217,N_2626,N_486);
and U10218 (N_10218,N_156,N_3103);
nand U10219 (N_10219,N_4108,N_2843);
or U10220 (N_10220,N_4935,N_2381);
and U10221 (N_10221,N_2016,N_4446);
nand U10222 (N_10222,N_5414,N_4331);
xnor U10223 (N_10223,N_2921,N_2939);
nor U10224 (N_10224,N_2567,N_4493);
nor U10225 (N_10225,N_306,N_2567);
nand U10226 (N_10226,N_1330,N_3760);
and U10227 (N_10227,N_2028,N_1157);
nand U10228 (N_10228,N_5380,N_1361);
nand U10229 (N_10229,N_5520,N_2451);
and U10230 (N_10230,N_1844,N_1278);
nor U10231 (N_10231,N_1959,N_2395);
or U10232 (N_10232,N_1563,N_2812);
nor U10233 (N_10233,N_4223,N_3957);
and U10234 (N_10234,N_4834,N_4351);
xnor U10235 (N_10235,N_4621,N_783);
nand U10236 (N_10236,N_1709,N_1964);
or U10237 (N_10237,N_4896,N_3452);
and U10238 (N_10238,N_5507,N_2846);
nor U10239 (N_10239,N_4041,N_1963);
nand U10240 (N_10240,N_2546,N_3101);
and U10241 (N_10241,N_120,N_5953);
and U10242 (N_10242,N_5001,N_1157);
nand U10243 (N_10243,N_1255,N_436);
and U10244 (N_10244,N_2105,N_1321);
and U10245 (N_10245,N_3582,N_117);
and U10246 (N_10246,N_2775,N_589);
nor U10247 (N_10247,N_5257,N_3667);
nand U10248 (N_10248,N_663,N_2935);
and U10249 (N_10249,N_1088,N_5276);
xor U10250 (N_10250,N_3043,N_3012);
nor U10251 (N_10251,N_2319,N_5370);
xnor U10252 (N_10252,N_3006,N_688);
and U10253 (N_10253,N_1671,N_1510);
nor U10254 (N_10254,N_3947,N_5577);
xnor U10255 (N_10255,N_4418,N_3896);
or U10256 (N_10256,N_3928,N_612);
or U10257 (N_10257,N_1695,N_5629);
nor U10258 (N_10258,N_4967,N_5182);
xnor U10259 (N_10259,N_4967,N_1243);
and U10260 (N_10260,N_5445,N_4432);
xor U10261 (N_10261,N_732,N_5970);
xnor U10262 (N_10262,N_1464,N_1551);
or U10263 (N_10263,N_3941,N_1752);
nor U10264 (N_10264,N_3081,N_5945);
nand U10265 (N_10265,N_1744,N_1716);
or U10266 (N_10266,N_3153,N_382);
nor U10267 (N_10267,N_4581,N_5214);
nand U10268 (N_10268,N_4961,N_5706);
and U10269 (N_10269,N_1735,N_3970);
nor U10270 (N_10270,N_3289,N_1335);
or U10271 (N_10271,N_3093,N_2384);
and U10272 (N_10272,N_4892,N_1636);
nand U10273 (N_10273,N_2303,N_2041);
or U10274 (N_10274,N_463,N_480);
and U10275 (N_10275,N_1982,N_4044);
nor U10276 (N_10276,N_511,N_3788);
or U10277 (N_10277,N_3684,N_2819);
or U10278 (N_10278,N_2783,N_1549);
or U10279 (N_10279,N_4792,N_4219);
or U10280 (N_10280,N_5604,N_1891);
and U10281 (N_10281,N_5377,N_3149);
nor U10282 (N_10282,N_5982,N_4787);
and U10283 (N_10283,N_2480,N_4448);
xnor U10284 (N_10284,N_3825,N_1058);
nand U10285 (N_10285,N_474,N_339);
nor U10286 (N_10286,N_424,N_749);
nand U10287 (N_10287,N_4311,N_2646);
and U10288 (N_10288,N_4265,N_1360);
and U10289 (N_10289,N_3982,N_5437);
or U10290 (N_10290,N_2803,N_1388);
xor U10291 (N_10291,N_5614,N_2592);
and U10292 (N_10292,N_2227,N_3422);
or U10293 (N_10293,N_1327,N_4437);
nor U10294 (N_10294,N_3630,N_4150);
nor U10295 (N_10295,N_3235,N_1864);
nand U10296 (N_10296,N_5676,N_247);
nand U10297 (N_10297,N_4826,N_2562);
and U10298 (N_10298,N_4261,N_4770);
nor U10299 (N_10299,N_1401,N_3720);
nor U10300 (N_10300,N_469,N_3512);
nor U10301 (N_10301,N_5514,N_3973);
nor U10302 (N_10302,N_3912,N_5789);
or U10303 (N_10303,N_3956,N_1288);
and U10304 (N_10304,N_4993,N_5146);
nand U10305 (N_10305,N_318,N_1434);
and U10306 (N_10306,N_2937,N_3989);
nand U10307 (N_10307,N_2875,N_4555);
or U10308 (N_10308,N_599,N_4961);
or U10309 (N_10309,N_3648,N_5989);
or U10310 (N_10310,N_3143,N_4847);
nand U10311 (N_10311,N_4807,N_1065);
nor U10312 (N_10312,N_5211,N_4442);
and U10313 (N_10313,N_99,N_2344);
xor U10314 (N_10314,N_4761,N_1691);
nand U10315 (N_10315,N_3048,N_347);
xor U10316 (N_10316,N_3943,N_559);
nor U10317 (N_10317,N_5096,N_1806);
xnor U10318 (N_10318,N_1174,N_776);
or U10319 (N_10319,N_2755,N_3810);
xor U10320 (N_10320,N_5179,N_315);
nor U10321 (N_10321,N_4210,N_5990);
or U10322 (N_10322,N_169,N_2326);
and U10323 (N_10323,N_1705,N_4910);
and U10324 (N_10324,N_3826,N_4637);
nor U10325 (N_10325,N_5650,N_1576);
nand U10326 (N_10326,N_3503,N_726);
or U10327 (N_10327,N_4504,N_4206);
nand U10328 (N_10328,N_300,N_1680);
and U10329 (N_10329,N_5981,N_1559);
or U10330 (N_10330,N_5035,N_542);
nor U10331 (N_10331,N_4177,N_2924);
or U10332 (N_10332,N_2466,N_589);
and U10333 (N_10333,N_2115,N_508);
or U10334 (N_10334,N_1965,N_1583);
nor U10335 (N_10335,N_4750,N_3371);
nand U10336 (N_10336,N_3532,N_2167);
and U10337 (N_10337,N_4428,N_1723);
nand U10338 (N_10338,N_1134,N_3631);
nand U10339 (N_10339,N_5389,N_5528);
and U10340 (N_10340,N_3612,N_4406);
xor U10341 (N_10341,N_3299,N_1462);
nand U10342 (N_10342,N_5084,N_5965);
nand U10343 (N_10343,N_4344,N_4466);
or U10344 (N_10344,N_211,N_2045);
nor U10345 (N_10345,N_3345,N_5950);
nand U10346 (N_10346,N_5613,N_1940);
nor U10347 (N_10347,N_252,N_2946);
nor U10348 (N_10348,N_3362,N_3694);
or U10349 (N_10349,N_5948,N_1382);
nor U10350 (N_10350,N_3705,N_1762);
nor U10351 (N_10351,N_15,N_3675);
nor U10352 (N_10352,N_356,N_2779);
and U10353 (N_10353,N_652,N_4044);
and U10354 (N_10354,N_616,N_3780);
nor U10355 (N_10355,N_1054,N_2339);
nor U10356 (N_10356,N_5935,N_1182);
nand U10357 (N_10357,N_4975,N_3286);
or U10358 (N_10358,N_1008,N_5772);
and U10359 (N_10359,N_3072,N_5570);
nand U10360 (N_10360,N_184,N_5054);
or U10361 (N_10361,N_1172,N_5684);
or U10362 (N_10362,N_1825,N_315);
nor U10363 (N_10363,N_5098,N_3448);
xnor U10364 (N_10364,N_5142,N_2031);
nand U10365 (N_10365,N_1274,N_1483);
nor U10366 (N_10366,N_1040,N_3923);
nand U10367 (N_10367,N_2270,N_1390);
and U10368 (N_10368,N_2029,N_2831);
nand U10369 (N_10369,N_75,N_478);
or U10370 (N_10370,N_28,N_898);
nor U10371 (N_10371,N_3599,N_1867);
nand U10372 (N_10372,N_1035,N_2937);
nor U10373 (N_10373,N_2606,N_1921);
nor U10374 (N_10374,N_3386,N_163);
or U10375 (N_10375,N_2637,N_2744);
nor U10376 (N_10376,N_618,N_3936);
and U10377 (N_10377,N_3935,N_4701);
or U10378 (N_10378,N_4167,N_3252);
nand U10379 (N_10379,N_1819,N_3718);
nand U10380 (N_10380,N_4802,N_5987);
nor U10381 (N_10381,N_2484,N_919);
or U10382 (N_10382,N_3525,N_2667);
and U10383 (N_10383,N_2933,N_422);
nor U10384 (N_10384,N_1107,N_44);
nor U10385 (N_10385,N_1061,N_1212);
and U10386 (N_10386,N_1488,N_989);
or U10387 (N_10387,N_1373,N_2143);
nand U10388 (N_10388,N_4748,N_2944);
or U10389 (N_10389,N_1455,N_1139);
nand U10390 (N_10390,N_4393,N_4960);
or U10391 (N_10391,N_1800,N_4923);
and U10392 (N_10392,N_5167,N_3606);
nand U10393 (N_10393,N_774,N_2776);
or U10394 (N_10394,N_3361,N_4988);
and U10395 (N_10395,N_1419,N_3431);
nor U10396 (N_10396,N_2117,N_4472);
and U10397 (N_10397,N_1161,N_1459);
nor U10398 (N_10398,N_8,N_4593);
nand U10399 (N_10399,N_2491,N_5771);
nor U10400 (N_10400,N_4479,N_70);
nor U10401 (N_10401,N_4359,N_5103);
nand U10402 (N_10402,N_1478,N_4087);
and U10403 (N_10403,N_4865,N_880);
nand U10404 (N_10404,N_5085,N_5874);
or U10405 (N_10405,N_3742,N_1265);
and U10406 (N_10406,N_382,N_2865);
or U10407 (N_10407,N_642,N_4551);
nand U10408 (N_10408,N_3177,N_3745);
nand U10409 (N_10409,N_4173,N_2011);
nand U10410 (N_10410,N_1349,N_3798);
nor U10411 (N_10411,N_4012,N_173);
nand U10412 (N_10412,N_3046,N_4515);
or U10413 (N_10413,N_5392,N_5493);
or U10414 (N_10414,N_5475,N_1252);
nand U10415 (N_10415,N_1205,N_5336);
xor U10416 (N_10416,N_4185,N_247);
nor U10417 (N_10417,N_3678,N_3024);
and U10418 (N_10418,N_696,N_3508);
or U10419 (N_10419,N_1686,N_4889);
or U10420 (N_10420,N_1759,N_5975);
nor U10421 (N_10421,N_680,N_3609);
or U10422 (N_10422,N_3045,N_5340);
nor U10423 (N_10423,N_3965,N_3945);
nand U10424 (N_10424,N_3902,N_5372);
or U10425 (N_10425,N_3990,N_5913);
nand U10426 (N_10426,N_2240,N_4114);
xor U10427 (N_10427,N_5202,N_842);
nor U10428 (N_10428,N_3472,N_80);
or U10429 (N_10429,N_1133,N_5437);
nand U10430 (N_10430,N_3815,N_1533);
xnor U10431 (N_10431,N_3358,N_4450);
or U10432 (N_10432,N_3496,N_5224);
and U10433 (N_10433,N_4526,N_4634);
xor U10434 (N_10434,N_5677,N_513);
and U10435 (N_10435,N_5084,N_4118);
or U10436 (N_10436,N_3674,N_1116);
nand U10437 (N_10437,N_4771,N_837);
nor U10438 (N_10438,N_5126,N_1429);
or U10439 (N_10439,N_88,N_2387);
xnor U10440 (N_10440,N_1363,N_2246);
nand U10441 (N_10441,N_2819,N_5287);
nand U10442 (N_10442,N_142,N_1913);
xnor U10443 (N_10443,N_3046,N_2763);
and U10444 (N_10444,N_5200,N_4756);
xor U10445 (N_10445,N_5008,N_4882);
nor U10446 (N_10446,N_4596,N_5317);
and U10447 (N_10447,N_811,N_3467);
or U10448 (N_10448,N_94,N_2977);
and U10449 (N_10449,N_4107,N_3314);
nor U10450 (N_10450,N_2288,N_1315);
and U10451 (N_10451,N_1612,N_2034);
and U10452 (N_10452,N_143,N_3253);
nor U10453 (N_10453,N_5918,N_5027);
xor U10454 (N_10454,N_4597,N_1747);
or U10455 (N_10455,N_4680,N_3135);
or U10456 (N_10456,N_755,N_4617);
or U10457 (N_10457,N_4529,N_1552);
nor U10458 (N_10458,N_895,N_856);
nand U10459 (N_10459,N_2029,N_5980);
xor U10460 (N_10460,N_4030,N_1681);
and U10461 (N_10461,N_5855,N_2324);
nand U10462 (N_10462,N_5109,N_344);
and U10463 (N_10463,N_5810,N_3276);
or U10464 (N_10464,N_1973,N_384);
nor U10465 (N_10465,N_3769,N_892);
nand U10466 (N_10466,N_4422,N_5118);
and U10467 (N_10467,N_2872,N_4594);
or U10468 (N_10468,N_169,N_3834);
and U10469 (N_10469,N_4537,N_2342);
or U10470 (N_10470,N_2560,N_103);
nor U10471 (N_10471,N_1566,N_1147);
nor U10472 (N_10472,N_369,N_3638);
nor U10473 (N_10473,N_3586,N_3380);
or U10474 (N_10474,N_1653,N_2642);
or U10475 (N_10475,N_5854,N_4878);
nor U10476 (N_10476,N_1519,N_105);
nand U10477 (N_10477,N_289,N_2518);
nand U10478 (N_10478,N_3575,N_3530);
or U10479 (N_10479,N_4572,N_1620);
nor U10480 (N_10480,N_5651,N_1119);
or U10481 (N_10481,N_4511,N_2864);
and U10482 (N_10482,N_2809,N_1907);
and U10483 (N_10483,N_4081,N_1930);
or U10484 (N_10484,N_974,N_2855);
nand U10485 (N_10485,N_1842,N_4426);
and U10486 (N_10486,N_1162,N_3753);
nand U10487 (N_10487,N_5148,N_1323);
xnor U10488 (N_10488,N_184,N_1439);
or U10489 (N_10489,N_5219,N_3467);
nor U10490 (N_10490,N_3811,N_5033);
and U10491 (N_10491,N_1005,N_1148);
or U10492 (N_10492,N_419,N_1529);
and U10493 (N_10493,N_2116,N_830);
nand U10494 (N_10494,N_588,N_2820);
or U10495 (N_10495,N_3778,N_3908);
and U10496 (N_10496,N_235,N_4182);
and U10497 (N_10497,N_2975,N_1798);
nand U10498 (N_10498,N_1969,N_1700);
and U10499 (N_10499,N_2485,N_5463);
or U10500 (N_10500,N_1400,N_55);
nand U10501 (N_10501,N_4996,N_1786);
or U10502 (N_10502,N_3972,N_4963);
and U10503 (N_10503,N_1815,N_4962);
nand U10504 (N_10504,N_5290,N_5243);
xnor U10505 (N_10505,N_3679,N_3196);
nor U10506 (N_10506,N_1621,N_4897);
and U10507 (N_10507,N_4633,N_5877);
or U10508 (N_10508,N_3584,N_3908);
and U10509 (N_10509,N_4101,N_5186);
and U10510 (N_10510,N_2720,N_5783);
and U10511 (N_10511,N_888,N_4612);
nor U10512 (N_10512,N_2067,N_2751);
or U10513 (N_10513,N_4399,N_872);
or U10514 (N_10514,N_3124,N_569);
xnor U10515 (N_10515,N_3268,N_1592);
nor U10516 (N_10516,N_4261,N_539);
or U10517 (N_10517,N_522,N_612);
nand U10518 (N_10518,N_2700,N_4467);
nand U10519 (N_10519,N_4804,N_888);
xnor U10520 (N_10520,N_4141,N_5955);
or U10521 (N_10521,N_5503,N_443);
nor U10522 (N_10522,N_4038,N_919);
nor U10523 (N_10523,N_4319,N_5233);
xor U10524 (N_10524,N_1518,N_4998);
and U10525 (N_10525,N_1259,N_3868);
nand U10526 (N_10526,N_1931,N_862);
nor U10527 (N_10527,N_3692,N_3772);
nand U10528 (N_10528,N_506,N_793);
nor U10529 (N_10529,N_944,N_3278);
nor U10530 (N_10530,N_62,N_74);
nor U10531 (N_10531,N_28,N_3960);
and U10532 (N_10532,N_2051,N_2015);
nor U10533 (N_10533,N_2679,N_104);
and U10534 (N_10534,N_3569,N_5551);
and U10535 (N_10535,N_1855,N_4177);
nand U10536 (N_10536,N_5184,N_4361);
and U10537 (N_10537,N_644,N_875);
and U10538 (N_10538,N_1001,N_2611);
nor U10539 (N_10539,N_2540,N_769);
nor U10540 (N_10540,N_1875,N_4122);
or U10541 (N_10541,N_3306,N_690);
nand U10542 (N_10542,N_4374,N_1217);
xnor U10543 (N_10543,N_3300,N_4636);
or U10544 (N_10544,N_3632,N_3920);
nand U10545 (N_10545,N_2164,N_5371);
nor U10546 (N_10546,N_404,N_3725);
nand U10547 (N_10547,N_1734,N_1409);
nand U10548 (N_10548,N_2658,N_759);
and U10549 (N_10549,N_4647,N_5603);
and U10550 (N_10550,N_3804,N_1362);
nand U10551 (N_10551,N_5674,N_4985);
and U10552 (N_10552,N_1392,N_2459);
nand U10553 (N_10553,N_2321,N_4469);
nor U10554 (N_10554,N_2910,N_4322);
nand U10555 (N_10555,N_154,N_4096);
nand U10556 (N_10556,N_1602,N_4701);
and U10557 (N_10557,N_4990,N_3227);
xor U10558 (N_10558,N_5803,N_1849);
xnor U10559 (N_10559,N_1840,N_1157);
nor U10560 (N_10560,N_2198,N_3630);
nand U10561 (N_10561,N_1681,N_4437);
or U10562 (N_10562,N_4462,N_3031);
nand U10563 (N_10563,N_5158,N_1893);
or U10564 (N_10564,N_5932,N_1043);
nor U10565 (N_10565,N_2342,N_5228);
nand U10566 (N_10566,N_1923,N_5568);
nand U10567 (N_10567,N_919,N_3639);
nor U10568 (N_10568,N_783,N_1174);
nor U10569 (N_10569,N_5671,N_2986);
or U10570 (N_10570,N_2228,N_3351);
nand U10571 (N_10571,N_1526,N_3144);
and U10572 (N_10572,N_604,N_819);
nand U10573 (N_10573,N_1248,N_3306);
nand U10574 (N_10574,N_5682,N_521);
and U10575 (N_10575,N_292,N_1288);
and U10576 (N_10576,N_3595,N_737);
nand U10577 (N_10577,N_5186,N_5794);
nand U10578 (N_10578,N_3968,N_2354);
nor U10579 (N_10579,N_2570,N_3147);
nand U10580 (N_10580,N_2850,N_2015);
and U10581 (N_10581,N_3258,N_2974);
nand U10582 (N_10582,N_4157,N_5556);
and U10583 (N_10583,N_5029,N_5474);
and U10584 (N_10584,N_5713,N_4174);
nand U10585 (N_10585,N_4023,N_4570);
nand U10586 (N_10586,N_1741,N_3061);
nor U10587 (N_10587,N_4467,N_3262);
or U10588 (N_10588,N_3715,N_4831);
nand U10589 (N_10589,N_1104,N_708);
or U10590 (N_10590,N_1839,N_823);
nand U10591 (N_10591,N_2464,N_524);
or U10592 (N_10592,N_2014,N_2675);
nand U10593 (N_10593,N_5107,N_2330);
nand U10594 (N_10594,N_5284,N_5613);
and U10595 (N_10595,N_4354,N_3891);
and U10596 (N_10596,N_3981,N_3497);
and U10597 (N_10597,N_3873,N_2429);
and U10598 (N_10598,N_1148,N_1149);
or U10599 (N_10599,N_3962,N_2090);
or U10600 (N_10600,N_5467,N_2073);
nand U10601 (N_10601,N_98,N_827);
and U10602 (N_10602,N_448,N_3258);
and U10603 (N_10603,N_3566,N_94);
and U10604 (N_10604,N_782,N_162);
and U10605 (N_10605,N_3890,N_1825);
or U10606 (N_10606,N_4480,N_2282);
and U10607 (N_10607,N_1012,N_5838);
nand U10608 (N_10608,N_3347,N_606);
nor U10609 (N_10609,N_3790,N_0);
nand U10610 (N_10610,N_3720,N_3575);
nand U10611 (N_10611,N_5544,N_1667);
and U10612 (N_10612,N_3875,N_2955);
nand U10613 (N_10613,N_151,N_2800);
nand U10614 (N_10614,N_5560,N_4441);
nand U10615 (N_10615,N_5200,N_4267);
and U10616 (N_10616,N_3392,N_5451);
nor U10617 (N_10617,N_2617,N_4838);
xnor U10618 (N_10618,N_1938,N_4055);
and U10619 (N_10619,N_1484,N_5114);
nor U10620 (N_10620,N_4870,N_5648);
nand U10621 (N_10621,N_4136,N_646);
or U10622 (N_10622,N_5903,N_4064);
nor U10623 (N_10623,N_4887,N_1095);
nand U10624 (N_10624,N_2399,N_5382);
or U10625 (N_10625,N_4736,N_5285);
nor U10626 (N_10626,N_4193,N_3253);
nand U10627 (N_10627,N_3334,N_4047);
and U10628 (N_10628,N_1710,N_809);
and U10629 (N_10629,N_4639,N_5214);
or U10630 (N_10630,N_3446,N_3335);
nor U10631 (N_10631,N_4137,N_3529);
and U10632 (N_10632,N_263,N_1628);
xnor U10633 (N_10633,N_2110,N_4300);
nor U10634 (N_10634,N_601,N_184);
nor U10635 (N_10635,N_2649,N_1268);
nor U10636 (N_10636,N_3207,N_2390);
nand U10637 (N_10637,N_2218,N_5352);
nor U10638 (N_10638,N_861,N_3877);
nor U10639 (N_10639,N_815,N_1242);
nand U10640 (N_10640,N_1530,N_2463);
nor U10641 (N_10641,N_1587,N_91);
and U10642 (N_10642,N_4342,N_4664);
xnor U10643 (N_10643,N_137,N_4043);
nand U10644 (N_10644,N_4324,N_3211);
or U10645 (N_10645,N_4763,N_5884);
nor U10646 (N_10646,N_5174,N_597);
nand U10647 (N_10647,N_4357,N_880);
xor U10648 (N_10648,N_2642,N_416);
nor U10649 (N_10649,N_3429,N_5712);
and U10650 (N_10650,N_3353,N_2417);
or U10651 (N_10651,N_1124,N_4904);
nor U10652 (N_10652,N_1647,N_1750);
nor U10653 (N_10653,N_1862,N_4286);
nor U10654 (N_10654,N_5429,N_3076);
xnor U10655 (N_10655,N_110,N_1613);
xor U10656 (N_10656,N_3962,N_5483);
or U10657 (N_10657,N_28,N_4781);
nand U10658 (N_10658,N_5066,N_1957);
nand U10659 (N_10659,N_1540,N_2161);
or U10660 (N_10660,N_4239,N_5853);
or U10661 (N_10661,N_3178,N_1376);
nor U10662 (N_10662,N_4,N_3271);
nor U10663 (N_10663,N_4230,N_1262);
nand U10664 (N_10664,N_926,N_4688);
and U10665 (N_10665,N_3711,N_2608);
or U10666 (N_10666,N_4936,N_709);
nand U10667 (N_10667,N_4780,N_5894);
nand U10668 (N_10668,N_2571,N_2499);
and U10669 (N_10669,N_3335,N_5828);
or U10670 (N_10670,N_5819,N_363);
nor U10671 (N_10671,N_417,N_2853);
nand U10672 (N_10672,N_603,N_2280);
nand U10673 (N_10673,N_5969,N_4590);
nor U10674 (N_10674,N_4578,N_1967);
nor U10675 (N_10675,N_2881,N_3111);
nand U10676 (N_10676,N_3169,N_1238);
or U10677 (N_10677,N_377,N_4779);
or U10678 (N_10678,N_2616,N_1558);
nor U10679 (N_10679,N_3465,N_1504);
xnor U10680 (N_10680,N_1781,N_2850);
or U10681 (N_10681,N_5267,N_2917);
nor U10682 (N_10682,N_77,N_3290);
and U10683 (N_10683,N_5944,N_1114);
and U10684 (N_10684,N_1400,N_580);
nor U10685 (N_10685,N_3720,N_1374);
nand U10686 (N_10686,N_2736,N_4997);
nor U10687 (N_10687,N_4125,N_5502);
nor U10688 (N_10688,N_4885,N_3376);
or U10689 (N_10689,N_700,N_3147);
and U10690 (N_10690,N_731,N_3701);
nor U10691 (N_10691,N_3202,N_1740);
nor U10692 (N_10692,N_5760,N_1149);
nor U10693 (N_10693,N_1311,N_4711);
and U10694 (N_10694,N_5045,N_3333);
nor U10695 (N_10695,N_1592,N_1688);
and U10696 (N_10696,N_3281,N_1677);
or U10697 (N_10697,N_2559,N_1229);
nor U10698 (N_10698,N_1303,N_3144);
and U10699 (N_10699,N_1866,N_3637);
nand U10700 (N_10700,N_3277,N_2685);
or U10701 (N_10701,N_1782,N_812);
and U10702 (N_10702,N_2455,N_5383);
nand U10703 (N_10703,N_274,N_2096);
or U10704 (N_10704,N_5228,N_2411);
nand U10705 (N_10705,N_1191,N_2194);
nor U10706 (N_10706,N_4963,N_803);
xor U10707 (N_10707,N_3038,N_4864);
or U10708 (N_10708,N_5808,N_35);
xnor U10709 (N_10709,N_1416,N_3570);
nor U10710 (N_10710,N_3397,N_555);
or U10711 (N_10711,N_5298,N_5608);
nor U10712 (N_10712,N_4501,N_4036);
xnor U10713 (N_10713,N_4782,N_121);
or U10714 (N_10714,N_2089,N_5404);
or U10715 (N_10715,N_2648,N_1140);
nor U10716 (N_10716,N_4910,N_229);
xor U10717 (N_10717,N_1020,N_5931);
nor U10718 (N_10718,N_1861,N_1757);
or U10719 (N_10719,N_5716,N_4055);
xor U10720 (N_10720,N_1471,N_3140);
nor U10721 (N_10721,N_4671,N_808);
or U10722 (N_10722,N_5303,N_143);
and U10723 (N_10723,N_2291,N_4906);
nor U10724 (N_10724,N_732,N_4368);
or U10725 (N_10725,N_581,N_2518);
xnor U10726 (N_10726,N_1273,N_3504);
nand U10727 (N_10727,N_2750,N_453);
and U10728 (N_10728,N_1730,N_2843);
xor U10729 (N_10729,N_1834,N_2220);
and U10730 (N_10730,N_1830,N_3980);
or U10731 (N_10731,N_2792,N_2989);
nand U10732 (N_10732,N_1818,N_5612);
nor U10733 (N_10733,N_2388,N_5641);
xor U10734 (N_10734,N_5685,N_5596);
nor U10735 (N_10735,N_5009,N_5011);
xnor U10736 (N_10736,N_995,N_3730);
xor U10737 (N_10737,N_364,N_2720);
or U10738 (N_10738,N_3668,N_4328);
nor U10739 (N_10739,N_2458,N_4146);
nand U10740 (N_10740,N_551,N_2943);
nor U10741 (N_10741,N_5528,N_5641);
nand U10742 (N_10742,N_3667,N_4451);
and U10743 (N_10743,N_3014,N_5220);
nor U10744 (N_10744,N_1011,N_5069);
nand U10745 (N_10745,N_5354,N_5800);
nor U10746 (N_10746,N_264,N_2979);
nand U10747 (N_10747,N_1937,N_4985);
xor U10748 (N_10748,N_5426,N_2463);
nand U10749 (N_10749,N_4442,N_70);
and U10750 (N_10750,N_5283,N_1522);
nand U10751 (N_10751,N_3448,N_692);
xnor U10752 (N_10752,N_4485,N_5785);
and U10753 (N_10753,N_5866,N_3681);
nand U10754 (N_10754,N_3292,N_456);
or U10755 (N_10755,N_1037,N_63);
nand U10756 (N_10756,N_5849,N_4036);
nand U10757 (N_10757,N_81,N_695);
and U10758 (N_10758,N_610,N_5886);
and U10759 (N_10759,N_5069,N_4808);
and U10760 (N_10760,N_3611,N_1506);
or U10761 (N_10761,N_1345,N_3146);
and U10762 (N_10762,N_5602,N_3019);
xnor U10763 (N_10763,N_310,N_4700);
or U10764 (N_10764,N_123,N_4820);
or U10765 (N_10765,N_5425,N_5626);
or U10766 (N_10766,N_4238,N_5311);
or U10767 (N_10767,N_1768,N_1296);
nor U10768 (N_10768,N_5143,N_2833);
nor U10769 (N_10769,N_700,N_5783);
nand U10770 (N_10770,N_4011,N_5880);
nand U10771 (N_10771,N_5315,N_1226);
and U10772 (N_10772,N_3614,N_155);
xnor U10773 (N_10773,N_4793,N_2843);
nand U10774 (N_10774,N_1034,N_4686);
and U10775 (N_10775,N_5288,N_3059);
and U10776 (N_10776,N_5865,N_5034);
nand U10777 (N_10777,N_679,N_5156);
or U10778 (N_10778,N_5923,N_5410);
xnor U10779 (N_10779,N_4926,N_961);
nor U10780 (N_10780,N_4571,N_4907);
nor U10781 (N_10781,N_1436,N_3002);
or U10782 (N_10782,N_1279,N_4413);
nand U10783 (N_10783,N_3069,N_3969);
xor U10784 (N_10784,N_2394,N_4022);
xnor U10785 (N_10785,N_437,N_1162);
nor U10786 (N_10786,N_2812,N_2170);
nand U10787 (N_10787,N_5127,N_4063);
nand U10788 (N_10788,N_5543,N_3600);
and U10789 (N_10789,N_3839,N_2703);
xor U10790 (N_10790,N_3767,N_3060);
or U10791 (N_10791,N_4912,N_3601);
or U10792 (N_10792,N_4149,N_1935);
xor U10793 (N_10793,N_4814,N_4423);
nand U10794 (N_10794,N_445,N_657);
xnor U10795 (N_10795,N_5884,N_558);
nand U10796 (N_10796,N_5323,N_282);
nand U10797 (N_10797,N_2015,N_4429);
nand U10798 (N_10798,N_4718,N_4101);
or U10799 (N_10799,N_1736,N_2744);
and U10800 (N_10800,N_1576,N_762);
or U10801 (N_10801,N_2436,N_930);
nor U10802 (N_10802,N_5050,N_4499);
or U10803 (N_10803,N_3096,N_4949);
xnor U10804 (N_10804,N_5186,N_3706);
or U10805 (N_10805,N_4261,N_460);
or U10806 (N_10806,N_208,N_3952);
or U10807 (N_10807,N_5984,N_5376);
nor U10808 (N_10808,N_4705,N_4487);
nand U10809 (N_10809,N_3235,N_5257);
and U10810 (N_10810,N_5118,N_3480);
or U10811 (N_10811,N_5076,N_62);
nor U10812 (N_10812,N_4440,N_4929);
and U10813 (N_10813,N_276,N_1814);
nor U10814 (N_10814,N_2771,N_4551);
or U10815 (N_10815,N_2123,N_5897);
nor U10816 (N_10816,N_4773,N_1310);
or U10817 (N_10817,N_1513,N_2394);
nand U10818 (N_10818,N_672,N_3284);
nand U10819 (N_10819,N_2861,N_753);
nand U10820 (N_10820,N_609,N_1525);
nand U10821 (N_10821,N_4342,N_2091);
and U10822 (N_10822,N_4642,N_2182);
nand U10823 (N_10823,N_3149,N_3279);
xor U10824 (N_10824,N_4057,N_3164);
xnor U10825 (N_10825,N_3463,N_1921);
and U10826 (N_10826,N_1013,N_568);
nor U10827 (N_10827,N_1097,N_865);
nand U10828 (N_10828,N_3855,N_3630);
nor U10829 (N_10829,N_5350,N_604);
xnor U10830 (N_10830,N_2146,N_3628);
or U10831 (N_10831,N_2758,N_2966);
xor U10832 (N_10832,N_3910,N_3101);
nor U10833 (N_10833,N_807,N_3189);
xnor U10834 (N_10834,N_4161,N_2780);
or U10835 (N_10835,N_4895,N_5488);
nor U10836 (N_10836,N_0,N_3191);
or U10837 (N_10837,N_4492,N_3005);
or U10838 (N_10838,N_1394,N_887);
nand U10839 (N_10839,N_2444,N_5066);
or U10840 (N_10840,N_5346,N_490);
nand U10841 (N_10841,N_3451,N_4672);
or U10842 (N_10842,N_2026,N_3432);
or U10843 (N_10843,N_5419,N_4536);
nor U10844 (N_10844,N_1120,N_2118);
nor U10845 (N_10845,N_1616,N_3980);
nand U10846 (N_10846,N_4819,N_62);
nand U10847 (N_10847,N_5344,N_4811);
or U10848 (N_10848,N_4506,N_1052);
nand U10849 (N_10849,N_2637,N_4796);
nor U10850 (N_10850,N_1086,N_4620);
or U10851 (N_10851,N_2289,N_1300);
or U10852 (N_10852,N_4075,N_742);
nand U10853 (N_10853,N_4553,N_1720);
nor U10854 (N_10854,N_852,N_718);
nor U10855 (N_10855,N_5567,N_2609);
and U10856 (N_10856,N_1514,N_4907);
or U10857 (N_10857,N_2655,N_4625);
xnor U10858 (N_10858,N_5869,N_1450);
nand U10859 (N_10859,N_4709,N_634);
nor U10860 (N_10860,N_1045,N_3853);
nand U10861 (N_10861,N_1839,N_4968);
nand U10862 (N_10862,N_2101,N_4865);
nor U10863 (N_10863,N_3823,N_50);
or U10864 (N_10864,N_3312,N_2731);
or U10865 (N_10865,N_4745,N_4085);
or U10866 (N_10866,N_3056,N_3589);
nand U10867 (N_10867,N_297,N_3159);
nand U10868 (N_10868,N_4936,N_3674);
xnor U10869 (N_10869,N_4176,N_4566);
nor U10870 (N_10870,N_5140,N_682);
or U10871 (N_10871,N_3568,N_3216);
nand U10872 (N_10872,N_2544,N_5693);
and U10873 (N_10873,N_133,N_2788);
xnor U10874 (N_10874,N_3030,N_769);
nand U10875 (N_10875,N_4451,N_2111);
or U10876 (N_10876,N_5096,N_664);
and U10877 (N_10877,N_2061,N_3887);
or U10878 (N_10878,N_1307,N_5304);
or U10879 (N_10879,N_1664,N_1417);
nor U10880 (N_10880,N_5845,N_2068);
and U10881 (N_10881,N_5040,N_5955);
xnor U10882 (N_10882,N_5595,N_5063);
or U10883 (N_10883,N_5243,N_3352);
nand U10884 (N_10884,N_3015,N_1894);
nand U10885 (N_10885,N_1795,N_2183);
nand U10886 (N_10886,N_4134,N_4069);
or U10887 (N_10887,N_3118,N_230);
nor U10888 (N_10888,N_3532,N_5518);
nand U10889 (N_10889,N_5647,N_2729);
nor U10890 (N_10890,N_1878,N_1117);
or U10891 (N_10891,N_2433,N_5607);
nand U10892 (N_10892,N_1860,N_3470);
or U10893 (N_10893,N_2000,N_535);
and U10894 (N_10894,N_1040,N_1330);
nand U10895 (N_10895,N_4109,N_4940);
nand U10896 (N_10896,N_5675,N_4862);
or U10897 (N_10897,N_3778,N_3347);
nand U10898 (N_10898,N_2856,N_537);
nor U10899 (N_10899,N_1872,N_4041);
xnor U10900 (N_10900,N_5859,N_4074);
nand U10901 (N_10901,N_4852,N_4838);
nor U10902 (N_10902,N_1088,N_4873);
or U10903 (N_10903,N_361,N_4486);
nand U10904 (N_10904,N_4824,N_1762);
and U10905 (N_10905,N_5907,N_4154);
xnor U10906 (N_10906,N_4222,N_5217);
nand U10907 (N_10907,N_4229,N_2344);
and U10908 (N_10908,N_1073,N_3116);
or U10909 (N_10909,N_2565,N_775);
nor U10910 (N_10910,N_2484,N_4828);
nand U10911 (N_10911,N_373,N_5293);
and U10912 (N_10912,N_5536,N_3005);
nand U10913 (N_10913,N_300,N_3661);
nor U10914 (N_10914,N_3696,N_2459);
nor U10915 (N_10915,N_252,N_55);
and U10916 (N_10916,N_2819,N_3832);
nor U10917 (N_10917,N_4445,N_2864);
xor U10918 (N_10918,N_2699,N_3326);
nand U10919 (N_10919,N_1016,N_5598);
nor U10920 (N_10920,N_5705,N_112);
nor U10921 (N_10921,N_1945,N_5688);
xor U10922 (N_10922,N_5199,N_5034);
or U10923 (N_10923,N_214,N_5514);
nor U10924 (N_10924,N_3655,N_3899);
nand U10925 (N_10925,N_205,N_3302);
nor U10926 (N_10926,N_1673,N_494);
or U10927 (N_10927,N_821,N_3232);
nor U10928 (N_10928,N_1762,N_3086);
or U10929 (N_10929,N_2113,N_22);
and U10930 (N_10930,N_2679,N_633);
or U10931 (N_10931,N_4355,N_5103);
and U10932 (N_10932,N_1353,N_2540);
nor U10933 (N_10933,N_3155,N_1225);
nand U10934 (N_10934,N_2693,N_3964);
and U10935 (N_10935,N_4915,N_1615);
xnor U10936 (N_10936,N_379,N_4134);
xor U10937 (N_10937,N_2249,N_2218);
and U10938 (N_10938,N_124,N_5280);
nand U10939 (N_10939,N_5027,N_2781);
nand U10940 (N_10940,N_1215,N_637);
or U10941 (N_10941,N_5003,N_5837);
nor U10942 (N_10942,N_5446,N_982);
and U10943 (N_10943,N_4235,N_693);
and U10944 (N_10944,N_1179,N_2735);
nor U10945 (N_10945,N_3627,N_5130);
xor U10946 (N_10946,N_4241,N_3159);
nor U10947 (N_10947,N_2948,N_3190);
nand U10948 (N_10948,N_5197,N_5410);
and U10949 (N_10949,N_840,N_4494);
and U10950 (N_10950,N_5161,N_1017);
and U10951 (N_10951,N_3894,N_2202);
and U10952 (N_10952,N_708,N_2741);
nor U10953 (N_10953,N_5437,N_64);
and U10954 (N_10954,N_1523,N_5124);
nand U10955 (N_10955,N_5551,N_5539);
nand U10956 (N_10956,N_2366,N_5770);
nand U10957 (N_10957,N_3535,N_5048);
nand U10958 (N_10958,N_3010,N_1332);
and U10959 (N_10959,N_4994,N_3921);
and U10960 (N_10960,N_3381,N_2170);
xnor U10961 (N_10961,N_1254,N_3963);
nand U10962 (N_10962,N_4213,N_1542);
and U10963 (N_10963,N_426,N_3711);
nor U10964 (N_10964,N_275,N_3378);
nand U10965 (N_10965,N_1402,N_4487);
nor U10966 (N_10966,N_2834,N_5739);
or U10967 (N_10967,N_3795,N_2772);
and U10968 (N_10968,N_870,N_2845);
nand U10969 (N_10969,N_5559,N_5775);
nor U10970 (N_10970,N_5346,N_1936);
and U10971 (N_10971,N_5851,N_1061);
nand U10972 (N_10972,N_3207,N_4290);
nor U10973 (N_10973,N_1842,N_3507);
nor U10974 (N_10974,N_2485,N_1712);
nor U10975 (N_10975,N_4902,N_4839);
nand U10976 (N_10976,N_2528,N_4999);
and U10977 (N_10977,N_380,N_4103);
and U10978 (N_10978,N_347,N_1452);
nor U10979 (N_10979,N_5470,N_3161);
or U10980 (N_10980,N_4748,N_3759);
and U10981 (N_10981,N_816,N_803);
and U10982 (N_10982,N_712,N_26);
nor U10983 (N_10983,N_4696,N_4925);
nand U10984 (N_10984,N_530,N_1185);
nor U10985 (N_10985,N_2324,N_372);
xor U10986 (N_10986,N_4819,N_5575);
or U10987 (N_10987,N_4688,N_3777);
and U10988 (N_10988,N_2743,N_2012);
or U10989 (N_10989,N_288,N_5100);
nor U10990 (N_10990,N_325,N_2923);
nor U10991 (N_10991,N_1925,N_3120);
xnor U10992 (N_10992,N_5509,N_5343);
and U10993 (N_10993,N_364,N_2331);
and U10994 (N_10994,N_1703,N_494);
nand U10995 (N_10995,N_4502,N_5116);
and U10996 (N_10996,N_677,N_2809);
nor U10997 (N_10997,N_2969,N_4702);
or U10998 (N_10998,N_5878,N_3341);
nand U10999 (N_10999,N_2923,N_3463);
or U11000 (N_11000,N_1796,N_2062);
nand U11001 (N_11001,N_4931,N_4305);
nand U11002 (N_11002,N_5182,N_3775);
and U11003 (N_11003,N_3249,N_5086);
nor U11004 (N_11004,N_3754,N_5969);
nor U11005 (N_11005,N_5899,N_4526);
nor U11006 (N_11006,N_5044,N_565);
nor U11007 (N_11007,N_1854,N_404);
and U11008 (N_11008,N_3601,N_4162);
and U11009 (N_11009,N_1406,N_1183);
and U11010 (N_11010,N_4411,N_3266);
nor U11011 (N_11011,N_257,N_5125);
nor U11012 (N_11012,N_4435,N_5116);
or U11013 (N_11013,N_254,N_5805);
nor U11014 (N_11014,N_2084,N_3907);
or U11015 (N_11015,N_2310,N_2761);
nand U11016 (N_11016,N_312,N_3564);
or U11017 (N_11017,N_2410,N_1077);
nor U11018 (N_11018,N_3065,N_1149);
nor U11019 (N_11019,N_2635,N_2331);
or U11020 (N_11020,N_5868,N_815);
nor U11021 (N_11021,N_2548,N_1154);
nor U11022 (N_11022,N_3025,N_4587);
or U11023 (N_11023,N_5660,N_3369);
or U11024 (N_11024,N_4338,N_4580);
xnor U11025 (N_11025,N_5828,N_288);
nor U11026 (N_11026,N_2789,N_1900);
xor U11027 (N_11027,N_2910,N_4715);
nand U11028 (N_11028,N_2682,N_1766);
nor U11029 (N_11029,N_2168,N_5574);
and U11030 (N_11030,N_1647,N_3352);
and U11031 (N_11031,N_2011,N_959);
and U11032 (N_11032,N_2103,N_302);
nor U11033 (N_11033,N_4559,N_106);
nand U11034 (N_11034,N_3345,N_2962);
nand U11035 (N_11035,N_432,N_5435);
or U11036 (N_11036,N_5324,N_104);
or U11037 (N_11037,N_3210,N_1766);
and U11038 (N_11038,N_4287,N_5105);
and U11039 (N_11039,N_1690,N_1458);
or U11040 (N_11040,N_1859,N_36);
nand U11041 (N_11041,N_3547,N_2683);
and U11042 (N_11042,N_579,N_395);
or U11043 (N_11043,N_3753,N_3420);
nand U11044 (N_11044,N_4330,N_639);
nand U11045 (N_11045,N_2560,N_5840);
nand U11046 (N_11046,N_2704,N_4693);
nor U11047 (N_11047,N_4771,N_458);
or U11048 (N_11048,N_5446,N_1617);
and U11049 (N_11049,N_2283,N_511);
or U11050 (N_11050,N_1973,N_3467);
or U11051 (N_11051,N_4217,N_5484);
xor U11052 (N_11052,N_5673,N_3848);
nor U11053 (N_11053,N_119,N_3618);
or U11054 (N_11054,N_5418,N_1251);
and U11055 (N_11055,N_575,N_3329);
nand U11056 (N_11056,N_2197,N_2730);
xnor U11057 (N_11057,N_3078,N_3311);
or U11058 (N_11058,N_1744,N_3742);
and U11059 (N_11059,N_3520,N_5016);
or U11060 (N_11060,N_3650,N_141);
nor U11061 (N_11061,N_1112,N_4789);
nand U11062 (N_11062,N_4328,N_2062);
nand U11063 (N_11063,N_2180,N_865);
and U11064 (N_11064,N_4795,N_938);
or U11065 (N_11065,N_2725,N_1225);
or U11066 (N_11066,N_1564,N_4050);
nand U11067 (N_11067,N_1709,N_3273);
nand U11068 (N_11068,N_20,N_2578);
and U11069 (N_11069,N_1134,N_2566);
nor U11070 (N_11070,N_118,N_4554);
and U11071 (N_11071,N_1305,N_4144);
nor U11072 (N_11072,N_3292,N_2129);
xor U11073 (N_11073,N_5232,N_4022);
and U11074 (N_11074,N_2524,N_705);
nor U11075 (N_11075,N_100,N_2298);
or U11076 (N_11076,N_5788,N_2323);
xor U11077 (N_11077,N_4846,N_1014);
nor U11078 (N_11078,N_2668,N_2132);
and U11079 (N_11079,N_4860,N_2342);
nor U11080 (N_11080,N_1403,N_2869);
and U11081 (N_11081,N_4409,N_4186);
nand U11082 (N_11082,N_5907,N_1132);
nand U11083 (N_11083,N_1261,N_745);
nor U11084 (N_11084,N_770,N_3473);
nor U11085 (N_11085,N_3379,N_5933);
nor U11086 (N_11086,N_4346,N_5370);
nor U11087 (N_11087,N_5400,N_3511);
and U11088 (N_11088,N_4398,N_1679);
xor U11089 (N_11089,N_3853,N_7);
nor U11090 (N_11090,N_5446,N_2340);
or U11091 (N_11091,N_1471,N_5635);
or U11092 (N_11092,N_3890,N_1933);
and U11093 (N_11093,N_2296,N_4596);
xnor U11094 (N_11094,N_4616,N_1825);
nand U11095 (N_11095,N_1135,N_593);
or U11096 (N_11096,N_4955,N_1876);
nor U11097 (N_11097,N_5084,N_807);
and U11098 (N_11098,N_3040,N_3795);
and U11099 (N_11099,N_2658,N_1078);
and U11100 (N_11100,N_5005,N_545);
nand U11101 (N_11101,N_2668,N_2351);
and U11102 (N_11102,N_3391,N_770);
or U11103 (N_11103,N_3023,N_5704);
nand U11104 (N_11104,N_3799,N_2742);
xor U11105 (N_11105,N_2636,N_4595);
xor U11106 (N_11106,N_87,N_5403);
nand U11107 (N_11107,N_1669,N_3635);
and U11108 (N_11108,N_5436,N_5189);
nand U11109 (N_11109,N_2933,N_5593);
or U11110 (N_11110,N_4894,N_215);
or U11111 (N_11111,N_1243,N_955);
nor U11112 (N_11112,N_4660,N_3898);
nand U11113 (N_11113,N_5674,N_618);
nor U11114 (N_11114,N_4992,N_5085);
nand U11115 (N_11115,N_1218,N_1743);
nor U11116 (N_11116,N_1912,N_1739);
or U11117 (N_11117,N_3691,N_1425);
xor U11118 (N_11118,N_3936,N_1471);
and U11119 (N_11119,N_1321,N_2871);
nand U11120 (N_11120,N_2936,N_1407);
or U11121 (N_11121,N_1565,N_5059);
and U11122 (N_11122,N_2513,N_2062);
nand U11123 (N_11123,N_2802,N_1522);
or U11124 (N_11124,N_4726,N_3852);
and U11125 (N_11125,N_2407,N_710);
or U11126 (N_11126,N_1542,N_1816);
and U11127 (N_11127,N_5002,N_4645);
or U11128 (N_11128,N_2843,N_477);
nand U11129 (N_11129,N_789,N_5887);
or U11130 (N_11130,N_1092,N_1411);
and U11131 (N_11131,N_3857,N_2114);
and U11132 (N_11132,N_5051,N_1549);
and U11133 (N_11133,N_3993,N_3059);
or U11134 (N_11134,N_1349,N_4140);
nor U11135 (N_11135,N_2048,N_3864);
and U11136 (N_11136,N_2785,N_1323);
or U11137 (N_11137,N_5849,N_1127);
and U11138 (N_11138,N_4612,N_2795);
nand U11139 (N_11139,N_1660,N_5731);
xnor U11140 (N_11140,N_1235,N_3699);
or U11141 (N_11141,N_4314,N_3190);
nor U11142 (N_11142,N_5713,N_4490);
or U11143 (N_11143,N_3692,N_84);
and U11144 (N_11144,N_2582,N_1757);
and U11145 (N_11145,N_541,N_1784);
nand U11146 (N_11146,N_5670,N_1089);
and U11147 (N_11147,N_4768,N_4680);
or U11148 (N_11148,N_433,N_997);
nand U11149 (N_11149,N_4292,N_1553);
nor U11150 (N_11150,N_4323,N_4939);
xor U11151 (N_11151,N_3200,N_1418);
xnor U11152 (N_11152,N_2025,N_2229);
nand U11153 (N_11153,N_2841,N_1487);
nor U11154 (N_11154,N_1684,N_2477);
or U11155 (N_11155,N_1432,N_925);
nor U11156 (N_11156,N_556,N_1284);
or U11157 (N_11157,N_265,N_4778);
or U11158 (N_11158,N_3276,N_3908);
or U11159 (N_11159,N_4590,N_4370);
nand U11160 (N_11160,N_1050,N_4114);
nor U11161 (N_11161,N_3021,N_3911);
nor U11162 (N_11162,N_2251,N_4704);
and U11163 (N_11163,N_5536,N_1788);
or U11164 (N_11164,N_5369,N_3474);
nand U11165 (N_11165,N_1146,N_3608);
nor U11166 (N_11166,N_5682,N_4969);
nand U11167 (N_11167,N_5910,N_3559);
nor U11168 (N_11168,N_1739,N_5279);
nand U11169 (N_11169,N_1809,N_4343);
nor U11170 (N_11170,N_4284,N_1537);
or U11171 (N_11171,N_3370,N_456);
nand U11172 (N_11172,N_1567,N_2354);
nor U11173 (N_11173,N_4304,N_1616);
nand U11174 (N_11174,N_1848,N_1203);
and U11175 (N_11175,N_5403,N_2658);
xnor U11176 (N_11176,N_4975,N_2836);
nor U11177 (N_11177,N_5696,N_4476);
and U11178 (N_11178,N_928,N_2402);
and U11179 (N_11179,N_5216,N_2540);
nand U11180 (N_11180,N_1059,N_1746);
nor U11181 (N_11181,N_5049,N_5717);
or U11182 (N_11182,N_5381,N_1821);
or U11183 (N_11183,N_2424,N_694);
nand U11184 (N_11184,N_5303,N_1222);
and U11185 (N_11185,N_5716,N_2338);
and U11186 (N_11186,N_4508,N_3897);
or U11187 (N_11187,N_1250,N_5382);
nor U11188 (N_11188,N_4445,N_123);
nand U11189 (N_11189,N_5348,N_4532);
or U11190 (N_11190,N_4404,N_1308);
nor U11191 (N_11191,N_5001,N_1810);
nand U11192 (N_11192,N_1901,N_5467);
or U11193 (N_11193,N_1748,N_2652);
and U11194 (N_11194,N_4278,N_2248);
nand U11195 (N_11195,N_4403,N_5364);
nor U11196 (N_11196,N_2540,N_3066);
nor U11197 (N_11197,N_2733,N_4117);
nand U11198 (N_11198,N_1263,N_5138);
or U11199 (N_11199,N_260,N_2632);
nor U11200 (N_11200,N_3842,N_3538);
nand U11201 (N_11201,N_1363,N_3558);
nand U11202 (N_11202,N_4861,N_5419);
nor U11203 (N_11203,N_150,N_970);
or U11204 (N_11204,N_639,N_2575);
xor U11205 (N_11205,N_5228,N_5044);
nor U11206 (N_11206,N_4035,N_675);
or U11207 (N_11207,N_4114,N_1082);
and U11208 (N_11208,N_2683,N_3626);
or U11209 (N_11209,N_5213,N_4111);
and U11210 (N_11210,N_5618,N_4696);
and U11211 (N_11211,N_1405,N_213);
or U11212 (N_11212,N_4630,N_193);
nand U11213 (N_11213,N_3795,N_2253);
and U11214 (N_11214,N_3879,N_5047);
nor U11215 (N_11215,N_3225,N_2517);
nor U11216 (N_11216,N_631,N_1196);
nand U11217 (N_11217,N_4140,N_2602);
nand U11218 (N_11218,N_746,N_3791);
or U11219 (N_11219,N_5099,N_2040);
and U11220 (N_11220,N_1839,N_4629);
and U11221 (N_11221,N_4061,N_726);
nand U11222 (N_11222,N_3523,N_4098);
or U11223 (N_11223,N_4763,N_678);
and U11224 (N_11224,N_2966,N_4559);
and U11225 (N_11225,N_3715,N_5843);
nor U11226 (N_11226,N_2469,N_2066);
xnor U11227 (N_11227,N_3922,N_426);
nor U11228 (N_11228,N_1244,N_5140);
and U11229 (N_11229,N_1078,N_2201);
nor U11230 (N_11230,N_3161,N_891);
and U11231 (N_11231,N_4936,N_5577);
or U11232 (N_11232,N_1104,N_2730);
and U11233 (N_11233,N_2727,N_1625);
nand U11234 (N_11234,N_3290,N_422);
or U11235 (N_11235,N_5719,N_3571);
nand U11236 (N_11236,N_5423,N_2081);
nor U11237 (N_11237,N_1293,N_2989);
nor U11238 (N_11238,N_2237,N_4204);
or U11239 (N_11239,N_1903,N_5930);
xor U11240 (N_11240,N_4812,N_233);
and U11241 (N_11241,N_5874,N_2957);
or U11242 (N_11242,N_3549,N_275);
nor U11243 (N_11243,N_3669,N_3191);
and U11244 (N_11244,N_5212,N_5874);
and U11245 (N_11245,N_2953,N_3878);
and U11246 (N_11246,N_2905,N_569);
and U11247 (N_11247,N_2817,N_5034);
and U11248 (N_11248,N_5881,N_3759);
or U11249 (N_11249,N_4901,N_1252);
xor U11250 (N_11250,N_2505,N_1547);
and U11251 (N_11251,N_1478,N_5035);
xor U11252 (N_11252,N_5178,N_4992);
nand U11253 (N_11253,N_4357,N_3330);
nor U11254 (N_11254,N_276,N_5287);
xnor U11255 (N_11255,N_5671,N_349);
and U11256 (N_11256,N_1425,N_5418);
or U11257 (N_11257,N_3025,N_4930);
and U11258 (N_11258,N_4298,N_3454);
nand U11259 (N_11259,N_4093,N_262);
xnor U11260 (N_11260,N_825,N_2845);
xor U11261 (N_11261,N_2893,N_2572);
and U11262 (N_11262,N_3229,N_4079);
or U11263 (N_11263,N_2300,N_2882);
and U11264 (N_11264,N_1966,N_1196);
nor U11265 (N_11265,N_447,N_1809);
nor U11266 (N_11266,N_314,N_4209);
and U11267 (N_11267,N_443,N_163);
nand U11268 (N_11268,N_51,N_2530);
xnor U11269 (N_11269,N_3476,N_5737);
nand U11270 (N_11270,N_5145,N_2068);
nor U11271 (N_11271,N_2647,N_3875);
nand U11272 (N_11272,N_5961,N_3495);
or U11273 (N_11273,N_1232,N_986);
and U11274 (N_11274,N_905,N_191);
nand U11275 (N_11275,N_248,N_1007);
xor U11276 (N_11276,N_3634,N_223);
and U11277 (N_11277,N_5688,N_3954);
and U11278 (N_11278,N_1935,N_999);
and U11279 (N_11279,N_2605,N_527);
nand U11280 (N_11280,N_3232,N_3148);
nand U11281 (N_11281,N_1500,N_589);
nor U11282 (N_11282,N_765,N_4087);
or U11283 (N_11283,N_2517,N_1696);
and U11284 (N_11284,N_4656,N_3810);
or U11285 (N_11285,N_4093,N_4918);
nand U11286 (N_11286,N_3793,N_350);
nand U11287 (N_11287,N_1161,N_3913);
or U11288 (N_11288,N_3695,N_501);
xnor U11289 (N_11289,N_3617,N_27);
nand U11290 (N_11290,N_1908,N_4583);
or U11291 (N_11291,N_2223,N_2507);
nand U11292 (N_11292,N_1276,N_4918);
nor U11293 (N_11293,N_2822,N_2716);
nor U11294 (N_11294,N_3117,N_4598);
and U11295 (N_11295,N_3815,N_10);
nand U11296 (N_11296,N_5895,N_4772);
xnor U11297 (N_11297,N_391,N_89);
nor U11298 (N_11298,N_3216,N_4216);
or U11299 (N_11299,N_2056,N_5534);
nand U11300 (N_11300,N_3441,N_1333);
nand U11301 (N_11301,N_1673,N_5150);
nor U11302 (N_11302,N_4025,N_1519);
and U11303 (N_11303,N_3301,N_3929);
or U11304 (N_11304,N_2972,N_5471);
nand U11305 (N_11305,N_5664,N_3530);
and U11306 (N_11306,N_730,N_1662);
or U11307 (N_11307,N_5367,N_1683);
or U11308 (N_11308,N_3263,N_3723);
and U11309 (N_11309,N_717,N_2701);
xor U11310 (N_11310,N_4281,N_3682);
and U11311 (N_11311,N_3397,N_1152);
nor U11312 (N_11312,N_2760,N_4185);
nand U11313 (N_11313,N_3508,N_3801);
nand U11314 (N_11314,N_1193,N_1332);
nor U11315 (N_11315,N_2800,N_4671);
nand U11316 (N_11316,N_3551,N_2159);
and U11317 (N_11317,N_2648,N_801);
nor U11318 (N_11318,N_2956,N_469);
nor U11319 (N_11319,N_763,N_2802);
and U11320 (N_11320,N_772,N_3714);
nor U11321 (N_11321,N_208,N_1190);
and U11322 (N_11322,N_2471,N_743);
and U11323 (N_11323,N_5626,N_4971);
nor U11324 (N_11324,N_3709,N_219);
xor U11325 (N_11325,N_3491,N_1888);
and U11326 (N_11326,N_4666,N_3342);
and U11327 (N_11327,N_5177,N_4478);
nand U11328 (N_11328,N_4468,N_4200);
nor U11329 (N_11329,N_501,N_1434);
nand U11330 (N_11330,N_4898,N_5753);
nor U11331 (N_11331,N_3734,N_1740);
nor U11332 (N_11332,N_547,N_5042);
nor U11333 (N_11333,N_5092,N_5910);
nand U11334 (N_11334,N_3484,N_5036);
or U11335 (N_11335,N_5778,N_2270);
nor U11336 (N_11336,N_2703,N_1759);
and U11337 (N_11337,N_396,N_4194);
nand U11338 (N_11338,N_102,N_1998);
nor U11339 (N_11339,N_3631,N_3166);
xor U11340 (N_11340,N_2633,N_4489);
or U11341 (N_11341,N_1925,N_247);
or U11342 (N_11342,N_3707,N_3019);
and U11343 (N_11343,N_799,N_5908);
nor U11344 (N_11344,N_3794,N_5777);
nor U11345 (N_11345,N_3245,N_3459);
xor U11346 (N_11346,N_3298,N_2981);
nor U11347 (N_11347,N_2442,N_882);
nor U11348 (N_11348,N_3749,N_3242);
xnor U11349 (N_11349,N_2183,N_4854);
and U11350 (N_11350,N_2688,N_1221);
nor U11351 (N_11351,N_2615,N_2359);
and U11352 (N_11352,N_1260,N_3084);
and U11353 (N_11353,N_4518,N_1547);
and U11354 (N_11354,N_4533,N_527);
or U11355 (N_11355,N_3352,N_5792);
and U11356 (N_11356,N_4217,N_5132);
and U11357 (N_11357,N_5745,N_570);
or U11358 (N_11358,N_4711,N_4791);
nor U11359 (N_11359,N_1744,N_4526);
nor U11360 (N_11360,N_4395,N_4686);
or U11361 (N_11361,N_2327,N_4947);
and U11362 (N_11362,N_786,N_3453);
and U11363 (N_11363,N_3966,N_5185);
nor U11364 (N_11364,N_3075,N_2425);
nor U11365 (N_11365,N_4910,N_5327);
nor U11366 (N_11366,N_3599,N_5409);
nand U11367 (N_11367,N_2429,N_2061);
and U11368 (N_11368,N_4806,N_3145);
or U11369 (N_11369,N_1494,N_915);
or U11370 (N_11370,N_2936,N_229);
and U11371 (N_11371,N_1585,N_410);
nor U11372 (N_11372,N_2966,N_341);
and U11373 (N_11373,N_5176,N_1009);
xor U11374 (N_11374,N_732,N_1757);
or U11375 (N_11375,N_1213,N_2656);
nor U11376 (N_11376,N_5612,N_1145);
and U11377 (N_11377,N_4660,N_4827);
nor U11378 (N_11378,N_1560,N_397);
nand U11379 (N_11379,N_3513,N_343);
xor U11380 (N_11380,N_4905,N_5982);
nand U11381 (N_11381,N_1765,N_5797);
nor U11382 (N_11382,N_2403,N_1842);
xor U11383 (N_11383,N_2704,N_2430);
or U11384 (N_11384,N_4996,N_3237);
nor U11385 (N_11385,N_859,N_3880);
and U11386 (N_11386,N_2798,N_4717);
nand U11387 (N_11387,N_3862,N_5920);
and U11388 (N_11388,N_4798,N_737);
and U11389 (N_11389,N_5460,N_4903);
xor U11390 (N_11390,N_3060,N_5771);
and U11391 (N_11391,N_5354,N_4038);
nand U11392 (N_11392,N_3978,N_1857);
and U11393 (N_11393,N_462,N_3345);
and U11394 (N_11394,N_3969,N_4442);
or U11395 (N_11395,N_3618,N_3151);
nor U11396 (N_11396,N_2160,N_1858);
nor U11397 (N_11397,N_4756,N_183);
nor U11398 (N_11398,N_2615,N_185);
and U11399 (N_11399,N_991,N_4341);
nor U11400 (N_11400,N_3387,N_2477);
nor U11401 (N_11401,N_4427,N_3576);
and U11402 (N_11402,N_5812,N_1);
or U11403 (N_11403,N_2963,N_612);
xor U11404 (N_11404,N_316,N_2428);
xor U11405 (N_11405,N_575,N_1950);
and U11406 (N_11406,N_3402,N_3701);
nand U11407 (N_11407,N_2135,N_116);
nor U11408 (N_11408,N_2779,N_170);
and U11409 (N_11409,N_4451,N_3328);
or U11410 (N_11410,N_4064,N_5460);
xnor U11411 (N_11411,N_4831,N_1967);
nand U11412 (N_11412,N_4797,N_4048);
nor U11413 (N_11413,N_3261,N_3089);
or U11414 (N_11414,N_4001,N_5772);
and U11415 (N_11415,N_2488,N_5164);
or U11416 (N_11416,N_1246,N_1557);
and U11417 (N_11417,N_5914,N_5037);
xnor U11418 (N_11418,N_4700,N_3332);
nand U11419 (N_11419,N_3525,N_5513);
xor U11420 (N_11420,N_4072,N_3118);
xnor U11421 (N_11421,N_4391,N_3262);
nand U11422 (N_11422,N_1255,N_4309);
nor U11423 (N_11423,N_679,N_261);
nand U11424 (N_11424,N_4084,N_4573);
and U11425 (N_11425,N_830,N_2585);
and U11426 (N_11426,N_2177,N_39);
and U11427 (N_11427,N_5122,N_451);
nand U11428 (N_11428,N_420,N_5749);
or U11429 (N_11429,N_3506,N_2412);
nand U11430 (N_11430,N_5574,N_306);
or U11431 (N_11431,N_5617,N_2928);
and U11432 (N_11432,N_3462,N_4820);
nand U11433 (N_11433,N_43,N_4715);
and U11434 (N_11434,N_575,N_271);
nand U11435 (N_11435,N_3963,N_4916);
nand U11436 (N_11436,N_4111,N_1845);
nor U11437 (N_11437,N_1897,N_5546);
nor U11438 (N_11438,N_1780,N_4705);
or U11439 (N_11439,N_4770,N_1964);
and U11440 (N_11440,N_3144,N_5381);
nand U11441 (N_11441,N_2768,N_4417);
nor U11442 (N_11442,N_1617,N_1835);
nand U11443 (N_11443,N_4024,N_3128);
or U11444 (N_11444,N_351,N_1564);
xor U11445 (N_11445,N_2005,N_4532);
or U11446 (N_11446,N_3211,N_1351);
nand U11447 (N_11447,N_2438,N_2819);
and U11448 (N_11448,N_4551,N_1915);
nor U11449 (N_11449,N_4270,N_3732);
nand U11450 (N_11450,N_2884,N_4784);
nor U11451 (N_11451,N_4527,N_2909);
xor U11452 (N_11452,N_2280,N_1954);
nor U11453 (N_11453,N_385,N_1685);
and U11454 (N_11454,N_5167,N_511);
nor U11455 (N_11455,N_3464,N_3621);
nor U11456 (N_11456,N_4271,N_5252);
nor U11457 (N_11457,N_4353,N_1138);
or U11458 (N_11458,N_2833,N_711);
nor U11459 (N_11459,N_1312,N_4078);
nor U11460 (N_11460,N_5197,N_2825);
nand U11461 (N_11461,N_5185,N_4965);
or U11462 (N_11462,N_5922,N_5602);
or U11463 (N_11463,N_1179,N_3418);
nand U11464 (N_11464,N_2078,N_5233);
or U11465 (N_11465,N_2269,N_4254);
and U11466 (N_11466,N_5187,N_3780);
or U11467 (N_11467,N_1141,N_283);
or U11468 (N_11468,N_139,N_2765);
or U11469 (N_11469,N_4458,N_3493);
nand U11470 (N_11470,N_1426,N_3206);
xor U11471 (N_11471,N_4988,N_3513);
xor U11472 (N_11472,N_29,N_2413);
nand U11473 (N_11473,N_2855,N_2220);
xor U11474 (N_11474,N_1624,N_1595);
or U11475 (N_11475,N_4825,N_2311);
nor U11476 (N_11476,N_3139,N_2343);
nand U11477 (N_11477,N_4134,N_682);
or U11478 (N_11478,N_5754,N_1653);
or U11479 (N_11479,N_3435,N_5175);
nand U11480 (N_11480,N_2784,N_4326);
or U11481 (N_11481,N_135,N_2407);
or U11482 (N_11482,N_3334,N_4265);
or U11483 (N_11483,N_1944,N_5688);
or U11484 (N_11484,N_1402,N_904);
nor U11485 (N_11485,N_3681,N_1521);
nand U11486 (N_11486,N_4749,N_5401);
or U11487 (N_11487,N_3258,N_3577);
and U11488 (N_11488,N_4688,N_3970);
and U11489 (N_11489,N_326,N_2235);
and U11490 (N_11490,N_803,N_1622);
and U11491 (N_11491,N_2183,N_4170);
or U11492 (N_11492,N_4157,N_1367);
nand U11493 (N_11493,N_1760,N_517);
or U11494 (N_11494,N_3307,N_3020);
and U11495 (N_11495,N_4282,N_1170);
or U11496 (N_11496,N_5593,N_4185);
xor U11497 (N_11497,N_440,N_1308);
nor U11498 (N_11498,N_5277,N_172);
and U11499 (N_11499,N_5748,N_3187);
nand U11500 (N_11500,N_2576,N_3225);
nor U11501 (N_11501,N_2861,N_4255);
or U11502 (N_11502,N_1643,N_632);
or U11503 (N_11503,N_1003,N_3908);
nand U11504 (N_11504,N_2847,N_4497);
or U11505 (N_11505,N_1914,N_54);
xnor U11506 (N_11506,N_5300,N_2457);
and U11507 (N_11507,N_2851,N_586);
and U11508 (N_11508,N_5791,N_2190);
and U11509 (N_11509,N_3841,N_4940);
nor U11510 (N_11510,N_2560,N_5882);
and U11511 (N_11511,N_3239,N_1069);
or U11512 (N_11512,N_1115,N_5149);
and U11513 (N_11513,N_3387,N_1512);
xnor U11514 (N_11514,N_319,N_2293);
xnor U11515 (N_11515,N_406,N_5401);
and U11516 (N_11516,N_1057,N_4173);
and U11517 (N_11517,N_470,N_4044);
xnor U11518 (N_11518,N_5192,N_5431);
or U11519 (N_11519,N_2652,N_3451);
or U11520 (N_11520,N_3589,N_3722);
xor U11521 (N_11521,N_884,N_1205);
nor U11522 (N_11522,N_280,N_755);
or U11523 (N_11523,N_5543,N_1116);
and U11524 (N_11524,N_2969,N_4402);
nand U11525 (N_11525,N_3939,N_4336);
xnor U11526 (N_11526,N_5143,N_3034);
or U11527 (N_11527,N_2998,N_4103);
and U11528 (N_11528,N_92,N_2447);
nand U11529 (N_11529,N_4729,N_2129);
and U11530 (N_11530,N_5179,N_3065);
and U11531 (N_11531,N_4414,N_2095);
and U11532 (N_11532,N_1864,N_5950);
nand U11533 (N_11533,N_5871,N_3703);
nor U11534 (N_11534,N_3504,N_2253);
and U11535 (N_11535,N_2855,N_5576);
or U11536 (N_11536,N_1497,N_3331);
nand U11537 (N_11537,N_5414,N_4435);
and U11538 (N_11538,N_5817,N_2610);
and U11539 (N_11539,N_977,N_914);
nand U11540 (N_11540,N_2999,N_390);
nand U11541 (N_11541,N_720,N_2600);
and U11542 (N_11542,N_4713,N_57);
and U11543 (N_11543,N_5920,N_4825);
and U11544 (N_11544,N_1289,N_738);
xnor U11545 (N_11545,N_1125,N_281);
nand U11546 (N_11546,N_5974,N_5077);
nor U11547 (N_11547,N_3239,N_1008);
nor U11548 (N_11548,N_2873,N_2662);
or U11549 (N_11549,N_3438,N_665);
xor U11550 (N_11550,N_4167,N_2040);
xnor U11551 (N_11551,N_4922,N_1086);
nor U11552 (N_11552,N_3011,N_5628);
nor U11553 (N_11553,N_2402,N_4728);
or U11554 (N_11554,N_4231,N_2920);
or U11555 (N_11555,N_3,N_4890);
nor U11556 (N_11556,N_3870,N_3837);
and U11557 (N_11557,N_5885,N_2367);
and U11558 (N_11558,N_3220,N_1561);
nor U11559 (N_11559,N_980,N_382);
and U11560 (N_11560,N_859,N_5319);
nor U11561 (N_11561,N_1149,N_3923);
nor U11562 (N_11562,N_5692,N_439);
and U11563 (N_11563,N_260,N_625);
or U11564 (N_11564,N_4647,N_3487);
nand U11565 (N_11565,N_2688,N_1676);
nor U11566 (N_11566,N_1453,N_574);
xor U11567 (N_11567,N_5277,N_2299);
nand U11568 (N_11568,N_1286,N_1368);
nand U11569 (N_11569,N_1517,N_536);
and U11570 (N_11570,N_5090,N_1970);
and U11571 (N_11571,N_331,N_3272);
xnor U11572 (N_11572,N_3229,N_5078);
nor U11573 (N_11573,N_2786,N_4947);
nor U11574 (N_11574,N_2606,N_2587);
xor U11575 (N_11575,N_4518,N_4358);
or U11576 (N_11576,N_405,N_2786);
nor U11577 (N_11577,N_5982,N_1869);
nor U11578 (N_11578,N_2279,N_143);
or U11579 (N_11579,N_1544,N_210);
and U11580 (N_11580,N_5544,N_4977);
and U11581 (N_11581,N_5035,N_3854);
nor U11582 (N_11582,N_1064,N_4190);
nor U11583 (N_11583,N_2815,N_5177);
nor U11584 (N_11584,N_1896,N_3975);
nor U11585 (N_11585,N_3736,N_4069);
or U11586 (N_11586,N_1935,N_926);
nor U11587 (N_11587,N_5857,N_595);
nor U11588 (N_11588,N_449,N_1664);
and U11589 (N_11589,N_4922,N_828);
xor U11590 (N_11590,N_1472,N_3163);
nor U11591 (N_11591,N_827,N_2592);
nor U11592 (N_11592,N_4357,N_4127);
and U11593 (N_11593,N_2943,N_1173);
nor U11594 (N_11594,N_4622,N_400);
and U11595 (N_11595,N_1069,N_3406);
and U11596 (N_11596,N_1801,N_879);
xnor U11597 (N_11597,N_1322,N_2720);
nand U11598 (N_11598,N_5581,N_4558);
and U11599 (N_11599,N_5862,N_2532);
xor U11600 (N_11600,N_4770,N_3807);
and U11601 (N_11601,N_2816,N_5938);
and U11602 (N_11602,N_2989,N_484);
xnor U11603 (N_11603,N_4629,N_3057);
and U11604 (N_11604,N_4918,N_1520);
and U11605 (N_11605,N_3909,N_1560);
xor U11606 (N_11606,N_262,N_1006);
or U11607 (N_11607,N_4156,N_5712);
and U11608 (N_11608,N_1063,N_1775);
xor U11609 (N_11609,N_721,N_4598);
nor U11610 (N_11610,N_5952,N_5111);
or U11611 (N_11611,N_202,N_4887);
nand U11612 (N_11612,N_5324,N_960);
nand U11613 (N_11613,N_1102,N_4071);
or U11614 (N_11614,N_896,N_1844);
nand U11615 (N_11615,N_5480,N_3707);
nand U11616 (N_11616,N_3529,N_1298);
or U11617 (N_11617,N_4572,N_2973);
nor U11618 (N_11618,N_2540,N_242);
or U11619 (N_11619,N_3758,N_3776);
or U11620 (N_11620,N_3390,N_4678);
nor U11621 (N_11621,N_3928,N_5295);
nor U11622 (N_11622,N_1635,N_5929);
nand U11623 (N_11623,N_1593,N_992);
nor U11624 (N_11624,N_63,N_1685);
and U11625 (N_11625,N_3548,N_5836);
and U11626 (N_11626,N_2366,N_2877);
nand U11627 (N_11627,N_1725,N_4206);
and U11628 (N_11628,N_19,N_3327);
xnor U11629 (N_11629,N_4487,N_4525);
or U11630 (N_11630,N_5523,N_1435);
nor U11631 (N_11631,N_1953,N_243);
nor U11632 (N_11632,N_374,N_5807);
nand U11633 (N_11633,N_842,N_614);
xnor U11634 (N_11634,N_856,N_4482);
or U11635 (N_11635,N_5719,N_2996);
or U11636 (N_11636,N_5014,N_1243);
nor U11637 (N_11637,N_778,N_1399);
and U11638 (N_11638,N_3924,N_3189);
nor U11639 (N_11639,N_5181,N_3177);
or U11640 (N_11640,N_3659,N_419);
nor U11641 (N_11641,N_2573,N_1034);
nand U11642 (N_11642,N_373,N_3949);
nor U11643 (N_11643,N_152,N_5094);
nand U11644 (N_11644,N_5652,N_3003);
or U11645 (N_11645,N_3333,N_5849);
nand U11646 (N_11646,N_3843,N_5066);
nor U11647 (N_11647,N_2629,N_1084);
or U11648 (N_11648,N_2902,N_1673);
nand U11649 (N_11649,N_3580,N_1147);
nor U11650 (N_11650,N_334,N_516);
and U11651 (N_11651,N_3699,N_276);
nand U11652 (N_11652,N_159,N_1118);
or U11653 (N_11653,N_3514,N_2309);
nand U11654 (N_11654,N_5434,N_4973);
or U11655 (N_11655,N_2337,N_2487);
nor U11656 (N_11656,N_516,N_5626);
and U11657 (N_11657,N_1706,N_3225);
nand U11658 (N_11658,N_2687,N_874);
nand U11659 (N_11659,N_4807,N_2788);
xor U11660 (N_11660,N_5414,N_26);
nor U11661 (N_11661,N_2130,N_5797);
or U11662 (N_11662,N_1499,N_259);
xnor U11663 (N_11663,N_1682,N_4606);
and U11664 (N_11664,N_1005,N_190);
or U11665 (N_11665,N_4695,N_5986);
and U11666 (N_11666,N_2486,N_1459);
and U11667 (N_11667,N_802,N_5410);
nand U11668 (N_11668,N_4674,N_910);
or U11669 (N_11669,N_175,N_797);
or U11670 (N_11670,N_1883,N_777);
nor U11671 (N_11671,N_2208,N_4178);
or U11672 (N_11672,N_685,N_1898);
or U11673 (N_11673,N_2190,N_3008);
nand U11674 (N_11674,N_3512,N_1766);
nand U11675 (N_11675,N_251,N_4378);
xnor U11676 (N_11676,N_3060,N_1383);
nand U11677 (N_11677,N_2186,N_5931);
and U11678 (N_11678,N_3524,N_5199);
nor U11679 (N_11679,N_1702,N_5699);
xnor U11680 (N_11680,N_4018,N_3530);
nor U11681 (N_11681,N_2492,N_5970);
nand U11682 (N_11682,N_3084,N_1863);
or U11683 (N_11683,N_118,N_2589);
nor U11684 (N_11684,N_5472,N_1702);
or U11685 (N_11685,N_290,N_444);
or U11686 (N_11686,N_5019,N_2307);
and U11687 (N_11687,N_4716,N_3340);
nand U11688 (N_11688,N_221,N_156);
or U11689 (N_11689,N_591,N_3167);
xor U11690 (N_11690,N_762,N_4339);
xor U11691 (N_11691,N_1170,N_5752);
nand U11692 (N_11692,N_3708,N_4012);
and U11693 (N_11693,N_2635,N_5311);
nand U11694 (N_11694,N_1498,N_27);
or U11695 (N_11695,N_5489,N_3508);
or U11696 (N_11696,N_1723,N_2456);
nor U11697 (N_11697,N_1190,N_5088);
and U11698 (N_11698,N_4216,N_5984);
and U11699 (N_11699,N_2402,N_3741);
and U11700 (N_11700,N_3726,N_4745);
xor U11701 (N_11701,N_2241,N_2224);
nand U11702 (N_11702,N_3607,N_581);
and U11703 (N_11703,N_3605,N_3293);
nand U11704 (N_11704,N_1534,N_325);
nor U11705 (N_11705,N_1143,N_5534);
nand U11706 (N_11706,N_4041,N_2172);
xnor U11707 (N_11707,N_5496,N_1891);
xor U11708 (N_11708,N_2316,N_3631);
or U11709 (N_11709,N_3878,N_1441);
or U11710 (N_11710,N_1411,N_5521);
nand U11711 (N_11711,N_2881,N_3852);
or U11712 (N_11712,N_3271,N_3989);
nor U11713 (N_11713,N_357,N_4981);
and U11714 (N_11714,N_2030,N_4332);
nand U11715 (N_11715,N_577,N_19);
and U11716 (N_11716,N_5674,N_3362);
nor U11717 (N_11717,N_5056,N_973);
nor U11718 (N_11718,N_1164,N_4176);
nand U11719 (N_11719,N_4441,N_4409);
xor U11720 (N_11720,N_1451,N_5521);
nor U11721 (N_11721,N_910,N_4196);
or U11722 (N_11722,N_1134,N_2995);
nand U11723 (N_11723,N_4802,N_147);
or U11724 (N_11724,N_2528,N_580);
or U11725 (N_11725,N_818,N_2526);
nand U11726 (N_11726,N_5494,N_2099);
or U11727 (N_11727,N_832,N_1291);
nand U11728 (N_11728,N_5601,N_4386);
nor U11729 (N_11729,N_76,N_1746);
nand U11730 (N_11730,N_2978,N_4746);
nand U11731 (N_11731,N_2446,N_1632);
and U11732 (N_11732,N_803,N_966);
xnor U11733 (N_11733,N_1390,N_3772);
or U11734 (N_11734,N_1756,N_1980);
nor U11735 (N_11735,N_3109,N_3190);
nor U11736 (N_11736,N_5600,N_2814);
and U11737 (N_11737,N_4610,N_922);
or U11738 (N_11738,N_4682,N_4870);
nand U11739 (N_11739,N_3787,N_3538);
or U11740 (N_11740,N_504,N_2361);
nor U11741 (N_11741,N_1672,N_4931);
or U11742 (N_11742,N_1763,N_601);
or U11743 (N_11743,N_3170,N_3949);
xor U11744 (N_11744,N_2005,N_4675);
nand U11745 (N_11745,N_1968,N_5111);
and U11746 (N_11746,N_1737,N_3292);
nor U11747 (N_11747,N_2572,N_1356);
and U11748 (N_11748,N_3520,N_2193);
nand U11749 (N_11749,N_4439,N_2540);
nand U11750 (N_11750,N_4394,N_455);
nand U11751 (N_11751,N_3839,N_100);
nand U11752 (N_11752,N_5469,N_4049);
nand U11753 (N_11753,N_5973,N_1721);
and U11754 (N_11754,N_1455,N_5769);
or U11755 (N_11755,N_966,N_4791);
nand U11756 (N_11756,N_281,N_4597);
nand U11757 (N_11757,N_3171,N_3599);
nor U11758 (N_11758,N_2703,N_4285);
nand U11759 (N_11759,N_3376,N_4911);
or U11760 (N_11760,N_752,N_4355);
nor U11761 (N_11761,N_3694,N_1046);
and U11762 (N_11762,N_1703,N_381);
or U11763 (N_11763,N_2125,N_1961);
or U11764 (N_11764,N_5034,N_49);
nand U11765 (N_11765,N_5617,N_1603);
nor U11766 (N_11766,N_3315,N_1388);
nand U11767 (N_11767,N_2304,N_594);
nor U11768 (N_11768,N_1352,N_1488);
and U11769 (N_11769,N_4806,N_2711);
or U11770 (N_11770,N_908,N_4286);
nand U11771 (N_11771,N_3006,N_1490);
and U11772 (N_11772,N_5388,N_2818);
nor U11773 (N_11773,N_4990,N_1552);
or U11774 (N_11774,N_3414,N_661);
nor U11775 (N_11775,N_2349,N_572);
nor U11776 (N_11776,N_3567,N_1037);
and U11777 (N_11777,N_5892,N_4759);
or U11778 (N_11778,N_4706,N_2387);
nand U11779 (N_11779,N_636,N_2132);
or U11780 (N_11780,N_1298,N_1036);
and U11781 (N_11781,N_4675,N_1152);
or U11782 (N_11782,N_5756,N_5182);
nand U11783 (N_11783,N_3670,N_1907);
nand U11784 (N_11784,N_4637,N_3558);
nor U11785 (N_11785,N_2577,N_4753);
nor U11786 (N_11786,N_3145,N_3971);
and U11787 (N_11787,N_3123,N_3282);
nor U11788 (N_11788,N_132,N_1078);
nand U11789 (N_11789,N_3521,N_2734);
nor U11790 (N_11790,N_763,N_2620);
or U11791 (N_11791,N_3044,N_199);
or U11792 (N_11792,N_575,N_4079);
and U11793 (N_11793,N_838,N_3731);
nand U11794 (N_11794,N_3883,N_3071);
and U11795 (N_11795,N_2863,N_4571);
nor U11796 (N_11796,N_1653,N_3847);
and U11797 (N_11797,N_2021,N_2272);
and U11798 (N_11798,N_4277,N_922);
or U11799 (N_11799,N_2293,N_670);
xor U11800 (N_11800,N_3035,N_2034);
or U11801 (N_11801,N_1604,N_825);
nor U11802 (N_11802,N_2264,N_4385);
nand U11803 (N_11803,N_3203,N_134);
nor U11804 (N_11804,N_236,N_3267);
or U11805 (N_11805,N_3545,N_1277);
nor U11806 (N_11806,N_5359,N_3920);
or U11807 (N_11807,N_2760,N_1186);
nor U11808 (N_11808,N_1708,N_274);
nor U11809 (N_11809,N_803,N_908);
nor U11810 (N_11810,N_3550,N_5753);
or U11811 (N_11811,N_1395,N_110);
and U11812 (N_11812,N_5981,N_893);
and U11813 (N_11813,N_3806,N_2054);
nor U11814 (N_11814,N_455,N_2234);
and U11815 (N_11815,N_1862,N_1358);
nand U11816 (N_11816,N_2781,N_4833);
or U11817 (N_11817,N_3640,N_3053);
or U11818 (N_11818,N_2529,N_90);
and U11819 (N_11819,N_5976,N_4855);
nand U11820 (N_11820,N_1334,N_1406);
nor U11821 (N_11821,N_4711,N_4280);
or U11822 (N_11822,N_3894,N_347);
and U11823 (N_11823,N_4809,N_562);
and U11824 (N_11824,N_274,N_5358);
nand U11825 (N_11825,N_3848,N_3835);
nor U11826 (N_11826,N_4593,N_529);
and U11827 (N_11827,N_5162,N_2423);
or U11828 (N_11828,N_67,N_1200);
nand U11829 (N_11829,N_2675,N_4589);
and U11830 (N_11830,N_1982,N_3277);
and U11831 (N_11831,N_2071,N_681);
and U11832 (N_11832,N_3869,N_4882);
nand U11833 (N_11833,N_2141,N_3092);
and U11834 (N_11834,N_1843,N_673);
or U11835 (N_11835,N_5913,N_3783);
nor U11836 (N_11836,N_1329,N_4946);
nor U11837 (N_11837,N_5938,N_2812);
nor U11838 (N_11838,N_2573,N_5511);
xnor U11839 (N_11839,N_2503,N_1238);
nand U11840 (N_11840,N_893,N_4077);
or U11841 (N_11841,N_3822,N_3546);
nor U11842 (N_11842,N_3128,N_4615);
nor U11843 (N_11843,N_2691,N_4461);
and U11844 (N_11844,N_5943,N_1503);
xnor U11845 (N_11845,N_3384,N_319);
and U11846 (N_11846,N_5836,N_5121);
or U11847 (N_11847,N_1916,N_2264);
xnor U11848 (N_11848,N_4292,N_4170);
nand U11849 (N_11849,N_359,N_467);
nand U11850 (N_11850,N_3550,N_1905);
nand U11851 (N_11851,N_272,N_2839);
nor U11852 (N_11852,N_2318,N_5156);
nor U11853 (N_11853,N_298,N_1304);
nand U11854 (N_11854,N_3483,N_2405);
nand U11855 (N_11855,N_1094,N_5380);
nand U11856 (N_11856,N_311,N_4649);
nor U11857 (N_11857,N_4270,N_2083);
nand U11858 (N_11858,N_682,N_3960);
or U11859 (N_11859,N_3901,N_4029);
xor U11860 (N_11860,N_2360,N_1160);
and U11861 (N_11861,N_4061,N_2631);
or U11862 (N_11862,N_614,N_4023);
and U11863 (N_11863,N_4800,N_2854);
or U11864 (N_11864,N_719,N_3343);
and U11865 (N_11865,N_1914,N_5928);
and U11866 (N_11866,N_5609,N_496);
nor U11867 (N_11867,N_1756,N_5676);
or U11868 (N_11868,N_5402,N_3248);
nand U11869 (N_11869,N_4370,N_1433);
xnor U11870 (N_11870,N_3074,N_4976);
nor U11871 (N_11871,N_451,N_359);
xor U11872 (N_11872,N_4564,N_4882);
xnor U11873 (N_11873,N_3140,N_3862);
nand U11874 (N_11874,N_1893,N_3270);
or U11875 (N_11875,N_589,N_5771);
nor U11876 (N_11876,N_4107,N_2947);
and U11877 (N_11877,N_5084,N_418);
xor U11878 (N_11878,N_1573,N_1559);
nor U11879 (N_11879,N_2354,N_529);
or U11880 (N_11880,N_3004,N_960);
or U11881 (N_11881,N_4799,N_3751);
nand U11882 (N_11882,N_5818,N_4523);
nand U11883 (N_11883,N_2375,N_4635);
nand U11884 (N_11884,N_3206,N_5066);
nand U11885 (N_11885,N_3652,N_3137);
and U11886 (N_11886,N_154,N_1866);
or U11887 (N_11887,N_213,N_2254);
nor U11888 (N_11888,N_1253,N_184);
nand U11889 (N_11889,N_2435,N_1119);
or U11890 (N_11890,N_581,N_3509);
nor U11891 (N_11891,N_4235,N_1012);
or U11892 (N_11892,N_1694,N_265);
and U11893 (N_11893,N_3140,N_4159);
nor U11894 (N_11894,N_4319,N_4402);
or U11895 (N_11895,N_2570,N_5833);
and U11896 (N_11896,N_1516,N_85);
nand U11897 (N_11897,N_144,N_1319);
nor U11898 (N_11898,N_1586,N_3860);
nor U11899 (N_11899,N_386,N_3788);
nand U11900 (N_11900,N_4937,N_1269);
or U11901 (N_11901,N_3997,N_3217);
nor U11902 (N_11902,N_795,N_5283);
nand U11903 (N_11903,N_679,N_1134);
or U11904 (N_11904,N_1632,N_1885);
and U11905 (N_11905,N_477,N_2009);
xnor U11906 (N_11906,N_1987,N_999);
xnor U11907 (N_11907,N_1763,N_3330);
or U11908 (N_11908,N_111,N_4635);
nor U11909 (N_11909,N_5680,N_5602);
or U11910 (N_11910,N_4960,N_5018);
or U11911 (N_11911,N_2722,N_5704);
or U11912 (N_11912,N_4082,N_5445);
and U11913 (N_11913,N_5139,N_3506);
and U11914 (N_11914,N_1990,N_874);
nand U11915 (N_11915,N_2195,N_1411);
nand U11916 (N_11916,N_448,N_2226);
nand U11917 (N_11917,N_2165,N_2004);
nand U11918 (N_11918,N_3881,N_5805);
and U11919 (N_11919,N_5983,N_736);
nand U11920 (N_11920,N_5548,N_1893);
or U11921 (N_11921,N_3147,N_2042);
xor U11922 (N_11922,N_5311,N_5789);
nor U11923 (N_11923,N_1585,N_3978);
and U11924 (N_11924,N_5231,N_3124);
nor U11925 (N_11925,N_1446,N_3609);
nand U11926 (N_11926,N_4964,N_677);
nor U11927 (N_11927,N_3183,N_2219);
nor U11928 (N_11928,N_5330,N_2748);
or U11929 (N_11929,N_1451,N_941);
or U11930 (N_11930,N_820,N_156);
or U11931 (N_11931,N_4683,N_2383);
or U11932 (N_11932,N_2806,N_5827);
xnor U11933 (N_11933,N_3236,N_1713);
and U11934 (N_11934,N_4543,N_4793);
xor U11935 (N_11935,N_5847,N_894);
nand U11936 (N_11936,N_4426,N_5937);
or U11937 (N_11937,N_5794,N_2046);
and U11938 (N_11938,N_3653,N_1717);
or U11939 (N_11939,N_5026,N_738);
and U11940 (N_11940,N_3967,N_3708);
nand U11941 (N_11941,N_4018,N_362);
xor U11942 (N_11942,N_3295,N_2417);
nor U11943 (N_11943,N_1302,N_4395);
nand U11944 (N_11944,N_4319,N_4142);
or U11945 (N_11945,N_1753,N_5161);
nand U11946 (N_11946,N_5785,N_278);
nor U11947 (N_11947,N_4751,N_4191);
xor U11948 (N_11948,N_285,N_3304);
or U11949 (N_11949,N_3236,N_5413);
or U11950 (N_11950,N_3708,N_3273);
and U11951 (N_11951,N_2906,N_854);
nor U11952 (N_11952,N_3215,N_3136);
or U11953 (N_11953,N_4535,N_3795);
nand U11954 (N_11954,N_615,N_4179);
nor U11955 (N_11955,N_602,N_1931);
or U11956 (N_11956,N_420,N_1386);
or U11957 (N_11957,N_1719,N_2217);
and U11958 (N_11958,N_557,N_4985);
or U11959 (N_11959,N_2401,N_518);
and U11960 (N_11960,N_2636,N_4553);
or U11961 (N_11961,N_4742,N_368);
nand U11962 (N_11962,N_662,N_2193);
or U11963 (N_11963,N_2089,N_1462);
or U11964 (N_11964,N_1773,N_812);
and U11965 (N_11965,N_1803,N_3928);
nand U11966 (N_11966,N_3256,N_459);
nand U11967 (N_11967,N_2827,N_4196);
nand U11968 (N_11968,N_5124,N_4187);
nor U11969 (N_11969,N_3421,N_707);
and U11970 (N_11970,N_3272,N_1299);
nor U11971 (N_11971,N_3268,N_190);
nand U11972 (N_11972,N_3983,N_3537);
or U11973 (N_11973,N_419,N_3963);
xnor U11974 (N_11974,N_870,N_4761);
or U11975 (N_11975,N_2986,N_105);
nand U11976 (N_11976,N_5458,N_998);
or U11977 (N_11977,N_5129,N_3308);
nand U11978 (N_11978,N_838,N_5157);
nand U11979 (N_11979,N_151,N_5367);
and U11980 (N_11980,N_2183,N_1671);
and U11981 (N_11981,N_1376,N_1354);
xnor U11982 (N_11982,N_3456,N_581);
nor U11983 (N_11983,N_2945,N_1216);
nand U11984 (N_11984,N_893,N_3439);
nand U11985 (N_11985,N_3926,N_3100);
or U11986 (N_11986,N_5464,N_812);
nor U11987 (N_11987,N_1093,N_5872);
xor U11988 (N_11988,N_1289,N_5694);
or U11989 (N_11989,N_5572,N_5607);
xnor U11990 (N_11990,N_5281,N_1864);
and U11991 (N_11991,N_1839,N_1938);
and U11992 (N_11992,N_4541,N_4538);
nor U11993 (N_11993,N_4019,N_3409);
or U11994 (N_11994,N_1378,N_5254);
nor U11995 (N_11995,N_4480,N_2068);
nor U11996 (N_11996,N_4145,N_4888);
and U11997 (N_11997,N_2140,N_3375);
nand U11998 (N_11998,N_521,N_3525);
xnor U11999 (N_11999,N_5590,N_592);
and U12000 (N_12000,N_9960,N_8599);
or U12001 (N_12001,N_9642,N_7085);
nand U12002 (N_12002,N_11354,N_7775);
nand U12003 (N_12003,N_9234,N_6796);
or U12004 (N_12004,N_8037,N_8107);
nor U12005 (N_12005,N_10252,N_8790);
nor U12006 (N_12006,N_7639,N_9916);
nand U12007 (N_12007,N_9955,N_9679);
and U12008 (N_12008,N_9295,N_11849);
and U12009 (N_12009,N_7511,N_10314);
or U12010 (N_12010,N_6354,N_9170);
and U12011 (N_12011,N_6438,N_9756);
and U12012 (N_12012,N_8303,N_8015);
xor U12013 (N_12013,N_7424,N_9020);
nand U12014 (N_12014,N_6131,N_9761);
nand U12015 (N_12015,N_8627,N_6530);
and U12016 (N_12016,N_11966,N_10051);
and U12017 (N_12017,N_6124,N_10349);
xnor U12018 (N_12018,N_10339,N_11525);
nand U12019 (N_12019,N_8464,N_11045);
nand U12020 (N_12020,N_8201,N_9653);
and U12021 (N_12021,N_6254,N_11147);
or U12022 (N_12022,N_11352,N_9276);
or U12023 (N_12023,N_10574,N_8002);
or U12024 (N_12024,N_11017,N_9751);
nand U12025 (N_12025,N_9786,N_7322);
or U12026 (N_12026,N_9497,N_11401);
and U12027 (N_12027,N_6920,N_10847);
and U12028 (N_12028,N_9816,N_9131);
nand U12029 (N_12029,N_7498,N_6763);
or U12030 (N_12030,N_7366,N_9190);
and U12031 (N_12031,N_10520,N_9980);
and U12032 (N_12032,N_11714,N_6099);
nand U12033 (N_12033,N_10709,N_11530);
nor U12034 (N_12034,N_7815,N_11566);
or U12035 (N_12035,N_10137,N_11360);
and U12036 (N_12036,N_6404,N_7169);
and U12037 (N_12037,N_7710,N_10729);
and U12038 (N_12038,N_8487,N_7555);
nor U12039 (N_12039,N_6273,N_7411);
and U12040 (N_12040,N_10103,N_11593);
nor U12041 (N_12041,N_8906,N_9403);
and U12042 (N_12042,N_10863,N_8331);
nor U12043 (N_12043,N_11144,N_11901);
nor U12044 (N_12044,N_10704,N_9535);
and U12045 (N_12045,N_6093,N_10287);
and U12046 (N_12046,N_9250,N_7230);
nor U12047 (N_12047,N_6483,N_11929);
xor U12048 (N_12048,N_9901,N_11029);
or U12049 (N_12049,N_11833,N_11513);
nand U12050 (N_12050,N_6921,N_11664);
xnor U12051 (N_12051,N_11280,N_7091);
or U12052 (N_12052,N_8795,N_9730);
nand U12053 (N_12053,N_6660,N_8441);
and U12054 (N_12054,N_7321,N_10482);
and U12055 (N_12055,N_8754,N_9668);
or U12056 (N_12056,N_11041,N_11063);
and U12057 (N_12057,N_7421,N_6814);
and U12058 (N_12058,N_7063,N_6659);
nor U12059 (N_12059,N_11660,N_7542);
and U12060 (N_12060,N_7677,N_8955);
and U12061 (N_12061,N_11392,N_7792);
and U12062 (N_12062,N_11866,N_7037);
and U12063 (N_12063,N_9870,N_10318);
and U12064 (N_12064,N_8761,N_9981);
or U12065 (N_12065,N_9006,N_6106);
or U12066 (N_12066,N_7353,N_7223);
xnor U12067 (N_12067,N_11223,N_6532);
nor U12068 (N_12068,N_7299,N_7712);
xnor U12069 (N_12069,N_9224,N_8071);
and U12070 (N_12070,N_6806,N_7401);
and U12071 (N_12071,N_8001,N_8456);
or U12072 (N_12072,N_9000,N_6815);
nand U12073 (N_12073,N_10901,N_6042);
or U12074 (N_12074,N_6421,N_11423);
nor U12075 (N_12075,N_7567,N_7144);
or U12076 (N_12076,N_11996,N_6703);
and U12077 (N_12077,N_11702,N_9284);
or U12078 (N_12078,N_11391,N_8908);
and U12079 (N_12079,N_7837,N_6210);
or U12080 (N_12080,N_6149,N_10861);
nand U12081 (N_12081,N_9483,N_7617);
and U12082 (N_12082,N_9289,N_7048);
nor U12083 (N_12083,N_8324,N_11773);
and U12084 (N_12084,N_10585,N_7630);
nand U12085 (N_12085,N_9147,N_8188);
and U12086 (N_12086,N_10175,N_8727);
and U12087 (N_12087,N_6973,N_6767);
and U12088 (N_12088,N_11947,N_8031);
nand U12089 (N_12089,N_9887,N_9713);
and U12090 (N_12090,N_7485,N_8405);
xnor U12091 (N_12091,N_9369,N_7900);
and U12092 (N_12092,N_10473,N_7975);
or U12093 (N_12093,N_11575,N_9512);
nor U12094 (N_12094,N_8447,N_11292);
nor U12095 (N_12095,N_11980,N_11272);
xnor U12096 (N_12096,N_8744,N_10122);
or U12097 (N_12097,N_11655,N_6558);
and U12098 (N_12098,N_6613,N_10794);
and U12099 (N_12099,N_7866,N_10059);
nand U12100 (N_12100,N_11690,N_9515);
nor U12101 (N_12101,N_9908,N_7013);
nand U12102 (N_12102,N_8218,N_6616);
nor U12103 (N_12103,N_10916,N_7875);
nand U12104 (N_12104,N_7281,N_7404);
xor U12105 (N_12105,N_9367,N_10423);
or U12106 (N_12106,N_10744,N_7842);
or U12107 (N_12107,N_9342,N_9691);
nand U12108 (N_12108,N_7006,N_9385);
nand U12109 (N_12109,N_11783,N_11739);
nand U12110 (N_12110,N_8788,N_11160);
xor U12111 (N_12111,N_10397,N_8609);
nand U12112 (N_12112,N_6259,N_6932);
nor U12113 (N_12113,N_9149,N_7676);
and U12114 (N_12114,N_7064,N_9759);
and U12115 (N_12115,N_7357,N_9805);
xnor U12116 (N_12116,N_11812,N_10911);
and U12117 (N_12117,N_10883,N_7448);
nor U12118 (N_12118,N_6875,N_9663);
and U12119 (N_12119,N_9658,N_7101);
or U12120 (N_12120,N_7583,N_9036);
nor U12121 (N_12121,N_6381,N_10081);
nor U12122 (N_12122,N_7440,N_10269);
or U12123 (N_12123,N_10271,N_8119);
nand U12124 (N_12124,N_7836,N_8753);
or U12125 (N_12125,N_6343,N_8704);
and U12126 (N_12126,N_11199,N_11761);
and U12127 (N_12127,N_10973,N_6489);
and U12128 (N_12128,N_11616,N_9776);
nor U12129 (N_12129,N_7827,N_7702);
nand U12130 (N_12130,N_11441,N_11168);
xnor U12131 (N_12131,N_9278,N_6067);
or U12132 (N_12132,N_6746,N_7500);
nor U12133 (N_12133,N_8115,N_9308);
and U12134 (N_12134,N_11411,N_6091);
or U12135 (N_12135,N_8596,N_11486);
or U12136 (N_12136,N_11084,N_8020);
and U12137 (N_12137,N_7286,N_10830);
nor U12138 (N_12138,N_8103,N_7878);
nor U12139 (N_12139,N_8675,N_7704);
and U12140 (N_12140,N_7205,N_9034);
or U12141 (N_12141,N_11804,N_9081);
nand U12142 (N_12142,N_9139,N_11046);
nand U12143 (N_12143,N_8543,N_10143);
nor U12144 (N_12144,N_11605,N_6205);
or U12145 (N_12145,N_7774,N_7474);
nor U12146 (N_12146,N_11619,N_9256);
xor U12147 (N_12147,N_11192,N_10112);
and U12148 (N_12148,N_11920,N_8863);
nor U12149 (N_12149,N_10549,N_11025);
and U12150 (N_12150,N_6615,N_6293);
nor U12151 (N_12151,N_10601,N_9069);
or U12152 (N_12152,N_11452,N_6694);
and U12153 (N_12153,N_10825,N_10995);
nor U12154 (N_12154,N_6678,N_9393);
nand U12155 (N_12155,N_11772,N_8547);
nand U12156 (N_12156,N_7125,N_11844);
nand U12157 (N_12157,N_11847,N_10722);
or U12158 (N_12158,N_9454,N_9014);
nand U12159 (N_12159,N_6445,N_8958);
nor U12160 (N_12160,N_7345,N_6211);
and U12161 (N_12161,N_8228,N_9845);
or U12162 (N_12162,N_11766,N_6538);
and U12163 (N_12163,N_11227,N_8875);
and U12164 (N_12164,N_11018,N_7591);
nand U12165 (N_12165,N_7059,N_10649);
xnor U12166 (N_12166,N_11538,N_6886);
nand U12167 (N_12167,N_8601,N_9425);
or U12168 (N_12168,N_7652,N_10238);
and U12169 (N_12169,N_11990,N_10413);
and U12170 (N_12170,N_9353,N_8118);
nand U12171 (N_12171,N_11485,N_7272);
xnor U12172 (N_12172,N_8409,N_6287);
and U12173 (N_12173,N_6598,N_11534);
nand U12174 (N_12174,N_7973,N_6656);
nand U12175 (N_12175,N_10904,N_7252);
nand U12176 (N_12176,N_7807,N_7834);
nor U12177 (N_12177,N_10121,N_6400);
nor U12178 (N_12178,N_9074,N_9809);
xor U12179 (N_12179,N_11681,N_8552);
or U12180 (N_12180,N_8408,N_11914);
nand U12181 (N_12181,N_8012,N_7147);
and U12182 (N_12182,N_8127,N_6079);
xnor U12183 (N_12183,N_9106,N_10371);
xor U12184 (N_12184,N_7671,N_8996);
nor U12185 (N_12185,N_10530,N_7342);
nand U12186 (N_12186,N_8975,N_8885);
and U12187 (N_12187,N_7516,N_8028);
nor U12188 (N_12188,N_7275,N_10948);
nor U12189 (N_12189,N_7871,N_10719);
xor U12190 (N_12190,N_9279,N_8310);
or U12191 (N_12191,N_11027,N_10996);
nand U12192 (N_12192,N_10002,N_6681);
or U12193 (N_12193,N_11611,N_7340);
xor U12194 (N_12194,N_8339,N_11562);
nand U12195 (N_12195,N_10650,N_8439);
and U12196 (N_12196,N_6959,N_11145);
nor U12197 (N_12197,N_11148,N_6208);
xnor U12198 (N_12198,N_9842,N_10934);
nor U12199 (N_12199,N_6983,N_11576);
xor U12200 (N_12200,N_7244,N_6851);
or U12201 (N_12201,N_6035,N_9184);
or U12202 (N_12202,N_10929,N_10640);
nor U12203 (N_12203,N_6166,N_11950);
nor U12204 (N_12204,N_9208,N_10355);
nor U12205 (N_12205,N_9134,N_6340);
nor U12206 (N_12206,N_8760,N_10485);
nand U12207 (N_12207,N_6611,N_10635);
nor U12208 (N_12208,N_7818,N_7817);
nand U12209 (N_12209,N_8555,N_9720);
and U12210 (N_12210,N_6213,N_11417);
nand U12211 (N_12211,N_9003,N_11234);
and U12212 (N_12212,N_11461,N_9118);
or U12213 (N_12213,N_8592,N_7713);
nor U12214 (N_12214,N_9101,N_8360);
nor U12215 (N_12215,N_9892,N_6178);
nor U12216 (N_12216,N_9741,N_9926);
and U12217 (N_12217,N_7435,N_9793);
nand U12218 (N_12218,N_9533,N_11474);
and U12219 (N_12219,N_7530,N_9522);
or U12220 (N_12220,N_9201,N_11735);
nor U12221 (N_12221,N_8433,N_9338);
or U12222 (N_12222,N_10582,N_11971);
xnor U12223 (N_12223,N_11725,N_7943);
and U12224 (N_12224,N_10716,N_10270);
xnor U12225 (N_12225,N_11995,N_7185);
nor U12226 (N_12226,N_11240,N_9007);
or U12227 (N_12227,N_10316,N_11344);
nand U12228 (N_12228,N_7663,N_7451);
nand U12229 (N_12229,N_9656,N_6915);
nor U12230 (N_12230,N_9912,N_11171);
nor U12231 (N_12231,N_11355,N_9817);
or U12232 (N_12232,N_6479,N_8137);
nor U12233 (N_12233,N_6800,N_6101);
and U12234 (N_12234,N_6177,N_11165);
or U12235 (N_12235,N_10256,N_6446);
or U12236 (N_12236,N_6114,N_9473);
nand U12237 (N_12237,N_6307,N_11905);
or U12238 (N_12238,N_9113,N_10148);
nor U12239 (N_12239,N_7739,N_7766);
or U12240 (N_12240,N_7649,N_8897);
or U12241 (N_12241,N_10259,N_6314);
nor U12242 (N_12242,N_7920,N_8700);
and U12243 (N_12243,N_11552,N_6368);
nor U12244 (N_12244,N_11036,N_8824);
and U12245 (N_12245,N_8748,N_9861);
nor U12246 (N_12246,N_7292,N_11093);
xor U12247 (N_12247,N_10764,N_7106);
or U12248 (N_12248,N_7280,N_7790);
nand U12249 (N_12249,N_8291,N_8842);
nand U12250 (N_12250,N_9815,N_8367);
xor U12251 (N_12251,N_10449,N_7670);
or U12252 (N_12252,N_11948,N_6735);
nor U12253 (N_12253,N_7250,N_8964);
and U12254 (N_12254,N_9600,N_10014);
and U12255 (N_12255,N_8535,N_10653);
or U12256 (N_12256,N_10898,N_8986);
xor U12257 (N_12257,N_11310,N_6926);
nand U12258 (N_12258,N_7527,N_7036);
nand U12259 (N_12259,N_6541,N_6691);
nor U12260 (N_12260,N_11998,N_8823);
nand U12261 (N_12261,N_7007,N_9066);
or U12262 (N_12262,N_6335,N_6914);
nand U12263 (N_12263,N_10933,N_6370);
or U12264 (N_12264,N_10732,N_6566);
nand U12265 (N_12265,N_8357,N_7150);
or U12266 (N_12266,N_9587,N_7637);
or U12267 (N_12267,N_7398,N_11055);
nor U12268 (N_12268,N_7112,N_9873);
or U12269 (N_12269,N_8486,N_6898);
or U12270 (N_12270,N_8892,N_10294);
or U12271 (N_12271,N_8517,N_11244);
nand U12272 (N_12272,N_6346,N_10641);
or U12273 (N_12273,N_6650,N_7860);
xor U12274 (N_12274,N_10124,N_9484);
nand U12275 (N_12275,N_10968,N_7763);
or U12276 (N_12276,N_7070,N_7999);
nor U12277 (N_12277,N_7202,N_9267);
xor U12278 (N_12278,N_9352,N_10931);
or U12279 (N_12279,N_9632,N_10645);
or U12280 (N_12280,N_8718,N_6462);
nor U12281 (N_12281,N_10874,N_7438);
xnor U12282 (N_12282,N_7277,N_7403);
nand U12283 (N_12283,N_8639,N_10576);
xor U12284 (N_12284,N_7130,N_11295);
and U12285 (N_12285,N_10171,N_7622);
or U12286 (N_12286,N_9551,N_10391);
nand U12287 (N_12287,N_11806,N_10389);
nand U12288 (N_12288,N_9123,N_9940);
nor U12289 (N_12289,N_9143,N_9331);
nand U12290 (N_12290,N_6553,N_10774);
nand U12291 (N_12291,N_11522,N_11710);
nor U12292 (N_12292,N_7953,N_7884);
xnor U12293 (N_12293,N_10840,N_9494);
nand U12294 (N_12294,N_9527,N_8004);
and U12295 (N_12295,N_9450,N_8340);
and U12296 (N_12296,N_8632,N_6029);
or U12297 (N_12297,N_8478,N_9410);
and U12298 (N_12298,N_8702,N_9307);
and U12299 (N_12299,N_9868,N_10627);
and U12300 (N_12300,N_6758,N_6285);
nand U12301 (N_12301,N_9025,N_9693);
and U12302 (N_12302,N_8334,N_11987);
xor U12303 (N_12303,N_6109,N_9365);
xnor U12304 (N_12304,N_8565,N_8140);
or U12305 (N_12305,N_9552,N_7109);
nor U12306 (N_12306,N_9951,N_11266);
nand U12307 (N_12307,N_6207,N_7972);
xor U12308 (N_12308,N_9579,N_6502);
and U12309 (N_12309,N_7563,N_7120);
and U12310 (N_12310,N_10040,N_8428);
nor U12311 (N_12311,N_6513,N_10153);
nand U12312 (N_12312,N_10317,N_9675);
and U12313 (N_12313,N_11054,N_8872);
or U12314 (N_12314,N_7584,N_7743);
and U12315 (N_12315,N_10999,N_11232);
nand U12316 (N_12316,N_8542,N_8177);
nor U12317 (N_12317,N_11173,N_9800);
nor U12318 (N_12318,N_10526,N_11953);
nand U12319 (N_12319,N_10958,N_11569);
xnor U12320 (N_12320,N_6963,N_10560);
and U12321 (N_12321,N_10481,N_9972);
nor U12322 (N_12322,N_8883,N_8173);
and U12323 (N_12323,N_10728,N_10105);
or U12324 (N_12324,N_7161,N_11560);
xnor U12325 (N_12325,N_9167,N_7862);
nor U12326 (N_12326,N_9159,N_6583);
nor U12327 (N_12327,N_6007,N_10400);
nor U12328 (N_12328,N_11645,N_6581);
or U12329 (N_12329,N_9890,N_11185);
nand U12330 (N_12330,N_10234,N_9945);
nor U12331 (N_12331,N_10388,N_8816);
and U12332 (N_12332,N_7010,N_10166);
or U12333 (N_12333,N_8796,N_7904);
and U12334 (N_12334,N_7441,N_11098);
and U12335 (N_12335,N_8396,N_7388);
nor U12336 (N_12336,N_10087,N_8490);
and U12337 (N_12337,N_7460,N_8633);
nand U12338 (N_12338,N_7127,N_8052);
and U12339 (N_12339,N_6154,N_11110);
and U12340 (N_12340,N_11840,N_10353);
and U12341 (N_12341,N_7648,N_8944);
or U12342 (N_12342,N_7408,N_7430);
nor U12343 (N_12343,N_8247,N_8029);
nand U12344 (N_12344,N_10325,N_7484);
nor U12345 (N_12345,N_10680,N_7727);
or U12346 (N_12346,N_6960,N_11500);
and U12347 (N_12347,N_9077,N_11925);
and U12348 (N_12348,N_8261,N_8735);
nand U12349 (N_12349,N_7658,N_7769);
nand U12350 (N_12350,N_6765,N_6118);
xnor U12351 (N_12351,N_10016,N_11418);
nand U12352 (N_12352,N_7825,N_11979);
nor U12353 (N_12353,N_11477,N_9602);
or U12354 (N_12354,N_10542,N_7318);
nor U12355 (N_12355,N_9462,N_8241);
or U12356 (N_12356,N_11465,N_10802);
or U12357 (N_12357,N_9644,N_6113);
or U12358 (N_12358,N_10424,N_9811);
nand U12359 (N_12359,N_8598,N_6874);
and U12360 (N_12360,N_9381,N_7672);
nor U12361 (N_12361,N_9993,N_6125);
xnor U12362 (N_12362,N_10899,N_7887);
or U12363 (N_12363,N_8981,N_11342);
xnor U12364 (N_12364,N_11737,N_7291);
nor U12365 (N_12365,N_9054,N_6153);
and U12366 (N_12366,N_8682,N_7279);
or U12367 (N_12367,N_8481,N_11789);
nor U12368 (N_12368,N_7011,N_8151);
nand U12369 (N_12369,N_10012,N_10429);
or U12370 (N_12370,N_9910,N_10804);
and U12371 (N_12371,N_7452,N_9701);
and U12372 (N_12372,N_6030,N_9914);
or U12373 (N_12373,N_11867,N_11573);
nand U12374 (N_12374,N_9347,N_11388);
xnor U12375 (N_12375,N_11546,N_10128);
nand U12376 (N_12376,N_11043,N_6321);
and U12377 (N_12377,N_8495,N_6700);
and U12378 (N_12378,N_6169,N_8407);
nand U12379 (N_12379,N_6721,N_8468);
nor U12380 (N_12380,N_9967,N_11805);
nand U12381 (N_12381,N_11832,N_9417);
and U12382 (N_12382,N_9323,N_8251);
nor U12383 (N_12383,N_8246,N_9029);
nand U12384 (N_12384,N_7428,N_10321);
nand U12385 (N_12385,N_11721,N_10363);
nor U12386 (N_12386,N_6225,N_8516);
or U12387 (N_12387,N_6821,N_11130);
nand U12388 (N_12388,N_11498,N_6373);
nand U12389 (N_12389,N_11122,N_8305);
nand U12390 (N_12390,N_6930,N_8924);
nor U12391 (N_12391,N_7754,N_7881);
or U12392 (N_12392,N_9599,N_9789);
nor U12393 (N_12393,N_7747,N_8726);
nor U12394 (N_12394,N_8315,N_9097);
or U12395 (N_12395,N_11624,N_9837);
nor U12396 (N_12396,N_7874,N_8677);
nand U12397 (N_12397,N_6740,N_9344);
nor U12398 (N_12398,N_7715,N_11913);
nor U12399 (N_12399,N_11437,N_8859);
nand U12400 (N_12400,N_11907,N_6745);
nor U12401 (N_12401,N_7638,N_11517);
and U12402 (N_12402,N_7575,N_8768);
or U12403 (N_12403,N_8782,N_8758);
nor U12404 (N_12404,N_6825,N_8778);
xor U12405 (N_12405,N_8553,N_7463);
or U12406 (N_12406,N_6041,N_6339);
nand U12407 (N_12407,N_9574,N_10214);
and U12408 (N_12408,N_8212,N_7897);
or U12409 (N_12409,N_7564,N_8581);
xor U12410 (N_12410,N_8227,N_10673);
and U12411 (N_12411,N_9893,N_6641);
nor U12412 (N_12412,N_11715,N_10445);
or U12413 (N_12413,N_10139,N_10426);
or U12414 (N_12414,N_6632,N_9812);
or U12415 (N_12415,N_6724,N_9750);
and U12416 (N_12416,N_7684,N_10084);
and U12417 (N_12417,N_9523,N_8836);
or U12418 (N_12418,N_10431,N_8838);
xor U12419 (N_12419,N_10989,N_11495);
nor U12420 (N_12420,N_6128,N_9188);
and U12421 (N_12421,N_8368,N_6998);
xor U12422 (N_12422,N_7016,N_10547);
or U12423 (N_12423,N_8443,N_8825);
and U12424 (N_12424,N_11440,N_6313);
and U12425 (N_12425,N_7962,N_7360);
and U12426 (N_12426,N_9853,N_8033);
and U12427 (N_12427,N_11396,N_8072);
nor U12428 (N_12428,N_11026,N_8962);
or U12429 (N_12429,N_8732,N_8733);
or U12430 (N_12430,N_8644,N_8578);
and U12431 (N_12431,N_7633,N_8057);
nand U12432 (N_12432,N_7008,N_9011);
or U12433 (N_12433,N_9948,N_9246);
or U12434 (N_12434,N_6204,N_10563);
or U12435 (N_12435,N_10647,N_11930);
and U12436 (N_12436,N_6320,N_9205);
and U12437 (N_12437,N_11410,N_10772);
nor U12438 (N_12438,N_11001,N_9846);
or U12439 (N_12439,N_11475,N_7406);
or U12440 (N_12440,N_11190,N_6475);
nor U12441 (N_12441,N_6907,N_11415);
and U12442 (N_12442,N_7420,N_9927);
nand U12443 (N_12443,N_11205,N_11073);
or U12444 (N_12444,N_11152,N_8570);
nor U12445 (N_12445,N_11170,N_7728);
xnor U12446 (N_12446,N_7651,N_10644);
and U12447 (N_12447,N_9624,N_10097);
nand U12448 (N_12448,N_10498,N_10187);
nor U12449 (N_12449,N_11813,N_6115);
or U12450 (N_12450,N_7764,N_10442);
nand U12451 (N_12451,N_7528,N_9364);
and U12452 (N_12452,N_6820,N_6794);
nand U12453 (N_12453,N_10031,N_7772);
and U12454 (N_12454,N_6890,N_9592);
or U12455 (N_12455,N_6328,N_9408);
nand U12456 (N_12456,N_9309,N_11894);
and U12457 (N_12457,N_8380,N_9095);
or U12458 (N_12458,N_6634,N_11997);
or U12459 (N_12459,N_10038,N_8138);
or U12460 (N_12460,N_11960,N_11121);
nor U12461 (N_12461,N_7949,N_6392);
or U12462 (N_12462,N_6485,N_9052);
nand U12463 (N_12463,N_8960,N_11182);
and U12464 (N_12464,N_10856,N_8411);
or U12465 (N_12465,N_8003,N_11897);
or U12466 (N_12466,N_11433,N_11123);
xnor U12467 (N_12467,N_9206,N_7311);
nor U12468 (N_12468,N_9835,N_6938);
xor U12469 (N_12469,N_11921,N_8783);
nor U12470 (N_12470,N_9770,N_7905);
nand U12471 (N_12471,N_6718,N_6858);
nor U12472 (N_12472,N_10872,N_11512);
and U12473 (N_12473,N_7447,N_9613);
or U12474 (N_12474,N_10245,N_11906);
nor U12475 (N_12475,N_6885,N_7802);
nand U12476 (N_12476,N_10337,N_8712);
xor U12477 (N_12477,N_9554,N_6636);
or U12478 (N_12478,N_6579,N_10028);
nor U12479 (N_12479,N_8301,N_11324);
and U12480 (N_12480,N_11153,N_11591);
nand U12481 (N_12481,N_10345,N_10086);
nor U12482 (N_12482,N_9917,N_8851);
or U12483 (N_12483,N_9176,N_8728);
nor U12484 (N_12484,N_8304,N_10991);
or U12485 (N_12485,N_7005,N_7938);
or U12486 (N_12486,N_8763,N_8323);
nand U12487 (N_12487,N_7134,N_11716);
and U12488 (N_12488,N_9705,N_7259);
or U12489 (N_12489,N_6793,N_8865);
and U12490 (N_12490,N_6709,N_8905);
nor U12491 (N_12491,N_10160,N_9528);
nand U12492 (N_12492,N_10428,N_6951);
nor U12493 (N_12493,N_9193,N_8657);
nor U12494 (N_12494,N_10420,N_9088);
nand U12495 (N_12495,N_7182,N_10466);
nand U12496 (N_12496,N_6185,N_9458);
or U12497 (N_12497,N_6470,N_11888);
and U12498 (N_12498,N_8868,N_10297);
and U12499 (N_12499,N_9611,N_11214);
xor U12500 (N_12500,N_8513,N_9690);
xnor U12501 (N_12501,N_10724,N_10438);
nand U12502 (N_12502,N_6474,N_11853);
or U12503 (N_12503,N_7114,N_7610);
or U12504 (N_12504,N_7236,N_8899);
nand U12505 (N_12505,N_10240,N_8116);
and U12506 (N_12506,N_7589,N_7614);
or U12507 (N_12507,N_11594,N_9313);
nand U12508 (N_12508,N_11134,N_7736);
nor U12509 (N_12509,N_9446,N_6602);
and U12510 (N_12510,N_7845,N_8496);
and U12511 (N_12511,N_11585,N_6270);
nor U12512 (N_12512,N_8484,N_9746);
xnor U12513 (N_12513,N_6011,N_7372);
nand U12514 (N_12514,N_8293,N_10730);
nor U12515 (N_12515,N_10718,N_9047);
or U12516 (N_12516,N_7669,N_11730);
nand U12517 (N_12517,N_7572,N_11225);
nand U12518 (N_12518,N_11803,N_11643);
xor U12519 (N_12519,N_8285,N_7910);
nand U12520 (N_12520,N_11941,N_6591);
nor U12521 (N_12521,N_9175,N_7267);
xnor U12522 (N_12522,N_11347,N_11821);
xor U12523 (N_12523,N_11072,N_10089);
nor U12524 (N_12524,N_9971,N_6216);
nor U12525 (N_12525,N_6341,N_8550);
xnor U12526 (N_12526,N_8837,N_9186);
or U12527 (N_12527,N_7214,N_9651);
nand U12528 (N_12528,N_8087,N_9553);
or U12529 (N_12529,N_7402,N_8773);
xor U12530 (N_12530,N_6058,N_6403);
and U12531 (N_12531,N_6624,N_9124);
nand U12532 (N_12532,N_9828,N_9918);
nor U12533 (N_12533,N_8299,N_8379);
nor U12534 (N_12534,N_8180,N_8548);
nor U12535 (N_12535,N_8410,N_9928);
nor U12536 (N_12536,N_7157,N_6174);
and U12537 (N_12537,N_8696,N_7674);
and U12538 (N_12538,N_6638,N_6565);
and U12539 (N_12539,N_9799,N_11038);
nor U12540 (N_12540,N_10282,N_11135);
and U12541 (N_12541,N_10665,N_10752);
nand U12542 (N_12542,N_7559,N_11974);
nor U12543 (N_12543,N_9731,N_9984);
and U12544 (N_12544,N_8337,N_6189);
nor U12545 (N_12545,N_8211,N_10298);
and U12546 (N_12546,N_8132,N_9886);
and U12547 (N_12547,N_10225,N_6977);
nor U12548 (N_12548,N_9315,N_10699);
nor U12549 (N_12549,N_7284,N_7066);
xor U12550 (N_12550,N_8390,N_8545);
and U12551 (N_12551,N_7162,N_11740);
nor U12552 (N_12552,N_9049,N_6221);
xnor U12553 (N_12553,N_6451,N_8911);
or U12554 (N_12554,N_8747,N_7912);
nand U12555 (N_12555,N_11506,N_11564);
xor U12556 (N_12556,N_7915,N_11949);
and U12557 (N_12557,N_9396,N_7359);
or U12558 (N_12558,N_8104,N_11712);
nand U12559 (N_12559,N_10561,N_8055);
nor U12560 (N_12560,N_6731,N_9862);
or U12561 (N_12561,N_10383,N_7253);
or U12562 (N_12562,N_6349,N_9838);
nand U12563 (N_12563,N_10876,N_11528);
nand U12564 (N_12564,N_11954,N_6102);
nor U12565 (N_12565,N_10066,N_10869);
xnor U12566 (N_12566,N_6843,N_7828);
and U12567 (N_12567,N_6132,N_9662);
nand U12568 (N_12568,N_8375,N_7877);
or U12569 (N_12569,N_6202,N_7180);
nand U12570 (N_12570,N_9299,N_7989);
nand U12571 (N_12571,N_10365,N_7165);
nand U12572 (N_12572,N_8111,N_10335);
nand U12573 (N_12573,N_11617,N_10177);
nand U12574 (N_12574,N_8877,N_10161);
or U12575 (N_12575,N_9027,N_10268);
nand U12576 (N_12576,N_7992,N_11279);
and U12577 (N_12577,N_11838,N_6463);
or U12578 (N_12578,N_7732,N_9615);
or U12579 (N_12579,N_10186,N_9511);
or U12580 (N_12580,N_8143,N_8306);
or U12581 (N_12581,N_6263,N_9894);
nor U12582 (N_12582,N_9779,N_7981);
nor U12583 (N_12583,N_11880,N_9964);
and U12584 (N_12584,N_10032,N_11330);
and U12585 (N_12585,N_9301,N_6364);
and U12586 (N_12586,N_7338,N_7439);
and U12587 (N_12587,N_11024,N_9305);
xnor U12588 (N_12588,N_7198,N_6434);
nor U12589 (N_12589,N_7183,N_11076);
and U12590 (N_12590,N_10799,N_11982);
nand U12591 (N_12591,N_9103,N_11315);
or U12592 (N_12592,N_6802,N_6835);
nand U12593 (N_12593,N_6606,N_8922);
nor U12594 (N_12594,N_6305,N_7786);
or U12595 (N_12595,N_8571,N_11215);
nor U12596 (N_12596,N_8818,N_10888);
or U12597 (N_12597,N_10299,N_10796);
and U12598 (N_12598,N_7823,N_9415);
nor U12599 (N_12599,N_9618,N_8343);
and U12600 (N_12600,N_6004,N_10592);
nor U12601 (N_12601,N_9712,N_8715);
nor U12602 (N_12602,N_11797,N_8083);
and U12603 (N_12603,N_11049,N_11903);
nor U12604 (N_12604,N_9764,N_7045);
nor U12605 (N_12605,N_10748,N_11322);
nor U12606 (N_12606,N_9844,N_10281);
or U12607 (N_12607,N_11652,N_11040);
nand U12608 (N_12608,N_7532,N_8152);
and U12609 (N_12609,N_11442,N_6516);
or U12610 (N_12610,N_11770,N_9280);
or U12611 (N_12611,N_8090,N_9563);
or U12612 (N_12612,N_10776,N_7028);
and U12613 (N_12613,N_7683,N_7108);
nor U12614 (N_12614,N_8497,N_8755);
nand U12615 (N_12615,N_6481,N_9032);
nand U12616 (N_12616,N_6807,N_11194);
nand U12617 (N_12617,N_7578,N_10663);
or U12618 (N_12618,N_7921,N_6297);
xnor U12619 (N_12619,N_11337,N_7700);
and U12620 (N_12620,N_9059,N_7305);
nor U12621 (N_12621,N_6394,N_10624);
nand U12622 (N_12622,N_6139,N_8769);
xor U12623 (N_12623,N_8102,N_11136);
and U12624 (N_12624,N_9685,N_7095);
nand U12625 (N_12625,N_11957,N_6706);
nand U12626 (N_12626,N_10470,N_7335);
nand U12627 (N_12627,N_8686,N_10157);
or U12628 (N_12628,N_9329,N_8853);
nand U12629 (N_12629,N_10377,N_8117);
and U12630 (N_12630,N_7699,N_8263);
nor U12631 (N_12631,N_7358,N_10250);
nor U12632 (N_12632,N_10085,N_11372);
and U12633 (N_12633,N_10711,N_10111);
and U12634 (N_12634,N_11691,N_8355);
xor U12635 (N_12635,N_7231,N_7324);
nor U12636 (N_12636,N_9112,N_9766);
nand U12637 (N_12637,N_11800,N_11733);
or U12638 (N_12638,N_6981,N_7675);
or U12639 (N_12639,N_11958,N_9076);
and U12640 (N_12640,N_10421,N_11254);
or U12641 (N_12641,N_9368,N_9218);
nor U12642 (N_12642,N_7840,N_8112);
and U12643 (N_12643,N_11207,N_8710);
and U12644 (N_12644,N_11945,N_7493);
nor U12645 (N_12645,N_6244,N_8329);
and U12646 (N_12646,N_9780,N_6791);
and U12647 (N_12647,N_6279,N_6044);
or U12648 (N_12648,N_10165,N_11235);
nor U12649 (N_12649,N_11118,N_9898);
nand U12650 (N_12650,N_9262,N_6988);
nand U12651 (N_12651,N_9128,N_9876);
and U12652 (N_12652,N_7520,N_7931);
and U12653 (N_12653,N_11250,N_11200);
or U12654 (N_12654,N_6797,N_7310);
nand U12655 (N_12655,N_10554,N_10669);
nor U12656 (N_12656,N_11532,N_6524);
and U12657 (N_12657,N_9355,N_10030);
or U12658 (N_12658,N_7856,N_8038);
and U12659 (N_12659,N_7319,N_6040);
or U12660 (N_12660,N_10584,N_11287);
or U12661 (N_12661,N_8879,N_9840);
nor U12662 (N_12662,N_8729,N_10857);
or U12663 (N_12663,N_10710,N_9700);
nand U12664 (N_12664,N_10902,N_10275);
nor U12665 (N_12665,N_9772,N_11233);
nand U12666 (N_12666,N_9909,N_9708);
nand U12667 (N_12667,N_11483,N_8646);
nand U12668 (N_12668,N_8011,N_9698);
or U12669 (N_12669,N_11241,N_6728);
or U12670 (N_12670,N_6830,N_9546);
or U12671 (N_12671,N_10763,N_8454);
nor U12672 (N_12672,N_6022,N_10306);
xnor U12673 (N_12673,N_9024,N_11686);
nand U12674 (N_12674,N_7102,N_6725);
or U12675 (N_12675,N_8183,N_6488);
nand U12676 (N_12676,N_10882,N_10338);
nand U12677 (N_12677,N_10932,N_8611);
nand U12678 (N_12678,N_10726,N_8684);
nand U12679 (N_12679,N_10350,N_7387);
nor U12680 (N_12680,N_10129,N_6312);
or U12681 (N_12681,N_9520,N_6855);
nand U12682 (N_12682,N_8121,N_9607);
nor U12683 (N_12683,N_7933,N_8316);
nor U12684 (N_12684,N_10701,N_7852);
nor U12685 (N_12685,N_7913,N_10501);
and U12686 (N_12686,N_7782,N_10960);
xor U12687 (N_12687,N_11722,N_8978);
or U12688 (N_12688,N_11434,N_6841);
nand U12689 (N_12689,N_8554,N_7156);
nand U12690 (N_12690,N_7596,N_11416);
or U12691 (N_12691,N_9728,N_6871);
nand U12692 (N_12692,N_9621,N_11748);
or U12693 (N_12693,N_6592,N_11767);
and U12694 (N_12694,N_8501,N_6943);
nor U12695 (N_12695,N_9716,N_7024);
nand U12696 (N_12696,N_10677,N_11896);
xnor U12697 (N_12697,N_8391,N_10994);
or U12698 (N_12698,N_9570,N_6607);
or U12699 (N_12699,N_10236,N_9684);
and U12700 (N_12700,N_7590,N_11060);
nand U12701 (N_12701,N_9225,N_6353);
nand U12702 (N_12702,N_10814,N_8053);
nand U12703 (N_12703,N_10054,N_9348);
nand U12704 (N_12704,N_7744,N_9545);
nand U12705 (N_12705,N_8237,N_10521);
or U12706 (N_12706,N_11758,N_10230);
nand U12707 (N_12707,N_7903,N_8990);
xor U12708 (N_12708,N_7607,N_6754);
and U12709 (N_12709,N_10536,N_9555);
nand U12710 (N_12710,N_8226,N_10749);
nor U12711 (N_12711,N_8736,N_6824);
or U12712 (N_12712,N_6883,N_11499);
or U12713 (N_12713,N_6899,N_9345);
and U12714 (N_12714,N_10525,N_6667);
or U12715 (N_12715,N_9031,N_9424);
nand U12716 (N_12716,N_8421,N_7082);
xor U12717 (N_12717,N_10731,N_8268);
or U12718 (N_12718,N_6644,N_9070);
or U12719 (N_12719,N_6967,N_7332);
or U12720 (N_12720,N_7051,N_8080);
or U12721 (N_12721,N_10723,N_9582);
nor U12722 (N_12722,N_8063,N_9151);
and U12723 (N_12723,N_8073,N_6409);
xor U12724 (N_12724,N_8219,N_8044);
nor U12725 (N_12725,N_7333,N_6359);
nand U12726 (N_12726,N_7552,N_6246);
nor U12727 (N_12727,N_7422,N_8889);
nand U12728 (N_12728,N_10096,N_8687);
and U12729 (N_12729,N_8970,N_8106);
or U12730 (N_12730,N_9488,N_9950);
nor U12731 (N_12731,N_7124,N_10020);
or U12732 (N_12732,N_10468,N_9376);
nand U12733 (N_12733,N_6054,N_11070);
xnor U12734 (N_12734,N_11431,N_6857);
or U12735 (N_12735,N_8196,N_11962);
or U12736 (N_12736,N_11717,N_10533);
or U12737 (N_12737,N_6471,N_11090);
xnor U12738 (N_12738,N_6075,N_8018);
or U12739 (N_12739,N_9387,N_9447);
nand U12740 (N_12740,N_8008,N_6256);
nor U12741 (N_12741,N_11924,N_6317);
xnor U12742 (N_12742,N_11587,N_6278);
and U12743 (N_12743,N_7839,N_7019);
nand U12744 (N_12744,N_11589,N_6127);
nor U12745 (N_12745,N_11259,N_10422);
xnor U12746 (N_12746,N_7612,N_6917);
nand U12747 (N_12747,N_9966,N_6089);
nor U12748 (N_12748,N_8455,N_9019);
or U12749 (N_12749,N_11099,N_11260);
and U12750 (N_12750,N_7661,N_9922);
nand U12751 (N_12751,N_10102,N_9290);
xnor U12752 (N_12752,N_9489,N_9518);
or U12753 (N_12753,N_10264,N_6017);
and U12754 (N_12754,N_7211,N_8099);
and U12755 (N_12755,N_11106,N_10714);
nand U12756 (N_12756,N_8077,N_6365);
nand U12757 (N_12757,N_10191,N_10529);
nor U12758 (N_12758,N_7526,N_8638);
nand U12759 (N_12759,N_6908,N_7087);
or U12760 (N_12760,N_8573,N_8400);
and U12761 (N_12761,N_8993,N_9213);
xor U12762 (N_12762,N_8683,N_9818);
xor U12763 (N_12763,N_8800,N_7696);
nand U12764 (N_12764,N_10454,N_6426);
nor U12765 (N_12765,N_10630,N_11726);
or U12766 (N_12766,N_7176,N_8154);
xnor U12767 (N_12767,N_7847,N_10207);
xor U12768 (N_12768,N_9854,N_7833);
nor U12769 (N_12769,N_11338,N_7383);
or U12770 (N_12770,N_9994,N_6922);
or U12771 (N_12771,N_10531,N_11659);
xor U12772 (N_12772,N_10024,N_11380);
or U12773 (N_12773,N_8403,N_11107);
nand U12774 (N_12774,N_11449,N_6049);
nor U12775 (N_12775,N_8968,N_9792);
and U12776 (N_12776,N_7343,N_6688);
and U12777 (N_12777,N_9135,N_10900);
and U12778 (N_12778,N_10133,N_7449);
xnor U12779 (N_12779,N_7673,N_6331);
and U12780 (N_12780,N_10193,N_10705);
and U12781 (N_12781,N_9942,N_11870);
or U12782 (N_12782,N_10944,N_6327);
nor U12783 (N_12783,N_8743,N_11680);
nand U12784 (N_12784,N_10344,N_7927);
nand U12785 (N_12785,N_7268,N_7203);
nand U12786 (N_12786,N_11842,N_11775);
nand U12787 (N_12787,N_10471,N_11505);
and U12788 (N_12788,N_10146,N_7967);
or U12789 (N_12789,N_11304,N_11724);
nand U12790 (N_12790,N_9028,N_11729);
and U12791 (N_12791,N_10398,N_9514);
nor U12792 (N_12792,N_8345,N_8047);
or U12793 (N_12793,N_8579,N_7709);
or U12794 (N_12794,N_8927,N_7468);
nand U12795 (N_12795,N_10410,N_11900);
xnor U12796 (N_12796,N_11379,N_9878);
or U12797 (N_12797,N_11062,N_7163);
and U12798 (N_12798,N_9536,N_9830);
nand U12799 (N_12799,N_8602,N_11407);
or U12800 (N_12800,N_6085,N_8187);
or U12801 (N_12801,N_8035,N_11425);
and U12802 (N_12802,N_10921,N_7427);
nand U12803 (N_12803,N_6924,N_11727);
or U12804 (N_12804,N_11749,N_10373);
nor U12805 (N_12805,N_10569,N_8491);
nor U12806 (N_12806,N_11830,N_9487);
nor U12807 (N_12807,N_6045,N_8381);
xor U12808 (N_12808,N_10436,N_7685);
and U12809 (N_12809,N_9211,N_8980);
and U12810 (N_12810,N_11264,N_9882);
nand U12811 (N_12811,N_8489,N_6288);
nor U12812 (N_12812,N_7803,N_7773);
nor U12813 (N_12813,N_8155,N_8904);
nor U12814 (N_12814,N_6183,N_7506);
nor U12815 (N_12815,N_7364,N_7141);
or U12816 (N_12816,N_10792,N_6575);
nor U12817 (N_12817,N_10144,N_10657);
or U12818 (N_12818,N_6990,N_11271);
nor U12819 (N_12819,N_6236,N_8942);
or U12820 (N_12820,N_9057,N_6925);
and U12821 (N_12821,N_11640,N_6495);
and U12822 (N_12822,N_6847,N_8672);
or U12823 (N_12823,N_6016,N_7432);
nand U12824 (N_12824,N_8048,N_11458);
and U12825 (N_12825,N_6987,N_10913);
and U12826 (N_12826,N_11628,N_6795);
or U12827 (N_12827,N_10612,N_10132);
or U12828 (N_12828,N_6473,N_8600);
and U12829 (N_12829,N_7175,N_6992);
and U12830 (N_12830,N_7232,N_9260);
and U12831 (N_12831,N_6219,N_6333);
and U12832 (N_12832,N_6173,N_6240);
nand U12833 (N_12833,N_10512,N_9590);
and U12834 (N_12834,N_9265,N_8253);
and U12835 (N_12835,N_7771,N_8150);
nor U12836 (N_12836,N_9531,N_10806);
xor U12837 (N_12837,N_10156,N_11567);
xor U12838 (N_12838,N_6577,N_10860);
or U12839 (N_12839,N_8802,N_7271);
and U12840 (N_12840,N_6217,N_8014);
and U12841 (N_12841,N_6787,N_8583);
nand U12842 (N_12842,N_8156,N_8311);
and U12843 (N_12843,N_6358,N_6310);
or U12844 (N_12844,N_9096,N_11142);
xnor U12845 (N_12845,N_8243,N_6491);
nand U12846 (N_12846,N_10356,N_8649);
xnor U12847 (N_12847,N_8234,N_8909);
and U12848 (N_12848,N_11610,N_10515);
nor U12849 (N_12849,N_9534,N_9222);
xor U12850 (N_12850,N_9444,N_6801);
nor U12851 (N_12851,N_10803,N_10467);
nand U12852 (N_12852,N_7587,N_11462);
and U12853 (N_12853,N_10519,N_10715);
nor U12854 (N_12854,N_11273,N_11212);
nor U12855 (N_12855,N_6543,N_7808);
nor U12856 (N_12856,N_9616,N_11184);
and U12857 (N_12857,N_10280,N_6621);
nor U12858 (N_12858,N_6628,N_7621);
nand U12859 (N_12859,N_6385,N_11595);
and U12860 (N_12860,N_8714,N_11819);
nor U12861 (N_12861,N_10393,N_8539);
and U12862 (N_12862,N_8377,N_11963);
nand U12863 (N_12863,N_9174,N_8371);
nand U12864 (N_12864,N_10817,N_6215);
or U12865 (N_12865,N_6069,N_11848);
nand U12866 (N_12866,N_9636,N_8009);
nor U12867 (N_12867,N_10196,N_6110);
nor U12868 (N_12868,N_9071,N_11698);
and U12869 (N_12869,N_11345,N_11649);
xor U12870 (N_12870,N_11364,N_6071);
and U12871 (N_12871,N_9625,N_11128);
or U12872 (N_12872,N_6864,N_11618);
or U12873 (N_12873,N_6736,N_6163);
and U12874 (N_12874,N_9575,N_7794);
or U12875 (N_12875,N_10272,N_6859);
nor U12876 (N_12876,N_11187,N_6486);
nand U12877 (N_12877,N_7140,N_6752);
or U12878 (N_12878,N_10970,N_7654);
nand U12879 (N_12879,N_11030,N_8900);
nor U12880 (N_12880,N_11771,N_6245);
or U12881 (N_12881,N_7896,N_10762);
xnor U12882 (N_12882,N_7000,N_6521);
nand U12883 (N_12883,N_8951,N_11786);
and U12884 (N_12884,N_6416,N_10249);
nor U12885 (N_12885,N_10866,N_6580);
or U12886 (N_12886,N_8587,N_10976);
and U12887 (N_12887,N_11255,N_11891);
nor U12888 (N_12888,N_8284,N_9099);
xnor U12889 (N_12889,N_6837,N_7539);
or U12890 (N_12890,N_10671,N_8867);
or U12891 (N_12891,N_10655,N_10367);
nor U12892 (N_12892,N_6799,N_11361);
xnor U12893 (N_12893,N_6087,N_10636);
nor U12894 (N_12894,N_7720,N_6284);
nand U12895 (N_12895,N_9742,N_10332);
and U12896 (N_12896,N_6950,N_6610);
and U12897 (N_12897,N_10990,N_11269);
or U12898 (N_12898,N_9362,N_8098);
or U12899 (N_12899,N_11989,N_6934);
nand U12900 (N_12900,N_10553,N_6573);
and U12901 (N_12901,N_7083,N_10822);
and U12902 (N_12902,N_7009,N_6116);
and U12903 (N_12903,N_11035,N_8973);
xor U12904 (N_12904,N_7425,N_6777);
xor U12905 (N_12905,N_11195,N_8425);
nor U12906 (N_12906,N_6053,N_9860);
nand U12907 (N_12907,N_11904,N_10596);
nand U12908 (N_12908,N_11466,N_11799);
nor U12909 (N_12909,N_10717,N_10646);
and U12910 (N_12910,N_10997,N_11554);
nand U12911 (N_12911,N_8167,N_6422);
and U12912 (N_12912,N_10205,N_10360);
and U12913 (N_12913,N_9482,N_9334);
and U12914 (N_12914,N_7450,N_11779);
nand U12915 (N_12915,N_9448,N_10348);
or U12916 (N_12916,N_7038,N_10517);
or U12917 (N_12917,N_6062,N_6894);
and U12918 (N_12918,N_8563,N_9442);
and U12919 (N_12919,N_11687,N_6982);
xnor U12920 (N_12920,N_9584,N_6048);
or U12921 (N_12921,N_8950,N_6697);
or U12922 (N_12922,N_9959,N_10093);
or U12923 (N_12923,N_11488,N_11818);
nand U12924 (N_12924,N_6501,N_11545);
nand U12925 (N_12925,N_7566,N_7624);
nor U12926 (N_12926,N_9429,N_6452);
nor U12927 (N_12927,N_10462,N_11362);
or U12928 (N_12928,N_9629,N_9672);
nand U12929 (N_12929,N_9241,N_7247);
nor U12930 (N_12930,N_11091,N_7459);
and U12931 (N_12931,N_11579,N_6904);
nand U12932 (N_12932,N_10403,N_6490);
and U12933 (N_12933,N_7665,N_6785);
or U12934 (N_12934,N_7846,N_8446);
or U12935 (N_12935,N_6712,N_6671);
or U12936 (N_12936,N_9490,N_10538);
nand U12937 (N_12937,N_9680,N_10000);
and U12938 (N_12938,N_11574,N_7655);
nor U12939 (N_12939,N_6838,N_7895);
or U12940 (N_12940,N_9093,N_8815);
and U12941 (N_12941,N_6569,N_6559);
nand U12942 (N_12942,N_7576,N_10439);
and U12943 (N_12943,N_10395,N_11993);
or U12944 (N_12944,N_6903,N_6507);
nand U12945 (N_12945,N_10935,N_11167);
or U12946 (N_12946,N_8202,N_10702);
and U12947 (N_12947,N_6431,N_10382);
nor U12948 (N_12948,N_10843,N_7942);
nand U12949 (N_12949,N_8192,N_8647);
nor U12950 (N_12950,N_6120,N_8576);
nand U12951 (N_12951,N_9238,N_9841);
xor U12952 (N_12952,N_8907,N_8266);
or U12953 (N_12953,N_9137,N_7868);
nand U12954 (N_12954,N_11701,N_6456);
nor U12955 (N_12955,N_8860,N_8625);
xnor U12956 (N_12956,N_11563,N_7128);
and U12957 (N_12957,N_6788,N_9126);
or U12958 (N_12958,N_10478,N_6266);
or U12959 (N_12959,N_7255,N_11868);
nor U12960 (N_12960,N_7984,N_10556);
nor U12961 (N_12961,N_6141,N_9919);
nor U12962 (N_12962,N_8660,N_6419);
and U12963 (N_12963,N_8472,N_8267);
and U12964 (N_12964,N_6013,N_7288);
and U12965 (N_12965,N_10745,N_7490);
and U12966 (N_12966,N_6097,N_11294);
and U12967 (N_12967,N_10278,N_6517);
nor U12968 (N_12968,N_11661,N_8257);
and U12969 (N_12969,N_7898,N_8533);
or U12970 (N_12970,N_7882,N_11209);
nor U12971 (N_12971,N_6545,N_7733);
nand U12972 (N_12972,N_7116,N_8544);
nand U12973 (N_12973,N_9787,N_8260);
or U12974 (N_12974,N_7393,N_7418);
or U12975 (N_12975,N_9836,N_6253);
and U12976 (N_12976,N_6230,N_8100);
xnor U12977 (N_12977,N_10686,N_10309);
or U12978 (N_12978,N_8781,N_7352);
nor U12979 (N_12979,N_8230,N_10524);
nor U12980 (N_12980,N_9907,N_10469);
nor U12981 (N_12981,N_10474,N_9091);
and U12982 (N_12982,N_7044,N_11646);
or U12983 (N_12983,N_10455,N_8937);
nor U12984 (N_12984,N_11258,N_6522);
or U12985 (N_12985,N_9783,N_10407);
nand U12986 (N_12986,N_11313,N_10116);
nor U12987 (N_12987,N_10879,N_6417);
or U12988 (N_12988,N_8423,N_10993);
xor U12989 (N_12989,N_8965,N_11261);
and U12990 (N_12990,N_8309,N_10380);
nand U12991 (N_12991,N_8762,N_9997);
or U12992 (N_12992,N_11159,N_11031);
nor U12993 (N_12993,N_7206,N_6384);
and U12994 (N_12994,N_10982,N_11460);
xor U12995 (N_12995,N_9165,N_9466);
nor U12996 (N_12996,N_8225,N_7582);
or U12997 (N_12997,N_8059,N_6786);
nor U12998 (N_12998,N_10925,N_9242);
nand U12999 (N_12999,N_8691,N_10602);
and U13000 (N_13000,N_10025,N_9640);
nand U13001 (N_13001,N_10179,N_7734);
or U13002 (N_13002,N_9969,N_8378);
and U13003 (N_13003,N_11471,N_10959);
or U13004 (N_13004,N_11636,N_9302);
xnor U13005 (N_13005,N_8256,N_9372);
nor U13006 (N_13006,N_7977,N_10476);
and U13007 (N_13007,N_11883,N_10465);
or U13008 (N_13008,N_8984,N_6034);
nor U13009 (N_13009,N_10246,N_9719);
or U13010 (N_13010,N_8656,N_6014);
nor U13011 (N_13011,N_6976,N_11470);
or U13012 (N_13012,N_6150,N_11201);
nand U13013 (N_13013,N_6375,N_8184);
nand U13014 (N_13014,N_11481,N_11400);
nand U13015 (N_13015,N_6729,N_9637);
or U13016 (N_13016,N_11245,N_7908);
or U13017 (N_13017,N_7939,N_10548);
and U13018 (N_13018,N_10231,N_10740);
and U13019 (N_13019,N_10727,N_9814);
xor U13020 (N_13020,N_11473,N_10537);
and U13021 (N_13021,N_8850,N_9240);
nand U13022 (N_13022,N_10131,N_6670);
nor U13023 (N_13023,N_6282,N_6818);
or U13024 (N_13024,N_6046,N_7482);
nand U13025 (N_13025,N_11745,N_8507);
and U13026 (N_13026,N_10019,N_7746);
nor U13027 (N_13027,N_9326,N_6957);
or U13028 (N_13028,N_6809,N_8398);
or U13029 (N_13029,N_9461,N_10340);
and U13030 (N_13030,N_7756,N_6995);
or U13031 (N_13031,N_9102,N_11231);
nor U13032 (N_13032,N_8988,N_8606);
nand U13033 (N_13033,N_11777,N_9435);
nand U13034 (N_13034,N_7216,N_8935);
nand U13035 (N_13035,N_11889,N_11928);
nand U13036 (N_13036,N_10951,N_10396);
or U13037 (N_13037,N_11289,N_10558);
and U13038 (N_13038,N_11268,N_9595);
or U13039 (N_13039,N_9704,N_10985);
or U13040 (N_13040,N_7497,N_7380);
or U13041 (N_13041,N_7641,N_7229);
nor U13042 (N_13042,N_11248,N_7145);
nand U13043 (N_13043,N_10035,N_6078);
and U13044 (N_13044,N_6056,N_9492);
and U13045 (N_13045,N_9832,N_7384);
xor U13046 (N_13046,N_7783,N_8204);
nor U13047 (N_13047,N_7221,N_7196);
xnor U13048 (N_13048,N_6738,N_9562);
nor U13049 (N_13049,N_8105,N_11688);
xor U13050 (N_13050,N_9604,N_9419);
nand U13051 (N_13051,N_6477,N_11353);
or U13052 (N_13052,N_9677,N_7721);
nor U13053 (N_13053,N_9687,N_6562);
nor U13054 (N_13054,N_7892,N_10300);
nor U13055 (N_13055,N_7894,N_7067);
or U13056 (N_13056,N_10805,N_7726);
nand U13057 (N_13057,N_9291,N_8457);
or U13058 (N_13058,N_10095,N_10691);
nor U13059 (N_13059,N_10964,N_8286);
xnor U13060 (N_13060,N_10354,N_7168);
nand U13061 (N_13061,N_6572,N_8040);
xor U13062 (N_13062,N_7233,N_11397);
and U13063 (N_13063,N_6298,N_11057);
nor U13064 (N_13064,N_11764,N_10826);
nor U13065 (N_13065,N_11367,N_6918);
or U13066 (N_13066,N_9774,N_10725);
nand U13067 (N_13067,N_8078,N_9804);
or U13068 (N_13068,N_7289,N_7434);
nor U13069 (N_13069,N_8536,N_11675);
or U13070 (N_13070,N_7534,N_7695);
nand U13071 (N_13071,N_11336,N_7429);
and U13072 (N_13072,N_7049,N_10842);
nand U13073 (N_13073,N_8141,N_6283);
or U13074 (N_13074,N_11484,N_10495);
nor U13075 (N_13075,N_11732,N_11936);
and U13076 (N_13076,N_10107,N_9351);
or U13077 (N_13077,N_9650,N_6138);
nand U13078 (N_13078,N_8961,N_11132);
and U13079 (N_13079,N_10163,N_8694);
and U13080 (N_13080,N_6402,N_9156);
and U13081 (N_13081,N_7605,N_8074);
nor U13082 (N_13082,N_6179,N_7386);
nand U13083 (N_13083,N_11923,N_7735);
nor U13084 (N_13084,N_10807,N_11520);
xnor U13085 (N_13085,N_6036,N_9455);
or U13086 (N_13086,N_7598,N_6234);
nand U13087 (N_13087,N_8692,N_11521);
nor U13088 (N_13088,N_8604,N_11104);
and U13089 (N_13089,N_6679,N_11535);
and U13090 (N_13090,N_6999,N_10311);
and U13091 (N_13091,N_10162,N_8477);
nand U13092 (N_13092,N_9214,N_7199);
or U13093 (N_13093,N_9571,N_6161);
or U13094 (N_13094,N_7540,N_7982);
or U13095 (N_13095,N_10679,N_8131);
nand U13096 (N_13096,N_11547,N_8036);
or U13097 (N_13097,N_6849,N_11623);
nand U13098 (N_13098,N_7550,N_6039);
or U13099 (N_13099,N_10244,N_7682);
or U13100 (N_13100,N_8561,N_10357);
and U13101 (N_13101,N_9501,N_11349);
and U13102 (N_13102,N_11283,N_6151);
and U13103 (N_13103,N_6568,N_7238);
nor U13104 (N_13104,N_6869,N_10446);
nor U13105 (N_13105,N_11220,N_9061);
nor U13106 (N_13106,N_11609,N_8385);
nor U13107 (N_13107,N_9923,N_9906);
nor U13108 (N_13108,N_10006,N_9330);
and U13109 (N_13109,N_9643,N_11644);
or U13110 (N_13110,N_6395,N_8459);
and U13111 (N_13111,N_10260,N_8282);
or U13112 (N_13112,N_7784,N_7246);
nand U13113 (N_13113,N_10660,N_11298);
or U13114 (N_13114,N_9583,N_10637);
or U13115 (N_13115,N_6094,N_11665);
nor U13116 (N_13116,N_11835,N_7966);
and U13117 (N_13117,N_7512,N_6181);
nand U13118 (N_13118,N_10113,N_11509);
xor U13119 (N_13119,N_11899,N_9319);
xnor U13120 (N_13120,N_9382,N_9226);
nor U13121 (N_13121,N_9439,N_7464);
xor U13122 (N_13122,N_8833,N_9084);
or U13123 (N_13123,N_11390,N_10573);
and U13124 (N_13124,N_11881,N_7225);
or U13125 (N_13125,N_7906,N_8706);
and U13126 (N_13126,N_7561,N_7601);
nor U13127 (N_13127,N_10914,N_9141);
and U13128 (N_13128,N_10288,N_9686);
nand U13129 (N_13129,N_9177,N_7315);
nand U13130 (N_13130,N_6055,N_6135);
or U13131 (N_13131,N_11052,N_10330);
nor U13132 (N_13132,N_11087,N_10819);
and U13133 (N_13133,N_8858,N_8943);
or U13134 (N_13134,N_10492,N_6018);
nor U13135 (N_13135,N_10832,N_9569);
xor U13136 (N_13136,N_6713,N_8734);
nor U13137 (N_13137,N_6891,N_11782);
and U13138 (N_13138,N_11478,N_8420);
and U13139 (N_13139,N_10789,N_6148);
or U13140 (N_13140,N_6220,N_8624);
nor U13141 (N_13141,N_9619,N_8841);
nand U13142 (N_13142,N_7107,N_6750);
and U13143 (N_13143,N_11956,N_6260);
nor U13144 (N_13144,N_9252,N_10815);
nand U13145 (N_13145,N_9434,N_6854);
nand U13146 (N_13146,N_9871,N_6715);
nand U13147 (N_13147,N_8081,N_7328);
nand U13148 (N_13148,N_11183,N_8209);
and U13149 (N_13149,N_6232,N_6948);
nor U13150 (N_13150,N_9674,N_11177);
nand U13151 (N_13151,N_10273,N_7046);
nor U13152 (N_13152,N_11542,N_10448);
nand U13153 (N_13153,N_7492,N_11912);
or U13154 (N_13154,N_7235,N_6810);
nor U13155 (N_13155,N_8991,N_9508);
nor U13156 (N_13156,N_9310,N_9808);
xor U13157 (N_13157,N_9373,N_10837);
nand U13158 (N_13158,N_9769,N_7029);
nor U13159 (N_13159,N_6070,N_11864);
and U13160 (N_13160,N_9395,N_10381);
xor U13161 (N_13161,N_8502,N_8200);
xor U13162 (N_13162,N_8998,N_6267);
nor U13163 (N_13163,N_8705,N_6909);
or U13164 (N_13164,N_9451,N_8890);
or U13165 (N_13165,N_10621,N_6027);
and U13166 (N_13166,N_9386,N_7623);
nor U13167 (N_13167,N_8325,N_11236);
nand U13168 (N_13168,N_7222,N_7052);
or U13169 (N_13169,N_8913,N_6057);
nand U13170 (N_13170,N_9048,N_7789);
nand U13171 (N_13171,N_6239,N_11895);
nand U13172 (N_13172,N_7537,N_10203);
or U13173 (N_13173,N_9136,N_8721);
nand U13174 (N_13174,N_11578,N_8475);
nor U13175 (N_13175,N_8178,N_10094);
or U13176 (N_13176,N_9182,N_9452);
and U13177 (N_13177,N_8461,N_10983);
and U13178 (N_13178,N_9915,N_8231);
and U13179 (N_13179,N_6812,N_8342);
nor U13180 (N_13180,N_9371,N_8369);
xor U13181 (N_13181,N_7804,N_8277);
or U13182 (N_13182,N_10138,N_11872);
or U13183 (N_13183,N_8689,N_8678);
or U13184 (N_13184,N_7400,N_7543);
and U13185 (N_13185,N_6556,N_8603);
nor U13186 (N_13186,N_10823,N_6732);
and U13187 (N_13187,N_6447,N_7806);
or U13188 (N_13188,N_7212,N_9920);
nor U13189 (N_13189,N_6635,N_6876);
and U13190 (N_13190,N_8404,N_6906);
nand U13191 (N_13191,N_8399,N_10079);
or U13192 (N_13192,N_8946,N_7891);
and U13193 (N_13193,N_9614,N_8703);
xor U13194 (N_13194,N_11639,N_8679);
nor U13195 (N_13195,N_8338,N_7800);
nand U13196 (N_13196,N_8397,N_11599);
nor U13197 (N_13197,N_6684,N_11968);
and U13198 (N_13198,N_9394,N_9296);
nand U13199 (N_13199,N_6769,N_7698);
or U13200 (N_13200,N_6309,N_7412);
nand U13201 (N_13201,N_11707,N_11836);
nor U13202 (N_13202,N_8848,N_7788);
and U13203 (N_13203,N_6143,N_6535);
or U13204 (N_13204,N_7911,N_9233);
nor U13205 (N_13205,N_11873,N_11627);
nor U13206 (N_13206,N_9251,N_7074);
and U13207 (N_13207,N_6433,N_6261);
nand U13208 (N_13208,N_6355,N_6021);
nor U13209 (N_13209,N_8326,N_7930);
and U13210 (N_13210,N_6570,N_8730);
nand U13211 (N_13211,N_11371,N_10954);
nor U13212 (N_13212,N_8242,N_7266);
nor U13213 (N_13213,N_7934,N_9827);
and U13214 (N_13214,N_11871,N_6994);
nor U13215 (N_13215,N_6866,N_10683);
nor U13216 (N_13216,N_10782,N_6229);
and U13217 (N_13217,N_7824,N_9203);
and U13218 (N_13218,N_11631,N_9941);
or U13219 (N_13219,N_9630,N_7208);
or U13220 (N_13220,N_7717,N_6257);
xnor U13221 (N_13221,N_8869,N_8665);
or U13222 (N_13222,N_7062,N_8832);
nand U13223 (N_13223,N_6618,N_8361);
and U13224 (N_13224,N_7996,N_8605);
xor U13225 (N_13225,N_6629,N_8392);
nand U13226 (N_13226,N_6302,N_11972);
or U13227 (N_13227,N_7611,N_6255);
nand U13228 (N_13228,N_7997,N_9513);
xnor U13229 (N_13229,N_9670,N_8884);
nor U13230 (N_13230,N_10510,N_6599);
nand U13231 (N_13231,N_6719,N_7901);
or U13232 (N_13232,N_6687,N_9635);
nand U13233 (N_13233,N_10384,N_10908);
nand U13234 (N_13234,N_11723,N_7136);
nor U13235 (N_13235,N_11670,N_9848);
nand U13236 (N_13236,N_6780,N_6834);
or U13237 (N_13237,N_10212,N_8352);
and U13238 (N_13238,N_7423,N_10897);
and U13239 (N_13239,N_7986,N_6816);
and U13240 (N_13240,N_8746,N_8482);
nand U13241 (N_13241,N_9580,N_6469);
xor U13242 (N_13242,N_7170,N_7629);
and U13243 (N_13243,N_9747,N_7349);
nor U13244 (N_13244,N_6537,N_11222);
nor U13245 (N_13245,N_8780,N_7508);
and U13246 (N_13246,N_6711,N_6388);
nand U13247 (N_13247,N_9021,N_8406);
nand U13248 (N_13248,N_6693,N_11065);
nand U13249 (N_13249,N_6956,N_10110);
nor U13250 (N_13250,N_10188,N_7002);
and U13251 (N_13251,N_7579,N_9192);
nor U13252 (N_13252,N_7983,N_6945);
nand U13253 (N_13253,N_11762,N_10594);
nand U13254 (N_13254,N_11841,N_10623);
nand U13255 (N_13255,N_7880,N_6839);
nand U13256 (N_13256,N_11007,N_8941);
and U13257 (N_13257,N_11420,N_6848);
or U13258 (N_13258,N_8480,N_7810);
and U13259 (N_13259,N_11642,N_10527);
xor U13260 (N_13260,N_9254,N_8870);
or U13261 (N_13261,N_10629,N_7541);
xor U13262 (N_13262,N_6414,N_6158);
nor U13263 (N_13263,N_8082,N_11066);
and U13264 (N_13264,N_8939,N_9078);
nand U13265 (N_13265,N_11114,N_8931);
or U13266 (N_13266,N_11531,N_8966);
and U13267 (N_13267,N_8521,N_8067);
nor U13268 (N_13268,N_9145,N_9589);
nor U13269 (N_13269,N_7971,N_7722);
nor U13270 (N_13270,N_9056,N_11334);
or U13271 (N_13271,N_8470,N_11719);
or U13272 (N_13272,N_11975,N_9379);
nor U13273 (N_13273,N_9877,N_7758);
nor U13274 (N_13274,N_6692,N_9519);
and U13275 (N_13275,N_11384,N_10626);
and U13276 (N_13276,N_10846,N_10399);
nor U13277 (N_13277,N_8936,N_7514);
nor U13278 (N_13278,N_11663,N_10940);
or U13279 (N_13279,N_10327,N_6371);
or U13280 (N_13280,N_10742,N_6620);
and U13281 (N_13281,N_11850,N_10616);
and U13282 (N_13282,N_8635,N_10896);
and U13283 (N_13283,N_10583,N_8250);
nor U13284 (N_13284,N_7137,N_10787);
and U13285 (N_13285,N_6682,N_6299);
nor U13286 (N_13286,N_6396,N_9255);
nand U13287 (N_13287,N_7138,N_8097);
and U13288 (N_13288,N_10437,N_10239);
and U13289 (N_13289,N_7184,N_9300);
and U13290 (N_13290,N_8070,N_8108);
xnor U13291 (N_13291,N_6831,N_9666);
nor U13292 (N_13292,N_9991,N_9956);
nand U13293 (N_13293,N_6702,N_9745);
and U13294 (N_13294,N_10361,N_6662);
nor U13295 (N_13295,N_9932,N_9114);
and U13296 (N_13296,N_8125,N_11728);
or U13297 (N_13297,N_6768,N_7486);
and U13298 (N_13298,N_9755,N_7748);
nor U13299 (N_13299,N_11308,N_7076);
and U13300 (N_13300,N_8153,N_7457);
or U13301 (N_13301,N_7118,N_11828);
and U13302 (N_13302,N_6111,N_6500);
or U13303 (N_13303,N_11703,N_10379);
nor U13304 (N_13304,N_9363,N_6122);
and U13305 (N_13305,N_9470,N_10408);
nand U13306 (N_13306,N_6561,N_9646);
nand U13307 (N_13307,N_9831,N_8785);
nor U13308 (N_13308,N_11529,N_11490);
and U13309 (N_13309,N_9127,N_8526);
or U13310 (N_13310,N_7378,N_10543);
nor U13311 (N_13311,N_9538,N_9426);
and U13312 (N_13312,N_7040,N_10484);
nor U13313 (N_13313,N_8992,N_8888);
nand U13314 (N_13314,N_8591,N_7103);
and U13315 (N_13315,N_10534,N_8779);
or U13316 (N_13316,N_11600,N_7491);
nand U13317 (N_13317,N_6760,N_9820);
nor U13318 (N_13318,N_8086,N_9933);
and U13319 (N_13319,N_11439,N_10173);
and U13320 (N_13320,N_7851,N_7166);
nand U13321 (N_13321,N_6165,N_9791);
or U13322 (N_13322,N_9317,N_8987);
and U13323 (N_13323,N_6544,N_10042);
nor U13324 (N_13324,N_7504,N_10464);
or U13325 (N_13325,N_9645,N_10242);
and U13326 (N_13326,N_9702,N_9053);
nand U13327 (N_13327,N_11370,N_7494);
and U13328 (N_13328,N_7351,N_11902);
or U13329 (N_13329,N_11000,N_9495);
and U13330 (N_13330,N_7200,N_8685);
nand U13331 (N_13331,N_10816,N_11459);
xnor U13332 (N_13332,N_10978,N_8947);
and U13333 (N_13333,N_10733,N_6608);
and U13334 (N_13334,N_7278,N_8921);
and U13335 (N_13335,N_6499,N_6753);
nand U13336 (N_13336,N_10433,N_8216);
nand U13337 (N_13337,N_11399,N_7080);
or U13338 (N_13338,N_10750,N_8751);
and U13339 (N_13339,N_9125,N_11238);
or U13340 (N_13340,N_7609,N_10597);
nor U13341 (N_13341,N_11666,N_6892);
nand U13342 (N_13342,N_7213,N_10835);
or U13343 (N_13343,N_7664,N_7968);
or U13344 (N_13344,N_10852,N_9421);
nand U13345 (N_13345,N_6301,N_11614);
nand U13346 (N_13346,N_7026,N_9788);
nor U13347 (N_13347,N_6201,N_7858);
xor U13348 (N_13348,N_7197,N_7731);
or U13349 (N_13349,N_6103,N_6387);
and U13350 (N_13350,N_10376,N_11539);
nor U13351 (N_13351,N_6739,N_7820);
xor U13352 (N_13352,N_9472,N_8166);
and U13353 (N_13353,N_7937,N_9464);
or U13354 (N_13354,N_11208,N_6146);
or U13355 (N_13355,N_8050,N_6714);
or U13356 (N_13356,N_10088,N_11856);
and U13357 (N_13357,N_6789,N_6964);
or U13358 (N_13358,N_11286,N_6733);
nand U13359 (N_13359,N_7777,N_7835);
nand U13360 (N_13360,N_11366,N_7816);
xor U13361 (N_13361,N_11339,N_9597);
nor U13362 (N_13362,N_8075,N_9733);
nor U13363 (N_13363,N_6184,N_7475);
or U13364 (N_13364,N_11855,N_7725);
nor U13365 (N_13365,N_10967,N_11752);
nand U13366 (N_13366,N_7811,N_11079);
nand U13367 (N_13367,N_6412,N_9407);
nor U13368 (N_13368,N_7688,N_8610);
nor U13369 (N_13369,N_10302,N_11288);
and U13370 (N_13370,N_10159,N_6156);
and U13371 (N_13371,N_11558,N_11650);
nand U13372 (N_13372,N_8176,N_7798);
and U13373 (N_13373,N_8757,N_11015);
xor U13374 (N_13374,N_7869,N_10909);
or U13375 (N_13375,N_6391,N_10104);
nor U13376 (N_13376,N_9617,N_9152);
or U13377 (N_13377,N_6363,N_10114);
and U13378 (N_13378,N_9253,N_9732);
nor U13379 (N_13379,N_11491,N_8881);
xnor U13380 (N_13380,N_6241,N_7153);
nor U13381 (N_13381,N_6804,N_6002);
nand U13382 (N_13382,N_8918,N_11125);
nor U13383 (N_13383,N_10108,N_8903);
nand U13384 (N_13384,N_8045,N_9961);
and U13385 (N_13385,N_8322,N_10417);
nor U13386 (N_13386,N_10551,N_10364);
xor U13387 (N_13387,N_6590,N_8235);
and U13388 (N_13388,N_9911,N_7632);
or U13389 (N_13389,N_6893,N_11243);
nor U13390 (N_13390,N_11092,N_9985);
nor U13391 (N_13391,N_6655,N_10027);
nor U13392 (N_13392,N_11075,N_7072);
or U13393 (N_13393,N_10046,N_11780);
xor U13394 (N_13394,N_11524,N_7395);
and U13395 (N_13395,N_9565,N_9328);
and U13396 (N_13396,N_9843,N_7691);
and U13397 (N_13397,N_6695,N_11359);
and U13398 (N_13398,N_9525,N_6294);
or U13399 (N_13399,N_11413,N_6190);
xnor U13400 (N_13400,N_10305,N_6472);
and U13401 (N_13401,N_10202,N_10785);
nand U13402 (N_13402,N_11204,N_8808);
nand U13403 (N_13403,N_10979,N_6361);
or U13404 (N_13404,N_11604,N_6304);
and U13405 (N_13405,N_10505,N_9060);
and U13406 (N_13406,N_11383,N_11247);
and U13407 (N_13407,N_8534,N_8129);
or U13408 (N_13408,N_6389,N_8383);
and U13409 (N_13409,N_10008,N_9335);
nor U13410 (N_13410,N_6325,N_10502);
nor U13411 (N_13411,N_10023,N_8597);
and U13412 (N_13412,N_8589,N_6552);
nor U13413 (N_13413,N_8205,N_10557);
nand U13414 (N_13414,N_6548,N_9022);
and U13415 (N_13415,N_7334,N_10368);
and U13416 (N_13416,N_11700,N_11293);
or U13417 (N_13417,N_7456,N_6941);
nor U13418 (N_13418,N_7171,N_11597);
or U13419 (N_13419,N_8887,N_7155);
and U13420 (N_13420,N_6609,N_9803);
and U13421 (N_13421,N_10756,N_11632);
or U13422 (N_13422,N_9982,N_8366);
nor U13423 (N_13423,N_10797,N_6515);
xnor U13424 (N_13424,N_9456,N_11669);
nor U13425 (N_13425,N_9965,N_11898);
nor U13426 (N_13426,N_10184,N_10065);
and U13427 (N_13427,N_9132,N_11986);
xnor U13428 (N_13428,N_7757,N_11186);
nor U13429 (N_13429,N_8060,N_11161);
nor U13430 (N_13430,N_10044,N_9785);
nor U13431 (N_13431,N_7679,N_11765);
nor U13432 (N_13432,N_9874,N_9717);
nor U13433 (N_13433,N_6326,N_6586);
or U13434 (N_13434,N_10753,N_9659);
nand U13435 (N_13435,N_7191,N_11751);
or U13436 (N_13436,N_10625,N_9855);
and U13437 (N_13437,N_8450,N_7368);
nor U13438 (N_13438,N_10265,N_7945);
nor U13439 (N_13439,N_11406,N_11219);
nand U13440 (N_13440,N_8716,N_6367);
or U13441 (N_13441,N_7367,N_11516);
xnor U13442 (N_13442,N_7859,N_8092);
and U13443 (N_13443,N_6969,N_6947);
or U13444 (N_13444,N_7481,N_11162);
and U13445 (N_13445,N_6037,N_6666);
nand U13446 (N_13446,N_10351,N_9973);
and U13447 (N_13447,N_11877,N_8902);
and U13448 (N_13448,N_8232,N_10237);
nand U13449 (N_13449,N_9833,N_6936);
and U13450 (N_13450,N_9107,N_8123);
or U13451 (N_13451,N_6868,N_7850);
and U13452 (N_13452,N_7478,N_8805);
and U13453 (N_13453,N_11606,N_9889);
and U13454 (N_13454,N_10041,N_9413);
or U13455 (N_13455,N_9567,N_8233);
nor U13456 (N_13456,N_8532,N_8051);
or U13457 (N_13457,N_9714,N_10942);
and U13458 (N_13458,N_9485,N_7568);
nand U13459 (N_13459,N_8527,N_11583);
nor U13460 (N_13460,N_7501,N_7970);
and U13461 (N_13461,N_7556,N_8976);
or U13462 (N_13462,N_6265,N_9550);
xnor U13463 (N_13463,N_10539,N_9610);
nand U13464 (N_13464,N_7854,N_9178);
xor U13465 (N_13465,N_10839,N_9936);
or U13466 (N_13466,N_10736,N_6197);
and U13467 (N_13467,N_10489,N_8871);
nand U13468 (N_13468,N_7635,N_10639);
xnor U13469 (N_13469,N_6550,N_10503);
nor U13470 (N_13470,N_8531,N_7832);
nand U13471 (N_13471,N_8643,N_11656);
nand U13472 (N_13472,N_6506,N_9813);
and U13473 (N_13473,N_6076,N_7944);
nor U13474 (N_13474,N_10821,N_9794);
and U13475 (N_13475,N_11047,N_9120);
or U13476 (N_13476,N_11541,N_6476);
or U13477 (N_13477,N_6319,N_10849);
nor U13478 (N_13478,N_7329,N_9183);
xor U13479 (N_13479,N_9822,N_8169);
or U13480 (N_13480,N_7902,N_10247);
or U13481 (N_13481,N_11039,N_8671);
and U13482 (N_13482,N_7012,N_8523);
nand U13483 (N_13483,N_6459,N_10461);
and U13484 (N_13484,N_8076,N_7298);
nor U13485 (N_13485,N_8770,N_10566);
xor U13486 (N_13486,N_6104,N_9378);
nand U13487 (N_13487,N_8101,N_7160);
and U13488 (N_13488,N_10759,N_8492);
nand U13489 (N_13489,N_8032,N_10402);
and U13490 (N_13490,N_10274,N_8688);
and U13491 (N_13491,N_11503,N_6642);
and U13492 (N_13492,N_7889,N_8133);
xor U13493 (N_13493,N_8061,N_10169);
and U13494 (N_13494,N_8673,N_10654);
nor U13495 (N_13495,N_8983,N_8427);
and U13496 (N_13496,N_9530,N_6432);
or U13497 (N_13497,N_10981,N_7142);
and U13498 (N_13498,N_9739,N_8676);
and U13499 (N_13499,N_8332,N_7405);
nand U13500 (N_13500,N_10998,N_6770);
xnor U13501 (N_13501,N_10060,N_7194);
nor U13502 (N_13502,N_11012,N_10155);
nand U13503 (N_13503,N_6478,N_6238);
or U13504 (N_13504,N_6449,N_8855);
or U13505 (N_13505,N_8442,N_6773);
nor U13506 (N_13506,N_9689,N_8896);
and U13507 (N_13507,N_10775,N_7602);
and U13508 (N_13508,N_8668,N_6986);
xor U13509 (N_13509,N_8776,N_9321);
nor U13510 (N_13510,N_8862,N_9939);
nor U13511 (N_13511,N_8010,N_9930);
and U13512 (N_13512,N_8054,N_10907);
or U13513 (N_13513,N_11126,N_6345);
or U13514 (N_13514,N_11382,N_8938);
or U13515 (N_13515,N_10927,N_7470);
nand U13516 (N_13516,N_8068,N_8122);
nand U13517 (N_13517,N_8917,N_11692);
or U13518 (N_13518,N_8429,N_6840);
and U13519 (N_13519,N_7426,N_10427);
xnor U13520 (N_13520,N_9480,N_7210);
or U13521 (N_13521,N_8812,N_10227);
or U13522 (N_13522,N_11375,N_9427);
nor U13523 (N_13523,N_11023,N_6206);
or U13524 (N_13524,N_8349,N_9013);
xor U13525 (N_13525,N_9952,N_9072);
nor U13526 (N_13526,N_11422,N_10241);
or U13527 (N_13527,N_9760,N_6531);
or U13528 (N_13528,N_11820,N_7258);
or U13529 (N_13529,N_10197,N_10618);
or U13530 (N_13530,N_9507,N_11480);
and U13531 (N_13531,N_7472,N_7615);
nand U13532 (N_13532,N_11016,N_6912);
and U13533 (N_13533,N_8163,N_9169);
nand U13534 (N_13534,N_6523,N_9867);
or U13535 (N_13535,N_10784,N_9987);
or U13536 (N_13536,N_9891,N_11882);
and U13537 (N_13537,N_9737,N_7961);
xnor U13538 (N_13538,N_7737,N_7879);
nand U13539 (N_13539,N_9903,N_8801);
or U13540 (N_13540,N_11179,N_8191);
or U13541 (N_13541,N_10200,N_11559);
or U13542 (N_13542,N_6059,N_9924);
xor U13543 (N_13543,N_6237,N_11419);
nand U13544 (N_13544,N_10036,N_11116);
nor U13545 (N_13545,N_8280,N_11237);
and U13546 (N_13546,N_8126,N_7313);
nand U13547 (N_13547,N_7041,N_6060);
and U13548 (N_13548,N_11787,N_11119);
nand U13549 (N_13549,N_6564,N_7640);
or U13550 (N_13550,N_8179,N_9181);
xor U13551 (N_13551,N_10118,N_11319);
nor U13552 (N_13552,N_8269,N_6649);
nand U13553 (N_13553,N_7581,N_7993);
and U13554 (N_13554,N_10078,N_7135);
nand U13555 (N_13555,N_8120,N_10885);
and U13556 (N_13556,N_8124,N_8608);
nor U13557 (N_13557,N_10319,N_6626);
and U13558 (N_13558,N_8895,N_8617);
nor U13559 (N_13559,N_7053,N_11321);
nand U13560 (N_13560,N_6819,N_7151);
nand U13561 (N_13561,N_7924,N_6464);
or U13562 (N_13562,N_8928,N_10936);
and U13563 (N_13563,N_7004,N_6741);
and U13564 (N_13564,N_8724,N_10279);
nor U13565 (N_13565,N_7599,N_11508);
or U13566 (N_13566,N_10223,N_10167);
or U13567 (N_13567,N_7950,N_8258);
and U13568 (N_13568,N_9115,N_11774);
nor U13569 (N_13569,N_7035,N_11010);
or U13570 (N_13570,N_8288,N_11253);
or U13571 (N_13571,N_7619,N_6098);
nor U13572 (N_13572,N_10045,N_8522);
and U13573 (N_13573,N_10026,N_6900);
nor U13574 (N_13574,N_9160,N_8880);
or U13575 (N_13575,N_8465,N_7890);
and U13576 (N_13576,N_10870,N_6833);
nor U13577 (N_13577,N_6074,N_9144);
and U13578 (N_13578,N_8817,N_11510);
and U13579 (N_13579,N_8244,N_10341);
or U13580 (N_13580,N_7152,N_10015);
and U13581 (N_13581,N_9243,N_10611);
nand U13582 (N_13582,N_6737,N_9633);
nor U13583 (N_13583,N_7285,N_9620);
nor U13584 (N_13584,N_6625,N_7094);
or U13585 (N_13585,N_10491,N_7948);
and U13586 (N_13586,N_11363,N_8007);
nand U13587 (N_13587,N_7479,N_8558);
or U13588 (N_13588,N_9346,N_11511);
nor U13589 (N_13589,N_9004,N_6710);
nand U13590 (N_13590,N_10058,N_10926);
nand U13591 (N_13591,N_9641,N_9990);
or U13592 (N_13592,N_8586,N_8645);
and U13593 (N_13593,N_6119,N_11651);
and U13594 (N_13594,N_11357,N_6247);
xor U13595 (N_13595,N_8661,N_8221);
and U13596 (N_13596,N_6708,N_11612);
and U13597 (N_13597,N_6783,N_10690);
nand U13598 (N_13598,N_10670,N_10619);
nand U13599 (N_13599,N_10450,N_11596);
or U13600 (N_13600,N_9634,N_6527);
nor U13601 (N_13601,N_6554,N_7237);
nor U13602 (N_13602,N_8949,N_10047);
nand U13603 (N_13603,N_10067,N_6600);
and U13604 (N_13604,N_6511,N_11543);
nand U13605 (N_13605,N_11493,N_6896);
and U13606 (N_13606,N_8623,N_10987);
nand U13607 (N_13607,N_10115,N_11155);
nand U13608 (N_13608,N_6047,N_9104);
nor U13609 (N_13609,N_10228,N_9825);
nand U13610 (N_13610,N_9202,N_7314);
or U13611 (N_13611,N_11927,N_10050);
and U13612 (N_13612,N_9179,N_8614);
nor U13613 (N_13613,N_7304,N_10738);
and U13614 (N_13614,N_10559,N_10588);
or U13615 (N_13615,N_7918,N_9083);
nor U13616 (N_13616,N_10253,N_6853);
nand U13617 (N_13617,N_11556,N_9573);
nor U13618 (N_13618,N_10313,N_8476);
and U13619 (N_13619,N_8094,N_10868);
nor U13620 (N_13620,N_11297,N_6303);
xnor U13621 (N_13621,N_10198,N_9354);
and U13622 (N_13622,N_9438,N_11695);
or U13623 (N_13623,N_8701,N_10963);
nand U13624 (N_13624,N_9017,N_10949);
nand U13625 (N_13625,N_9657,N_7529);
nand U13626 (N_13626,N_6514,N_9161);
nor U13627 (N_13627,N_10836,N_10322);
or U13628 (N_13628,N_6805,N_7487);
and U13629 (N_13629,N_10447,N_8440);
xnor U13630 (N_13630,N_6296,N_11755);
nand U13631 (N_13631,N_10043,N_6243);
and U13632 (N_13632,N_9778,N_6274);
nand U13633 (N_13633,N_6798,N_10506);
xor U13634 (N_13634,N_9859,N_7133);
nand U13635 (N_13635,N_6654,N_8722);
and U13636 (N_13636,N_8874,N_11101);
xor U13637 (N_13637,N_7940,N_7295);
xnor U13638 (N_13638,N_11120,N_8275);
or U13639 (N_13639,N_8005,N_10707);
nor U13640 (N_13640,N_7126,N_10828);
or U13641 (N_13641,N_9055,N_11955);
nand U13642 (N_13642,N_8831,N_8786);
nand U13643 (N_13643,N_7376,N_7375);
nor U13644 (N_13644,N_6025,N_7331);
nand U13645 (N_13645,N_6332,N_11141);
nand U13646 (N_13646,N_9272,N_11402);
and U13647 (N_13647,N_6594,N_11203);
or U13648 (N_13648,N_11414,N_7018);
nand U13649 (N_13649,N_8630,N_10608);
and U13650 (N_13650,N_9628,N_11369);
nor U13651 (N_13651,N_10493,N_7995);
and U13652 (N_13652,N_9795,N_8826);
and U13653 (N_13653,N_10048,N_7657);
or U13654 (N_13654,N_10190,N_11252);
nand U13655 (N_13655,N_8725,N_11078);
nor U13656 (N_13656,N_7893,N_7730);
or U13657 (N_13657,N_9050,N_11311);
nand U13658 (N_13658,N_6762,N_8982);
nor U13659 (N_13659,N_11922,N_8819);
nand U13660 (N_13660,N_9437,N_10766);
and U13661 (N_13661,N_8787,N_8720);
and U13662 (N_13662,N_10152,N_10813);
nor U13663 (N_13663,N_7362,N_8181);
nor U13664 (N_13664,N_9479,N_7119);
or U13665 (N_13665,N_6443,N_6897);
nand U13666 (N_13666,N_8445,N_8198);
or U13667 (N_13667,N_9762,N_6734);
nand U13668 (N_13668,N_9895,N_8954);
nor U13669 (N_13669,N_10834,N_6157);
xnor U13670 (N_13670,N_7022,N_8650);
and U13671 (N_13671,N_7753,N_7826);
nand U13672 (N_13672,N_8174,N_9392);
and U13673 (N_13673,N_6175,N_7952);
nor U13674 (N_13674,N_7207,N_10224);
nand U13675 (N_13675,N_10628,N_6378);
or U13676 (N_13676,N_9111,N_11009);
and U13677 (N_13677,N_10232,N_10011);
nand U13678 (N_13678,N_6108,N_10544);
and U13679 (N_13679,N_6200,N_6440);
nand U13680 (N_13680,N_7381,N_8358);
and U13681 (N_13681,N_10443,N_7830);
nor U13682 (N_13682,N_9681,N_10829);
or U13683 (N_13683,N_7377,N_10550);
nor U13684 (N_13684,N_8372,N_10378);
and U13685 (N_13685,N_11570,N_10209);
or U13686 (N_13686,N_8170,N_11910);
nand U13687 (N_13687,N_11428,N_9884);
or U13688 (N_13688,N_7522,N_11408);
and U13689 (N_13689,N_11350,N_11679);
and U13690 (N_13690,N_9449,N_11329);
nand U13691 (N_13691,N_8845,N_10780);
or U13692 (N_13692,N_7154,N_9467);
nor U13693 (N_13693,N_6465,N_11859);
and U13694 (N_13694,N_11988,N_11822);
nor U13695 (N_13695,N_8395,N_8416);
or U13696 (N_13696,N_9223,N_11456);
nand U13697 (N_13697,N_9129,N_6315);
xor U13698 (N_13698,N_6722,N_6884);
nor U13699 (N_13699,N_10208,N_6648);
nand U13700 (N_13700,N_7795,N_7573);
and U13701 (N_13701,N_11744,N_9333);
and U13702 (N_13702,N_9727,N_8631);
nand U13703 (N_13703,N_9603,N_8452);
or U13704 (N_13704,N_6155,N_7533);
xor U13705 (N_13705,N_6482,N_8843);
or U13706 (N_13706,N_8341,N_7536);
nor U13707 (N_13707,N_10684,N_9337);
nand U13708 (N_13708,N_6901,N_7462);
nand U13709 (N_13709,N_10441,N_6584);
or U13710 (N_13710,N_9866,N_10056);
nand U13711 (N_13711,N_9857,N_9502);
or U13712 (N_13712,N_8064,N_11332);
nand U13713 (N_13713,N_6450,N_7344);
nor U13714 (N_13714,N_10532,N_8387);
xor U13715 (N_13715,N_7355,N_6803);
nor U13716 (N_13716,N_10575,N_6979);
and U13717 (N_13717,N_8925,N_9572);
nor U13718 (N_13718,N_10941,N_11317);
nand U13719 (N_13719,N_11693,N_6160);
or U13720 (N_13720,N_11890,N_11778);
nand U13721 (N_13721,N_9722,N_6975);
and U13722 (N_13722,N_11373,N_10370);
or U13723 (N_13723,N_9465,N_10333);
nor U13724 (N_13724,N_10219,N_10695);
and U13725 (N_13725,N_8362,N_7385);
and U13726 (N_13726,N_11951,N_9397);
nand U13727 (N_13727,N_6366,N_7369);
nor U13728 (N_13728,N_6126,N_11117);
nand U13729 (N_13729,N_6172,N_9306);
nor U13730 (N_13730,N_9593,N_7686);
and U13731 (N_13731,N_6350,N_10158);
nor U13732 (N_13732,N_7031,N_9026);
xor U13733 (N_13733,N_10069,N_7872);
and U13734 (N_13734,N_9963,N_10867);
or U13735 (N_13735,N_9782,N_7265);
xor U13736 (N_13736,N_11648,N_6923);
or U13737 (N_13737,N_7964,N_8272);
nor U13738 (N_13738,N_7925,N_9200);
and U13739 (N_13739,N_6435,N_9983);
and U13740 (N_13740,N_8245,N_6407);
nor U13741 (N_13741,N_7812,N_8049);
or U13742 (N_13742,N_9244,N_8882);
nand U13743 (N_13743,N_8794,N_9209);
nor U13744 (N_13744,N_11865,N_6593);
and U13745 (N_13745,N_10180,N_9925);
nand U13746 (N_13746,N_8749,N_8281);
or U13747 (N_13747,N_11769,N_11626);
and U13748 (N_13748,N_6604,N_8731);
and U13749 (N_13749,N_6117,N_9275);
or U13750 (N_13750,N_9978,N_8109);
or U13751 (N_13751,N_9155,N_8295);
nor U13752 (N_13752,N_11854,N_11163);
xor U13753 (N_13753,N_8386,N_9957);
nand U13754 (N_13754,N_6176,N_7853);
nand U13755 (N_13755,N_9398,N_8289);
and U13756 (N_13756,N_6235,N_9405);
and U13757 (N_13757,N_7306,N_11876);
and U13758 (N_13758,N_10589,N_8473);
and U13759 (N_13759,N_6974,N_10791);
and U13760 (N_13760,N_11553,N_10962);
and U13761 (N_13761,N_8365,N_11377);
nor U13762 (N_13762,N_8479,N_11166);
or U13763 (N_13763,N_6348,N_9325);
and U13764 (N_13764,N_6646,N_8161);
nand U13765 (N_13765,N_8940,N_6262);
nor U13766 (N_13766,N_11518,N_11059);
nand U13767 (N_13767,N_10106,N_10915);
nor U13768 (N_13768,N_6003,N_7287);
nand U13769 (N_13769,N_6689,N_11108);
or U13770 (N_13770,N_6454,N_7588);
nand U13771 (N_13771,N_7759,N_11637);
and U13772 (N_13772,N_7524,N_10698);
nor U13773 (N_13773,N_10359,N_10168);
nand U13774 (N_13774,N_10565,N_8920);
and U13775 (N_13775,N_7716,N_10135);
xor U13776 (N_13776,N_11216,N_9897);
nor U13777 (N_13777,N_10634,N_7796);
and U13778 (N_13778,N_10838,N_7580);
nand U13779 (N_13779,N_9079,N_11263);
and U13780 (N_13780,N_7643,N_7263);
nand U13781 (N_13781,N_10486,N_8662);
nor U13782 (N_13782,N_7273,N_10984);
nand U13783 (N_13783,N_9133,N_7509);
or U13784 (N_13784,N_7098,N_9503);
nand U13785 (N_13785,N_8926,N_9865);
xnor U13786 (N_13786,N_6023,N_7667);
and U13787 (N_13787,N_8590,N_11911);
nor U13788 (N_13788,N_6276,N_9341);
or U13789 (N_13789,N_9561,N_6829);
or U13790 (N_13790,N_9736,N_10312);
xor U13791 (N_13791,N_8025,N_8994);
nand U13792 (N_13792,N_9297,N_8828);
or U13793 (N_13793,N_8969,N_8389);
nor U13794 (N_13794,N_9883,N_7557);
nor U13795 (N_13795,N_6742,N_8607);
nor U13796 (N_13796,N_10523,N_11754);
nand U13797 (N_13797,N_7976,N_7361);
and U13798 (N_13798,N_6984,N_6528);
nand U13799 (N_13799,N_9433,N_9725);
and U13800 (N_13800,N_10425,N_8364);
nor U13801 (N_13801,N_8811,N_9001);
nand U13802 (N_13802,N_7569,N_7797);
xor U13803 (N_13803,N_11064,N_11969);
nand U13804 (N_13804,N_10864,N_10662);
nand U13805 (N_13805,N_10779,N_7480);
nor U13806 (N_13806,N_11817,N_6466);
nor U13807 (N_13807,N_6032,N_9648);
nand U13808 (N_13808,N_9639,N_11682);
nor U13809 (N_13809,N_6228,N_11051);
or U13810 (N_13810,N_7799,N_10812);
nand U13811 (N_13811,N_9361,N_9431);
and U13812 (N_13812,N_11788,N_6105);
nand U13813 (N_13813,N_7374,N_11398);
nor U13814 (N_13814,N_7186,N_8813);
and U13815 (N_13815,N_11435,N_8799);
nor U13816 (N_13816,N_8766,N_10737);
and U13817 (N_13817,N_6505,N_9560);
xor U13818 (N_13818,N_6191,N_9558);
and U13819 (N_13819,N_11217,N_9457);
or U13820 (N_13820,N_8529,N_9682);
or U13821 (N_13821,N_7177,N_11211);
or U13822 (N_13822,N_10004,N_9237);
or U13823 (N_13823,N_11792,N_10696);
or U13824 (N_13824,N_9082,N_9064);
or U13825 (N_13825,N_10504,N_10937);
nor U13826 (N_13826,N_6772,N_6623);
nand U13827 (N_13827,N_8929,N_7571);
and U13828 (N_13828,N_10444,N_6028);
nor U13829 (N_13829,N_6441,N_11022);
and U13830 (N_13830,N_7061,N_8566);
and U13831 (N_13831,N_9524,N_10487);
and U13832 (N_13832,N_9863,N_8839);
or U13833 (N_13833,N_7994,N_8852);
or U13834 (N_13834,N_11285,N_6192);
or U13835 (N_13835,N_8287,N_7653);
or U13836 (N_13836,N_9767,N_8658);
xnor U13837 (N_13837,N_11781,N_8930);
and U13838 (N_13838,N_7916,N_8414);
xnor U13839 (N_13839,N_6026,N_8834);
nor U13840 (N_13840,N_8873,N_7681);
nor U13841 (N_13841,N_6637,N_11565);
or U13842 (N_13842,N_9239,N_10769);
or U13843 (N_13843,N_8159,N_7631);
nor U13844 (N_13844,N_7363,N_10528);
or U13845 (N_13845,N_10961,N_10432);
nor U13846 (N_13846,N_9744,N_9377);
nor U13847 (N_13847,N_8999,N_6418);
nor U13848 (N_13848,N_11251,N_9282);
nand U13849 (N_13849,N_7634,N_11668);
nand U13850 (N_13850,N_11718,N_6683);
and U13851 (N_13851,N_8510,N_11137);
nor U13852 (N_13852,N_9834,N_10201);
nor U13853 (N_13853,N_10809,N_10195);
or U13854 (N_13854,N_9998,N_11568);
nand U13855 (N_13855,N_6406,N_8239);
nor U13856 (N_13856,N_9217,N_6784);
nor U13857 (N_13857,N_6000,N_8084);
xnor U13858 (N_13858,N_6645,N_10712);
nor U13859 (N_13859,N_11935,N_6536);
or U13860 (N_13860,N_6258,N_11738);
or U13861 (N_13861,N_9477,N_9436);
and U13862 (N_13862,N_10366,N_7178);
xor U13863 (N_13863,N_7765,N_6222);
and U13864 (N_13864,N_10411,N_11395);
or U13865 (N_13865,N_6672,N_8575);
nand U13866 (N_13866,N_6910,N_6272);
nor U13867 (N_13867,N_11464,N_8621);
or U13868 (N_13868,N_8213,N_11736);
nor U13869 (N_13869,N_8750,N_10617);
nand U13870 (N_13870,N_11807,N_10578);
nor U13871 (N_13871,N_9947,N_10005);
nor U13872 (N_13872,N_11300,N_11768);
and U13873 (N_13873,N_9068,N_11312);
nand U13874 (N_13874,N_7323,N_6761);
nand U13875 (N_13875,N_10675,N_7159);
nand U13876 (N_13876,N_7346,N_6944);
and U13877 (N_13877,N_11892,N_9931);
or U13878 (N_13878,N_6574,N_9087);
and U13879 (N_13879,N_10878,N_9509);
nand U13880 (N_13880,N_11734,N_11622);
and U13881 (N_13881,N_9905,N_7768);
and U13882 (N_13882,N_7146,N_10562);
and U13883 (N_13883,N_10192,N_6295);
nand U13884 (N_13884,N_8636,N_6966);
nand U13885 (N_13885,N_10405,N_7787);
or U13886 (N_13886,N_7662,N_9678);
nor U13887 (N_13887,N_8648,N_6467);
nand U13888 (N_13888,N_10946,N_10552);
or U13889 (N_13889,N_7689,N_8210);
nor U13890 (N_13890,N_11641,N_10746);
or U13891 (N_13891,N_11829,N_9532);
xor U13892 (N_13892,N_10210,N_8217);
nand U13893 (N_13893,N_9566,N_10213);
or U13894 (N_13894,N_9647,N_6850);
and U13895 (N_13895,N_11582,N_9801);
or U13896 (N_13896,N_11002,N_6533);
or U13897 (N_13897,N_7594,N_11095);
or U13898 (N_13898,N_7086,N_6497);
or U13899 (N_13899,N_7069,N_10887);
xor U13900 (N_13900,N_6430,N_10858);
or U13901 (N_13901,N_10877,N_6140);
or U13902 (N_13902,N_11704,N_9231);
nand U13903 (N_13903,N_10101,N_8854);
or U13904 (N_13904,N_10415,N_10622);
nor U13905 (N_13905,N_6775,N_8651);
nor U13906 (N_13906,N_10564,N_10037);
or U13907 (N_13907,N_7761,N_6597);
xor U13908 (N_13908,N_10329,N_6647);
nor U13909 (N_13909,N_6444,N_10824);
nand U13910 (N_13910,N_7453,N_10092);
xor U13911 (N_13911,N_11430,N_10229);
nor U13912 (N_13912,N_11316,N_6630);
or U13913 (N_13913,N_9040,N_6397);
xor U13914 (N_13914,N_11970,N_10324);
and U13915 (N_13915,N_10906,N_6144);
nor U13916 (N_13916,N_11105,N_9724);
or U13917 (N_13917,N_7857,N_9937);
nor U13918 (N_13918,N_10416,N_10980);
nor U13919 (N_13919,N_10682,N_8932);
nand U13920 (N_13920,N_7864,N_9875);
nor U13921 (N_13921,N_9158,N_8528);
nor U13922 (N_13922,N_11537,N_8893);
nor U13923 (N_13923,N_7523,N_6130);
xnor U13924 (N_13924,N_6589,N_10938);
and U13925 (N_13925,N_8901,N_9612);
nand U13926 (N_13926,N_10323,N_9110);
or U13927 (N_13927,N_6955,N_8197);
xnor U13928 (N_13928,N_11633,N_11634);
xnor U13929 (N_13929,N_7123,N_8415);
and U13930 (N_13930,N_8559,N_11994);
or U13931 (N_13931,N_7444,N_9517);
xor U13932 (N_13932,N_8189,N_9318);
xor U13933 (N_13933,N_10090,N_11457);
and U13934 (N_13934,N_6123,N_11793);
or U13935 (N_13935,N_10497,N_6439);
and U13936 (N_13936,N_11191,N_8674);
nand U13937 (N_13937,N_10735,N_10071);
nor U13938 (N_13938,N_8469,N_6008);
or U13939 (N_13939,N_9498,N_10659);
and U13940 (N_13940,N_8222,N_8709);
xor U13941 (N_13941,N_6640,N_7001);
nor U13942 (N_13942,N_10947,N_9496);
and U13943 (N_13943,N_8525,N_10988);
xor U13944 (N_13944,N_11226,N_11667);
xnor U13945 (N_13945,N_8026,N_9340);
xnor U13946 (N_13946,N_7957,N_10514);
nor U13947 (N_13947,N_8572,N_11801);
nor U13948 (N_13948,N_9664,N_9977);
nor U13949 (N_13949,N_9065,N_7467);
and U13950 (N_13950,N_11284,N_11555);
nor U13951 (N_13951,N_10154,N_7844);
and U13952 (N_13952,N_8488,N_6249);
nor U13953 (N_13953,N_7391,N_10613);
and U13954 (N_13954,N_7538,N_9247);
and U13955 (N_13955,N_8171,N_9493);
nand U13956 (N_13956,N_8549,N_11647);
nor U13957 (N_13957,N_8034,N_10434);
or U13958 (N_13958,N_9292,N_7885);
nand U13959 (N_13959,N_7914,N_9839);
and U13960 (N_13960,N_6978,N_7848);
nand U13961 (N_13961,N_7701,N_11291);
and U13962 (N_13962,N_8756,N_9850);
or U13963 (N_13963,N_7668,N_9180);
or U13964 (N_13964,N_8861,N_8438);
or U13965 (N_13965,N_11705,N_8145);
or U13966 (N_13966,N_11677,N_11915);
and U13967 (N_13967,N_9526,N_9826);
and U13968 (N_13968,N_6425,N_9350);
or U13969 (N_13969,N_7586,N_6492);
xnor U13970 (N_13970,N_8207,N_8666);
or U13971 (N_13971,N_7505,N_9899);
nand U13972 (N_13972,N_8878,N_10419);
nand U13973 (N_13973,N_8772,N_11620);
nor U13974 (N_13974,N_9266,N_10034);
nor U13975 (N_13975,N_9748,N_6019);
xnor U13976 (N_13976,N_6673,N_8580);
or U13977 (N_13977,N_9706,N_7068);
or U13978 (N_13978,N_11662,N_6614);
nor U13979 (N_13979,N_8110,N_6588);
and U13980 (N_13980,N_9869,N_9002);
nand U13981 (N_13981,N_9542,N_11306);
nor U13982 (N_13982,N_7121,N_11759);
nand U13983 (N_13983,N_6275,N_11884);
nor U13984 (N_13984,N_10172,N_8158);
nand U13985 (N_13985,N_8146,N_8637);
and U13986 (N_13986,N_10850,N_6696);
xnor U13987 (N_13987,N_6334,N_10567);
or U13988 (N_13988,N_6749,N_9194);
and U13989 (N_13989,N_7560,N_8283);
xnor U13990 (N_13990,N_6578,N_9665);
xnor U13991 (N_13991,N_9974,N_11333);
nand U13992 (N_13992,N_11193,N_6152);
and U13993 (N_13993,N_8147,N_9229);
nand U13994 (N_13994,N_8312,N_11151);
and U13995 (N_13995,N_8934,N_9585);
xor U13996 (N_13996,N_10643,N_7217);
and U13997 (N_13997,N_8363,N_7293);
and U13998 (N_13998,N_10235,N_10783);
xnor U13999 (N_13999,N_10216,N_9018);
nand U14000 (N_14000,N_11068,N_11102);
and U14001 (N_14001,N_8989,N_6748);
or U14002 (N_14002,N_11374,N_6031);
nor U14003 (N_14003,N_6063,N_9943);
or U14004 (N_14004,N_7660,N_6751);
or U14005 (N_14005,N_6774,N_9189);
nor U14006 (N_14006,N_10522,N_11527);
and U14007 (N_14007,N_11393,N_10326);
nand U14008 (N_14008,N_11874,N_6658);
nor U14009 (N_14009,N_11158,N_9157);
nand U14010 (N_14010,N_10952,N_8430);
nand U14011 (N_14011,N_11328,N_10693);
and U14012 (N_14012,N_11878,N_6080);
nand U14013 (N_14013,N_7047,N_10459);
nor U14014 (N_14014,N_8085,N_7510);
or U14015 (N_14015,N_9549,N_7320);
nand U14016 (N_14016,N_10267,N_10039);
or U14017 (N_14017,N_10296,N_9236);
or U14018 (N_14018,N_9288,N_6842);
or U14019 (N_14019,N_11861,N_6277);
and U14020 (N_14020,N_7300,N_10945);
nand U14021 (N_14021,N_10083,N_8091);
and U14022 (N_14022,N_8458,N_8693);
or U14023 (N_14023,N_11455,N_10199);
and U14024 (N_14024,N_9819,N_10507);
or U14025 (N_14025,N_9499,N_7030);
nor U14026 (N_14026,N_9771,N_8350);
and U14027 (N_14027,N_7088,N_10375);
nand U14028 (N_14028,N_8435,N_10342);
or U14029 (N_14029,N_10091,N_8669);
nor U14030 (N_14030,N_9988,N_11299);
and U14031 (N_14031,N_9441,N_8847);
nand U14032 (N_14032,N_9257,N_10854);
nor U14033 (N_14033,N_7636,N_7139);
xor U14034 (N_14034,N_7888,N_6889);
nand U14035 (N_14035,N_9491,N_10130);
nor U14036 (N_14036,N_6744,N_10757);
xnor U14037 (N_14037,N_7394,N_11697);
nand U14038 (N_14038,N_9781,N_9913);
nand U14039 (N_14039,N_8504,N_8096);
nor U14040 (N_14040,N_10540,N_6159);
xor U14041 (N_14041,N_11305,N_11446);
and U14042 (N_14042,N_6180,N_10788);
and U14043 (N_14043,N_11603,N_8467);
or U14044 (N_14044,N_7570,N_8359);
nand U14045 (N_14045,N_8742,N_9445);
xor U14046 (N_14046,N_8248,N_11823);
or U14047 (N_14047,N_6860,N_8255);
xor U14048 (N_14048,N_9880,N_10721);
xor U14049 (N_14049,N_9150,N_11746);
nand U14050 (N_14050,N_11139,N_9695);
or U14051 (N_14051,N_11005,N_6145);
nand U14052 (N_14052,N_6551,N_8821);
and U14053 (N_14053,N_11946,N_7433);
and U14054 (N_14054,N_6300,N_8039);
nand U14055 (N_14055,N_10176,N_11335);
nand U14056 (N_14056,N_6813,N_9773);
nor U14057 (N_14057,N_9191,N_10957);
or U14058 (N_14058,N_7339,N_11940);
nand U14059 (N_14059,N_11376,N_6006);
and U14060 (N_14060,N_11180,N_9743);
and U14061 (N_14061,N_10808,N_6686);
or U14062 (N_14062,N_9856,N_11150);
and U14063 (N_14063,N_9443,N_11003);
and U14064 (N_14064,N_7399,N_8451);
or U14065 (N_14065,N_8759,N_8846);
nand U14066 (N_14066,N_10939,N_11741);
or U14067 (N_14067,N_9544,N_6555);
nor U14068 (N_14068,N_10336,N_7829);
nor U14069 (N_14069,N_6088,N_10692);
or U14070 (N_14070,N_11834,N_8912);
or U14071 (N_14071,N_10123,N_9075);
nand U14072 (N_14072,N_7416,N_11533);
nor U14073 (N_14073,N_11673,N_11602);
xor U14074 (N_14074,N_11412,N_10765);
nand U14075 (N_14075,N_6916,N_7692);
nand U14076 (N_14076,N_9418,N_7257);
or U14077 (N_14077,N_7779,N_6082);
xor U14078 (N_14078,N_6549,N_7861);
or U14079 (N_14079,N_10496,N_6073);
nor U14080 (N_14080,N_11405,N_10049);
nor U14081 (N_14081,N_8948,N_9384);
nor U14082 (N_14082,N_7301,N_6764);
nand U14083 (N_14083,N_10307,N_7079);
nand U14084 (N_14084,N_7521,N_8374);
and U14085 (N_14085,N_9198,N_8698);
nor U14086 (N_14086,N_7172,N_11157);
nand U14087 (N_14087,N_9726,N_8069);
nand U14088 (N_14088,N_8967,N_6362);
and U14089 (N_14089,N_11112,N_9171);
nor U14090 (N_14090,N_7317,N_7483);
nand U14091 (N_14091,N_11965,N_6622);
nand U14092 (N_14092,N_6757,N_8016);
nand U14093 (N_14093,N_11654,N_10661);
nor U14094 (N_14094,N_10007,N_10871);
xnor U14095 (N_14095,N_7959,N_11450);
nand U14096 (N_14096,N_7104,N_9578);
or U14097 (N_14097,N_11176,N_9823);
and U14098 (N_14098,N_11825,N_10372);
or U14099 (N_14099,N_6846,N_6852);
and U14100 (N_14100,N_7562,N_7873);
and U14101 (N_14101,N_11346,N_7055);
nor U14102 (N_14102,N_11577,N_6164);
and U14103 (N_14103,N_10029,N_9098);
nor U14104 (N_14104,N_10170,N_6420);
and U14105 (N_14105,N_11785,N_7723);
or U14106 (N_14106,N_7477,N_8952);
and U14107 (N_14107,N_9187,N_7290);
xor U14108 (N_14108,N_6823,N_7585);
and U14109 (N_14109,N_7922,N_6888);
and U14110 (N_14110,N_7987,N_9197);
or U14111 (N_14111,N_8667,N_8784);
and U14112 (N_14112,N_9219,N_9849);
nor U14113 (N_14113,N_10266,N_10142);
nand U14114 (N_14114,N_10790,N_11678);
and U14115 (N_14115,N_8318,N_10930);
nand U14116 (N_14116,N_11852,N_10218);
or U14117 (N_14117,N_11689,N_6509);
and U14118 (N_14118,N_11984,N_9358);
nor U14119 (N_14119,N_9500,N_9688);
xor U14120 (N_14120,N_11931,N_8959);
and U14121 (N_14121,N_10480,N_6224);
nand U14122 (N_14122,N_6717,N_9605);
nand U14123 (N_14123,N_9707,N_8356);
or U14124 (N_14124,N_6337,N_7650);
xor U14125 (N_14125,N_9504,N_11810);
nor U14126 (N_14126,N_11436,N_8149);
nor U14127 (N_14127,N_10546,N_6324);
or U14128 (N_14128,N_9954,N_10720);
nand U14129 (N_14129,N_10178,N_11389);
and U14130 (N_14130,N_10760,N_6567);
or U14131 (N_14131,N_10781,N_9119);
and U14132 (N_14132,N_10362,N_7354);
nand U14133 (N_14133,N_8898,N_8613);
or U14134 (N_14134,N_7234,N_7220);
nand U14135 (N_14135,N_6879,N_10739);
nor U14136 (N_14136,N_10074,N_9797);
nand U14137 (N_14137,N_11044,N_10595);
nand U14138 (N_14138,N_11699,N_10600);
nand U14139 (N_14139,N_10768,N_6529);
or U14140 (N_14140,N_8708,N_11939);
nor U14141 (N_14141,N_8436,N_10134);
xnor U14142 (N_14142,N_7951,N_11708);
nor U14143 (N_14143,N_10590,N_9460);
and U14144 (N_14144,N_9588,N_10064);
nor U14145 (N_14145,N_11625,N_11590);
or U14146 (N_14146,N_10463,N_9109);
and U14147 (N_14147,N_8540,N_7703);
or U14148 (N_14148,N_9968,N_6701);
nand U14149 (N_14149,N_7600,N_10845);
or U14150 (N_14150,N_6195,N_6619);
or U14151 (N_14151,N_10886,N_9303);
nor U14152 (N_14152,N_6970,N_11006);
nand U14153 (N_14153,N_10688,N_11977);
nand U14154 (N_14154,N_7075,N_7415);
and U14155 (N_14155,N_6933,N_8330);
nand U14156 (N_14156,N_7694,N_8186);
or U14157 (N_14157,N_8910,N_11514);
or U14158 (N_14158,N_8208,N_10820);
or U14159 (N_14159,N_11496,N_7956);
or U14160 (N_14160,N_7436,N_7060);
and U14161 (N_14161,N_10052,N_11303);
nand U14162 (N_14162,N_8319,N_8022);
nand U14163 (N_14163,N_8577,N_7410);
xor U14164 (N_14164,N_6413,N_9758);
nand U14165 (N_14165,N_9245,N_6336);
and U14166 (N_14166,N_8829,N_7577);
xnor U14167 (N_14167,N_8193,N_6251);
nand U14168 (N_14168,N_8707,N_10283);
and U14169 (N_14169,N_9073,N_8298);
or U14170 (N_14170,N_6186,N_8134);
nor U14171 (N_14171,N_8628,N_10062);
nor U14172 (N_14172,N_10220,N_10793);
nand U14173 (N_14173,N_6937,N_10800);
or U14174 (N_14174,N_9216,N_6504);
and U14175 (N_14175,N_9228,N_8224);
nor U14176 (N_14176,N_9999,N_9975);
and U14177 (N_14177,N_11290,N_8426);
nand U14178 (N_14178,N_7073,N_6372);
and U14179 (N_14179,N_11684,N_8160);
nand U14180 (N_14180,N_10605,N_10890);
nand U14181 (N_14181,N_9235,N_10580);
or U14182 (N_14182,N_11811,N_7867);
nand U14183 (N_14183,N_6252,N_8557);
nor U14184 (N_14184,N_11004,N_6290);
nor U14185 (N_14185,N_6954,N_7392);
nand U14186 (N_14186,N_11816,N_7919);
nand U14187 (N_14187,N_10986,N_9851);
and U14188 (N_14188,N_10221,N_6631);
nand U14189 (N_14189,N_10098,N_8738);
nand U14190 (N_14190,N_8327,N_7226);
and U14191 (N_14191,N_7515,N_11983);
nor U14192 (N_14192,N_9506,N_11893);
xnor U14193 (N_14193,N_7625,N_6756);
nor U14194 (N_14194,N_11451,N_10678);
or U14195 (N_14195,N_9594,N_7980);
nor U14196 (N_14196,N_10290,N_6880);
and U14197 (N_14197,N_8135,N_9949);
and U14198 (N_14198,N_9463,N_11635);
and U14199 (N_14199,N_6993,N_7627);
xnor U14200 (N_14200,N_8019,N_6508);
or U14201 (N_14201,N_8663,N_6411);
nor U14202 (N_14202,N_8530,N_7174);
and U14203 (N_14203,N_11544,N_7189);
or U14204 (N_14204,N_10606,N_6665);
nor U14205 (N_14205,N_7642,N_7618);
nand U14206 (N_14206,N_10347,N_7690);
xor U14207 (N_14207,N_8024,N_7738);
nand U14208 (N_14208,N_7307,N_8791);
nand U14209 (N_14209,N_9402,N_9383);
xor U14210 (N_14210,N_10656,N_6919);
or U14211 (N_14211,N_10700,N_6680);
and U14212 (N_14212,N_6386,N_7693);
and U14213 (N_14213,N_8302,N_11198);
or U14214 (N_14214,N_6617,N_11706);
or U14215 (N_14215,N_9609,N_8659);
xnor U14216 (N_14216,N_9312,N_10204);
or U14217 (N_14217,N_9210,N_10013);
nor U14218 (N_14218,N_9718,N_10773);
and U14219 (N_14219,N_7519,N_7705);
nand U14220 (N_14220,N_11763,N_10125);
nand U14221 (N_14221,N_7092,N_8739);
nor U14222 (N_14222,N_11630,N_10668);
and U14223 (N_14223,N_7760,N_10277);
nand U14224 (N_14224,N_7330,N_11561);
nand U14225 (N_14225,N_6664,N_10508);
xor U14226 (N_14226,N_11519,N_11613);
nor U14227 (N_14227,N_8444,N_8418);
and U14228 (N_14228,N_9375,N_6005);
xnor U14229 (N_14229,N_6730,N_6929);
nand U14230 (N_14230,N_7711,N_7513);
or U14231 (N_14231,N_10070,N_11149);
and U14232 (N_14232,N_7469,N_8238);
and U14233 (N_14233,N_10490,N_11443);
nand U14234 (N_14234,N_6643,N_8820);
or U14235 (N_14235,N_11467,N_6171);
nor U14236 (N_14236,N_9829,N_8792);
and U14237 (N_14237,N_6399,N_11747);
or U14238 (N_14238,N_6887,N_9935);
nand U14239 (N_14239,N_8737,N_10194);
and U14240 (N_14240,N_6311,N_11615);
nand U14241 (N_14241,N_8401,N_11246);
or U14242 (N_14242,N_11917,N_8803);
nand U14243 (N_14243,N_7597,N_8023);
or U14244 (N_14244,N_6415,N_6512);
xnor U14245 (N_14245,N_7132,N_8626);
or U14246 (N_14246,N_8634,N_11713);
and U14247 (N_14247,N_11909,N_11421);
or U14248 (N_14248,N_10292,N_8797);
nor U14249 (N_14249,N_11096,N_10666);
nand U14250 (N_14250,N_6072,N_7870);
nand U14251 (N_14251,N_11694,N_7461);
or U14252 (N_14252,N_11720,N_9390);
xnor U14253 (N_14253,N_11100,N_7947);
or U14254 (N_14254,N_9086,N_11448);
nand U14255 (N_14255,N_8042,N_11601);
nand U14256 (N_14256,N_6134,N_7096);
nand U14257 (N_14257,N_11368,N_8640);
nand U14258 (N_14258,N_9163,N_10577);
nor U14259 (N_14259,N_6856,N_7042);
nand U14260 (N_14260,N_8652,N_10895);
or U14261 (N_14261,N_8653,N_9671);
or U14262 (N_14262,N_10082,N_10811);
or U14263 (N_14263,N_9044,N_6133);
nand U14264 (N_14264,N_9304,N_11607);
or U14265 (N_14265,N_11301,N_10545);
or U14266 (N_14266,N_8972,N_9166);
and U14267 (N_14267,N_7793,N_10452);
nor U14268 (N_14268,N_9775,N_7296);
or U14269 (N_14269,N_9475,N_10258);
or U14270 (N_14270,N_11453,N_11497);
nand U14271 (N_14271,N_6068,N_7454);
and U14272 (N_14272,N_7023,N_9539);
and U14273 (N_14273,N_11127,N_9622);
and U14274 (N_14274,N_10262,N_11083);
nand U14275 (N_14275,N_8494,N_7025);
or U14276 (N_14276,N_6935,N_10017);
nand U14277 (N_14277,N_9008,N_10440);
nor U14278 (N_14278,N_7032,N_11492);
and U14279 (N_14279,N_10642,N_10917);
xor U14280 (N_14280,N_9872,N_7242);
nand U14281 (N_14281,N_9359,N_9327);
nand U14282 (N_14282,N_11053,N_8560);
or U14283 (N_14283,N_11756,N_6081);
or U14284 (N_14284,N_8515,N_8518);
xor U14285 (N_14285,N_6242,N_10189);
xnor U14286 (N_14286,N_8585,N_11685);
nor U14287 (N_14287,N_7941,N_8856);
xor U14288 (N_14288,N_9320,N_11325);
xor U14289 (N_14289,N_11857,N_9080);
nor U14290 (N_14290,N_10992,N_11942);
or U14291 (N_14291,N_10777,N_11230);
xor U14292 (N_14292,N_6390,N_11174);
or U14293 (N_14293,N_8474,N_11256);
or U14294 (N_14294,N_8252,N_7356);
nand U14295 (N_14295,N_7187,N_7547);
or U14296 (N_14296,N_7489,N_10075);
nand U14297 (N_14297,N_9314,N_7781);
and U14298 (N_14298,N_9274,N_7592);
or U14299 (N_14299,N_11638,N_7767);
nand U14300 (N_14300,N_10848,N_9058);
or U14301 (N_14301,N_11674,N_11489);
nand U14302 (N_14302,N_11908,N_6958);
or U14303 (N_14303,N_10414,N_10579);
and U14304 (N_14304,N_7960,N_10795);
and U14305 (N_14305,N_9349,N_10841);
or U14306 (N_14306,N_10593,N_10859);
or U14307 (N_14307,N_10664,N_11580);
or U14308 (N_14308,N_11069,N_8142);
and U14309 (N_14309,N_11314,N_7958);
and U14310 (N_14310,N_10458,N_10953);
or U14311 (N_14311,N_8384,N_8827);
or U14312 (N_14312,N_8789,N_11444);
or U14313 (N_14313,N_11385,N_7327);
xnor U14314 (N_14314,N_9979,N_7465);
or U14315 (N_14315,N_8168,N_10291);
nor U14316 (N_14316,N_11469,N_8641);
nand U14317 (N_14317,N_8229,N_11318);
nor U14318 (N_14318,N_6902,N_10587);
nor U14319 (N_14319,N_11037,N_11796);
or U14320 (N_14320,N_7963,N_7365);
and U14321 (N_14321,N_10217,N_7819);
and U14322 (N_14322,N_10001,N_10599);
or U14323 (N_14323,N_6010,N_6268);
or U14324 (N_14324,N_9806,N_9900);
or U14325 (N_14325,N_9486,N_7926);
and U14326 (N_14326,N_9298,N_9749);
nor U14327 (N_14327,N_10633,N_8419);
nor U14328 (N_14328,N_8448,N_7020);
xor U14329 (N_14329,N_10243,N_11549);
or U14330 (N_14330,N_7204,N_6546);
or U14331 (N_14331,N_7969,N_7337);
or U14332 (N_14332,N_8333,N_7714);
or U14333 (N_14333,N_10255,N_6518);
nor U14334 (N_14334,N_7282,N_6121);
or U14335 (N_14335,N_9559,N_9564);
nand U14336 (N_14336,N_10477,N_9042);
nand U14337 (N_14337,N_11445,N_6698);
xor U14338 (N_14338,N_11358,N_9469);
and U14339 (N_14339,N_9100,N_8699);
and U14340 (N_14340,N_7603,N_8471);
or U14341 (N_14341,N_11008,N_10211);
or U14342 (N_14342,N_10881,N_11463);
and U14343 (N_14343,N_6484,N_8798);
or U14344 (N_14344,N_8977,N_9285);
or U14345 (N_14345,N_10061,N_7488);
and U14346 (N_14346,N_6280,N_9038);
and U14347 (N_14347,N_10174,N_7502);
nand U14348 (N_14348,N_7251,N_9938);
and U14349 (N_14349,N_7297,N_7974);
nor U14350 (N_14350,N_6214,N_9881);
nand U14351 (N_14351,N_10672,N_6836);
and U14352 (N_14352,N_7985,N_9709);
nand U14353 (N_14353,N_11862,N_9989);
and U14354 (N_14354,N_11221,N_9703);
or U14355 (N_14355,N_9271,N_6199);
and U14356 (N_14356,N_10912,N_10891);
or U14357 (N_14357,N_6292,N_10708);
or U14358 (N_14358,N_7740,N_11973);
or U14359 (N_14359,N_6289,N_8670);
or U14360 (N_14360,N_10435,N_7770);
nand U14361 (N_14361,N_10080,N_8144);
and U14362 (N_14362,N_7476,N_6379);
or U14363 (N_14363,N_8711,N_8840);
or U14364 (N_14364,N_7039,N_11265);
and U14365 (N_14365,N_8264,N_6187);
and U14366 (N_14366,N_6357,N_8953);
and U14367 (N_14367,N_8767,N_11858);
or U14368 (N_14368,N_8979,N_9230);
nand U14369 (N_14369,N_6095,N_8128);
or U14370 (N_14370,N_9195,N_8916);
xnor U14371 (N_14371,N_9108,N_11468);
nor U14372 (N_14372,N_7517,N_7131);
nor U14373 (N_14373,N_10905,N_6895);
nand U14374 (N_14374,N_10226,N_8588);
or U14375 (N_14375,N_10950,N_6576);
nor U14376 (N_14376,N_9738,N_7276);
nand U14377 (N_14377,N_7431,N_8089);
or U14378 (N_14378,N_10631,N_6822);
nor U14379 (N_14379,N_10303,N_6458);
nor U14380 (N_14380,N_8723,N_8041);
nand U14381 (N_14381,N_10010,N_11795);
nor U14382 (N_14382,N_7081,N_8971);
nand U14383 (N_14383,N_7863,N_9992);
nor U14384 (N_14384,N_7243,N_8271);
nand U14385 (N_14385,N_9468,N_11671);
or U14386 (N_14386,N_7419,N_7455);
nor U14387 (N_14387,N_6699,N_6382);
nand U14388 (N_14388,N_11926,N_6827);
nand U14389 (N_14389,N_7923,N_6347);
or U14390 (N_14390,N_9332,N_9416);
nand U14391 (N_14391,N_7417,N_7752);
nand U14392 (N_14392,N_9063,N_7604);
or U14393 (N_14393,N_10401,N_8351);
or U14394 (N_14394,N_11331,N_7707);
or U14395 (N_14395,N_8417,N_11309);
nand U14396 (N_14396,N_11757,N_9105);
nor U14397 (N_14397,N_8680,N_6498);
nor U14398 (N_14398,N_8541,N_9360);
xnor U14399 (N_14399,N_9283,N_6033);
or U14400 (N_14400,N_8963,N_10818);
xnor U14401 (N_14401,N_10077,N_10053);
or U14402 (N_14402,N_6996,N_10966);
nand U14403 (N_14403,N_7308,N_7750);
or U14404 (N_14404,N_6534,N_7551);
nor U14405 (N_14405,N_6882,N_8567);
nand U14406 (N_14406,N_10833,N_8300);
or U14407 (N_14407,N_8249,N_9414);
and U14408 (N_14408,N_10374,N_10831);
nand U14409 (N_14409,N_9440,N_8506);
nand U14410 (N_14410,N_6453,N_8206);
nor U14411 (N_14411,N_8695,N_10185);
nand U14412 (N_14412,N_9807,N_10072);
nand U14413 (N_14413,N_10955,N_7805);
or U14414 (N_14414,N_10801,N_9212);
and U14415 (N_14415,N_8432,N_8000);
nor U14416 (N_14416,N_7260,N_10920);
xor U14417 (N_14417,N_8388,N_11094);
nor U14418 (N_14418,N_7442,N_8622);
nand U14419 (N_14419,N_10334,N_11824);
nor U14420 (N_14420,N_6457,N_11189);
or U14421 (N_14421,N_6808,N_6142);
or U14422 (N_14422,N_11932,N_7928);
or U14423 (N_14423,N_10109,N_10681);
nand U14424 (N_14424,N_7003,N_10284);
nand U14425 (N_14425,N_10689,N_7228);
nand U14426 (N_14426,N_6188,N_11959);
nand U14427 (N_14427,N_11381,N_9138);
and U14428 (N_14428,N_7050,N_6193);
and U14429 (N_14429,N_11242,N_10535);
nor U14430 (N_14430,N_11213,N_8466);
nand U14431 (N_14431,N_7099,N_8809);
xnor U14432 (N_14432,N_7499,N_11981);
nand U14433 (N_14433,N_6526,N_11034);
and U14434 (N_14434,N_7117,N_8562);
or U14435 (N_14435,N_7616,N_8556);
or U14436 (N_14436,N_8136,N_11178);
xor U14437 (N_14437,N_6940,N_7396);
nand U14438 (N_14438,N_11985,N_8043);
xnor U14439 (N_14439,N_11494,N_6015);
and U14440 (N_14440,N_7755,N_7209);
or U14441 (N_14441,N_10603,N_6905);
and U14442 (N_14442,N_9196,N_9148);
nor U14443 (N_14443,N_8629,N_7988);
nor U14444 (N_14444,N_10149,N_9045);
or U14445 (N_14445,N_11140,N_6844);
or U14446 (N_14446,N_9356,N_9631);
nor U14447 (N_14447,N_9623,N_7058);
nor U14448 (N_14448,N_11504,N_11088);
and U14449 (N_14449,N_8462,N_9946);
nand U14450 (N_14450,N_8995,N_11164);
nor U14451 (N_14451,N_11387,N_11447);
or U14452 (N_14452,N_11776,N_6639);
or U14453 (N_14453,N_9430,N_7409);
xnor U14454 (N_14454,N_6669,N_6442);
nand U14455 (N_14455,N_7687,N_11019);
nor U14456 (N_14456,N_8619,N_8519);
or U14457 (N_14457,N_6653,N_11827);
nand U14458 (N_14458,N_9858,N_7865);
nand U14459 (N_14459,N_9043,N_7917);
xnor U14460 (N_14460,N_7056,N_11944);
and U14461 (N_14461,N_8974,N_6863);
or U14462 (N_14462,N_11048,N_6668);
or U14463 (N_14463,N_8453,N_10965);
nor U14464 (N_14464,N_8642,N_9324);
nand U14465 (N_14465,N_10390,N_6766);
nor U14466 (N_14466,N_6480,N_6716);
xnor U14467 (N_14467,N_10687,N_9153);
nor U14468 (N_14468,N_6790,N_11378);
nor U14469 (N_14469,N_7219,N_6627);
and U14470 (N_14470,N_11540,N_11224);
and U14471 (N_14471,N_11082,N_9958);
nor U14472 (N_14472,N_11218,N_11050);
and U14473 (N_14473,N_9735,N_11808);
or U14474 (N_14474,N_7742,N_10392);
and U14475 (N_14475,N_7656,N_10697);
nor U14476 (N_14476,N_7978,N_9734);
nor U14477 (N_14477,N_8278,N_10910);
xor U14478 (N_14478,N_9962,N_10404);
and U14479 (N_14479,N_9409,N_7239);
and U14480 (N_14480,N_6865,N_7341);
nand U14481 (N_14481,N_8203,N_8538);
and U14482 (N_14482,N_7553,N_6271);
xor U14483 (N_14483,N_6493,N_10571);
or U14484 (N_14484,N_10798,N_8194);
nand U14485 (N_14485,N_7227,N_9765);
or U14486 (N_14486,N_8511,N_10488);
nor U14487 (N_14487,N_8503,N_10586);
xor U14488 (N_14488,N_6633,N_9293);
nor U14489 (N_14489,N_9215,N_7181);
nor U14490 (N_14490,N_8793,N_6832);
and U14491 (N_14491,N_10068,N_10222);
nor U14492 (N_14492,N_6308,N_11536);
and U14493 (N_14493,N_8172,N_10685);
and U14494 (N_14494,N_8182,N_7303);
xnor U14495 (N_14495,N_9204,N_8382);
nor U14496 (N_14496,N_8564,N_10880);
xnor U14497 (N_14497,N_11196,N_11501);
or U14498 (N_14498,N_8584,N_10021);
or U14499 (N_14499,N_7270,N_6112);
nand U14500 (N_14500,N_10483,N_11584);
or U14501 (N_14501,N_7437,N_9652);
nor U14502 (N_14502,N_9790,N_7057);
nor U14503 (N_14503,N_10516,N_7574);
nand U14504 (N_14504,N_9740,N_7813);
nand U14505 (N_14505,N_10974,N_11143);
nor U14506 (N_14506,N_7218,N_7644);
or U14507 (N_14507,N_9370,N_9037);
xor U14508 (N_14508,N_7855,N_11482);
and U14509 (N_14509,N_6828,N_9016);
or U14510 (N_14510,N_7719,N_11658);
and U14511 (N_14511,N_11014,N_10293);
nor U14512 (N_14512,N_11169,N_8655);
xnor U14513 (N_14513,N_9543,N_11978);
nand U14514 (N_14514,N_7348,N_9090);
and U14515 (N_14515,N_11598,N_10151);
and U14516 (N_14516,N_8822,N_6137);
or U14517 (N_14517,N_7525,N_10346);
or U14518 (N_14518,N_8830,N_11206);
xnor U14519 (N_14519,N_7545,N_6086);
and U14520 (N_14520,N_11394,N_9412);
xor U14521 (N_14521,N_8437,N_9576);
and U14522 (N_14522,N_7843,N_10494);
nor U14523 (N_14523,N_11278,N_6374);
nand U14524 (N_14524,N_8027,N_10851);
nor U14525 (N_14525,N_8317,N_8308);
nor U14526 (N_14526,N_6657,N_10460);
nor U14527 (N_14527,N_9428,N_7373);
nor U14528 (N_14528,N_9577,N_8616);
and U14529 (N_14529,N_6949,N_7113);
or U14530 (N_14530,N_10761,N_11067);
or U14531 (N_14531,N_8279,N_6393);
and U14532 (N_14532,N_9162,N_7148);
or U14533 (N_14533,N_11281,N_11131);
or U14534 (N_14534,N_9864,N_8353);
nor U14535 (N_14535,N_10827,N_11424);
or U14536 (N_14536,N_7302,N_6330);
nor U14537 (N_14537,N_8891,N_6972);
nand U14538 (N_14538,N_10610,N_7929);
or U14539 (N_14539,N_6250,N_8485);
xor U14540 (N_14540,N_9824,N_9232);
nand U14541 (N_14541,N_8088,N_6652);
and U14542 (N_14542,N_8373,N_9311);
and U14543 (N_14543,N_11020,N_7565);
nand U14544 (N_14544,N_10343,N_6427);
and U14545 (N_14545,N_9294,N_7264);
or U14546 (N_14546,N_7034,N_7100);
nor U14547 (N_14547,N_9009,N_9986);
nor U14548 (N_14548,N_11302,N_6968);
nand U14549 (N_14549,N_9516,N_7935);
nand U14550 (N_14550,N_9401,N_8719);
nor U14551 (N_14551,N_9343,N_11919);
and U14552 (N_14552,N_11089,N_9270);
and U14553 (N_14553,N_11839,N_6227);
nor U14554 (N_14554,N_7613,N_9117);
and U14555 (N_14555,N_7946,N_9116);
nor U14556 (N_14556,N_8079,N_9199);
nand U14557 (N_14557,N_7089,N_11365);
or U14558 (N_14558,N_9715,N_10541);
nand U14559 (N_14559,N_10771,N_6991);
nand U14560 (N_14560,N_11181,N_9929);
and U14561 (N_14561,N_8537,N_11794);
and U14562 (N_14562,N_8066,N_7751);
or U14563 (N_14563,N_6248,N_6878);
or U14564 (N_14564,N_10248,N_11550);
and U14565 (N_14565,N_7718,N_11676);
or U14566 (N_14566,N_6461,N_8162);
nor U14567 (N_14567,N_8697,N_11790);
nand U14568 (N_14568,N_7549,N_9453);
nor U14569 (N_14569,N_10889,N_8681);
or U14570 (N_14570,N_8370,N_9581);
nor U14571 (N_14571,N_9626,N_6231);
nand U14572 (N_14572,N_11487,N_6269);
nand U14573 (N_14573,N_11526,N_7256);
nand U14574 (N_14574,N_9879,N_10500);
nor U14575 (N_14575,N_6540,N_7269);
nand U14576 (N_14576,N_9970,N_10406);
and U14577 (N_14577,N_9660,N_8618);
nor U14578 (N_14578,N_10614,N_10513);
and U14579 (N_14579,N_10412,N_10286);
nand U14580 (N_14580,N_10499,N_8320);
nor U14581 (N_14581,N_8849,N_8771);
nand U14582 (N_14582,N_10457,N_6989);
or U14583 (N_14583,N_6913,N_9902);
and U14584 (N_14584,N_9638,N_8130);
nor U14585 (N_14585,N_9400,N_8460);
xor U14586 (N_14586,N_8664,N_8236);
and U14587 (N_14587,N_7084,N_8508);
or U14588 (N_14588,N_9168,N_9896);
nor U14589 (N_14589,N_9142,N_8612);
nand U14590 (N_14590,N_6496,N_6587);
or U14591 (N_14591,N_6817,N_7606);
nor U14592 (N_14592,N_10972,N_10315);
nand U14593 (N_14593,N_6226,N_10120);
nand U14594 (N_14594,N_6405,N_6677);
nand U14595 (N_14595,N_8314,N_7458);
and U14596 (N_14596,N_10581,N_11523);
nand U14597 (N_14597,N_9521,N_7706);
and U14598 (N_14598,N_7021,N_9339);
nand U14599 (N_14599,N_7316,N_6107);
nand U14600 (N_14600,N_8810,N_6603);
or U14601 (N_14601,N_9336,N_9654);
or U14602 (N_14602,N_6408,N_11323);
nand U14603 (N_14603,N_9753,N_11403);
or U14604 (N_14604,N_11146,N_9281);
or U14605 (N_14605,N_7336,N_7780);
xor U14606 (N_14606,N_10903,N_11086);
nand U14607 (N_14607,N_11952,N_7065);
or U14608 (N_14608,N_6429,N_11479);
nand U14609 (N_14609,N_7149,N_10453);
xnor U14610 (N_14610,N_9423,N_9810);
or U14611 (N_14611,N_6601,N_6870);
or U14612 (N_14612,N_6077,N_7379);
nand U14613 (N_14613,N_7979,N_11743);
nor U14614 (N_14614,N_8745,N_11133);
nor U14615 (N_14615,N_10033,N_8290);
nand U14616 (N_14616,N_11074,N_6605);
nor U14617 (N_14617,N_8223,N_11249);
nand U14618 (N_14618,N_8864,N_7254);
nor U14619 (N_14619,N_9322,N_11071);
or U14620 (N_14620,N_7821,N_9510);
or U14621 (N_14621,N_7466,N_6064);
or U14622 (N_14622,N_10893,N_7620);
or U14623 (N_14623,N_8814,N_9094);
or U14624 (N_14624,N_6448,N_9888);
or U14625 (N_14625,N_11964,N_10164);
and U14626 (N_14626,N_11197,N_7033);
xnor U14627 (N_14627,N_11210,N_6747);
or U14628 (N_14628,N_8764,N_10150);
nor U14629 (N_14629,N_8804,N_10215);
and U14630 (N_14630,N_8933,N_11502);
or U14631 (N_14631,N_9173,N_10430);
and U14632 (N_14632,N_9711,N_10320);
or U14633 (N_14633,N_9821,N_11916);
nor U14634 (N_14634,N_8594,N_10145);
nor U14635 (N_14635,N_7646,N_9478);
and U14636 (N_14636,N_10747,N_11188);
nand U14637 (N_14637,N_8582,N_6723);
or U14638 (N_14638,N_6685,N_9227);
nor U14639 (N_14639,N_8148,N_8498);
or U14640 (N_14640,N_7886,N_11154);
and U14641 (N_14641,N_11172,N_6663);
nand U14642 (N_14642,N_8307,N_6170);
and U14643 (N_14643,N_10786,N_11386);
nor U14644 (N_14644,N_6872,N_6084);
nor U14645 (N_14645,N_8344,N_9976);
nor U14646 (N_14646,N_6557,N_6233);
nand U14647 (N_14647,N_8139,N_10409);
or U14648 (N_14648,N_6571,N_10884);
nand U14649 (N_14649,N_10755,N_7167);
nand U14650 (N_14650,N_6782,N_6428);
and U14651 (N_14651,N_10638,N_10741);
nor U14652 (N_14652,N_9263,N_11814);
or U14653 (N_14653,N_7876,N_9261);
and U14654 (N_14654,N_11426,N_9548);
nor U14655 (N_14655,N_7370,N_11085);
nor U14656 (N_14656,N_10251,N_6369);
and U14657 (N_14657,N_6980,N_6494);
nand U14658 (N_14658,N_7507,N_6651);
or U14659 (N_14659,N_9540,N_10694);
or U14660 (N_14660,N_6792,N_11307);
and U14661 (N_14661,N_7122,N_9035);
or U14662 (N_14662,N_8876,N_10263);
xor U14663 (N_14663,N_11267,N_11592);
and U14664 (N_14664,N_9606,N_11629);
xnor U14665 (N_14665,N_9529,N_11557);
nand U14666 (N_14666,N_6962,N_11999);
nor U14667 (N_14667,N_7347,N_11885);
nor U14668 (N_14668,N_11340,N_7014);
nand U14669 (N_14669,N_7110,N_8412);
xor U14670 (N_14670,N_9051,N_10285);
or U14671 (N_14671,N_8276,N_8190);
nor U14672 (N_14672,N_6100,N_9784);
or U14673 (N_14673,N_6961,N_7778);
or U14674 (N_14674,N_9422,N_8240);
nor U14675 (N_14675,N_7071,N_8195);
and U14676 (N_14676,N_11013,N_9505);
or U14677 (N_14677,N_7389,N_9046);
nor U14678 (N_14678,N_6001,N_6861);
nor U14679 (N_14679,N_8985,N_9316);
nand U14680 (N_14680,N_8593,N_9404);
or U14681 (N_14681,N_8273,N_11791);
nand U14682 (N_14682,N_6043,N_6582);
and U14683 (N_14683,N_7294,N_7708);
nand U14684 (N_14684,N_9568,N_6398);
and U14685 (N_14685,N_6024,N_9388);
or U14686 (N_14686,N_10892,N_11802);
and U14687 (N_14687,N_9399,N_10703);
and U14688 (N_14688,N_9406,N_8262);
or U14689 (N_14689,N_9763,N_8093);
nand U14690 (N_14690,N_8402,N_6931);
and U14691 (N_14691,N_7608,N_6020);
and U14692 (N_14692,N_10943,N_7936);
and U14693 (N_14693,N_8215,N_10328);
or U14694 (N_14694,N_11784,N_11124);
xor U14695 (N_14695,N_9067,N_8376);
nand U14696 (N_14696,N_10969,N_9411);
xor U14697 (N_14697,N_8620,N_8493);
nor U14698 (N_14698,N_10301,N_8394);
and U14699 (N_14699,N_9557,N_8297);
or U14700 (N_14700,N_9140,N_9699);
xor U14701 (N_14701,N_7261,N_8919);
nor U14702 (N_14702,N_8483,N_9752);
or U14703 (N_14703,N_11887,N_7015);
nand U14704 (N_14704,N_11961,N_10233);
nand U14705 (N_14705,N_10667,N_9033);
and U14706 (N_14706,N_7593,N_8449);
nand U14707 (N_14707,N_10369,N_11937);
or U14708 (N_14708,N_11476,N_7473);
nand U14709 (N_14709,N_6129,N_8568);
nor U14710 (N_14710,N_7093,N_6223);
nand U14711 (N_14711,N_7647,N_10604);
and U14712 (N_14712,N_10509,N_6560);
and U14713 (N_14713,N_11472,N_8422);
or U14714 (N_14714,N_10751,N_9852);
or U14715 (N_14715,N_9692,N_6318);
and U14716 (N_14716,N_6539,N_8046);
xor U14717 (N_14717,N_6510,N_11021);
and U14718 (N_14718,N_11277,N_8551);
nor U14719 (N_14719,N_6726,N_6881);
and U14720 (N_14720,N_8270,N_10119);
and U14721 (N_14721,N_8313,N_10385);
nand U14722 (N_14722,N_8114,N_8056);
nor U14723 (N_14723,N_10387,N_10620);
and U14724 (N_14724,N_6167,N_6286);
or U14725 (N_14725,N_7043,N_7762);
nand U14726 (N_14726,N_7749,N_10304);
or U14727 (N_14727,N_8113,N_9172);
nor U14728 (N_14728,N_8777,N_9904);
nand U14729 (N_14729,N_8807,N_9547);
nand U14730 (N_14730,N_6877,N_9798);
and U14731 (N_14731,N_7849,N_7248);
and U14732 (N_14732,N_7809,N_9661);
and U14733 (N_14733,N_10418,N_8424);
xor U14734 (N_14734,N_9796,N_6338);
nor U14735 (N_14735,N_9389,N_11229);
xor U14736 (N_14736,N_8058,N_11080);
nor U14737 (N_14737,N_7173,N_10479);
or U14738 (N_14738,N_8006,N_9729);
or U14739 (N_14739,N_7909,N_8017);
nor U14740 (N_14740,N_10865,N_10743);
nand U14741 (N_14741,N_8336,N_9030);
nand U14742 (N_14742,N_9683,N_7446);
nand U14743 (N_14743,N_8175,N_7309);
or U14744 (N_14744,N_7445,N_7503);
nor U14745 (N_14745,N_6759,N_9541);
nand U14746 (N_14746,N_8945,N_9556);
nand U14747 (N_14747,N_7531,N_11837);
nand U14748 (N_14748,N_7990,N_6468);
xnor U14749 (N_14749,N_11239,N_6092);
nand U14750 (N_14750,N_7776,N_6779);
or U14751 (N_14751,N_9391,N_7078);
and U14752 (N_14752,N_11875,N_11326);
and U14753 (N_14753,N_9207,N_10063);
nor U14754 (N_14754,N_6038,N_6218);
nor U14755 (N_14755,N_11061,N_7188);
nand U14756 (N_14756,N_6965,N_6755);
nor U14757 (N_14757,N_10358,N_7932);
and U14758 (N_14758,N_11809,N_9154);
nand U14759 (N_14759,N_7998,N_7678);
nand U14760 (N_14760,N_10674,N_10003);
and U14761 (N_14761,N_6360,N_9655);
nand U14762 (N_14762,N_6012,N_10568);
and U14763 (N_14763,N_6423,N_10648);
and U14764 (N_14764,N_9696,N_10894);
nand U14765 (N_14765,N_10778,N_10182);
nand U14766 (N_14766,N_11934,N_9259);
or U14767 (N_14767,N_9374,N_8434);
or U14768 (N_14768,N_7201,N_8894);
and U14769 (N_14769,N_9121,N_7554);
nor U14770 (N_14770,N_10456,N_6997);
nand U14771 (N_14771,N_7077,N_11551);
xnor U14772 (N_14772,N_9723,N_6707);
or U14773 (N_14773,N_8741,N_10651);
xnor U14774 (N_14774,N_6595,N_7274);
and U14775 (N_14775,N_8348,N_6342);
and U14776 (N_14776,N_9012,N_6826);
xnor U14777 (N_14777,N_9122,N_10310);
nor U14778 (N_14778,N_7129,N_6985);
nand U14779 (N_14779,N_9268,N_8254);
xor U14780 (N_14780,N_8765,N_7215);
nor U14781 (N_14781,N_6351,N_8354);
nand U14782 (N_14782,N_11653,N_10706);
nand U14783 (N_14783,N_6356,N_8505);
and U14784 (N_14784,N_8431,N_7724);
or U14785 (N_14785,N_7626,N_7115);
nand U14786 (N_14786,N_11228,N_9420);
or U14787 (N_14787,N_10758,N_8740);
nor U14788 (N_14788,N_8296,N_10853);
nor U14789 (N_14789,N_9694,N_7111);
nand U14790 (N_14790,N_7190,N_10591);
or U14791 (N_14791,N_6291,N_10386);
and U14792 (N_14792,N_11175,N_11427);
and U14793 (N_14793,N_7831,N_6563);
xnor U14794 (N_14794,N_7090,N_6743);
nand U14795 (N_14795,N_6083,N_11262);
nand U14796 (N_14796,N_6194,N_11115);
or U14797 (N_14797,N_11672,N_11709);
or U14798 (N_14798,N_10136,N_10956);
nand U14799 (N_14799,N_7595,N_10183);
xnor U14800 (N_14800,N_7443,N_7164);
nor U14801 (N_14801,N_7414,N_10975);
xor U14802 (N_14802,N_9934,N_11129);
xnor U14803 (N_14803,N_9777,N_6953);
nand U14804 (N_14804,N_10924,N_11320);
nor U14805 (N_14805,N_11432,N_10147);
and U14806 (N_14806,N_7105,N_11429);
or U14807 (N_14807,N_10658,N_11608);
or U14808 (N_14808,N_9248,N_8157);
or U14809 (N_14809,N_8499,N_8013);
nand U14810 (N_14810,N_8220,N_8574);
and U14811 (N_14811,N_6674,N_7249);
nand U14812 (N_14812,N_7645,N_7883);
nor U14813 (N_14813,N_10977,N_8500);
and U14814 (N_14814,N_10254,N_9258);
and U14815 (N_14815,N_8774,N_10100);
or U14816 (N_14816,N_10289,N_9221);
and U14817 (N_14817,N_8328,N_7179);
and U14818 (N_14818,N_8199,N_6720);
nand U14819 (N_14819,N_7245,N_11058);
nor U14820 (N_14820,N_10607,N_7899);
and U14821 (N_14821,N_9264,N_7192);
nand U14822 (N_14822,N_11507,N_11274);
and U14823 (N_14823,N_6845,N_7326);
nor U14824 (N_14824,N_7548,N_7697);
nor U14825 (N_14825,N_6596,N_10609);
nand U14826 (N_14826,N_11976,N_8690);
nor U14827 (N_14827,N_8062,N_6182);
nor U14828 (N_14828,N_9601,N_10923);
and U14829 (N_14829,N_9944,N_10475);
nor U14830 (N_14830,N_6436,N_11879);
nand U14831 (N_14831,N_11404,N_11276);
and U14832 (N_14832,N_6873,N_11753);
nand U14833 (N_14833,N_9481,N_6066);
or U14834 (N_14834,N_11138,N_6168);
nor U14835 (N_14835,N_9471,N_6329);
or U14836 (N_14836,N_10022,N_9669);
nor U14837 (N_14837,N_10971,N_11869);
nor U14838 (N_14838,N_10919,N_7907);
or U14839 (N_14839,N_9273,N_10918);
nor U14840 (N_14840,N_11296,N_7496);
nand U14841 (N_14841,N_6704,N_7954);
nand U14842 (N_14842,N_9286,N_7741);
nor U14843 (N_14843,N_6811,N_7495);
and U14844 (N_14844,N_7841,N_10518);
xnor U14845 (N_14845,N_6090,N_7407);
nor U14846 (N_14846,N_10076,N_7471);
nand U14847 (N_14847,N_10057,N_11343);
nand U14848 (N_14848,N_11548,N_8923);
or U14849 (N_14849,N_9721,N_9537);
nand U14850 (N_14850,N_10873,N_6383);
or U14851 (N_14851,N_8886,N_6776);
or U14852 (N_14852,N_6971,N_8524);
and U14853 (N_14853,N_9432,N_11109);
xnor U14854 (N_14854,N_10652,N_8514);
nand U14855 (N_14855,N_10844,N_6690);
nor U14856 (N_14856,N_10713,N_6487);
nor U14857 (N_14857,N_7350,N_11077);
nand U14858 (N_14858,N_10451,N_6377);
or U14859 (N_14859,N_11033,N_8520);
nor U14860 (N_14860,N_11943,N_7027);
nand U14861 (N_14861,N_6675,N_6306);
or U14862 (N_14862,N_7518,N_9673);
nand U14863 (N_14863,N_7240,N_11588);
nand U14864 (N_14864,N_6322,N_10570);
nor U14865 (N_14865,N_8463,N_10206);
nand U14866 (N_14866,N_11991,N_6380);
xor U14867 (N_14867,N_9005,N_10073);
or U14868 (N_14868,N_8717,N_6661);
and U14869 (N_14869,N_7241,N_6344);
nor U14870 (N_14870,N_10810,N_10308);
nand U14871 (N_14871,N_9380,N_8857);
xnor U14872 (N_14872,N_8914,N_8713);
or U14873 (N_14873,N_10099,N_8321);
xor U14874 (N_14874,N_10261,N_8835);
nor U14875 (N_14875,N_11851,N_10734);
nand U14876 (N_14876,N_11111,N_6928);
or U14877 (N_14877,N_6547,N_8265);
or U14878 (N_14878,N_7814,N_9995);
nand U14879 (N_14879,N_10055,N_6503);
nand U14880 (N_14880,N_11581,N_10862);
or U14881 (N_14881,N_8294,N_9015);
nor U14882 (N_14882,N_11886,N_9996);
nand U14883 (N_14883,N_10276,N_11992);
and U14884 (N_14884,N_7745,N_9802);
nor U14885 (N_14885,N_6009,N_9459);
nor U14886 (N_14886,N_7801,N_8185);
nor U14887 (N_14887,N_7371,N_6542);
nor U14888 (N_14888,N_6911,N_10928);
and U14889 (N_14889,N_8214,N_10331);
or U14890 (N_14890,N_8274,N_7097);
and U14891 (N_14891,N_6942,N_10140);
xnor U14892 (N_14892,N_9062,N_11798);
xor U14893 (N_14893,N_11933,N_10257);
nor U14894 (N_14894,N_11831,N_11571);
nand U14895 (N_14895,N_11275,N_8957);
nand U14896 (N_14896,N_8292,N_7017);
or U14897 (N_14897,N_11202,N_7143);
nor U14898 (N_14898,N_10615,N_10117);
xor U14899 (N_14899,N_11815,N_8615);
and U14900 (N_14900,N_10472,N_7991);
nor U14901 (N_14901,N_11327,N_10127);
nand U14902 (N_14902,N_9757,N_8866);
or U14903 (N_14903,N_9357,N_10754);
and U14904 (N_14904,N_11156,N_9608);
nor U14905 (N_14905,N_6136,N_11621);
or U14906 (N_14906,N_8030,N_7666);
xor U14907 (N_14907,N_10767,N_6946);
nor U14908 (N_14908,N_6061,N_6525);
nand U14909 (N_14909,N_6051,N_11938);
nand U14910 (N_14910,N_7838,N_8512);
nand U14911 (N_14911,N_9627,N_11454);
or U14912 (N_14912,N_7390,N_7382);
nor U14913 (N_14913,N_11351,N_10009);
nor U14914 (N_14914,N_7397,N_9010);
nor U14915 (N_14915,N_11572,N_6585);
or U14916 (N_14916,N_8915,N_11657);
nor U14917 (N_14917,N_7195,N_9039);
or U14918 (N_14918,N_9146,N_11097);
xnor U14919 (N_14919,N_11270,N_6455);
nand U14920 (N_14920,N_8413,N_11711);
nor U14921 (N_14921,N_8095,N_11843);
nor U14922 (N_14922,N_6727,N_8844);
nand U14923 (N_14923,N_7413,N_11042);
and U14924 (N_14924,N_11356,N_9130);
or U14925 (N_14925,N_6460,N_6771);
nor U14926 (N_14926,N_8164,N_7791);
or U14927 (N_14927,N_6196,N_8346);
xnor U14928 (N_14928,N_9474,N_7224);
and U14929 (N_14929,N_6862,N_6065);
or U14930 (N_14930,N_9220,N_9697);
xnor U14931 (N_14931,N_9023,N_6705);
nor U14932 (N_14932,N_9041,N_11257);
or U14933 (N_14933,N_11846,N_8259);
nand U14934 (N_14934,N_7628,N_10511);
or U14935 (N_14935,N_11731,N_9676);
nand U14936 (N_14936,N_6209,N_7312);
nand U14937 (N_14937,N_11586,N_9287);
nor U14938 (N_14938,N_11056,N_7283);
nor U14939 (N_14939,N_6264,N_7544);
nand U14940 (N_14940,N_11032,N_6778);
nand U14941 (N_14941,N_6096,N_6198);
nor U14942 (N_14942,N_9591,N_11438);
and U14943 (N_14943,N_10555,N_10598);
and U14944 (N_14944,N_6401,N_7193);
or U14945 (N_14945,N_9710,N_8065);
or U14946 (N_14946,N_8997,N_11696);
xnor U14947 (N_14947,N_6437,N_9885);
and U14948 (N_14948,N_10181,N_11113);
nor U14949 (N_14949,N_9667,N_8569);
xor U14950 (N_14950,N_8165,N_9476);
nand U14951 (N_14951,N_6052,N_6781);
or U14952 (N_14952,N_8775,N_11742);
xnor U14953 (N_14953,N_8806,N_7785);
nand U14954 (N_14954,N_11011,N_6212);
nor U14955 (N_14955,N_6410,N_11409);
nor U14956 (N_14956,N_11918,N_10770);
nand U14957 (N_14957,N_6162,N_11826);
or U14958 (N_14958,N_10676,N_6424);
or U14959 (N_14959,N_11028,N_9921);
nor U14960 (N_14960,N_6316,N_6147);
nand U14961 (N_14961,N_8021,N_10295);
nor U14962 (N_14962,N_7158,N_6927);
and U14963 (N_14963,N_8546,N_10855);
or U14964 (N_14964,N_9953,N_11967);
nand U14965 (N_14965,N_8752,N_9249);
xor U14966 (N_14966,N_7054,N_9269);
xor U14967 (N_14967,N_10126,N_11282);
nand U14968 (N_14968,N_11750,N_10018);
and U14969 (N_14969,N_10352,N_9596);
or U14970 (N_14970,N_11348,N_10922);
nor U14971 (N_14971,N_9089,N_7965);
nor U14972 (N_14972,N_7680,N_10632);
or U14973 (N_14973,N_7558,N_9847);
nor U14974 (N_14974,N_6676,N_6050);
nor U14975 (N_14975,N_9092,N_11341);
and U14976 (N_14976,N_10875,N_10141);
or U14977 (N_14977,N_7659,N_7262);
or U14978 (N_14978,N_9754,N_8956);
or U14979 (N_14979,N_11081,N_9185);
or U14980 (N_14980,N_6520,N_11515);
nor U14981 (N_14981,N_7535,N_8654);
nand U14982 (N_14982,N_9768,N_7546);
nand U14983 (N_14983,N_9598,N_10572);
and U14984 (N_14984,N_9366,N_8393);
and U14985 (N_14985,N_10394,N_6939);
nand U14986 (N_14986,N_8335,N_9649);
nor U14987 (N_14987,N_7955,N_11860);
and U14988 (N_14988,N_6323,N_6352);
or U14989 (N_14989,N_9085,N_7822);
and U14990 (N_14990,N_6952,N_8347);
and U14991 (N_14991,N_9164,N_6203);
nor U14992 (N_14992,N_9277,N_6612);
nor U14993 (N_14993,N_8509,N_6867);
nand U14994 (N_14994,N_6376,N_7729);
nand U14995 (N_14995,N_11845,N_7325);
and U14996 (N_14996,N_11760,N_6519);
nand U14997 (N_14997,N_8595,N_11103);
nand U14998 (N_14998,N_6281,N_11863);
nand U14999 (N_14999,N_9586,N_11683);
nor U15000 (N_15000,N_10812,N_7951);
or U15001 (N_15001,N_6420,N_8014);
nand U15002 (N_15002,N_6851,N_6553);
nand U15003 (N_15003,N_11252,N_6437);
nand U15004 (N_15004,N_11230,N_9975);
nor U15005 (N_15005,N_11851,N_11452);
nand U15006 (N_15006,N_10614,N_9671);
nand U15007 (N_15007,N_7138,N_6246);
nor U15008 (N_15008,N_8740,N_6116);
and U15009 (N_15009,N_7462,N_6012);
nor U15010 (N_15010,N_9166,N_10187);
and U15011 (N_15011,N_11429,N_9463);
or U15012 (N_15012,N_9100,N_10943);
nor U15013 (N_15013,N_11143,N_7074);
nor U15014 (N_15014,N_9368,N_9059);
nor U15015 (N_15015,N_7848,N_6820);
and U15016 (N_15016,N_10766,N_6584);
nand U15017 (N_15017,N_8095,N_8391);
xnor U15018 (N_15018,N_9226,N_7358);
and U15019 (N_15019,N_10488,N_6078);
nor U15020 (N_15020,N_11652,N_11293);
or U15021 (N_15021,N_10291,N_6276);
nor U15022 (N_15022,N_9059,N_9353);
and U15023 (N_15023,N_9615,N_9287);
nor U15024 (N_15024,N_10144,N_10607);
nor U15025 (N_15025,N_10195,N_11965);
nor U15026 (N_15026,N_10030,N_9338);
or U15027 (N_15027,N_6846,N_8076);
xor U15028 (N_15028,N_8175,N_11372);
nor U15029 (N_15029,N_6565,N_7265);
or U15030 (N_15030,N_6481,N_8484);
nand U15031 (N_15031,N_7797,N_9745);
nand U15032 (N_15032,N_8356,N_10089);
or U15033 (N_15033,N_11190,N_11757);
or U15034 (N_15034,N_10663,N_9033);
or U15035 (N_15035,N_9099,N_8793);
and U15036 (N_15036,N_10008,N_7252);
and U15037 (N_15037,N_8180,N_10453);
or U15038 (N_15038,N_10863,N_6843);
and U15039 (N_15039,N_8571,N_8123);
xnor U15040 (N_15040,N_10538,N_11878);
nor U15041 (N_15041,N_7118,N_7632);
nor U15042 (N_15042,N_7447,N_10756);
or U15043 (N_15043,N_11607,N_11367);
or U15044 (N_15044,N_6521,N_9944);
nand U15045 (N_15045,N_7567,N_7563);
or U15046 (N_15046,N_11294,N_7605);
or U15047 (N_15047,N_9398,N_11454);
nand U15048 (N_15048,N_6243,N_9411);
and U15049 (N_15049,N_7111,N_9722);
nor U15050 (N_15050,N_10240,N_10960);
or U15051 (N_15051,N_7619,N_9230);
or U15052 (N_15052,N_8828,N_7105);
xor U15053 (N_15053,N_8567,N_9457);
nand U15054 (N_15054,N_10462,N_11759);
or U15055 (N_15055,N_11519,N_9501);
nor U15056 (N_15056,N_10275,N_9062);
and U15057 (N_15057,N_11377,N_9818);
xnor U15058 (N_15058,N_9023,N_6433);
xor U15059 (N_15059,N_9099,N_9773);
or U15060 (N_15060,N_10386,N_6829);
and U15061 (N_15061,N_7965,N_9499);
nor U15062 (N_15062,N_8254,N_9511);
or U15063 (N_15063,N_6599,N_10063);
xnor U15064 (N_15064,N_11882,N_10904);
or U15065 (N_15065,N_6430,N_11099);
nor U15066 (N_15066,N_6649,N_8497);
nand U15067 (N_15067,N_10539,N_9568);
nand U15068 (N_15068,N_11708,N_9589);
and U15069 (N_15069,N_9570,N_9291);
and U15070 (N_15070,N_10563,N_10316);
or U15071 (N_15071,N_6764,N_7208);
or U15072 (N_15072,N_9130,N_7938);
or U15073 (N_15073,N_8076,N_9379);
and U15074 (N_15074,N_7516,N_10937);
nand U15075 (N_15075,N_11472,N_6751);
xor U15076 (N_15076,N_11908,N_8767);
or U15077 (N_15077,N_9418,N_7249);
and U15078 (N_15078,N_6508,N_9410);
or U15079 (N_15079,N_10930,N_8981);
nand U15080 (N_15080,N_10058,N_7250);
nor U15081 (N_15081,N_6886,N_9453);
nor U15082 (N_15082,N_6982,N_7309);
nand U15083 (N_15083,N_6894,N_9467);
nand U15084 (N_15084,N_6838,N_9779);
nand U15085 (N_15085,N_8542,N_7443);
or U15086 (N_15086,N_10422,N_10053);
and U15087 (N_15087,N_11051,N_7087);
nor U15088 (N_15088,N_8081,N_8284);
nor U15089 (N_15089,N_6753,N_10456);
nor U15090 (N_15090,N_8491,N_11099);
or U15091 (N_15091,N_10375,N_6536);
nand U15092 (N_15092,N_11271,N_7335);
nor U15093 (N_15093,N_9601,N_8311);
nand U15094 (N_15094,N_7116,N_7802);
or U15095 (N_15095,N_7765,N_10991);
nand U15096 (N_15096,N_9549,N_9079);
nand U15097 (N_15097,N_8439,N_9922);
and U15098 (N_15098,N_11047,N_9253);
and U15099 (N_15099,N_11566,N_9484);
or U15100 (N_15100,N_6450,N_8448);
xor U15101 (N_15101,N_6737,N_7657);
or U15102 (N_15102,N_8945,N_10219);
nor U15103 (N_15103,N_11564,N_6193);
or U15104 (N_15104,N_9255,N_11249);
nand U15105 (N_15105,N_7684,N_8275);
or U15106 (N_15106,N_11256,N_7890);
or U15107 (N_15107,N_6368,N_6916);
or U15108 (N_15108,N_11049,N_7684);
nor U15109 (N_15109,N_8790,N_8846);
or U15110 (N_15110,N_9381,N_8686);
and U15111 (N_15111,N_10860,N_8485);
nor U15112 (N_15112,N_10180,N_11599);
nor U15113 (N_15113,N_10667,N_10921);
and U15114 (N_15114,N_9700,N_6327);
xnor U15115 (N_15115,N_7583,N_11010);
nor U15116 (N_15116,N_8136,N_10245);
xnor U15117 (N_15117,N_6792,N_9895);
xor U15118 (N_15118,N_6447,N_11431);
nor U15119 (N_15119,N_8332,N_6178);
and U15120 (N_15120,N_8457,N_11665);
and U15121 (N_15121,N_10003,N_8282);
nand U15122 (N_15122,N_7070,N_10035);
xor U15123 (N_15123,N_7291,N_7055);
and U15124 (N_15124,N_10221,N_8358);
and U15125 (N_15125,N_8981,N_10212);
and U15126 (N_15126,N_10878,N_7143);
and U15127 (N_15127,N_9540,N_6768);
or U15128 (N_15128,N_6338,N_6132);
or U15129 (N_15129,N_7825,N_8358);
nand U15130 (N_15130,N_6599,N_10332);
nor U15131 (N_15131,N_6912,N_7065);
nor U15132 (N_15132,N_8752,N_6489);
and U15133 (N_15133,N_7259,N_9377);
and U15134 (N_15134,N_8155,N_11009);
nand U15135 (N_15135,N_8085,N_11706);
nor U15136 (N_15136,N_9159,N_10510);
nor U15137 (N_15137,N_8999,N_7956);
or U15138 (N_15138,N_10415,N_9551);
nor U15139 (N_15139,N_7927,N_8188);
and U15140 (N_15140,N_8865,N_9904);
xor U15141 (N_15141,N_6098,N_9900);
or U15142 (N_15142,N_10381,N_7369);
nor U15143 (N_15143,N_9748,N_9292);
and U15144 (N_15144,N_9660,N_11664);
or U15145 (N_15145,N_8608,N_8937);
nor U15146 (N_15146,N_9942,N_8712);
nor U15147 (N_15147,N_6872,N_8976);
or U15148 (N_15148,N_11589,N_8593);
nand U15149 (N_15149,N_6015,N_10222);
xnor U15150 (N_15150,N_10256,N_11324);
and U15151 (N_15151,N_9189,N_11577);
nor U15152 (N_15152,N_9783,N_11809);
nand U15153 (N_15153,N_7119,N_6529);
or U15154 (N_15154,N_10345,N_9492);
and U15155 (N_15155,N_6947,N_7524);
nand U15156 (N_15156,N_10619,N_8863);
nand U15157 (N_15157,N_11071,N_6404);
nand U15158 (N_15158,N_8395,N_8430);
nor U15159 (N_15159,N_7684,N_6602);
xor U15160 (N_15160,N_6639,N_11757);
and U15161 (N_15161,N_10834,N_6232);
xnor U15162 (N_15162,N_8724,N_11331);
nand U15163 (N_15163,N_11836,N_6083);
or U15164 (N_15164,N_6968,N_11196);
or U15165 (N_15165,N_11823,N_10751);
and U15166 (N_15166,N_9330,N_8011);
nand U15167 (N_15167,N_11656,N_7017);
nor U15168 (N_15168,N_7343,N_8790);
nor U15169 (N_15169,N_11673,N_8872);
xor U15170 (N_15170,N_11716,N_9319);
nor U15171 (N_15171,N_9240,N_8408);
nand U15172 (N_15172,N_10739,N_7592);
nand U15173 (N_15173,N_8213,N_10752);
nor U15174 (N_15174,N_8995,N_6450);
nor U15175 (N_15175,N_11453,N_10487);
and U15176 (N_15176,N_11207,N_8061);
nand U15177 (N_15177,N_7270,N_7829);
and U15178 (N_15178,N_9306,N_8960);
nor U15179 (N_15179,N_8403,N_7294);
and U15180 (N_15180,N_10285,N_10609);
xnor U15181 (N_15181,N_6222,N_7987);
and U15182 (N_15182,N_9223,N_7436);
and U15183 (N_15183,N_9835,N_10530);
nor U15184 (N_15184,N_11116,N_10178);
nand U15185 (N_15185,N_8775,N_6631);
nand U15186 (N_15186,N_10676,N_11031);
nand U15187 (N_15187,N_8264,N_7052);
or U15188 (N_15188,N_10872,N_9629);
nor U15189 (N_15189,N_9941,N_9448);
nand U15190 (N_15190,N_9960,N_10876);
or U15191 (N_15191,N_8687,N_8953);
or U15192 (N_15192,N_10144,N_8957);
and U15193 (N_15193,N_8200,N_7487);
nor U15194 (N_15194,N_6445,N_10482);
or U15195 (N_15195,N_6484,N_10638);
and U15196 (N_15196,N_10098,N_11527);
or U15197 (N_15197,N_7428,N_9671);
or U15198 (N_15198,N_9861,N_10373);
or U15199 (N_15199,N_7095,N_8565);
or U15200 (N_15200,N_7300,N_8023);
or U15201 (N_15201,N_6543,N_9725);
nor U15202 (N_15202,N_9309,N_8084);
nor U15203 (N_15203,N_7584,N_10052);
nand U15204 (N_15204,N_8408,N_8625);
or U15205 (N_15205,N_8107,N_6062);
or U15206 (N_15206,N_10235,N_11617);
xnor U15207 (N_15207,N_8574,N_6599);
nor U15208 (N_15208,N_10169,N_8871);
nand U15209 (N_15209,N_10086,N_9439);
xnor U15210 (N_15210,N_9800,N_6919);
and U15211 (N_15211,N_9314,N_10165);
and U15212 (N_15212,N_6947,N_8325);
and U15213 (N_15213,N_8435,N_8287);
nand U15214 (N_15214,N_9633,N_6390);
xor U15215 (N_15215,N_10311,N_6896);
nand U15216 (N_15216,N_8138,N_8309);
nand U15217 (N_15217,N_11062,N_8996);
nand U15218 (N_15218,N_8671,N_8634);
xnor U15219 (N_15219,N_9948,N_8518);
nand U15220 (N_15220,N_11986,N_8176);
or U15221 (N_15221,N_6009,N_7289);
xnor U15222 (N_15222,N_6772,N_8007);
nand U15223 (N_15223,N_11793,N_7124);
nor U15224 (N_15224,N_11111,N_10553);
and U15225 (N_15225,N_6611,N_11682);
nor U15226 (N_15226,N_7713,N_6074);
or U15227 (N_15227,N_8131,N_7545);
or U15228 (N_15228,N_10558,N_10807);
xor U15229 (N_15229,N_9325,N_6556);
nand U15230 (N_15230,N_9948,N_11980);
and U15231 (N_15231,N_10522,N_10826);
nor U15232 (N_15232,N_6580,N_10761);
xor U15233 (N_15233,N_6770,N_11886);
or U15234 (N_15234,N_8005,N_6957);
nand U15235 (N_15235,N_6139,N_9666);
or U15236 (N_15236,N_7556,N_7850);
nand U15237 (N_15237,N_6268,N_8354);
xor U15238 (N_15238,N_9180,N_10855);
nor U15239 (N_15239,N_9558,N_9743);
nor U15240 (N_15240,N_10958,N_8709);
and U15241 (N_15241,N_10792,N_7933);
and U15242 (N_15242,N_10681,N_10641);
or U15243 (N_15243,N_6502,N_6624);
or U15244 (N_15244,N_7553,N_11298);
nor U15245 (N_15245,N_10185,N_7961);
nor U15246 (N_15246,N_7624,N_11087);
nor U15247 (N_15247,N_8812,N_7282);
nand U15248 (N_15248,N_6838,N_10909);
or U15249 (N_15249,N_9134,N_8809);
nor U15250 (N_15250,N_11375,N_8020);
nand U15251 (N_15251,N_11325,N_7984);
xor U15252 (N_15252,N_6870,N_9394);
or U15253 (N_15253,N_8534,N_10650);
xor U15254 (N_15254,N_9087,N_11896);
nor U15255 (N_15255,N_7016,N_11801);
xnor U15256 (N_15256,N_6748,N_7424);
nor U15257 (N_15257,N_6832,N_9986);
nand U15258 (N_15258,N_8631,N_8359);
or U15259 (N_15259,N_6974,N_10611);
or U15260 (N_15260,N_6997,N_9442);
and U15261 (N_15261,N_8526,N_7670);
and U15262 (N_15262,N_10250,N_9106);
and U15263 (N_15263,N_7237,N_9537);
and U15264 (N_15264,N_10095,N_7527);
nand U15265 (N_15265,N_9305,N_6495);
or U15266 (N_15266,N_9174,N_7625);
nand U15267 (N_15267,N_8946,N_10965);
or U15268 (N_15268,N_8326,N_11760);
nand U15269 (N_15269,N_7918,N_7998);
xor U15270 (N_15270,N_9771,N_9118);
or U15271 (N_15271,N_10551,N_11324);
and U15272 (N_15272,N_9750,N_9807);
nand U15273 (N_15273,N_8841,N_8087);
and U15274 (N_15274,N_11386,N_8270);
xor U15275 (N_15275,N_7731,N_11865);
xor U15276 (N_15276,N_6293,N_6614);
or U15277 (N_15277,N_6706,N_8280);
nor U15278 (N_15278,N_6122,N_9806);
and U15279 (N_15279,N_7517,N_6975);
nand U15280 (N_15280,N_10170,N_8024);
or U15281 (N_15281,N_6685,N_7507);
and U15282 (N_15282,N_8382,N_7770);
and U15283 (N_15283,N_9528,N_9634);
and U15284 (N_15284,N_9889,N_6138);
nand U15285 (N_15285,N_6942,N_7269);
and U15286 (N_15286,N_9311,N_6792);
nor U15287 (N_15287,N_9303,N_9404);
nand U15288 (N_15288,N_10349,N_7381);
or U15289 (N_15289,N_10491,N_8362);
xor U15290 (N_15290,N_10203,N_7215);
or U15291 (N_15291,N_10679,N_6922);
and U15292 (N_15292,N_7850,N_6783);
nor U15293 (N_15293,N_11349,N_10471);
nor U15294 (N_15294,N_10756,N_11424);
and U15295 (N_15295,N_8377,N_9170);
xor U15296 (N_15296,N_11390,N_7629);
nand U15297 (N_15297,N_11103,N_7394);
and U15298 (N_15298,N_9412,N_9768);
xnor U15299 (N_15299,N_7266,N_11154);
nand U15300 (N_15300,N_8727,N_6223);
or U15301 (N_15301,N_6904,N_7935);
nor U15302 (N_15302,N_6523,N_8047);
and U15303 (N_15303,N_6425,N_11220);
and U15304 (N_15304,N_7452,N_8876);
and U15305 (N_15305,N_6537,N_7387);
nor U15306 (N_15306,N_6527,N_7569);
and U15307 (N_15307,N_8512,N_8931);
nand U15308 (N_15308,N_8053,N_7399);
or U15309 (N_15309,N_9594,N_7226);
nand U15310 (N_15310,N_7791,N_7985);
or U15311 (N_15311,N_7590,N_9947);
and U15312 (N_15312,N_9312,N_8537);
or U15313 (N_15313,N_9167,N_11448);
nand U15314 (N_15314,N_9933,N_8187);
nor U15315 (N_15315,N_6271,N_8243);
or U15316 (N_15316,N_8447,N_7936);
nor U15317 (N_15317,N_9700,N_7904);
nor U15318 (N_15318,N_7027,N_11714);
or U15319 (N_15319,N_8780,N_11420);
nor U15320 (N_15320,N_9168,N_9805);
nand U15321 (N_15321,N_8360,N_6327);
or U15322 (N_15322,N_9649,N_6203);
or U15323 (N_15323,N_6765,N_8905);
xnor U15324 (N_15324,N_7279,N_6893);
xnor U15325 (N_15325,N_10888,N_6383);
or U15326 (N_15326,N_7306,N_10588);
and U15327 (N_15327,N_9540,N_7029);
or U15328 (N_15328,N_7853,N_9607);
or U15329 (N_15329,N_11279,N_8516);
nand U15330 (N_15330,N_8279,N_10545);
xor U15331 (N_15331,N_11394,N_10110);
nor U15332 (N_15332,N_6214,N_9956);
and U15333 (N_15333,N_11527,N_8560);
and U15334 (N_15334,N_9294,N_9512);
and U15335 (N_15335,N_6251,N_11460);
and U15336 (N_15336,N_9020,N_6816);
nand U15337 (N_15337,N_7694,N_9323);
or U15338 (N_15338,N_9894,N_7348);
nand U15339 (N_15339,N_8104,N_9404);
nor U15340 (N_15340,N_10256,N_10586);
or U15341 (N_15341,N_9351,N_11083);
nor U15342 (N_15342,N_6108,N_10853);
or U15343 (N_15343,N_6790,N_6086);
or U15344 (N_15344,N_8265,N_9322);
or U15345 (N_15345,N_9701,N_10483);
nor U15346 (N_15346,N_8093,N_10825);
nor U15347 (N_15347,N_8202,N_11221);
or U15348 (N_15348,N_8803,N_8723);
and U15349 (N_15349,N_6241,N_8036);
or U15350 (N_15350,N_7363,N_11453);
and U15351 (N_15351,N_6802,N_8989);
or U15352 (N_15352,N_11687,N_6419);
and U15353 (N_15353,N_11211,N_9706);
and U15354 (N_15354,N_10914,N_6045);
nor U15355 (N_15355,N_9704,N_11945);
xor U15356 (N_15356,N_10525,N_7477);
nand U15357 (N_15357,N_8868,N_6118);
nor U15358 (N_15358,N_10231,N_10385);
or U15359 (N_15359,N_11574,N_6567);
nand U15360 (N_15360,N_7037,N_11024);
or U15361 (N_15361,N_11078,N_9168);
nor U15362 (N_15362,N_10203,N_7534);
nor U15363 (N_15363,N_7043,N_8288);
nor U15364 (N_15364,N_7797,N_9943);
or U15365 (N_15365,N_10254,N_9979);
or U15366 (N_15366,N_7124,N_9406);
and U15367 (N_15367,N_11868,N_6202);
xnor U15368 (N_15368,N_10509,N_9394);
nand U15369 (N_15369,N_6909,N_10639);
or U15370 (N_15370,N_8171,N_7689);
nand U15371 (N_15371,N_9107,N_11673);
nor U15372 (N_15372,N_10820,N_6354);
and U15373 (N_15373,N_8823,N_7498);
nor U15374 (N_15374,N_10422,N_6844);
nand U15375 (N_15375,N_11859,N_7839);
nand U15376 (N_15376,N_9524,N_8933);
xor U15377 (N_15377,N_11261,N_10269);
or U15378 (N_15378,N_11502,N_11889);
and U15379 (N_15379,N_9239,N_9744);
or U15380 (N_15380,N_6494,N_6162);
nand U15381 (N_15381,N_8780,N_6041);
nor U15382 (N_15382,N_8601,N_9445);
and U15383 (N_15383,N_10991,N_7827);
or U15384 (N_15384,N_11651,N_10522);
nor U15385 (N_15385,N_11772,N_7176);
xor U15386 (N_15386,N_11627,N_10593);
and U15387 (N_15387,N_6698,N_11419);
and U15388 (N_15388,N_9276,N_8212);
and U15389 (N_15389,N_10384,N_11508);
and U15390 (N_15390,N_9542,N_8142);
nor U15391 (N_15391,N_9076,N_9071);
nand U15392 (N_15392,N_8979,N_9188);
nand U15393 (N_15393,N_8119,N_8697);
nand U15394 (N_15394,N_6222,N_7721);
and U15395 (N_15395,N_7714,N_11788);
nand U15396 (N_15396,N_11247,N_10714);
xor U15397 (N_15397,N_9558,N_9745);
nor U15398 (N_15398,N_7873,N_9071);
and U15399 (N_15399,N_11762,N_10531);
nand U15400 (N_15400,N_11509,N_7442);
xnor U15401 (N_15401,N_8401,N_10525);
and U15402 (N_15402,N_7061,N_6055);
xor U15403 (N_15403,N_11137,N_10596);
and U15404 (N_15404,N_11134,N_7682);
and U15405 (N_15405,N_7458,N_6244);
nand U15406 (N_15406,N_7713,N_11750);
xnor U15407 (N_15407,N_9058,N_6511);
nor U15408 (N_15408,N_10805,N_7359);
and U15409 (N_15409,N_8635,N_11820);
nand U15410 (N_15410,N_11344,N_11583);
nand U15411 (N_15411,N_10427,N_7592);
and U15412 (N_15412,N_9999,N_6654);
nor U15413 (N_15413,N_7507,N_11860);
xor U15414 (N_15414,N_6501,N_7887);
nand U15415 (N_15415,N_11272,N_8381);
and U15416 (N_15416,N_6383,N_10437);
xor U15417 (N_15417,N_7247,N_11282);
nor U15418 (N_15418,N_7112,N_10562);
and U15419 (N_15419,N_7044,N_6625);
nand U15420 (N_15420,N_7761,N_9662);
nand U15421 (N_15421,N_8543,N_7453);
and U15422 (N_15422,N_6462,N_9804);
nor U15423 (N_15423,N_6023,N_7263);
and U15424 (N_15424,N_10304,N_10846);
or U15425 (N_15425,N_10476,N_10249);
and U15426 (N_15426,N_8155,N_10413);
or U15427 (N_15427,N_10608,N_8206);
and U15428 (N_15428,N_7880,N_9547);
or U15429 (N_15429,N_10133,N_9953);
nor U15430 (N_15430,N_6070,N_10630);
nor U15431 (N_15431,N_10376,N_7991);
or U15432 (N_15432,N_9468,N_8008);
and U15433 (N_15433,N_9497,N_9219);
xor U15434 (N_15434,N_9567,N_6608);
or U15435 (N_15435,N_11003,N_7271);
or U15436 (N_15436,N_6009,N_9491);
and U15437 (N_15437,N_8255,N_6266);
xor U15438 (N_15438,N_10001,N_11118);
nand U15439 (N_15439,N_6362,N_7259);
nand U15440 (N_15440,N_11317,N_8623);
nand U15441 (N_15441,N_10922,N_7420);
nor U15442 (N_15442,N_7983,N_11570);
nor U15443 (N_15443,N_10336,N_11937);
and U15444 (N_15444,N_11335,N_8799);
nor U15445 (N_15445,N_8783,N_7236);
nor U15446 (N_15446,N_11322,N_11262);
nand U15447 (N_15447,N_10617,N_10922);
xnor U15448 (N_15448,N_6481,N_6013);
nor U15449 (N_15449,N_6077,N_8488);
nor U15450 (N_15450,N_11027,N_8290);
and U15451 (N_15451,N_11808,N_11933);
or U15452 (N_15452,N_6118,N_9196);
nand U15453 (N_15453,N_9380,N_6369);
nand U15454 (N_15454,N_9930,N_6176);
or U15455 (N_15455,N_10264,N_7766);
nand U15456 (N_15456,N_10610,N_9608);
nor U15457 (N_15457,N_7155,N_11860);
and U15458 (N_15458,N_7862,N_7008);
nand U15459 (N_15459,N_6057,N_9906);
or U15460 (N_15460,N_7635,N_7844);
and U15461 (N_15461,N_7016,N_7949);
nor U15462 (N_15462,N_8654,N_6695);
and U15463 (N_15463,N_6613,N_9306);
and U15464 (N_15464,N_7803,N_8798);
or U15465 (N_15465,N_8118,N_8683);
or U15466 (N_15466,N_8434,N_6981);
nand U15467 (N_15467,N_10107,N_7349);
and U15468 (N_15468,N_6739,N_8835);
and U15469 (N_15469,N_7663,N_8792);
and U15470 (N_15470,N_7579,N_11854);
nor U15471 (N_15471,N_8192,N_11618);
or U15472 (N_15472,N_8011,N_10515);
or U15473 (N_15473,N_7405,N_8486);
or U15474 (N_15474,N_8532,N_10018);
nand U15475 (N_15475,N_10979,N_6531);
or U15476 (N_15476,N_11168,N_8114);
nor U15477 (N_15477,N_8792,N_11097);
nand U15478 (N_15478,N_7349,N_10215);
nor U15479 (N_15479,N_9696,N_10879);
nand U15480 (N_15480,N_9515,N_7907);
and U15481 (N_15481,N_9556,N_10043);
nand U15482 (N_15482,N_6625,N_6048);
xnor U15483 (N_15483,N_9333,N_11552);
or U15484 (N_15484,N_11054,N_9561);
xor U15485 (N_15485,N_10959,N_6609);
nand U15486 (N_15486,N_8462,N_10313);
and U15487 (N_15487,N_10890,N_7255);
nand U15488 (N_15488,N_7134,N_11207);
and U15489 (N_15489,N_11763,N_9056);
and U15490 (N_15490,N_11992,N_7328);
xnor U15491 (N_15491,N_9741,N_7080);
nand U15492 (N_15492,N_7082,N_7612);
xor U15493 (N_15493,N_9594,N_7279);
nand U15494 (N_15494,N_11762,N_6331);
nand U15495 (N_15495,N_11679,N_11395);
nor U15496 (N_15496,N_10659,N_7324);
and U15497 (N_15497,N_8554,N_7128);
nor U15498 (N_15498,N_7688,N_9959);
xor U15499 (N_15499,N_9065,N_9089);
nand U15500 (N_15500,N_6072,N_11323);
nand U15501 (N_15501,N_6648,N_6007);
or U15502 (N_15502,N_8500,N_10265);
xor U15503 (N_15503,N_10564,N_10889);
and U15504 (N_15504,N_11432,N_8205);
nor U15505 (N_15505,N_6525,N_10353);
nand U15506 (N_15506,N_11191,N_9557);
and U15507 (N_15507,N_11170,N_10583);
and U15508 (N_15508,N_6644,N_6559);
nand U15509 (N_15509,N_7627,N_9772);
and U15510 (N_15510,N_6395,N_6289);
or U15511 (N_15511,N_10784,N_7103);
xnor U15512 (N_15512,N_9591,N_7395);
or U15513 (N_15513,N_8494,N_11000);
or U15514 (N_15514,N_9055,N_7093);
xnor U15515 (N_15515,N_9268,N_11606);
and U15516 (N_15516,N_11358,N_11429);
nor U15517 (N_15517,N_8294,N_9388);
nor U15518 (N_15518,N_6535,N_6733);
nand U15519 (N_15519,N_8436,N_11912);
nand U15520 (N_15520,N_9894,N_8667);
and U15521 (N_15521,N_6192,N_8199);
nor U15522 (N_15522,N_6521,N_11419);
nand U15523 (N_15523,N_7793,N_7787);
or U15524 (N_15524,N_9131,N_8766);
nor U15525 (N_15525,N_8900,N_6758);
or U15526 (N_15526,N_7423,N_10588);
or U15527 (N_15527,N_10503,N_6557);
nor U15528 (N_15528,N_11638,N_8083);
nand U15529 (N_15529,N_9663,N_10094);
and U15530 (N_15530,N_8782,N_7390);
xor U15531 (N_15531,N_6378,N_11593);
and U15532 (N_15532,N_10106,N_9751);
or U15533 (N_15533,N_8303,N_9756);
nand U15534 (N_15534,N_6476,N_9182);
nand U15535 (N_15535,N_6085,N_7847);
xor U15536 (N_15536,N_9395,N_7826);
xor U15537 (N_15537,N_6482,N_7659);
nand U15538 (N_15538,N_7660,N_11928);
or U15539 (N_15539,N_6173,N_9609);
nand U15540 (N_15540,N_9750,N_8964);
or U15541 (N_15541,N_10261,N_6291);
or U15542 (N_15542,N_9047,N_8918);
nor U15543 (N_15543,N_6343,N_11613);
and U15544 (N_15544,N_6270,N_6555);
nand U15545 (N_15545,N_6657,N_6937);
nor U15546 (N_15546,N_8172,N_11255);
xor U15547 (N_15547,N_11374,N_6782);
or U15548 (N_15548,N_7225,N_10581);
nand U15549 (N_15549,N_8914,N_10444);
nand U15550 (N_15550,N_7377,N_6316);
nor U15551 (N_15551,N_7563,N_10547);
or U15552 (N_15552,N_8484,N_7403);
nand U15553 (N_15553,N_11334,N_6460);
nand U15554 (N_15554,N_7115,N_9495);
nand U15555 (N_15555,N_8102,N_9603);
and U15556 (N_15556,N_11864,N_10216);
xnor U15557 (N_15557,N_10498,N_6100);
and U15558 (N_15558,N_10381,N_10648);
or U15559 (N_15559,N_9065,N_9387);
or U15560 (N_15560,N_6650,N_10618);
nand U15561 (N_15561,N_11496,N_6575);
and U15562 (N_15562,N_9586,N_11275);
or U15563 (N_15563,N_6933,N_10981);
nand U15564 (N_15564,N_9764,N_8814);
nand U15565 (N_15565,N_9493,N_11270);
nor U15566 (N_15566,N_10173,N_8719);
or U15567 (N_15567,N_11773,N_10181);
and U15568 (N_15568,N_6244,N_6969);
and U15569 (N_15569,N_9921,N_11614);
nor U15570 (N_15570,N_11923,N_7609);
nand U15571 (N_15571,N_7929,N_9766);
or U15572 (N_15572,N_7422,N_7406);
and U15573 (N_15573,N_7859,N_8665);
and U15574 (N_15574,N_6606,N_10466);
nand U15575 (N_15575,N_11651,N_10377);
or U15576 (N_15576,N_10575,N_7897);
and U15577 (N_15577,N_9911,N_11164);
or U15578 (N_15578,N_11858,N_9408);
and U15579 (N_15579,N_6402,N_10436);
or U15580 (N_15580,N_10237,N_10703);
nor U15581 (N_15581,N_8945,N_11130);
nand U15582 (N_15582,N_9946,N_7076);
nor U15583 (N_15583,N_11596,N_8046);
or U15584 (N_15584,N_11460,N_8838);
nor U15585 (N_15585,N_10509,N_6754);
nor U15586 (N_15586,N_10286,N_11474);
nand U15587 (N_15587,N_6188,N_6415);
or U15588 (N_15588,N_7367,N_9022);
and U15589 (N_15589,N_9936,N_11647);
nor U15590 (N_15590,N_7929,N_6897);
xnor U15591 (N_15591,N_7604,N_8736);
xor U15592 (N_15592,N_10054,N_8975);
xnor U15593 (N_15593,N_6869,N_8437);
and U15594 (N_15594,N_11355,N_7897);
xnor U15595 (N_15595,N_10114,N_8835);
or U15596 (N_15596,N_11607,N_9136);
nand U15597 (N_15597,N_8907,N_6879);
nand U15598 (N_15598,N_7984,N_9880);
nand U15599 (N_15599,N_9189,N_9990);
nor U15600 (N_15600,N_6038,N_7020);
or U15601 (N_15601,N_6669,N_6208);
nor U15602 (N_15602,N_9732,N_7367);
nand U15603 (N_15603,N_10368,N_10243);
and U15604 (N_15604,N_9276,N_9809);
nor U15605 (N_15605,N_7790,N_9377);
nor U15606 (N_15606,N_7772,N_10550);
or U15607 (N_15607,N_7575,N_7972);
nand U15608 (N_15608,N_10183,N_10955);
or U15609 (N_15609,N_6082,N_8104);
and U15610 (N_15610,N_10545,N_11714);
and U15611 (N_15611,N_11379,N_11490);
nor U15612 (N_15612,N_6976,N_7987);
xor U15613 (N_15613,N_6267,N_10552);
and U15614 (N_15614,N_9442,N_8667);
xnor U15615 (N_15615,N_7689,N_9903);
nand U15616 (N_15616,N_8837,N_9062);
and U15617 (N_15617,N_9704,N_6957);
or U15618 (N_15618,N_7500,N_8920);
nand U15619 (N_15619,N_10063,N_8341);
and U15620 (N_15620,N_7331,N_7684);
nor U15621 (N_15621,N_7190,N_7410);
nor U15622 (N_15622,N_6768,N_6432);
nor U15623 (N_15623,N_8300,N_10123);
and U15624 (N_15624,N_6778,N_11853);
or U15625 (N_15625,N_11119,N_8962);
nor U15626 (N_15626,N_11827,N_7867);
and U15627 (N_15627,N_11215,N_11740);
or U15628 (N_15628,N_7560,N_7826);
nor U15629 (N_15629,N_7768,N_9593);
nand U15630 (N_15630,N_8135,N_6755);
nor U15631 (N_15631,N_8302,N_7153);
nand U15632 (N_15632,N_7216,N_6847);
nor U15633 (N_15633,N_8653,N_10745);
or U15634 (N_15634,N_6027,N_9563);
nor U15635 (N_15635,N_11825,N_9217);
nor U15636 (N_15636,N_7716,N_8916);
and U15637 (N_15637,N_7488,N_11265);
nand U15638 (N_15638,N_8111,N_10467);
xnor U15639 (N_15639,N_8412,N_9420);
or U15640 (N_15640,N_11834,N_11975);
xor U15641 (N_15641,N_6580,N_8488);
nand U15642 (N_15642,N_8651,N_6273);
xor U15643 (N_15643,N_10726,N_8357);
or U15644 (N_15644,N_11428,N_7162);
nand U15645 (N_15645,N_10721,N_8465);
or U15646 (N_15646,N_10547,N_6743);
xnor U15647 (N_15647,N_10353,N_11255);
and U15648 (N_15648,N_6232,N_11228);
or U15649 (N_15649,N_8197,N_9548);
nor U15650 (N_15650,N_7253,N_11506);
or U15651 (N_15651,N_9756,N_9165);
or U15652 (N_15652,N_9238,N_7184);
and U15653 (N_15653,N_8896,N_7461);
nand U15654 (N_15654,N_8031,N_6499);
xor U15655 (N_15655,N_7390,N_8540);
and U15656 (N_15656,N_10238,N_11278);
or U15657 (N_15657,N_8327,N_6600);
or U15658 (N_15658,N_8522,N_10482);
nor U15659 (N_15659,N_10592,N_6562);
xnor U15660 (N_15660,N_6873,N_9713);
nor U15661 (N_15661,N_8757,N_10242);
or U15662 (N_15662,N_9193,N_6379);
xnor U15663 (N_15663,N_9685,N_8984);
nand U15664 (N_15664,N_10400,N_8756);
or U15665 (N_15665,N_7753,N_9397);
and U15666 (N_15666,N_6691,N_9529);
and U15667 (N_15667,N_10914,N_10821);
or U15668 (N_15668,N_8410,N_10185);
nor U15669 (N_15669,N_8228,N_10846);
and U15670 (N_15670,N_8575,N_10834);
and U15671 (N_15671,N_11405,N_11103);
nand U15672 (N_15672,N_9482,N_6746);
nor U15673 (N_15673,N_8234,N_6092);
and U15674 (N_15674,N_9549,N_8048);
xor U15675 (N_15675,N_11716,N_7392);
xor U15676 (N_15676,N_11439,N_9699);
nand U15677 (N_15677,N_10368,N_11060);
and U15678 (N_15678,N_10265,N_6356);
nand U15679 (N_15679,N_11166,N_9174);
or U15680 (N_15680,N_7381,N_9495);
nand U15681 (N_15681,N_7933,N_6863);
nor U15682 (N_15682,N_10085,N_9287);
nand U15683 (N_15683,N_6358,N_9580);
nor U15684 (N_15684,N_10165,N_11598);
nand U15685 (N_15685,N_7326,N_7234);
xor U15686 (N_15686,N_10936,N_7152);
nor U15687 (N_15687,N_10476,N_11399);
nor U15688 (N_15688,N_10216,N_10659);
nand U15689 (N_15689,N_7784,N_8914);
and U15690 (N_15690,N_10062,N_11442);
nand U15691 (N_15691,N_11687,N_7911);
and U15692 (N_15692,N_9012,N_10698);
nor U15693 (N_15693,N_6184,N_11691);
nor U15694 (N_15694,N_6769,N_7439);
xnor U15695 (N_15695,N_10974,N_6622);
and U15696 (N_15696,N_8960,N_11717);
and U15697 (N_15697,N_10527,N_6027);
or U15698 (N_15698,N_6068,N_8309);
and U15699 (N_15699,N_10041,N_7616);
and U15700 (N_15700,N_10350,N_9173);
nand U15701 (N_15701,N_9364,N_6777);
or U15702 (N_15702,N_9136,N_9813);
and U15703 (N_15703,N_6205,N_7248);
and U15704 (N_15704,N_8795,N_9941);
nand U15705 (N_15705,N_10670,N_9439);
or U15706 (N_15706,N_7890,N_6780);
and U15707 (N_15707,N_7036,N_8040);
nand U15708 (N_15708,N_6205,N_7444);
or U15709 (N_15709,N_6922,N_10179);
or U15710 (N_15710,N_6388,N_6767);
nand U15711 (N_15711,N_6018,N_6477);
and U15712 (N_15712,N_7440,N_6474);
nand U15713 (N_15713,N_9523,N_6372);
xor U15714 (N_15714,N_8021,N_7878);
nand U15715 (N_15715,N_7122,N_7113);
nand U15716 (N_15716,N_9707,N_6152);
and U15717 (N_15717,N_6436,N_10380);
nor U15718 (N_15718,N_10723,N_11058);
nor U15719 (N_15719,N_9064,N_8983);
or U15720 (N_15720,N_10363,N_11849);
and U15721 (N_15721,N_9672,N_9454);
and U15722 (N_15722,N_6598,N_9400);
or U15723 (N_15723,N_11407,N_6451);
and U15724 (N_15724,N_9624,N_9079);
nor U15725 (N_15725,N_9588,N_7079);
nand U15726 (N_15726,N_10420,N_8131);
nand U15727 (N_15727,N_10571,N_8670);
or U15728 (N_15728,N_6111,N_10822);
nor U15729 (N_15729,N_11605,N_10383);
or U15730 (N_15730,N_9303,N_9877);
and U15731 (N_15731,N_11743,N_9495);
nand U15732 (N_15732,N_11900,N_10569);
nor U15733 (N_15733,N_7136,N_10290);
xor U15734 (N_15734,N_10901,N_7440);
nand U15735 (N_15735,N_7679,N_10200);
or U15736 (N_15736,N_6987,N_7522);
or U15737 (N_15737,N_8035,N_8467);
and U15738 (N_15738,N_10201,N_7244);
and U15739 (N_15739,N_9252,N_10911);
or U15740 (N_15740,N_8706,N_6612);
xor U15741 (N_15741,N_8974,N_7700);
xnor U15742 (N_15742,N_6554,N_11805);
xnor U15743 (N_15743,N_8002,N_6904);
nand U15744 (N_15744,N_11655,N_11108);
and U15745 (N_15745,N_11482,N_6100);
and U15746 (N_15746,N_10990,N_6246);
and U15747 (N_15747,N_9845,N_8048);
nand U15748 (N_15748,N_10619,N_10092);
nor U15749 (N_15749,N_11777,N_7192);
or U15750 (N_15750,N_7578,N_6906);
and U15751 (N_15751,N_7520,N_7687);
and U15752 (N_15752,N_8305,N_6059);
and U15753 (N_15753,N_9819,N_6753);
xor U15754 (N_15754,N_7106,N_9298);
and U15755 (N_15755,N_11992,N_6277);
nor U15756 (N_15756,N_11970,N_8064);
nor U15757 (N_15757,N_8057,N_6339);
nand U15758 (N_15758,N_10249,N_6765);
or U15759 (N_15759,N_11535,N_6068);
nor U15760 (N_15760,N_7617,N_7150);
nor U15761 (N_15761,N_10431,N_9529);
and U15762 (N_15762,N_10549,N_9953);
and U15763 (N_15763,N_9952,N_7907);
and U15764 (N_15764,N_7988,N_7995);
and U15765 (N_15765,N_9371,N_10225);
or U15766 (N_15766,N_7086,N_6346);
xnor U15767 (N_15767,N_9242,N_7118);
nand U15768 (N_15768,N_7847,N_11230);
or U15769 (N_15769,N_9161,N_8038);
and U15770 (N_15770,N_8763,N_6888);
xnor U15771 (N_15771,N_7140,N_7156);
nand U15772 (N_15772,N_8152,N_7655);
xnor U15773 (N_15773,N_11966,N_10941);
xnor U15774 (N_15774,N_9501,N_11417);
nor U15775 (N_15775,N_8528,N_9780);
or U15776 (N_15776,N_9165,N_8198);
nand U15777 (N_15777,N_10223,N_10594);
nand U15778 (N_15778,N_11606,N_10351);
and U15779 (N_15779,N_10251,N_11246);
or U15780 (N_15780,N_6055,N_11327);
nand U15781 (N_15781,N_9727,N_9535);
and U15782 (N_15782,N_8518,N_10733);
and U15783 (N_15783,N_10919,N_8471);
nor U15784 (N_15784,N_6488,N_11926);
xnor U15785 (N_15785,N_11269,N_11033);
or U15786 (N_15786,N_10273,N_7715);
nor U15787 (N_15787,N_11959,N_7304);
or U15788 (N_15788,N_6124,N_10513);
nor U15789 (N_15789,N_11153,N_7627);
nor U15790 (N_15790,N_10573,N_6465);
and U15791 (N_15791,N_10071,N_6213);
nand U15792 (N_15792,N_7170,N_8450);
or U15793 (N_15793,N_6583,N_11237);
nor U15794 (N_15794,N_7898,N_11036);
nor U15795 (N_15795,N_7490,N_8987);
nor U15796 (N_15796,N_6473,N_6055);
nand U15797 (N_15797,N_11596,N_9175);
or U15798 (N_15798,N_10912,N_10585);
and U15799 (N_15799,N_6175,N_8275);
or U15800 (N_15800,N_7467,N_6248);
nor U15801 (N_15801,N_6984,N_10924);
xnor U15802 (N_15802,N_9612,N_10152);
and U15803 (N_15803,N_8215,N_6191);
xnor U15804 (N_15804,N_11088,N_11397);
or U15805 (N_15805,N_10991,N_9994);
xnor U15806 (N_15806,N_10786,N_10454);
nand U15807 (N_15807,N_8923,N_9503);
nor U15808 (N_15808,N_6162,N_9652);
nand U15809 (N_15809,N_10836,N_7351);
nand U15810 (N_15810,N_8009,N_11253);
nor U15811 (N_15811,N_6255,N_7889);
nor U15812 (N_15812,N_10793,N_11396);
and U15813 (N_15813,N_9635,N_8218);
and U15814 (N_15814,N_9048,N_9591);
nor U15815 (N_15815,N_9478,N_6196);
nand U15816 (N_15816,N_6232,N_10238);
xnor U15817 (N_15817,N_7510,N_11013);
and U15818 (N_15818,N_7680,N_10876);
or U15819 (N_15819,N_7586,N_8763);
and U15820 (N_15820,N_9370,N_7065);
nor U15821 (N_15821,N_7152,N_10732);
xor U15822 (N_15822,N_9084,N_8894);
nand U15823 (N_15823,N_8625,N_11620);
and U15824 (N_15824,N_7009,N_11086);
xnor U15825 (N_15825,N_7861,N_10842);
xnor U15826 (N_15826,N_10695,N_7858);
nor U15827 (N_15827,N_9052,N_11361);
nand U15828 (N_15828,N_7834,N_7647);
and U15829 (N_15829,N_7779,N_11591);
or U15830 (N_15830,N_8949,N_6270);
or U15831 (N_15831,N_7925,N_8739);
or U15832 (N_15832,N_11645,N_10321);
or U15833 (N_15833,N_7116,N_9839);
or U15834 (N_15834,N_8552,N_8494);
and U15835 (N_15835,N_7739,N_8378);
and U15836 (N_15836,N_9771,N_10493);
and U15837 (N_15837,N_10879,N_10381);
or U15838 (N_15838,N_9554,N_10240);
nand U15839 (N_15839,N_6017,N_10122);
or U15840 (N_15840,N_9864,N_11544);
nand U15841 (N_15841,N_6719,N_11697);
and U15842 (N_15842,N_11967,N_6758);
nor U15843 (N_15843,N_8597,N_8636);
nand U15844 (N_15844,N_10647,N_11924);
nand U15845 (N_15845,N_10090,N_8442);
or U15846 (N_15846,N_10227,N_7386);
nor U15847 (N_15847,N_9186,N_7222);
or U15848 (N_15848,N_8111,N_6672);
nor U15849 (N_15849,N_9063,N_9421);
nand U15850 (N_15850,N_6222,N_8096);
nor U15851 (N_15851,N_7002,N_10634);
nand U15852 (N_15852,N_11624,N_6714);
and U15853 (N_15853,N_8136,N_11416);
nor U15854 (N_15854,N_9285,N_11550);
nor U15855 (N_15855,N_6434,N_11364);
and U15856 (N_15856,N_9633,N_11684);
nand U15857 (N_15857,N_11772,N_11731);
nand U15858 (N_15858,N_9114,N_6256);
xnor U15859 (N_15859,N_9385,N_9938);
nand U15860 (N_15860,N_6913,N_10925);
and U15861 (N_15861,N_10803,N_9292);
or U15862 (N_15862,N_6702,N_10127);
nand U15863 (N_15863,N_7488,N_6594);
xnor U15864 (N_15864,N_7795,N_8190);
xnor U15865 (N_15865,N_9496,N_7394);
nor U15866 (N_15866,N_10771,N_10779);
or U15867 (N_15867,N_11628,N_11519);
or U15868 (N_15868,N_7735,N_7797);
nor U15869 (N_15869,N_6478,N_7067);
nor U15870 (N_15870,N_9618,N_7435);
xnor U15871 (N_15871,N_8019,N_11757);
or U15872 (N_15872,N_9748,N_8812);
nand U15873 (N_15873,N_9611,N_11135);
nor U15874 (N_15874,N_7216,N_6066);
and U15875 (N_15875,N_9924,N_6612);
nand U15876 (N_15876,N_9526,N_10347);
or U15877 (N_15877,N_10844,N_9876);
and U15878 (N_15878,N_10486,N_8857);
nand U15879 (N_15879,N_8599,N_9326);
or U15880 (N_15880,N_6277,N_6574);
nand U15881 (N_15881,N_11103,N_7773);
nor U15882 (N_15882,N_8622,N_11634);
nand U15883 (N_15883,N_11342,N_7642);
and U15884 (N_15884,N_9057,N_8784);
and U15885 (N_15885,N_11834,N_10067);
or U15886 (N_15886,N_8012,N_9448);
xor U15887 (N_15887,N_10892,N_10452);
nand U15888 (N_15888,N_11807,N_11539);
nand U15889 (N_15889,N_6542,N_7572);
nor U15890 (N_15890,N_11811,N_7631);
and U15891 (N_15891,N_11793,N_7474);
and U15892 (N_15892,N_8337,N_8160);
nand U15893 (N_15893,N_7984,N_10190);
and U15894 (N_15894,N_6926,N_8641);
nor U15895 (N_15895,N_10433,N_11192);
nor U15896 (N_15896,N_6432,N_7742);
nor U15897 (N_15897,N_11480,N_11442);
nand U15898 (N_15898,N_8344,N_7291);
xor U15899 (N_15899,N_10132,N_10937);
nor U15900 (N_15900,N_8530,N_9521);
nor U15901 (N_15901,N_8830,N_11158);
nand U15902 (N_15902,N_7473,N_8186);
or U15903 (N_15903,N_6891,N_7452);
xnor U15904 (N_15904,N_10263,N_7932);
and U15905 (N_15905,N_9427,N_10360);
nand U15906 (N_15906,N_8618,N_7260);
or U15907 (N_15907,N_7962,N_7979);
nor U15908 (N_15908,N_6818,N_9970);
nor U15909 (N_15909,N_7032,N_9005);
and U15910 (N_15910,N_7594,N_11933);
nor U15911 (N_15911,N_9889,N_10155);
or U15912 (N_15912,N_10253,N_7003);
nor U15913 (N_15913,N_9937,N_11220);
nor U15914 (N_15914,N_9258,N_11935);
and U15915 (N_15915,N_6980,N_11940);
nand U15916 (N_15916,N_6031,N_10770);
or U15917 (N_15917,N_6249,N_7922);
nand U15918 (N_15918,N_7455,N_9066);
xor U15919 (N_15919,N_9258,N_9589);
xnor U15920 (N_15920,N_11176,N_11737);
xor U15921 (N_15921,N_8983,N_7146);
xnor U15922 (N_15922,N_6447,N_8080);
or U15923 (N_15923,N_8610,N_9422);
nand U15924 (N_15924,N_7198,N_11012);
nand U15925 (N_15925,N_8869,N_10333);
and U15926 (N_15926,N_8417,N_11682);
or U15927 (N_15927,N_10432,N_10155);
nor U15928 (N_15928,N_10018,N_8435);
xor U15929 (N_15929,N_11620,N_11323);
and U15930 (N_15930,N_11504,N_11276);
xor U15931 (N_15931,N_7636,N_9307);
nor U15932 (N_15932,N_10248,N_9717);
nand U15933 (N_15933,N_8895,N_10259);
nor U15934 (N_15934,N_10068,N_7637);
xnor U15935 (N_15935,N_8214,N_8250);
and U15936 (N_15936,N_6346,N_9653);
nand U15937 (N_15937,N_10736,N_8679);
or U15938 (N_15938,N_6002,N_9874);
xnor U15939 (N_15939,N_11836,N_11099);
nand U15940 (N_15940,N_7987,N_8394);
nor U15941 (N_15941,N_10893,N_10203);
or U15942 (N_15942,N_8561,N_7998);
nand U15943 (N_15943,N_9953,N_10952);
or U15944 (N_15944,N_7615,N_7852);
nor U15945 (N_15945,N_9876,N_6149);
or U15946 (N_15946,N_9470,N_7463);
nor U15947 (N_15947,N_7622,N_9290);
and U15948 (N_15948,N_7283,N_10764);
and U15949 (N_15949,N_11199,N_11353);
nand U15950 (N_15950,N_8740,N_10859);
or U15951 (N_15951,N_10532,N_9128);
xor U15952 (N_15952,N_8374,N_8162);
xor U15953 (N_15953,N_11179,N_8153);
nand U15954 (N_15954,N_10637,N_6037);
and U15955 (N_15955,N_8541,N_8611);
nand U15956 (N_15956,N_11198,N_11864);
nand U15957 (N_15957,N_10825,N_9971);
or U15958 (N_15958,N_9225,N_6021);
or U15959 (N_15959,N_9209,N_11552);
or U15960 (N_15960,N_11782,N_8812);
and U15961 (N_15961,N_7201,N_6645);
and U15962 (N_15962,N_6386,N_11182);
nand U15963 (N_15963,N_8779,N_6992);
xor U15964 (N_15964,N_7007,N_8232);
and U15965 (N_15965,N_6676,N_6289);
xnor U15966 (N_15966,N_10393,N_10428);
or U15967 (N_15967,N_11554,N_7498);
nand U15968 (N_15968,N_11814,N_6726);
nand U15969 (N_15969,N_11067,N_9771);
nand U15970 (N_15970,N_8204,N_10284);
and U15971 (N_15971,N_6724,N_11097);
or U15972 (N_15972,N_11554,N_8609);
nand U15973 (N_15973,N_9546,N_8339);
and U15974 (N_15974,N_9567,N_10147);
or U15975 (N_15975,N_8626,N_8904);
nand U15976 (N_15976,N_6891,N_10229);
and U15977 (N_15977,N_9736,N_10385);
or U15978 (N_15978,N_8775,N_10059);
nor U15979 (N_15979,N_7326,N_6769);
and U15980 (N_15980,N_6474,N_10716);
and U15981 (N_15981,N_9403,N_9079);
nor U15982 (N_15982,N_6620,N_7814);
and U15983 (N_15983,N_8906,N_6992);
and U15984 (N_15984,N_11538,N_11294);
or U15985 (N_15985,N_8454,N_9324);
nand U15986 (N_15986,N_8257,N_7987);
nand U15987 (N_15987,N_7540,N_11555);
or U15988 (N_15988,N_8459,N_11394);
or U15989 (N_15989,N_7175,N_6882);
nand U15990 (N_15990,N_6810,N_10202);
nor U15991 (N_15991,N_8843,N_7059);
and U15992 (N_15992,N_8753,N_7026);
or U15993 (N_15993,N_11774,N_11866);
or U15994 (N_15994,N_8714,N_10831);
xnor U15995 (N_15995,N_6360,N_6153);
nor U15996 (N_15996,N_7752,N_9344);
nor U15997 (N_15997,N_7969,N_8012);
nand U15998 (N_15998,N_10532,N_8029);
xor U15999 (N_15999,N_8410,N_10629);
xnor U16000 (N_16000,N_11504,N_9241);
nand U16001 (N_16001,N_10741,N_6290);
and U16002 (N_16002,N_10914,N_8310);
nor U16003 (N_16003,N_11266,N_7702);
or U16004 (N_16004,N_11407,N_7079);
and U16005 (N_16005,N_9708,N_7478);
or U16006 (N_16006,N_10364,N_9324);
and U16007 (N_16007,N_8204,N_10341);
nor U16008 (N_16008,N_6537,N_6435);
nand U16009 (N_16009,N_10221,N_10342);
and U16010 (N_16010,N_11191,N_8572);
nand U16011 (N_16011,N_8946,N_9574);
or U16012 (N_16012,N_9325,N_9693);
or U16013 (N_16013,N_11579,N_6091);
and U16014 (N_16014,N_9122,N_7401);
and U16015 (N_16015,N_6993,N_6653);
nand U16016 (N_16016,N_6966,N_8946);
xnor U16017 (N_16017,N_10562,N_6771);
and U16018 (N_16018,N_10355,N_11975);
nand U16019 (N_16019,N_7177,N_7851);
nor U16020 (N_16020,N_9296,N_6008);
xor U16021 (N_16021,N_8199,N_11051);
and U16022 (N_16022,N_7649,N_11497);
nand U16023 (N_16023,N_6190,N_7188);
nand U16024 (N_16024,N_10147,N_8746);
nor U16025 (N_16025,N_9110,N_6061);
xor U16026 (N_16026,N_10492,N_6667);
nor U16027 (N_16027,N_10523,N_10714);
or U16028 (N_16028,N_11699,N_10995);
nor U16029 (N_16029,N_8844,N_7435);
and U16030 (N_16030,N_7903,N_7525);
or U16031 (N_16031,N_10808,N_11482);
nor U16032 (N_16032,N_9957,N_6061);
or U16033 (N_16033,N_9817,N_9542);
and U16034 (N_16034,N_6309,N_11571);
nor U16035 (N_16035,N_9921,N_6677);
xor U16036 (N_16036,N_9993,N_11801);
or U16037 (N_16037,N_6604,N_6964);
nand U16038 (N_16038,N_10950,N_6960);
nor U16039 (N_16039,N_10612,N_7487);
or U16040 (N_16040,N_8511,N_9480);
and U16041 (N_16041,N_6645,N_10263);
nor U16042 (N_16042,N_7841,N_8295);
nand U16043 (N_16043,N_6813,N_10256);
nor U16044 (N_16044,N_8386,N_8803);
and U16045 (N_16045,N_11488,N_6667);
nand U16046 (N_16046,N_10217,N_7864);
nor U16047 (N_16047,N_7330,N_11942);
nor U16048 (N_16048,N_6282,N_7951);
nand U16049 (N_16049,N_10633,N_8934);
and U16050 (N_16050,N_7495,N_10304);
nor U16051 (N_16051,N_9028,N_6105);
and U16052 (N_16052,N_7159,N_8940);
or U16053 (N_16053,N_10538,N_7889);
or U16054 (N_16054,N_9849,N_9036);
xor U16055 (N_16055,N_8820,N_6306);
nor U16056 (N_16056,N_6158,N_7257);
nor U16057 (N_16057,N_8892,N_7984);
xor U16058 (N_16058,N_8811,N_8135);
xor U16059 (N_16059,N_6563,N_6284);
nand U16060 (N_16060,N_10064,N_9112);
or U16061 (N_16061,N_10171,N_8072);
nand U16062 (N_16062,N_10092,N_6714);
and U16063 (N_16063,N_7574,N_10789);
or U16064 (N_16064,N_6681,N_6949);
nor U16065 (N_16065,N_7797,N_9987);
and U16066 (N_16066,N_6831,N_8241);
nor U16067 (N_16067,N_11142,N_10392);
or U16068 (N_16068,N_6145,N_6348);
or U16069 (N_16069,N_11694,N_11883);
xnor U16070 (N_16070,N_8800,N_6011);
nand U16071 (N_16071,N_7597,N_9299);
and U16072 (N_16072,N_7753,N_8510);
nand U16073 (N_16073,N_11830,N_8183);
nand U16074 (N_16074,N_9143,N_9060);
and U16075 (N_16075,N_8410,N_7959);
nor U16076 (N_16076,N_10056,N_8650);
and U16077 (N_16077,N_6418,N_11030);
nand U16078 (N_16078,N_9257,N_7460);
xnor U16079 (N_16079,N_7592,N_6484);
xor U16080 (N_16080,N_6153,N_8383);
nor U16081 (N_16081,N_10001,N_11174);
nor U16082 (N_16082,N_8019,N_11520);
nand U16083 (N_16083,N_8372,N_7214);
nor U16084 (N_16084,N_6074,N_11681);
and U16085 (N_16085,N_11030,N_10760);
and U16086 (N_16086,N_7895,N_6205);
and U16087 (N_16087,N_9552,N_9006);
and U16088 (N_16088,N_10156,N_8481);
nand U16089 (N_16089,N_10619,N_11305);
or U16090 (N_16090,N_10160,N_9715);
nor U16091 (N_16091,N_8391,N_10350);
xor U16092 (N_16092,N_11763,N_9036);
nor U16093 (N_16093,N_10150,N_7888);
nor U16094 (N_16094,N_6722,N_10708);
nand U16095 (N_16095,N_10683,N_8905);
and U16096 (N_16096,N_7154,N_9478);
and U16097 (N_16097,N_8306,N_8880);
xor U16098 (N_16098,N_11001,N_8759);
or U16099 (N_16099,N_6715,N_10811);
nor U16100 (N_16100,N_7208,N_7935);
nor U16101 (N_16101,N_11261,N_6538);
and U16102 (N_16102,N_7626,N_8377);
xnor U16103 (N_16103,N_9634,N_7349);
or U16104 (N_16104,N_8698,N_9195);
or U16105 (N_16105,N_7470,N_8229);
nand U16106 (N_16106,N_11348,N_10969);
and U16107 (N_16107,N_8175,N_7371);
nand U16108 (N_16108,N_7552,N_8071);
or U16109 (N_16109,N_6963,N_8424);
xnor U16110 (N_16110,N_10581,N_7902);
nand U16111 (N_16111,N_8202,N_11483);
and U16112 (N_16112,N_7971,N_9194);
and U16113 (N_16113,N_7795,N_9282);
and U16114 (N_16114,N_9600,N_11156);
nor U16115 (N_16115,N_10055,N_6397);
and U16116 (N_16116,N_11321,N_9970);
nor U16117 (N_16117,N_9820,N_7241);
nor U16118 (N_16118,N_9764,N_10614);
or U16119 (N_16119,N_10615,N_6240);
nand U16120 (N_16120,N_6062,N_9363);
nor U16121 (N_16121,N_10381,N_11653);
and U16122 (N_16122,N_10231,N_6568);
or U16123 (N_16123,N_9036,N_8650);
nand U16124 (N_16124,N_9894,N_11111);
and U16125 (N_16125,N_11222,N_7813);
or U16126 (N_16126,N_9332,N_6630);
nand U16127 (N_16127,N_7492,N_7513);
nor U16128 (N_16128,N_11219,N_7790);
nand U16129 (N_16129,N_9383,N_6690);
nor U16130 (N_16130,N_10905,N_10747);
nor U16131 (N_16131,N_6790,N_10024);
or U16132 (N_16132,N_9246,N_7693);
or U16133 (N_16133,N_10839,N_11726);
or U16134 (N_16134,N_11266,N_10387);
xnor U16135 (N_16135,N_7209,N_8912);
nand U16136 (N_16136,N_11254,N_7051);
or U16137 (N_16137,N_7300,N_7401);
or U16138 (N_16138,N_7159,N_8407);
or U16139 (N_16139,N_7314,N_9066);
or U16140 (N_16140,N_11291,N_7518);
or U16141 (N_16141,N_11702,N_6808);
nand U16142 (N_16142,N_7850,N_6757);
nor U16143 (N_16143,N_9144,N_11832);
nand U16144 (N_16144,N_9225,N_7304);
xnor U16145 (N_16145,N_10429,N_9200);
nand U16146 (N_16146,N_8807,N_6412);
and U16147 (N_16147,N_8050,N_7041);
and U16148 (N_16148,N_6601,N_11975);
xnor U16149 (N_16149,N_10463,N_8080);
nor U16150 (N_16150,N_6116,N_7519);
nor U16151 (N_16151,N_11725,N_9155);
nand U16152 (N_16152,N_6922,N_6047);
nand U16153 (N_16153,N_11153,N_8071);
xnor U16154 (N_16154,N_10850,N_6446);
or U16155 (N_16155,N_6547,N_8909);
nand U16156 (N_16156,N_9880,N_10245);
or U16157 (N_16157,N_10254,N_7672);
and U16158 (N_16158,N_11168,N_10441);
and U16159 (N_16159,N_6825,N_6735);
and U16160 (N_16160,N_6250,N_7711);
or U16161 (N_16161,N_9483,N_9889);
nor U16162 (N_16162,N_11671,N_11326);
and U16163 (N_16163,N_6953,N_6466);
nand U16164 (N_16164,N_11373,N_7645);
xor U16165 (N_16165,N_8200,N_6177);
and U16166 (N_16166,N_11282,N_8651);
xor U16167 (N_16167,N_6893,N_7867);
and U16168 (N_16168,N_9604,N_11467);
nand U16169 (N_16169,N_11115,N_8737);
nor U16170 (N_16170,N_11115,N_7935);
nand U16171 (N_16171,N_7711,N_6362);
nand U16172 (N_16172,N_11479,N_7298);
nand U16173 (N_16173,N_11523,N_8215);
or U16174 (N_16174,N_9569,N_9660);
xor U16175 (N_16175,N_10012,N_11978);
and U16176 (N_16176,N_7608,N_11629);
or U16177 (N_16177,N_7939,N_6682);
or U16178 (N_16178,N_8098,N_8075);
nor U16179 (N_16179,N_11701,N_11334);
nand U16180 (N_16180,N_11104,N_7897);
or U16181 (N_16181,N_10126,N_11921);
and U16182 (N_16182,N_9033,N_11883);
or U16183 (N_16183,N_7372,N_9952);
nor U16184 (N_16184,N_7812,N_11364);
and U16185 (N_16185,N_10852,N_8393);
or U16186 (N_16186,N_7077,N_8618);
or U16187 (N_16187,N_7854,N_9779);
nor U16188 (N_16188,N_10487,N_11696);
xnor U16189 (N_16189,N_7813,N_10208);
nand U16190 (N_16190,N_11474,N_7580);
and U16191 (N_16191,N_11753,N_6786);
nor U16192 (N_16192,N_10567,N_6430);
and U16193 (N_16193,N_6443,N_8422);
xnor U16194 (N_16194,N_6177,N_6352);
nand U16195 (N_16195,N_7918,N_11001);
and U16196 (N_16196,N_11757,N_9315);
or U16197 (N_16197,N_9818,N_6335);
nor U16198 (N_16198,N_11326,N_6030);
xor U16199 (N_16199,N_8471,N_7919);
and U16200 (N_16200,N_8297,N_9725);
or U16201 (N_16201,N_9782,N_11022);
xnor U16202 (N_16202,N_7205,N_9823);
nand U16203 (N_16203,N_9483,N_10229);
nor U16204 (N_16204,N_9784,N_11155);
nor U16205 (N_16205,N_8895,N_8055);
xor U16206 (N_16206,N_11003,N_11260);
or U16207 (N_16207,N_10392,N_9511);
nor U16208 (N_16208,N_7994,N_10254);
nand U16209 (N_16209,N_6707,N_6601);
or U16210 (N_16210,N_6364,N_10331);
or U16211 (N_16211,N_11522,N_9031);
xnor U16212 (N_16212,N_8805,N_8926);
nand U16213 (N_16213,N_9186,N_9768);
or U16214 (N_16214,N_10196,N_7364);
or U16215 (N_16215,N_7484,N_6574);
nand U16216 (N_16216,N_11549,N_7503);
nand U16217 (N_16217,N_6500,N_11844);
or U16218 (N_16218,N_8239,N_6065);
nand U16219 (N_16219,N_11260,N_8840);
nor U16220 (N_16220,N_9572,N_7584);
nor U16221 (N_16221,N_7215,N_11500);
and U16222 (N_16222,N_10311,N_7150);
xor U16223 (N_16223,N_8370,N_11577);
nor U16224 (N_16224,N_6377,N_9278);
and U16225 (N_16225,N_9631,N_9959);
and U16226 (N_16226,N_10891,N_9055);
nor U16227 (N_16227,N_8346,N_8413);
xor U16228 (N_16228,N_10688,N_9511);
nor U16229 (N_16229,N_10424,N_8953);
nor U16230 (N_16230,N_11818,N_9975);
or U16231 (N_16231,N_6598,N_8466);
nand U16232 (N_16232,N_11338,N_6886);
and U16233 (N_16233,N_8850,N_9953);
nor U16234 (N_16234,N_7994,N_7531);
nor U16235 (N_16235,N_11456,N_8936);
and U16236 (N_16236,N_7732,N_9861);
and U16237 (N_16237,N_7192,N_11753);
and U16238 (N_16238,N_10599,N_8494);
nor U16239 (N_16239,N_6292,N_10316);
nand U16240 (N_16240,N_8562,N_10864);
nor U16241 (N_16241,N_9956,N_7590);
or U16242 (N_16242,N_6587,N_6137);
nand U16243 (N_16243,N_6202,N_9610);
nor U16244 (N_16244,N_6939,N_11569);
nand U16245 (N_16245,N_7470,N_6408);
nor U16246 (N_16246,N_8412,N_10876);
nor U16247 (N_16247,N_6926,N_6689);
and U16248 (N_16248,N_7940,N_8922);
and U16249 (N_16249,N_7425,N_10283);
nand U16250 (N_16250,N_8749,N_7809);
or U16251 (N_16251,N_11462,N_11334);
or U16252 (N_16252,N_8498,N_6248);
xnor U16253 (N_16253,N_10946,N_10979);
or U16254 (N_16254,N_11535,N_7696);
or U16255 (N_16255,N_6233,N_6511);
nand U16256 (N_16256,N_10415,N_8029);
xor U16257 (N_16257,N_8219,N_9556);
nor U16258 (N_16258,N_7758,N_9947);
and U16259 (N_16259,N_10523,N_7153);
or U16260 (N_16260,N_10303,N_8287);
or U16261 (N_16261,N_6018,N_10800);
or U16262 (N_16262,N_8359,N_9173);
nand U16263 (N_16263,N_11794,N_8076);
and U16264 (N_16264,N_6258,N_10553);
nand U16265 (N_16265,N_10137,N_9804);
nand U16266 (N_16266,N_6428,N_6631);
and U16267 (N_16267,N_8950,N_8425);
and U16268 (N_16268,N_11566,N_10584);
nor U16269 (N_16269,N_11396,N_11516);
nor U16270 (N_16270,N_9711,N_11201);
nor U16271 (N_16271,N_6430,N_10140);
nor U16272 (N_16272,N_7809,N_9090);
nand U16273 (N_16273,N_9235,N_8540);
or U16274 (N_16274,N_7385,N_8053);
and U16275 (N_16275,N_10187,N_11980);
and U16276 (N_16276,N_7791,N_6903);
nor U16277 (N_16277,N_9300,N_10303);
or U16278 (N_16278,N_7954,N_8681);
nand U16279 (N_16279,N_10248,N_9986);
and U16280 (N_16280,N_10251,N_11001);
or U16281 (N_16281,N_9333,N_6523);
nand U16282 (N_16282,N_8625,N_8883);
and U16283 (N_16283,N_9666,N_8894);
nor U16284 (N_16284,N_6681,N_10439);
nand U16285 (N_16285,N_11540,N_8589);
or U16286 (N_16286,N_11160,N_10411);
xor U16287 (N_16287,N_10133,N_7875);
nor U16288 (N_16288,N_6882,N_7949);
and U16289 (N_16289,N_6072,N_9754);
or U16290 (N_16290,N_11566,N_11651);
nor U16291 (N_16291,N_11761,N_7049);
nor U16292 (N_16292,N_10357,N_11123);
or U16293 (N_16293,N_8151,N_6529);
and U16294 (N_16294,N_9087,N_9119);
and U16295 (N_16295,N_6952,N_8513);
and U16296 (N_16296,N_10322,N_6304);
nor U16297 (N_16297,N_11189,N_9583);
nand U16298 (N_16298,N_8314,N_11396);
nand U16299 (N_16299,N_9450,N_10522);
nor U16300 (N_16300,N_8953,N_10283);
nand U16301 (N_16301,N_11488,N_7895);
and U16302 (N_16302,N_10272,N_10105);
nor U16303 (N_16303,N_7157,N_9813);
xnor U16304 (N_16304,N_11200,N_11625);
and U16305 (N_16305,N_6505,N_7956);
and U16306 (N_16306,N_9889,N_8804);
and U16307 (N_16307,N_8224,N_11514);
nand U16308 (N_16308,N_9477,N_6461);
xor U16309 (N_16309,N_11152,N_11350);
or U16310 (N_16310,N_7293,N_11310);
or U16311 (N_16311,N_6399,N_7300);
and U16312 (N_16312,N_11981,N_6694);
or U16313 (N_16313,N_6239,N_11377);
or U16314 (N_16314,N_11633,N_9476);
and U16315 (N_16315,N_9998,N_11743);
nor U16316 (N_16316,N_7619,N_11623);
and U16317 (N_16317,N_8182,N_8810);
xnor U16318 (N_16318,N_7350,N_8803);
nand U16319 (N_16319,N_7134,N_6733);
xor U16320 (N_16320,N_8361,N_9263);
and U16321 (N_16321,N_7971,N_9005);
and U16322 (N_16322,N_7238,N_11804);
or U16323 (N_16323,N_9057,N_7421);
nand U16324 (N_16324,N_11968,N_9228);
and U16325 (N_16325,N_8667,N_6154);
nand U16326 (N_16326,N_11387,N_10131);
nor U16327 (N_16327,N_10134,N_11283);
nand U16328 (N_16328,N_9256,N_8037);
and U16329 (N_16329,N_11769,N_10198);
or U16330 (N_16330,N_11895,N_7376);
nand U16331 (N_16331,N_9015,N_6145);
xnor U16332 (N_16332,N_8807,N_8289);
nor U16333 (N_16333,N_8913,N_9026);
xnor U16334 (N_16334,N_6469,N_8049);
nand U16335 (N_16335,N_8583,N_10778);
nand U16336 (N_16336,N_6774,N_11374);
nor U16337 (N_16337,N_9244,N_6597);
and U16338 (N_16338,N_9310,N_7411);
and U16339 (N_16339,N_6423,N_9855);
xor U16340 (N_16340,N_10040,N_10423);
nor U16341 (N_16341,N_7623,N_8724);
and U16342 (N_16342,N_6722,N_7867);
or U16343 (N_16343,N_11402,N_11810);
and U16344 (N_16344,N_8246,N_6638);
nand U16345 (N_16345,N_10815,N_7174);
nor U16346 (N_16346,N_11620,N_10865);
nand U16347 (N_16347,N_8573,N_8789);
xor U16348 (N_16348,N_11093,N_7421);
nand U16349 (N_16349,N_11291,N_11797);
xor U16350 (N_16350,N_11535,N_8804);
nand U16351 (N_16351,N_7013,N_8563);
nor U16352 (N_16352,N_7901,N_11728);
xor U16353 (N_16353,N_11108,N_8408);
nand U16354 (N_16354,N_11986,N_11734);
nor U16355 (N_16355,N_10151,N_6444);
nor U16356 (N_16356,N_9189,N_8233);
or U16357 (N_16357,N_10683,N_10282);
nor U16358 (N_16358,N_6100,N_11460);
nand U16359 (N_16359,N_11496,N_10350);
nor U16360 (N_16360,N_9847,N_8512);
and U16361 (N_16361,N_10434,N_9678);
or U16362 (N_16362,N_6000,N_9516);
nand U16363 (N_16363,N_8767,N_8197);
or U16364 (N_16364,N_10996,N_7308);
nor U16365 (N_16365,N_9736,N_11137);
xor U16366 (N_16366,N_10931,N_6048);
nor U16367 (N_16367,N_7419,N_6716);
nor U16368 (N_16368,N_6768,N_8101);
nor U16369 (N_16369,N_10257,N_7890);
nor U16370 (N_16370,N_7342,N_6972);
nor U16371 (N_16371,N_6021,N_6789);
nand U16372 (N_16372,N_8900,N_11292);
nand U16373 (N_16373,N_9397,N_11784);
nor U16374 (N_16374,N_11819,N_10496);
and U16375 (N_16375,N_9960,N_10862);
nand U16376 (N_16376,N_10607,N_8933);
and U16377 (N_16377,N_6252,N_8772);
or U16378 (N_16378,N_11664,N_10639);
and U16379 (N_16379,N_6963,N_6845);
and U16380 (N_16380,N_9962,N_10230);
nand U16381 (N_16381,N_9160,N_7963);
nand U16382 (N_16382,N_10471,N_10210);
nor U16383 (N_16383,N_10053,N_11601);
or U16384 (N_16384,N_8278,N_8929);
xnor U16385 (N_16385,N_7010,N_11445);
or U16386 (N_16386,N_11317,N_9175);
or U16387 (N_16387,N_10311,N_11671);
nor U16388 (N_16388,N_11023,N_6856);
and U16389 (N_16389,N_8991,N_8967);
nor U16390 (N_16390,N_10569,N_6862);
and U16391 (N_16391,N_9193,N_10995);
or U16392 (N_16392,N_11293,N_6936);
nand U16393 (N_16393,N_8466,N_8149);
or U16394 (N_16394,N_11160,N_8504);
nand U16395 (N_16395,N_10018,N_7902);
nor U16396 (N_16396,N_9271,N_9071);
and U16397 (N_16397,N_9034,N_8979);
nand U16398 (N_16398,N_9805,N_10032);
and U16399 (N_16399,N_11793,N_11246);
nor U16400 (N_16400,N_11003,N_7740);
and U16401 (N_16401,N_6238,N_11658);
or U16402 (N_16402,N_9688,N_9607);
and U16403 (N_16403,N_7603,N_6194);
xor U16404 (N_16404,N_9836,N_10977);
nand U16405 (N_16405,N_9049,N_10519);
nand U16406 (N_16406,N_11569,N_7016);
nand U16407 (N_16407,N_10397,N_7260);
nor U16408 (N_16408,N_7221,N_11650);
nand U16409 (N_16409,N_9014,N_6288);
or U16410 (N_16410,N_10396,N_10357);
nor U16411 (N_16411,N_9019,N_10003);
nor U16412 (N_16412,N_10917,N_8152);
or U16413 (N_16413,N_9377,N_10873);
nor U16414 (N_16414,N_10813,N_11221);
and U16415 (N_16415,N_8117,N_9264);
xnor U16416 (N_16416,N_9721,N_6101);
nor U16417 (N_16417,N_6792,N_11064);
nor U16418 (N_16418,N_8541,N_10421);
nand U16419 (N_16419,N_9914,N_6715);
or U16420 (N_16420,N_10074,N_7092);
and U16421 (N_16421,N_10854,N_11880);
nor U16422 (N_16422,N_11322,N_10783);
and U16423 (N_16423,N_8897,N_8259);
xor U16424 (N_16424,N_6054,N_6498);
and U16425 (N_16425,N_11062,N_8494);
nand U16426 (N_16426,N_8872,N_9054);
and U16427 (N_16427,N_9457,N_11751);
or U16428 (N_16428,N_8955,N_10702);
and U16429 (N_16429,N_11987,N_6009);
nor U16430 (N_16430,N_10340,N_10629);
xnor U16431 (N_16431,N_7201,N_7443);
xnor U16432 (N_16432,N_10010,N_9022);
or U16433 (N_16433,N_6742,N_6572);
nor U16434 (N_16434,N_7638,N_8956);
nor U16435 (N_16435,N_11704,N_10824);
and U16436 (N_16436,N_10349,N_7170);
xnor U16437 (N_16437,N_7581,N_10156);
xnor U16438 (N_16438,N_6353,N_11268);
and U16439 (N_16439,N_7439,N_8567);
or U16440 (N_16440,N_7346,N_8460);
nand U16441 (N_16441,N_7394,N_10436);
or U16442 (N_16442,N_10134,N_6421);
or U16443 (N_16443,N_8569,N_11168);
nor U16444 (N_16444,N_9393,N_6274);
or U16445 (N_16445,N_6490,N_7230);
and U16446 (N_16446,N_7257,N_8886);
nor U16447 (N_16447,N_7298,N_7279);
nor U16448 (N_16448,N_9321,N_9464);
or U16449 (N_16449,N_9479,N_11284);
nand U16450 (N_16450,N_6081,N_9500);
xor U16451 (N_16451,N_11399,N_6915);
and U16452 (N_16452,N_6068,N_7189);
nand U16453 (N_16453,N_8422,N_8805);
nor U16454 (N_16454,N_8578,N_9565);
nor U16455 (N_16455,N_11562,N_8427);
xor U16456 (N_16456,N_7283,N_7313);
nand U16457 (N_16457,N_8663,N_8836);
and U16458 (N_16458,N_10786,N_6125);
nor U16459 (N_16459,N_9363,N_7335);
xor U16460 (N_16460,N_6901,N_7687);
nor U16461 (N_16461,N_8477,N_9681);
and U16462 (N_16462,N_9031,N_6924);
nor U16463 (N_16463,N_8138,N_10859);
nor U16464 (N_16464,N_6045,N_10942);
and U16465 (N_16465,N_7684,N_7698);
or U16466 (N_16466,N_11144,N_9770);
nand U16467 (N_16467,N_9149,N_6293);
nor U16468 (N_16468,N_8690,N_7843);
nor U16469 (N_16469,N_10052,N_8403);
nor U16470 (N_16470,N_9525,N_11349);
xor U16471 (N_16471,N_7052,N_8108);
nand U16472 (N_16472,N_7760,N_9927);
and U16473 (N_16473,N_8144,N_7790);
or U16474 (N_16474,N_10061,N_11758);
nand U16475 (N_16475,N_8155,N_9456);
xor U16476 (N_16476,N_9124,N_11561);
nand U16477 (N_16477,N_9663,N_11975);
or U16478 (N_16478,N_10335,N_8916);
or U16479 (N_16479,N_11374,N_9871);
and U16480 (N_16480,N_11737,N_11487);
nor U16481 (N_16481,N_9520,N_8007);
or U16482 (N_16482,N_6346,N_8618);
nor U16483 (N_16483,N_6087,N_7007);
or U16484 (N_16484,N_7672,N_9580);
nor U16485 (N_16485,N_6292,N_8964);
and U16486 (N_16486,N_8990,N_8982);
nor U16487 (N_16487,N_10491,N_6214);
or U16488 (N_16488,N_11828,N_10827);
nand U16489 (N_16489,N_6989,N_7007);
or U16490 (N_16490,N_11047,N_10524);
nand U16491 (N_16491,N_6252,N_11489);
and U16492 (N_16492,N_7722,N_10637);
nand U16493 (N_16493,N_11177,N_10224);
nor U16494 (N_16494,N_10971,N_10426);
nor U16495 (N_16495,N_11976,N_8490);
nand U16496 (N_16496,N_7941,N_9171);
or U16497 (N_16497,N_8431,N_7521);
nor U16498 (N_16498,N_10591,N_11876);
xnor U16499 (N_16499,N_9936,N_9383);
and U16500 (N_16500,N_8162,N_11398);
nand U16501 (N_16501,N_8805,N_8140);
or U16502 (N_16502,N_7922,N_8442);
nor U16503 (N_16503,N_11839,N_11470);
nor U16504 (N_16504,N_6868,N_10227);
nand U16505 (N_16505,N_11968,N_11989);
or U16506 (N_16506,N_9804,N_7902);
or U16507 (N_16507,N_7100,N_6304);
nand U16508 (N_16508,N_10238,N_6996);
xnor U16509 (N_16509,N_8533,N_7285);
nor U16510 (N_16510,N_6850,N_9865);
nand U16511 (N_16511,N_8396,N_6419);
nor U16512 (N_16512,N_10494,N_9333);
or U16513 (N_16513,N_9033,N_7916);
and U16514 (N_16514,N_9877,N_7486);
nor U16515 (N_16515,N_11096,N_8148);
and U16516 (N_16516,N_8742,N_8647);
nand U16517 (N_16517,N_11804,N_6620);
and U16518 (N_16518,N_7723,N_7039);
nand U16519 (N_16519,N_9727,N_9038);
and U16520 (N_16520,N_7178,N_11762);
nor U16521 (N_16521,N_7257,N_10900);
nor U16522 (N_16522,N_6089,N_8911);
or U16523 (N_16523,N_8442,N_7002);
nand U16524 (N_16524,N_6268,N_11127);
nor U16525 (N_16525,N_9029,N_7242);
and U16526 (N_16526,N_10762,N_8391);
and U16527 (N_16527,N_8808,N_6445);
and U16528 (N_16528,N_10630,N_11589);
or U16529 (N_16529,N_10955,N_6952);
and U16530 (N_16530,N_9730,N_9696);
nand U16531 (N_16531,N_9432,N_6945);
xnor U16532 (N_16532,N_6320,N_10322);
nand U16533 (N_16533,N_6954,N_8567);
xor U16534 (N_16534,N_6949,N_7706);
and U16535 (N_16535,N_9675,N_10117);
xor U16536 (N_16536,N_10118,N_6352);
nand U16537 (N_16537,N_8525,N_6106);
xor U16538 (N_16538,N_11603,N_7614);
nand U16539 (N_16539,N_9164,N_7825);
nand U16540 (N_16540,N_9604,N_7507);
or U16541 (N_16541,N_11254,N_10195);
xnor U16542 (N_16542,N_10819,N_10277);
and U16543 (N_16543,N_8166,N_9984);
nand U16544 (N_16544,N_7395,N_11812);
nand U16545 (N_16545,N_7221,N_10176);
or U16546 (N_16546,N_6134,N_6633);
nand U16547 (N_16547,N_11141,N_9030);
nor U16548 (N_16548,N_10381,N_11331);
nand U16549 (N_16549,N_6694,N_7655);
or U16550 (N_16550,N_7916,N_10554);
xnor U16551 (N_16551,N_6462,N_8747);
nor U16552 (N_16552,N_11923,N_11993);
nand U16553 (N_16553,N_8080,N_7597);
nor U16554 (N_16554,N_8403,N_7579);
nor U16555 (N_16555,N_11797,N_7717);
nand U16556 (N_16556,N_11774,N_7026);
nand U16557 (N_16557,N_11512,N_10516);
nand U16558 (N_16558,N_11501,N_7353);
xor U16559 (N_16559,N_11647,N_8379);
and U16560 (N_16560,N_7541,N_10933);
xnor U16561 (N_16561,N_11966,N_8422);
xnor U16562 (N_16562,N_9493,N_11645);
or U16563 (N_16563,N_7233,N_11257);
nor U16564 (N_16564,N_7331,N_6476);
xnor U16565 (N_16565,N_7884,N_9022);
xor U16566 (N_16566,N_7597,N_8142);
nor U16567 (N_16567,N_11325,N_10565);
nor U16568 (N_16568,N_10234,N_7503);
and U16569 (N_16569,N_6706,N_9737);
nor U16570 (N_16570,N_6064,N_7801);
nor U16571 (N_16571,N_6176,N_7282);
nor U16572 (N_16572,N_7726,N_6662);
or U16573 (N_16573,N_7257,N_10109);
nand U16574 (N_16574,N_7607,N_10502);
or U16575 (N_16575,N_9268,N_6352);
or U16576 (N_16576,N_6482,N_10586);
or U16577 (N_16577,N_6325,N_8279);
or U16578 (N_16578,N_9093,N_8154);
and U16579 (N_16579,N_6738,N_10023);
and U16580 (N_16580,N_6928,N_9620);
nor U16581 (N_16581,N_9835,N_10928);
nor U16582 (N_16582,N_10211,N_9068);
and U16583 (N_16583,N_9921,N_9663);
or U16584 (N_16584,N_9504,N_8400);
nor U16585 (N_16585,N_11599,N_10342);
or U16586 (N_16586,N_6361,N_7478);
and U16587 (N_16587,N_10414,N_8812);
or U16588 (N_16588,N_10942,N_8250);
and U16589 (N_16589,N_8604,N_11400);
nor U16590 (N_16590,N_9908,N_7469);
nor U16591 (N_16591,N_10778,N_11494);
and U16592 (N_16592,N_7807,N_10549);
xnor U16593 (N_16593,N_10184,N_6313);
xor U16594 (N_16594,N_11572,N_11853);
and U16595 (N_16595,N_11307,N_10654);
and U16596 (N_16596,N_6352,N_9698);
nand U16597 (N_16597,N_10138,N_11183);
nor U16598 (N_16598,N_8925,N_9822);
nor U16599 (N_16599,N_9684,N_10209);
nand U16600 (N_16600,N_8283,N_7173);
nor U16601 (N_16601,N_7326,N_11318);
nor U16602 (N_16602,N_11703,N_6036);
xnor U16603 (N_16603,N_10655,N_10054);
nor U16604 (N_16604,N_9820,N_7708);
nor U16605 (N_16605,N_11403,N_11702);
nand U16606 (N_16606,N_8822,N_7942);
nor U16607 (N_16607,N_6524,N_8687);
nor U16608 (N_16608,N_10762,N_11018);
and U16609 (N_16609,N_9313,N_6062);
nand U16610 (N_16610,N_7724,N_7514);
and U16611 (N_16611,N_10181,N_6267);
nor U16612 (N_16612,N_7433,N_9012);
nor U16613 (N_16613,N_8245,N_6754);
and U16614 (N_16614,N_11769,N_6824);
nor U16615 (N_16615,N_10595,N_7893);
nor U16616 (N_16616,N_11951,N_6273);
or U16617 (N_16617,N_8267,N_9281);
or U16618 (N_16618,N_9504,N_7474);
nand U16619 (N_16619,N_9109,N_7369);
xor U16620 (N_16620,N_10768,N_10166);
nor U16621 (N_16621,N_6970,N_9138);
and U16622 (N_16622,N_9132,N_7760);
nand U16623 (N_16623,N_10326,N_10864);
nor U16624 (N_16624,N_11931,N_9384);
or U16625 (N_16625,N_8005,N_8147);
or U16626 (N_16626,N_8205,N_8467);
xnor U16627 (N_16627,N_11735,N_9287);
xor U16628 (N_16628,N_8680,N_6510);
nor U16629 (N_16629,N_9291,N_11210);
nand U16630 (N_16630,N_8285,N_8677);
nand U16631 (N_16631,N_8205,N_10466);
xor U16632 (N_16632,N_7396,N_8915);
xnor U16633 (N_16633,N_10827,N_6641);
or U16634 (N_16634,N_10889,N_8792);
xnor U16635 (N_16635,N_6070,N_8436);
and U16636 (N_16636,N_9587,N_11957);
xnor U16637 (N_16637,N_10244,N_11938);
nor U16638 (N_16638,N_9620,N_7150);
nor U16639 (N_16639,N_6671,N_9045);
nand U16640 (N_16640,N_11067,N_8402);
and U16641 (N_16641,N_10616,N_6593);
and U16642 (N_16642,N_6249,N_9407);
nand U16643 (N_16643,N_10854,N_6602);
and U16644 (N_16644,N_7677,N_8004);
xnor U16645 (N_16645,N_8784,N_11979);
or U16646 (N_16646,N_6733,N_7711);
nor U16647 (N_16647,N_11317,N_9073);
or U16648 (N_16648,N_6760,N_11669);
xor U16649 (N_16649,N_10432,N_8488);
or U16650 (N_16650,N_6484,N_6162);
nor U16651 (N_16651,N_7547,N_6650);
nand U16652 (N_16652,N_10139,N_6409);
and U16653 (N_16653,N_8027,N_8044);
and U16654 (N_16654,N_9184,N_11382);
and U16655 (N_16655,N_10954,N_7635);
or U16656 (N_16656,N_10299,N_7017);
and U16657 (N_16657,N_10083,N_8417);
nand U16658 (N_16658,N_6875,N_10440);
nand U16659 (N_16659,N_10189,N_11825);
or U16660 (N_16660,N_6826,N_9418);
nor U16661 (N_16661,N_11275,N_7020);
and U16662 (N_16662,N_11076,N_7532);
or U16663 (N_16663,N_8436,N_11173);
nor U16664 (N_16664,N_6717,N_8763);
nor U16665 (N_16665,N_10106,N_8154);
nand U16666 (N_16666,N_10492,N_8500);
and U16667 (N_16667,N_11350,N_8253);
or U16668 (N_16668,N_7499,N_6547);
or U16669 (N_16669,N_9210,N_10318);
or U16670 (N_16670,N_9700,N_9740);
nor U16671 (N_16671,N_8757,N_9712);
nor U16672 (N_16672,N_8403,N_10239);
nor U16673 (N_16673,N_7876,N_8010);
nor U16674 (N_16674,N_7744,N_9795);
and U16675 (N_16675,N_10516,N_6124);
nor U16676 (N_16676,N_8511,N_7478);
xor U16677 (N_16677,N_7003,N_6925);
or U16678 (N_16678,N_11595,N_11602);
and U16679 (N_16679,N_6735,N_8464);
nand U16680 (N_16680,N_10383,N_11295);
nor U16681 (N_16681,N_11394,N_6982);
nor U16682 (N_16682,N_11263,N_9084);
or U16683 (N_16683,N_11892,N_11296);
nand U16684 (N_16684,N_10583,N_10335);
or U16685 (N_16685,N_11530,N_8928);
nand U16686 (N_16686,N_7369,N_8194);
nor U16687 (N_16687,N_9699,N_10889);
nand U16688 (N_16688,N_6873,N_8783);
or U16689 (N_16689,N_7423,N_9147);
or U16690 (N_16690,N_9545,N_6931);
and U16691 (N_16691,N_7995,N_10740);
or U16692 (N_16692,N_9896,N_6455);
or U16693 (N_16693,N_10578,N_6332);
nand U16694 (N_16694,N_10188,N_11862);
and U16695 (N_16695,N_11275,N_7184);
nand U16696 (N_16696,N_7013,N_6832);
and U16697 (N_16697,N_9037,N_10199);
xor U16698 (N_16698,N_10335,N_11801);
nand U16699 (N_16699,N_11589,N_6512);
xor U16700 (N_16700,N_11909,N_9026);
and U16701 (N_16701,N_8267,N_11205);
or U16702 (N_16702,N_8355,N_8306);
and U16703 (N_16703,N_11480,N_10303);
nor U16704 (N_16704,N_11901,N_10409);
and U16705 (N_16705,N_6887,N_11246);
nor U16706 (N_16706,N_9321,N_9789);
nand U16707 (N_16707,N_10203,N_9109);
or U16708 (N_16708,N_7800,N_10129);
or U16709 (N_16709,N_10664,N_9324);
and U16710 (N_16710,N_9117,N_6368);
nor U16711 (N_16711,N_9813,N_9885);
nand U16712 (N_16712,N_9581,N_9939);
and U16713 (N_16713,N_8344,N_6123);
and U16714 (N_16714,N_11286,N_8294);
xor U16715 (N_16715,N_7304,N_11603);
xnor U16716 (N_16716,N_10816,N_7744);
nand U16717 (N_16717,N_9960,N_7244);
and U16718 (N_16718,N_6379,N_6883);
nor U16719 (N_16719,N_9804,N_6091);
nor U16720 (N_16720,N_8387,N_6130);
and U16721 (N_16721,N_11914,N_7799);
xnor U16722 (N_16722,N_7850,N_8616);
nand U16723 (N_16723,N_7258,N_11875);
nor U16724 (N_16724,N_6757,N_9617);
and U16725 (N_16725,N_11753,N_11351);
and U16726 (N_16726,N_9103,N_7639);
xor U16727 (N_16727,N_6510,N_7314);
nand U16728 (N_16728,N_7987,N_10885);
nor U16729 (N_16729,N_8468,N_10320);
and U16730 (N_16730,N_6882,N_11160);
and U16731 (N_16731,N_11587,N_10697);
and U16732 (N_16732,N_7019,N_8137);
nor U16733 (N_16733,N_8946,N_9784);
xnor U16734 (N_16734,N_11580,N_8592);
nand U16735 (N_16735,N_9314,N_9312);
and U16736 (N_16736,N_7614,N_9954);
nor U16737 (N_16737,N_11414,N_6450);
and U16738 (N_16738,N_7310,N_7485);
nor U16739 (N_16739,N_7194,N_9571);
and U16740 (N_16740,N_10799,N_10550);
nand U16741 (N_16741,N_6281,N_10043);
nand U16742 (N_16742,N_11155,N_8320);
nor U16743 (N_16743,N_8388,N_10114);
or U16744 (N_16744,N_6506,N_9661);
xnor U16745 (N_16745,N_10391,N_10004);
nor U16746 (N_16746,N_11368,N_7619);
and U16747 (N_16747,N_10616,N_10617);
nor U16748 (N_16748,N_11546,N_7674);
nor U16749 (N_16749,N_6433,N_9928);
or U16750 (N_16750,N_7737,N_11634);
nand U16751 (N_16751,N_7823,N_6405);
or U16752 (N_16752,N_7820,N_8091);
or U16753 (N_16753,N_6921,N_7985);
nand U16754 (N_16754,N_11057,N_9658);
or U16755 (N_16755,N_8830,N_8516);
nand U16756 (N_16756,N_11861,N_11909);
nor U16757 (N_16757,N_9941,N_10556);
or U16758 (N_16758,N_7709,N_8183);
nor U16759 (N_16759,N_8111,N_8156);
nand U16760 (N_16760,N_7441,N_8331);
nand U16761 (N_16761,N_11247,N_9734);
or U16762 (N_16762,N_10591,N_11778);
and U16763 (N_16763,N_11723,N_10627);
or U16764 (N_16764,N_9431,N_9747);
xor U16765 (N_16765,N_10763,N_8495);
or U16766 (N_16766,N_7590,N_9922);
nand U16767 (N_16767,N_10722,N_10650);
and U16768 (N_16768,N_11680,N_6287);
or U16769 (N_16769,N_8836,N_7743);
nor U16770 (N_16770,N_9851,N_8789);
or U16771 (N_16771,N_9297,N_7135);
or U16772 (N_16772,N_6155,N_6546);
nand U16773 (N_16773,N_6915,N_7520);
or U16774 (N_16774,N_8758,N_11328);
nor U16775 (N_16775,N_11500,N_10529);
nor U16776 (N_16776,N_6673,N_6048);
nor U16777 (N_16777,N_7157,N_8940);
nor U16778 (N_16778,N_9112,N_8607);
nor U16779 (N_16779,N_8700,N_10618);
nand U16780 (N_16780,N_11545,N_6766);
xnor U16781 (N_16781,N_9134,N_10647);
nand U16782 (N_16782,N_9560,N_8331);
nor U16783 (N_16783,N_7658,N_8389);
and U16784 (N_16784,N_8825,N_8606);
and U16785 (N_16785,N_6959,N_7796);
or U16786 (N_16786,N_8953,N_11282);
and U16787 (N_16787,N_9384,N_9253);
nand U16788 (N_16788,N_11987,N_11753);
nand U16789 (N_16789,N_7671,N_6206);
xnor U16790 (N_16790,N_8422,N_8889);
and U16791 (N_16791,N_8852,N_11284);
nand U16792 (N_16792,N_9344,N_6107);
nor U16793 (N_16793,N_8522,N_9002);
and U16794 (N_16794,N_10814,N_9241);
nor U16795 (N_16795,N_11465,N_10415);
nand U16796 (N_16796,N_11464,N_7424);
nand U16797 (N_16797,N_7082,N_11329);
and U16798 (N_16798,N_9754,N_8915);
xor U16799 (N_16799,N_8862,N_10008);
or U16800 (N_16800,N_9733,N_8497);
or U16801 (N_16801,N_9112,N_6687);
xnor U16802 (N_16802,N_11483,N_8469);
nand U16803 (N_16803,N_7333,N_10894);
or U16804 (N_16804,N_10621,N_10241);
nor U16805 (N_16805,N_8057,N_6968);
and U16806 (N_16806,N_11190,N_7126);
and U16807 (N_16807,N_10530,N_9470);
nor U16808 (N_16808,N_11484,N_7412);
nand U16809 (N_16809,N_10409,N_8686);
or U16810 (N_16810,N_7560,N_9018);
or U16811 (N_16811,N_10409,N_6168);
xor U16812 (N_16812,N_6250,N_7037);
nand U16813 (N_16813,N_7259,N_9665);
nand U16814 (N_16814,N_8831,N_7554);
or U16815 (N_16815,N_7239,N_7922);
nand U16816 (N_16816,N_11447,N_11144);
and U16817 (N_16817,N_6170,N_11140);
xor U16818 (N_16818,N_8362,N_6690);
nor U16819 (N_16819,N_11609,N_11422);
nand U16820 (N_16820,N_9257,N_7629);
nor U16821 (N_16821,N_8770,N_6195);
nand U16822 (N_16822,N_10443,N_11198);
and U16823 (N_16823,N_9269,N_9721);
nor U16824 (N_16824,N_9434,N_10864);
nor U16825 (N_16825,N_11657,N_6402);
and U16826 (N_16826,N_6358,N_6785);
and U16827 (N_16827,N_7115,N_9274);
nand U16828 (N_16828,N_8441,N_10459);
nand U16829 (N_16829,N_11897,N_7886);
or U16830 (N_16830,N_11219,N_11085);
nand U16831 (N_16831,N_10935,N_7833);
and U16832 (N_16832,N_8279,N_11577);
or U16833 (N_16833,N_6693,N_9039);
nand U16834 (N_16834,N_7698,N_9337);
and U16835 (N_16835,N_9086,N_10482);
nand U16836 (N_16836,N_10671,N_6938);
nor U16837 (N_16837,N_11296,N_11947);
nor U16838 (N_16838,N_7904,N_8751);
nor U16839 (N_16839,N_7369,N_8489);
and U16840 (N_16840,N_9753,N_10391);
nand U16841 (N_16841,N_6884,N_6809);
nand U16842 (N_16842,N_6516,N_7252);
or U16843 (N_16843,N_9142,N_9173);
nor U16844 (N_16844,N_9272,N_8005);
nand U16845 (N_16845,N_6756,N_10312);
and U16846 (N_16846,N_9818,N_9020);
and U16847 (N_16847,N_10621,N_8148);
nor U16848 (N_16848,N_7009,N_7881);
and U16849 (N_16849,N_6123,N_8659);
nor U16850 (N_16850,N_9286,N_10001);
nor U16851 (N_16851,N_7224,N_7676);
or U16852 (N_16852,N_11566,N_11408);
nor U16853 (N_16853,N_9356,N_9479);
or U16854 (N_16854,N_7206,N_7877);
and U16855 (N_16855,N_7324,N_10087);
and U16856 (N_16856,N_11150,N_9645);
or U16857 (N_16857,N_9462,N_9148);
nand U16858 (N_16858,N_9230,N_10393);
or U16859 (N_16859,N_9867,N_11762);
nand U16860 (N_16860,N_7118,N_11508);
nand U16861 (N_16861,N_7907,N_10327);
nand U16862 (N_16862,N_7734,N_10146);
nor U16863 (N_16863,N_6311,N_11002);
nand U16864 (N_16864,N_7560,N_10809);
or U16865 (N_16865,N_7801,N_11977);
and U16866 (N_16866,N_6156,N_7674);
and U16867 (N_16867,N_8645,N_8991);
and U16868 (N_16868,N_9616,N_8909);
nand U16869 (N_16869,N_9688,N_8068);
xor U16870 (N_16870,N_6873,N_8031);
nand U16871 (N_16871,N_9846,N_8192);
nor U16872 (N_16872,N_9229,N_10023);
or U16873 (N_16873,N_7124,N_7599);
nand U16874 (N_16874,N_6277,N_7161);
nor U16875 (N_16875,N_7643,N_9744);
and U16876 (N_16876,N_10186,N_6985);
nor U16877 (N_16877,N_11922,N_10172);
or U16878 (N_16878,N_6662,N_10997);
nor U16879 (N_16879,N_6953,N_6036);
and U16880 (N_16880,N_7929,N_10089);
and U16881 (N_16881,N_7733,N_8298);
or U16882 (N_16882,N_7723,N_9944);
or U16883 (N_16883,N_8983,N_10046);
and U16884 (N_16884,N_10835,N_7631);
nor U16885 (N_16885,N_7101,N_7698);
or U16886 (N_16886,N_11209,N_6984);
and U16887 (N_16887,N_6939,N_8692);
nand U16888 (N_16888,N_11647,N_9226);
nand U16889 (N_16889,N_8325,N_11310);
nor U16890 (N_16890,N_10507,N_7094);
and U16891 (N_16891,N_11712,N_10068);
and U16892 (N_16892,N_8521,N_7865);
nand U16893 (N_16893,N_9321,N_8302);
or U16894 (N_16894,N_8729,N_7530);
nor U16895 (N_16895,N_10325,N_9059);
or U16896 (N_16896,N_9981,N_10270);
or U16897 (N_16897,N_8483,N_7052);
or U16898 (N_16898,N_9946,N_6009);
nand U16899 (N_16899,N_11789,N_7557);
nor U16900 (N_16900,N_10624,N_7383);
and U16901 (N_16901,N_6405,N_6854);
or U16902 (N_16902,N_8364,N_9198);
and U16903 (N_16903,N_8077,N_10185);
nand U16904 (N_16904,N_11015,N_6763);
and U16905 (N_16905,N_8856,N_11452);
nand U16906 (N_16906,N_7252,N_11669);
or U16907 (N_16907,N_9246,N_8523);
nor U16908 (N_16908,N_10727,N_6302);
and U16909 (N_16909,N_7038,N_7923);
nor U16910 (N_16910,N_9478,N_7454);
and U16911 (N_16911,N_11534,N_7704);
or U16912 (N_16912,N_11628,N_11061);
or U16913 (N_16913,N_9848,N_6820);
nand U16914 (N_16914,N_7991,N_10121);
and U16915 (N_16915,N_8851,N_8617);
and U16916 (N_16916,N_9893,N_7451);
nand U16917 (N_16917,N_9866,N_9618);
nor U16918 (N_16918,N_6529,N_10577);
nor U16919 (N_16919,N_10866,N_7470);
xor U16920 (N_16920,N_10693,N_6826);
nor U16921 (N_16921,N_6400,N_11629);
and U16922 (N_16922,N_10498,N_6637);
nor U16923 (N_16923,N_6593,N_11938);
nor U16924 (N_16924,N_6124,N_7052);
or U16925 (N_16925,N_7027,N_10205);
and U16926 (N_16926,N_11940,N_7691);
nand U16927 (N_16927,N_10947,N_10781);
nand U16928 (N_16928,N_8206,N_11990);
and U16929 (N_16929,N_8222,N_8972);
or U16930 (N_16930,N_8887,N_8170);
or U16931 (N_16931,N_11743,N_10568);
nand U16932 (N_16932,N_10799,N_8630);
nor U16933 (N_16933,N_9008,N_9218);
and U16934 (N_16934,N_9042,N_9309);
or U16935 (N_16935,N_7361,N_7731);
nand U16936 (N_16936,N_11086,N_9259);
nor U16937 (N_16937,N_10444,N_7135);
and U16938 (N_16938,N_7685,N_9095);
and U16939 (N_16939,N_9684,N_8758);
nand U16940 (N_16940,N_6422,N_8007);
or U16941 (N_16941,N_6980,N_11213);
nand U16942 (N_16942,N_8882,N_7068);
nor U16943 (N_16943,N_10600,N_11170);
xnor U16944 (N_16944,N_6627,N_7555);
nand U16945 (N_16945,N_6758,N_11022);
nor U16946 (N_16946,N_9166,N_9704);
and U16947 (N_16947,N_11250,N_11772);
and U16948 (N_16948,N_11557,N_7012);
nor U16949 (N_16949,N_9299,N_7720);
nand U16950 (N_16950,N_11684,N_10952);
or U16951 (N_16951,N_10681,N_9795);
or U16952 (N_16952,N_7418,N_9568);
nand U16953 (N_16953,N_7231,N_9475);
or U16954 (N_16954,N_10724,N_7462);
xor U16955 (N_16955,N_10257,N_6573);
xnor U16956 (N_16956,N_8420,N_9554);
and U16957 (N_16957,N_11503,N_7244);
or U16958 (N_16958,N_10549,N_7894);
nor U16959 (N_16959,N_7797,N_7956);
and U16960 (N_16960,N_11650,N_6692);
and U16961 (N_16961,N_7068,N_7570);
nand U16962 (N_16962,N_9567,N_10602);
nor U16963 (N_16963,N_9697,N_9055);
and U16964 (N_16964,N_11123,N_11561);
nor U16965 (N_16965,N_11039,N_8263);
or U16966 (N_16966,N_11470,N_11701);
or U16967 (N_16967,N_11895,N_11731);
nand U16968 (N_16968,N_6756,N_8032);
xor U16969 (N_16969,N_9138,N_10669);
nand U16970 (N_16970,N_7475,N_8827);
or U16971 (N_16971,N_6036,N_7296);
nand U16972 (N_16972,N_7295,N_6828);
nor U16973 (N_16973,N_10280,N_10207);
or U16974 (N_16974,N_7596,N_10407);
or U16975 (N_16975,N_8356,N_9830);
or U16976 (N_16976,N_10098,N_6106);
or U16977 (N_16977,N_9621,N_8280);
or U16978 (N_16978,N_11298,N_9934);
or U16979 (N_16979,N_10051,N_8744);
or U16980 (N_16980,N_9958,N_9154);
nor U16981 (N_16981,N_6971,N_7239);
xor U16982 (N_16982,N_8245,N_11667);
nand U16983 (N_16983,N_8050,N_10699);
nor U16984 (N_16984,N_7126,N_7849);
nor U16985 (N_16985,N_10144,N_8447);
nor U16986 (N_16986,N_9906,N_8774);
and U16987 (N_16987,N_7141,N_8142);
nor U16988 (N_16988,N_7087,N_7827);
and U16989 (N_16989,N_7539,N_6770);
nand U16990 (N_16990,N_10561,N_8937);
and U16991 (N_16991,N_8869,N_7072);
nand U16992 (N_16992,N_7784,N_6429);
nand U16993 (N_16993,N_11290,N_7466);
and U16994 (N_16994,N_11340,N_7465);
and U16995 (N_16995,N_10615,N_6071);
and U16996 (N_16996,N_6771,N_11628);
xor U16997 (N_16997,N_10775,N_11706);
nand U16998 (N_16998,N_7896,N_6470);
or U16999 (N_16999,N_10367,N_9280);
nor U17000 (N_17000,N_9058,N_10300);
or U17001 (N_17001,N_10797,N_11714);
nand U17002 (N_17002,N_9218,N_8056);
and U17003 (N_17003,N_8675,N_6873);
and U17004 (N_17004,N_9055,N_11272);
or U17005 (N_17005,N_11494,N_6075);
nand U17006 (N_17006,N_7288,N_7148);
and U17007 (N_17007,N_10157,N_7499);
nor U17008 (N_17008,N_6037,N_7676);
nor U17009 (N_17009,N_7245,N_10217);
xor U17010 (N_17010,N_7423,N_10167);
nor U17011 (N_17011,N_6724,N_11245);
and U17012 (N_17012,N_7376,N_9146);
or U17013 (N_17013,N_11614,N_6753);
nor U17014 (N_17014,N_8692,N_9922);
nand U17015 (N_17015,N_10847,N_9441);
nand U17016 (N_17016,N_10240,N_9452);
or U17017 (N_17017,N_9273,N_6552);
nor U17018 (N_17018,N_10301,N_9667);
nand U17019 (N_17019,N_10593,N_11318);
and U17020 (N_17020,N_11328,N_11002);
nor U17021 (N_17021,N_7906,N_7542);
and U17022 (N_17022,N_10244,N_11978);
or U17023 (N_17023,N_7986,N_7079);
or U17024 (N_17024,N_8247,N_7258);
and U17025 (N_17025,N_10680,N_10959);
nand U17026 (N_17026,N_6844,N_9471);
or U17027 (N_17027,N_8195,N_6729);
nand U17028 (N_17028,N_9948,N_6197);
nand U17029 (N_17029,N_7896,N_11818);
and U17030 (N_17030,N_9896,N_8804);
nand U17031 (N_17031,N_7214,N_9905);
nand U17032 (N_17032,N_9672,N_10993);
or U17033 (N_17033,N_11816,N_10251);
and U17034 (N_17034,N_10421,N_7452);
xor U17035 (N_17035,N_6224,N_9738);
and U17036 (N_17036,N_6076,N_10726);
or U17037 (N_17037,N_11502,N_11481);
or U17038 (N_17038,N_10879,N_6209);
nand U17039 (N_17039,N_6090,N_10910);
or U17040 (N_17040,N_6631,N_8178);
and U17041 (N_17041,N_9738,N_11068);
or U17042 (N_17042,N_10361,N_9555);
or U17043 (N_17043,N_8171,N_9376);
nor U17044 (N_17044,N_11326,N_7300);
or U17045 (N_17045,N_11593,N_6083);
nand U17046 (N_17046,N_8259,N_7435);
nor U17047 (N_17047,N_8117,N_6164);
nor U17048 (N_17048,N_10132,N_11965);
nor U17049 (N_17049,N_10872,N_8103);
nor U17050 (N_17050,N_9314,N_11414);
nor U17051 (N_17051,N_7503,N_10629);
or U17052 (N_17052,N_8293,N_10341);
and U17053 (N_17053,N_9795,N_10951);
nand U17054 (N_17054,N_11828,N_9817);
xor U17055 (N_17055,N_6272,N_11810);
nand U17056 (N_17056,N_9531,N_9701);
nor U17057 (N_17057,N_9807,N_6071);
or U17058 (N_17058,N_8181,N_11135);
or U17059 (N_17059,N_11657,N_7157);
xor U17060 (N_17060,N_9565,N_6735);
nand U17061 (N_17061,N_10983,N_8371);
xnor U17062 (N_17062,N_7367,N_7514);
nand U17063 (N_17063,N_11024,N_11986);
nand U17064 (N_17064,N_7690,N_10349);
or U17065 (N_17065,N_11497,N_11209);
and U17066 (N_17066,N_7619,N_10767);
nor U17067 (N_17067,N_10767,N_10666);
xnor U17068 (N_17068,N_11896,N_8481);
and U17069 (N_17069,N_11678,N_6082);
nand U17070 (N_17070,N_11184,N_7870);
nand U17071 (N_17071,N_9187,N_6967);
nor U17072 (N_17072,N_10248,N_6438);
xor U17073 (N_17073,N_7397,N_11509);
nand U17074 (N_17074,N_7341,N_10191);
nor U17075 (N_17075,N_6540,N_7896);
nand U17076 (N_17076,N_7850,N_11463);
nor U17077 (N_17077,N_7417,N_6230);
and U17078 (N_17078,N_11191,N_8423);
or U17079 (N_17079,N_7770,N_7577);
nor U17080 (N_17080,N_6184,N_10438);
and U17081 (N_17081,N_7928,N_7041);
or U17082 (N_17082,N_10573,N_11873);
and U17083 (N_17083,N_7664,N_9329);
and U17084 (N_17084,N_9004,N_10356);
xnor U17085 (N_17085,N_8880,N_11812);
and U17086 (N_17086,N_11626,N_7044);
and U17087 (N_17087,N_11424,N_7435);
nor U17088 (N_17088,N_6875,N_6891);
xnor U17089 (N_17089,N_8396,N_8475);
or U17090 (N_17090,N_10828,N_9368);
nand U17091 (N_17091,N_8675,N_11784);
and U17092 (N_17092,N_8994,N_10382);
nor U17093 (N_17093,N_7711,N_6363);
xnor U17094 (N_17094,N_8138,N_7809);
and U17095 (N_17095,N_11140,N_7859);
nand U17096 (N_17096,N_8714,N_11451);
and U17097 (N_17097,N_11281,N_9873);
nand U17098 (N_17098,N_10396,N_8515);
and U17099 (N_17099,N_7869,N_6781);
or U17100 (N_17100,N_8680,N_6676);
nand U17101 (N_17101,N_7839,N_8533);
and U17102 (N_17102,N_9066,N_10696);
and U17103 (N_17103,N_8501,N_6082);
nor U17104 (N_17104,N_9888,N_9632);
and U17105 (N_17105,N_8359,N_6808);
and U17106 (N_17106,N_7111,N_8208);
nand U17107 (N_17107,N_9662,N_8020);
and U17108 (N_17108,N_11477,N_10398);
xnor U17109 (N_17109,N_9332,N_6328);
and U17110 (N_17110,N_11020,N_8924);
or U17111 (N_17111,N_6368,N_7121);
nand U17112 (N_17112,N_6634,N_9440);
nand U17113 (N_17113,N_8763,N_8528);
and U17114 (N_17114,N_10931,N_7711);
nor U17115 (N_17115,N_10401,N_11849);
xor U17116 (N_17116,N_9641,N_9114);
or U17117 (N_17117,N_9308,N_11228);
and U17118 (N_17118,N_6954,N_6556);
xor U17119 (N_17119,N_8356,N_10878);
nor U17120 (N_17120,N_8001,N_10101);
xor U17121 (N_17121,N_8166,N_10226);
or U17122 (N_17122,N_8294,N_6546);
and U17123 (N_17123,N_9241,N_11194);
and U17124 (N_17124,N_6335,N_9661);
nor U17125 (N_17125,N_8737,N_10409);
or U17126 (N_17126,N_11449,N_9571);
and U17127 (N_17127,N_9885,N_7997);
xor U17128 (N_17128,N_9055,N_6345);
and U17129 (N_17129,N_11285,N_6109);
nor U17130 (N_17130,N_11876,N_7358);
or U17131 (N_17131,N_7166,N_8905);
nor U17132 (N_17132,N_7224,N_7001);
xnor U17133 (N_17133,N_10518,N_7847);
nand U17134 (N_17134,N_7430,N_9221);
nand U17135 (N_17135,N_7047,N_6011);
xnor U17136 (N_17136,N_9647,N_10780);
nand U17137 (N_17137,N_6707,N_10770);
and U17138 (N_17138,N_7517,N_8764);
and U17139 (N_17139,N_7938,N_8219);
nand U17140 (N_17140,N_7470,N_11554);
nand U17141 (N_17141,N_9125,N_10388);
nor U17142 (N_17142,N_8445,N_9567);
xor U17143 (N_17143,N_6021,N_7831);
or U17144 (N_17144,N_10598,N_11101);
or U17145 (N_17145,N_11335,N_6080);
nor U17146 (N_17146,N_6903,N_10263);
and U17147 (N_17147,N_7491,N_10491);
nand U17148 (N_17148,N_7386,N_10834);
or U17149 (N_17149,N_9281,N_6358);
or U17150 (N_17150,N_11873,N_8152);
nand U17151 (N_17151,N_8375,N_11734);
nor U17152 (N_17152,N_7276,N_11978);
and U17153 (N_17153,N_10584,N_8444);
and U17154 (N_17154,N_9624,N_6669);
xnor U17155 (N_17155,N_11784,N_6794);
and U17156 (N_17156,N_9367,N_10388);
or U17157 (N_17157,N_11199,N_11685);
xor U17158 (N_17158,N_6437,N_11494);
xnor U17159 (N_17159,N_7965,N_9415);
nand U17160 (N_17160,N_9149,N_9432);
nor U17161 (N_17161,N_9698,N_6896);
nor U17162 (N_17162,N_6980,N_11559);
and U17163 (N_17163,N_9024,N_8424);
or U17164 (N_17164,N_8947,N_9725);
or U17165 (N_17165,N_7530,N_7080);
nor U17166 (N_17166,N_7253,N_10998);
and U17167 (N_17167,N_6453,N_7212);
nand U17168 (N_17168,N_10977,N_7235);
and U17169 (N_17169,N_6080,N_8019);
or U17170 (N_17170,N_6743,N_11919);
and U17171 (N_17171,N_9107,N_10824);
nor U17172 (N_17172,N_9957,N_7992);
nand U17173 (N_17173,N_11679,N_7021);
or U17174 (N_17174,N_10529,N_11930);
or U17175 (N_17175,N_11922,N_6492);
or U17176 (N_17176,N_7087,N_7193);
nor U17177 (N_17177,N_10200,N_7645);
or U17178 (N_17178,N_9269,N_11335);
nand U17179 (N_17179,N_10243,N_9597);
xnor U17180 (N_17180,N_6983,N_7043);
nor U17181 (N_17181,N_8915,N_6780);
nand U17182 (N_17182,N_10099,N_10472);
nor U17183 (N_17183,N_6634,N_11869);
nand U17184 (N_17184,N_11888,N_9010);
nand U17185 (N_17185,N_10459,N_6413);
and U17186 (N_17186,N_7864,N_8068);
nand U17187 (N_17187,N_10330,N_8644);
and U17188 (N_17188,N_10472,N_10244);
nand U17189 (N_17189,N_7609,N_11447);
xnor U17190 (N_17190,N_11555,N_9955);
or U17191 (N_17191,N_10591,N_8016);
or U17192 (N_17192,N_9075,N_10634);
nand U17193 (N_17193,N_9269,N_11039);
and U17194 (N_17194,N_7846,N_9586);
nand U17195 (N_17195,N_10001,N_7798);
or U17196 (N_17196,N_7707,N_7563);
nand U17197 (N_17197,N_9939,N_6423);
or U17198 (N_17198,N_7097,N_8379);
nor U17199 (N_17199,N_9152,N_7311);
or U17200 (N_17200,N_11750,N_6188);
or U17201 (N_17201,N_9062,N_9647);
or U17202 (N_17202,N_10912,N_10269);
and U17203 (N_17203,N_9442,N_6155);
or U17204 (N_17204,N_7128,N_6594);
or U17205 (N_17205,N_8133,N_7429);
or U17206 (N_17206,N_11424,N_11435);
and U17207 (N_17207,N_8796,N_10136);
or U17208 (N_17208,N_8061,N_11605);
and U17209 (N_17209,N_7483,N_10992);
xor U17210 (N_17210,N_8874,N_9015);
and U17211 (N_17211,N_10205,N_9766);
nor U17212 (N_17212,N_8804,N_9663);
and U17213 (N_17213,N_9389,N_8460);
or U17214 (N_17214,N_9217,N_8974);
or U17215 (N_17215,N_10640,N_6976);
or U17216 (N_17216,N_8094,N_11317);
or U17217 (N_17217,N_8003,N_10869);
and U17218 (N_17218,N_10088,N_10431);
nand U17219 (N_17219,N_9890,N_9609);
nor U17220 (N_17220,N_8297,N_8153);
or U17221 (N_17221,N_6724,N_9306);
nor U17222 (N_17222,N_8571,N_10049);
xnor U17223 (N_17223,N_10191,N_9024);
nor U17224 (N_17224,N_7345,N_6805);
xnor U17225 (N_17225,N_11047,N_9024);
xnor U17226 (N_17226,N_11401,N_8897);
and U17227 (N_17227,N_10321,N_11531);
or U17228 (N_17228,N_9085,N_10318);
nand U17229 (N_17229,N_7806,N_6024);
nor U17230 (N_17230,N_11214,N_8136);
nand U17231 (N_17231,N_9096,N_9557);
or U17232 (N_17232,N_6124,N_9019);
nand U17233 (N_17233,N_9235,N_9831);
and U17234 (N_17234,N_9523,N_11458);
and U17235 (N_17235,N_8132,N_8987);
and U17236 (N_17236,N_11290,N_11996);
or U17237 (N_17237,N_10157,N_11880);
xnor U17238 (N_17238,N_9301,N_10248);
nor U17239 (N_17239,N_8779,N_11977);
nor U17240 (N_17240,N_6482,N_8007);
or U17241 (N_17241,N_11251,N_9257);
and U17242 (N_17242,N_8743,N_8262);
nor U17243 (N_17243,N_8810,N_8282);
nor U17244 (N_17244,N_7867,N_10623);
and U17245 (N_17245,N_7359,N_9597);
or U17246 (N_17246,N_9161,N_7589);
or U17247 (N_17247,N_10426,N_9586);
xor U17248 (N_17248,N_6902,N_8134);
nand U17249 (N_17249,N_10890,N_11060);
or U17250 (N_17250,N_8897,N_6295);
and U17251 (N_17251,N_6701,N_9802);
and U17252 (N_17252,N_9813,N_10608);
or U17253 (N_17253,N_6682,N_11616);
nor U17254 (N_17254,N_8430,N_8092);
or U17255 (N_17255,N_7650,N_7338);
xnor U17256 (N_17256,N_10473,N_10651);
nor U17257 (N_17257,N_8423,N_6958);
nand U17258 (N_17258,N_10528,N_10379);
nand U17259 (N_17259,N_11697,N_8095);
or U17260 (N_17260,N_9084,N_10572);
nand U17261 (N_17261,N_7202,N_7568);
nor U17262 (N_17262,N_8018,N_11445);
nand U17263 (N_17263,N_11451,N_8787);
nor U17264 (N_17264,N_8309,N_9285);
or U17265 (N_17265,N_7757,N_10037);
nor U17266 (N_17266,N_8526,N_6303);
or U17267 (N_17267,N_9464,N_11616);
nor U17268 (N_17268,N_7367,N_7120);
and U17269 (N_17269,N_9194,N_7476);
nor U17270 (N_17270,N_10435,N_7331);
nor U17271 (N_17271,N_7019,N_11836);
nand U17272 (N_17272,N_6194,N_10012);
nor U17273 (N_17273,N_10715,N_9188);
nand U17274 (N_17274,N_11603,N_8272);
or U17275 (N_17275,N_11502,N_10280);
or U17276 (N_17276,N_8523,N_9894);
nand U17277 (N_17277,N_10941,N_7905);
xnor U17278 (N_17278,N_10793,N_9383);
or U17279 (N_17279,N_11549,N_11724);
xor U17280 (N_17280,N_6717,N_9943);
nand U17281 (N_17281,N_11230,N_8550);
nor U17282 (N_17282,N_7769,N_10184);
nand U17283 (N_17283,N_10369,N_6113);
nand U17284 (N_17284,N_11485,N_9749);
nand U17285 (N_17285,N_9760,N_11396);
xnor U17286 (N_17286,N_11884,N_7329);
or U17287 (N_17287,N_9767,N_10118);
nand U17288 (N_17288,N_9505,N_8039);
and U17289 (N_17289,N_11630,N_9298);
nor U17290 (N_17290,N_11850,N_8303);
and U17291 (N_17291,N_9442,N_9662);
nand U17292 (N_17292,N_9469,N_7309);
or U17293 (N_17293,N_6649,N_8571);
or U17294 (N_17294,N_11466,N_7895);
xor U17295 (N_17295,N_7122,N_8225);
xnor U17296 (N_17296,N_11244,N_8157);
or U17297 (N_17297,N_9955,N_11953);
xnor U17298 (N_17298,N_6160,N_9809);
xor U17299 (N_17299,N_7234,N_8560);
and U17300 (N_17300,N_7462,N_10589);
xnor U17301 (N_17301,N_6233,N_9809);
nand U17302 (N_17302,N_9972,N_9271);
or U17303 (N_17303,N_6403,N_10703);
nand U17304 (N_17304,N_11747,N_11015);
xnor U17305 (N_17305,N_10649,N_8285);
or U17306 (N_17306,N_6808,N_7144);
nor U17307 (N_17307,N_7996,N_7201);
nor U17308 (N_17308,N_11594,N_11330);
nand U17309 (N_17309,N_7104,N_7375);
nor U17310 (N_17310,N_6906,N_6615);
or U17311 (N_17311,N_8765,N_11951);
nand U17312 (N_17312,N_8011,N_6759);
nand U17313 (N_17313,N_8423,N_11284);
xor U17314 (N_17314,N_11011,N_11024);
or U17315 (N_17315,N_8755,N_9790);
nand U17316 (N_17316,N_9997,N_10572);
nor U17317 (N_17317,N_11582,N_8387);
nor U17318 (N_17318,N_11384,N_10736);
nor U17319 (N_17319,N_7073,N_6301);
nor U17320 (N_17320,N_10053,N_8460);
or U17321 (N_17321,N_6440,N_11231);
nor U17322 (N_17322,N_7326,N_10325);
or U17323 (N_17323,N_11216,N_6784);
nand U17324 (N_17324,N_6939,N_11653);
and U17325 (N_17325,N_10703,N_8785);
nand U17326 (N_17326,N_11344,N_11408);
or U17327 (N_17327,N_10381,N_9615);
nand U17328 (N_17328,N_6706,N_6411);
or U17329 (N_17329,N_8502,N_6240);
nand U17330 (N_17330,N_8304,N_6249);
and U17331 (N_17331,N_7573,N_6118);
or U17332 (N_17332,N_7254,N_8009);
xnor U17333 (N_17333,N_11502,N_9724);
nand U17334 (N_17334,N_11614,N_8794);
nand U17335 (N_17335,N_10522,N_10098);
and U17336 (N_17336,N_6021,N_10102);
nor U17337 (N_17337,N_9749,N_10724);
nor U17338 (N_17338,N_7457,N_7802);
nor U17339 (N_17339,N_9177,N_9164);
or U17340 (N_17340,N_10277,N_6167);
and U17341 (N_17341,N_6783,N_6435);
nand U17342 (N_17342,N_6205,N_9994);
and U17343 (N_17343,N_8863,N_11982);
nand U17344 (N_17344,N_11000,N_11966);
nand U17345 (N_17345,N_10794,N_7922);
or U17346 (N_17346,N_7797,N_8449);
and U17347 (N_17347,N_11230,N_11232);
and U17348 (N_17348,N_7427,N_11730);
and U17349 (N_17349,N_11029,N_11838);
or U17350 (N_17350,N_6731,N_6704);
or U17351 (N_17351,N_8468,N_8661);
xnor U17352 (N_17352,N_11039,N_8868);
nor U17353 (N_17353,N_10724,N_9608);
and U17354 (N_17354,N_8979,N_11132);
or U17355 (N_17355,N_9847,N_7339);
nand U17356 (N_17356,N_10205,N_9908);
and U17357 (N_17357,N_9129,N_6161);
and U17358 (N_17358,N_11558,N_6980);
and U17359 (N_17359,N_9966,N_6552);
nor U17360 (N_17360,N_7623,N_9012);
and U17361 (N_17361,N_7965,N_8748);
nand U17362 (N_17362,N_8702,N_11204);
nor U17363 (N_17363,N_9646,N_8339);
nor U17364 (N_17364,N_8633,N_6386);
nor U17365 (N_17365,N_9619,N_8435);
xnor U17366 (N_17366,N_11252,N_9163);
nor U17367 (N_17367,N_7582,N_11260);
nor U17368 (N_17368,N_8017,N_7835);
nand U17369 (N_17369,N_7115,N_10812);
nand U17370 (N_17370,N_11437,N_6203);
nor U17371 (N_17371,N_11431,N_10290);
or U17372 (N_17372,N_11413,N_7654);
or U17373 (N_17373,N_11982,N_11769);
and U17374 (N_17374,N_11345,N_8355);
or U17375 (N_17375,N_7943,N_10927);
xnor U17376 (N_17376,N_11811,N_6772);
and U17377 (N_17377,N_9659,N_7965);
or U17378 (N_17378,N_9140,N_10117);
or U17379 (N_17379,N_11997,N_10007);
nor U17380 (N_17380,N_9402,N_7667);
xnor U17381 (N_17381,N_11076,N_9009);
and U17382 (N_17382,N_11046,N_11030);
or U17383 (N_17383,N_11530,N_7348);
or U17384 (N_17384,N_6041,N_11108);
or U17385 (N_17385,N_10275,N_11775);
and U17386 (N_17386,N_8202,N_8366);
and U17387 (N_17387,N_7953,N_9443);
and U17388 (N_17388,N_11725,N_6809);
nor U17389 (N_17389,N_7629,N_8077);
nor U17390 (N_17390,N_7299,N_10799);
and U17391 (N_17391,N_7458,N_7256);
or U17392 (N_17392,N_9246,N_11848);
or U17393 (N_17393,N_6227,N_8577);
xnor U17394 (N_17394,N_6800,N_8685);
and U17395 (N_17395,N_10349,N_6900);
and U17396 (N_17396,N_10139,N_8176);
xor U17397 (N_17397,N_7675,N_11618);
xor U17398 (N_17398,N_10459,N_10364);
nor U17399 (N_17399,N_11136,N_11472);
nor U17400 (N_17400,N_10294,N_9557);
and U17401 (N_17401,N_7316,N_10516);
or U17402 (N_17402,N_11286,N_8649);
nand U17403 (N_17403,N_10019,N_10091);
nand U17404 (N_17404,N_8195,N_7960);
xnor U17405 (N_17405,N_11086,N_10440);
nand U17406 (N_17406,N_10199,N_10695);
and U17407 (N_17407,N_6289,N_6252);
nand U17408 (N_17408,N_9887,N_8163);
xnor U17409 (N_17409,N_6264,N_11664);
or U17410 (N_17410,N_11638,N_10249);
xnor U17411 (N_17411,N_10611,N_9684);
xor U17412 (N_17412,N_8799,N_9301);
nor U17413 (N_17413,N_11716,N_9163);
and U17414 (N_17414,N_7686,N_6049);
nor U17415 (N_17415,N_7320,N_10599);
nand U17416 (N_17416,N_11027,N_10275);
xor U17417 (N_17417,N_10570,N_6546);
and U17418 (N_17418,N_10586,N_6805);
nor U17419 (N_17419,N_11273,N_11328);
nor U17420 (N_17420,N_9882,N_10636);
xnor U17421 (N_17421,N_8993,N_6324);
or U17422 (N_17422,N_7321,N_11221);
or U17423 (N_17423,N_10395,N_10537);
or U17424 (N_17424,N_9787,N_7506);
or U17425 (N_17425,N_11485,N_7855);
or U17426 (N_17426,N_6449,N_11777);
and U17427 (N_17427,N_11751,N_7714);
xor U17428 (N_17428,N_9453,N_8651);
nor U17429 (N_17429,N_10102,N_11984);
and U17430 (N_17430,N_10066,N_9403);
nand U17431 (N_17431,N_9887,N_6110);
nand U17432 (N_17432,N_9955,N_9823);
and U17433 (N_17433,N_11557,N_11337);
or U17434 (N_17434,N_11603,N_11019);
and U17435 (N_17435,N_8663,N_11157);
nand U17436 (N_17436,N_10482,N_11601);
nand U17437 (N_17437,N_9233,N_7814);
or U17438 (N_17438,N_8235,N_6975);
and U17439 (N_17439,N_6856,N_9637);
or U17440 (N_17440,N_9759,N_11762);
or U17441 (N_17441,N_11687,N_9920);
xnor U17442 (N_17442,N_8617,N_7451);
nor U17443 (N_17443,N_11329,N_7608);
and U17444 (N_17444,N_7481,N_6071);
and U17445 (N_17445,N_8677,N_11180);
or U17446 (N_17446,N_11671,N_11025);
nor U17447 (N_17447,N_9421,N_9883);
or U17448 (N_17448,N_10624,N_11948);
nor U17449 (N_17449,N_6371,N_10503);
and U17450 (N_17450,N_6652,N_11140);
nor U17451 (N_17451,N_9458,N_11184);
nor U17452 (N_17452,N_6917,N_7437);
or U17453 (N_17453,N_7927,N_9690);
or U17454 (N_17454,N_6748,N_8829);
nand U17455 (N_17455,N_7477,N_11272);
or U17456 (N_17456,N_6518,N_6534);
xor U17457 (N_17457,N_7631,N_6716);
or U17458 (N_17458,N_6968,N_8229);
nand U17459 (N_17459,N_11346,N_6259);
or U17460 (N_17460,N_8055,N_8863);
nand U17461 (N_17461,N_8860,N_10272);
or U17462 (N_17462,N_10822,N_6309);
nor U17463 (N_17463,N_7472,N_8982);
nand U17464 (N_17464,N_11539,N_8552);
xor U17465 (N_17465,N_11254,N_8400);
nor U17466 (N_17466,N_11977,N_6911);
nand U17467 (N_17467,N_9748,N_8459);
nand U17468 (N_17468,N_11767,N_10668);
nor U17469 (N_17469,N_10848,N_9337);
nor U17470 (N_17470,N_10187,N_11651);
nand U17471 (N_17471,N_10951,N_11179);
xnor U17472 (N_17472,N_11200,N_7304);
or U17473 (N_17473,N_9923,N_10313);
or U17474 (N_17474,N_9645,N_10465);
xnor U17475 (N_17475,N_9785,N_6668);
or U17476 (N_17476,N_7269,N_10163);
and U17477 (N_17477,N_8527,N_9179);
and U17478 (N_17478,N_10150,N_11839);
nor U17479 (N_17479,N_8307,N_7330);
or U17480 (N_17480,N_6945,N_10744);
or U17481 (N_17481,N_10087,N_11221);
nand U17482 (N_17482,N_6643,N_7382);
xor U17483 (N_17483,N_6282,N_6092);
xnor U17484 (N_17484,N_11014,N_8209);
nand U17485 (N_17485,N_9573,N_10409);
xor U17486 (N_17486,N_10774,N_6804);
nand U17487 (N_17487,N_11715,N_6411);
xnor U17488 (N_17488,N_7615,N_6725);
nor U17489 (N_17489,N_6736,N_6314);
and U17490 (N_17490,N_7145,N_11498);
nand U17491 (N_17491,N_6130,N_8561);
or U17492 (N_17492,N_8080,N_9419);
or U17493 (N_17493,N_6349,N_11175);
and U17494 (N_17494,N_7120,N_6085);
nor U17495 (N_17495,N_10592,N_8556);
and U17496 (N_17496,N_11991,N_9194);
and U17497 (N_17497,N_9863,N_6304);
or U17498 (N_17498,N_7289,N_9757);
nor U17499 (N_17499,N_10183,N_9361);
and U17500 (N_17500,N_7824,N_9261);
and U17501 (N_17501,N_11507,N_8836);
xor U17502 (N_17502,N_8421,N_11402);
and U17503 (N_17503,N_8605,N_7127);
and U17504 (N_17504,N_6770,N_6903);
and U17505 (N_17505,N_9709,N_8448);
nand U17506 (N_17506,N_7409,N_6447);
or U17507 (N_17507,N_9966,N_9114);
nor U17508 (N_17508,N_11639,N_10680);
nand U17509 (N_17509,N_7806,N_6528);
and U17510 (N_17510,N_6105,N_11966);
nor U17511 (N_17511,N_9574,N_11826);
nor U17512 (N_17512,N_8113,N_11127);
and U17513 (N_17513,N_11556,N_8351);
nor U17514 (N_17514,N_9775,N_9730);
or U17515 (N_17515,N_8257,N_8903);
nor U17516 (N_17516,N_9501,N_11095);
and U17517 (N_17517,N_11036,N_11804);
nand U17518 (N_17518,N_7950,N_11131);
nand U17519 (N_17519,N_9417,N_6016);
nand U17520 (N_17520,N_6688,N_11605);
and U17521 (N_17521,N_8021,N_9037);
nor U17522 (N_17522,N_9298,N_10954);
xor U17523 (N_17523,N_10793,N_6694);
and U17524 (N_17524,N_11197,N_6943);
nand U17525 (N_17525,N_10215,N_8093);
nor U17526 (N_17526,N_9186,N_7399);
xor U17527 (N_17527,N_6647,N_8389);
xnor U17528 (N_17528,N_9233,N_11211);
nand U17529 (N_17529,N_11392,N_10933);
and U17530 (N_17530,N_9110,N_9846);
nor U17531 (N_17531,N_6465,N_10771);
and U17532 (N_17532,N_9441,N_6593);
nor U17533 (N_17533,N_10395,N_11942);
xor U17534 (N_17534,N_6636,N_10398);
xnor U17535 (N_17535,N_10509,N_7650);
nand U17536 (N_17536,N_8397,N_9125);
or U17537 (N_17537,N_10750,N_10304);
or U17538 (N_17538,N_10043,N_6324);
nand U17539 (N_17539,N_10955,N_10945);
nor U17540 (N_17540,N_9699,N_6983);
nor U17541 (N_17541,N_10846,N_7636);
or U17542 (N_17542,N_7077,N_8026);
or U17543 (N_17543,N_10989,N_11741);
nand U17544 (N_17544,N_7427,N_8130);
xnor U17545 (N_17545,N_10382,N_9193);
xnor U17546 (N_17546,N_8019,N_6418);
xnor U17547 (N_17547,N_6443,N_8401);
or U17548 (N_17548,N_8254,N_10208);
nand U17549 (N_17549,N_7807,N_7141);
xor U17550 (N_17550,N_9303,N_11694);
and U17551 (N_17551,N_11303,N_11793);
xor U17552 (N_17552,N_6830,N_9504);
xor U17553 (N_17553,N_10784,N_8747);
nor U17554 (N_17554,N_8592,N_10759);
nand U17555 (N_17555,N_11644,N_7394);
nor U17556 (N_17556,N_7106,N_9521);
or U17557 (N_17557,N_11740,N_8743);
nor U17558 (N_17558,N_8818,N_7800);
or U17559 (N_17559,N_10136,N_8377);
or U17560 (N_17560,N_10082,N_8046);
nand U17561 (N_17561,N_7253,N_8184);
and U17562 (N_17562,N_11974,N_7942);
or U17563 (N_17563,N_10374,N_10468);
and U17564 (N_17564,N_8114,N_6894);
or U17565 (N_17565,N_10282,N_8588);
nor U17566 (N_17566,N_9277,N_11563);
or U17567 (N_17567,N_10058,N_6211);
xor U17568 (N_17568,N_7464,N_11292);
or U17569 (N_17569,N_10908,N_9639);
xnor U17570 (N_17570,N_11416,N_9854);
nand U17571 (N_17571,N_11969,N_9675);
and U17572 (N_17572,N_7457,N_11625);
nand U17573 (N_17573,N_7557,N_9517);
and U17574 (N_17574,N_11484,N_6114);
nor U17575 (N_17575,N_8375,N_9050);
or U17576 (N_17576,N_10861,N_10033);
nand U17577 (N_17577,N_10907,N_11898);
or U17578 (N_17578,N_11639,N_11788);
nand U17579 (N_17579,N_7407,N_10243);
or U17580 (N_17580,N_9452,N_6211);
nor U17581 (N_17581,N_11133,N_8178);
and U17582 (N_17582,N_7572,N_8389);
nor U17583 (N_17583,N_6250,N_11403);
nand U17584 (N_17584,N_6209,N_10490);
nor U17585 (N_17585,N_8499,N_9505);
nor U17586 (N_17586,N_6430,N_7514);
or U17587 (N_17587,N_8937,N_10570);
xnor U17588 (N_17588,N_9759,N_6036);
nand U17589 (N_17589,N_11785,N_10237);
and U17590 (N_17590,N_11993,N_6584);
and U17591 (N_17591,N_8632,N_9339);
nand U17592 (N_17592,N_7066,N_10744);
or U17593 (N_17593,N_7753,N_6835);
xnor U17594 (N_17594,N_7587,N_8789);
and U17595 (N_17595,N_6154,N_8378);
nand U17596 (N_17596,N_9472,N_11328);
nand U17597 (N_17597,N_10826,N_11214);
nand U17598 (N_17598,N_10893,N_7746);
and U17599 (N_17599,N_10123,N_7803);
nand U17600 (N_17600,N_7325,N_11703);
nand U17601 (N_17601,N_8801,N_11927);
nor U17602 (N_17602,N_9238,N_7087);
xnor U17603 (N_17603,N_10306,N_6147);
nand U17604 (N_17604,N_9689,N_8370);
nand U17605 (N_17605,N_7896,N_6115);
or U17606 (N_17606,N_9425,N_11628);
xor U17607 (N_17607,N_6853,N_7932);
xor U17608 (N_17608,N_11025,N_11057);
nand U17609 (N_17609,N_7825,N_10970);
nor U17610 (N_17610,N_11775,N_6864);
nand U17611 (N_17611,N_8812,N_9824);
nand U17612 (N_17612,N_10796,N_7297);
or U17613 (N_17613,N_11031,N_6906);
nand U17614 (N_17614,N_11165,N_6474);
nor U17615 (N_17615,N_11591,N_8132);
or U17616 (N_17616,N_11418,N_10974);
and U17617 (N_17617,N_7911,N_8853);
and U17618 (N_17618,N_7543,N_10616);
and U17619 (N_17619,N_11660,N_6995);
and U17620 (N_17620,N_11259,N_6549);
xnor U17621 (N_17621,N_8866,N_7107);
and U17622 (N_17622,N_8582,N_7892);
nand U17623 (N_17623,N_8422,N_10901);
and U17624 (N_17624,N_6977,N_11896);
nor U17625 (N_17625,N_8392,N_10393);
nor U17626 (N_17626,N_7970,N_9037);
or U17627 (N_17627,N_8967,N_7656);
nor U17628 (N_17628,N_7357,N_8137);
or U17629 (N_17629,N_10145,N_11365);
xor U17630 (N_17630,N_6502,N_6836);
or U17631 (N_17631,N_10192,N_7243);
nand U17632 (N_17632,N_10136,N_10932);
or U17633 (N_17633,N_8776,N_10280);
and U17634 (N_17634,N_10503,N_6895);
or U17635 (N_17635,N_11463,N_6284);
and U17636 (N_17636,N_11316,N_9447);
and U17637 (N_17637,N_6519,N_10026);
and U17638 (N_17638,N_10218,N_10030);
nor U17639 (N_17639,N_8490,N_9677);
and U17640 (N_17640,N_9004,N_9090);
nand U17641 (N_17641,N_11302,N_9063);
and U17642 (N_17642,N_6794,N_11366);
nor U17643 (N_17643,N_9724,N_8835);
xnor U17644 (N_17644,N_6558,N_7460);
or U17645 (N_17645,N_11760,N_9026);
xor U17646 (N_17646,N_11130,N_7566);
xor U17647 (N_17647,N_10500,N_9408);
or U17648 (N_17648,N_6115,N_8160);
nor U17649 (N_17649,N_9020,N_6439);
and U17650 (N_17650,N_7663,N_8976);
nand U17651 (N_17651,N_6057,N_6688);
xor U17652 (N_17652,N_6812,N_9589);
nand U17653 (N_17653,N_7676,N_10201);
nor U17654 (N_17654,N_11561,N_7053);
nand U17655 (N_17655,N_7614,N_9980);
or U17656 (N_17656,N_6286,N_9782);
or U17657 (N_17657,N_7459,N_6695);
nor U17658 (N_17658,N_10706,N_7553);
nand U17659 (N_17659,N_11191,N_10432);
xnor U17660 (N_17660,N_10524,N_8016);
or U17661 (N_17661,N_8015,N_6697);
nand U17662 (N_17662,N_9060,N_9622);
or U17663 (N_17663,N_8663,N_9635);
nand U17664 (N_17664,N_11481,N_10797);
and U17665 (N_17665,N_8639,N_9541);
nand U17666 (N_17666,N_9153,N_10435);
xor U17667 (N_17667,N_11551,N_9642);
and U17668 (N_17668,N_11176,N_10480);
nand U17669 (N_17669,N_7609,N_9163);
nor U17670 (N_17670,N_11376,N_10552);
nand U17671 (N_17671,N_11197,N_11568);
nand U17672 (N_17672,N_11677,N_8290);
and U17673 (N_17673,N_8945,N_7197);
xnor U17674 (N_17674,N_7711,N_10678);
nor U17675 (N_17675,N_7162,N_10977);
nor U17676 (N_17676,N_10608,N_8641);
or U17677 (N_17677,N_6392,N_6798);
nor U17678 (N_17678,N_6303,N_10909);
or U17679 (N_17679,N_9146,N_7478);
nor U17680 (N_17680,N_10950,N_10152);
nand U17681 (N_17681,N_7725,N_10392);
and U17682 (N_17682,N_9983,N_6229);
or U17683 (N_17683,N_9693,N_9966);
nand U17684 (N_17684,N_11602,N_11667);
or U17685 (N_17685,N_6029,N_6627);
nor U17686 (N_17686,N_8895,N_7823);
xnor U17687 (N_17687,N_11330,N_9311);
xor U17688 (N_17688,N_11348,N_7855);
and U17689 (N_17689,N_9652,N_11067);
or U17690 (N_17690,N_11549,N_9787);
and U17691 (N_17691,N_11187,N_10572);
or U17692 (N_17692,N_11701,N_9647);
nand U17693 (N_17693,N_6330,N_8090);
nor U17694 (N_17694,N_11918,N_6791);
or U17695 (N_17695,N_6842,N_10064);
nand U17696 (N_17696,N_10528,N_10454);
nand U17697 (N_17697,N_9878,N_9105);
nand U17698 (N_17698,N_11040,N_6235);
nor U17699 (N_17699,N_9191,N_8816);
and U17700 (N_17700,N_11497,N_10745);
and U17701 (N_17701,N_7242,N_11576);
or U17702 (N_17702,N_10417,N_6199);
nor U17703 (N_17703,N_9727,N_11288);
or U17704 (N_17704,N_9469,N_7136);
and U17705 (N_17705,N_6158,N_11003);
and U17706 (N_17706,N_10315,N_7351);
xnor U17707 (N_17707,N_6910,N_9466);
nor U17708 (N_17708,N_6762,N_7843);
and U17709 (N_17709,N_8837,N_11467);
nand U17710 (N_17710,N_11618,N_8802);
nor U17711 (N_17711,N_10400,N_10801);
and U17712 (N_17712,N_10755,N_7144);
nor U17713 (N_17713,N_6774,N_9571);
nand U17714 (N_17714,N_8498,N_11517);
and U17715 (N_17715,N_10523,N_11387);
and U17716 (N_17716,N_8611,N_7610);
xor U17717 (N_17717,N_10043,N_11728);
and U17718 (N_17718,N_6634,N_10533);
or U17719 (N_17719,N_10094,N_10182);
and U17720 (N_17720,N_9062,N_11340);
and U17721 (N_17721,N_8114,N_8416);
and U17722 (N_17722,N_7811,N_9367);
and U17723 (N_17723,N_10040,N_10660);
or U17724 (N_17724,N_7703,N_9744);
nor U17725 (N_17725,N_7845,N_11499);
and U17726 (N_17726,N_10031,N_8860);
or U17727 (N_17727,N_11819,N_7653);
xor U17728 (N_17728,N_11421,N_7191);
and U17729 (N_17729,N_6856,N_9579);
nand U17730 (N_17730,N_11126,N_11191);
nor U17731 (N_17731,N_6553,N_10765);
and U17732 (N_17732,N_9996,N_11341);
or U17733 (N_17733,N_9446,N_6738);
and U17734 (N_17734,N_11485,N_10083);
nand U17735 (N_17735,N_6962,N_10958);
or U17736 (N_17736,N_10174,N_11493);
nor U17737 (N_17737,N_7914,N_9343);
or U17738 (N_17738,N_7273,N_9452);
nand U17739 (N_17739,N_10646,N_8635);
and U17740 (N_17740,N_10487,N_7203);
nor U17741 (N_17741,N_11142,N_11125);
and U17742 (N_17742,N_7506,N_9067);
and U17743 (N_17743,N_8281,N_11582);
nand U17744 (N_17744,N_6198,N_11325);
or U17745 (N_17745,N_7502,N_7428);
nor U17746 (N_17746,N_10979,N_7664);
nand U17747 (N_17747,N_7355,N_6395);
and U17748 (N_17748,N_7402,N_6953);
nor U17749 (N_17749,N_10983,N_6936);
or U17750 (N_17750,N_11088,N_7971);
nand U17751 (N_17751,N_6826,N_6342);
or U17752 (N_17752,N_9453,N_11177);
and U17753 (N_17753,N_8341,N_11895);
xor U17754 (N_17754,N_10765,N_11250);
nand U17755 (N_17755,N_10578,N_11276);
and U17756 (N_17756,N_7775,N_6362);
and U17757 (N_17757,N_9376,N_8769);
and U17758 (N_17758,N_11136,N_10806);
nand U17759 (N_17759,N_11363,N_7365);
or U17760 (N_17760,N_8279,N_7792);
nand U17761 (N_17761,N_7445,N_11946);
or U17762 (N_17762,N_7100,N_9981);
and U17763 (N_17763,N_8340,N_6350);
and U17764 (N_17764,N_11205,N_8757);
or U17765 (N_17765,N_7115,N_9024);
xnor U17766 (N_17766,N_8056,N_10616);
xnor U17767 (N_17767,N_7492,N_11635);
nand U17768 (N_17768,N_7151,N_8361);
nand U17769 (N_17769,N_8435,N_11408);
or U17770 (N_17770,N_11681,N_9213);
nor U17771 (N_17771,N_10540,N_7098);
or U17772 (N_17772,N_10477,N_11838);
or U17773 (N_17773,N_6785,N_7914);
nor U17774 (N_17774,N_8423,N_9604);
nand U17775 (N_17775,N_9890,N_6487);
or U17776 (N_17776,N_10666,N_10486);
or U17777 (N_17777,N_7005,N_9328);
xor U17778 (N_17778,N_7462,N_8599);
or U17779 (N_17779,N_11420,N_10168);
nor U17780 (N_17780,N_7936,N_8585);
or U17781 (N_17781,N_7122,N_11345);
xnor U17782 (N_17782,N_9553,N_6315);
or U17783 (N_17783,N_6070,N_10570);
nand U17784 (N_17784,N_6359,N_8892);
or U17785 (N_17785,N_7489,N_7534);
and U17786 (N_17786,N_10476,N_8888);
nand U17787 (N_17787,N_8310,N_9810);
nand U17788 (N_17788,N_10254,N_6201);
nor U17789 (N_17789,N_10685,N_11168);
nor U17790 (N_17790,N_7558,N_6915);
xor U17791 (N_17791,N_11574,N_8508);
xnor U17792 (N_17792,N_6275,N_9636);
nand U17793 (N_17793,N_10509,N_6175);
nand U17794 (N_17794,N_6296,N_9697);
or U17795 (N_17795,N_11995,N_8311);
xnor U17796 (N_17796,N_10127,N_10774);
xnor U17797 (N_17797,N_11918,N_10572);
and U17798 (N_17798,N_9971,N_11877);
or U17799 (N_17799,N_6922,N_9671);
nor U17800 (N_17800,N_7537,N_9107);
or U17801 (N_17801,N_10075,N_9794);
or U17802 (N_17802,N_6070,N_8303);
and U17803 (N_17803,N_8941,N_10822);
or U17804 (N_17804,N_10072,N_11091);
or U17805 (N_17805,N_8775,N_10405);
nor U17806 (N_17806,N_8284,N_6182);
nor U17807 (N_17807,N_6431,N_7175);
nor U17808 (N_17808,N_6135,N_8314);
and U17809 (N_17809,N_10616,N_10411);
and U17810 (N_17810,N_10343,N_6725);
nor U17811 (N_17811,N_9930,N_8593);
or U17812 (N_17812,N_8235,N_7917);
and U17813 (N_17813,N_8387,N_8840);
nor U17814 (N_17814,N_9999,N_7135);
and U17815 (N_17815,N_10266,N_11390);
and U17816 (N_17816,N_9180,N_7720);
or U17817 (N_17817,N_8755,N_6928);
xnor U17818 (N_17818,N_11644,N_6996);
or U17819 (N_17819,N_11797,N_8389);
nand U17820 (N_17820,N_8677,N_10491);
and U17821 (N_17821,N_10969,N_10550);
and U17822 (N_17822,N_11990,N_11763);
nor U17823 (N_17823,N_10769,N_10577);
nand U17824 (N_17824,N_6695,N_7181);
or U17825 (N_17825,N_6835,N_8202);
and U17826 (N_17826,N_11095,N_8299);
xnor U17827 (N_17827,N_10019,N_9265);
and U17828 (N_17828,N_10784,N_11591);
nand U17829 (N_17829,N_8532,N_6014);
nor U17830 (N_17830,N_6938,N_8084);
or U17831 (N_17831,N_7635,N_9321);
or U17832 (N_17832,N_7897,N_6216);
nor U17833 (N_17833,N_11939,N_11922);
nor U17834 (N_17834,N_7207,N_7063);
nand U17835 (N_17835,N_10058,N_9151);
or U17836 (N_17836,N_6364,N_9109);
and U17837 (N_17837,N_6031,N_6684);
nor U17838 (N_17838,N_6529,N_7244);
nor U17839 (N_17839,N_9959,N_11825);
nand U17840 (N_17840,N_6208,N_8562);
xnor U17841 (N_17841,N_10138,N_10769);
nor U17842 (N_17842,N_9336,N_6853);
nand U17843 (N_17843,N_6363,N_9986);
and U17844 (N_17844,N_7822,N_9067);
xor U17845 (N_17845,N_11985,N_7693);
or U17846 (N_17846,N_11788,N_11687);
and U17847 (N_17847,N_8782,N_7444);
or U17848 (N_17848,N_8291,N_8777);
nand U17849 (N_17849,N_9540,N_6856);
or U17850 (N_17850,N_6259,N_10383);
and U17851 (N_17851,N_11245,N_10662);
or U17852 (N_17852,N_11701,N_9576);
or U17853 (N_17853,N_7008,N_8714);
or U17854 (N_17854,N_9930,N_10826);
xor U17855 (N_17855,N_6848,N_7525);
nand U17856 (N_17856,N_7188,N_8021);
or U17857 (N_17857,N_10626,N_9673);
or U17858 (N_17858,N_7907,N_11104);
nand U17859 (N_17859,N_6779,N_7340);
or U17860 (N_17860,N_9704,N_9342);
nand U17861 (N_17861,N_7484,N_11364);
and U17862 (N_17862,N_9031,N_8743);
nand U17863 (N_17863,N_10325,N_10861);
nand U17864 (N_17864,N_10843,N_8822);
nor U17865 (N_17865,N_11788,N_7029);
nor U17866 (N_17866,N_6546,N_11697);
nor U17867 (N_17867,N_9147,N_10602);
nand U17868 (N_17868,N_7287,N_6768);
or U17869 (N_17869,N_9466,N_7943);
nor U17870 (N_17870,N_6347,N_6999);
or U17871 (N_17871,N_8194,N_7838);
xor U17872 (N_17872,N_6193,N_8037);
and U17873 (N_17873,N_10000,N_9432);
nand U17874 (N_17874,N_9646,N_10786);
and U17875 (N_17875,N_7032,N_7871);
or U17876 (N_17876,N_9904,N_9091);
xor U17877 (N_17877,N_9666,N_7356);
xor U17878 (N_17878,N_10649,N_8380);
nor U17879 (N_17879,N_7838,N_8121);
nand U17880 (N_17880,N_9042,N_7322);
and U17881 (N_17881,N_9752,N_6001);
nor U17882 (N_17882,N_10471,N_10397);
nor U17883 (N_17883,N_7138,N_7139);
nor U17884 (N_17884,N_10495,N_10662);
or U17885 (N_17885,N_9248,N_9312);
and U17886 (N_17886,N_10039,N_11960);
nand U17887 (N_17887,N_11922,N_6006);
and U17888 (N_17888,N_10993,N_10187);
nand U17889 (N_17889,N_8178,N_9472);
xnor U17890 (N_17890,N_8797,N_11432);
and U17891 (N_17891,N_8146,N_6814);
and U17892 (N_17892,N_7688,N_10813);
nor U17893 (N_17893,N_7888,N_8959);
nand U17894 (N_17894,N_10737,N_10276);
xor U17895 (N_17895,N_9945,N_10444);
nand U17896 (N_17896,N_9887,N_10827);
and U17897 (N_17897,N_9992,N_11403);
nor U17898 (N_17898,N_11471,N_8024);
nand U17899 (N_17899,N_10296,N_8544);
nor U17900 (N_17900,N_11978,N_11550);
or U17901 (N_17901,N_8665,N_6108);
nor U17902 (N_17902,N_10440,N_10410);
nor U17903 (N_17903,N_10141,N_9825);
and U17904 (N_17904,N_11215,N_9071);
nand U17905 (N_17905,N_11495,N_6787);
nand U17906 (N_17906,N_9765,N_11358);
nand U17907 (N_17907,N_10709,N_11779);
xnor U17908 (N_17908,N_7224,N_11549);
and U17909 (N_17909,N_8914,N_6700);
or U17910 (N_17910,N_6068,N_6673);
xnor U17911 (N_17911,N_9571,N_9462);
nor U17912 (N_17912,N_11861,N_9153);
xnor U17913 (N_17913,N_7990,N_11601);
nor U17914 (N_17914,N_10123,N_9374);
and U17915 (N_17915,N_8423,N_9771);
nor U17916 (N_17916,N_9203,N_10863);
nor U17917 (N_17917,N_11982,N_7684);
or U17918 (N_17918,N_9060,N_7592);
or U17919 (N_17919,N_9445,N_7849);
and U17920 (N_17920,N_10868,N_6745);
nor U17921 (N_17921,N_10154,N_11020);
or U17922 (N_17922,N_10743,N_7556);
and U17923 (N_17923,N_7276,N_6570);
and U17924 (N_17924,N_9613,N_6388);
and U17925 (N_17925,N_9209,N_9783);
nor U17926 (N_17926,N_10266,N_8519);
nand U17927 (N_17927,N_7277,N_9510);
xnor U17928 (N_17928,N_8831,N_8076);
and U17929 (N_17929,N_6452,N_6883);
nor U17930 (N_17930,N_9697,N_11787);
or U17931 (N_17931,N_11131,N_11946);
xor U17932 (N_17932,N_8473,N_11490);
and U17933 (N_17933,N_8569,N_10624);
or U17934 (N_17934,N_11538,N_8476);
and U17935 (N_17935,N_9233,N_7527);
or U17936 (N_17936,N_6373,N_6849);
or U17937 (N_17937,N_7693,N_11703);
and U17938 (N_17938,N_10169,N_9755);
or U17939 (N_17939,N_8187,N_9870);
nand U17940 (N_17940,N_7996,N_8698);
nor U17941 (N_17941,N_6589,N_7696);
or U17942 (N_17942,N_10486,N_8859);
or U17943 (N_17943,N_9826,N_6596);
and U17944 (N_17944,N_8438,N_9450);
nand U17945 (N_17945,N_11541,N_10305);
nand U17946 (N_17946,N_7849,N_11131);
nand U17947 (N_17947,N_7925,N_9398);
nand U17948 (N_17948,N_10836,N_9398);
or U17949 (N_17949,N_9216,N_7182);
nand U17950 (N_17950,N_9612,N_6885);
nor U17951 (N_17951,N_7278,N_11017);
xnor U17952 (N_17952,N_6919,N_6642);
nand U17953 (N_17953,N_8869,N_11678);
and U17954 (N_17954,N_9618,N_8287);
nand U17955 (N_17955,N_6621,N_11465);
or U17956 (N_17956,N_11469,N_8491);
or U17957 (N_17957,N_9536,N_8535);
or U17958 (N_17958,N_6155,N_11493);
and U17959 (N_17959,N_9784,N_7279);
nor U17960 (N_17960,N_8657,N_9966);
nor U17961 (N_17961,N_7210,N_8981);
or U17962 (N_17962,N_11133,N_8470);
nand U17963 (N_17963,N_6995,N_8560);
nand U17964 (N_17964,N_7415,N_10447);
nand U17965 (N_17965,N_8364,N_8687);
or U17966 (N_17966,N_8819,N_11039);
nor U17967 (N_17967,N_8306,N_9250);
nor U17968 (N_17968,N_7435,N_9460);
or U17969 (N_17969,N_11490,N_10465);
or U17970 (N_17970,N_10045,N_10060);
nor U17971 (N_17971,N_10688,N_10122);
and U17972 (N_17972,N_8272,N_8150);
or U17973 (N_17973,N_8489,N_6854);
and U17974 (N_17974,N_8122,N_6113);
nor U17975 (N_17975,N_10399,N_9039);
and U17976 (N_17976,N_10612,N_10941);
or U17977 (N_17977,N_6424,N_7209);
or U17978 (N_17978,N_7031,N_10742);
or U17979 (N_17979,N_8160,N_11854);
or U17980 (N_17980,N_7329,N_9555);
xor U17981 (N_17981,N_11378,N_10297);
xnor U17982 (N_17982,N_6117,N_7751);
nor U17983 (N_17983,N_10113,N_11995);
and U17984 (N_17984,N_8161,N_11935);
nand U17985 (N_17985,N_7938,N_8708);
nor U17986 (N_17986,N_7139,N_8400);
xor U17987 (N_17987,N_11647,N_7134);
nand U17988 (N_17988,N_7244,N_9187);
or U17989 (N_17989,N_6037,N_11003);
nor U17990 (N_17990,N_10073,N_10743);
xor U17991 (N_17991,N_8410,N_10061);
and U17992 (N_17992,N_8740,N_7924);
or U17993 (N_17993,N_6791,N_7708);
nand U17994 (N_17994,N_7840,N_8610);
nor U17995 (N_17995,N_9053,N_11784);
nor U17996 (N_17996,N_7364,N_9919);
or U17997 (N_17997,N_8747,N_11217);
xor U17998 (N_17998,N_6490,N_9813);
and U17999 (N_17999,N_7290,N_10543);
nor U18000 (N_18000,N_13035,N_12522);
and U18001 (N_18001,N_12112,N_13268);
nand U18002 (N_18002,N_12089,N_16031);
and U18003 (N_18003,N_13996,N_12540);
or U18004 (N_18004,N_13616,N_13100);
or U18005 (N_18005,N_14528,N_14911);
or U18006 (N_18006,N_16991,N_14546);
nor U18007 (N_18007,N_14814,N_15825);
and U18008 (N_18008,N_17797,N_15218);
or U18009 (N_18009,N_16121,N_17839);
nand U18010 (N_18010,N_16332,N_14271);
or U18011 (N_18011,N_13610,N_16523);
or U18012 (N_18012,N_13811,N_16637);
or U18013 (N_18013,N_14909,N_13861);
nand U18014 (N_18014,N_16139,N_16351);
or U18015 (N_18015,N_12763,N_15383);
and U18016 (N_18016,N_12663,N_12789);
nor U18017 (N_18017,N_15120,N_15592);
or U18018 (N_18018,N_16621,N_14358);
nor U18019 (N_18019,N_16609,N_14202);
nor U18020 (N_18020,N_12185,N_15221);
nor U18021 (N_18021,N_17953,N_16159);
and U18022 (N_18022,N_16452,N_17090);
or U18023 (N_18023,N_14779,N_16221);
and U18024 (N_18024,N_13865,N_15616);
or U18025 (N_18025,N_15308,N_14997);
nand U18026 (N_18026,N_13767,N_16875);
nor U18027 (N_18027,N_12672,N_17507);
and U18028 (N_18028,N_16883,N_15949);
xor U18029 (N_18029,N_16404,N_14153);
and U18030 (N_18030,N_13603,N_15016);
nor U18031 (N_18031,N_17144,N_14910);
nand U18032 (N_18032,N_14018,N_15496);
or U18033 (N_18033,N_17021,N_17730);
nor U18034 (N_18034,N_14119,N_16175);
and U18035 (N_18035,N_12684,N_17429);
and U18036 (N_18036,N_17273,N_16367);
nor U18037 (N_18037,N_17221,N_13226);
nor U18038 (N_18038,N_12733,N_15943);
and U18039 (N_18039,N_16636,N_12719);
nand U18040 (N_18040,N_12421,N_15320);
or U18041 (N_18041,N_16516,N_15623);
or U18042 (N_18042,N_12065,N_16323);
nor U18043 (N_18043,N_12157,N_14255);
and U18044 (N_18044,N_13870,N_15959);
xor U18045 (N_18045,N_13698,N_17950);
or U18046 (N_18046,N_16957,N_12600);
nor U18047 (N_18047,N_12989,N_17177);
nor U18048 (N_18048,N_16830,N_15967);
xor U18049 (N_18049,N_15673,N_16925);
nor U18050 (N_18050,N_12103,N_17163);
or U18051 (N_18051,N_15029,N_12251);
and U18052 (N_18052,N_12514,N_16937);
or U18053 (N_18053,N_13313,N_12200);
xor U18054 (N_18054,N_16580,N_13793);
and U18055 (N_18055,N_17464,N_17160);
nor U18056 (N_18056,N_16115,N_13998);
xor U18057 (N_18057,N_12494,N_12113);
and U18058 (N_18058,N_17012,N_15651);
and U18059 (N_18059,N_14575,N_14876);
or U18060 (N_18060,N_14306,N_14195);
or U18061 (N_18061,N_12452,N_17552);
or U18062 (N_18062,N_12381,N_12035);
or U18063 (N_18063,N_15947,N_17959);
nor U18064 (N_18064,N_15377,N_17463);
and U18065 (N_18065,N_15887,N_13392);
or U18066 (N_18066,N_16095,N_12750);
and U18067 (N_18067,N_15505,N_15071);
xnor U18068 (N_18068,N_14444,N_14748);
and U18069 (N_18069,N_16357,N_12637);
nand U18070 (N_18070,N_17395,N_16951);
xor U18071 (N_18071,N_15174,N_12690);
nor U18072 (N_18072,N_14985,N_15873);
nor U18073 (N_18073,N_14366,N_15529);
or U18074 (N_18074,N_17592,N_17087);
nor U18075 (N_18075,N_14936,N_16709);
or U18076 (N_18076,N_17046,N_14436);
nor U18077 (N_18077,N_15039,N_12956);
or U18078 (N_18078,N_17248,N_13263);
nand U18079 (N_18079,N_14058,N_15042);
and U18080 (N_18080,N_17741,N_14125);
nor U18081 (N_18081,N_16807,N_12705);
nand U18082 (N_18082,N_12068,N_17536);
and U18083 (N_18083,N_15695,N_15667);
nor U18084 (N_18084,N_16873,N_16038);
nand U18085 (N_18085,N_13476,N_12077);
and U18086 (N_18086,N_17212,N_17722);
or U18087 (N_18087,N_16395,N_15040);
nor U18088 (N_18088,N_13242,N_16559);
nand U18089 (N_18089,N_15437,N_17166);
xnor U18090 (N_18090,N_16331,N_14784);
nand U18091 (N_18091,N_13790,N_17649);
and U18092 (N_18092,N_14378,N_14389);
nand U18093 (N_18093,N_15010,N_15208);
nor U18094 (N_18094,N_12498,N_17532);
or U18095 (N_18095,N_16407,N_15580);
nor U18096 (N_18096,N_17339,N_14821);
or U18097 (N_18097,N_12471,N_14216);
nand U18098 (N_18098,N_14536,N_14923);
nand U18099 (N_18099,N_14386,N_15332);
and U18100 (N_18100,N_17267,N_13430);
or U18101 (N_18101,N_13097,N_15192);
xor U18102 (N_18102,N_16945,N_12550);
and U18103 (N_18103,N_15017,N_17140);
and U18104 (N_18104,N_15735,N_12899);
and U18105 (N_18105,N_13301,N_17566);
or U18106 (N_18106,N_12781,N_14360);
and U18107 (N_18107,N_16203,N_14327);
or U18108 (N_18108,N_12530,N_15966);
or U18109 (N_18109,N_15605,N_16555);
or U18110 (N_18110,N_14233,N_13349);
xnor U18111 (N_18111,N_12512,N_15474);
nor U18112 (N_18112,N_17199,N_13716);
or U18113 (N_18113,N_15155,N_15343);
or U18114 (N_18114,N_15544,N_14867);
nor U18115 (N_18115,N_13890,N_17089);
nand U18116 (N_18116,N_16895,N_14663);
and U18117 (N_18117,N_16693,N_15691);
and U18118 (N_18118,N_16504,N_15900);
nand U18119 (N_18119,N_14231,N_14213);
nand U18120 (N_18120,N_12225,N_16800);
and U18121 (N_18121,N_16855,N_14486);
nand U18122 (N_18122,N_13773,N_15729);
xor U18123 (N_18123,N_12734,N_17157);
nor U18124 (N_18124,N_14291,N_16836);
xnor U18125 (N_18125,N_12983,N_14700);
xnor U18126 (N_18126,N_15225,N_15807);
nand U18127 (N_18127,N_12335,N_15003);
nor U18128 (N_18128,N_17695,N_16814);
nor U18129 (N_18129,N_12838,N_12007);
or U18130 (N_18130,N_16944,N_12660);
nor U18131 (N_18131,N_12912,N_15122);
xnor U18132 (N_18132,N_16243,N_15407);
or U18133 (N_18133,N_15043,N_16804);
xnor U18134 (N_18134,N_16839,N_15431);
xor U18135 (N_18135,N_15455,N_16400);
or U18136 (N_18136,N_12428,N_12563);
nand U18137 (N_18137,N_13534,N_13553);
and U18138 (N_18138,N_15266,N_15709);
nor U18139 (N_18139,N_17268,N_13224);
nor U18140 (N_18140,N_14890,N_12859);
nand U18141 (N_18141,N_14014,N_14168);
nor U18142 (N_18142,N_13960,N_17851);
and U18143 (N_18143,N_14505,N_15446);
nor U18144 (N_18144,N_15141,N_13387);
and U18145 (N_18145,N_13023,N_15164);
and U18146 (N_18146,N_17848,N_16669);
or U18147 (N_18147,N_14975,N_12150);
and U18148 (N_18148,N_16554,N_12831);
nor U18149 (N_18149,N_13351,N_15892);
and U18150 (N_18150,N_13500,N_12067);
or U18151 (N_18151,N_14674,N_17644);
nor U18152 (N_18152,N_17294,N_15121);
and U18153 (N_18153,N_14706,N_17018);
and U18154 (N_18154,N_12223,N_13883);
nand U18155 (N_18155,N_14289,N_13763);
and U18156 (N_18156,N_13347,N_13673);
and U18157 (N_18157,N_17970,N_15538);
or U18158 (N_18158,N_17580,N_15823);
or U18159 (N_18159,N_17300,N_14384);
nand U18160 (N_18160,N_12994,N_17826);
or U18161 (N_18161,N_16885,N_17436);
and U18162 (N_18162,N_13194,N_12279);
and U18163 (N_18163,N_16168,N_14776);
nand U18164 (N_18164,N_16756,N_17745);
or U18165 (N_18165,N_13486,N_13501);
nor U18166 (N_18166,N_14065,N_17051);
and U18167 (N_18167,N_15798,N_17636);
and U18168 (N_18168,N_14833,N_15999);
and U18169 (N_18169,N_14376,N_12709);
or U18170 (N_18170,N_17265,N_15273);
and U18171 (N_18171,N_13297,N_12726);
or U18172 (N_18172,N_12119,N_12454);
nand U18173 (N_18173,N_14007,N_13970);
nor U18174 (N_18174,N_13646,N_17215);
and U18175 (N_18175,N_16443,N_14917);
nor U18176 (N_18176,N_13593,N_13897);
or U18177 (N_18177,N_14090,N_13241);
nand U18178 (N_18178,N_14357,N_15636);
nor U18179 (N_18179,N_15844,N_14355);
nand U18180 (N_18180,N_17928,N_13852);
nand U18181 (N_18181,N_17669,N_15187);
or U18182 (N_18182,N_13468,N_16787);
nor U18183 (N_18183,N_17861,N_13190);
nand U18184 (N_18184,N_14515,N_13722);
or U18185 (N_18185,N_15613,N_15188);
nand U18186 (N_18186,N_12212,N_14320);
nand U18187 (N_18187,N_15771,N_15049);
xor U18188 (N_18188,N_16252,N_14173);
nor U18189 (N_18189,N_14801,N_14749);
nand U18190 (N_18190,N_15297,N_17183);
or U18191 (N_18191,N_12260,N_16929);
nor U18192 (N_18192,N_17443,N_12560);
and U18193 (N_18193,N_13532,N_12960);
xor U18194 (N_18194,N_15839,N_13346);
nor U18195 (N_18195,N_16356,N_14217);
nand U18196 (N_18196,N_14276,N_16440);
or U18197 (N_18197,N_16717,N_13580);
xor U18198 (N_18198,N_15766,N_15097);
and U18199 (N_18199,N_15952,N_14495);
and U18200 (N_18200,N_16600,N_14336);
nor U18201 (N_18201,N_15159,N_16042);
and U18202 (N_18202,N_17086,N_13528);
or U18203 (N_18203,N_12674,N_16973);
or U18204 (N_18204,N_17800,N_16565);
nand U18205 (N_18205,N_13664,N_17107);
nor U18206 (N_18206,N_13055,N_14569);
nor U18207 (N_18207,N_14503,N_17486);
nand U18208 (N_18208,N_15813,N_14507);
or U18209 (N_18209,N_16808,N_13115);
nand U18210 (N_18210,N_14193,N_12451);
nand U18211 (N_18211,N_13391,N_14682);
nor U18212 (N_18212,N_13658,N_13676);
nor U18213 (N_18213,N_16892,N_12622);
nor U18214 (N_18214,N_12860,N_14281);
or U18215 (N_18215,N_13704,N_14548);
nand U18216 (N_18216,N_16930,N_13257);
nor U18217 (N_18217,N_16143,N_12356);
and U18218 (N_18218,N_15539,N_15520);
xnor U18219 (N_18219,N_12677,N_12752);
and U18220 (N_18220,N_16623,N_12032);
or U18221 (N_18221,N_16100,N_12747);
nor U18222 (N_18222,N_14619,N_16321);
xnor U18223 (N_18223,N_17736,N_15404);
xor U18224 (N_18224,N_17158,N_13582);
or U18225 (N_18225,N_17358,N_17099);
or U18226 (N_18226,N_17804,N_13556);
nor U18227 (N_18227,N_15657,N_13045);
and U18228 (N_18228,N_13344,N_17511);
nor U18229 (N_18229,N_15650,N_14547);
or U18230 (N_18230,N_12244,N_16428);
and U18231 (N_18231,N_17923,N_13130);
and U18232 (N_18232,N_13508,N_15819);
nand U18233 (N_18233,N_16272,N_16575);
nand U18234 (N_18234,N_17266,N_17870);
xor U18235 (N_18235,N_13419,N_14309);
and U18236 (N_18236,N_14511,N_17972);
xnor U18237 (N_18237,N_16998,N_13940);
or U18238 (N_18238,N_16087,N_14981);
xnor U18239 (N_18239,N_14310,N_14613);
xnor U18240 (N_18240,N_17508,N_16550);
and U18241 (N_18241,N_16616,N_17392);
nor U18242 (N_18242,N_15290,N_16269);
or U18243 (N_18243,N_14356,N_12780);
and U18244 (N_18244,N_12430,N_17220);
nand U18245 (N_18245,N_16140,N_14282);
nand U18246 (N_18246,N_17312,N_17834);
xor U18247 (N_18247,N_16292,N_14907);
or U18248 (N_18248,N_15974,N_12256);
or U18249 (N_18249,N_17001,N_17407);
and U18250 (N_18250,N_12608,N_14257);
nor U18251 (N_18251,N_13641,N_14442);
nor U18252 (N_18252,N_13353,N_16674);
nand U18253 (N_18253,N_17825,N_13250);
nor U18254 (N_18254,N_16904,N_16587);
nor U18255 (N_18255,N_15843,N_14154);
xnor U18256 (N_18256,N_16799,N_16455);
and U18257 (N_18257,N_17355,N_13173);
nand U18258 (N_18258,N_14599,N_15731);
and U18259 (N_18259,N_14425,N_16234);
xor U18260 (N_18260,N_16411,N_15091);
nor U18261 (N_18261,N_15961,N_17269);
xor U18262 (N_18262,N_12576,N_14326);
nand U18263 (N_18263,N_15791,N_14071);
nor U18264 (N_18264,N_13657,N_13164);
nor U18265 (N_18265,N_14052,N_13845);
nor U18266 (N_18266,N_12629,N_13216);
nor U18267 (N_18267,N_16166,N_14038);
nand U18268 (N_18268,N_17942,N_14432);
and U18269 (N_18269,N_14210,N_12958);
nand U18270 (N_18270,N_16826,N_12375);
and U18271 (N_18271,N_12346,N_17143);
and U18272 (N_18272,N_15341,N_15513);
xnor U18273 (N_18273,N_14820,N_16491);
and U18274 (N_18274,N_16134,N_17706);
nand U18275 (N_18275,N_12334,N_12390);
nor U18276 (N_18276,N_16336,N_16903);
nand U18277 (N_18277,N_17381,N_13458);
and U18278 (N_18278,N_14246,N_14369);
nor U18279 (N_18279,N_12382,N_13921);
or U18280 (N_18280,N_15555,N_13374);
xnor U18281 (N_18281,N_14886,N_17216);
nor U18282 (N_18282,N_17367,N_16771);
nor U18283 (N_18283,N_17313,N_14864);
nand U18284 (N_18284,N_16970,N_17638);
and U18285 (N_18285,N_14417,N_14013);
nor U18286 (N_18286,N_12299,N_17354);
nor U18287 (N_18287,N_13733,N_15591);
or U18288 (N_18288,N_12500,N_16278);
and U18289 (N_18289,N_13195,N_14460);
and U18290 (N_18290,N_14269,N_13814);
or U18291 (N_18291,N_13215,N_16192);
or U18292 (N_18292,N_15270,N_14677);
nand U18293 (N_18293,N_12144,N_17662);
nand U18294 (N_18294,N_14318,N_14262);
nor U18295 (N_18295,N_17694,N_14298);
nand U18296 (N_18296,N_12946,N_16760);
nand U18297 (N_18297,N_15160,N_15727);
and U18298 (N_18298,N_12016,N_15272);
nor U18299 (N_18299,N_15009,N_15621);
or U18300 (N_18300,N_16412,N_15182);
and U18301 (N_18301,N_13197,N_12025);
or U18302 (N_18302,N_16853,N_17147);
or U18303 (N_18303,N_16186,N_16309);
nor U18304 (N_18304,N_14681,N_15235);
nand U18305 (N_18305,N_13207,N_16436);
or U18306 (N_18306,N_15023,N_16479);
or U18307 (N_18307,N_12728,N_15792);
nand U18308 (N_18308,N_13804,N_14448);
and U18309 (N_18309,N_12121,N_14147);
and U18310 (N_18310,N_14483,N_17139);
nor U18311 (N_18311,N_16920,N_14330);
nor U18312 (N_18312,N_15133,N_16313);
nand U18313 (N_18313,N_14238,N_15213);
xor U18314 (N_18314,N_13398,N_14328);
nor U18315 (N_18315,N_17752,N_13587);
and U18316 (N_18316,N_15161,N_13723);
or U18317 (N_18317,N_15686,N_17622);
nor U18318 (N_18318,N_13361,N_12126);
and U18319 (N_18319,N_13544,N_16641);
nor U18320 (N_18320,N_13399,N_16703);
or U18321 (N_18321,N_16796,N_16975);
xor U18322 (N_18322,N_14343,N_15794);
and U18323 (N_18323,N_16739,N_17047);
or U18324 (N_18324,N_14521,N_16349);
and U18325 (N_18325,N_14322,N_12171);
or U18326 (N_18326,N_12557,N_15903);
nor U18327 (N_18327,N_13525,N_12701);
nand U18328 (N_18328,N_12919,N_17128);
nor U18329 (N_18329,N_15503,N_17779);
or U18330 (N_18330,N_14443,N_14106);
or U18331 (N_18331,N_12080,N_12193);
or U18332 (N_18332,N_15850,N_17759);
nand U18333 (N_18333,N_13254,N_12468);
or U18334 (N_18334,N_16795,N_13548);
nor U18335 (N_18335,N_16268,N_12605);
or U18336 (N_18336,N_17180,N_15124);
and U18337 (N_18337,N_14070,N_12991);
nor U18338 (N_18338,N_12499,N_14169);
or U18339 (N_18339,N_13323,N_14691);
or U18340 (N_18340,N_13266,N_12646);
and U18341 (N_18341,N_13415,N_13234);
or U18342 (N_18342,N_12511,N_15630);
nand U18343 (N_18343,N_15190,N_14032);
nand U18344 (N_18344,N_13373,N_14347);
and U18345 (N_18345,N_16144,N_13070);
and U18346 (N_18346,N_13154,N_16802);
xnor U18347 (N_18347,N_14720,N_12883);
and U18348 (N_18348,N_14782,N_16818);
nand U18349 (N_18349,N_13423,N_15024);
nand U18350 (N_18350,N_16276,N_13341);
and U18351 (N_18351,N_16364,N_13686);
and U18352 (N_18352,N_13005,N_12207);
and U18353 (N_18353,N_17224,N_16563);
and U18354 (N_18354,N_12152,N_15781);
nor U18355 (N_18355,N_17004,N_17737);
and U18356 (N_18356,N_13849,N_16206);
nand U18357 (N_18357,N_14179,N_16880);
or U18358 (N_18358,N_12643,N_12350);
and U18359 (N_18359,N_13752,N_13455);
nor U18360 (N_18360,N_14571,N_17547);
or U18361 (N_18361,N_16135,N_13796);
nor U18362 (N_18362,N_12389,N_13188);
nand U18363 (N_18363,N_15851,N_12475);
and U18364 (N_18364,N_16230,N_14969);
xor U18365 (N_18365,N_15109,N_13911);
or U18366 (N_18366,N_12572,N_17013);
xor U18367 (N_18367,N_13731,N_13251);
nor U18368 (N_18368,N_12866,N_12014);
xor U18369 (N_18369,N_17445,N_17746);
and U18370 (N_18370,N_17259,N_14746);
nor U18371 (N_18371,N_15713,N_17304);
and U18372 (N_18372,N_17491,N_16431);
or U18373 (N_18373,N_16173,N_12783);
nand U18374 (N_18374,N_17005,N_15902);
nand U18375 (N_18375,N_14803,N_17109);
nand U18376 (N_18376,N_16255,N_16982);
nor U18377 (N_18377,N_13860,N_15963);
nor U18378 (N_18378,N_13143,N_16105);
nor U18379 (N_18379,N_17346,N_17587);
and U18380 (N_18380,N_13933,N_16061);
nand U18381 (N_18381,N_13627,N_14144);
nand U18382 (N_18382,N_13677,N_13880);
or U18383 (N_18383,N_12263,N_15107);
xnor U18384 (N_18384,N_16456,N_17353);
nor U18385 (N_18385,N_13329,N_14739);
or U18386 (N_18386,N_12470,N_12008);
and U18387 (N_18387,N_14512,N_14897);
xnor U18388 (N_18388,N_13208,N_12533);
nand U18389 (N_18389,N_17850,N_15051);
and U18390 (N_18390,N_13111,N_12174);
nor U18391 (N_18391,N_14753,N_16153);
nor U18392 (N_18392,N_17809,N_16626);
nand U18393 (N_18393,N_17891,N_13309);
nor U18394 (N_18394,N_17831,N_15284);
nand U18395 (N_18395,N_12493,N_16645);
or U18396 (N_18396,N_14802,N_16696);
or U18397 (N_18397,N_13795,N_12827);
nand U18398 (N_18398,N_17028,N_15359);
nand U18399 (N_18399,N_17666,N_13778);
or U18400 (N_18400,N_12175,N_13404);
xnor U18401 (N_18401,N_13617,N_16029);
nand U18402 (N_18402,N_16544,N_16156);
or U18403 (N_18403,N_13535,N_14260);
and U18404 (N_18404,N_17727,N_17461);
nand U18405 (N_18405,N_13975,N_17836);
xor U18406 (N_18406,N_16235,N_15973);
or U18407 (N_18407,N_14604,N_17119);
nand U18408 (N_18408,N_16767,N_17434);
or U18409 (N_18409,N_15214,N_16040);
nand U18410 (N_18410,N_12180,N_15327);
xor U18411 (N_18411,N_17871,N_16274);
and U18412 (N_18412,N_14411,N_12039);
xnor U18413 (N_18413,N_14423,N_16705);
or U18414 (N_18414,N_13298,N_16145);
nand U18415 (N_18415,N_13024,N_14516);
nand U18416 (N_18416,N_17898,N_14945);
or U18417 (N_18417,N_14733,N_12926);
and U18418 (N_18418,N_12597,N_14471);
nor U18419 (N_18419,N_15550,N_12137);
and U18420 (N_18420,N_15302,N_16147);
xor U18421 (N_18421,N_12809,N_15595);
xor U18422 (N_18422,N_16577,N_15594);
and U18423 (N_18423,N_16299,N_17738);
nand U18424 (N_18424,N_13537,N_17169);
nor U18425 (N_18425,N_13016,N_15779);
nand U18426 (N_18426,N_16414,N_17814);
or U18427 (N_18427,N_13915,N_13966);
or U18428 (N_18428,N_13333,N_12074);
or U18429 (N_18429,N_12768,N_12415);
nor U18430 (N_18430,N_12010,N_14489);
or U18431 (N_18431,N_15292,N_14073);
nor U18432 (N_18432,N_17561,N_17331);
or U18433 (N_18433,N_13262,N_17921);
nand U18434 (N_18434,N_13775,N_17802);
xor U18435 (N_18435,N_16392,N_13739);
or U18436 (N_18436,N_14451,N_16605);
nand U18437 (N_18437,N_17875,N_12241);
and U18438 (N_18438,N_12894,N_17074);
nand U18439 (N_18439,N_14829,N_12354);
or U18440 (N_18440,N_13409,N_15413);
and U18441 (N_18441,N_13956,N_14526);
nor U18442 (N_18442,N_16989,N_15674);
xor U18443 (N_18443,N_12440,N_17103);
or U18444 (N_18444,N_13439,N_14069);
or U18445 (N_18445,N_15914,N_17975);
and U18446 (N_18446,N_16646,N_16160);
nor U18447 (N_18447,N_12913,N_16701);
nor U18448 (N_18448,N_17717,N_13381);
nand U18449 (N_18449,N_13365,N_17148);
or U18450 (N_18450,N_15699,N_17557);
nor U18451 (N_18451,N_13978,N_15940);
nor U18452 (N_18452,N_16076,N_15955);
nand U18453 (N_18453,N_17444,N_13674);
xnor U18454 (N_18454,N_13276,N_16311);
and U18455 (N_18455,N_16766,N_17543);
and U18456 (N_18456,N_17612,N_15363);
and U18457 (N_18457,N_14822,N_13974);
and U18458 (N_18458,N_13269,N_13819);
nand U18459 (N_18459,N_13284,N_13103);
nand U18460 (N_18460,N_14824,N_17778);
or U18461 (N_18461,N_15501,N_15833);
nor U18462 (N_18462,N_14990,N_13871);
nor U18463 (N_18463,N_13252,N_17022);
or U18464 (N_18464,N_13245,N_12638);
nor U18465 (N_18465,N_13780,N_14948);
xor U18466 (N_18466,N_12036,N_14063);
and U18467 (N_18467,N_14484,N_14364);
xor U18468 (N_18468,N_16542,N_13924);
nand U18469 (N_18469,N_17306,N_12448);
xnor U18470 (N_18470,N_14041,N_16191);
nand U18471 (N_18471,N_14405,N_16288);
and U18472 (N_18472,N_14670,N_16813);
and U18473 (N_18473,N_13182,N_14053);
nor U18474 (N_18474,N_14609,N_12749);
nor U18475 (N_18475,N_14178,N_12096);
or U18476 (N_18476,N_15954,N_14253);
xnor U18477 (N_18477,N_13302,N_15768);
xor U18478 (N_18478,N_15842,N_14190);
nand U18479 (N_18479,N_17805,N_17941);
nand U18480 (N_18480,N_12274,N_14797);
or U18481 (N_18481,N_17165,N_14970);
or U18482 (N_18482,N_16439,N_15325);
and U18483 (N_18483,N_16028,N_15484);
nand U18484 (N_18484,N_14049,N_16379);
and U18485 (N_18485,N_13163,N_16784);
and U18486 (N_18486,N_16869,N_16141);
and U18487 (N_18487,N_16627,N_15965);
and U18488 (N_18488,N_13908,N_17493);
and U18489 (N_18489,N_15658,N_12122);
nor U18490 (N_18490,N_13138,N_15546);
nor U18491 (N_18491,N_12811,N_16026);
nand U18492 (N_18492,N_13759,N_15635);
xor U18493 (N_18493,N_17788,N_13813);
xor U18494 (N_18494,N_15547,N_15475);
nor U18495 (N_18495,N_14350,N_17112);
nand U18496 (N_18496,N_15465,N_16898);
and U18497 (N_18497,N_13126,N_13895);
or U18498 (N_18498,N_14046,N_15719);
and U18499 (N_18499,N_14553,N_14592);
nor U18500 (N_18500,N_15867,N_12665);
nand U18501 (N_18501,N_12053,N_12182);
or U18502 (N_18502,N_13136,N_16675);
nor U18503 (N_18503,N_16886,N_15527);
and U18504 (N_18504,N_12484,N_13105);
nor U18505 (N_18505,N_16539,N_15783);
and U18506 (N_18506,N_15622,N_12617);
nand U18507 (N_18507,N_17780,N_16689);
nand U18508 (N_18508,N_16908,N_13411);
and U18509 (N_18509,N_14767,N_14109);
and U18510 (N_18510,N_14894,N_14794);
or U18511 (N_18511,N_15656,N_12153);
nor U18512 (N_18512,N_17155,N_13081);
and U18513 (N_18513,N_13095,N_16004);
and U18514 (N_18514,N_16934,N_17883);
nor U18515 (N_18515,N_12105,N_17991);
xor U18516 (N_18516,N_15294,N_12073);
and U18517 (N_18517,N_14919,N_17280);
and U18518 (N_18518,N_16517,N_14447);
or U18519 (N_18519,N_12323,N_16682);
nor U18520 (N_18520,N_13573,N_15767);
nor U18521 (N_18521,N_12407,N_16840);
or U18522 (N_18522,N_17417,N_15577);
nor U18523 (N_18523,N_12358,N_12710);
nor U18524 (N_18524,N_14114,N_17524);
nor U18525 (N_18525,N_17235,N_17934);
nor U18526 (N_18526,N_16535,N_14137);
and U18527 (N_18527,N_13934,N_13651);
and U18528 (N_18528,N_13020,N_14439);
and U18529 (N_18529,N_14935,N_12867);
nor U18530 (N_18530,N_16481,N_17696);
or U18531 (N_18531,N_14621,N_17541);
or U18532 (N_18532,N_16429,N_12967);
nor U18533 (N_18533,N_12614,N_16861);
nor U18534 (N_18534,N_12490,N_12170);
or U18535 (N_18535,N_12235,N_14398);
or U18536 (N_18536,N_17520,N_14514);
nand U18537 (N_18537,N_15370,N_16845);
or U18538 (N_18538,N_15126,N_14678);
or U18539 (N_18539,N_16453,N_12116);
and U18540 (N_18540,N_17402,N_17209);
and U18541 (N_18541,N_12107,N_16205);
xor U18542 (N_18542,N_13491,N_13655);
nor U18543 (N_18543,N_15425,N_13388);
xor U18544 (N_18544,N_12020,N_12296);
or U18545 (N_18545,N_16218,N_17404);
or U18546 (N_18546,N_16497,N_16859);
nand U18547 (N_18547,N_12215,N_16533);
nand U18548 (N_18548,N_12562,N_12775);
or U18549 (N_18549,N_15210,N_14245);
nand U18550 (N_18550,N_17329,N_14224);
and U18551 (N_18551,N_15930,N_17560);
nor U18552 (N_18552,N_16667,N_15316);
or U18553 (N_18553,N_14946,N_15714);
nor U18554 (N_18554,N_14696,N_17902);
and U18555 (N_18555,N_15884,N_15941);
and U18556 (N_18556,N_15113,N_15811);
nor U18557 (N_18557,N_15131,N_12250);
xnor U18558 (N_18558,N_15036,N_15847);
nor U18559 (N_18559,N_16935,N_13666);
and U18560 (N_18560,N_14028,N_16372);
nor U18561 (N_18561,N_13529,N_15923);
and U18562 (N_18562,N_16393,N_12839);
or U18563 (N_18563,N_17065,N_16547);
nand U18564 (N_18564,N_12851,N_14593);
nor U18565 (N_18565,N_13256,N_12195);
nor U18566 (N_18566,N_14450,N_15898);
nor U18567 (N_18567,N_13253,N_13267);
or U18568 (N_18568,N_16619,N_13031);
nor U18569 (N_18569,N_13776,N_15597);
nor U18570 (N_18570,N_15429,N_13010);
and U18571 (N_18571,N_15393,N_17968);
or U18572 (N_18572,N_15692,N_17734);
or U18573 (N_18573,N_15293,N_15560);
nor U18574 (N_18574,N_15780,N_13086);
nand U18575 (N_18575,N_17205,N_15426);
nand U18576 (N_18576,N_14139,N_16936);
and U18577 (N_18577,N_16154,N_14500);
nor U18578 (N_18578,N_15603,N_12070);
xnor U18579 (N_18579,N_17015,N_13570);
nand U18580 (N_18580,N_14457,N_17763);
nor U18581 (N_18581,N_13828,N_15770);
nor U18582 (N_18582,N_15706,N_15005);
and U18583 (N_18583,N_15250,N_15072);
nand U18584 (N_18584,N_14170,N_15335);
nand U18585 (N_18585,N_12050,N_14286);
nand U18586 (N_18586,N_15864,N_15322);
nand U18587 (N_18587,N_17455,N_17326);
and U18588 (N_18588,N_14698,N_15611);
nor U18589 (N_18589,N_15816,N_17314);
or U18590 (N_18590,N_13239,N_14266);
nor U18591 (N_18591,N_12968,N_15764);
or U18592 (N_18592,N_14818,N_13511);
and U18593 (N_18593,N_17364,N_16918);
nor U18594 (N_18594,N_17878,N_15830);
or U18595 (N_18595,N_17892,N_15946);
and U18596 (N_18596,N_12676,N_17900);
nand U18597 (N_18597,N_17389,N_14134);
or U18598 (N_18598,N_17751,N_12847);
nor U18599 (N_18599,N_15749,N_13850);
nor U18600 (N_18600,N_15763,N_12849);
or U18601 (N_18601,N_16879,N_15100);
nor U18602 (N_18602,N_16197,N_15321);
nor U18603 (N_18603,N_14305,N_12276);
xor U18604 (N_18604,N_13675,N_13069);
xor U18605 (N_18605,N_15608,N_17609);
nand U18606 (N_18606,N_14382,N_15606);
nand U18607 (N_18607,N_13769,N_15566);
xnor U18608 (N_18608,N_12298,N_15241);
nand U18609 (N_18609,N_13406,N_12516);
nand U18610 (N_18610,N_17952,N_16915);
or U18611 (N_18611,N_14734,N_13555);
nor U18612 (N_18612,N_15128,N_12474);
and U18613 (N_18613,N_15534,N_16229);
nor U18614 (N_18614,N_16995,N_13585);
or U18615 (N_18615,N_13987,N_13132);
nor U18616 (N_18616,N_13495,N_15876);
and U18617 (N_18617,N_16104,N_14345);
and U18618 (N_18618,N_16996,N_13509);
nand U18619 (N_18619,N_14819,N_13041);
nor U18620 (N_18620,N_16971,N_17213);
or U18621 (N_18621,N_15185,N_15263);
xor U18622 (N_18622,N_16521,N_17400);
nor U18623 (N_18623,N_13701,N_13331);
and U18624 (N_18624,N_14497,N_14697);
xnor U18625 (N_18625,N_13464,N_17024);
nand U18626 (N_18626,N_16490,N_14591);
or U18627 (N_18627,N_15001,N_17011);
and U18628 (N_18628,N_13560,N_12848);
and U18629 (N_18629,N_13859,N_12214);
or U18630 (N_18630,N_16571,N_13094);
and U18631 (N_18631,N_16190,N_15531);
nor U18632 (N_18632,N_13785,N_17468);
nor U18633 (N_18633,N_12264,N_13893);
and U18634 (N_18634,N_12102,N_15193);
nand U18635 (N_18635,N_12973,N_13597);
or U18636 (N_18636,N_13988,N_16953);
nor U18637 (N_18637,N_12104,N_15666);
and U18638 (N_18638,N_17880,N_17671);
nor U18639 (N_18639,N_13390,N_15329);
nor U18640 (N_18640,N_14072,N_14397);
and U18641 (N_18641,N_12097,N_14695);
and U18642 (N_18642,N_16743,N_13211);
nor U18643 (N_18643,N_12247,N_14810);
nand U18644 (N_18644,N_17689,N_16376);
nand U18645 (N_18645,N_15810,N_15257);
and U18646 (N_18646,N_12978,N_14949);
xnor U18647 (N_18647,N_12376,N_13470);
nand U18648 (N_18648,N_15443,N_12741);
nor U18649 (N_18649,N_14718,N_13687);
and U18650 (N_18650,N_14413,N_12717);
or U18651 (N_18651,N_17170,N_13074);
and U18652 (N_18652,N_17083,N_16763);
or U18653 (N_18653,N_15863,N_17685);
nor U18654 (N_18654,N_17299,N_17260);
and U18655 (N_18655,N_17988,N_17571);
and U18656 (N_18656,N_16240,N_17371);
nor U18657 (N_18657,N_13345,N_12554);
or U18658 (N_18658,N_16174,N_16486);
and U18659 (N_18659,N_13036,N_14261);
and U18660 (N_18660,N_12515,N_12508);
nand U18661 (N_18661,N_17192,N_12670);
nor U18662 (N_18662,N_17100,N_13109);
or U18663 (N_18663,N_15919,N_13789);
and U18664 (N_18664,N_13127,N_16488);
xnor U18665 (N_18665,N_16713,N_13884);
nor U18666 (N_18666,N_13170,N_15145);
nand U18667 (N_18667,N_13142,N_15707);
nor U18668 (N_18668,N_13873,N_14554);
nor U18669 (N_18669,N_15401,N_15556);
or U18670 (N_18670,N_16657,N_16074);
or U18671 (N_18671,N_14307,N_15201);
and U18672 (N_18672,N_13389,N_13564);
nor U18673 (N_18673,N_16365,N_14579);
nand U18674 (N_18674,N_14564,N_16136);
and U18675 (N_18675,N_15701,N_12852);
nand U18676 (N_18676,N_15751,N_15716);
and U18677 (N_18677,N_14212,N_12396);
and U18678 (N_18678,N_16591,N_17393);
nand U18679 (N_18679,N_15567,N_13835);
nand U18680 (N_18680,N_12159,N_14264);
or U18681 (N_18681,N_12364,N_16677);
xnor U18682 (N_18682,N_12374,N_17523);
or U18683 (N_18683,N_12972,N_12785);
nor U18684 (N_18684,N_16334,N_14319);
xnor U18685 (N_18685,N_12723,N_13292);
and U18686 (N_18686,N_13450,N_16803);
nor U18687 (N_18687,N_14081,N_12921);
nand U18688 (N_18688,N_13113,N_12422);
or U18689 (N_18689,N_17704,N_17263);
or U18690 (N_18690,N_14277,N_15697);
and U18691 (N_18691,N_17359,N_12664);
and U18692 (N_18692,N_16858,N_15398);
nor U18693 (N_18693,N_16058,N_16708);
nor U18694 (N_18694,N_15098,N_14311);
nor U18695 (N_18695,N_12856,N_16036);
and U18696 (N_18696,N_16341,N_14206);
nand U18697 (N_18697,N_15306,N_16169);
or U18698 (N_18698,N_13414,N_16672);
nor U18699 (N_18699,N_16769,N_15360);
and U18700 (N_18700,N_17688,N_13968);
nor U18701 (N_18701,N_12965,N_13885);
and U18702 (N_18702,N_13906,N_17106);
nand U18703 (N_18703,N_17980,N_13485);
nor U18704 (N_18704,N_17929,N_15179);
or U18705 (N_18705,N_12801,N_15925);
nor U18706 (N_18706,N_12947,N_16772);
nor U18707 (N_18707,N_17098,N_14252);
and U18708 (N_18708,N_13363,N_14762);
and U18709 (N_18709,N_17503,N_13155);
nand U18710 (N_18710,N_17237,N_13581);
xnor U18711 (N_18711,N_12294,N_13905);
nand U18712 (N_18712,N_16196,N_15904);
xor U18713 (N_18713,N_12953,N_14117);
and U18714 (N_18714,N_17351,N_12527);
and U18715 (N_18715,N_13649,N_14996);
or U18716 (N_18716,N_17865,N_15627);
nor U18717 (N_18717,N_16724,N_12314);
nor U18718 (N_18718,N_15168,N_15136);
nor U18719 (N_18719,N_16241,N_17120);
nand U18720 (N_18720,N_12551,N_13247);
nand U18721 (N_18721,N_15046,N_13829);
nand U18722 (N_18722,N_14741,N_15416);
nand U18723 (N_18723,N_17422,N_16955);
nand U18724 (N_18724,N_16167,N_17595);
nand U18725 (N_18725,N_12133,N_13214);
xor U18726 (N_18726,N_14415,N_13713);
xor U18727 (N_18727,N_16078,N_17913);
and U18728 (N_18728,N_17616,N_14796);
nor U18729 (N_18729,N_12587,N_15415);
or U18730 (N_18730,N_13523,N_15158);
and U18731 (N_18731,N_16790,N_13550);
nor U18732 (N_18732,N_15761,N_12196);
nand U18733 (N_18733,N_13243,N_13076);
nand U18734 (N_18734,N_16279,N_17495);
nand U18735 (N_18735,N_17352,N_12117);
nand U18736 (N_18736,N_12595,N_13360);
nand U18737 (N_18737,N_14275,N_17519);
nand U18738 (N_18738,N_16825,N_12253);
xor U18739 (N_18739,N_12659,N_14723);
or U18740 (N_18740,N_12478,N_17575);
and U18741 (N_18741,N_14431,N_17888);
and U18742 (N_18742,N_15102,N_13437);
nand U18743 (N_18743,N_15521,N_15818);
nand U18744 (N_18744,N_14928,N_14921);
and U18745 (N_18745,N_13186,N_12844);
or U18746 (N_18746,N_14177,N_14589);
or U18747 (N_18747,N_15890,N_14557);
nand U18748 (N_18748,N_12940,N_16465);
nand U18749 (N_18749,N_12525,N_16089);
nor U18750 (N_18750,N_17282,N_17101);
or U18751 (N_18751,N_13071,N_17742);
or U18752 (N_18752,N_14469,N_17081);
nor U18753 (N_18753,N_12770,N_14964);
nand U18754 (N_18754,N_12488,N_16758);
or U18755 (N_18755,N_12132,N_15129);
or U18756 (N_18756,N_17327,N_16653);
xnor U18757 (N_18757,N_12406,N_16239);
or U18758 (N_18758,N_12347,N_13383);
or U18759 (N_18759,N_15957,N_14414);
and U18760 (N_18760,N_17659,N_14690);
nand U18761 (N_18761,N_15964,N_15523);
nand U18762 (N_18762,N_14400,N_14412);
nand U18763 (N_18763,N_16044,N_16640);
nand U18764 (N_18764,N_14644,N_13599);
or U18765 (N_18765,N_14680,N_16224);
xnor U18766 (N_18766,N_16094,N_15574);
nand U18767 (N_18767,N_16165,N_16537);
nor U18768 (N_18768,N_12128,N_17989);
nor U18769 (N_18769,N_16294,N_12986);
and U18770 (N_18770,N_12661,N_17225);
xor U18771 (N_18771,N_17360,N_13656);
nand U18772 (N_18772,N_12078,N_15905);
nand U18773 (N_18773,N_17171,N_12079);
xnor U18774 (N_18774,N_17832,N_16860);
nor U18775 (N_18775,N_16471,N_15245);
nor U18776 (N_18776,N_12877,N_15998);
nand U18777 (N_18777,N_14934,N_13156);
or U18778 (N_18778,N_14775,N_15869);
nand U18779 (N_18779,N_15790,N_14338);
nor U18780 (N_18780,N_15387,N_14730);
or U18781 (N_18781,N_14428,N_15328);
or U18782 (N_18782,N_15644,N_16602);
nand U18783 (N_18783,N_12004,N_17061);
and U18784 (N_18784,N_14390,N_16266);
nor U18785 (N_18785,N_15215,N_17998);
nand U18786 (N_18786,N_13510,N_12523);
or U18787 (N_18787,N_16976,N_14952);
nand U18788 (N_18788,N_14214,N_12935);
xor U18789 (N_18789,N_12944,N_16774);
nor U18790 (N_18790,N_12549,N_14669);
and U18791 (N_18791,N_13177,N_15231);
nor U18792 (N_18792,N_12696,N_13452);
xor U18793 (N_18793,N_12857,N_13330);
nor U18794 (N_18794,N_17739,N_14381);
nand U18795 (N_18795,N_13079,N_14606);
or U18796 (N_18796,N_17332,N_15917);
nand U18797 (N_18797,N_13538,N_14854);
nor U18798 (N_18798,N_12767,N_17241);
or U18799 (N_18799,N_13891,N_13447);
nand U18800 (N_18800,N_12615,N_12198);
and U18801 (N_18801,N_14927,N_14672);
and U18802 (N_18802,N_14692,N_13947);
nor U18803 (N_18803,N_12630,N_12158);
and U18804 (N_18804,N_14590,N_14751);
or U18805 (N_18805,N_12273,N_13643);
or U18806 (N_18806,N_15910,N_17513);
and U18807 (N_18807,N_12463,N_14863);
and U18808 (N_18808,N_15369,N_13578);
nand U18809 (N_18809,N_17550,N_13431);
and U18810 (N_18810,N_15324,N_12013);
nor U18811 (N_18811,N_17281,N_17377);
nor U18812 (N_18812,N_13913,N_12803);
xor U18813 (N_18813,N_15517,N_13521);
nor U18814 (N_18814,N_15162,N_16071);
or U18815 (N_18815,N_15637,N_17076);
xnor U18816 (N_18816,N_17948,N_12923);
nor U18817 (N_18817,N_17605,N_16967);
nand U18818 (N_18818,N_13514,N_13642);
nor U18819 (N_18819,N_13567,N_15804);
nor U18820 (N_18820,N_17122,N_16933);
or U18821 (N_18821,N_16633,N_17127);
nor U18822 (N_18822,N_14588,N_15067);
nand U18823 (N_18823,N_14540,N_14226);
or U18824 (N_18824,N_14758,N_16628);
and U18825 (N_18825,N_13231,N_13801);
nand U18826 (N_18826,N_17677,N_14042);
xnor U18827 (N_18827,N_16980,N_12141);
xor U18828 (N_18828,N_17031,N_14019);
and U18829 (N_18829,N_12539,N_15724);
nand U18830 (N_18830,N_12042,N_15371);
and U18831 (N_18831,N_15228,N_17369);
nand U18832 (N_18832,N_15909,N_14635);
nor U18833 (N_18833,N_15389,N_15648);
and U18834 (N_18834,N_16843,N_17145);
or U18835 (N_18835,N_16213,N_14963);
nor U18836 (N_18836,N_15696,N_14344);
nand U18837 (N_18837,N_13412,N_14054);
nor U18838 (N_18838,N_16110,N_17946);
nand U18839 (N_18839,N_14773,N_12071);
nor U18840 (N_18840,N_15870,N_12835);
or U18841 (N_18841,N_12574,N_15033);
nand U18842 (N_18842,N_17771,N_12698);
nor U18843 (N_18843,N_14441,N_14025);
and U18844 (N_18844,N_17675,N_12821);
nand U18845 (N_18845,N_15725,N_16069);
nand U18846 (N_18846,N_14375,N_16878);
nand U18847 (N_18847,N_16833,N_15702);
nand U18848 (N_18848,N_16263,N_16469);
nand U18849 (N_18849,N_17808,N_14348);
nor U18850 (N_18850,N_13936,N_13117);
nand U18851 (N_18851,N_13366,N_15736);
or U18852 (N_18852,N_12419,N_14947);
nand U18853 (N_18853,N_16187,N_15659);
nand U18854 (N_18854,N_17765,N_15082);
or U18855 (N_18855,N_17630,N_13786);
and U18856 (N_18856,N_12023,N_17480);
or U18857 (N_18857,N_16352,N_14105);
nor U18858 (N_18858,N_15252,N_16699);
nor U18859 (N_18859,N_14200,N_17747);
nand U18860 (N_18860,N_17886,N_15104);
nand U18861 (N_18861,N_14652,N_13935);
or U18862 (N_18862,N_15717,N_14102);
or U18863 (N_18863,N_14625,N_15106);
nor U18864 (N_18864,N_16634,N_16613);
and U18865 (N_18865,N_14239,N_17650);
nor U18866 (N_18866,N_14891,N_13337);
nor U18867 (N_18867,N_13920,N_13061);
and U18868 (N_18868,N_12243,N_13889);
nand U18869 (N_18869,N_15386,N_15537);
and U18870 (N_18870,N_15177,N_13459);
or U18871 (N_18871,N_14410,N_12716);
nand U18872 (N_18872,N_13034,N_15852);
and U18873 (N_18873,N_12885,N_16900);
nand U18874 (N_18874,N_17126,N_13512);
nand U18875 (N_18875,N_12414,N_12834);
and U18876 (N_18876,N_14743,N_12290);
nor U18877 (N_18877,N_14781,N_15075);
nor U18878 (N_18878,N_13157,N_13018);
and U18879 (N_18879,N_12905,N_17621);
and U18880 (N_18880,N_12693,N_13275);
nor U18881 (N_18881,N_13979,N_14847);
nand U18882 (N_18882,N_16695,N_13151);
xnor U18883 (N_18883,N_13557,N_12903);
nand U18884 (N_18884,N_15286,N_12729);
nor U18885 (N_18885,N_14258,N_13691);
and U18886 (N_18886,N_16835,N_16893);
xnor U18887 (N_18887,N_14908,N_12999);
or U18888 (N_18888,N_13837,N_12233);
nand U18889 (N_18889,N_14148,N_15906);
or U18890 (N_18890,N_13991,N_14754);
nor U18891 (N_18891,N_17413,N_14284);
and U18892 (N_18892,N_15478,N_14597);
and U18893 (N_18893,N_12743,N_17064);
nor U18894 (N_18894,N_15824,N_12027);
or U18895 (N_18895,N_13492,N_17292);
nor U18896 (N_18896,N_14458,N_16448);
nor U18897 (N_18897,N_17243,N_12802);
nor U18898 (N_18898,N_15522,N_15035);
nand U18899 (N_18899,N_17819,N_15493);
and U18900 (N_18900,N_17222,N_16070);
and U18901 (N_18901,N_17995,N_16610);
xor U18902 (N_18902,N_16086,N_16033);
nor U18903 (N_18903,N_12520,N_15034);
or U18904 (N_18904,N_14368,N_17384);
or U18905 (N_18905,N_16177,N_13604);
or U18906 (N_18906,N_12222,N_17162);
or U18907 (N_18907,N_15908,N_14596);
nand U18908 (N_18908,N_17295,N_17729);
or U18909 (N_18909,N_15817,N_13295);
and U18910 (N_18910,N_14161,N_17376);
xor U18911 (N_18911,N_17617,N_16081);
nand U18912 (N_18912,N_15988,N_13407);
and U18913 (N_18913,N_13596,N_15586);
xnor U18914 (N_18914,N_15194,N_17319);
nor U18915 (N_18915,N_12439,N_12455);
or U18916 (N_18916,N_14082,N_13288);
nand U18917 (N_18917,N_17700,N_15746);
or U18918 (N_18918,N_12395,N_15260);
nand U18919 (N_18919,N_12762,N_12598);
or U18920 (N_18920,N_14068,N_17007);
or U18921 (N_18921,N_15339,N_17014);
or U18922 (N_18922,N_16590,N_14843);
nor U18923 (N_18923,N_17640,N_13622);
and U18924 (N_18924,N_16005,N_13008);
and U18925 (N_18925,N_16923,N_16084);
and U18926 (N_18926,N_17897,N_15617);
nor U18927 (N_18927,N_13927,N_15525);
nor U18928 (N_18928,N_15103,N_15099);
or U18929 (N_18929,N_13064,N_16583);
nor U18930 (N_18930,N_12284,N_16848);
xor U18931 (N_18931,N_14660,N_16483);
nor U18932 (N_18932,N_16270,N_16343);
nor U18933 (N_18933,N_16882,N_14993);
or U18934 (N_18934,N_17582,N_13503);
nand U18935 (N_18935,N_17471,N_17499);
xor U18936 (N_18936,N_17456,N_15271);
or U18937 (N_18937,N_12992,N_16914);
or U18938 (N_18938,N_12648,N_16280);
nor U18939 (N_18939,N_15111,N_17606);
xnor U18940 (N_18940,N_14702,N_14643);
or U18941 (N_18941,N_16178,N_16569);
or U18942 (N_18942,N_17567,N_15803);
and U18943 (N_18943,N_16214,N_15795);
and U18944 (N_18944,N_15911,N_13427);
xnor U18945 (N_18945,N_12401,N_12727);
or U18946 (N_18946,N_13626,N_14011);
nor U18947 (N_18947,N_16997,N_14736);
or U18948 (N_18948,N_13393,N_14542);
nor U18949 (N_18949,N_16326,N_17697);
or U18950 (N_18950,N_15929,N_15808);
xnor U18951 (N_18951,N_13743,N_16714);
nor U18952 (N_18952,N_14435,N_16329);
or U18953 (N_18953,N_16185,N_13343);
or U18954 (N_18954,N_15081,N_15242);
or U18955 (N_18955,N_13043,N_13432);
nand U18956 (N_18956,N_16593,N_16423);
nor U18957 (N_18957,N_14882,N_15571);
nand U18958 (N_18958,N_13073,N_17305);
nand U18959 (N_18959,N_15796,N_16335);
nor U18960 (N_18960,N_17938,N_17506);
or U18961 (N_18961,N_12397,N_12427);
nor U18962 (N_18962,N_16731,N_17223);
nand U18963 (N_18963,N_14563,N_14464);
or U18964 (N_18964,N_15687,N_16347);
or U18965 (N_18965,N_17438,N_16489);
and U18966 (N_18966,N_16660,N_12203);
or U18967 (N_18967,N_13841,N_13006);
nand U18968 (N_18968,N_14648,N_13102);
and U18969 (N_18969,N_15524,N_14580);
and U18970 (N_18970,N_15588,N_13227);
nor U18971 (N_18971,N_15381,N_16122);
or U18972 (N_18972,N_14349,N_16874);
or U18973 (N_18973,N_13145,N_12888);
nand U18974 (N_18974,N_12343,N_17502);
or U18975 (N_18975,N_15738,N_17019);
nor U18976 (N_18976,N_14601,N_12570);
nor U18977 (N_18977,N_15261,N_12702);
and U18978 (N_18978,N_16405,N_15855);
nor U18979 (N_18979,N_15408,N_12480);
and U18980 (N_18980,N_17356,N_15624);
and U18981 (N_18981,N_15255,N_13116);
and U18982 (N_18982,N_17194,N_16437);
xor U18983 (N_18983,N_16655,N_15063);
and U18984 (N_18984,N_13563,N_17731);
and U18985 (N_18985,N_16207,N_12384);
or U18986 (N_18986,N_16777,N_15384);
xor U18987 (N_18987,N_16704,N_16050);
nand U18988 (N_18988,N_12504,N_15202);
and U18989 (N_18989,N_14629,N_13119);
and U18990 (N_18990,N_14488,N_12804);
or U18991 (N_18991,N_16688,N_14649);
and U18992 (N_18992,N_14830,N_13729);
or U18993 (N_18993,N_15317,N_12645);
nor U18994 (N_18994,N_16416,N_16781);
nor U18995 (N_18995,N_13140,N_15467);
nand U18996 (N_18996,N_16021,N_12517);
xor U18997 (N_18997,N_12057,N_17341);
or U18998 (N_18998,N_12623,N_16595);
or U18999 (N_18999,N_14141,N_15353);
nand U19000 (N_19000,N_16260,N_16644);
or U19001 (N_19001,N_16810,N_16242);
xor U19002 (N_19002,N_15653,N_17408);
or U19003 (N_19003,N_17187,N_14888);
or U19004 (N_19004,N_12555,N_12040);
and U19005 (N_19005,N_16999,N_13708);
or U19006 (N_19006,N_17423,N_13420);
and U19007 (N_19007,N_13684,N_12639);
or U19008 (N_19008,N_12300,N_14159);
nor U19009 (N_19009,N_17068,N_15175);
or U19010 (N_19010,N_14201,N_13854);
or U19011 (N_19011,N_12730,N_17615);
nor U19012 (N_19012,N_16137,N_13726);
nand U19013 (N_19013,N_12981,N_16259);
or U19014 (N_19014,N_15165,N_17190);
and U19015 (N_19015,N_16007,N_17940);
or U19016 (N_19016,N_17905,N_17714);
nand U19017 (N_19017,N_17874,N_14030);
nor U19018 (N_19018,N_13258,N_14302);
nor U19019 (N_19019,N_17573,N_13766);
and U19020 (N_19020,N_15356,N_12594);
nor U19021 (N_19021,N_16204,N_15277);
xnor U19022 (N_19022,N_16723,N_15861);
or U19023 (N_19023,N_17175,N_13265);
and U19024 (N_19024,N_15853,N_13614);
and U19025 (N_19025,N_17247,N_12509);
nor U19026 (N_19026,N_14509,N_14594);
nand U19027 (N_19027,N_12192,N_12846);
nand U19028 (N_19028,N_15115,N_17317);
and U19029 (N_19029,N_13473,N_16608);
nor U19030 (N_19030,N_15388,N_15314);
nor U19031 (N_19031,N_15395,N_12037);
and U19032 (N_19032,N_13522,N_12892);
and U19033 (N_19033,N_16747,N_14617);
or U19034 (N_19034,N_17728,N_15048);
xor U19035 (N_19035,N_12058,N_15229);
nand U19036 (N_19036,N_17056,N_16247);
nand U19037 (N_19037,N_15312,N_15303);
and U19038 (N_19038,N_16194,N_14558);
nand U19039 (N_19039,N_13379,N_14408);
or U19040 (N_19040,N_17048,N_15108);
nor U19041 (N_19041,N_14725,N_17899);
and U19042 (N_19042,N_14939,N_12518);
or U19043 (N_19043,N_12135,N_13304);
and U19044 (N_19044,N_16310,N_16952);
and U19045 (N_19045,N_16460,N_15858);
nor U19046 (N_19046,N_13084,N_13755);
or U19047 (N_19047,N_15800,N_14881);
or U19048 (N_19048,N_13545,N_13971);
and U19049 (N_19049,N_16527,N_14502);
nand U19050 (N_19050,N_17654,N_17293);
and U19051 (N_19051,N_16432,N_13653);
nor U19052 (N_19052,N_13171,N_14465);
nor U19053 (N_19053,N_15453,N_14209);
xnor U19054 (N_19054,N_14905,N_12959);
or U19055 (N_19055,N_12711,N_12204);
or U19056 (N_19056,N_12546,N_14017);
and U19057 (N_19057,N_16789,N_15922);
nand U19058 (N_19058,N_12757,N_17613);
nand U19059 (N_19059,N_14031,N_17039);
or U19060 (N_19060,N_16729,N_13124);
xnor U19061 (N_19061,N_12392,N_17977);
or U19062 (N_19062,N_12776,N_14961);
or U19063 (N_19063,N_16403,N_15362);
nor U19064 (N_19064,N_17379,N_17919);
and U19065 (N_19065,N_14527,N_13807);
xor U19066 (N_19066,N_17882,N_14362);
nand U19067 (N_19067,N_14988,N_13342);
nor U19068 (N_19068,N_15938,N_17858);
or U19069 (N_19069,N_15829,N_12229);
nor U19070 (N_19070,N_17678,N_17075);
and U19071 (N_19071,N_12528,N_16589);
or U19072 (N_19072,N_12049,N_16552);
and U19073 (N_19073,N_17211,N_17246);
and U19074 (N_19074,N_14616,N_15230);
or U19075 (N_19075,N_13318,N_12920);
nand U19076 (N_19076,N_16846,N_13791);
xor U19077 (N_19077,N_17962,N_13377);
nor U19078 (N_19078,N_17842,N_12173);
nand U19079 (N_19079,N_14995,N_17828);
and U19080 (N_19080,N_16461,N_12378);
nand U19081 (N_19081,N_16473,N_17924);
xor U19082 (N_19082,N_13128,N_13152);
nand U19083 (N_19083,N_15602,N_12686);
or U19084 (N_19084,N_13044,N_16863);
or U19085 (N_19085,N_13271,N_16208);
nand U19086 (N_19086,N_15095,N_12029);
nand U19087 (N_19087,N_13436,N_15309);
and U19088 (N_19088,N_13378,N_14029);
or U19089 (N_19089,N_15211,N_15745);
nand U19090 (N_19090,N_16046,N_12360);
or U19091 (N_19091,N_17176,N_16283);
or U19092 (N_19092,N_17594,N_15979);
and U19093 (N_19093,N_12322,N_14651);
or U19094 (N_19094,N_12218,N_15330);
nand U19095 (N_19095,N_15554,N_13168);
and U19096 (N_19096,N_13607,N_17008);
and U19097 (N_19097,N_16720,N_15032);
or U19098 (N_19098,N_17534,N_17555);
and U19099 (N_19099,N_17135,N_13600);
nand U19100 (N_19100,N_15625,N_13527);
and U19101 (N_19101,N_15265,N_17776);
or U19102 (N_19102,N_14094,N_17753);
or U19103 (N_19103,N_16716,N_17608);
or U19104 (N_19104,N_14664,N_14015);
xor U19105 (N_19105,N_13321,N_17816);
nand U19106 (N_19106,N_15117,N_13507);
and U19107 (N_19107,N_14050,N_17390);
and U19108 (N_19108,N_13446,N_17957);
nor U19109 (N_19109,N_17933,N_12784);
nand U19110 (N_19110,N_15094,N_14827);
nand U19111 (N_19111,N_16685,N_16618);
nor U19112 (N_19112,N_13203,N_15753);
or U19113 (N_19113,N_12139,N_14426);
or U19114 (N_19114,N_12338,N_15865);
and U19115 (N_19115,N_17108,N_16475);
nand U19116 (N_19116,N_14519,N_13065);
or U19117 (N_19117,N_17994,N_17415);
and U19118 (N_19118,N_14874,N_14399);
nor U19119 (N_19119,N_16261,N_12774);
or U19120 (N_19120,N_14060,N_13640);
nand U19121 (N_19121,N_16267,N_14116);
or U19122 (N_19122,N_12771,N_13479);
nand U19123 (N_19123,N_13945,N_13059);
nand U19124 (N_19124,N_12453,N_15447);
nand U19125 (N_19125,N_12202,N_16034);
xnor U19126 (N_19126,N_12018,N_17197);
and U19127 (N_19127,N_15021,N_17110);
and U19128 (N_19128,N_16974,N_14204);
nor U19129 (N_19129,N_12578,N_12062);
and U19130 (N_19130,N_12377,N_16536);
nor U19131 (N_19131,N_15655,N_17624);
or U19132 (N_19132,N_14640,N_12850);
and U19133 (N_19133,N_13418,N_16960);
and U19134 (N_19134,N_14764,N_16572);
and U19135 (N_19135,N_17619,N_17482);
nor U19136 (N_19136,N_13605,N_12446);
xnor U19137 (N_19137,N_16396,N_15654);
nand U19138 (N_19138,N_14602,N_13628);
and U19139 (N_19139,N_14478,N_15442);
or U19140 (N_19140,N_12778,N_16683);
or U19141 (N_19141,N_14335,N_14760);
nand U19142 (N_19142,N_14353,N_17362);
and U19143 (N_19143,N_15772,N_14146);
or U19144 (N_19144,N_16377,N_15671);
nand U19145 (N_19145,N_12628,N_16130);
or U19146 (N_19146,N_17864,N_16322);
or U19147 (N_19147,N_14228,N_13727);
nand U19148 (N_19148,N_12442,N_15311);
xor U19149 (N_19149,N_14962,N_15848);
nor U19150 (N_19150,N_14622,N_16910);
xnor U19151 (N_19151,N_16812,N_12895);
and U19152 (N_19152,N_17854,N_13498);
and U19153 (N_19153,N_15646,N_17058);
nand U19154 (N_19154,N_17810,N_16079);
nor U19155 (N_19155,N_15840,N_15059);
nand U19156 (N_19156,N_17680,N_14978);
nor U19157 (N_19157,N_12889,N_14893);
and U19158 (N_19158,N_16508,N_16106);
nor U19159 (N_19159,N_17754,N_15712);
and U19160 (N_19160,N_14920,N_16732);
and U19161 (N_19161,N_14008,N_16361);
nor U19162 (N_19162,N_12118,N_14249);
nand U19163 (N_19163,N_13989,N_14098);
or U19164 (N_19164,N_14761,N_12385);
nand U19165 (N_19165,N_16986,N_17563);
and U19166 (N_19166,N_14694,N_15993);
nor U19167 (N_19167,N_17895,N_15217);
xnor U19168 (N_19168,N_13350,N_17931);
nor U19169 (N_19169,N_12231,N_14279);
nand U19170 (N_19170,N_17233,N_17927);
and U19171 (N_19171,N_16520,N_15011);
xor U19172 (N_19172,N_17052,N_13327);
and U19173 (N_19173,N_12724,N_14162);
nor U19174 (N_19174,N_14265,N_12798);
nand U19175 (N_19175,N_13816,N_17599);
or U19176 (N_19176,N_15291,N_15156);
or U19177 (N_19177,N_15196,N_16415);
xor U19178 (N_19178,N_14768,N_16827);
or U19179 (N_19179,N_12868,N_13715);
or U19180 (N_19180,N_17660,N_15733);
and U19181 (N_19181,N_13384,N_17693);
or U19182 (N_19182,N_15726,N_13133);
and U19183 (N_19183,N_16671,N_17845);
nand U19184 (N_19184,N_12445,N_14133);
or U19185 (N_19185,N_12982,N_17986);
nand U19186 (N_19186,N_12242,N_17040);
nand U19187 (N_19187,N_15614,N_12721);
nor U19188 (N_19188,N_16424,N_15913);
nor U19189 (N_19189,N_17807,N_12086);
or U19190 (N_19190,N_15289,N_15834);
and U19191 (N_19191,N_17658,N_12505);
nand U19192 (N_19192,N_17029,N_17308);
nand U19193 (N_19193,N_12147,N_14872);
xnor U19194 (N_19194,N_12980,N_12368);
nor U19195 (N_19195,N_14614,N_16155);
and U19196 (N_19196,N_14951,N_12246);
nand U19197 (N_19197,N_16834,N_17072);
nand U19198 (N_19198,N_15661,N_17501);
nor U19199 (N_19199,N_16324,N_13408);
and U19200 (N_19200,N_17427,N_17618);
nor U19201 (N_19201,N_12875,N_14729);
and U19202 (N_19202,N_16098,N_13165);
or U19203 (N_19203,N_15989,N_15758);
nor U19204 (N_19204,N_14361,N_13179);
nor U19205 (N_19205,N_16073,N_13056);
nand U19206 (N_19206,N_13909,N_14845);
nand U19207 (N_19207,N_12795,N_16838);
nand U19208 (N_19208,N_17604,N_13526);
xnor U19209 (N_19209,N_17556,N_12625);
nor U19210 (N_19210,N_14941,N_16947);
nor U19211 (N_19211,N_16127,N_17357);
nor U19212 (N_19212,N_16380,N_13876);
xor U19213 (N_19213,N_17189,N_12420);
nand U19214 (N_19214,N_12041,N_17505);
and U19215 (N_19215,N_17982,N_16131);
xor U19216 (N_19216,N_16728,N_13489);
or U19217 (N_19217,N_12283,N_16801);
nor U19218 (N_19218,N_15007,N_15056);
and U19219 (N_19219,N_14122,N_13574);
xnor U19220 (N_19220,N_16690,N_16531);
nor U19221 (N_19221,N_13608,N_15754);
and U19222 (N_19222,N_16354,N_14250);
nor U19223 (N_19223,N_12532,N_12742);
nor U19224 (N_19224,N_16107,N_17525);
xor U19225 (N_19225,N_13291,N_17965);
or U19226 (N_19226,N_13212,N_15703);
nor U19227 (N_19227,N_12160,N_14299);
nand U19228 (N_19228,N_16765,N_14892);
and U19229 (N_19229,N_12995,N_17460);
nor U19230 (N_19230,N_17442,N_16419);
and U19231 (N_19231,N_12148,N_12869);
xor U19232 (N_19232,N_17711,N_15027);
nor U19233 (N_19233,N_17433,N_15510);
nor U19234 (N_19234,N_16047,N_15013);
nand U19235 (N_19235,N_13737,N_14904);
or U19236 (N_19236,N_17466,N_14676);
xnor U19237 (N_19237,N_12473,N_14205);
nor U19238 (N_19238,N_14111,N_12313);
or U19239 (N_19239,N_13517,N_12418);
nand U19240 (N_19240,N_15062,N_14992);
and U19241 (N_19241,N_12731,N_15212);
nor U19242 (N_19242,N_12072,N_12220);
or U19243 (N_19243,N_16223,N_13518);
nand U19244 (N_19244,N_13689,N_14048);
and U19245 (N_19245,N_13118,N_17806);
or U19246 (N_19246,N_17418,N_13621);
nor U19247 (N_19247,N_16458,N_14316);
nor U19248 (N_19248,N_12115,N_16867);
nand U19249 (N_19249,N_14524,N_15881);
nand U19250 (N_19250,N_16866,N_13013);
and U19251 (N_19251,N_16692,N_16108);
nand U19252 (N_19252,N_16776,N_15828);
xnor U19253 (N_19253,N_15765,N_17053);
nor U19254 (N_19254,N_14687,N_15750);
and U19255 (N_19255,N_17432,N_17549);
and U19256 (N_19256,N_12601,N_13300);
nand U19257 (N_19257,N_12281,N_13471);
nor U19258 (N_19258,N_17620,N_17026);
nand U19259 (N_19259,N_14241,N_14914);
nand U19260 (N_19260,N_17133,N_16090);
xor U19261 (N_19261,N_17916,N_12394);
nand U19262 (N_19262,N_12937,N_16012);
and U19263 (N_19263,N_15530,N_13531);
or U19264 (N_19264,N_13356,N_12066);
nor U19265 (N_19265,N_16342,N_12915);
nor U19266 (N_19266,N_13277,N_14815);
nand U19267 (N_19267,N_12922,N_12732);
nand U19268 (N_19268,N_13092,N_13864);
and U19269 (N_19269,N_14838,N_17121);
and U19270 (N_19270,N_12984,N_13192);
and U19271 (N_19271,N_16824,N_15189);
nor U19272 (N_19272,N_16459,N_16638);
and U19273 (N_19273,N_12492,N_16518);
nor U19274 (N_19274,N_16712,N_15871);
xor U19275 (N_19275,N_13907,N_14079);
and U19276 (N_19276,N_15809,N_13475);
or U19277 (N_19277,N_16468,N_17918);
and U19278 (N_19278,N_12929,N_16358);
and U19279 (N_19279,N_17123,N_12607);
and U19280 (N_19280,N_15240,N_12321);
nor U19281 (N_19281,N_16546,N_13937);
nor U19282 (N_19282,N_14136,N_15679);
and U19283 (N_19283,N_14826,N_14986);
or U19284 (N_19284,N_15123,N_12813);
nor U19285 (N_19285,N_17625,N_12434);
or U19286 (N_19286,N_13466,N_14194);
or U19287 (N_19287,N_12536,N_14363);
and U19288 (N_19288,N_14984,N_17849);
and U19289 (N_19289,N_14713,N_12333);
nand U19290 (N_19290,N_17783,N_17510);
or U19291 (N_19291,N_17803,N_13147);
and U19292 (N_19292,N_12786,N_16666);
and U19293 (N_19293,N_15080,N_15088);
and U19294 (N_19294,N_15553,N_14005);
nor U19295 (N_19295,N_14714,N_13949);
and U19296 (N_19296,N_13497,N_13606);
nand U19297 (N_19297,N_13842,N_15346);
xnor U19298 (N_19298,N_14304,N_13919);
and U19299 (N_19299,N_16503,N_14623);
and U19300 (N_19300,N_12123,N_15610);
nand U19301 (N_19301,N_13762,N_12553);
nand U19302 (N_19302,N_16650,N_17515);
nand U19303 (N_19303,N_15403,N_14263);
or U19304 (N_19304,N_13855,N_13202);
or U19305 (N_19305,N_13504,N_14491);
or U19306 (N_19306,N_17494,N_12178);
nor U19307 (N_19307,N_15704,N_17479);
and U19308 (N_19308,N_16413,N_13463);
nor U19309 (N_19309,N_15374,N_12655);
and U19310 (N_19310,N_16604,N_15274);
or U19311 (N_19311,N_17579,N_15223);
or U19312 (N_19312,N_17820,N_13950);
or U19313 (N_19313,N_15462,N_12815);
or U19314 (N_19314,N_17242,N_17474);
nor U19315 (N_19315,N_15045,N_15806);
nand U19316 (N_19316,N_16648,N_17077);
nor U19317 (N_19317,N_17042,N_13575);
or U19318 (N_19318,N_12146,N_16374);
or U19319 (N_19319,N_15564,N_14215);
or U19320 (N_19320,N_14726,N_16548);
or U19321 (N_19321,N_14115,N_13783);
and U19322 (N_19322,N_12423,N_13697);
or U19323 (N_19323,N_14581,N_12272);
or U19324 (N_19324,N_17954,N_14957);
nand U19325 (N_19325,N_12753,N_14851);
or U19326 (N_19326,N_12187,N_16315);
nand U19327 (N_19327,N_12367,N_17182);
or U19328 (N_19328,N_17932,N_15645);
nor U19329 (N_19329,N_16157,N_16607);
nor U19330 (N_19330,N_13030,N_13078);
or U19331 (N_19331,N_17449,N_12489);
nor U19332 (N_19332,N_13205,N_12341);
nor U19333 (N_19333,N_12024,N_13280);
nor U19334 (N_19334,N_13364,N_15167);
xnor U19335 (N_19335,N_17334,N_12075);
and U19336 (N_19336,N_14043,N_13939);
and U19337 (N_19337,N_16238,N_16711);
and U19338 (N_19338,N_13325,N_17338);
and U19339 (N_19339,N_15737,N_17572);
and U19340 (N_19340,N_16507,N_13898);
nor U19341 (N_19341,N_14288,N_17562);
or U19342 (N_19342,N_13062,N_13946);
nor U19343 (N_19343,N_14332,N_17652);
nand U19344 (N_19344,N_17769,N_12275);
nand U19345 (N_19345,N_13057,N_12845);
or U19346 (N_19346,N_15665,N_17748);
xor U19347 (N_19347,N_17603,N_16199);
and U19348 (N_19348,N_17890,N_15984);
or U19349 (N_19349,N_14230,N_16897);
nand U19350 (N_19350,N_17311,N_15600);
xor U19351 (N_19351,N_15444,N_14545);
and U19352 (N_19352,N_14709,N_14938);
and U19353 (N_19353,N_12405,N_12854);
and U19354 (N_19354,N_14367,N_15427);
xnor U19355 (N_19355,N_15191,N_17639);
and U19356 (N_19356,N_17484,N_12325);
or U19357 (N_19357,N_16101,N_15545);
and U19358 (N_19358,N_15456,N_15147);
nor U19359 (N_19359,N_12925,N_12125);
nand U19360 (N_19360,N_15090,N_14844);
and U19361 (N_19361,N_17629,N_12270);
nor U19362 (N_19362,N_16151,N_17884);
or U19363 (N_19363,N_12383,N_16525);
and U19364 (N_19364,N_13110,N_15288);
nor U19365 (N_19365,N_15166,N_17447);
and U19366 (N_19366,N_16216,N_12502);
nand U19367 (N_19367,N_15281,N_17577);
nand U19368 (N_19368,N_14954,N_12592);
nand U19369 (N_19369,N_14805,N_17815);
or U19370 (N_19370,N_15789,N_16958);
nand U19371 (N_19371,N_17600,N_13630);
xor U19372 (N_19372,N_14365,N_13480);
nand U19373 (N_19373,N_13777,N_13230);
or U19374 (N_19374,N_12647,N_14240);
and U19375 (N_19375,N_17492,N_14466);
nand U19376 (N_19376,N_13493,N_13744);
xor U19377 (N_19377,N_16183,N_13577);
and U19378 (N_19378,N_16009,N_12706);
nand U19379 (N_19379,N_16543,N_16778);
and U19380 (N_19380,N_15508,N_12361);
nand U19381 (N_19381,N_13965,N_16401);
and U19382 (N_19382,N_14499,N_17231);
or U19383 (N_19383,N_16792,N_16681);
nand U19384 (N_19384,N_12513,N_15301);
xor U19385 (N_19385,N_12683,N_17857);
and U19386 (N_19386,N_13394,N_17702);
or U19387 (N_19387,N_16099,N_17154);
or U19388 (N_19388,N_16985,N_15139);
and U19389 (N_19389,N_16055,N_12669);
nor U19390 (N_19390,N_12745,N_17206);
nor U19391 (N_19391,N_16679,N_17219);
nand U19392 (N_19392,N_16562,N_17399);
or U19393 (N_19393,N_14842,N_16320);
or U19394 (N_19394,N_13469,N_16018);
nor U19395 (N_19395,N_17264,N_14485);
nor U19396 (N_19396,N_13075,N_13312);
or U19397 (N_19397,N_12519,N_12569);
nor U19398 (N_19398,N_16663,N_16510);
nor U19399 (N_19399,N_17092,N_14044);
and U19400 (N_19400,N_14823,N_17533);
and U19401 (N_19401,N_14712,N_12871);
and U19402 (N_19402,N_16841,N_16938);
and U19403 (N_19403,N_15030,N_15786);
nor U19404 (N_19404,N_12932,N_14237);
nor U19405 (N_19405,N_13976,N_16330);
or U19406 (N_19406,N_15573,N_15684);
xnor U19407 (N_19407,N_15634,N_16138);
nand U19408 (N_19408,N_12328,N_16301);
xnor U19409 (N_19409,N_13781,N_17151);
xnor U19410 (N_19410,N_17114,N_15020);
nor U19411 (N_19411,N_16463,N_17218);
or U19412 (N_19412,N_17458,N_13943);
nor U19413 (N_19413,N_13874,N_13033);
and U19414 (N_19414,N_13792,N_16387);
or U19415 (N_19415,N_13225,N_17607);
or U19416 (N_19416,N_17838,N_12194);
and U19417 (N_19417,N_12584,N_12606);
or U19418 (N_19418,N_16494,N_17691);
nand U19419 (N_19419,N_12955,N_16522);
and U19420 (N_19420,N_12006,N_17129);
nand U19421 (N_19421,N_12823,N_14438);
and U19422 (N_19422,N_12034,N_15345);
or U19423 (N_19423,N_12329,N_14668);
or U19424 (N_19424,N_17554,N_14742);
and U19425 (N_19425,N_14800,N_14383);
or U19426 (N_19426,N_16931,N_17467);
and U19427 (N_19427,N_14671,N_17038);
nor U19428 (N_19428,N_15101,N_13799);
nand U19429 (N_19429,N_13661,N_12640);
nor U19430 (N_19430,N_13264,N_17601);
xor U19431 (N_19431,N_14705,N_13645);
or U19432 (N_19432,N_16000,N_14956);
nand U19433 (N_19433,N_14732,N_17297);
xor U19434 (N_19434,N_17782,N_17230);
nor U19435 (N_19435,N_14084,N_14163);
nor U19436 (N_19436,N_17963,N_12291);
xor U19437 (N_19437,N_13449,N_12101);
xnor U19438 (N_19438,N_16954,N_13009);
or U19439 (N_19439,N_17214,N_13339);
or U19440 (N_19440,N_12872,N_14506);
nor U19441 (N_19441,N_15008,N_17344);
nand U19442 (N_19442,N_15837,N_14871);
or U19443 (N_19443,N_12507,N_16697);
and U19444 (N_19444,N_14523,N_14903);
nor U19445 (N_19445,N_14654,N_16478);
nand U19446 (N_19446,N_17156,N_17509);
xor U19447 (N_19447,N_16791,N_17472);
xor U19448 (N_19448,N_15907,N_12408);
xor U19449 (N_19449,N_13012,N_16594);
xor U19450 (N_19450,N_12098,N_16512);
or U19451 (N_19451,N_17333,N_17173);
and U19452 (N_19452,N_14752,N_17134);
xnor U19453 (N_19453,N_15685,N_13053);
and U19454 (N_19454,N_16752,N_12232);
and U19455 (N_19455,N_15782,N_17961);
nand U19456 (N_19456,N_13682,N_12238);
or U19457 (N_19457,N_13690,N_15232);
nand U19458 (N_19458,N_15532,N_13096);
xor U19459 (N_19459,N_15140,N_17030);
or U19460 (N_19460,N_17682,N_16397);
xor U19461 (N_19461,N_16823,N_13615);
nor U19462 (N_19462,N_16418,N_17610);
or U19463 (N_19463,N_17673,N_12737);
nand U19464 (N_19464,N_13805,N_12069);
nor U19465 (N_19465,N_16030,N_12510);
and U19466 (N_19466,N_17301,N_14463);
xnor U19467 (N_19467,N_14010,N_17060);
or U19468 (N_19468,N_14715,N_13923);
and U19469 (N_19469,N_12095,N_17679);
or U19470 (N_19470,N_17526,N_12950);
nor U19471 (N_19471,N_16466,N_13639);
xor U19472 (N_19472,N_15459,N_14686);
nor U19473 (N_19473,N_13083,N_13977);
nand U19474 (N_19474,N_15137,N_13568);
nand U19475 (N_19475,N_14274,N_13201);
nor U19476 (N_19476,N_15587,N_16755);
xnor U19477 (N_19477,N_12644,N_14846);
or U19478 (N_19478,N_12472,N_17020);
and U19479 (N_19479,N_15342,N_13144);
nor U19480 (N_19480,N_15968,N_12111);
nor U19481 (N_19481,N_13917,N_16770);
or U19482 (N_19482,N_15134,N_12881);
nand U19483 (N_19483,N_13282,N_14421);
xor U19484 (N_19484,N_17483,N_17879);
or U19485 (N_19485,N_15244,N_17238);
or U19486 (N_19486,N_12344,N_12221);
and U19487 (N_19487,N_12044,N_14092);
or U19488 (N_19488,N_15854,N_17179);
nor U19489 (N_19489,N_13335,N_17032);
or U19490 (N_19490,N_13355,N_17795);
and U19491 (N_19491,N_14189,N_14247);
nor U19492 (N_19492,N_16719,N_15373);
and U19493 (N_19493,N_16264,N_12788);
and U19494 (N_19494,N_15280,N_15734);
nand U19495 (N_19495,N_15151,N_17153);
and U19496 (N_19496,N_15351,N_16348);
nor U19497 (N_19497,N_17896,N_12136);
and U19498 (N_19498,N_16016,N_13892);
nor U19499 (N_19499,N_17569,N_17764);
and U19500 (N_19500,N_12240,N_15238);
nand U19501 (N_19501,N_13720,N_14639);
nand U19502 (N_19502,N_17787,N_13750);
nor U19503 (N_19503,N_15975,N_17833);
xor U19504 (N_19504,N_17174,N_15528);
and U19505 (N_19505,N_15543,N_15163);
and U19506 (N_19506,N_13217,N_12352);
or U19507 (N_19507,N_16232,N_16588);
nor U19508 (N_19508,N_15149,N_16963);
nor U19509 (N_19509,N_12443,N_15251);
nand U19510 (N_19510,N_12501,N_17470);
nor U19511 (N_19511,N_16586,N_15448);
nand U19512 (N_19512,N_14929,N_12310);
xor U19513 (N_19513,N_15514,N_15460);
nor U19514 (N_19514,N_14051,N_12596);
nor U19515 (N_19515,N_12312,N_17593);
xnor U19516 (N_19516,N_13825,N_15076);
nand U19517 (N_19517,N_16889,N_17406);
nor U19518 (N_19518,N_14323,N_16805);
and U19519 (N_19519,N_17756,N_17036);
nor U19520 (N_19520,N_12819,N_14906);
xor U19521 (N_19521,N_12426,N_12547);
or U19522 (N_19522,N_15895,N_14292);
or U19523 (N_19523,N_17196,N_17960);
nor U19524 (N_19524,N_17847,N_14804);
or U19525 (N_19525,N_16406,N_14925);
or U19526 (N_19526,N_12289,N_17490);
nor U19527 (N_19527,N_14061,N_17125);
nor U19528 (N_19528,N_17172,N_15841);
nand U19529 (N_19529,N_17586,N_17085);
nor U19530 (N_19530,N_16389,N_16734);
xor U19531 (N_19531,N_17841,N_16652);
or U19532 (N_19532,N_16451,N_16353);
and U19533 (N_19533,N_12259,N_12467);
nor U19534 (N_19534,N_15953,N_12810);
nor U19535 (N_19535,N_12901,N_17307);
nor U19536 (N_19536,N_14342,N_14135);
nor U19537 (N_19537,N_14883,N_13812);
and U19538 (N_19538,N_13047,N_15470);
nor U19539 (N_19539,N_15944,N_17564);
nand U19540 (N_19540,N_17762,N_14661);
and U19541 (N_19541,N_12131,N_12911);
and U19542 (N_19542,N_13579,N_16195);
nor U19543 (N_19543,N_13957,N_14000);
nand U19544 (N_19544,N_17925,N_16402);
xor U19545 (N_19545,N_15146,N_13918);
or U19546 (N_19546,N_17781,N_17137);
nand U19547 (N_19547,N_15458,N_12028);
or U19548 (N_19548,N_17539,N_14401);
and U19549 (N_19549,N_15561,N_17000);
nor U19550 (N_19550,N_13683,N_16246);
or U19551 (N_19551,N_17912,N_15801);
nor U19552 (N_19552,N_16284,N_14121);
nor U19553 (N_19553,N_17006,N_13983);
and U19554 (N_19554,N_12033,N_14091);
and U19555 (N_19555,N_14325,N_14385);
and U19556 (N_19556,N_16245,N_17518);
xor U19557 (N_19557,N_14056,N_17283);
and U19558 (N_19558,N_14379,N_17315);
or U19559 (N_19559,N_16630,N_13223);
and U19560 (N_19560,N_17372,N_16736);
xor U19561 (N_19561,N_17309,N_16308);
nand U19562 (N_19562,N_16434,N_12833);
and U19563 (N_19563,N_15970,N_17590);
and U19564 (N_19564,N_13260,N_16062);
and U19565 (N_19565,N_17469,N_13090);
nor U19566 (N_19566,N_14067,N_13546);
and U19567 (N_19567,N_12997,N_14157);
or U19568 (N_19568,N_13340,N_15144);
and U19569 (N_19569,N_13370,N_12537);
or U19570 (N_19570,N_13438,N_12918);
or U19571 (N_19571,N_15198,N_17258);
xor U19572 (N_19572,N_13206,N_14055);
xor U19573 (N_19573,N_17452,N_15357);
or U19574 (N_19574,N_14388,N_15835);
xnor U19575 (N_19575,N_17073,N_15582);
nor U19576 (N_19576,N_17348,N_14522);
xnor U19577 (N_19577,N_13131,N_17363);
nor U19578 (N_19578,N_16053,N_12280);
or U19579 (N_19579,N_15400,N_12268);
or U19580 (N_19580,N_17255,N_13213);
and U19581 (N_19581,N_15956,N_14454);
nand U19582 (N_19582,N_16312,N_15355);
and U19583 (N_19583,N_13803,N_16656);
and U19584 (N_19584,N_15950,N_16472);
or U19585 (N_19585,N_17596,N_15096);
nor U19586 (N_19586,N_14243,N_12998);
or U19587 (N_19587,N_16096,N_17718);
and U19588 (N_19588,N_15708,N_14197);
or U19589 (N_19589,N_17647,N_13719);
and U19590 (N_19590,N_12399,N_14967);
nor U19591 (N_19591,N_16133,N_17091);
nor U19592 (N_19592,N_15264,N_15065);
and U19593 (N_19593,N_13286,N_17387);
or U19594 (N_19594,N_16741,N_15557);
or U19595 (N_19595,N_16083,N_17676);
nor U19596 (N_19596,N_12151,N_13663);
nand U19597 (N_19597,N_13681,N_16528);
xnor U19598 (N_19598,N_15669,N_14520);
xor U19599 (N_19599,N_16979,N_13114);
nor U19600 (N_19600,N_15396,N_15154);
nand U19601 (N_19601,N_12544,N_16304);
and U19602 (N_19602,N_16226,N_17628);
nor U19603 (N_19603,N_12996,N_14835);
nor U19604 (N_19604,N_14254,N_15304);
nand U19605 (N_19605,N_17997,N_15497);
nand U19606 (N_19606,N_16916,N_15340);
or U19607 (N_19607,N_17069,N_17936);
and U19608 (N_19608,N_15248,N_12939);
nor U19609 (N_19609,N_13307,N_13838);
and U19610 (N_19610,N_15815,N_16257);
or U19611 (N_19611,N_17388,N_13085);
nand U19612 (N_19612,N_12000,N_17512);
nand U19613 (N_19613,N_16847,N_17591);
and U19614 (N_19614,N_15563,N_16378);
nor U19615 (N_19615,N_16093,N_15732);
and U19616 (N_19616,N_16969,N_12791);
or U19617 (N_19617,N_14297,N_15315);
and U19618 (N_19618,N_13671,N_15380);
xor U19619 (N_19619,N_13941,N_12496);
xor U19620 (N_19620,N_14538,N_15058);
nand U19621 (N_19621,N_12524,N_13877);
and U19622 (N_19622,N_12814,N_12928);
or U19623 (N_19623,N_17347,N_16793);
nand U19624 (N_19624,N_12337,N_15410);
nand U19625 (N_19625,N_16687,N_13530);
and U19626 (N_19626,N_14494,N_17383);
or U19627 (N_19627,N_17188,N_12864);
nor U19628 (N_19628,N_12305,N_13710);
nand U19629 (N_19629,N_16574,N_13938);
nand U19630 (N_19630,N_12164,N_12154);
or U19631 (N_19631,N_13831,N_16492);
nand U19632 (N_19632,N_17674,N_12177);
and U19633 (N_19633,N_13612,N_13738);
and U19634 (N_19634,N_13718,N_16545);
nor U19635 (N_19635,N_14270,N_17885);
and U19636 (N_19636,N_14149,N_13358);
nor U19637 (N_19637,N_15414,N_13488);
and U19638 (N_19638,N_12138,N_15114);
nand U19639 (N_19639,N_16297,N_14987);
nand U19640 (N_19640,N_16001,N_14424);
nand U19641 (N_19641,N_15463,N_17310);
nor U19642 (N_19642,N_16198,N_15551);
and U19643 (N_19643,N_15037,N_16385);
nand U19644 (N_19644,N_15348,N_16828);
or U19645 (N_19645,N_16911,N_12588);
or U19646 (N_19646,N_13395,N_14477);
or U19647 (N_19647,N_17130,N_17298);
nand U19648 (N_19648,N_17278,N_15972);
nor U19649 (N_19649,N_12282,N_13944);
nor U19650 (N_19650,N_14040,N_12870);
and U19651 (N_19651,N_15678,N_16597);
or U19652 (N_19652,N_13153,N_17279);
or U19653 (N_19653,N_12015,N_15812);
and U19654 (N_19654,N_12561,N_14624);
or U19655 (N_19655,N_12969,N_13494);
or U19656 (N_19656,N_17275,N_14339);
nor U19657 (N_19657,N_15762,N_14229);
nand U19658 (N_19658,N_14222,N_17701);
or U19659 (N_19659,N_12449,N_15457);
or U19660 (N_19660,N_16722,N_15689);
or U19661 (N_19661,N_17497,N_12694);
or U19662 (N_19662,N_12657,N_16779);
xor U19663 (N_19663,N_16856,N_12800);
xnor U19664 (N_19664,N_13405,N_12271);
or U19665 (N_19665,N_13014,N_12817);
nand U19666 (N_19666,N_14900,N_16068);
nand U19667 (N_19667,N_17236,N_17947);
nand U19668 (N_19668,N_12248,N_17844);
or U19669 (N_19669,N_17951,N_13707);
and U19670 (N_19670,N_12181,N_13594);
nand U19671 (N_19671,N_17583,N_14118);
and U19672 (N_19672,N_14955,N_17755);
or U19673 (N_19673,N_13551,N_17274);
nor U19674 (N_19674,N_15642,N_14020);
nor U19675 (N_19675,N_13798,N_15633);
xor U19676 (N_19676,N_16624,N_15295);
and U19677 (N_19677,N_17152,N_13706);
nand U19678 (N_19678,N_16295,N_16219);
or U19679 (N_19679,N_13435,N_17760);
and U19680 (N_19680,N_14267,N_16691);
and U19681 (N_19681,N_17522,N_13490);
nand U19682 (N_19682,N_13029,N_12975);
nand U19683 (N_19683,N_16981,N_12806);
nand U19684 (N_19684,N_17016,N_12345);
and U19685 (N_19685,N_16114,N_17641);
nor U19686 (N_19686,N_17817,N_13995);
xnor U19687 (N_19687,N_13961,N_16629);
nor U19688 (N_19688,N_15744,N_17827);
or U19689 (N_19689,N_15720,N_17303);
nand U19690 (N_19690,N_13730,N_12604);
xor U19691 (N_19691,N_14429,N_15969);
xnor U19692 (N_19692,N_13063,N_14185);
nor U19693 (N_19693,N_16425,N_16338);
and U19694 (N_19694,N_15305,N_15995);
nand U19695 (N_19695,N_13477,N_16864);
nand U19696 (N_19696,N_12633,N_13541);
or U19697 (N_19697,N_16164,N_14708);
or U19698 (N_19698,N_17136,N_13369);
and U19699 (N_19699,N_14120,N_15085);
and U19700 (N_19700,N_12897,N_15640);
or U19701 (N_19701,N_15364,N_12002);
nor U19702 (N_19702,N_13705,N_14901);
or U19703 (N_19703,N_16573,N_14167);
nor U19704 (N_19704,N_15026,N_15777);
nor U19705 (N_19705,N_13150,N_17558);
or U19706 (N_19706,N_12667,N_17860);
or U19707 (N_19707,N_15477,N_14089);
nand U19708 (N_19708,N_12085,N_16271);
nor U19709 (N_19709,N_14387,N_12045);
and U19710 (N_19710,N_16556,N_17421);
nor U19711 (N_19711,N_17244,N_14293);
nor U19712 (N_19712,N_16738,N_17686);
or U19713 (N_19713,N_15976,N_12796);
or U19714 (N_19714,N_15441,N_13052);
and U19715 (N_19715,N_15494,N_15552);
or U19716 (N_19716,N_15931,N_14828);
nand U19717 (N_19717,N_13765,N_13289);
or U19718 (N_19718,N_12156,N_17598);
and U19719 (N_19719,N_16761,N_17863);
nor U19720 (N_19720,N_14437,N_17335);
nor U19721 (N_19721,N_17904,N_17757);
nand U19722 (N_19722,N_16003,N_14607);
nor U19723 (N_19723,N_14012,N_15540);
nor U19724 (N_19724,N_15466,N_15204);
nor U19725 (N_19725,N_17322,N_16251);
nor U19726 (N_19726,N_16293,N_17521);
nand U19727 (N_19727,N_16615,N_16598);
or U19728 (N_19728,N_12410,N_12552);
nand U19729 (N_19729,N_13332,N_14731);
nand U19730 (N_19730,N_17964,N_13146);
and U19731 (N_19731,N_16567,N_16553);
or U19732 (N_19732,N_12370,N_12715);
nand U19733 (N_19733,N_12829,N_15559);
nor U19734 (N_19734,N_14675,N_14839);
nor U19735 (N_19735,N_12458,N_17034);
and U19736 (N_19736,N_13569,N_14487);
or U19737 (N_19737,N_17210,N_14561);
nor U19738 (N_19738,N_13050,N_17204);
xor U19739 (N_19739,N_14915,N_15506);
nand U19740 (N_19740,N_17240,N_17876);
or U19741 (N_19741,N_16884,N_16248);
nor U19742 (N_19742,N_12371,N_16733);
and U19743 (N_19743,N_13758,N_15479);
or U19744 (N_19744,N_14841,N_13334);
and U19745 (N_19745,N_13625,N_12257);
or U19746 (N_19746,N_15439,N_12799);
xnor U19747 (N_19747,N_16526,N_15236);
nand U19748 (N_19748,N_16118,N_12577);
nand U19749 (N_19749,N_13354,N_17286);
or U19750 (N_19750,N_16496,N_16236);
nor U19751 (N_19751,N_16849,N_13782);
nor U19752 (N_19752,N_17627,N_15660);
and U19753 (N_19753,N_17462,N_17181);
or U19754 (N_19754,N_12890,N_16132);
nor U19755 (N_19755,N_16091,N_13425);
and U19756 (N_19756,N_16727,N_12580);
nor U19757 (N_19757,N_13754,N_12535);
and U19758 (N_19758,N_15935,N_14703);
and U19759 (N_19759,N_12722,N_16676);
and U19760 (N_19760,N_16972,N_12339);
and U19761 (N_19761,N_14647,N_12011);
or U19762 (N_19762,N_15533,N_16788);
nor U19763 (N_19763,N_14657,N_12878);
or U19764 (N_19764,N_16664,N_14268);
and U19765 (N_19765,N_14740,N_15411);
nor U19766 (N_19766,N_12130,N_12265);
or U19767 (N_19767,N_15601,N_12586);
or U19768 (N_19768,N_17102,N_16564);
nand U19769 (N_19769,N_16088,N_13141);
or U19770 (N_19770,N_14108,N_13054);
xor U19771 (N_19771,N_13098,N_12979);
or U19772 (N_19772,N_16906,N_12627);
and U19773 (N_19773,N_14583,N_12977);
and U19774 (N_19774,N_14933,N_14340);
and U19775 (N_19775,N_13148,N_16363);
nor U19776 (N_19776,N_16499,N_15206);
nand U19777 (N_19777,N_13554,N_14789);
or U19778 (N_19778,N_12924,N_12916);
xnor U19779 (N_19779,N_12003,N_17093);
and U19780 (N_19780,N_13740,N_13159);
xor U19781 (N_19781,N_13178,N_13362);
nor U19782 (N_19782,N_14567,N_14354);
or U19783 (N_19783,N_16730,N_17981);
nand U19784 (N_19784,N_16961,N_14960);
nand U19785 (N_19785,N_12087,N_15916);
nand U19786 (N_19786,N_17794,N_13533);
nand U19787 (N_19787,N_16919,N_16289);
nand U19788 (N_19788,N_17656,N_12201);
or U19789 (N_19789,N_12064,N_17993);
nand U19790 (N_19790,N_15641,N_13916);
nor U19791 (N_19791,N_12254,N_16557);
xor U19792 (N_19792,N_13964,N_17911);
nor U19793 (N_19793,N_17859,N_12526);
xnor U19794 (N_19794,N_17478,N_17350);
and U19795 (N_19795,N_17703,N_12654);
nand U19796 (N_19796,N_14757,N_17320);
nor U19797 (N_19797,N_16820,N_15418);
xnor U19798 (N_19798,N_13703,N_15694);
nand U19799 (N_19799,N_14737,N_17229);
and U19800 (N_19800,N_14817,N_15596);
xnor U19801 (N_19801,N_13862,N_16558);
and U19802 (N_19802,N_13809,N_15176);
xor U19803 (N_19803,N_17868,N_14086);
or U19804 (N_19804,N_14508,N_13000);
and U19805 (N_19805,N_15728,N_13571);
nand U19806 (N_19806,N_14074,N_15578);
or U19807 (N_19807,N_15267,N_15987);
or U19808 (N_19808,N_13851,N_15259);
nand U19809 (N_19809,N_14392,N_13751);
nor U19810 (N_19810,N_12252,N_17067);
or U19811 (N_19811,N_14472,N_12100);
nand U19812 (N_19812,N_16888,N_12140);
nor U19813 (N_19813,N_16941,N_16457);
nand U19814 (N_19814,N_15978,N_12917);
nand U19815 (N_19815,N_13576,N_15756);
nor U19816 (N_19816,N_14780,N_16887);
or U19817 (N_19817,N_14140,N_12261);
nor U19818 (N_19818,N_17276,N_17435);
nand U19819 (N_19819,N_12566,N_14860);
or U19820 (N_19820,N_13692,N_16188);
nand U19821 (N_19821,N_16119,N_12573);
nand U19822 (N_19822,N_17822,N_15996);
nand U19823 (N_19823,N_15821,N_12744);
nand U19824 (N_19824,N_13840,N_16612);
xor U19825 (N_19825,N_12603,N_12635);
or U19826 (N_19826,N_12363,N_16737);
or U19827 (N_19827,N_16253,N_15670);
nand U19828 (N_19828,N_16250,N_15604);
or U19829 (N_19829,N_13281,N_15319);
nor U19830 (N_19830,N_12914,N_16797);
nor U19831 (N_19831,N_14039,N_16048);
nand U19832 (N_19832,N_16146,N_16832);
or U19833 (N_19833,N_13629,N_12288);
nand U19834 (N_19834,N_14188,N_12707);
or U19835 (N_19835,N_15390,N_16541);
and U19836 (N_19836,N_13741,N_17559);
or U19837 (N_19837,N_12219,N_14626);
and U19838 (N_19838,N_15461,N_16668);
nor U19839 (N_19839,N_13542,N_17643);
and U19840 (N_19840,N_16158,N_15180);
nor U19841 (N_19841,N_13196,N_17631);
and U19842 (N_19842,N_16398,N_16302);
or U19843 (N_19843,N_16319,N_14541);
or U19844 (N_19844,N_17124,N_14578);
xor U19845 (N_19845,N_14924,N_15334);
nor U19846 (N_19846,N_16894,N_17451);
nor U19847 (N_19847,N_13632,N_15607);
nor U19848 (N_19848,N_16785,N_16149);
or U19849 (N_19849,N_14475,N_17937);
nand U19850 (N_19850,N_13299,N_14273);
nand U19851 (N_19851,N_13261,N_14899);
xnor U19852 (N_19852,N_16909,N_14037);
nand U19853 (N_19853,N_17553,N_13496);
nand U19854 (N_19854,N_14402,N_15990);
or U19855 (N_19855,N_12658,N_15055);
nand U19856 (N_19856,N_12765,N_15422);
or U19857 (N_19857,N_13702,N_17829);
nand U19858 (N_19858,N_14735,N_12236);
and U19859 (N_19859,N_13669,N_13306);
nor U19860 (N_19860,N_13601,N_15542);
nand U19861 (N_19861,N_16056,N_17710);
xor U19862 (N_19862,N_17692,N_13963);
or U19863 (N_19863,N_16065,N_13832);
nand U19864 (N_19864,N_12206,N_12764);
or U19865 (N_19865,N_16152,N_12746);
nand U19866 (N_19866,N_12699,N_16881);
nand U19867 (N_19867,N_16113,N_13969);
nor U19868 (N_19868,N_14314,N_15866);
or U19869 (N_19869,N_12056,N_13952);
and U19870 (N_19870,N_14837,N_12841);
nand U19871 (N_19871,N_12963,N_12308);
or U19872 (N_19872,N_17473,N_12191);
nor U19873 (N_19873,N_14433,N_12738);
nand U19874 (N_19874,N_17328,N_12351);
nor U19875 (N_19875,N_14552,N_12019);
or U19876 (N_19876,N_15318,N_14001);
nand U19877 (N_19877,N_17611,N_12495);
nand U19878 (N_19878,N_12703,N_17966);
nand U19879 (N_19879,N_17683,N_12779);
nand U19880 (N_19880,N_16611,N_12359);
nand U19881 (N_19881,N_17057,N_13853);
or U19882 (N_19882,N_15619,N_13293);
xor U19883 (N_19883,N_16209,N_12840);
and U19884 (N_19884,N_16603,N_13505);
or U19885 (N_19885,N_12197,N_12217);
nor U19886 (N_19886,N_14940,N_12082);
and U19887 (N_19887,N_15195,N_16534);
and U19888 (N_19888,N_15222,N_15934);
nor U19889 (N_19889,N_13806,N_16968);
xnor U19890 (N_19890,N_14862,N_14473);
nand U19891 (N_19891,N_15536,N_16161);
nand U19892 (N_19892,N_16162,N_13863);
nor U19893 (N_19893,N_15173,N_12714);
or U19894 (N_19894,N_15489,N_13990);
and U19895 (N_19895,N_14317,N_13101);
or U19896 (N_19896,N_14869,N_17774);
nand U19897 (N_19897,N_12143,N_14683);
and U19898 (N_19898,N_13402,N_14533);
or U19899 (N_19899,N_15583,N_17059);
and U19900 (N_19900,N_13189,N_17945);
nand U19901 (N_19901,N_14573,N_15239);
nand U19902 (N_19902,N_14662,N_12830);
nor U19903 (N_19903,N_13824,N_14501);
nand U19904 (N_19904,N_13326,N_13410);
nor U19905 (N_19905,N_16317,N_13462);
and U19906 (N_19906,N_13696,N_12541);
and U19907 (N_19907,N_13487,N_15143);
xor U19908 (N_19908,N_15487,N_13817);
and U19909 (N_19909,N_14290,N_16505);
or U19910 (N_19910,N_15572,N_15015);
and U19911 (N_19911,N_13930,N_17116);
xor U19912 (N_19912,N_17699,N_13068);
and U19913 (N_19913,N_14750,N_15200);
or U19914 (N_19914,N_12438,N_13129);
and U19915 (N_19915,N_15482,N_13072);
nor U19916 (N_19916,N_17459,N_12902);
or U19917 (N_19917,N_16570,N_16540);
nor U19918 (N_19918,N_14798,N_12927);
nor U19919 (N_19919,N_17707,N_16006);
nand U19920 (N_19920,N_14922,N_15862);
or U19921 (N_19921,N_16433,N_16622);
nor U19922 (N_19922,N_15344,N_17431);
nand U19923 (N_19923,N_16877,N_13328);
xnor U19924 (N_19924,N_12976,N_13994);
and U19925 (N_19925,N_16576,N_15152);
nor U19926 (N_19926,N_17385,N_14889);
or U19927 (N_19927,N_15278,N_15889);
nand U19928 (N_19928,N_17201,N_14778);
and U19929 (N_19929,N_13609,N_15084);
nor U19930 (N_19930,N_17178,N_14295);
or U19931 (N_19931,N_17063,N_14184);
nand U19932 (N_19932,N_14816,N_13986);
or U19933 (N_19933,N_15199,N_15629);
and U19934 (N_19934,N_14719,N_16179);
and U19935 (N_19935,N_12653,N_13385);
nand U19936 (N_19936,N_17043,N_12485);
nand U19937 (N_19937,N_12797,N_16524);
nor U19938 (N_19938,N_16410,N_17375);
or U19939 (N_19939,N_15632,N_12679);
nor U19940 (N_19940,N_13502,N_16449);
nor U19941 (N_19941,N_16829,N_17528);
xor U19942 (N_19942,N_14807,N_14016);
nor U19943 (N_19943,N_12285,N_13274);
or U19944 (N_19944,N_15385,N_12216);
and U19945 (N_19945,N_17088,N_17398);
nand U19946 (N_19946,N_13654,N_12725);
nor U19947 (N_19947,N_17908,N_15269);
or U19948 (N_19948,N_16300,N_13087);
nand U19949 (N_19949,N_13002,N_16566);
nor U19950 (N_19950,N_15997,N_13220);
or U19951 (N_19951,N_12211,N_13830);
nand U19952 (N_19952,N_14155,N_16420);
nor U19953 (N_19953,N_17096,N_17645);
nand U19954 (N_19954,N_17570,N_12948);
nand U19955 (N_19955,N_12816,N_17250);
xnor U19956 (N_19956,N_17903,N_14278);
nor U19957 (N_19957,N_16698,N_15432);
and U19958 (N_19958,N_12286,N_16265);
xnor U19959 (N_19959,N_12167,N_16014);
and U19960 (N_19960,N_13736,N_17840);
and U19961 (N_19961,N_15153,N_16948);
nand U19962 (N_19962,N_14637,N_17565);
and U19963 (N_19963,N_16117,N_14861);
nand U19964 (N_19964,N_17793,N_12169);
xnor U19965 (N_19965,N_16686,N_14918);
nand U19966 (N_19966,N_15171,N_14568);
and U19967 (N_19967,N_15896,N_14532);
nand U19968 (N_19968,N_15548,N_17537);
nor U19969 (N_19969,N_14087,N_13184);
nor U19970 (N_19970,N_17234,N_14595);
and U19971 (N_19971,N_12618,N_14636);
xor U19972 (N_19972,N_16370,N_13091);
or U19973 (N_19973,N_13623,N_16482);
or U19974 (N_19974,N_15170,N_15471);
or U19975 (N_19975,N_15721,N_17544);
nor U19976 (N_19976,N_13547,N_17987);
or U19977 (N_19977,N_15575,N_13380);
nand U19978 (N_19978,N_14449,N_16212);
or U19979 (N_19979,N_17185,N_14172);
or U19980 (N_19980,N_17374,N_14334);
nor U19981 (N_19981,N_15018,N_16382);
and U19982 (N_19982,N_15436,N_17668);
nor U19983 (N_19983,N_16994,N_15367);
nand U19984 (N_19984,N_12990,N_13650);
or U19985 (N_19985,N_17200,N_15382);
nand U19986 (N_19986,N_14808,N_12938);
nor U19987 (N_19987,N_14717,N_17412);
and U19988 (N_19988,N_16477,N_13233);
nor U19989 (N_19989,N_17426,N_12503);
or U19990 (N_19990,N_16561,N_13099);
or U19991 (N_19991,N_14510,N_17409);
and U19992 (N_19992,N_13810,N_12149);
nand U19993 (N_19993,N_14492,N_13633);
and U19994 (N_19994,N_13888,N_16509);
nor U19995 (N_19995,N_16651,N_15138);
nand U19996 (N_19996,N_14026,N_14099);
nand U19997 (N_19997,N_15609,N_15093);
nand U19998 (N_19998,N_14576,N_15739);
and U19999 (N_19999,N_17050,N_12697);
nor U20000 (N_20000,N_12879,N_17690);
nor U20001 (N_20001,N_14983,N_17796);
nand U20002 (N_20002,N_14701,N_16851);
or U20003 (N_20003,N_12575,N_14977);
nand U20004 (N_20004,N_17545,N_17118);
and U20005 (N_20005,N_14747,N_12534);
xnor U20006 (N_20006,N_16581,N_14097);
and U20007 (N_20007,N_15372,N_13240);
or U20008 (N_20008,N_13802,N_13753);
nand U20009 (N_20009,N_14896,N_15125);
nand U20010 (N_20010,N_16222,N_14107);
or U20011 (N_20011,N_14980,N_12620);
nand U20012 (N_20012,N_13210,N_12326);
and U20013 (N_20013,N_13088,N_14482);
xnor U20014 (N_20014,N_13204,N_14679);
nand U20015 (N_20015,N_17584,N_15130);
nand U20016 (N_20016,N_14430,N_13843);
nand U20017 (N_20017,N_12876,N_15626);
and U20018 (N_20018,N_17405,N_16786);
and U20019 (N_20019,N_15338,N_15951);
or U20020 (N_20020,N_15899,N_17440);
or U20021 (N_20021,N_15927,N_17856);
and U20022 (N_20022,N_17094,N_16109);
or U20023 (N_20023,N_13959,N_13172);
nand U20024 (N_20024,N_12773,N_16642);
or U20025 (N_20025,N_16530,N_14831);
nor U20026 (N_20026,N_17944,N_15366);
and U20027 (N_20027,N_16182,N_17271);
nand U20028 (N_20028,N_14513,N_16742);
nand U20029 (N_20029,N_13721,N_17003);
nand U20030 (N_20030,N_14132,N_16142);
nand U20031 (N_20031,N_15354,N_13443);
and U20032 (N_20032,N_13910,N_15643);
and U20033 (N_20033,N_17391,N_14033);
or U20034 (N_20034,N_12437,N_12120);
nand U20035 (N_20035,N_13026,N_12237);
nand U20036 (N_20036,N_15491,N_17790);
and U20037 (N_20037,N_14009,N_15116);
or U20038 (N_20038,N_17217,N_13294);
or U20039 (N_20039,N_16435,N_15127);
nor U20040 (N_20040,N_13559,N_16262);
xnor U20041 (N_20041,N_15897,N_15299);
xnor U20042 (N_20042,N_12766,N_17365);
nor U20043 (N_20043,N_15237,N_16654);
or U20044 (N_20044,N_16092,N_15576);
nand U20045 (N_20045,N_14693,N_13166);
nand U20046 (N_20046,N_15379,N_12842);
or U20047 (N_20047,N_17161,N_13858);
and U20048 (N_20048,N_15615,N_17585);
nor U20049 (N_20049,N_17457,N_17732);
nor U20050 (N_20050,N_13520,N_17453);
or U20051 (N_20051,N_17958,N_14006);
nand U20052 (N_20052,N_12558,N_17698);
and U20053 (N_20053,N_14711,N_14836);
and U20054 (N_20054,N_14953,N_16966);
nand U20055 (N_20055,N_16487,N_12369);
xnor U20056 (N_20056,N_12807,N_14023);
or U20057 (N_20057,N_17330,N_14002);
or U20058 (N_20058,N_13598,N_13648);
or U20059 (N_20059,N_13248,N_14455);
or U20060 (N_20060,N_14395,N_12579);
nand U20061 (N_20061,N_16798,N_14584);
nor U20062 (N_20062,N_17893,N_12951);
nand U20063 (N_20063,N_14459,N_13872);
nand U20064 (N_20064,N_17227,N_12464);
nand U20065 (N_20065,N_16643,N_16978);
xor U20066 (N_20066,N_15041,N_17743);
or U20067 (N_20067,N_14666,N_14562);
nand U20068 (N_20068,N_14628,N_17403);
nor U20069 (N_20069,N_12491,N_15971);
and U20070 (N_20070,N_12124,N_14877);
nand U20071 (N_20071,N_14556,N_13158);
nor U20072 (N_20072,N_15397,N_14346);
and U20073 (N_20073,N_13613,N_12413);
nand U20074 (N_20074,N_13543,N_15352);
nor U20075 (N_20075,N_15958,N_14937);
or U20076 (N_20076,N_16470,N_16515);
or U20077 (N_20077,N_15499,N_16579);
nor U20078 (N_20078,N_12411,N_15207);
xor U20079 (N_20079,N_16220,N_12682);
nand U20080 (N_20080,N_12837,N_13244);
nand U20081 (N_20081,N_14850,N_14393);
and U20082 (N_20082,N_17670,N_15452);
and U20083 (N_20083,N_12287,N_15894);
xor U20084 (N_20084,N_16011,N_16373);
and U20085 (N_20085,N_12061,N_12190);
nor U20086 (N_20086,N_13058,N_12487);
xnor U20087 (N_20087,N_12417,N_16256);
or U20088 (N_20088,N_14452,N_17725);
nor U20089 (N_20089,N_16661,N_12739);
and U20090 (N_20090,N_16027,N_13191);
and U20091 (N_20091,N_14974,N_12094);
nand U20092 (N_20092,N_12324,N_14112);
nor U20093 (N_20093,N_14187,N_14296);
nor U20094 (N_20094,N_16417,N_14866);
and U20095 (N_20095,N_17735,N_13472);
nand U20096 (N_20096,N_13454,N_13955);
nand U20097 (N_20097,N_14285,N_12055);
xor U20098 (N_20098,N_12213,N_17514);
nand U20099 (N_20099,N_17894,N_16064);
nand U20100 (N_20100,N_13397,N_14227);
and U20101 (N_20101,N_15205,N_16870);
or U20102 (N_20102,N_13693,N_13484);
and U20103 (N_20103,N_17740,N_12556);
and U20104 (N_20104,N_14792,N_13246);
or U20105 (N_20105,N_14998,N_16150);
and U20106 (N_20106,N_12320,N_16939);
nand U20107 (N_20107,N_12258,N_12166);
nor U20108 (N_20108,N_12093,N_14419);
nor U20109 (N_20109,N_13338,N_14610);
nand U20110 (N_20110,N_17146,N_14638);
nand U20111 (N_20111,N_14312,N_15473);
xnor U20112 (N_20112,N_14879,N_16639);
or U20113 (N_20113,N_12589,N_12483);
nand U20114 (N_20114,N_14329,N_17935);
nor U20115 (N_20115,N_16052,N_16057);
nand U20116 (N_20116,N_16102,N_15483);
and U20117 (N_20117,N_17568,N_13121);
and U20118 (N_20118,N_12718,N_16511);
nand U20119 (N_20119,N_13028,N_15723);
and U20120 (N_20120,N_16180,N_16513);
or U20121 (N_20121,N_12900,N_12161);
or U20122 (N_20122,N_12832,N_12129);
nor U20123 (N_20123,N_12673,N_13403);
nor U20124 (N_20124,N_15052,N_16172);
nor U20125 (N_20125,N_12355,N_12304);
nor U20126 (N_20126,N_13066,N_12812);
nor U20127 (N_20127,N_13038,N_15652);
or U20128 (N_20128,N_13022,N_17380);
xor U20129 (N_20129,N_17633,N_12529);
nand U20130 (N_20130,N_12949,N_16718);
nor U20131 (N_20131,N_14440,N_13319);
nand U20132 (N_20132,N_12616,N_17846);
nand U20133 (N_20133,N_15797,N_12186);
and U20134 (N_20134,N_15991,N_14308);
nor U20135 (N_20135,N_16659,N_13027);
nor U20136 (N_20136,N_12671,N_12349);
nand U20137 (N_20137,N_16926,N_12818);
nor U20138 (N_20138,N_15857,N_17291);
nand U20139 (N_20139,N_12641,N_17687);
and U20140 (N_20140,N_12568,N_15631);
or U20141 (N_20141,N_16447,N_12188);
and U20142 (N_20142,N_16244,N_16844);
xor U20143 (N_20143,N_15347,N_15822);
or U20144 (N_20144,N_14544,N_14221);
or U20145 (N_20145,N_14313,N_17750);
nor U20146 (N_20146,N_14192,N_12624);
nor U20147 (N_20147,N_15025,N_14689);
or U20148 (N_20148,N_14530,N_12893);
or U20149 (N_20149,N_15333,N_15856);
and U20150 (N_20150,N_14667,N_15664);
and U20151 (N_20151,N_12987,N_14999);
or U20152 (N_20152,N_17866,N_12820);
nor U20153 (N_20153,N_13400,N_12297);
and U20154 (N_20154,N_16599,N_15053);
nor U20155 (N_20155,N_15562,N_17915);
nor U20156 (N_20156,N_17251,N_17713);
nor U20157 (N_20157,N_15877,N_16217);
or U20158 (N_20158,N_13667,N_15888);
and U20159 (N_20159,N_13972,N_15061);
nor U20160 (N_20160,N_12542,N_16233);
and U20161 (N_20161,N_14685,N_15150);
or U20162 (N_20162,N_16097,N_14416);
and U20163 (N_20163,N_12559,N_13882);
nor U20164 (N_20164,N_16582,N_15589);
nand U20165 (N_20165,N_17663,N_17316);
xor U20166 (N_20166,N_16049,N_13757);
xor U20167 (N_20167,N_14551,N_13619);
nor U20168 (N_20168,N_16298,N_13359);
and U20169 (N_20169,N_15994,N_17430);
or U20170 (N_20170,N_12059,N_15675);
nand U20171 (N_20171,N_14958,N_14550);
nor U20172 (N_20172,N_14912,N_14618);
nand U20173 (N_20173,N_17195,N_14225);
nor U20174 (N_20174,N_14394,N_14704);
or U20175 (N_20175,N_12612,N_15490);
or U20176 (N_20176,N_16842,N_17773);
and U20177 (N_20177,N_15365,N_15983);
or U20178 (N_20178,N_17901,N_16454);
or U20179 (N_20179,N_15518,N_15361);
and U20180 (N_20180,N_16066,N_12720);
nand U20181 (N_20181,N_14047,N_15722);
and U20182 (N_20182,N_14145,N_15087);
or U20183 (N_20183,N_13922,N_15438);
nor U20184 (N_20184,N_14156,N_12882);
nand U20185 (N_20185,N_15883,N_17887);
nand U20186 (N_20186,N_13011,N_13426);
and U20187 (N_20187,N_16498,N_17009);
or U20188 (N_20188,N_12301,N_12543);
nand U20189 (N_20189,N_14138,N_16450);
and U20190 (N_20190,N_15326,N_16023);
and U20191 (N_20191,N_14075,N_16303);
nor U20192 (N_20192,N_13259,N_12165);
and U20193 (N_20193,N_16103,N_14370);
or U20194 (N_20194,N_14633,N_16063);
and U20195 (N_20195,N_12906,N_16445);
xor U20196 (N_20196,N_13001,N_17071);
nand U20197 (N_20197,N_17653,N_14966);
nor U20198 (N_20198,N_15787,N_14566);
xnor U20199 (N_20199,N_16394,N_14034);
and U20200 (N_20200,N_12311,N_14727);
or U20201 (N_20201,N_12402,N_12052);
nand U20202 (N_20202,N_16421,N_13376);
or U20203 (N_20203,N_14427,N_17626);
nor U20204 (N_20204,N_12708,N_12582);
and U20205 (N_20205,N_15031,N_13926);
or U20206 (N_20206,N_13912,N_14434);
nand U20207 (N_20207,N_14036,N_13209);
and U20208 (N_20208,N_16171,N_12431);
xnor U20209 (N_20209,N_15672,N_16578);
nand U20210 (N_20210,N_17132,N_14982);
and U20211 (N_20211,N_12751,N_15112);
or U20212 (N_20212,N_14234,N_16120);
nor U20213 (N_20213,N_13699,N_14968);
or U20214 (N_20214,N_13175,N_15558);
nand U20215 (N_20215,N_17111,N_14403);
nand U20216 (N_20216,N_14462,N_15618);
and U20217 (N_20217,N_16273,N_12142);
xnor U20218 (N_20218,N_17340,N_15256);
or U20219 (N_20219,N_16082,N_12666);
and U20220 (N_20220,N_12331,N_15275);
and U20221 (N_20221,N_12168,N_17835);
nand U20222 (N_20222,N_16932,N_13382);
nor U20223 (N_20223,N_13869,N_13761);
and U20224 (N_20224,N_12424,N_12971);
nand U20225 (N_20225,N_16426,N_16754);
or U20226 (N_20226,N_15073,N_17079);
or U20227 (N_20227,N_17535,N_15169);
or U20228 (N_20228,N_16125,N_15526);
and U20229 (N_20229,N_12896,N_15820);
and U20230 (N_20230,N_16441,N_15832);
or U20231 (N_20231,N_13104,N_14208);
nor U20232 (N_20232,N_15268,N_16281);
and U20233 (N_20233,N_14642,N_17985);
or U20234 (N_20234,N_14849,N_17906);
or U20235 (N_20235,N_13760,N_16080);
nand U20236 (N_20236,N_12293,N_15700);
nor U20237 (N_20237,N_15880,N_17684);
or U20238 (N_20238,N_14759,N_17635);
nand U20239 (N_20239,N_14418,N_17664);
and U20240 (N_20240,N_15759,N_17239);
nor U20241 (N_20241,N_15004,N_15451);
nor U20242 (N_20242,N_17138,N_16984);
nand U20243 (N_20243,N_13219,N_14799);
and U20244 (N_20244,N_15310,N_12429);
or U20245 (N_20245,N_17485,N_17672);
or U20246 (N_20246,N_13929,N_17708);
xnor U20247 (N_20247,N_15495,N_17055);
or U20248 (N_20248,N_14634,N_12340);
and U20249 (N_20249,N_15296,N_17792);
and U20250 (N_20250,N_16759,N_13007);
or U20251 (N_20251,N_15945,N_14785);
nand U20252 (N_20252,N_16202,N_14994);
nand U20253 (N_20253,N_17768,N_17272);
or U20254 (N_20254,N_14220,N_12904);
nor U20255 (N_20255,N_13161,N_12457);
xor U20256 (N_20256,N_12172,N_15519);
nor U20257 (N_20257,N_13506,N_14834);
or U20258 (N_20258,N_15581,N_13562);
or U20259 (N_20259,N_15399,N_13160);
nor U20260 (N_20260,N_17428,N_15599);
nor U20261 (N_20261,N_15074,N_17853);
or U20262 (N_20262,N_15628,N_14244);
nand U20263 (N_20263,N_14976,N_13818);
and U20264 (N_20264,N_15565,N_13631);
nand U20265 (N_20265,N_12388,N_13901);
or U20266 (N_20266,N_12825,N_12155);
and U20267 (N_20267,N_15773,N_16762);
or U20268 (N_20268,N_13060,N_17228);
nand U20269 (N_20269,N_15698,N_12372);
or U20270 (N_20270,N_17289,N_12907);
xor U20271 (N_20271,N_16749,N_13037);
nand U20272 (N_20272,N_13942,N_15258);
and U20273 (N_20273,N_14630,N_12398);
or U20274 (N_20274,N_15054,N_15710);
xor U20275 (N_20275,N_16715,N_13951);
and U20276 (N_20276,N_16551,N_15668);
or U20277 (N_20277,N_14176,N_15203);
xnor U20278 (N_20278,N_12689,N_16782);
nor U20279 (N_20279,N_13981,N_17632);
nor U20280 (N_20280,N_16635,N_14605);
nor U20281 (N_20281,N_12267,N_12755);
xnor U20282 (N_20282,N_17080,N_17637);
nor U20283 (N_20283,N_16181,N_16993);
nand U20284 (N_20284,N_15743,N_14211);
nand U20285 (N_20285,N_14024,N_14171);
nor U20286 (N_20286,N_17476,N_15424);
nor U20287 (N_20287,N_13200,N_14359);
nor U20288 (N_20288,N_17095,N_16126);
nand U20289 (N_20289,N_17113,N_15747);
xnor U20290 (N_20290,N_15086,N_12828);
nor U20291 (N_20291,N_13183,N_15376);
or U20292 (N_20292,N_14468,N_12632);
nand U20293 (N_20293,N_16189,N_15157);
or U20294 (N_20294,N_15246,N_13881);
nor U20295 (N_20295,N_14608,N_14371);
or U20296 (N_20296,N_16990,N_15243);
or U20297 (N_20297,N_17949,N_17801);
or U20298 (N_20298,N_13857,N_14926);
nand U20299 (N_20299,N_16391,N_12662);
xnor U20300 (N_20300,N_13886,N_16956);
nor U20301 (N_20301,N_14738,N_16485);
and U20302 (N_20302,N_15504,N_14632);
nand U20303 (N_20303,N_14795,N_15711);
and U20304 (N_20304,N_15882,N_13348);
nor U20305 (N_20305,N_17914,N_16116);
or U20306 (N_20306,N_13314,N_12685);
or U20307 (N_20307,N_17705,N_16275);
or U20308 (N_20308,N_13457,N_13904);
or U20309 (N_20309,N_13887,N_17542);
nand U20310 (N_20310,N_16002,N_12048);
or U20311 (N_20311,N_14884,N_16817);
and U20312 (N_20312,N_16277,N_17715);
nor U20313 (N_20313,N_14160,N_14913);
or U20314 (N_20314,N_17926,N_17824);
or U20315 (N_20315,N_17186,N_15831);
nor U20316 (N_20316,N_13445,N_16249);
nand U20317 (N_20317,N_15069,N_12736);
or U20318 (N_20318,N_12602,N_17002);
xor U20319 (N_20319,N_17983,N_17967);
and U20320 (N_20320,N_15535,N_17321);
nor U20321 (N_20321,N_12134,N_14763);
nand U20322 (N_20322,N_13735,N_13125);
nor U20323 (N_20323,N_17546,N_16680);
or U20324 (N_20324,N_17984,N_12891);
nand U20325 (N_20325,N_14855,N_13712);
or U20326 (N_20326,N_16822,N_15662);
and U20327 (N_20327,N_17325,N_13176);
xnor U20328 (N_20328,N_16816,N_15262);
xor U20329 (N_20329,N_15620,N_16211);
nor U20330 (N_20330,N_14470,N_13962);
and U20331 (N_20331,N_14811,N_15406);
xnor U20332 (N_20332,N_16059,N_14287);
xnor U20333 (N_20333,N_16112,N_14535);
xnor U20334 (N_20334,N_16318,N_13953);
or U20335 (N_20335,N_16474,N_14959);
xor U20336 (N_20336,N_14865,N_13659);
or U20337 (N_20337,N_12357,N_16476);
nor U20338 (N_20338,N_17749,N_14555);
and U20339 (N_20339,N_17253,N_12403);
nor U20340 (N_20340,N_13368,N_15285);
or U20341 (N_20341,N_17719,N_13324);
nand U20342 (N_20342,N_12441,N_13635);
nand U20343 (N_20343,N_13441,N_16519);
and U20344 (N_20344,N_15083,N_17489);
and U20345 (N_20345,N_14445,N_12943);
or U20346 (N_20346,N_16054,N_16200);
and U20347 (N_20347,N_12262,N_14646);
and U20348 (N_20348,N_13558,N_17922);
nand U20349 (N_20349,N_17252,N_13290);
nor U20350 (N_20350,N_17943,N_13771);
nand U20351 (N_20351,N_16658,N_16678);
or U20352 (N_20352,N_14825,N_15077);
or U20353 (N_20353,N_14480,N_15449);
nor U20354 (N_20354,N_13108,N_13992);
and U20355 (N_20355,N_17105,N_13283);
nor U20356 (N_20356,N_14103,N_13474);
and U20357 (N_20357,N_12365,N_14406);
and U20358 (N_20358,N_16987,N_13311);
xnor U20359 (N_20359,N_16024,N_12700);
or U20360 (N_20360,N_13592,N_15939);
xnor U20361 (N_20361,N_17655,N_14673);
or U20362 (N_20362,N_13900,N_12183);
xnor U20363 (N_20363,N_12793,N_16584);
or U20364 (N_20364,N_12425,N_17425);
or U20365 (N_20365,N_13481,N_12985);
or U20366 (N_20366,N_12735,N_17574);
nand U20367 (N_20367,N_14165,N_16942);
or U20368 (N_20368,N_12760,N_12209);
xnor U20369 (N_20369,N_14724,N_13714);
or U20370 (N_20370,N_15507,N_16480);
xnor U20371 (N_20371,N_15874,N_12084);
or U20372 (N_20372,N_12051,N_12966);
nand U20373 (N_20373,N_13602,N_17104);
and U20374 (N_20374,N_15891,N_17651);
nor U20375 (N_20375,N_13107,N_17766);
and U20376 (N_20376,N_15066,N_12162);
or U20377 (N_20377,N_13499,N_17465);
or U20378 (N_20378,N_15440,N_15358);
nand U20379 (N_20379,N_16529,N_14142);
nor U20380 (N_20380,N_12858,N_14391);
nand U20381 (N_20381,N_13624,N_17366);
nor U20382 (N_20382,N_14688,N_17540);
or U20383 (N_20383,N_15002,N_12210);
or U20384 (N_20384,N_12109,N_15172);
nand U20385 (N_20385,N_16625,N_13588);
or U20386 (N_20386,N_12479,N_15774);
xnor U20387 (N_20387,N_13928,N_17450);
nor U20388 (N_20388,N_15693,N_17448);
or U20389 (N_20389,N_12108,N_17475);
nand U20390 (N_20390,N_12366,N_15313);
nand U20391 (N_20391,N_14973,N_16163);
and U20392 (N_20392,N_14256,N_17257);
nand U20393 (N_20393,N_13089,N_16368);
or U20394 (N_20394,N_15409,N_17027);
or U20395 (N_20395,N_17207,N_15375);
nor U20396 (N_20396,N_17974,N_16943);
nor U20397 (N_20397,N_14180,N_15683);
and U20398 (N_20398,N_16495,N_12336);
and U20399 (N_20399,N_13728,N_15937);
and U20400 (N_20400,N_15119,N_14991);
nand U20401 (N_20401,N_12506,N_14374);
nand U20402 (N_20402,N_14461,N_15181);
nor U20403 (N_20403,N_17578,N_13899);
or U20404 (N_20404,N_14684,N_13375);
or U20405 (N_20405,N_16359,N_12599);
nand U20406 (N_20406,N_12873,N_14916);
xor U20407 (N_20407,N_15197,N_12898);
xnor U20408 (N_20408,N_16964,N_17411);
nand U20409 (N_20409,N_15715,N_17744);
nand U20410 (N_20410,N_13779,N_14931);
xnor U20411 (N_20411,N_14650,N_14315);
and U20412 (N_20412,N_14812,N_12460);
or U20413 (N_20413,N_17487,N_16438);
and U20414 (N_20414,N_13652,N_17720);
and U20415 (N_20415,N_16768,N_16706);
nand U20416 (N_20416,N_14598,N_13051);
nand U20417 (N_20417,N_16831,N_16422);
and U20418 (N_20418,N_15511,N_16924);
nor U20419 (N_20419,N_17045,N_14577);
xor U20420 (N_20420,N_14022,N_12650);
or U20421 (N_20421,N_17996,N_17437);
nor U20422 (N_20422,N_13875,N_15276);
nand U20423 (N_20423,N_14756,N_15183);
nor U20424 (N_20424,N_15512,N_14787);
and U20425 (N_20425,N_13839,N_12808);
or U20426 (N_20426,N_13967,N_16852);
nor U20427 (N_20427,N_15845,N_16010);
nand U20428 (N_20428,N_13668,N_12386);
or U20429 (N_20429,N_12391,N_15893);
nor U20430 (N_20430,N_12348,N_14611);
or U20431 (N_20431,N_15680,N_13046);
nor U20432 (N_20432,N_16008,N_14665);
or U20433 (N_20433,N_15740,N_12874);
or U20434 (N_20434,N_12277,N_13973);
nand U20435 (N_20435,N_13218,N_12447);
and U20436 (N_20436,N_17589,N_14722);
nor U20437 (N_20437,N_14699,N_16170);
or U20438 (N_20438,N_12179,N_16307);
or U20439 (N_20439,N_12964,N_12691);
or U20440 (N_20440,N_16753,N_17872);
nand U20441 (N_20441,N_12076,N_15568);
nor U20442 (N_20442,N_16254,N_16381);
xnor U20443 (N_20443,N_12043,N_13421);
or U20444 (N_20444,N_14979,N_13748);
and U20445 (N_20445,N_15509,N_13482);
xnor U20446 (N_20446,N_14236,N_12404);
and U20447 (N_20447,N_13647,N_12046);
and U20448 (N_20448,N_14793,N_13272);
nand U20449 (N_20449,N_16210,N_14481);
nor U20450 (N_20450,N_15948,N_17716);
and U20451 (N_20451,N_15434,N_15638);
nor U20452 (N_20452,N_13483,N_12083);
or U20453 (N_20453,N_15516,N_12092);
xor U20454 (N_20454,N_17386,N_13746);
and U20455 (N_20455,N_13742,N_13925);
or U20456 (N_20456,N_17500,N_13688);
and U20457 (N_20457,N_13734,N_14612);
xnor U20458 (N_20458,N_17323,N_16231);
xnor U20459 (N_20459,N_15915,N_15209);
xnor U20460 (N_20460,N_13287,N_15006);
nand U20461 (N_20461,N_13317,N_17772);
nor U20462 (N_20462,N_15445,N_16408);
nand U20463 (N_20463,N_12782,N_17973);
nand U20464 (N_20464,N_14895,N_12681);
and U20465 (N_20465,N_15838,N_15498);
nand U20466 (N_20466,N_14902,N_16532);
or U20467 (N_20467,N_14517,N_15423);
nor U20468 (N_20468,N_14027,N_12249);
nand U20469 (N_20469,N_17837,N_13308);
or U20470 (N_20470,N_16067,N_17623);
and U20471 (N_20471,N_16350,N_14942);
xnor U20472 (N_20472,N_12942,N_16306);
or U20473 (N_20473,N_13017,N_14943);
nor U20474 (N_20474,N_14186,N_15730);
xnor U20475 (N_20475,N_12145,N_15368);
xnor U20476 (N_20476,N_17262,N_12687);
nand U20477 (N_20477,N_14707,N_15742);
or U20478 (N_20478,N_12538,N_14324);
or U20479 (N_20479,N_15057,N_16360);
and U20480 (N_20480,N_17910,N_15132);
nor U20481 (N_20481,N_14587,N_13931);
nand U20482 (N_20482,N_12642,N_13080);
or U20483 (N_20483,N_13434,N_13003);
nor U20484 (N_20484,N_12302,N_17414);
nor U20485 (N_20485,N_12393,N_13371);
nor U20486 (N_20486,N_14965,N_15776);
or U20487 (N_20487,N_17277,N_16290);
nand U20488 (N_20488,N_14887,N_16215);
and U20489 (N_20489,N_13440,N_14174);
nor U20490 (N_20490,N_17634,N_13903);
nor U20491 (N_20491,N_17642,N_17726);
and U20492 (N_20492,N_15579,N_12230);
and U20493 (N_20493,N_14600,N_15985);
nor U20494 (N_20494,N_17149,N_12861);
and U20495 (N_20495,N_13169,N_12974);
nand U20496 (N_20496,N_14127,N_15283);
or U20497 (N_20497,N_13914,N_14422);
and U20498 (N_20498,N_15757,N_12239);
or U20499 (N_20499,N_14856,N_13413);
nand U20500 (N_20500,N_12675,N_13788);
and U20501 (N_20501,N_14352,N_15331);
nand U20502 (N_20502,N_12001,N_16043);
and U20503 (N_20503,N_12954,N_12176);
nand U20504 (N_20504,N_16899,N_17813);
nor U20505 (N_20505,N_16032,N_14972);
nor U20506 (N_20506,N_16430,N_14129);
xnor U20507 (N_20507,N_14496,N_17723);
nand U20508 (N_20508,N_17168,N_14182);
or U20509 (N_20509,N_17159,N_13833);
xnor U20510 (N_20510,N_15647,N_14868);
nor U20511 (N_20511,N_14771,N_12740);
xnor U20512 (N_20512,N_15663,N_15219);
and U20513 (N_20513,N_15793,N_17249);
xnor U20514 (N_20514,N_13296,N_13821);
nor U20515 (N_20515,N_13303,N_12941);
and U20516 (N_20516,N_16193,N_13620);
nand U20517 (N_20517,N_17193,N_16371);
and U20518 (N_20518,N_14088,N_15775);
nand U20519 (N_20519,N_13444,N_13238);
nand U20520 (N_20520,N_15480,N_16493);
nor U20521 (N_20521,N_17368,N_14631);
or U20522 (N_20522,N_17041,N_12787);
nand U20523 (N_20523,N_13797,N_15933);
xnor U20524 (N_20524,N_15977,N_12327);
and U20525 (N_20525,N_15836,N_13120);
and U20526 (N_20526,N_16129,N_15718);
and U20527 (N_20527,N_12957,N_15502);
or U20528 (N_20528,N_12945,N_17410);
or U20529 (N_20529,N_17990,N_16399);
or U20530 (N_20530,N_13367,N_13982);
or U20531 (N_20531,N_14294,N_12486);
nor U20532 (N_20532,N_15962,N_15875);
nor U20533 (N_20533,N_16649,N_12038);
nor U20534 (N_20534,N_16601,N_15918);
or U20535 (N_20535,N_15300,N_14407);
and U20536 (N_20536,N_13135,N_17712);
xor U20537 (N_20537,N_13794,N_12934);
nor U20538 (N_20538,N_14083,N_13451);
nand U20539 (N_20539,N_14301,N_12880);
and U20540 (N_20540,N_17191,N_12754);
xor U20541 (N_20541,N_15778,N_16811);
nand U20542 (N_20542,N_17873,N_13756);
xor U20543 (N_20543,N_14479,N_12063);
xnor U20544 (N_20544,N_14653,N_15981);
or U20545 (N_20545,N_15690,N_14283);
nor U20546 (N_20546,N_13336,N_15468);
nand U20547 (N_20547,N_13590,N_14337);
and U20548 (N_20548,N_17142,N_16735);
xnor U20549 (N_20549,N_16850,N_16725);
xnor U20550 (N_20550,N_15569,N_17054);
nand U20551 (N_20551,N_13236,N_12855);
nor U20552 (N_20552,N_15019,N_17049);
or U20553 (N_20553,N_17382,N_15247);
or U20554 (N_20554,N_14766,N_13139);
nor U20555 (N_20555,N_17527,N_15254);
and U20556 (N_20556,N_13586,N_12482);
nor U20557 (N_20557,N_17270,N_13004);
xor U20558 (N_20558,N_16369,N_13552);
or U20559 (N_20559,N_15419,N_13847);
or U20560 (N_20560,N_14898,N_14989);
nor U20561 (N_20561,N_13315,N_12590);
nor U20562 (N_20562,N_15469,N_16327);
and U20563 (N_20563,N_13235,N_17812);
and U20564 (N_20564,N_16744,N_16019);
nand U20565 (N_20565,N_17044,N_14076);
or U20566 (N_20566,N_15878,N_12805);
nand U20567 (N_20567,N_12634,N_15799);
and U20568 (N_20568,N_15068,N_17208);
and U20569 (N_20569,N_14396,N_13174);
or U20570 (N_20570,N_16060,N_14531);
and U20571 (N_20571,N_17454,N_12790);
and U20572 (N_20572,N_17588,N_16592);
nor U20573 (N_20573,N_17167,N_15282);
nand U20574 (N_20574,N_17420,N_12863);
nor U20575 (N_20575,N_12610,N_15584);
and U20576 (N_20576,N_13372,N_14218);
nand U20577 (N_20577,N_17976,N_14303);
and U20578 (N_20578,N_16921,N_13199);
and U20579 (N_20579,N_17284,N_12110);
nor U20580 (N_20580,N_12651,N_12022);
and U20581 (N_20581,N_12047,N_16500);
or U20582 (N_20582,N_16854,N_13122);
nand U20583 (N_20583,N_12712,N_17862);
or U20584 (N_20584,N_15323,N_13185);
nor U20585 (N_20585,N_16560,N_16227);
or U20586 (N_20586,N_13700,N_15118);
nor U20587 (N_20587,N_12853,N_16585);
nor U20588 (N_20588,N_17798,N_16296);
or U20589 (N_20589,N_14004,N_17010);
nand U20590 (N_20590,N_16959,N_15741);
nand U20591 (N_20591,N_14078,N_15681);
or U20592 (N_20592,N_13584,N_12317);
xnor U20593 (N_20593,N_14790,N_13316);
nor U20594 (N_20594,N_17504,N_16927);
nor U20595 (N_20595,N_12318,N_14096);
or U20596 (N_20596,N_12205,N_17035);
or U20597 (N_20597,N_16388,N_17017);
and U20598 (N_20598,N_16442,N_13868);
nor U20599 (N_20599,N_17117,N_15038);
and U20600 (N_20600,N_14873,N_12886);
and U20601 (N_20601,N_15012,N_13467);
nor U20602 (N_20602,N_17296,N_17396);
or U20603 (N_20603,N_17498,N_12962);
nor U20604 (N_20604,N_16775,N_13724);
xnor U20605 (N_20605,N_13401,N_17198);
nand U20606 (N_20606,N_15220,N_14059);
nor U20607 (N_20607,N_13137,N_12794);
nand U20608 (N_20608,N_16383,N_17648);
nand U20609 (N_20609,N_13221,N_12021);
nor U20610 (N_20610,N_13082,N_17337);
nand U20611 (N_20611,N_12009,N_16673);
or U20612 (N_20612,N_14870,N_17920);
nor U20613 (N_20613,N_14769,N_16902);
and U20614 (N_20614,N_12379,N_17370);
nand U20615 (N_20615,N_15912,N_13513);
or U20616 (N_20616,N_15402,N_15394);
nor U20617 (N_20617,N_16035,N_14066);
nand U20618 (N_20618,N_16201,N_12993);
nand U20619 (N_20619,N_14603,N_15412);
nand U20620 (N_20620,N_12026,N_16707);
and U20621 (N_20621,N_14223,N_16344);
or U20622 (N_20622,N_15639,N_17164);
or U20623 (N_20623,N_14774,N_13747);
and U20624 (N_20624,N_16225,N_14659);
and U20625 (N_20625,N_17516,N_16325);
or U20626 (N_20626,N_15186,N_17602);
and U20627 (N_20627,N_16037,N_15885);
nor U20628 (N_20628,N_14166,N_13456);
xnor U20629 (N_20629,N_14537,N_14101);
or U20630 (N_20630,N_14813,N_17597);
and U20631 (N_20631,N_17992,N_16745);
nor U20632 (N_20632,N_12930,N_12704);
and U20633 (N_20633,N_16258,N_15336);
or U20634 (N_20634,N_15060,N_14093);
and U20635 (N_20635,N_13077,N_13040);
and U20636 (N_20636,N_17288,N_12769);
or U20637 (N_20637,N_16891,N_12908);
or U20638 (N_20638,N_14615,N_17548);
nand U20639 (N_20639,N_16965,N_16514);
or U20640 (N_20640,N_16871,N_17037);
and U20641 (N_20641,N_15089,N_14880);
nor U20642 (N_20642,N_14280,N_17877);
and U20643 (N_20643,N_14333,N_17889);
xnor U20644 (N_20644,N_14875,N_14755);
and U20645 (N_20645,N_17078,N_12887);
nor U20646 (N_20646,N_12988,N_13067);
nor U20647 (N_20647,N_13429,N_16085);
and U20648 (N_20648,N_13549,N_12822);
xnor U20649 (N_20649,N_14131,N_14853);
and U20650 (N_20650,N_15178,N_15705);
or U20651 (N_20651,N_14151,N_16857);
nand U20652 (N_20652,N_12292,N_12088);
nand U20653 (N_20653,N_13516,N_14490);
xnor U20654 (N_20654,N_15760,N_14235);
and U20655 (N_20655,N_12884,N_13448);
nand U20656 (N_20656,N_14057,N_17917);
nor U20657 (N_20657,N_17867,N_14126);
or U20658 (N_20658,N_16794,N_16750);
nand U20659 (N_20659,N_13025,N_15593);
or U20660 (N_20660,N_14064,N_15105);
nor U20661 (N_20661,N_13800,N_13999);
nand U20662 (N_20662,N_16502,N_15000);
and U20663 (N_20663,N_17786,N_15279);
nor U20664 (N_20664,N_14300,N_13826);
or U20665 (N_20665,N_16444,N_17758);
nand U20666 (N_20666,N_16345,N_14627);
nor U20667 (N_20667,N_15879,N_14586);
nor U20668 (N_20668,N_16386,N_17203);
or U20669 (N_20669,N_12531,N_14164);
or U20670 (N_20670,N_14351,N_13352);
and U20671 (N_20671,N_15110,N_16346);
nor U20672 (N_20672,N_15307,N_16670);
and U20673 (N_20673,N_15802,N_17439);
or U20674 (N_20674,N_14721,N_13822);
nand U20675 (N_20675,N_14219,N_12332);
nand U20676 (N_20676,N_16128,N_17416);
xnor U20677 (N_20677,N_16780,N_16462);
and U20678 (N_20678,N_14857,N_17318);
nand U20679 (N_20679,N_13879,N_16896);
nand U20680 (N_20680,N_12909,N_15253);
nand U20681 (N_20681,N_14110,N_13198);
nor U20682 (N_20682,N_16694,N_13539);
nand U20683 (N_20683,N_15886,N_12163);
nor U20684 (N_20684,N_17811,N_17373);
and U20685 (N_20685,N_16286,N_17349);
or U20686 (N_20686,N_12199,N_13422);
nor U20687 (N_20687,N_14848,N_15249);
or U20688 (N_20688,N_13958,N_15079);
nand U20689 (N_20689,N_16337,N_15920);
nor U20690 (N_20690,N_16148,N_12012);
nor U20691 (N_20691,N_13320,N_15392);
and U20692 (N_20692,N_16446,N_16905);
nand U20693 (N_20693,N_17969,N_17097);
xor U20694 (N_20694,N_12836,N_16077);
nor U20695 (N_20695,N_13310,N_12409);
xnor U20696 (N_20696,N_12465,N_17709);
or U20697 (N_20697,N_16176,N_14565);
and U20698 (N_20698,N_16748,N_15942);
nor U20699 (N_20699,N_14404,N_13019);
xnor U20700 (N_20700,N_14656,N_17141);
or U20701 (N_20701,N_15142,N_15298);
nor U20702 (N_20702,N_12400,N_12609);
or U20703 (N_20703,N_16726,N_15826);
or U20704 (N_20704,N_14525,N_12353);
nor U20705 (N_20705,N_14104,N_13273);
and U20706 (N_20706,N_16184,N_16757);
or U20707 (N_20707,N_13848,N_12565);
xor U20708 (N_20708,N_12450,N_14539);
nor U20709 (N_20709,N_17066,N_13618);
xor U20710 (N_20710,N_16339,N_16051);
or U20711 (N_20711,N_15435,N_16287);
nand U20712 (N_20712,N_14077,N_12099);
or U20713 (N_20713,N_12652,N_16568);
nand U20714 (N_20714,N_13985,N_13015);
or U20715 (N_20715,N_16124,N_12636);
nor U20716 (N_20716,N_14373,N_16237);
nand U20717 (N_20717,N_12695,N_17033);
and U20718 (N_20718,N_13660,N_13424);
and U20719 (N_20719,N_16620,N_17232);
nand U20720 (N_20720,N_16316,N_12619);
and U20721 (N_20721,N_12432,N_15677);
or U20722 (N_20722,N_15485,N_13524);
nor U20723 (N_20723,N_12469,N_14772);
nor U20724 (N_20724,N_17956,N_13461);
and U20725 (N_20725,N_13039,N_13021);
xor U20726 (N_20726,N_15492,N_14380);
and U20727 (N_20727,N_13279,N_13784);
or U20728 (N_20728,N_12466,N_15216);
and U20729 (N_20729,N_14123,N_15234);
xnor U20730 (N_20730,N_13679,N_17529);
or U20731 (N_20731,N_12581,N_14409);
and U20732 (N_20732,N_15682,N_14570);
xnor U20733 (N_20733,N_13583,N_12228);
nor U20734 (N_20734,N_15337,N_15928);
or U20735 (N_20735,N_14971,N_16355);
or U20736 (N_20736,N_16746,N_17285);
and U20737 (N_20737,N_16039,N_12688);
or U20738 (N_20738,N_13193,N_17823);
or U20739 (N_20739,N_14446,N_16865);
nand U20740 (N_20740,N_15570,N_12865);
nor U20741 (N_20741,N_16384,N_13123);
nor U20742 (N_20742,N_13285,N_15755);
nor U20743 (N_20743,N_12777,N_12412);
xnor U20744 (N_20744,N_13954,N_12106);
and U20745 (N_20745,N_15827,N_15515);
nand U20746 (N_20746,N_13453,N_15549);
and U20747 (N_20747,N_15676,N_14770);
nor U20748 (N_20748,N_12456,N_12380);
nand U20749 (N_20749,N_17657,N_17843);
and U20750 (N_20750,N_12315,N_16285);
nand U20751 (N_20751,N_12295,N_14809);
and U20752 (N_20752,N_17761,N_16988);
or U20753 (N_20753,N_17131,N_14560);
or U20754 (N_20754,N_13902,N_16632);
nand U20755 (N_20755,N_15960,N_13815);
nand U20756 (N_20756,N_15047,N_15148);
nand U20757 (N_20757,N_16949,N_15472);
and U20758 (N_20758,N_16710,N_13662);
nand U20759 (N_20759,N_17777,N_14950);
nor U20760 (N_20760,N_16596,N_15788);
nand U20761 (N_20761,N_16700,N_12031);
nand U20762 (N_20762,N_14765,N_15784);
or U20763 (N_20763,N_15014,N_17202);
or U20764 (N_20764,N_14518,N_15486);
nand U20765 (N_20765,N_15859,N_13417);
nor U20766 (N_20766,N_16819,N_13774);
xnor U20767 (N_20767,N_13709,N_13732);
and U20768 (N_20768,N_14783,N_17724);
nor U20769 (N_20769,N_13386,N_16962);
or U20770 (N_20770,N_14710,N_12481);
nand U20771 (N_20771,N_13772,N_14045);
nor U20772 (N_20772,N_17667,N_14331);
nand U20773 (N_20773,N_14242,N_14199);
or U20774 (N_20774,N_17394,N_12303);
and U20775 (N_20775,N_15092,N_13032);
nor U20776 (N_20776,N_16928,N_12583);
xor U20777 (N_20777,N_15992,N_17062);
nor U20778 (N_20778,N_16041,N_14878);
nand U20779 (N_20779,N_13770,N_13694);
nor U20780 (N_20780,N_13181,N_16484);
and U20781 (N_20781,N_13637,N_16614);
and U20782 (N_20782,N_16806,N_13536);
nor U20783 (N_20783,N_16940,N_12952);
and U20784 (N_20784,N_16721,N_12307);
and U20785 (N_20785,N_15769,N_16045);
nor U20786 (N_20786,N_16549,N_15849);
and U20787 (N_20787,N_12309,N_13948);
nor U20788 (N_20788,N_13768,N_16467);
or U20789 (N_20789,N_17576,N_12936);
or U20790 (N_20790,N_17978,N_17789);
and U20791 (N_20791,N_17971,N_15421);
nand U20792 (N_20792,N_13237,N_15454);
or U20793 (N_20793,N_15224,N_13678);
or U20794 (N_20794,N_13565,N_14062);
and U20795 (N_20795,N_14534,N_14003);
nor U20796 (N_20796,N_16025,N_15986);
nand U20797 (N_20797,N_13856,N_13878);
or U20798 (N_20798,N_14832,N_15350);
nor U20799 (N_20799,N_12081,N_17290);
nor U20800 (N_20800,N_14474,N_17184);
nand U20801 (N_20801,N_16917,N_12756);
or U20802 (N_20802,N_12224,N_15135);
nor U20803 (N_20803,N_16606,N_17150);
and U20804 (N_20804,N_15752,N_15349);
nor U20805 (N_20805,N_16647,N_14559);
xor U20806 (N_20806,N_13428,N_16538);
or U20807 (N_20807,N_14504,N_15488);
nand U20808 (N_20808,N_17336,N_14932);
xnor U20809 (N_20809,N_12444,N_15070);
nand U20810 (N_20810,N_13442,N_14080);
nand U20811 (N_20811,N_14251,N_15649);
xnor U20812 (N_20812,N_12564,N_16862);
nor U20813 (N_20813,N_15078,N_14852);
xor U20814 (N_20814,N_16950,N_14248);
nand U20815 (N_20815,N_12060,N_12626);
nand U20816 (N_20816,N_17397,N_13112);
xor U20817 (N_20817,N_14152,N_12005);
or U20818 (N_20818,N_14456,N_16015);
or U20819 (N_20819,N_15428,N_13515);
or U20820 (N_20820,N_14196,N_12459);
or U20821 (N_20821,N_12266,N_16075);
and U20822 (N_20822,N_15064,N_14124);
nor U20823 (N_20823,N_12189,N_15430);
and U20824 (N_20824,N_16022,N_12621);
xor U20825 (N_20825,N_12362,N_17775);
nor U20826 (N_20826,N_12931,N_12477);
or U20827 (N_20827,N_13322,N_12054);
nand U20828 (N_20828,N_12933,N_17115);
nand U20829 (N_20829,N_17551,N_15541);
nand U20830 (N_20830,N_12585,N_16013);
and U20831 (N_20831,N_15433,N_12114);
nand U20832 (N_20832,N_17665,N_12127);
and U20833 (N_20833,N_17342,N_15585);
xnor U20834 (N_20834,N_12319,N_14791);
and U20835 (N_20835,N_13460,N_16773);
or U20836 (N_20836,N_14572,N_13249);
or U20837 (N_20837,N_12571,N_16907);
nor U20838 (N_20838,N_12278,N_12545);
nor U20839 (N_20839,N_12713,N_16913);
and U20840 (N_20840,N_16837,N_13433);
nor U20841 (N_20841,N_16946,N_14658);
and U20842 (N_20842,N_17025,N_13093);
nand U20843 (N_20843,N_13228,N_14529);
nor U20844 (N_20844,N_17245,N_17733);
and U20845 (N_20845,N_14175,N_14858);
or U20846 (N_20846,N_16291,N_14543);
nor U20847 (N_20847,N_15860,N_13187);
and U20848 (N_20848,N_15590,N_16783);
and U20849 (N_20849,N_12656,N_13993);
nor U20850 (N_20850,N_17324,N_15924);
or U20851 (N_20851,N_14158,N_17681);
xnor U20852 (N_20852,N_12090,N_15420);
and U20853 (N_20853,N_14585,N_15391);
nor U20854 (N_20854,N_17378,N_14582);
and U20855 (N_20855,N_14944,N_17855);
or U20856 (N_20856,N_13465,N_16228);
nor U20857 (N_20857,N_17477,N_13540);
nand U20858 (N_20858,N_12649,N_13149);
and U20859 (N_20859,N_15481,N_14259);
and U20860 (N_20860,N_14143,N_14191);
and U20861 (N_20861,N_16872,N_16366);
nand U20862 (N_20862,N_17830,N_13717);
xor U20863 (N_20863,N_17955,N_12255);
xnor U20864 (N_20864,N_14232,N_13270);
nor U20865 (N_20865,N_14341,N_16617);
and U20866 (N_20866,N_13894,N_12306);
xor U20867 (N_20867,N_16362,N_13167);
or U20868 (N_20868,N_13638,N_16751);
nor U20869 (N_20869,N_12761,N_13589);
or U20870 (N_20870,N_14100,N_14777);
and U20871 (N_20871,N_12611,N_13566);
nand U20872 (N_20872,N_15044,N_12208);
or U20873 (N_20873,N_14207,N_17419);
and U20874 (N_20874,N_12824,N_12227);
and U20875 (N_20875,N_15926,N_16922);
or U20876 (N_20876,N_13932,N_14930);
nand U20877 (N_20877,N_15612,N_13846);
nand U20878 (N_20878,N_14645,N_13611);
and U20879 (N_20879,N_17361,N_12017);
nor U20880 (N_20880,N_16684,N_12591);
nor U20881 (N_20881,N_13808,N_12330);
nor U20882 (N_20882,N_12772,N_13670);
nor U20883 (N_20883,N_14840,N_12387);
xor U20884 (N_20884,N_13711,N_17799);
nor U20885 (N_20885,N_17721,N_16314);
and U20886 (N_20886,N_16328,N_14085);
xor U20887 (N_20887,N_14788,N_14744);
and U20888 (N_20888,N_12416,N_16017);
or U20889 (N_20889,N_12678,N_13357);
xor U20890 (N_20890,N_16123,N_13836);
or U20891 (N_20891,N_14321,N_14420);
and U20892 (N_20892,N_12567,N_12826);
xnor U20893 (N_20893,N_16340,N_15872);
nor U20894 (N_20894,N_12792,N_15921);
and U20895 (N_20895,N_12692,N_15785);
and U20896 (N_20896,N_14377,N_17082);
or U20897 (N_20897,N_17256,N_14021);
nand U20898 (N_20898,N_16764,N_17023);
or U20899 (N_20899,N_13844,N_13787);
nand U20900 (N_20900,N_12961,N_15233);
or U20901 (N_20901,N_16501,N_17481);
nor U20902 (N_20902,N_17538,N_13222);
nor U20903 (N_20903,N_12433,N_13416);
nand U20904 (N_20904,N_17770,N_13106);
and U20905 (N_20905,N_12668,N_17084);
and U20906 (N_20906,N_17531,N_12521);
and U20907 (N_20907,N_14113,N_17785);
or U20908 (N_20908,N_16662,N_13725);
or U20909 (N_20909,N_14128,N_14574);
nor U20910 (N_20910,N_12759,N_16890);
nand U20911 (N_20911,N_12910,N_15050);
and U20912 (N_20912,N_16665,N_13180);
xnor U20913 (N_20913,N_14183,N_16901);
nand U20914 (N_20914,N_13636,N_12862);
or U20915 (N_20915,N_14453,N_16390);
xnor U20916 (N_20916,N_13278,N_16464);
nor U20917 (N_20917,N_17646,N_16868);
or U20918 (N_20918,N_14806,N_13042);
nand U20919 (N_20919,N_17261,N_12184);
and U20920 (N_20920,N_16072,N_14493);
xor U20921 (N_20921,N_16815,N_16111);
or U20922 (N_20922,N_13672,N_16375);
or U20923 (N_20923,N_15378,N_17852);
and U20924 (N_20924,N_12462,N_13572);
xor U20925 (N_20925,N_14716,N_14198);
nor U20926 (N_20926,N_12631,N_15405);
and U20927 (N_20927,N_12970,N_17881);
or U20928 (N_20928,N_17446,N_16992);
nand U20929 (N_20929,N_17661,N_14498);
or U20930 (N_20930,N_15932,N_14203);
nand U20931 (N_20931,N_15598,N_14885);
or U20932 (N_20932,N_17930,N_16876);
nand U20933 (N_20933,N_17784,N_12091);
xor U20934 (N_20934,N_15464,N_13827);
nor U20935 (N_20935,N_15227,N_12316);
nand U20936 (N_20936,N_14095,N_12269);
nor U20937 (N_20937,N_13680,N_14620);
xnor U20938 (N_20938,N_12226,N_14272);
or U20939 (N_20939,N_13396,N_15805);
nor U20940 (N_20940,N_17530,N_17488);
and U20941 (N_20941,N_17070,N_13229);
xor U20942 (N_20942,N_15688,N_15226);
xor U20943 (N_20943,N_12436,N_16821);
nor U20944 (N_20944,N_13745,N_15450);
nand U20945 (N_20945,N_17869,N_13048);
and U20946 (N_20946,N_13232,N_16631);
nand U20947 (N_20947,N_16305,N_16409);
and U20948 (N_20948,N_17496,N_17441);
nand U20949 (N_20949,N_12548,N_12245);
nand U20950 (N_20950,N_17979,N_15814);
nor U20951 (N_20951,N_12680,N_17343);
or U20952 (N_20952,N_16912,N_13591);
nor U20953 (N_20953,N_16333,N_17254);
nand U20954 (N_20954,N_17907,N_17287);
nand U20955 (N_20955,N_15982,N_15500);
nor U20956 (N_20956,N_16020,N_16740);
and U20957 (N_20957,N_17517,N_15028);
and U20958 (N_20958,N_13834,N_12613);
xnor U20959 (N_20959,N_13764,N_16809);
or U20960 (N_20960,N_14549,N_16506);
and U20961 (N_20961,N_14641,N_15980);
nand U20962 (N_20962,N_14728,N_13644);
nand U20963 (N_20963,N_17581,N_15287);
nand U20964 (N_20964,N_13695,N_12234);
and U20965 (N_20965,N_15184,N_17818);
xor U20966 (N_20966,N_14859,N_13595);
and U20967 (N_20967,N_15417,N_14467);
nor U20968 (N_20968,N_17821,N_17939);
nor U20969 (N_20969,N_16702,N_15936);
or U20970 (N_20970,N_17424,N_13255);
xnor U20971 (N_20971,N_14181,N_13820);
xor U20972 (N_20972,N_13561,N_13997);
nor U20973 (N_20973,N_13305,N_14476);
nor U20974 (N_20974,N_12030,N_12748);
and U20975 (N_20975,N_12593,N_16983);
nor U20976 (N_20976,N_17791,N_14130);
and U20977 (N_20977,N_13867,N_17909);
and U20978 (N_20978,N_15022,N_13665);
nand U20979 (N_20979,N_13162,N_13749);
nor U20980 (N_20980,N_16977,N_15748);
nand U20981 (N_20981,N_15901,N_14372);
and U20982 (N_20982,N_12497,N_12758);
and U20983 (N_20983,N_17614,N_13866);
or U20984 (N_20984,N_13984,N_12373);
nand U20985 (N_20985,N_13823,N_17999);
xor U20986 (N_20986,N_13980,N_15846);
nand U20987 (N_20987,N_14150,N_13049);
and U20988 (N_20988,N_13519,N_12843);
or U20989 (N_20989,N_14745,N_17401);
and U20990 (N_20990,N_13134,N_13478);
or U20991 (N_20991,N_14786,N_14655);
nand U20992 (N_20992,N_12476,N_16427);
nand U20993 (N_20993,N_16282,N_17302);
or U20994 (N_20994,N_17345,N_12461);
and U20995 (N_20995,N_13685,N_13634);
nor U20996 (N_20996,N_17226,N_12435);
and U20997 (N_20997,N_12342,N_15868);
and U20998 (N_20998,N_13896,N_14035);
nor U20999 (N_20999,N_15476,N_17767);
and U21000 (N_21000,N_13802,N_16015);
or U21001 (N_21001,N_14097,N_14678);
nand U21002 (N_21002,N_14328,N_12893);
nand U21003 (N_21003,N_13706,N_13758);
or U21004 (N_21004,N_13993,N_16756);
nor U21005 (N_21005,N_12758,N_13953);
xor U21006 (N_21006,N_14594,N_17715);
nor U21007 (N_21007,N_16090,N_15074);
xnor U21008 (N_21008,N_15726,N_17713);
or U21009 (N_21009,N_14974,N_16973);
nor U21010 (N_21010,N_16915,N_16393);
and U21011 (N_21011,N_13422,N_16503);
or U21012 (N_21012,N_16708,N_16860);
xnor U21013 (N_21013,N_17391,N_15942);
xor U21014 (N_21014,N_12499,N_17182);
nand U21015 (N_21015,N_17693,N_14970);
nor U21016 (N_21016,N_14048,N_14464);
nor U21017 (N_21017,N_16565,N_12155);
or U21018 (N_21018,N_16103,N_13580);
xnor U21019 (N_21019,N_16579,N_12887);
and U21020 (N_21020,N_16549,N_17435);
nand U21021 (N_21021,N_14422,N_15874);
and U21022 (N_21022,N_17893,N_16906);
or U21023 (N_21023,N_14600,N_13569);
nand U21024 (N_21024,N_14641,N_17534);
and U21025 (N_21025,N_17168,N_13854);
and U21026 (N_21026,N_14912,N_12158);
nor U21027 (N_21027,N_12336,N_12467);
or U21028 (N_21028,N_13864,N_12255);
and U21029 (N_21029,N_15530,N_15236);
and U21030 (N_21030,N_12361,N_14332);
xor U21031 (N_21031,N_16656,N_16846);
or U21032 (N_21032,N_14829,N_12322);
nand U21033 (N_21033,N_14681,N_12501);
nor U21034 (N_21034,N_16884,N_12386);
or U21035 (N_21035,N_16974,N_17317);
or U21036 (N_21036,N_16646,N_16773);
xor U21037 (N_21037,N_14191,N_13717);
and U21038 (N_21038,N_15994,N_14581);
nor U21039 (N_21039,N_12003,N_12422);
nor U21040 (N_21040,N_16957,N_16006);
nor U21041 (N_21041,N_14371,N_17035);
and U21042 (N_21042,N_13413,N_13895);
and U21043 (N_21043,N_14979,N_12426);
or U21044 (N_21044,N_15609,N_13660);
nor U21045 (N_21045,N_13376,N_12943);
nand U21046 (N_21046,N_16383,N_15339);
nor U21047 (N_21047,N_15674,N_12411);
or U21048 (N_21048,N_14365,N_16639);
nor U21049 (N_21049,N_13581,N_12888);
or U21050 (N_21050,N_17052,N_12671);
and U21051 (N_21051,N_17394,N_16792);
nor U21052 (N_21052,N_12753,N_15205);
nand U21053 (N_21053,N_13342,N_15187);
nand U21054 (N_21054,N_12596,N_17509);
and U21055 (N_21055,N_12299,N_15701);
nor U21056 (N_21056,N_13387,N_17082);
nand U21057 (N_21057,N_15642,N_12438);
nor U21058 (N_21058,N_12241,N_17582);
nor U21059 (N_21059,N_16710,N_12928);
nor U21060 (N_21060,N_16862,N_14743);
nand U21061 (N_21061,N_13719,N_13436);
nor U21062 (N_21062,N_12966,N_17917);
or U21063 (N_21063,N_15657,N_17045);
xnor U21064 (N_21064,N_13866,N_12661);
or U21065 (N_21065,N_17741,N_17867);
nand U21066 (N_21066,N_15796,N_17864);
or U21067 (N_21067,N_13613,N_14777);
nor U21068 (N_21068,N_14190,N_14806);
nor U21069 (N_21069,N_13655,N_15169);
nand U21070 (N_21070,N_15892,N_12605);
nand U21071 (N_21071,N_16788,N_12391);
and U21072 (N_21072,N_12791,N_17190);
nand U21073 (N_21073,N_12956,N_17858);
nor U21074 (N_21074,N_17639,N_13794);
and U21075 (N_21075,N_16802,N_17054);
and U21076 (N_21076,N_12087,N_12783);
and U21077 (N_21077,N_14133,N_14319);
and U21078 (N_21078,N_15335,N_16800);
nand U21079 (N_21079,N_12606,N_13150);
and U21080 (N_21080,N_17109,N_17201);
nor U21081 (N_21081,N_12984,N_17827);
nand U21082 (N_21082,N_13241,N_13629);
or U21083 (N_21083,N_17139,N_15439);
nand U21084 (N_21084,N_16813,N_16065);
nand U21085 (N_21085,N_13384,N_15051);
nor U21086 (N_21086,N_14033,N_15891);
nor U21087 (N_21087,N_17489,N_16354);
nand U21088 (N_21088,N_13798,N_12589);
nor U21089 (N_21089,N_12980,N_17396);
or U21090 (N_21090,N_15402,N_15078);
nor U21091 (N_21091,N_15108,N_17006);
nor U21092 (N_21092,N_14707,N_14452);
and U21093 (N_21093,N_12033,N_14507);
xnor U21094 (N_21094,N_14149,N_13923);
xor U21095 (N_21095,N_15264,N_16154);
or U21096 (N_21096,N_13591,N_14842);
or U21097 (N_21097,N_15790,N_15762);
nor U21098 (N_21098,N_13427,N_12326);
xor U21099 (N_21099,N_12920,N_16322);
nor U21100 (N_21100,N_13470,N_17988);
or U21101 (N_21101,N_15358,N_14220);
or U21102 (N_21102,N_12888,N_12200);
or U21103 (N_21103,N_14353,N_17717);
nand U21104 (N_21104,N_14206,N_12280);
or U21105 (N_21105,N_16238,N_12304);
or U21106 (N_21106,N_17507,N_15882);
nor U21107 (N_21107,N_12103,N_14475);
or U21108 (N_21108,N_15158,N_13728);
xor U21109 (N_21109,N_13012,N_15142);
nor U21110 (N_21110,N_16676,N_12477);
and U21111 (N_21111,N_14939,N_13829);
or U21112 (N_21112,N_15803,N_15505);
nor U21113 (N_21113,N_17994,N_13045);
and U21114 (N_21114,N_15747,N_13777);
nand U21115 (N_21115,N_15141,N_14715);
xnor U21116 (N_21116,N_14694,N_13416);
and U21117 (N_21117,N_12111,N_17587);
and U21118 (N_21118,N_12023,N_15416);
nand U21119 (N_21119,N_12074,N_16973);
or U21120 (N_21120,N_16534,N_12280);
nand U21121 (N_21121,N_15032,N_14861);
or U21122 (N_21122,N_12569,N_13651);
and U21123 (N_21123,N_13894,N_17125);
and U21124 (N_21124,N_17053,N_15577);
nor U21125 (N_21125,N_13594,N_14259);
nor U21126 (N_21126,N_17998,N_14043);
nand U21127 (N_21127,N_15760,N_16404);
nand U21128 (N_21128,N_14706,N_16346);
nor U21129 (N_21129,N_14752,N_13933);
or U21130 (N_21130,N_13882,N_14519);
or U21131 (N_21131,N_17026,N_12091);
nor U21132 (N_21132,N_16924,N_12414);
xor U21133 (N_21133,N_13803,N_13332);
nor U21134 (N_21134,N_15379,N_12617);
and U21135 (N_21135,N_16351,N_15039);
or U21136 (N_21136,N_13494,N_13912);
nand U21137 (N_21137,N_14892,N_16092);
nand U21138 (N_21138,N_16884,N_15180);
and U21139 (N_21139,N_15672,N_14838);
and U21140 (N_21140,N_15455,N_14076);
or U21141 (N_21141,N_17842,N_15153);
or U21142 (N_21142,N_12573,N_14818);
xor U21143 (N_21143,N_17282,N_16514);
xor U21144 (N_21144,N_16456,N_13471);
and U21145 (N_21145,N_13754,N_12734);
nand U21146 (N_21146,N_14349,N_13264);
nor U21147 (N_21147,N_12415,N_16477);
or U21148 (N_21148,N_13681,N_14399);
nor U21149 (N_21149,N_15486,N_14782);
nor U21150 (N_21150,N_16547,N_12976);
and U21151 (N_21151,N_14816,N_14080);
nand U21152 (N_21152,N_13838,N_13357);
or U21153 (N_21153,N_12752,N_15033);
nor U21154 (N_21154,N_14474,N_16902);
nor U21155 (N_21155,N_16128,N_17556);
or U21156 (N_21156,N_13571,N_14754);
or U21157 (N_21157,N_17447,N_17107);
xor U21158 (N_21158,N_12655,N_16324);
nor U21159 (N_21159,N_15035,N_17941);
xnor U21160 (N_21160,N_17998,N_17579);
and U21161 (N_21161,N_12145,N_16704);
nand U21162 (N_21162,N_12881,N_14731);
xor U21163 (N_21163,N_16884,N_14958);
nand U21164 (N_21164,N_13306,N_17402);
and U21165 (N_21165,N_17756,N_17022);
xnor U21166 (N_21166,N_15654,N_15676);
and U21167 (N_21167,N_12312,N_12461);
nand U21168 (N_21168,N_14455,N_12716);
nand U21169 (N_21169,N_14223,N_14373);
nor U21170 (N_21170,N_16752,N_16479);
nand U21171 (N_21171,N_15712,N_16029);
nor U21172 (N_21172,N_15745,N_12516);
xnor U21173 (N_21173,N_15735,N_17004);
or U21174 (N_21174,N_12532,N_15041);
and U21175 (N_21175,N_13433,N_13840);
or U21176 (N_21176,N_15904,N_14732);
nand U21177 (N_21177,N_14999,N_15755);
or U21178 (N_21178,N_15050,N_14194);
xnor U21179 (N_21179,N_16191,N_15837);
nand U21180 (N_21180,N_14930,N_17719);
or U21181 (N_21181,N_16112,N_13342);
or U21182 (N_21182,N_16992,N_12853);
and U21183 (N_21183,N_12338,N_17692);
or U21184 (N_21184,N_13580,N_17467);
nor U21185 (N_21185,N_17394,N_13947);
nand U21186 (N_21186,N_17704,N_13396);
or U21187 (N_21187,N_17249,N_15666);
or U21188 (N_21188,N_12511,N_17663);
nand U21189 (N_21189,N_15122,N_14833);
and U21190 (N_21190,N_14937,N_17999);
and U21191 (N_21191,N_14031,N_14769);
or U21192 (N_21192,N_16935,N_14440);
or U21193 (N_21193,N_14727,N_14087);
nor U21194 (N_21194,N_12661,N_14658);
nor U21195 (N_21195,N_14363,N_12952);
nand U21196 (N_21196,N_13883,N_17284);
nand U21197 (N_21197,N_17677,N_12186);
xnor U21198 (N_21198,N_16867,N_17155);
and U21199 (N_21199,N_13543,N_13991);
and U21200 (N_21200,N_17697,N_12886);
or U21201 (N_21201,N_15091,N_17323);
and U21202 (N_21202,N_16481,N_13080);
nor U21203 (N_21203,N_15719,N_17742);
nand U21204 (N_21204,N_14091,N_15198);
or U21205 (N_21205,N_15660,N_15081);
or U21206 (N_21206,N_14774,N_15824);
or U21207 (N_21207,N_17710,N_15619);
nand U21208 (N_21208,N_16317,N_17447);
or U21209 (N_21209,N_12573,N_16349);
nand U21210 (N_21210,N_12940,N_17376);
or U21211 (N_21211,N_12361,N_12666);
nand U21212 (N_21212,N_17624,N_13964);
and U21213 (N_21213,N_16924,N_15836);
and U21214 (N_21214,N_13078,N_14956);
nor U21215 (N_21215,N_15073,N_13607);
nor U21216 (N_21216,N_16095,N_15624);
nor U21217 (N_21217,N_13670,N_14091);
nor U21218 (N_21218,N_17360,N_14654);
or U21219 (N_21219,N_13426,N_17747);
or U21220 (N_21220,N_16971,N_14510);
and U21221 (N_21221,N_12909,N_12741);
nand U21222 (N_21222,N_16140,N_13700);
nand U21223 (N_21223,N_16286,N_14575);
nor U21224 (N_21224,N_12765,N_17366);
nand U21225 (N_21225,N_15744,N_13084);
or U21226 (N_21226,N_12124,N_14767);
nand U21227 (N_21227,N_16053,N_15198);
or U21228 (N_21228,N_16692,N_17219);
or U21229 (N_21229,N_16633,N_16405);
or U21230 (N_21230,N_17174,N_16878);
xor U21231 (N_21231,N_14208,N_13706);
xor U21232 (N_21232,N_16031,N_14786);
nand U21233 (N_21233,N_16764,N_13817);
xnor U21234 (N_21234,N_14120,N_12552);
nand U21235 (N_21235,N_15054,N_15900);
nand U21236 (N_21236,N_12352,N_13407);
and U21237 (N_21237,N_16197,N_15058);
nand U21238 (N_21238,N_13554,N_14661);
or U21239 (N_21239,N_16389,N_13218);
xor U21240 (N_21240,N_15426,N_16139);
xnor U21241 (N_21241,N_15629,N_16964);
nand U21242 (N_21242,N_12485,N_13175);
nand U21243 (N_21243,N_12602,N_17103);
or U21244 (N_21244,N_15207,N_13700);
and U21245 (N_21245,N_14968,N_12396);
xor U21246 (N_21246,N_14824,N_17066);
and U21247 (N_21247,N_12614,N_17410);
nor U21248 (N_21248,N_13068,N_13211);
nand U21249 (N_21249,N_14662,N_12741);
or U21250 (N_21250,N_14066,N_17070);
nand U21251 (N_21251,N_15783,N_15231);
nand U21252 (N_21252,N_17906,N_15766);
and U21253 (N_21253,N_14597,N_14144);
or U21254 (N_21254,N_14269,N_12531);
or U21255 (N_21255,N_13692,N_13604);
and U21256 (N_21256,N_16168,N_12723);
or U21257 (N_21257,N_12538,N_13103);
nand U21258 (N_21258,N_16553,N_12223);
nand U21259 (N_21259,N_16287,N_14873);
and U21260 (N_21260,N_15678,N_17906);
and U21261 (N_21261,N_13599,N_15441);
and U21262 (N_21262,N_14883,N_17820);
and U21263 (N_21263,N_13027,N_17294);
nor U21264 (N_21264,N_15655,N_15949);
or U21265 (N_21265,N_14586,N_14716);
and U21266 (N_21266,N_16976,N_12684);
or U21267 (N_21267,N_13081,N_15511);
nand U21268 (N_21268,N_16140,N_12032);
nand U21269 (N_21269,N_16909,N_16299);
and U21270 (N_21270,N_12058,N_12540);
or U21271 (N_21271,N_14346,N_14979);
nor U21272 (N_21272,N_17673,N_12437);
nand U21273 (N_21273,N_16568,N_15089);
nand U21274 (N_21274,N_12263,N_17547);
nand U21275 (N_21275,N_15857,N_16434);
and U21276 (N_21276,N_13000,N_16648);
and U21277 (N_21277,N_13501,N_16118);
nand U21278 (N_21278,N_15837,N_17650);
xnor U21279 (N_21279,N_17622,N_15674);
and U21280 (N_21280,N_12782,N_12750);
or U21281 (N_21281,N_12714,N_13234);
xor U21282 (N_21282,N_13546,N_14775);
nor U21283 (N_21283,N_14891,N_13667);
and U21284 (N_21284,N_12417,N_14824);
nor U21285 (N_21285,N_15672,N_15373);
and U21286 (N_21286,N_13556,N_14183);
or U21287 (N_21287,N_12462,N_14833);
or U21288 (N_21288,N_13472,N_12836);
nand U21289 (N_21289,N_12741,N_16999);
and U21290 (N_21290,N_16256,N_13114);
nor U21291 (N_21291,N_13044,N_14170);
nor U21292 (N_21292,N_13147,N_12508);
nor U21293 (N_21293,N_16955,N_14978);
nor U21294 (N_21294,N_14632,N_16661);
and U21295 (N_21295,N_14572,N_12791);
or U21296 (N_21296,N_14488,N_13912);
xor U21297 (N_21297,N_12727,N_15768);
or U21298 (N_21298,N_13633,N_15133);
and U21299 (N_21299,N_12360,N_14187);
or U21300 (N_21300,N_14250,N_13815);
nor U21301 (N_21301,N_13858,N_13413);
or U21302 (N_21302,N_16423,N_17490);
nand U21303 (N_21303,N_13724,N_15729);
or U21304 (N_21304,N_12800,N_15948);
xor U21305 (N_21305,N_17273,N_13945);
or U21306 (N_21306,N_15310,N_13038);
nor U21307 (N_21307,N_14024,N_17259);
nor U21308 (N_21308,N_13306,N_16187);
nor U21309 (N_21309,N_16143,N_14727);
or U21310 (N_21310,N_13024,N_16509);
nand U21311 (N_21311,N_17230,N_13356);
and U21312 (N_21312,N_16923,N_14903);
nor U21313 (N_21313,N_13981,N_17904);
nand U21314 (N_21314,N_16337,N_17652);
xnor U21315 (N_21315,N_14814,N_17076);
or U21316 (N_21316,N_13801,N_16388);
nor U21317 (N_21317,N_15362,N_14322);
nor U21318 (N_21318,N_12581,N_16447);
xor U21319 (N_21319,N_12811,N_13464);
nand U21320 (N_21320,N_12927,N_16806);
and U21321 (N_21321,N_17648,N_15182);
xor U21322 (N_21322,N_12158,N_14179);
and U21323 (N_21323,N_16289,N_14395);
and U21324 (N_21324,N_16357,N_14742);
or U21325 (N_21325,N_16983,N_17220);
or U21326 (N_21326,N_13118,N_13559);
nor U21327 (N_21327,N_16285,N_17762);
xor U21328 (N_21328,N_15039,N_13113);
xnor U21329 (N_21329,N_17383,N_15143);
nor U21330 (N_21330,N_15338,N_16556);
nor U21331 (N_21331,N_15113,N_16746);
and U21332 (N_21332,N_14379,N_12116);
nand U21333 (N_21333,N_12527,N_14030);
nand U21334 (N_21334,N_12699,N_14446);
xnor U21335 (N_21335,N_13445,N_15078);
xor U21336 (N_21336,N_14845,N_13771);
or U21337 (N_21337,N_12047,N_13144);
and U21338 (N_21338,N_16669,N_14733);
nor U21339 (N_21339,N_15521,N_12884);
nand U21340 (N_21340,N_15107,N_16373);
or U21341 (N_21341,N_15699,N_14594);
and U21342 (N_21342,N_17058,N_15619);
or U21343 (N_21343,N_12905,N_14814);
nand U21344 (N_21344,N_15390,N_15615);
and U21345 (N_21345,N_13529,N_13837);
nor U21346 (N_21346,N_15470,N_16159);
nor U21347 (N_21347,N_17434,N_16397);
and U21348 (N_21348,N_13873,N_15781);
or U21349 (N_21349,N_16346,N_15499);
nand U21350 (N_21350,N_17620,N_15826);
xnor U21351 (N_21351,N_15040,N_14195);
nor U21352 (N_21352,N_15480,N_17161);
nand U21353 (N_21353,N_17647,N_15581);
and U21354 (N_21354,N_12008,N_15213);
nand U21355 (N_21355,N_16695,N_16180);
nor U21356 (N_21356,N_12956,N_12456);
nand U21357 (N_21357,N_15145,N_13117);
or U21358 (N_21358,N_16686,N_15414);
xnor U21359 (N_21359,N_14143,N_12957);
nand U21360 (N_21360,N_12523,N_15528);
or U21361 (N_21361,N_12939,N_17306);
xor U21362 (N_21362,N_12929,N_14134);
nand U21363 (N_21363,N_15822,N_13768);
and U21364 (N_21364,N_16562,N_12952);
and U21365 (N_21365,N_13295,N_16095);
or U21366 (N_21366,N_13954,N_15361);
nand U21367 (N_21367,N_14134,N_13187);
xnor U21368 (N_21368,N_15177,N_12570);
nand U21369 (N_21369,N_12744,N_14828);
xor U21370 (N_21370,N_13796,N_15338);
nand U21371 (N_21371,N_13241,N_17315);
nor U21372 (N_21372,N_13231,N_14628);
nor U21373 (N_21373,N_12710,N_16241);
and U21374 (N_21374,N_12870,N_14007);
and U21375 (N_21375,N_16545,N_12328);
or U21376 (N_21376,N_16275,N_12556);
nor U21377 (N_21377,N_17709,N_15925);
nor U21378 (N_21378,N_16481,N_16341);
xor U21379 (N_21379,N_15060,N_17340);
nor U21380 (N_21380,N_17136,N_12634);
or U21381 (N_21381,N_15525,N_14017);
nand U21382 (N_21382,N_14294,N_13049);
xor U21383 (N_21383,N_17087,N_12260);
or U21384 (N_21384,N_13146,N_15463);
nor U21385 (N_21385,N_15105,N_14195);
nor U21386 (N_21386,N_13615,N_16936);
nand U21387 (N_21387,N_14733,N_17787);
and U21388 (N_21388,N_16263,N_12388);
nor U21389 (N_21389,N_15553,N_14918);
nand U21390 (N_21390,N_17296,N_16082);
xor U21391 (N_21391,N_17632,N_15085);
or U21392 (N_21392,N_14443,N_15748);
nor U21393 (N_21393,N_12791,N_17007);
nor U21394 (N_21394,N_15667,N_15911);
and U21395 (N_21395,N_14418,N_13626);
and U21396 (N_21396,N_13935,N_12922);
nand U21397 (N_21397,N_13362,N_16673);
and U21398 (N_21398,N_15036,N_12514);
nand U21399 (N_21399,N_12179,N_17222);
nor U21400 (N_21400,N_13186,N_16643);
nor U21401 (N_21401,N_16748,N_12087);
nor U21402 (N_21402,N_13933,N_14897);
and U21403 (N_21403,N_12852,N_16460);
and U21404 (N_21404,N_12771,N_17026);
or U21405 (N_21405,N_15854,N_12014);
nor U21406 (N_21406,N_13716,N_16146);
nand U21407 (N_21407,N_14921,N_16021);
or U21408 (N_21408,N_12562,N_15278);
xnor U21409 (N_21409,N_17375,N_14435);
xnor U21410 (N_21410,N_15781,N_15833);
nand U21411 (N_21411,N_12624,N_13232);
or U21412 (N_21412,N_12246,N_15230);
xnor U21413 (N_21413,N_14297,N_12896);
xor U21414 (N_21414,N_15887,N_15234);
nand U21415 (N_21415,N_16395,N_13231);
nor U21416 (N_21416,N_16637,N_14871);
and U21417 (N_21417,N_13317,N_13413);
nand U21418 (N_21418,N_15688,N_14807);
or U21419 (N_21419,N_12091,N_12122);
xor U21420 (N_21420,N_16534,N_14078);
nand U21421 (N_21421,N_12932,N_16267);
and U21422 (N_21422,N_12797,N_14150);
nor U21423 (N_21423,N_12615,N_14299);
or U21424 (N_21424,N_14228,N_15522);
or U21425 (N_21425,N_15496,N_16421);
xor U21426 (N_21426,N_14905,N_15588);
or U21427 (N_21427,N_13113,N_15255);
nor U21428 (N_21428,N_13477,N_17442);
and U21429 (N_21429,N_13451,N_13092);
nor U21430 (N_21430,N_12139,N_12786);
and U21431 (N_21431,N_17160,N_17657);
and U21432 (N_21432,N_16501,N_14162);
or U21433 (N_21433,N_14723,N_13498);
or U21434 (N_21434,N_12183,N_14950);
or U21435 (N_21435,N_17368,N_16094);
or U21436 (N_21436,N_14041,N_15530);
nand U21437 (N_21437,N_15629,N_17278);
nand U21438 (N_21438,N_12486,N_17186);
nand U21439 (N_21439,N_16025,N_13485);
xnor U21440 (N_21440,N_14851,N_14853);
nor U21441 (N_21441,N_17553,N_16317);
and U21442 (N_21442,N_16435,N_14433);
nor U21443 (N_21443,N_15725,N_17544);
or U21444 (N_21444,N_17031,N_12112);
or U21445 (N_21445,N_12117,N_15581);
or U21446 (N_21446,N_15770,N_15778);
xnor U21447 (N_21447,N_17428,N_14758);
xnor U21448 (N_21448,N_13608,N_12717);
or U21449 (N_21449,N_13457,N_12751);
xor U21450 (N_21450,N_12374,N_16499);
nor U21451 (N_21451,N_14262,N_17380);
nor U21452 (N_21452,N_14174,N_16088);
nor U21453 (N_21453,N_15550,N_16463);
and U21454 (N_21454,N_13495,N_13136);
and U21455 (N_21455,N_15350,N_14698);
or U21456 (N_21456,N_13690,N_14740);
or U21457 (N_21457,N_17937,N_17319);
and U21458 (N_21458,N_17495,N_14415);
and U21459 (N_21459,N_12242,N_12745);
and U21460 (N_21460,N_14064,N_12061);
or U21461 (N_21461,N_14174,N_15675);
nand U21462 (N_21462,N_12997,N_13486);
or U21463 (N_21463,N_12623,N_17403);
and U21464 (N_21464,N_15877,N_15640);
and U21465 (N_21465,N_17622,N_14490);
and U21466 (N_21466,N_15963,N_17588);
and U21467 (N_21467,N_15078,N_16952);
or U21468 (N_21468,N_17836,N_13891);
or U21469 (N_21469,N_15166,N_15041);
or U21470 (N_21470,N_17448,N_16347);
or U21471 (N_21471,N_14512,N_12053);
nand U21472 (N_21472,N_15471,N_14225);
or U21473 (N_21473,N_16088,N_14400);
or U21474 (N_21474,N_13138,N_16529);
xor U21475 (N_21475,N_12453,N_17779);
and U21476 (N_21476,N_15181,N_17332);
nor U21477 (N_21477,N_13390,N_14600);
nand U21478 (N_21478,N_15162,N_12628);
and U21479 (N_21479,N_12509,N_12367);
nor U21480 (N_21480,N_13329,N_16694);
and U21481 (N_21481,N_13831,N_17867);
nand U21482 (N_21482,N_13947,N_12742);
or U21483 (N_21483,N_17751,N_12055);
nand U21484 (N_21484,N_17525,N_15415);
xor U21485 (N_21485,N_15980,N_12577);
nand U21486 (N_21486,N_13995,N_14149);
nand U21487 (N_21487,N_17233,N_16221);
or U21488 (N_21488,N_14478,N_15014);
and U21489 (N_21489,N_17817,N_13936);
xnor U21490 (N_21490,N_14056,N_16289);
and U21491 (N_21491,N_14105,N_12748);
nand U21492 (N_21492,N_17313,N_12135);
and U21493 (N_21493,N_15169,N_13947);
nor U21494 (N_21494,N_16541,N_13505);
or U21495 (N_21495,N_15059,N_13146);
xnor U21496 (N_21496,N_12310,N_14840);
xor U21497 (N_21497,N_12566,N_13235);
or U21498 (N_21498,N_13383,N_14562);
or U21499 (N_21499,N_17084,N_13195);
or U21500 (N_21500,N_16046,N_15679);
xor U21501 (N_21501,N_16727,N_16886);
xor U21502 (N_21502,N_12048,N_14024);
nand U21503 (N_21503,N_17574,N_16495);
nor U21504 (N_21504,N_12566,N_12291);
xnor U21505 (N_21505,N_17199,N_15249);
nor U21506 (N_21506,N_15273,N_13531);
and U21507 (N_21507,N_12997,N_16992);
nor U21508 (N_21508,N_13017,N_12802);
or U21509 (N_21509,N_14486,N_16743);
nand U21510 (N_21510,N_15733,N_16730);
nor U21511 (N_21511,N_17042,N_15320);
nand U21512 (N_21512,N_13341,N_12634);
and U21513 (N_21513,N_15944,N_14946);
or U21514 (N_21514,N_12091,N_16512);
and U21515 (N_21515,N_14490,N_17296);
nand U21516 (N_21516,N_16831,N_12671);
and U21517 (N_21517,N_15596,N_17030);
or U21518 (N_21518,N_12012,N_14173);
nor U21519 (N_21519,N_16192,N_16915);
nand U21520 (N_21520,N_15061,N_16790);
and U21521 (N_21521,N_16590,N_14211);
nand U21522 (N_21522,N_14017,N_15019);
and U21523 (N_21523,N_12324,N_13516);
or U21524 (N_21524,N_17914,N_15243);
nor U21525 (N_21525,N_14902,N_13902);
or U21526 (N_21526,N_16241,N_13121);
nor U21527 (N_21527,N_16770,N_12622);
or U21528 (N_21528,N_15265,N_17983);
nand U21529 (N_21529,N_12900,N_12620);
or U21530 (N_21530,N_15756,N_12075);
nand U21531 (N_21531,N_13518,N_12183);
or U21532 (N_21532,N_14337,N_12183);
nand U21533 (N_21533,N_15229,N_15693);
or U21534 (N_21534,N_17437,N_15194);
or U21535 (N_21535,N_13978,N_13179);
and U21536 (N_21536,N_15041,N_13912);
nand U21537 (N_21537,N_14223,N_15103);
and U21538 (N_21538,N_13376,N_15213);
xor U21539 (N_21539,N_12025,N_16417);
nand U21540 (N_21540,N_17666,N_12561);
xor U21541 (N_21541,N_15658,N_17827);
xor U21542 (N_21542,N_17722,N_13250);
and U21543 (N_21543,N_17368,N_17879);
or U21544 (N_21544,N_13244,N_17593);
nand U21545 (N_21545,N_15154,N_12561);
nand U21546 (N_21546,N_15763,N_17570);
nand U21547 (N_21547,N_17657,N_14063);
nor U21548 (N_21548,N_13899,N_16861);
nand U21549 (N_21549,N_13181,N_12331);
nand U21550 (N_21550,N_12641,N_13643);
nand U21551 (N_21551,N_14600,N_17196);
nand U21552 (N_21552,N_16733,N_12518);
nor U21553 (N_21553,N_16697,N_14960);
nor U21554 (N_21554,N_16471,N_15937);
or U21555 (N_21555,N_17631,N_16026);
nor U21556 (N_21556,N_12634,N_13488);
xor U21557 (N_21557,N_15697,N_16892);
xor U21558 (N_21558,N_16602,N_15508);
xor U21559 (N_21559,N_12586,N_16719);
or U21560 (N_21560,N_13237,N_15407);
nand U21561 (N_21561,N_16946,N_16865);
and U21562 (N_21562,N_12559,N_17046);
or U21563 (N_21563,N_12380,N_17491);
nand U21564 (N_21564,N_15140,N_14372);
nand U21565 (N_21565,N_15938,N_13435);
nor U21566 (N_21566,N_16399,N_16885);
and U21567 (N_21567,N_17865,N_15579);
nor U21568 (N_21568,N_15896,N_13301);
or U21569 (N_21569,N_16926,N_12442);
nand U21570 (N_21570,N_16086,N_15119);
nand U21571 (N_21571,N_16172,N_17170);
xor U21572 (N_21572,N_13457,N_14179);
xor U21573 (N_21573,N_12073,N_12160);
and U21574 (N_21574,N_14108,N_12120);
nand U21575 (N_21575,N_16335,N_12484);
xnor U21576 (N_21576,N_12158,N_17088);
and U21577 (N_21577,N_13648,N_13181);
nor U21578 (N_21578,N_16417,N_14545);
nor U21579 (N_21579,N_14904,N_12840);
nor U21580 (N_21580,N_17618,N_16067);
nand U21581 (N_21581,N_16902,N_13677);
or U21582 (N_21582,N_12956,N_15925);
nand U21583 (N_21583,N_15316,N_15613);
nor U21584 (N_21584,N_12726,N_14946);
nand U21585 (N_21585,N_17975,N_12994);
nand U21586 (N_21586,N_17846,N_12996);
or U21587 (N_21587,N_14276,N_14030);
nand U21588 (N_21588,N_16910,N_17470);
nand U21589 (N_21589,N_12565,N_17637);
nor U21590 (N_21590,N_14434,N_15025);
nand U21591 (N_21591,N_17831,N_17742);
nand U21592 (N_21592,N_12663,N_17411);
and U21593 (N_21593,N_17394,N_16946);
or U21594 (N_21594,N_17598,N_16685);
or U21595 (N_21595,N_12384,N_17024);
nand U21596 (N_21596,N_16667,N_14005);
nor U21597 (N_21597,N_13768,N_12137);
nor U21598 (N_21598,N_12730,N_16356);
or U21599 (N_21599,N_17791,N_12223);
nand U21600 (N_21600,N_17977,N_16424);
or U21601 (N_21601,N_17032,N_15245);
nand U21602 (N_21602,N_13636,N_16708);
xnor U21603 (N_21603,N_12295,N_13065);
and U21604 (N_21604,N_13942,N_13948);
and U21605 (N_21605,N_14054,N_17719);
xnor U21606 (N_21606,N_12771,N_17478);
or U21607 (N_21607,N_13881,N_13666);
nor U21608 (N_21608,N_17005,N_14835);
nand U21609 (N_21609,N_12733,N_14123);
xor U21610 (N_21610,N_13998,N_13992);
xor U21611 (N_21611,N_15910,N_13824);
xor U21612 (N_21612,N_15531,N_14659);
nand U21613 (N_21613,N_17925,N_16775);
nand U21614 (N_21614,N_13523,N_16039);
nand U21615 (N_21615,N_17110,N_13845);
nand U21616 (N_21616,N_16475,N_12352);
nand U21617 (N_21617,N_13023,N_17755);
and U21618 (N_21618,N_13190,N_13411);
or U21619 (N_21619,N_16452,N_13875);
or U21620 (N_21620,N_15542,N_16249);
nor U21621 (N_21621,N_14601,N_14312);
nor U21622 (N_21622,N_12224,N_15457);
nor U21623 (N_21623,N_17019,N_16031);
xor U21624 (N_21624,N_12907,N_13902);
or U21625 (N_21625,N_12537,N_15508);
nor U21626 (N_21626,N_16389,N_12446);
nand U21627 (N_21627,N_12090,N_16304);
nor U21628 (N_21628,N_15668,N_14723);
or U21629 (N_21629,N_14729,N_12556);
and U21630 (N_21630,N_15077,N_13619);
and U21631 (N_21631,N_12280,N_17493);
or U21632 (N_21632,N_15669,N_12561);
nor U21633 (N_21633,N_15912,N_15222);
nor U21634 (N_21634,N_14317,N_16523);
or U21635 (N_21635,N_14418,N_14172);
xor U21636 (N_21636,N_13452,N_12661);
and U21637 (N_21637,N_12147,N_16625);
or U21638 (N_21638,N_16529,N_15133);
xor U21639 (N_21639,N_14980,N_14837);
xnor U21640 (N_21640,N_16392,N_17796);
or U21641 (N_21641,N_16415,N_16347);
or U21642 (N_21642,N_16424,N_17834);
and U21643 (N_21643,N_13568,N_13153);
nor U21644 (N_21644,N_17363,N_13695);
nand U21645 (N_21645,N_14316,N_15569);
or U21646 (N_21646,N_17769,N_15684);
nor U21647 (N_21647,N_14949,N_12303);
or U21648 (N_21648,N_13709,N_13766);
nor U21649 (N_21649,N_12202,N_16010);
xor U21650 (N_21650,N_14810,N_15748);
nor U21651 (N_21651,N_14472,N_14235);
xor U21652 (N_21652,N_17951,N_16439);
or U21653 (N_21653,N_16371,N_12292);
nor U21654 (N_21654,N_16255,N_12866);
nor U21655 (N_21655,N_16248,N_16556);
and U21656 (N_21656,N_12360,N_13198);
nor U21657 (N_21657,N_17347,N_17336);
nor U21658 (N_21658,N_12387,N_17801);
xor U21659 (N_21659,N_12247,N_15417);
nand U21660 (N_21660,N_13676,N_15403);
nand U21661 (N_21661,N_17058,N_12160);
and U21662 (N_21662,N_17728,N_12295);
nand U21663 (N_21663,N_17400,N_16921);
or U21664 (N_21664,N_15615,N_15877);
or U21665 (N_21665,N_16870,N_15808);
or U21666 (N_21666,N_14215,N_12220);
and U21667 (N_21667,N_12350,N_15312);
and U21668 (N_21668,N_13247,N_16272);
nor U21669 (N_21669,N_14695,N_17488);
xor U21670 (N_21670,N_12515,N_15821);
or U21671 (N_21671,N_16131,N_12694);
nand U21672 (N_21672,N_12225,N_17954);
and U21673 (N_21673,N_15796,N_16084);
or U21674 (N_21674,N_17254,N_14327);
and U21675 (N_21675,N_16603,N_13276);
or U21676 (N_21676,N_13012,N_16290);
nand U21677 (N_21677,N_16842,N_15541);
nor U21678 (N_21678,N_14773,N_14072);
or U21679 (N_21679,N_14080,N_13827);
nand U21680 (N_21680,N_12036,N_15055);
and U21681 (N_21681,N_14607,N_14788);
nor U21682 (N_21682,N_16859,N_15165);
nor U21683 (N_21683,N_17332,N_12738);
nand U21684 (N_21684,N_14548,N_17146);
or U21685 (N_21685,N_12512,N_17536);
nand U21686 (N_21686,N_12820,N_13934);
or U21687 (N_21687,N_13761,N_15014);
nor U21688 (N_21688,N_16647,N_14272);
nor U21689 (N_21689,N_14487,N_15816);
and U21690 (N_21690,N_12632,N_12222);
nand U21691 (N_21691,N_12385,N_13946);
or U21692 (N_21692,N_12791,N_15649);
nor U21693 (N_21693,N_16708,N_17824);
or U21694 (N_21694,N_15764,N_12608);
or U21695 (N_21695,N_13123,N_13673);
nand U21696 (N_21696,N_15629,N_15597);
or U21697 (N_21697,N_17605,N_14392);
or U21698 (N_21698,N_12272,N_12727);
nand U21699 (N_21699,N_13611,N_15469);
or U21700 (N_21700,N_14813,N_13136);
and U21701 (N_21701,N_17587,N_15202);
and U21702 (N_21702,N_16904,N_13093);
xor U21703 (N_21703,N_13734,N_12486);
or U21704 (N_21704,N_16858,N_12394);
or U21705 (N_21705,N_16347,N_12925);
nor U21706 (N_21706,N_12983,N_12677);
and U21707 (N_21707,N_17699,N_13934);
and U21708 (N_21708,N_14133,N_15487);
or U21709 (N_21709,N_14177,N_13006);
nor U21710 (N_21710,N_17699,N_15630);
and U21711 (N_21711,N_12694,N_13178);
nand U21712 (N_21712,N_17580,N_16740);
or U21713 (N_21713,N_15377,N_15944);
nor U21714 (N_21714,N_16512,N_14370);
or U21715 (N_21715,N_13764,N_14386);
and U21716 (N_21716,N_12898,N_16174);
nand U21717 (N_21717,N_12628,N_13323);
nor U21718 (N_21718,N_14113,N_16959);
and U21719 (N_21719,N_16551,N_17462);
nor U21720 (N_21720,N_16546,N_14404);
or U21721 (N_21721,N_14391,N_14477);
xor U21722 (N_21722,N_16654,N_14154);
nor U21723 (N_21723,N_17102,N_15304);
nand U21724 (N_21724,N_16455,N_14801);
nor U21725 (N_21725,N_17302,N_17024);
xor U21726 (N_21726,N_14662,N_17600);
or U21727 (N_21727,N_17142,N_17845);
xor U21728 (N_21728,N_12854,N_14982);
or U21729 (N_21729,N_16059,N_15192);
nand U21730 (N_21730,N_16493,N_17645);
nor U21731 (N_21731,N_15027,N_17742);
or U21732 (N_21732,N_12666,N_12453);
nand U21733 (N_21733,N_12613,N_15317);
nand U21734 (N_21734,N_12124,N_15566);
nand U21735 (N_21735,N_12410,N_16181);
xnor U21736 (N_21736,N_15989,N_14219);
nand U21737 (N_21737,N_13819,N_15935);
xor U21738 (N_21738,N_14910,N_16976);
nor U21739 (N_21739,N_14080,N_14231);
nand U21740 (N_21740,N_15111,N_12205);
and U21741 (N_21741,N_16297,N_16073);
nor U21742 (N_21742,N_17829,N_14830);
nor U21743 (N_21743,N_14594,N_16400);
nand U21744 (N_21744,N_12846,N_16028);
and U21745 (N_21745,N_17841,N_13952);
nor U21746 (N_21746,N_17514,N_17070);
nand U21747 (N_21747,N_13137,N_16271);
nor U21748 (N_21748,N_14421,N_14458);
xor U21749 (N_21749,N_16711,N_14793);
and U21750 (N_21750,N_15153,N_14227);
nand U21751 (N_21751,N_16786,N_12460);
or U21752 (N_21752,N_16977,N_17073);
nand U21753 (N_21753,N_16314,N_14890);
nor U21754 (N_21754,N_16350,N_13052);
and U21755 (N_21755,N_15296,N_12496);
nor U21756 (N_21756,N_14660,N_17866);
xnor U21757 (N_21757,N_16200,N_14727);
or U21758 (N_21758,N_13002,N_14119);
nor U21759 (N_21759,N_14222,N_17469);
and U21760 (N_21760,N_13166,N_12921);
and U21761 (N_21761,N_12414,N_13498);
nand U21762 (N_21762,N_12680,N_14691);
nand U21763 (N_21763,N_13127,N_14817);
xor U21764 (N_21764,N_16766,N_15910);
and U21765 (N_21765,N_15242,N_13294);
or U21766 (N_21766,N_12955,N_12593);
xor U21767 (N_21767,N_12959,N_12128);
and U21768 (N_21768,N_17120,N_15479);
nand U21769 (N_21769,N_16098,N_13801);
and U21770 (N_21770,N_16797,N_12062);
nand U21771 (N_21771,N_13204,N_17453);
nor U21772 (N_21772,N_14067,N_17576);
or U21773 (N_21773,N_15206,N_14517);
and U21774 (N_21774,N_14161,N_16811);
xnor U21775 (N_21775,N_16635,N_12955);
nand U21776 (N_21776,N_14087,N_14713);
nor U21777 (N_21777,N_13734,N_13969);
nand U21778 (N_21778,N_15643,N_16408);
or U21779 (N_21779,N_16301,N_12661);
and U21780 (N_21780,N_14413,N_16668);
nor U21781 (N_21781,N_17199,N_12929);
nor U21782 (N_21782,N_14157,N_17627);
nand U21783 (N_21783,N_12820,N_13044);
nand U21784 (N_21784,N_13622,N_16290);
and U21785 (N_21785,N_13461,N_17508);
or U21786 (N_21786,N_12239,N_14644);
xnor U21787 (N_21787,N_16406,N_16403);
and U21788 (N_21788,N_14289,N_16206);
nor U21789 (N_21789,N_15952,N_17099);
nand U21790 (N_21790,N_13344,N_12687);
or U21791 (N_21791,N_13044,N_14864);
xnor U21792 (N_21792,N_15819,N_17963);
nand U21793 (N_21793,N_14623,N_13581);
nand U21794 (N_21794,N_12122,N_15942);
nor U21795 (N_21795,N_16711,N_15465);
and U21796 (N_21796,N_14995,N_14769);
or U21797 (N_21797,N_14441,N_13304);
nor U21798 (N_21798,N_12446,N_13308);
or U21799 (N_21799,N_12461,N_13313);
xnor U21800 (N_21800,N_17490,N_16204);
nand U21801 (N_21801,N_17181,N_17033);
or U21802 (N_21802,N_13103,N_13573);
and U21803 (N_21803,N_14633,N_15927);
or U21804 (N_21804,N_16132,N_12724);
and U21805 (N_21805,N_15611,N_12571);
or U21806 (N_21806,N_16205,N_16634);
nor U21807 (N_21807,N_15222,N_14757);
nand U21808 (N_21808,N_16599,N_13319);
and U21809 (N_21809,N_12468,N_12264);
xor U21810 (N_21810,N_15198,N_16630);
and U21811 (N_21811,N_14984,N_13215);
nand U21812 (N_21812,N_15456,N_12916);
nand U21813 (N_21813,N_15992,N_12187);
and U21814 (N_21814,N_14948,N_13460);
nand U21815 (N_21815,N_16733,N_13600);
or U21816 (N_21816,N_13616,N_12798);
nand U21817 (N_21817,N_13677,N_12048);
nand U21818 (N_21818,N_14133,N_12528);
nand U21819 (N_21819,N_15834,N_15296);
nor U21820 (N_21820,N_12512,N_13546);
nand U21821 (N_21821,N_13845,N_13238);
and U21822 (N_21822,N_15715,N_12863);
or U21823 (N_21823,N_14477,N_12536);
nor U21824 (N_21824,N_14857,N_17696);
xnor U21825 (N_21825,N_15857,N_17690);
xnor U21826 (N_21826,N_14811,N_14559);
nor U21827 (N_21827,N_12425,N_16762);
xnor U21828 (N_21828,N_16131,N_14800);
and U21829 (N_21829,N_17562,N_16212);
or U21830 (N_21830,N_13932,N_16944);
nor U21831 (N_21831,N_14361,N_17534);
nor U21832 (N_21832,N_12220,N_13828);
xnor U21833 (N_21833,N_12068,N_16322);
nor U21834 (N_21834,N_14620,N_14683);
nand U21835 (N_21835,N_15761,N_14695);
and U21836 (N_21836,N_12388,N_13783);
and U21837 (N_21837,N_12132,N_12627);
and U21838 (N_21838,N_14851,N_17340);
nand U21839 (N_21839,N_15738,N_16801);
or U21840 (N_21840,N_14485,N_17817);
nand U21841 (N_21841,N_17354,N_13079);
nand U21842 (N_21842,N_16874,N_15805);
nand U21843 (N_21843,N_12768,N_12627);
nor U21844 (N_21844,N_13378,N_17749);
nand U21845 (N_21845,N_12938,N_16820);
or U21846 (N_21846,N_14837,N_12721);
nand U21847 (N_21847,N_13678,N_12362);
nand U21848 (N_21848,N_17235,N_13448);
or U21849 (N_21849,N_14937,N_15229);
and U21850 (N_21850,N_16323,N_15083);
and U21851 (N_21851,N_16409,N_16480);
nand U21852 (N_21852,N_14505,N_17206);
nor U21853 (N_21853,N_13472,N_16092);
or U21854 (N_21854,N_15731,N_15573);
and U21855 (N_21855,N_16329,N_13150);
nor U21856 (N_21856,N_13340,N_15737);
nand U21857 (N_21857,N_13812,N_14018);
nand U21858 (N_21858,N_16995,N_15110);
nor U21859 (N_21859,N_13110,N_13735);
or U21860 (N_21860,N_13556,N_14635);
nand U21861 (N_21861,N_15860,N_14465);
nand U21862 (N_21862,N_17720,N_12777);
and U21863 (N_21863,N_12947,N_12345);
nand U21864 (N_21864,N_14802,N_13479);
nor U21865 (N_21865,N_17683,N_17107);
nand U21866 (N_21866,N_16764,N_14842);
nor U21867 (N_21867,N_13531,N_12369);
nor U21868 (N_21868,N_15368,N_14098);
nor U21869 (N_21869,N_13418,N_15826);
or U21870 (N_21870,N_17158,N_14679);
nor U21871 (N_21871,N_13995,N_16347);
nand U21872 (N_21872,N_15315,N_16490);
nor U21873 (N_21873,N_12282,N_16271);
or U21874 (N_21874,N_14066,N_15183);
and U21875 (N_21875,N_13685,N_17072);
xnor U21876 (N_21876,N_16059,N_12809);
or U21877 (N_21877,N_14029,N_13842);
and U21878 (N_21878,N_14632,N_15819);
and U21879 (N_21879,N_13549,N_13218);
and U21880 (N_21880,N_15917,N_17090);
nor U21881 (N_21881,N_13488,N_15837);
or U21882 (N_21882,N_12367,N_17550);
and U21883 (N_21883,N_14442,N_12483);
and U21884 (N_21884,N_15333,N_12122);
or U21885 (N_21885,N_16295,N_12782);
or U21886 (N_21886,N_16452,N_15428);
and U21887 (N_21887,N_15226,N_12847);
and U21888 (N_21888,N_14526,N_14004);
nor U21889 (N_21889,N_12144,N_15856);
or U21890 (N_21890,N_12703,N_14803);
nand U21891 (N_21891,N_13759,N_14386);
or U21892 (N_21892,N_14845,N_15850);
and U21893 (N_21893,N_14291,N_15108);
and U21894 (N_21894,N_14055,N_15611);
nand U21895 (N_21895,N_16626,N_15159);
nand U21896 (N_21896,N_16233,N_14025);
nor U21897 (N_21897,N_15035,N_13338);
nand U21898 (N_21898,N_14267,N_16755);
and U21899 (N_21899,N_17602,N_12540);
or U21900 (N_21900,N_14347,N_13332);
nand U21901 (N_21901,N_15205,N_16524);
nor U21902 (N_21902,N_13466,N_15543);
nor U21903 (N_21903,N_17921,N_16731);
nand U21904 (N_21904,N_17645,N_17610);
nand U21905 (N_21905,N_17355,N_16048);
and U21906 (N_21906,N_14458,N_15834);
and U21907 (N_21907,N_16918,N_12489);
and U21908 (N_21908,N_14265,N_14849);
or U21909 (N_21909,N_13159,N_15935);
nor U21910 (N_21910,N_16090,N_13971);
or U21911 (N_21911,N_17182,N_15364);
or U21912 (N_21912,N_14934,N_14383);
or U21913 (N_21913,N_14770,N_14856);
and U21914 (N_21914,N_13220,N_16649);
nor U21915 (N_21915,N_17440,N_15333);
nor U21916 (N_21916,N_14083,N_16139);
nor U21917 (N_21917,N_13350,N_12454);
or U21918 (N_21918,N_15705,N_13076);
nor U21919 (N_21919,N_16520,N_13110);
nand U21920 (N_21920,N_14958,N_12244);
nor U21921 (N_21921,N_16902,N_17566);
xor U21922 (N_21922,N_14555,N_16585);
xor U21923 (N_21923,N_12571,N_16458);
and U21924 (N_21924,N_13943,N_14644);
and U21925 (N_21925,N_16654,N_13528);
and U21926 (N_21926,N_17640,N_14571);
xnor U21927 (N_21927,N_14883,N_12557);
nor U21928 (N_21928,N_14507,N_14918);
nor U21929 (N_21929,N_12424,N_17990);
nand U21930 (N_21930,N_15884,N_15397);
nand U21931 (N_21931,N_17421,N_17218);
nand U21932 (N_21932,N_12954,N_12161);
xor U21933 (N_21933,N_17676,N_17141);
xor U21934 (N_21934,N_15264,N_12573);
or U21935 (N_21935,N_17763,N_14240);
or U21936 (N_21936,N_13064,N_15585);
nor U21937 (N_21937,N_12830,N_17937);
and U21938 (N_21938,N_17205,N_15574);
or U21939 (N_21939,N_15055,N_15537);
or U21940 (N_21940,N_17490,N_14336);
or U21941 (N_21941,N_17355,N_12004);
or U21942 (N_21942,N_16265,N_13630);
and U21943 (N_21943,N_16783,N_16436);
and U21944 (N_21944,N_14400,N_17213);
nand U21945 (N_21945,N_12438,N_14789);
and U21946 (N_21946,N_13964,N_17511);
or U21947 (N_21947,N_16648,N_16664);
nand U21948 (N_21948,N_12102,N_15548);
or U21949 (N_21949,N_16210,N_13270);
and U21950 (N_21950,N_13577,N_17448);
or U21951 (N_21951,N_16175,N_16406);
xor U21952 (N_21952,N_15468,N_13100);
nor U21953 (N_21953,N_17433,N_12373);
nand U21954 (N_21954,N_15418,N_12394);
nor U21955 (N_21955,N_12531,N_16800);
xor U21956 (N_21956,N_15151,N_16120);
nor U21957 (N_21957,N_16741,N_14006);
nand U21958 (N_21958,N_12500,N_14496);
or U21959 (N_21959,N_16294,N_17141);
nand U21960 (N_21960,N_16454,N_16329);
and U21961 (N_21961,N_12912,N_17293);
nor U21962 (N_21962,N_12934,N_13460);
nand U21963 (N_21963,N_12976,N_15411);
or U21964 (N_21964,N_13362,N_15957);
nand U21965 (N_21965,N_17442,N_14053);
nand U21966 (N_21966,N_14615,N_14309);
nor U21967 (N_21967,N_16601,N_14053);
nand U21968 (N_21968,N_14518,N_12141);
nand U21969 (N_21969,N_12615,N_14625);
or U21970 (N_21970,N_15782,N_16257);
nor U21971 (N_21971,N_17924,N_13681);
or U21972 (N_21972,N_15686,N_14720);
or U21973 (N_21973,N_15752,N_12531);
nand U21974 (N_21974,N_16733,N_15314);
or U21975 (N_21975,N_13291,N_15792);
and U21976 (N_21976,N_15907,N_17629);
nand U21977 (N_21977,N_17082,N_16153);
and U21978 (N_21978,N_14526,N_15446);
or U21979 (N_21979,N_15893,N_14320);
or U21980 (N_21980,N_16429,N_16954);
or U21981 (N_21981,N_13372,N_15146);
or U21982 (N_21982,N_14057,N_14016);
or U21983 (N_21983,N_14787,N_12444);
and U21984 (N_21984,N_13139,N_12961);
nand U21985 (N_21985,N_15921,N_15419);
nor U21986 (N_21986,N_13031,N_17485);
or U21987 (N_21987,N_13284,N_13042);
nand U21988 (N_21988,N_12566,N_13278);
or U21989 (N_21989,N_15204,N_17557);
nand U21990 (N_21990,N_13493,N_12133);
or U21991 (N_21991,N_15423,N_16094);
or U21992 (N_21992,N_13012,N_15531);
xor U21993 (N_21993,N_12709,N_12499);
or U21994 (N_21994,N_12323,N_15070);
and U21995 (N_21995,N_14631,N_15782);
nand U21996 (N_21996,N_15984,N_16141);
and U21997 (N_21997,N_12934,N_16910);
or U21998 (N_21998,N_15585,N_15000);
or U21999 (N_21999,N_14115,N_15288);
and U22000 (N_22000,N_13708,N_14982);
nor U22001 (N_22001,N_15655,N_12018);
nand U22002 (N_22002,N_16932,N_13440);
or U22003 (N_22003,N_12869,N_17497);
or U22004 (N_22004,N_17844,N_14754);
nand U22005 (N_22005,N_14704,N_14218);
nor U22006 (N_22006,N_16618,N_15187);
or U22007 (N_22007,N_17536,N_12402);
nand U22008 (N_22008,N_16608,N_14396);
and U22009 (N_22009,N_13655,N_16633);
nor U22010 (N_22010,N_14536,N_14421);
or U22011 (N_22011,N_12576,N_14126);
nor U22012 (N_22012,N_12045,N_12844);
nor U22013 (N_22013,N_14472,N_14049);
xor U22014 (N_22014,N_13809,N_15429);
nor U22015 (N_22015,N_13551,N_13222);
nand U22016 (N_22016,N_17767,N_14138);
and U22017 (N_22017,N_12410,N_15697);
xnor U22018 (N_22018,N_15969,N_17889);
or U22019 (N_22019,N_15078,N_16932);
nor U22020 (N_22020,N_13809,N_16456);
and U22021 (N_22021,N_14247,N_15137);
or U22022 (N_22022,N_13398,N_13568);
or U22023 (N_22023,N_16417,N_16027);
and U22024 (N_22024,N_16794,N_15756);
xnor U22025 (N_22025,N_14229,N_16601);
and U22026 (N_22026,N_16930,N_16846);
and U22027 (N_22027,N_16780,N_12136);
or U22028 (N_22028,N_16595,N_13796);
and U22029 (N_22029,N_17773,N_12596);
nor U22030 (N_22030,N_14845,N_16649);
nor U22031 (N_22031,N_14599,N_13663);
xnor U22032 (N_22032,N_12081,N_17060);
nand U22033 (N_22033,N_12339,N_15743);
and U22034 (N_22034,N_16578,N_12731);
or U22035 (N_22035,N_16784,N_17510);
nand U22036 (N_22036,N_14876,N_16049);
nor U22037 (N_22037,N_14669,N_13294);
nand U22038 (N_22038,N_12899,N_13354);
nor U22039 (N_22039,N_16557,N_13334);
and U22040 (N_22040,N_14108,N_13782);
nor U22041 (N_22041,N_14155,N_12518);
nor U22042 (N_22042,N_15214,N_12063);
nand U22043 (N_22043,N_12331,N_17037);
and U22044 (N_22044,N_15660,N_13966);
nand U22045 (N_22045,N_14838,N_13529);
and U22046 (N_22046,N_15795,N_16219);
nand U22047 (N_22047,N_17158,N_13629);
and U22048 (N_22048,N_16645,N_12402);
nor U22049 (N_22049,N_12505,N_16767);
or U22050 (N_22050,N_12162,N_17471);
or U22051 (N_22051,N_12104,N_15118);
nand U22052 (N_22052,N_13414,N_17105);
and U22053 (N_22053,N_12133,N_17535);
or U22054 (N_22054,N_14368,N_15693);
nand U22055 (N_22055,N_14555,N_14413);
nand U22056 (N_22056,N_13820,N_13503);
or U22057 (N_22057,N_12388,N_17286);
nand U22058 (N_22058,N_14398,N_12732);
nor U22059 (N_22059,N_16750,N_12069);
nor U22060 (N_22060,N_14653,N_15374);
and U22061 (N_22061,N_14834,N_12126);
or U22062 (N_22062,N_17857,N_17484);
and U22063 (N_22063,N_15916,N_15508);
and U22064 (N_22064,N_13586,N_13837);
xnor U22065 (N_22065,N_14141,N_12960);
and U22066 (N_22066,N_17260,N_17204);
or U22067 (N_22067,N_13296,N_17711);
or U22068 (N_22068,N_13074,N_14930);
nor U22069 (N_22069,N_13757,N_14104);
nor U22070 (N_22070,N_15491,N_15967);
nor U22071 (N_22071,N_16003,N_14292);
or U22072 (N_22072,N_17643,N_16882);
nor U22073 (N_22073,N_12843,N_13115);
nor U22074 (N_22074,N_15982,N_12974);
or U22075 (N_22075,N_12301,N_17953);
and U22076 (N_22076,N_13163,N_16390);
and U22077 (N_22077,N_15114,N_12197);
nor U22078 (N_22078,N_15940,N_17179);
or U22079 (N_22079,N_16818,N_15016);
or U22080 (N_22080,N_13381,N_13627);
and U22081 (N_22081,N_12208,N_16891);
nor U22082 (N_22082,N_17677,N_13113);
nand U22083 (N_22083,N_12400,N_15392);
nand U22084 (N_22084,N_13970,N_15889);
and U22085 (N_22085,N_16196,N_12299);
and U22086 (N_22086,N_12797,N_14053);
nand U22087 (N_22087,N_12165,N_13618);
nor U22088 (N_22088,N_17328,N_15089);
nand U22089 (N_22089,N_13988,N_16239);
or U22090 (N_22090,N_12775,N_14061);
nand U22091 (N_22091,N_15079,N_15279);
xnor U22092 (N_22092,N_17683,N_17045);
nor U22093 (N_22093,N_17278,N_15214);
or U22094 (N_22094,N_13563,N_17129);
nand U22095 (N_22095,N_12973,N_12744);
nor U22096 (N_22096,N_12186,N_12102);
nand U22097 (N_22097,N_12634,N_12804);
nand U22098 (N_22098,N_13983,N_17131);
nor U22099 (N_22099,N_13502,N_12439);
and U22100 (N_22100,N_16126,N_12250);
nor U22101 (N_22101,N_17999,N_15062);
xnor U22102 (N_22102,N_14137,N_15261);
nand U22103 (N_22103,N_17013,N_17570);
and U22104 (N_22104,N_14758,N_15311);
and U22105 (N_22105,N_13935,N_13865);
or U22106 (N_22106,N_12007,N_14843);
nor U22107 (N_22107,N_14610,N_13874);
or U22108 (N_22108,N_17638,N_12870);
nand U22109 (N_22109,N_13610,N_17788);
nor U22110 (N_22110,N_17623,N_17542);
xnor U22111 (N_22111,N_17525,N_16984);
and U22112 (N_22112,N_13120,N_12222);
or U22113 (N_22113,N_15475,N_15584);
nand U22114 (N_22114,N_17908,N_12076);
nor U22115 (N_22115,N_15551,N_17412);
and U22116 (N_22116,N_14867,N_16562);
or U22117 (N_22117,N_17245,N_15306);
nor U22118 (N_22118,N_15583,N_12269);
and U22119 (N_22119,N_14635,N_14754);
and U22120 (N_22120,N_16200,N_12159);
nand U22121 (N_22121,N_17986,N_12933);
or U22122 (N_22122,N_14610,N_16186);
or U22123 (N_22123,N_16502,N_17959);
xnor U22124 (N_22124,N_17818,N_16747);
and U22125 (N_22125,N_17697,N_12469);
or U22126 (N_22126,N_12248,N_12808);
and U22127 (N_22127,N_15894,N_14504);
nor U22128 (N_22128,N_15511,N_17404);
and U22129 (N_22129,N_12584,N_16381);
or U22130 (N_22130,N_13792,N_16993);
nand U22131 (N_22131,N_17956,N_14054);
nor U22132 (N_22132,N_17184,N_16891);
nor U22133 (N_22133,N_15708,N_13044);
nor U22134 (N_22134,N_17444,N_13027);
and U22135 (N_22135,N_12443,N_16382);
nand U22136 (N_22136,N_16005,N_16061);
or U22137 (N_22137,N_15465,N_15342);
and U22138 (N_22138,N_13289,N_14550);
or U22139 (N_22139,N_17472,N_16712);
and U22140 (N_22140,N_12663,N_16065);
and U22141 (N_22141,N_17133,N_13332);
nand U22142 (N_22142,N_13186,N_17245);
or U22143 (N_22143,N_16914,N_14563);
nand U22144 (N_22144,N_14803,N_14988);
nor U22145 (N_22145,N_16221,N_13921);
nor U22146 (N_22146,N_16869,N_17761);
or U22147 (N_22147,N_13553,N_17777);
or U22148 (N_22148,N_16415,N_17487);
and U22149 (N_22149,N_17006,N_14215);
or U22150 (N_22150,N_12582,N_12601);
or U22151 (N_22151,N_16536,N_12913);
or U22152 (N_22152,N_12996,N_16356);
xnor U22153 (N_22153,N_17118,N_16947);
nand U22154 (N_22154,N_17692,N_15856);
and U22155 (N_22155,N_13770,N_17011);
nor U22156 (N_22156,N_13801,N_12901);
nand U22157 (N_22157,N_12374,N_12123);
xnor U22158 (N_22158,N_15480,N_16780);
or U22159 (N_22159,N_13753,N_13726);
and U22160 (N_22160,N_12323,N_15826);
nor U22161 (N_22161,N_12232,N_15695);
and U22162 (N_22162,N_14003,N_12346);
nand U22163 (N_22163,N_17061,N_13162);
xor U22164 (N_22164,N_15951,N_16939);
nor U22165 (N_22165,N_13058,N_17206);
or U22166 (N_22166,N_13262,N_12819);
xnor U22167 (N_22167,N_12064,N_15142);
nor U22168 (N_22168,N_15213,N_14208);
nand U22169 (N_22169,N_13841,N_13940);
nor U22170 (N_22170,N_14461,N_17810);
nor U22171 (N_22171,N_15296,N_12163);
nand U22172 (N_22172,N_12455,N_12634);
or U22173 (N_22173,N_13602,N_16680);
nor U22174 (N_22174,N_17062,N_13562);
nand U22175 (N_22175,N_16036,N_13161);
nand U22176 (N_22176,N_12371,N_17890);
and U22177 (N_22177,N_17831,N_12476);
and U22178 (N_22178,N_15824,N_12508);
and U22179 (N_22179,N_14674,N_15374);
or U22180 (N_22180,N_12875,N_16402);
or U22181 (N_22181,N_13588,N_13717);
and U22182 (N_22182,N_12207,N_14531);
nor U22183 (N_22183,N_17911,N_15824);
nand U22184 (N_22184,N_14340,N_16296);
nand U22185 (N_22185,N_15842,N_13620);
nand U22186 (N_22186,N_15045,N_12096);
nor U22187 (N_22187,N_12603,N_17582);
nor U22188 (N_22188,N_15259,N_13289);
or U22189 (N_22189,N_15366,N_16912);
nor U22190 (N_22190,N_14149,N_14337);
xor U22191 (N_22191,N_13831,N_13196);
and U22192 (N_22192,N_17243,N_12334);
nor U22193 (N_22193,N_12627,N_13784);
or U22194 (N_22194,N_14386,N_14300);
and U22195 (N_22195,N_17253,N_16734);
nor U22196 (N_22196,N_12071,N_13651);
or U22197 (N_22197,N_13367,N_13147);
and U22198 (N_22198,N_13244,N_15882);
nor U22199 (N_22199,N_12475,N_13663);
nor U22200 (N_22200,N_14880,N_12190);
or U22201 (N_22201,N_13472,N_14745);
nor U22202 (N_22202,N_16886,N_17513);
nor U22203 (N_22203,N_13368,N_17031);
nand U22204 (N_22204,N_16328,N_15364);
nor U22205 (N_22205,N_15114,N_15083);
or U22206 (N_22206,N_17107,N_15320);
or U22207 (N_22207,N_17056,N_15649);
nor U22208 (N_22208,N_16516,N_14204);
nand U22209 (N_22209,N_16100,N_17381);
nor U22210 (N_22210,N_17110,N_16123);
and U22211 (N_22211,N_17156,N_12646);
nor U22212 (N_22212,N_16071,N_13721);
xnor U22213 (N_22213,N_17416,N_17221);
nand U22214 (N_22214,N_12953,N_12907);
nor U22215 (N_22215,N_14722,N_13108);
nor U22216 (N_22216,N_14214,N_14357);
xor U22217 (N_22217,N_14496,N_15365);
nand U22218 (N_22218,N_17703,N_15943);
nand U22219 (N_22219,N_16817,N_15762);
and U22220 (N_22220,N_13696,N_12621);
and U22221 (N_22221,N_15748,N_13115);
xor U22222 (N_22222,N_17155,N_16195);
nor U22223 (N_22223,N_17992,N_16481);
and U22224 (N_22224,N_12570,N_13790);
nor U22225 (N_22225,N_12977,N_16928);
xnor U22226 (N_22226,N_17696,N_12444);
and U22227 (N_22227,N_12933,N_15000);
nor U22228 (N_22228,N_12489,N_17609);
and U22229 (N_22229,N_12691,N_14329);
xnor U22230 (N_22230,N_17155,N_15518);
xor U22231 (N_22231,N_16087,N_17398);
nor U22232 (N_22232,N_15610,N_16038);
nand U22233 (N_22233,N_12140,N_16708);
xor U22234 (N_22234,N_13454,N_16802);
nand U22235 (N_22235,N_12840,N_12548);
and U22236 (N_22236,N_14317,N_12918);
and U22237 (N_22237,N_14794,N_12465);
or U22238 (N_22238,N_13374,N_15522);
or U22239 (N_22239,N_14364,N_12376);
nand U22240 (N_22240,N_14286,N_12152);
nor U22241 (N_22241,N_17819,N_12787);
and U22242 (N_22242,N_17730,N_14272);
xnor U22243 (N_22243,N_16845,N_17450);
nor U22244 (N_22244,N_13887,N_16651);
nand U22245 (N_22245,N_14080,N_14992);
nor U22246 (N_22246,N_15553,N_17902);
nand U22247 (N_22247,N_17517,N_17525);
or U22248 (N_22248,N_13989,N_17796);
or U22249 (N_22249,N_12591,N_16441);
and U22250 (N_22250,N_14061,N_16648);
xnor U22251 (N_22251,N_13095,N_15150);
nor U22252 (N_22252,N_14382,N_13425);
and U22253 (N_22253,N_15902,N_12900);
and U22254 (N_22254,N_17011,N_15673);
nand U22255 (N_22255,N_14876,N_17088);
nor U22256 (N_22256,N_16076,N_17587);
xnor U22257 (N_22257,N_17646,N_12174);
nor U22258 (N_22258,N_12225,N_14517);
or U22259 (N_22259,N_17508,N_17209);
xor U22260 (N_22260,N_15256,N_12233);
and U22261 (N_22261,N_16569,N_13777);
xnor U22262 (N_22262,N_12700,N_14584);
and U22263 (N_22263,N_16257,N_17078);
and U22264 (N_22264,N_15969,N_14435);
or U22265 (N_22265,N_12060,N_12524);
xnor U22266 (N_22266,N_12479,N_13552);
and U22267 (N_22267,N_13196,N_14480);
or U22268 (N_22268,N_12882,N_14693);
nor U22269 (N_22269,N_12128,N_14551);
xor U22270 (N_22270,N_15453,N_14567);
or U22271 (N_22271,N_13851,N_17820);
nor U22272 (N_22272,N_15479,N_15290);
nor U22273 (N_22273,N_13901,N_15344);
nor U22274 (N_22274,N_14619,N_15280);
nand U22275 (N_22275,N_13391,N_15315);
xnor U22276 (N_22276,N_12424,N_16086);
or U22277 (N_22277,N_12885,N_16968);
or U22278 (N_22278,N_16845,N_16121);
nor U22279 (N_22279,N_15566,N_17436);
nor U22280 (N_22280,N_16475,N_16347);
and U22281 (N_22281,N_16751,N_14379);
nor U22282 (N_22282,N_17380,N_17108);
and U22283 (N_22283,N_15161,N_14612);
nand U22284 (N_22284,N_12617,N_16299);
nor U22285 (N_22285,N_13785,N_12598);
or U22286 (N_22286,N_12016,N_16607);
and U22287 (N_22287,N_17617,N_17336);
and U22288 (N_22288,N_12985,N_15137);
nand U22289 (N_22289,N_13738,N_13598);
nor U22290 (N_22290,N_13789,N_17969);
nor U22291 (N_22291,N_17212,N_16820);
nor U22292 (N_22292,N_12102,N_15549);
nor U22293 (N_22293,N_12070,N_16821);
nor U22294 (N_22294,N_13263,N_13596);
and U22295 (N_22295,N_13199,N_14055);
or U22296 (N_22296,N_12938,N_16433);
xor U22297 (N_22297,N_17184,N_13974);
nand U22298 (N_22298,N_16988,N_15936);
nor U22299 (N_22299,N_16375,N_13004);
or U22300 (N_22300,N_12732,N_16875);
nand U22301 (N_22301,N_17478,N_13044);
nand U22302 (N_22302,N_12462,N_17998);
nand U22303 (N_22303,N_17284,N_14448);
nand U22304 (N_22304,N_14101,N_16961);
or U22305 (N_22305,N_14155,N_16108);
or U22306 (N_22306,N_12914,N_13323);
nor U22307 (N_22307,N_13331,N_12428);
or U22308 (N_22308,N_12280,N_13364);
or U22309 (N_22309,N_17908,N_15826);
nand U22310 (N_22310,N_16590,N_14484);
and U22311 (N_22311,N_15723,N_17851);
nor U22312 (N_22312,N_14526,N_13762);
xnor U22313 (N_22313,N_15713,N_12390);
xnor U22314 (N_22314,N_15044,N_14880);
or U22315 (N_22315,N_14331,N_13951);
nand U22316 (N_22316,N_13908,N_13752);
or U22317 (N_22317,N_12500,N_12926);
nand U22318 (N_22318,N_16049,N_16635);
nor U22319 (N_22319,N_15171,N_12464);
nor U22320 (N_22320,N_14357,N_14775);
xnor U22321 (N_22321,N_15928,N_15264);
or U22322 (N_22322,N_12912,N_14096);
xnor U22323 (N_22323,N_14748,N_15844);
nand U22324 (N_22324,N_14908,N_16655);
or U22325 (N_22325,N_16754,N_15576);
and U22326 (N_22326,N_16853,N_16655);
and U22327 (N_22327,N_13548,N_14071);
and U22328 (N_22328,N_13322,N_15294);
nand U22329 (N_22329,N_16447,N_12832);
nand U22330 (N_22330,N_12783,N_14653);
nand U22331 (N_22331,N_16959,N_16623);
or U22332 (N_22332,N_16660,N_15312);
nand U22333 (N_22333,N_13639,N_12157);
xnor U22334 (N_22334,N_14749,N_17829);
nand U22335 (N_22335,N_14742,N_16650);
or U22336 (N_22336,N_13102,N_15663);
nor U22337 (N_22337,N_16757,N_16457);
nand U22338 (N_22338,N_15857,N_12386);
and U22339 (N_22339,N_12917,N_15617);
xnor U22340 (N_22340,N_12398,N_15138);
nand U22341 (N_22341,N_15004,N_16142);
and U22342 (N_22342,N_16410,N_15346);
and U22343 (N_22343,N_17716,N_15844);
nand U22344 (N_22344,N_14092,N_12583);
nor U22345 (N_22345,N_17591,N_12731);
nor U22346 (N_22346,N_16978,N_13500);
nand U22347 (N_22347,N_14447,N_16955);
and U22348 (N_22348,N_12339,N_15456);
xor U22349 (N_22349,N_15308,N_14563);
or U22350 (N_22350,N_16261,N_14245);
or U22351 (N_22351,N_12152,N_14018);
xnor U22352 (N_22352,N_13263,N_16408);
and U22353 (N_22353,N_14956,N_17182);
nand U22354 (N_22354,N_13322,N_12418);
nand U22355 (N_22355,N_15057,N_12586);
nand U22356 (N_22356,N_15172,N_17040);
nor U22357 (N_22357,N_14799,N_15667);
or U22358 (N_22358,N_15890,N_13244);
nor U22359 (N_22359,N_12450,N_13819);
nor U22360 (N_22360,N_12980,N_15421);
nand U22361 (N_22361,N_13967,N_16725);
nand U22362 (N_22362,N_15931,N_15719);
and U22363 (N_22363,N_14981,N_12672);
xnor U22364 (N_22364,N_17847,N_16662);
or U22365 (N_22365,N_15101,N_15337);
xnor U22366 (N_22366,N_17540,N_16744);
and U22367 (N_22367,N_15702,N_13135);
xnor U22368 (N_22368,N_16398,N_15418);
or U22369 (N_22369,N_13181,N_16524);
nor U22370 (N_22370,N_14572,N_14737);
and U22371 (N_22371,N_15147,N_17894);
nor U22372 (N_22372,N_13471,N_12263);
or U22373 (N_22373,N_17728,N_16604);
nand U22374 (N_22374,N_15120,N_15872);
nand U22375 (N_22375,N_15338,N_13510);
nand U22376 (N_22376,N_16245,N_16767);
or U22377 (N_22377,N_16013,N_17722);
nand U22378 (N_22378,N_12049,N_12795);
xnor U22379 (N_22379,N_16869,N_12376);
nor U22380 (N_22380,N_12406,N_14624);
xnor U22381 (N_22381,N_15865,N_17310);
xor U22382 (N_22382,N_13068,N_13957);
nand U22383 (N_22383,N_14583,N_16782);
nor U22384 (N_22384,N_17798,N_14783);
or U22385 (N_22385,N_13331,N_16846);
nor U22386 (N_22386,N_16097,N_13848);
nand U22387 (N_22387,N_15135,N_17955);
and U22388 (N_22388,N_17597,N_14328);
nor U22389 (N_22389,N_12887,N_17913);
or U22390 (N_22390,N_16164,N_15601);
or U22391 (N_22391,N_13381,N_16566);
nor U22392 (N_22392,N_15626,N_17283);
nand U22393 (N_22393,N_17117,N_16986);
or U22394 (N_22394,N_13468,N_14801);
nor U22395 (N_22395,N_14853,N_13274);
or U22396 (N_22396,N_16818,N_12592);
or U22397 (N_22397,N_12914,N_13128);
and U22398 (N_22398,N_16796,N_12911);
and U22399 (N_22399,N_16773,N_15458);
and U22400 (N_22400,N_17955,N_16779);
or U22401 (N_22401,N_12673,N_15288);
and U22402 (N_22402,N_12253,N_16886);
nor U22403 (N_22403,N_16303,N_16776);
and U22404 (N_22404,N_16050,N_15264);
and U22405 (N_22405,N_14252,N_13771);
nor U22406 (N_22406,N_16731,N_12599);
nor U22407 (N_22407,N_16570,N_15841);
xnor U22408 (N_22408,N_17952,N_14365);
nand U22409 (N_22409,N_17523,N_17793);
nand U22410 (N_22410,N_16894,N_16356);
and U22411 (N_22411,N_14731,N_12014);
nand U22412 (N_22412,N_12134,N_15232);
nand U22413 (N_22413,N_15590,N_16757);
nor U22414 (N_22414,N_14733,N_12195);
nand U22415 (N_22415,N_16498,N_17145);
nor U22416 (N_22416,N_12731,N_14369);
and U22417 (N_22417,N_13001,N_13204);
or U22418 (N_22418,N_16760,N_13557);
xor U22419 (N_22419,N_14483,N_12995);
nand U22420 (N_22420,N_14050,N_15404);
nor U22421 (N_22421,N_17534,N_16006);
xor U22422 (N_22422,N_14303,N_17950);
nor U22423 (N_22423,N_16914,N_14017);
nor U22424 (N_22424,N_16602,N_14133);
nor U22425 (N_22425,N_12706,N_15643);
nand U22426 (N_22426,N_17245,N_13465);
nand U22427 (N_22427,N_12864,N_15121);
nor U22428 (N_22428,N_17770,N_14511);
and U22429 (N_22429,N_13222,N_14833);
nand U22430 (N_22430,N_17488,N_16166);
and U22431 (N_22431,N_15826,N_14603);
or U22432 (N_22432,N_13737,N_14477);
nor U22433 (N_22433,N_15935,N_12919);
and U22434 (N_22434,N_13572,N_12522);
nand U22435 (N_22435,N_12553,N_16495);
nor U22436 (N_22436,N_14920,N_13080);
xor U22437 (N_22437,N_17735,N_17351);
xor U22438 (N_22438,N_17601,N_12280);
and U22439 (N_22439,N_12786,N_16079);
and U22440 (N_22440,N_12976,N_15058);
and U22441 (N_22441,N_16749,N_15667);
or U22442 (N_22442,N_15101,N_14733);
and U22443 (N_22443,N_16769,N_14572);
nand U22444 (N_22444,N_12543,N_12551);
nor U22445 (N_22445,N_16804,N_12799);
or U22446 (N_22446,N_16991,N_16844);
and U22447 (N_22447,N_12501,N_13978);
nor U22448 (N_22448,N_13481,N_16520);
and U22449 (N_22449,N_13070,N_15587);
nand U22450 (N_22450,N_14596,N_13579);
nor U22451 (N_22451,N_16852,N_13014);
nor U22452 (N_22452,N_16744,N_16028);
nor U22453 (N_22453,N_16134,N_13296);
and U22454 (N_22454,N_15441,N_12555);
and U22455 (N_22455,N_17527,N_16076);
or U22456 (N_22456,N_14343,N_14737);
and U22457 (N_22457,N_15012,N_12261);
or U22458 (N_22458,N_16091,N_17645);
nand U22459 (N_22459,N_17951,N_17191);
nand U22460 (N_22460,N_16063,N_16721);
nor U22461 (N_22461,N_17017,N_15894);
nor U22462 (N_22462,N_17290,N_12834);
xnor U22463 (N_22463,N_14768,N_13914);
or U22464 (N_22464,N_14699,N_16257);
nor U22465 (N_22465,N_12680,N_17997);
and U22466 (N_22466,N_12805,N_17238);
or U22467 (N_22467,N_17984,N_15900);
nor U22468 (N_22468,N_12702,N_13406);
nor U22469 (N_22469,N_13385,N_16888);
nor U22470 (N_22470,N_15114,N_13484);
nand U22471 (N_22471,N_14699,N_13293);
and U22472 (N_22472,N_13538,N_14135);
nor U22473 (N_22473,N_17529,N_16996);
nor U22474 (N_22474,N_15878,N_15549);
or U22475 (N_22475,N_13174,N_15528);
nor U22476 (N_22476,N_12508,N_15549);
and U22477 (N_22477,N_14677,N_14339);
nand U22478 (N_22478,N_12235,N_15389);
nand U22479 (N_22479,N_17345,N_15804);
and U22480 (N_22480,N_15400,N_12620);
nor U22481 (N_22481,N_17019,N_14559);
or U22482 (N_22482,N_13344,N_16559);
and U22483 (N_22483,N_17724,N_15534);
nor U22484 (N_22484,N_14865,N_17349);
nand U22485 (N_22485,N_12981,N_15721);
xnor U22486 (N_22486,N_12995,N_16365);
and U22487 (N_22487,N_16603,N_13792);
and U22488 (N_22488,N_13121,N_17395);
or U22489 (N_22489,N_14557,N_16921);
or U22490 (N_22490,N_16008,N_13942);
and U22491 (N_22491,N_15023,N_15126);
nand U22492 (N_22492,N_12299,N_15814);
or U22493 (N_22493,N_16741,N_16224);
nand U22494 (N_22494,N_13869,N_16225);
nand U22495 (N_22495,N_14381,N_13705);
and U22496 (N_22496,N_13195,N_12403);
or U22497 (N_22497,N_17070,N_12693);
nor U22498 (N_22498,N_14414,N_12409);
nand U22499 (N_22499,N_17073,N_17585);
nand U22500 (N_22500,N_16964,N_13128);
nor U22501 (N_22501,N_13981,N_12038);
or U22502 (N_22502,N_14626,N_15602);
or U22503 (N_22503,N_13332,N_16059);
nor U22504 (N_22504,N_17220,N_14696);
nor U22505 (N_22505,N_15101,N_12778);
or U22506 (N_22506,N_15650,N_14724);
nand U22507 (N_22507,N_13602,N_14971);
or U22508 (N_22508,N_12934,N_15274);
xnor U22509 (N_22509,N_14365,N_15834);
and U22510 (N_22510,N_12321,N_12897);
and U22511 (N_22511,N_17536,N_14979);
nand U22512 (N_22512,N_13506,N_14542);
nor U22513 (N_22513,N_12924,N_13145);
or U22514 (N_22514,N_12817,N_17045);
nand U22515 (N_22515,N_12982,N_12213);
or U22516 (N_22516,N_16984,N_13093);
nor U22517 (N_22517,N_15875,N_17486);
xnor U22518 (N_22518,N_16342,N_16985);
and U22519 (N_22519,N_13242,N_15730);
nand U22520 (N_22520,N_15215,N_12603);
nor U22521 (N_22521,N_13433,N_13995);
or U22522 (N_22522,N_14605,N_13800);
nand U22523 (N_22523,N_15486,N_13859);
or U22524 (N_22524,N_17962,N_16276);
xor U22525 (N_22525,N_14501,N_17067);
nand U22526 (N_22526,N_12399,N_13879);
nor U22527 (N_22527,N_15040,N_12724);
nand U22528 (N_22528,N_14227,N_15325);
and U22529 (N_22529,N_14195,N_14918);
and U22530 (N_22530,N_14774,N_14866);
or U22531 (N_22531,N_17702,N_16711);
and U22532 (N_22532,N_16206,N_17465);
and U22533 (N_22533,N_15095,N_12871);
and U22534 (N_22534,N_16745,N_16603);
nand U22535 (N_22535,N_13786,N_12902);
nand U22536 (N_22536,N_15976,N_12586);
nand U22537 (N_22537,N_15990,N_12072);
nand U22538 (N_22538,N_17889,N_17972);
nand U22539 (N_22539,N_12357,N_13941);
nor U22540 (N_22540,N_17749,N_15416);
nand U22541 (N_22541,N_12258,N_12464);
xor U22542 (N_22542,N_14203,N_13781);
nand U22543 (N_22543,N_16149,N_13709);
or U22544 (N_22544,N_16947,N_15914);
nor U22545 (N_22545,N_14598,N_13948);
nand U22546 (N_22546,N_13411,N_15978);
nor U22547 (N_22547,N_13510,N_14022);
and U22548 (N_22548,N_15070,N_12481);
or U22549 (N_22549,N_14553,N_16760);
nand U22550 (N_22550,N_13187,N_15327);
or U22551 (N_22551,N_14354,N_17554);
nand U22552 (N_22552,N_16989,N_17577);
nor U22553 (N_22553,N_15595,N_14138);
nor U22554 (N_22554,N_17120,N_14464);
and U22555 (N_22555,N_13040,N_15293);
nor U22556 (N_22556,N_17480,N_17515);
and U22557 (N_22557,N_13187,N_14289);
nand U22558 (N_22558,N_15136,N_15837);
and U22559 (N_22559,N_15492,N_13005);
nor U22560 (N_22560,N_14418,N_15164);
and U22561 (N_22561,N_16087,N_14929);
or U22562 (N_22562,N_17010,N_15274);
nor U22563 (N_22563,N_14022,N_13219);
nand U22564 (N_22564,N_16905,N_16038);
nor U22565 (N_22565,N_15341,N_16151);
nor U22566 (N_22566,N_13075,N_14430);
or U22567 (N_22567,N_17668,N_15826);
nand U22568 (N_22568,N_16617,N_12556);
nand U22569 (N_22569,N_12209,N_13118);
and U22570 (N_22570,N_13129,N_15904);
nor U22571 (N_22571,N_15592,N_15401);
or U22572 (N_22572,N_16681,N_15870);
xor U22573 (N_22573,N_15308,N_12349);
and U22574 (N_22574,N_12203,N_16771);
or U22575 (N_22575,N_16859,N_12804);
and U22576 (N_22576,N_12679,N_12544);
or U22577 (N_22577,N_17033,N_16314);
nand U22578 (N_22578,N_17480,N_15342);
or U22579 (N_22579,N_12495,N_13352);
and U22580 (N_22580,N_12378,N_13582);
and U22581 (N_22581,N_17287,N_12041);
nand U22582 (N_22582,N_12992,N_12423);
xor U22583 (N_22583,N_16871,N_14470);
nand U22584 (N_22584,N_12263,N_12440);
xnor U22585 (N_22585,N_17702,N_12535);
or U22586 (N_22586,N_12901,N_16668);
nor U22587 (N_22587,N_13736,N_14614);
and U22588 (N_22588,N_12248,N_13391);
and U22589 (N_22589,N_15524,N_12393);
nor U22590 (N_22590,N_15469,N_12587);
xnor U22591 (N_22591,N_14553,N_15876);
or U22592 (N_22592,N_15576,N_14667);
nor U22593 (N_22593,N_15410,N_14557);
and U22594 (N_22594,N_16125,N_12768);
nand U22595 (N_22595,N_13040,N_13678);
or U22596 (N_22596,N_14191,N_16798);
nand U22597 (N_22597,N_15671,N_15184);
or U22598 (N_22598,N_13983,N_13353);
and U22599 (N_22599,N_15260,N_14292);
nand U22600 (N_22600,N_17014,N_13800);
and U22601 (N_22601,N_15806,N_15167);
and U22602 (N_22602,N_14400,N_12877);
and U22603 (N_22603,N_14238,N_14537);
nor U22604 (N_22604,N_14199,N_17835);
nor U22605 (N_22605,N_14835,N_12185);
nor U22606 (N_22606,N_16673,N_14571);
nand U22607 (N_22607,N_15043,N_13577);
nand U22608 (N_22608,N_16173,N_17355);
xor U22609 (N_22609,N_13592,N_17362);
nand U22610 (N_22610,N_15325,N_17440);
or U22611 (N_22611,N_16962,N_13786);
nor U22612 (N_22612,N_15194,N_12143);
xor U22613 (N_22613,N_16680,N_17303);
nand U22614 (N_22614,N_13043,N_13681);
or U22615 (N_22615,N_17197,N_13555);
nor U22616 (N_22616,N_15454,N_17622);
or U22617 (N_22617,N_13802,N_14645);
nor U22618 (N_22618,N_14548,N_16310);
nor U22619 (N_22619,N_12949,N_16215);
nor U22620 (N_22620,N_15225,N_17735);
and U22621 (N_22621,N_14826,N_17928);
or U22622 (N_22622,N_17241,N_17097);
nand U22623 (N_22623,N_12398,N_17980);
nand U22624 (N_22624,N_12193,N_13506);
or U22625 (N_22625,N_15478,N_17199);
nand U22626 (N_22626,N_16948,N_12572);
or U22627 (N_22627,N_13054,N_14141);
nor U22628 (N_22628,N_15330,N_15107);
nand U22629 (N_22629,N_12837,N_16197);
nand U22630 (N_22630,N_17206,N_17284);
and U22631 (N_22631,N_14311,N_16024);
and U22632 (N_22632,N_17013,N_12299);
and U22633 (N_22633,N_16935,N_16909);
or U22634 (N_22634,N_13602,N_12894);
or U22635 (N_22635,N_14550,N_17434);
nand U22636 (N_22636,N_14697,N_14293);
nor U22637 (N_22637,N_16603,N_12305);
xor U22638 (N_22638,N_13488,N_14500);
nand U22639 (N_22639,N_14804,N_14430);
nand U22640 (N_22640,N_14016,N_13766);
xor U22641 (N_22641,N_14466,N_16097);
nor U22642 (N_22642,N_14046,N_17446);
xor U22643 (N_22643,N_12045,N_16978);
xnor U22644 (N_22644,N_14424,N_16356);
nand U22645 (N_22645,N_17845,N_13481);
and U22646 (N_22646,N_15970,N_17524);
nand U22647 (N_22647,N_14115,N_13811);
or U22648 (N_22648,N_14045,N_12260);
and U22649 (N_22649,N_17602,N_13094);
and U22650 (N_22650,N_15418,N_16092);
nor U22651 (N_22651,N_17761,N_15726);
nor U22652 (N_22652,N_13538,N_17710);
and U22653 (N_22653,N_17179,N_15931);
xnor U22654 (N_22654,N_14132,N_14982);
nand U22655 (N_22655,N_15564,N_16845);
or U22656 (N_22656,N_12285,N_15866);
and U22657 (N_22657,N_15672,N_14692);
or U22658 (N_22658,N_13881,N_17617);
nor U22659 (N_22659,N_16350,N_13911);
xnor U22660 (N_22660,N_13938,N_15287);
or U22661 (N_22661,N_14906,N_12777);
nand U22662 (N_22662,N_12637,N_12188);
or U22663 (N_22663,N_16460,N_15979);
or U22664 (N_22664,N_15174,N_13653);
nor U22665 (N_22665,N_17123,N_16580);
or U22666 (N_22666,N_15024,N_17830);
or U22667 (N_22667,N_17376,N_13265);
xor U22668 (N_22668,N_15095,N_13608);
nand U22669 (N_22669,N_17910,N_13372);
nor U22670 (N_22670,N_14118,N_15725);
and U22671 (N_22671,N_15951,N_15965);
nor U22672 (N_22672,N_13633,N_13641);
or U22673 (N_22673,N_14767,N_16107);
xnor U22674 (N_22674,N_16624,N_15629);
nand U22675 (N_22675,N_14778,N_12910);
nor U22676 (N_22676,N_12957,N_16859);
and U22677 (N_22677,N_14234,N_16388);
xor U22678 (N_22678,N_13530,N_16512);
and U22679 (N_22679,N_17394,N_16051);
nand U22680 (N_22680,N_15503,N_12746);
or U22681 (N_22681,N_15464,N_12886);
nand U22682 (N_22682,N_17634,N_12735);
or U22683 (N_22683,N_16094,N_12653);
nand U22684 (N_22684,N_14449,N_12760);
xor U22685 (N_22685,N_16844,N_12430);
nor U22686 (N_22686,N_12635,N_15459);
nand U22687 (N_22687,N_14833,N_16905);
nor U22688 (N_22688,N_15545,N_16297);
nor U22689 (N_22689,N_17718,N_13128);
nor U22690 (N_22690,N_12495,N_13672);
xor U22691 (N_22691,N_16986,N_14082);
or U22692 (N_22692,N_14434,N_17233);
nor U22693 (N_22693,N_13162,N_14806);
nor U22694 (N_22694,N_17922,N_12014);
and U22695 (N_22695,N_16902,N_17098);
nor U22696 (N_22696,N_16004,N_15326);
or U22697 (N_22697,N_17780,N_17183);
xnor U22698 (N_22698,N_14621,N_16938);
nand U22699 (N_22699,N_14276,N_12076);
nor U22700 (N_22700,N_15566,N_17529);
and U22701 (N_22701,N_13742,N_17570);
and U22702 (N_22702,N_13047,N_12697);
or U22703 (N_22703,N_15099,N_14724);
or U22704 (N_22704,N_16754,N_17826);
nand U22705 (N_22705,N_15542,N_12822);
and U22706 (N_22706,N_13341,N_12616);
nor U22707 (N_22707,N_16442,N_17900);
nand U22708 (N_22708,N_17442,N_16567);
or U22709 (N_22709,N_16277,N_12563);
or U22710 (N_22710,N_12308,N_13602);
and U22711 (N_22711,N_16369,N_16218);
and U22712 (N_22712,N_15699,N_15053);
and U22713 (N_22713,N_16534,N_16185);
nand U22714 (N_22714,N_14030,N_15349);
or U22715 (N_22715,N_14698,N_15547);
and U22716 (N_22716,N_13598,N_16004);
xnor U22717 (N_22717,N_12511,N_12024);
or U22718 (N_22718,N_17606,N_13289);
nand U22719 (N_22719,N_12624,N_17107);
nand U22720 (N_22720,N_17395,N_13338);
nand U22721 (N_22721,N_16948,N_13084);
nor U22722 (N_22722,N_17904,N_14114);
or U22723 (N_22723,N_12843,N_14119);
and U22724 (N_22724,N_15659,N_17633);
or U22725 (N_22725,N_14288,N_15505);
or U22726 (N_22726,N_17767,N_13473);
nor U22727 (N_22727,N_13231,N_15323);
or U22728 (N_22728,N_15018,N_13283);
and U22729 (N_22729,N_17422,N_14472);
nand U22730 (N_22730,N_16335,N_15928);
or U22731 (N_22731,N_16944,N_15317);
or U22732 (N_22732,N_13851,N_15773);
xnor U22733 (N_22733,N_12757,N_14641);
and U22734 (N_22734,N_13303,N_12954);
nand U22735 (N_22735,N_17990,N_17691);
nand U22736 (N_22736,N_15864,N_15442);
nand U22737 (N_22737,N_12446,N_13375);
nor U22738 (N_22738,N_13956,N_13116);
or U22739 (N_22739,N_16355,N_15132);
and U22740 (N_22740,N_13140,N_16241);
nor U22741 (N_22741,N_12438,N_16552);
xor U22742 (N_22742,N_12388,N_17202);
or U22743 (N_22743,N_14420,N_16926);
or U22744 (N_22744,N_12667,N_13156);
and U22745 (N_22745,N_15973,N_14137);
and U22746 (N_22746,N_14816,N_17453);
and U22747 (N_22747,N_12393,N_12884);
or U22748 (N_22748,N_14473,N_13850);
nand U22749 (N_22749,N_17142,N_13269);
nor U22750 (N_22750,N_16654,N_14723);
nor U22751 (N_22751,N_17618,N_14085);
nand U22752 (N_22752,N_16054,N_16222);
nor U22753 (N_22753,N_17107,N_14468);
and U22754 (N_22754,N_15628,N_16499);
or U22755 (N_22755,N_15964,N_13529);
and U22756 (N_22756,N_14584,N_16599);
or U22757 (N_22757,N_15647,N_13238);
and U22758 (N_22758,N_15458,N_17427);
nand U22759 (N_22759,N_13131,N_16638);
and U22760 (N_22760,N_12839,N_14046);
and U22761 (N_22761,N_15447,N_13684);
and U22762 (N_22762,N_16281,N_15979);
xnor U22763 (N_22763,N_17605,N_17192);
xnor U22764 (N_22764,N_12984,N_13103);
nor U22765 (N_22765,N_17036,N_17045);
and U22766 (N_22766,N_17784,N_15924);
and U22767 (N_22767,N_12632,N_15464);
or U22768 (N_22768,N_17968,N_16690);
and U22769 (N_22769,N_13119,N_14801);
and U22770 (N_22770,N_13072,N_17345);
nor U22771 (N_22771,N_16882,N_13578);
nor U22772 (N_22772,N_12984,N_15253);
nor U22773 (N_22773,N_16587,N_14888);
xnor U22774 (N_22774,N_16772,N_12015);
or U22775 (N_22775,N_16963,N_13385);
nand U22776 (N_22776,N_17106,N_13497);
or U22777 (N_22777,N_16760,N_15847);
and U22778 (N_22778,N_14625,N_17686);
nor U22779 (N_22779,N_14690,N_16960);
and U22780 (N_22780,N_14111,N_16805);
nand U22781 (N_22781,N_16603,N_15849);
nand U22782 (N_22782,N_12148,N_13822);
and U22783 (N_22783,N_14518,N_17081);
or U22784 (N_22784,N_17568,N_13677);
xor U22785 (N_22785,N_14600,N_12103);
nor U22786 (N_22786,N_15009,N_13496);
and U22787 (N_22787,N_12034,N_17358);
nand U22788 (N_22788,N_14146,N_16576);
xnor U22789 (N_22789,N_16476,N_13443);
nand U22790 (N_22790,N_14565,N_15574);
or U22791 (N_22791,N_16909,N_13496);
and U22792 (N_22792,N_12521,N_16875);
or U22793 (N_22793,N_15645,N_12464);
or U22794 (N_22794,N_14754,N_13195);
nor U22795 (N_22795,N_12553,N_12523);
nand U22796 (N_22796,N_12657,N_15735);
and U22797 (N_22797,N_12562,N_14769);
or U22798 (N_22798,N_12695,N_13449);
and U22799 (N_22799,N_12561,N_12139);
nand U22800 (N_22800,N_12956,N_16571);
and U22801 (N_22801,N_13042,N_13362);
or U22802 (N_22802,N_16376,N_15563);
nor U22803 (N_22803,N_13574,N_17460);
nor U22804 (N_22804,N_16344,N_13969);
nand U22805 (N_22805,N_17689,N_16380);
nand U22806 (N_22806,N_17777,N_13293);
nand U22807 (N_22807,N_12376,N_17819);
and U22808 (N_22808,N_15266,N_15699);
nand U22809 (N_22809,N_12752,N_15908);
nand U22810 (N_22810,N_16348,N_13182);
nand U22811 (N_22811,N_16407,N_16899);
nand U22812 (N_22812,N_12864,N_15557);
or U22813 (N_22813,N_17720,N_16963);
nand U22814 (N_22814,N_15802,N_13156);
or U22815 (N_22815,N_14990,N_13295);
or U22816 (N_22816,N_12681,N_14440);
and U22817 (N_22817,N_13687,N_12029);
xnor U22818 (N_22818,N_15202,N_16021);
or U22819 (N_22819,N_13170,N_15930);
or U22820 (N_22820,N_17787,N_12885);
xor U22821 (N_22821,N_15870,N_15690);
nand U22822 (N_22822,N_16123,N_13580);
nor U22823 (N_22823,N_17423,N_14802);
or U22824 (N_22824,N_15146,N_12791);
and U22825 (N_22825,N_17951,N_17989);
nor U22826 (N_22826,N_14981,N_14235);
and U22827 (N_22827,N_17821,N_16801);
nor U22828 (N_22828,N_15291,N_17505);
nor U22829 (N_22829,N_15528,N_13157);
and U22830 (N_22830,N_15197,N_16329);
xnor U22831 (N_22831,N_17339,N_16143);
or U22832 (N_22832,N_12861,N_17887);
and U22833 (N_22833,N_15022,N_14705);
nor U22834 (N_22834,N_17009,N_16014);
or U22835 (N_22835,N_16802,N_14899);
or U22836 (N_22836,N_16197,N_14246);
and U22837 (N_22837,N_16521,N_12285);
nand U22838 (N_22838,N_14778,N_16298);
or U22839 (N_22839,N_14763,N_16327);
or U22840 (N_22840,N_17565,N_17988);
and U22841 (N_22841,N_12243,N_13114);
or U22842 (N_22842,N_14404,N_15088);
xor U22843 (N_22843,N_13222,N_15552);
nand U22844 (N_22844,N_13790,N_17343);
nand U22845 (N_22845,N_15972,N_13057);
nand U22846 (N_22846,N_12600,N_16658);
nor U22847 (N_22847,N_16842,N_12735);
nand U22848 (N_22848,N_12123,N_16241);
or U22849 (N_22849,N_12555,N_15168);
nor U22850 (N_22850,N_14214,N_15115);
or U22851 (N_22851,N_12559,N_14751);
nor U22852 (N_22852,N_17529,N_17394);
nand U22853 (N_22853,N_13576,N_17270);
nand U22854 (N_22854,N_14588,N_12989);
and U22855 (N_22855,N_12928,N_16727);
and U22856 (N_22856,N_14535,N_16351);
or U22857 (N_22857,N_15455,N_14767);
or U22858 (N_22858,N_17810,N_14441);
nand U22859 (N_22859,N_12597,N_13342);
xor U22860 (N_22860,N_16843,N_12172);
nor U22861 (N_22861,N_14521,N_12378);
or U22862 (N_22862,N_12830,N_17683);
nand U22863 (N_22863,N_12566,N_16542);
or U22864 (N_22864,N_15094,N_17955);
or U22865 (N_22865,N_14838,N_14809);
xor U22866 (N_22866,N_17683,N_15312);
nand U22867 (N_22867,N_17484,N_17698);
or U22868 (N_22868,N_13549,N_15386);
or U22869 (N_22869,N_13091,N_14753);
or U22870 (N_22870,N_12371,N_12944);
nor U22871 (N_22871,N_16969,N_16507);
xor U22872 (N_22872,N_15506,N_13057);
xor U22873 (N_22873,N_14153,N_13945);
xnor U22874 (N_22874,N_13314,N_12622);
and U22875 (N_22875,N_12939,N_17111);
nand U22876 (N_22876,N_12324,N_16356);
xnor U22877 (N_22877,N_13233,N_16757);
nor U22878 (N_22878,N_12787,N_17898);
nand U22879 (N_22879,N_15903,N_14160);
xor U22880 (N_22880,N_15764,N_13172);
and U22881 (N_22881,N_17981,N_13408);
nand U22882 (N_22882,N_16395,N_12364);
or U22883 (N_22883,N_15797,N_14428);
nor U22884 (N_22884,N_17191,N_15674);
or U22885 (N_22885,N_15072,N_12397);
or U22886 (N_22886,N_15413,N_13147);
nor U22887 (N_22887,N_17330,N_12757);
nor U22888 (N_22888,N_15103,N_13412);
xor U22889 (N_22889,N_15891,N_16012);
nor U22890 (N_22890,N_13356,N_14474);
or U22891 (N_22891,N_17619,N_13143);
nand U22892 (N_22892,N_16220,N_15089);
or U22893 (N_22893,N_17204,N_17197);
nor U22894 (N_22894,N_16939,N_12804);
nor U22895 (N_22895,N_14512,N_16851);
nor U22896 (N_22896,N_17932,N_17816);
nand U22897 (N_22897,N_14002,N_15911);
nand U22898 (N_22898,N_15916,N_14240);
nand U22899 (N_22899,N_15229,N_16366);
nand U22900 (N_22900,N_13031,N_14304);
xnor U22901 (N_22901,N_15914,N_17368);
nor U22902 (N_22902,N_14888,N_14651);
or U22903 (N_22903,N_17849,N_13914);
nor U22904 (N_22904,N_15805,N_12770);
nor U22905 (N_22905,N_13133,N_16880);
nor U22906 (N_22906,N_17727,N_16242);
and U22907 (N_22907,N_14670,N_12115);
nand U22908 (N_22908,N_12698,N_17623);
nor U22909 (N_22909,N_15218,N_12254);
and U22910 (N_22910,N_15497,N_12372);
or U22911 (N_22911,N_12049,N_13002);
nand U22912 (N_22912,N_13679,N_14990);
and U22913 (N_22913,N_16404,N_13929);
nand U22914 (N_22914,N_13073,N_15198);
nand U22915 (N_22915,N_14420,N_14596);
or U22916 (N_22916,N_14932,N_17188);
nor U22917 (N_22917,N_16363,N_12269);
nor U22918 (N_22918,N_12205,N_17168);
nor U22919 (N_22919,N_16412,N_13965);
nand U22920 (N_22920,N_16610,N_15108);
nor U22921 (N_22921,N_16249,N_14207);
or U22922 (N_22922,N_13510,N_15130);
xor U22923 (N_22923,N_14447,N_14921);
nor U22924 (N_22924,N_12320,N_15501);
and U22925 (N_22925,N_17038,N_15372);
and U22926 (N_22926,N_15026,N_12679);
and U22927 (N_22927,N_16470,N_16608);
or U22928 (N_22928,N_13103,N_13716);
nor U22929 (N_22929,N_14508,N_15662);
and U22930 (N_22930,N_12887,N_16266);
nor U22931 (N_22931,N_15562,N_16637);
nand U22932 (N_22932,N_13805,N_16279);
nor U22933 (N_22933,N_16376,N_16522);
nor U22934 (N_22934,N_14199,N_17892);
and U22935 (N_22935,N_17142,N_16731);
nand U22936 (N_22936,N_14457,N_14426);
nand U22937 (N_22937,N_16114,N_14516);
xor U22938 (N_22938,N_16676,N_14035);
or U22939 (N_22939,N_13250,N_13218);
and U22940 (N_22940,N_12073,N_17984);
xor U22941 (N_22941,N_13814,N_12448);
nand U22942 (N_22942,N_12629,N_15857);
and U22943 (N_22943,N_17842,N_13763);
nand U22944 (N_22944,N_15348,N_13069);
and U22945 (N_22945,N_17157,N_16819);
nand U22946 (N_22946,N_14424,N_15483);
nand U22947 (N_22947,N_15319,N_15068);
nor U22948 (N_22948,N_17222,N_16043);
or U22949 (N_22949,N_12085,N_15463);
and U22950 (N_22950,N_17058,N_12772);
nor U22951 (N_22951,N_17025,N_16159);
xor U22952 (N_22952,N_17715,N_15113);
xor U22953 (N_22953,N_14610,N_17676);
nand U22954 (N_22954,N_17401,N_15256);
nand U22955 (N_22955,N_16102,N_16420);
and U22956 (N_22956,N_15630,N_12453);
or U22957 (N_22957,N_13865,N_13027);
xnor U22958 (N_22958,N_14423,N_14926);
and U22959 (N_22959,N_14048,N_15153);
nor U22960 (N_22960,N_17405,N_15351);
and U22961 (N_22961,N_12027,N_12059);
or U22962 (N_22962,N_14631,N_13370);
xor U22963 (N_22963,N_16180,N_15763);
nor U22964 (N_22964,N_14946,N_15332);
or U22965 (N_22965,N_17029,N_16250);
and U22966 (N_22966,N_16197,N_14631);
or U22967 (N_22967,N_14628,N_13377);
nand U22968 (N_22968,N_13378,N_13587);
nor U22969 (N_22969,N_14392,N_12273);
and U22970 (N_22970,N_12490,N_17990);
nor U22971 (N_22971,N_17865,N_12516);
nand U22972 (N_22972,N_17053,N_16936);
and U22973 (N_22973,N_16981,N_15163);
nor U22974 (N_22974,N_16691,N_13293);
nand U22975 (N_22975,N_15930,N_13580);
and U22976 (N_22976,N_12785,N_14773);
or U22977 (N_22977,N_14653,N_16281);
nand U22978 (N_22978,N_17389,N_15332);
and U22979 (N_22979,N_14177,N_17390);
and U22980 (N_22980,N_16216,N_16546);
and U22981 (N_22981,N_14758,N_13895);
and U22982 (N_22982,N_13223,N_17990);
xnor U22983 (N_22983,N_13797,N_17352);
and U22984 (N_22984,N_17192,N_12276);
or U22985 (N_22985,N_15488,N_13785);
xnor U22986 (N_22986,N_17767,N_16794);
and U22987 (N_22987,N_15078,N_14724);
nor U22988 (N_22988,N_15752,N_14856);
nor U22989 (N_22989,N_14869,N_15089);
nor U22990 (N_22990,N_16460,N_13561);
or U22991 (N_22991,N_13299,N_13162);
xor U22992 (N_22992,N_16705,N_14697);
and U22993 (N_22993,N_13330,N_13875);
or U22994 (N_22994,N_14096,N_14721);
and U22995 (N_22995,N_12829,N_13269);
nor U22996 (N_22996,N_15504,N_13307);
or U22997 (N_22997,N_14556,N_15158);
nor U22998 (N_22998,N_12445,N_13271);
or U22999 (N_22999,N_16920,N_17823);
or U23000 (N_23000,N_13256,N_17311);
and U23001 (N_23001,N_16706,N_16042);
or U23002 (N_23002,N_17246,N_16724);
nor U23003 (N_23003,N_14611,N_14907);
and U23004 (N_23004,N_15879,N_15162);
nor U23005 (N_23005,N_16598,N_17890);
or U23006 (N_23006,N_13967,N_14916);
and U23007 (N_23007,N_14238,N_12098);
nor U23008 (N_23008,N_14914,N_17847);
and U23009 (N_23009,N_15479,N_15128);
xor U23010 (N_23010,N_16671,N_12079);
nor U23011 (N_23011,N_14642,N_16079);
nor U23012 (N_23012,N_14348,N_17520);
and U23013 (N_23013,N_16886,N_16213);
or U23014 (N_23014,N_17956,N_13178);
nor U23015 (N_23015,N_15704,N_14891);
and U23016 (N_23016,N_16381,N_17384);
nand U23017 (N_23017,N_15512,N_14651);
or U23018 (N_23018,N_16430,N_13263);
or U23019 (N_23019,N_15294,N_16929);
nor U23020 (N_23020,N_15041,N_14029);
xnor U23021 (N_23021,N_13518,N_13941);
or U23022 (N_23022,N_16982,N_16516);
or U23023 (N_23023,N_17848,N_13729);
xor U23024 (N_23024,N_17269,N_15260);
or U23025 (N_23025,N_12201,N_16692);
nor U23026 (N_23026,N_17179,N_13727);
nor U23027 (N_23027,N_15839,N_13456);
and U23028 (N_23028,N_16615,N_17050);
nand U23029 (N_23029,N_15704,N_17322);
nor U23030 (N_23030,N_14173,N_14867);
and U23031 (N_23031,N_17947,N_15012);
nand U23032 (N_23032,N_12292,N_16834);
and U23033 (N_23033,N_13547,N_12719);
nor U23034 (N_23034,N_16162,N_14668);
or U23035 (N_23035,N_17592,N_14280);
nand U23036 (N_23036,N_14135,N_12013);
nor U23037 (N_23037,N_15733,N_16125);
or U23038 (N_23038,N_17150,N_13986);
and U23039 (N_23039,N_16102,N_13550);
and U23040 (N_23040,N_16081,N_13870);
or U23041 (N_23041,N_13768,N_14255);
nand U23042 (N_23042,N_13117,N_14889);
nand U23043 (N_23043,N_17416,N_14000);
or U23044 (N_23044,N_16979,N_14873);
and U23045 (N_23045,N_15516,N_15984);
or U23046 (N_23046,N_16227,N_17596);
nor U23047 (N_23047,N_17131,N_15955);
nor U23048 (N_23048,N_17700,N_15418);
nor U23049 (N_23049,N_15971,N_17984);
xnor U23050 (N_23050,N_15816,N_13815);
or U23051 (N_23051,N_14923,N_16386);
nand U23052 (N_23052,N_17515,N_14809);
nor U23053 (N_23053,N_16865,N_14362);
and U23054 (N_23054,N_12632,N_13317);
or U23055 (N_23055,N_17764,N_13484);
or U23056 (N_23056,N_16698,N_17515);
and U23057 (N_23057,N_15576,N_16318);
and U23058 (N_23058,N_12861,N_12656);
or U23059 (N_23059,N_16058,N_15847);
and U23060 (N_23060,N_17353,N_16950);
and U23061 (N_23061,N_14462,N_13399);
nor U23062 (N_23062,N_17299,N_13949);
nor U23063 (N_23063,N_14146,N_16996);
nor U23064 (N_23064,N_16310,N_16521);
or U23065 (N_23065,N_12254,N_16373);
nand U23066 (N_23066,N_14649,N_13864);
nor U23067 (N_23067,N_14153,N_14790);
and U23068 (N_23068,N_17652,N_12494);
nor U23069 (N_23069,N_15293,N_17180);
nor U23070 (N_23070,N_16783,N_17662);
nand U23071 (N_23071,N_16438,N_16270);
nor U23072 (N_23072,N_16367,N_16181);
and U23073 (N_23073,N_15942,N_12119);
and U23074 (N_23074,N_14693,N_15730);
nand U23075 (N_23075,N_17267,N_13014);
nand U23076 (N_23076,N_14729,N_12275);
nor U23077 (N_23077,N_13093,N_15595);
and U23078 (N_23078,N_16965,N_12907);
or U23079 (N_23079,N_16342,N_15945);
or U23080 (N_23080,N_14474,N_16752);
and U23081 (N_23081,N_17847,N_13318);
xnor U23082 (N_23082,N_13546,N_12833);
nand U23083 (N_23083,N_13076,N_14662);
and U23084 (N_23084,N_14158,N_16148);
and U23085 (N_23085,N_14667,N_15799);
or U23086 (N_23086,N_16368,N_17143);
and U23087 (N_23087,N_14300,N_16359);
and U23088 (N_23088,N_15263,N_13703);
and U23089 (N_23089,N_12168,N_16296);
or U23090 (N_23090,N_12457,N_13804);
and U23091 (N_23091,N_12888,N_12229);
or U23092 (N_23092,N_14124,N_16273);
or U23093 (N_23093,N_17355,N_17288);
or U23094 (N_23094,N_13860,N_16987);
nor U23095 (N_23095,N_15855,N_12319);
or U23096 (N_23096,N_13670,N_16086);
or U23097 (N_23097,N_16910,N_14198);
or U23098 (N_23098,N_16667,N_14953);
and U23099 (N_23099,N_17530,N_14244);
nand U23100 (N_23100,N_15417,N_15276);
or U23101 (N_23101,N_13121,N_15092);
or U23102 (N_23102,N_14518,N_15846);
and U23103 (N_23103,N_15546,N_13247);
or U23104 (N_23104,N_13646,N_14956);
nor U23105 (N_23105,N_17450,N_14346);
or U23106 (N_23106,N_15010,N_17098);
nand U23107 (N_23107,N_15534,N_13434);
xnor U23108 (N_23108,N_13622,N_13704);
and U23109 (N_23109,N_14932,N_15091);
nand U23110 (N_23110,N_12160,N_15100);
xnor U23111 (N_23111,N_17396,N_14337);
or U23112 (N_23112,N_12118,N_14388);
and U23113 (N_23113,N_17494,N_14755);
and U23114 (N_23114,N_17143,N_17636);
nand U23115 (N_23115,N_17233,N_16787);
nor U23116 (N_23116,N_16172,N_15150);
or U23117 (N_23117,N_16947,N_15270);
nand U23118 (N_23118,N_12019,N_17561);
or U23119 (N_23119,N_15988,N_12462);
and U23120 (N_23120,N_16638,N_13086);
nand U23121 (N_23121,N_12456,N_15901);
or U23122 (N_23122,N_12132,N_17312);
xor U23123 (N_23123,N_14759,N_13602);
and U23124 (N_23124,N_16259,N_14707);
nor U23125 (N_23125,N_14302,N_16859);
xnor U23126 (N_23126,N_15123,N_14412);
nor U23127 (N_23127,N_12958,N_14889);
or U23128 (N_23128,N_17062,N_17516);
nand U23129 (N_23129,N_13517,N_14731);
or U23130 (N_23130,N_14135,N_14166);
nand U23131 (N_23131,N_16048,N_12210);
xnor U23132 (N_23132,N_16560,N_13034);
nand U23133 (N_23133,N_15951,N_13311);
nor U23134 (N_23134,N_17430,N_14000);
and U23135 (N_23135,N_12266,N_12208);
nand U23136 (N_23136,N_12937,N_15741);
nor U23137 (N_23137,N_14291,N_16146);
or U23138 (N_23138,N_13448,N_12438);
nor U23139 (N_23139,N_17111,N_16685);
and U23140 (N_23140,N_16369,N_17496);
nand U23141 (N_23141,N_13472,N_15964);
or U23142 (N_23142,N_12287,N_13523);
nor U23143 (N_23143,N_13201,N_17378);
nor U23144 (N_23144,N_17122,N_17322);
and U23145 (N_23145,N_14730,N_12218);
or U23146 (N_23146,N_16533,N_17560);
nor U23147 (N_23147,N_12308,N_13196);
and U23148 (N_23148,N_16227,N_17787);
nor U23149 (N_23149,N_16096,N_12845);
nor U23150 (N_23150,N_12703,N_16768);
nand U23151 (N_23151,N_13968,N_12079);
and U23152 (N_23152,N_15593,N_16642);
or U23153 (N_23153,N_13428,N_16243);
nand U23154 (N_23154,N_12884,N_12499);
nor U23155 (N_23155,N_14662,N_13522);
nand U23156 (N_23156,N_14039,N_14786);
or U23157 (N_23157,N_15702,N_17343);
nand U23158 (N_23158,N_13478,N_17919);
nand U23159 (N_23159,N_14268,N_17235);
and U23160 (N_23160,N_13960,N_12957);
nand U23161 (N_23161,N_14752,N_17418);
or U23162 (N_23162,N_15925,N_14477);
or U23163 (N_23163,N_17614,N_17140);
and U23164 (N_23164,N_13413,N_16816);
and U23165 (N_23165,N_13523,N_12294);
nor U23166 (N_23166,N_16824,N_17724);
and U23167 (N_23167,N_16425,N_13199);
xor U23168 (N_23168,N_14430,N_12560);
or U23169 (N_23169,N_15160,N_17138);
or U23170 (N_23170,N_14973,N_15144);
and U23171 (N_23171,N_16464,N_13886);
and U23172 (N_23172,N_17474,N_13795);
nand U23173 (N_23173,N_13621,N_16456);
and U23174 (N_23174,N_17501,N_15218);
nand U23175 (N_23175,N_12507,N_13018);
xnor U23176 (N_23176,N_16317,N_12093);
or U23177 (N_23177,N_17950,N_14015);
or U23178 (N_23178,N_15283,N_14875);
xor U23179 (N_23179,N_15032,N_17391);
or U23180 (N_23180,N_12836,N_13747);
nand U23181 (N_23181,N_17374,N_16624);
xor U23182 (N_23182,N_17259,N_14912);
nand U23183 (N_23183,N_15290,N_14327);
xnor U23184 (N_23184,N_17695,N_17411);
nor U23185 (N_23185,N_15709,N_17066);
xnor U23186 (N_23186,N_14197,N_16197);
xnor U23187 (N_23187,N_12352,N_13128);
and U23188 (N_23188,N_15711,N_12246);
or U23189 (N_23189,N_14593,N_12138);
or U23190 (N_23190,N_14728,N_12551);
and U23191 (N_23191,N_14446,N_12905);
nand U23192 (N_23192,N_17124,N_13679);
nor U23193 (N_23193,N_14611,N_14089);
or U23194 (N_23194,N_14689,N_13236);
or U23195 (N_23195,N_14098,N_16123);
nand U23196 (N_23196,N_16299,N_15904);
and U23197 (N_23197,N_12571,N_14291);
nand U23198 (N_23198,N_13809,N_13939);
nand U23199 (N_23199,N_16594,N_16035);
and U23200 (N_23200,N_14567,N_13026);
nor U23201 (N_23201,N_13438,N_14788);
and U23202 (N_23202,N_17876,N_15407);
nand U23203 (N_23203,N_16928,N_13921);
and U23204 (N_23204,N_15897,N_16337);
nand U23205 (N_23205,N_17209,N_16822);
nor U23206 (N_23206,N_16662,N_17584);
xor U23207 (N_23207,N_12982,N_15112);
and U23208 (N_23208,N_13642,N_16342);
or U23209 (N_23209,N_17786,N_14608);
nor U23210 (N_23210,N_13288,N_16391);
and U23211 (N_23211,N_15714,N_12574);
nor U23212 (N_23212,N_14712,N_16675);
or U23213 (N_23213,N_16006,N_14770);
nand U23214 (N_23214,N_15766,N_14929);
or U23215 (N_23215,N_15498,N_13711);
nor U23216 (N_23216,N_17088,N_14193);
and U23217 (N_23217,N_13598,N_12657);
nand U23218 (N_23218,N_13591,N_17937);
nor U23219 (N_23219,N_17731,N_16169);
xnor U23220 (N_23220,N_14155,N_15525);
nor U23221 (N_23221,N_14146,N_17956);
and U23222 (N_23222,N_12643,N_16624);
and U23223 (N_23223,N_17954,N_12633);
nand U23224 (N_23224,N_17928,N_15615);
and U23225 (N_23225,N_14250,N_16802);
or U23226 (N_23226,N_13907,N_15228);
xor U23227 (N_23227,N_16213,N_17947);
xnor U23228 (N_23228,N_12968,N_13263);
nor U23229 (N_23229,N_12538,N_15149);
xnor U23230 (N_23230,N_12236,N_17246);
or U23231 (N_23231,N_17768,N_13090);
nor U23232 (N_23232,N_17209,N_14678);
or U23233 (N_23233,N_16991,N_12374);
nand U23234 (N_23234,N_14170,N_13069);
and U23235 (N_23235,N_12865,N_15542);
and U23236 (N_23236,N_15501,N_15291);
nand U23237 (N_23237,N_15150,N_12740);
nand U23238 (N_23238,N_14586,N_16068);
nand U23239 (N_23239,N_17954,N_14523);
nor U23240 (N_23240,N_15582,N_15387);
nand U23241 (N_23241,N_12471,N_15554);
or U23242 (N_23242,N_13028,N_15446);
nand U23243 (N_23243,N_15602,N_12262);
nand U23244 (N_23244,N_12180,N_17121);
xor U23245 (N_23245,N_16583,N_14343);
nand U23246 (N_23246,N_17955,N_13057);
xnor U23247 (N_23247,N_13349,N_17658);
nand U23248 (N_23248,N_12608,N_14342);
nor U23249 (N_23249,N_12753,N_12352);
and U23250 (N_23250,N_17740,N_12538);
or U23251 (N_23251,N_15037,N_14438);
nand U23252 (N_23252,N_13907,N_15611);
or U23253 (N_23253,N_16925,N_12662);
or U23254 (N_23254,N_16927,N_17819);
and U23255 (N_23255,N_16752,N_16932);
and U23256 (N_23256,N_14560,N_17586);
or U23257 (N_23257,N_13126,N_13204);
nor U23258 (N_23258,N_12950,N_13129);
or U23259 (N_23259,N_12396,N_13600);
and U23260 (N_23260,N_13237,N_13829);
and U23261 (N_23261,N_15980,N_16462);
and U23262 (N_23262,N_16567,N_13546);
or U23263 (N_23263,N_15975,N_14885);
or U23264 (N_23264,N_12843,N_12765);
or U23265 (N_23265,N_16416,N_14190);
nor U23266 (N_23266,N_16725,N_14185);
nand U23267 (N_23267,N_12819,N_12927);
nand U23268 (N_23268,N_15122,N_12010);
xnor U23269 (N_23269,N_14439,N_16513);
nand U23270 (N_23270,N_14124,N_12510);
and U23271 (N_23271,N_14812,N_12818);
nand U23272 (N_23272,N_15135,N_13425);
nor U23273 (N_23273,N_14626,N_16029);
and U23274 (N_23274,N_16002,N_16372);
xnor U23275 (N_23275,N_16004,N_14057);
nor U23276 (N_23276,N_15320,N_12933);
nor U23277 (N_23277,N_13188,N_14538);
nor U23278 (N_23278,N_15796,N_17241);
nand U23279 (N_23279,N_14637,N_16049);
or U23280 (N_23280,N_12902,N_14399);
nand U23281 (N_23281,N_13468,N_12723);
nor U23282 (N_23282,N_15958,N_15695);
or U23283 (N_23283,N_12026,N_17906);
nand U23284 (N_23284,N_15612,N_12770);
nand U23285 (N_23285,N_14765,N_13195);
or U23286 (N_23286,N_16694,N_13044);
or U23287 (N_23287,N_15540,N_13179);
and U23288 (N_23288,N_13451,N_17378);
and U23289 (N_23289,N_17957,N_12048);
nand U23290 (N_23290,N_13328,N_12211);
nand U23291 (N_23291,N_12410,N_13415);
and U23292 (N_23292,N_14511,N_15402);
xor U23293 (N_23293,N_12966,N_16163);
nand U23294 (N_23294,N_13602,N_13423);
or U23295 (N_23295,N_17154,N_14138);
nor U23296 (N_23296,N_13456,N_13846);
nor U23297 (N_23297,N_16260,N_16330);
nand U23298 (N_23298,N_12808,N_13820);
nor U23299 (N_23299,N_12316,N_13078);
or U23300 (N_23300,N_13007,N_17554);
and U23301 (N_23301,N_12510,N_16220);
xor U23302 (N_23302,N_14729,N_17075);
and U23303 (N_23303,N_15993,N_12858);
nor U23304 (N_23304,N_15305,N_17618);
or U23305 (N_23305,N_12995,N_12884);
xnor U23306 (N_23306,N_12462,N_14964);
or U23307 (N_23307,N_13321,N_13835);
or U23308 (N_23308,N_15260,N_16022);
nor U23309 (N_23309,N_12105,N_14874);
or U23310 (N_23310,N_13623,N_15909);
xor U23311 (N_23311,N_16797,N_16623);
nand U23312 (N_23312,N_15556,N_15266);
or U23313 (N_23313,N_17211,N_17537);
nand U23314 (N_23314,N_13563,N_12200);
xnor U23315 (N_23315,N_13760,N_16141);
xnor U23316 (N_23316,N_12829,N_13558);
nor U23317 (N_23317,N_12304,N_16216);
nand U23318 (N_23318,N_15216,N_12927);
nor U23319 (N_23319,N_13687,N_12432);
xor U23320 (N_23320,N_15839,N_15298);
nand U23321 (N_23321,N_16307,N_16552);
nor U23322 (N_23322,N_13628,N_12131);
or U23323 (N_23323,N_16001,N_13966);
and U23324 (N_23324,N_12028,N_17158);
nor U23325 (N_23325,N_16922,N_12993);
nor U23326 (N_23326,N_15368,N_14157);
nand U23327 (N_23327,N_16346,N_16103);
nor U23328 (N_23328,N_12465,N_17472);
nand U23329 (N_23329,N_13164,N_13110);
or U23330 (N_23330,N_15674,N_12511);
and U23331 (N_23331,N_16167,N_16470);
and U23332 (N_23332,N_13745,N_15651);
xor U23333 (N_23333,N_14288,N_12885);
nor U23334 (N_23334,N_15762,N_17654);
or U23335 (N_23335,N_14094,N_15718);
and U23336 (N_23336,N_16738,N_16318);
and U23337 (N_23337,N_14881,N_12311);
nand U23338 (N_23338,N_13578,N_15979);
and U23339 (N_23339,N_15481,N_12286);
xor U23340 (N_23340,N_17228,N_13760);
or U23341 (N_23341,N_13975,N_15029);
or U23342 (N_23342,N_14404,N_12161);
and U23343 (N_23343,N_16922,N_14439);
or U23344 (N_23344,N_14031,N_15953);
and U23345 (N_23345,N_13627,N_13576);
xor U23346 (N_23346,N_16395,N_17423);
nor U23347 (N_23347,N_16869,N_16598);
or U23348 (N_23348,N_13446,N_13003);
and U23349 (N_23349,N_13069,N_17646);
or U23350 (N_23350,N_12143,N_14025);
nor U23351 (N_23351,N_15239,N_15697);
and U23352 (N_23352,N_16104,N_13614);
nor U23353 (N_23353,N_12027,N_17482);
and U23354 (N_23354,N_13526,N_12419);
nand U23355 (N_23355,N_16910,N_14556);
and U23356 (N_23356,N_17752,N_17969);
nor U23357 (N_23357,N_16249,N_17681);
and U23358 (N_23358,N_15959,N_12389);
nor U23359 (N_23359,N_16794,N_14317);
xnor U23360 (N_23360,N_13668,N_17766);
nor U23361 (N_23361,N_13799,N_13342);
xnor U23362 (N_23362,N_12045,N_12709);
xor U23363 (N_23363,N_13121,N_16459);
and U23364 (N_23364,N_12085,N_14008);
or U23365 (N_23365,N_16426,N_12968);
nor U23366 (N_23366,N_17510,N_17272);
nand U23367 (N_23367,N_14009,N_16240);
nor U23368 (N_23368,N_14486,N_15511);
or U23369 (N_23369,N_12906,N_15926);
and U23370 (N_23370,N_17471,N_15765);
and U23371 (N_23371,N_13683,N_15374);
or U23372 (N_23372,N_13886,N_12860);
nor U23373 (N_23373,N_17127,N_17969);
and U23374 (N_23374,N_12839,N_13936);
and U23375 (N_23375,N_17061,N_17440);
or U23376 (N_23376,N_16843,N_14535);
or U23377 (N_23377,N_17440,N_17543);
nand U23378 (N_23378,N_15061,N_14909);
and U23379 (N_23379,N_14387,N_17454);
or U23380 (N_23380,N_12117,N_17148);
or U23381 (N_23381,N_15982,N_12760);
nor U23382 (N_23382,N_16277,N_13548);
nand U23383 (N_23383,N_14716,N_12701);
nand U23384 (N_23384,N_14380,N_13412);
or U23385 (N_23385,N_12857,N_12814);
nand U23386 (N_23386,N_15806,N_14785);
nand U23387 (N_23387,N_15539,N_13886);
and U23388 (N_23388,N_14687,N_15115);
nand U23389 (N_23389,N_17034,N_12946);
or U23390 (N_23390,N_12951,N_13786);
nand U23391 (N_23391,N_12807,N_14219);
and U23392 (N_23392,N_14314,N_17816);
or U23393 (N_23393,N_15791,N_14121);
nand U23394 (N_23394,N_16467,N_16086);
nor U23395 (N_23395,N_13986,N_13040);
nor U23396 (N_23396,N_16099,N_14730);
and U23397 (N_23397,N_15283,N_12650);
or U23398 (N_23398,N_16682,N_16006);
and U23399 (N_23399,N_12787,N_14576);
nand U23400 (N_23400,N_17122,N_13230);
and U23401 (N_23401,N_15117,N_16941);
nor U23402 (N_23402,N_15278,N_12129);
nand U23403 (N_23403,N_15458,N_15825);
or U23404 (N_23404,N_13562,N_17685);
and U23405 (N_23405,N_12626,N_15272);
or U23406 (N_23406,N_14900,N_16773);
and U23407 (N_23407,N_13050,N_17804);
or U23408 (N_23408,N_12635,N_12673);
or U23409 (N_23409,N_16207,N_16246);
nand U23410 (N_23410,N_12696,N_17960);
nor U23411 (N_23411,N_16256,N_12987);
nor U23412 (N_23412,N_15290,N_13087);
nor U23413 (N_23413,N_14932,N_17913);
xnor U23414 (N_23414,N_14473,N_15460);
and U23415 (N_23415,N_17193,N_15979);
xnor U23416 (N_23416,N_12160,N_14123);
and U23417 (N_23417,N_12872,N_14509);
nand U23418 (N_23418,N_15553,N_13571);
and U23419 (N_23419,N_17741,N_16445);
nor U23420 (N_23420,N_16700,N_16374);
or U23421 (N_23421,N_15558,N_17233);
nor U23422 (N_23422,N_13240,N_13723);
nor U23423 (N_23423,N_15201,N_12004);
or U23424 (N_23424,N_14646,N_16115);
or U23425 (N_23425,N_16486,N_17027);
nand U23426 (N_23426,N_15798,N_13027);
nand U23427 (N_23427,N_16319,N_14294);
nor U23428 (N_23428,N_12777,N_17890);
xor U23429 (N_23429,N_16477,N_13198);
nor U23430 (N_23430,N_15485,N_13420);
and U23431 (N_23431,N_17135,N_15075);
and U23432 (N_23432,N_17666,N_13885);
or U23433 (N_23433,N_14466,N_16320);
or U23434 (N_23434,N_14017,N_16273);
xnor U23435 (N_23435,N_12839,N_13295);
and U23436 (N_23436,N_14978,N_17023);
xnor U23437 (N_23437,N_13302,N_15615);
xor U23438 (N_23438,N_16084,N_14357);
nand U23439 (N_23439,N_13190,N_17931);
and U23440 (N_23440,N_13246,N_13548);
nor U23441 (N_23441,N_15203,N_15945);
nor U23442 (N_23442,N_17672,N_17808);
nor U23443 (N_23443,N_14003,N_13459);
nand U23444 (N_23444,N_17248,N_14508);
and U23445 (N_23445,N_12078,N_12584);
nand U23446 (N_23446,N_14303,N_14949);
nor U23447 (N_23447,N_17333,N_12953);
nor U23448 (N_23448,N_16130,N_14047);
nor U23449 (N_23449,N_14896,N_13265);
nor U23450 (N_23450,N_14328,N_15598);
xnor U23451 (N_23451,N_15949,N_12725);
and U23452 (N_23452,N_12687,N_12612);
nor U23453 (N_23453,N_12220,N_13727);
and U23454 (N_23454,N_12417,N_17674);
and U23455 (N_23455,N_17390,N_13799);
nand U23456 (N_23456,N_15258,N_16270);
nand U23457 (N_23457,N_14411,N_17394);
nor U23458 (N_23458,N_13432,N_16646);
xnor U23459 (N_23459,N_15319,N_17748);
or U23460 (N_23460,N_15828,N_17675);
nand U23461 (N_23461,N_14000,N_14789);
or U23462 (N_23462,N_14814,N_14461);
nand U23463 (N_23463,N_17439,N_16906);
or U23464 (N_23464,N_16880,N_15278);
and U23465 (N_23465,N_15867,N_16662);
nand U23466 (N_23466,N_16716,N_13592);
and U23467 (N_23467,N_12025,N_16996);
and U23468 (N_23468,N_13102,N_12935);
or U23469 (N_23469,N_14275,N_15706);
xor U23470 (N_23470,N_16627,N_15176);
xnor U23471 (N_23471,N_17801,N_16071);
nand U23472 (N_23472,N_16105,N_16303);
nand U23473 (N_23473,N_16458,N_13409);
and U23474 (N_23474,N_16732,N_12227);
nor U23475 (N_23475,N_13519,N_12263);
xor U23476 (N_23476,N_17398,N_16192);
and U23477 (N_23477,N_14962,N_17908);
or U23478 (N_23478,N_17829,N_16283);
or U23479 (N_23479,N_14642,N_12808);
or U23480 (N_23480,N_17782,N_14749);
xnor U23481 (N_23481,N_17315,N_16236);
nand U23482 (N_23482,N_15066,N_15886);
or U23483 (N_23483,N_15602,N_12834);
and U23484 (N_23484,N_17869,N_15078);
and U23485 (N_23485,N_15102,N_17820);
or U23486 (N_23486,N_15022,N_16040);
and U23487 (N_23487,N_17095,N_12737);
xnor U23488 (N_23488,N_16526,N_12147);
nand U23489 (N_23489,N_16315,N_15523);
and U23490 (N_23490,N_17177,N_12713);
or U23491 (N_23491,N_16898,N_14744);
nand U23492 (N_23492,N_13457,N_15992);
nor U23493 (N_23493,N_13570,N_12264);
or U23494 (N_23494,N_17048,N_16604);
and U23495 (N_23495,N_12771,N_15952);
and U23496 (N_23496,N_15347,N_17091);
nand U23497 (N_23497,N_15384,N_15287);
or U23498 (N_23498,N_14482,N_13897);
nor U23499 (N_23499,N_14907,N_13626);
or U23500 (N_23500,N_17235,N_16270);
nor U23501 (N_23501,N_17533,N_12034);
xnor U23502 (N_23502,N_17275,N_15077);
xor U23503 (N_23503,N_13640,N_14468);
xnor U23504 (N_23504,N_12407,N_15303);
and U23505 (N_23505,N_16115,N_12233);
nand U23506 (N_23506,N_17690,N_17169);
and U23507 (N_23507,N_12082,N_14854);
and U23508 (N_23508,N_13439,N_16437);
and U23509 (N_23509,N_15021,N_13363);
or U23510 (N_23510,N_13190,N_15939);
and U23511 (N_23511,N_17605,N_14230);
or U23512 (N_23512,N_12739,N_16413);
nand U23513 (N_23513,N_13166,N_14216);
nor U23514 (N_23514,N_15360,N_16010);
or U23515 (N_23515,N_15238,N_17574);
or U23516 (N_23516,N_12802,N_15723);
or U23517 (N_23517,N_12101,N_17500);
and U23518 (N_23518,N_15070,N_12878);
nor U23519 (N_23519,N_17334,N_14341);
or U23520 (N_23520,N_12659,N_16628);
nor U23521 (N_23521,N_14888,N_14587);
nor U23522 (N_23522,N_17796,N_15320);
or U23523 (N_23523,N_15697,N_13832);
nand U23524 (N_23524,N_16977,N_17475);
or U23525 (N_23525,N_17038,N_15484);
or U23526 (N_23526,N_16771,N_12262);
xor U23527 (N_23527,N_13525,N_13648);
and U23528 (N_23528,N_16358,N_13100);
nor U23529 (N_23529,N_12913,N_17671);
and U23530 (N_23530,N_17922,N_13801);
nand U23531 (N_23531,N_15525,N_17804);
or U23532 (N_23532,N_13972,N_12814);
and U23533 (N_23533,N_15123,N_16526);
xnor U23534 (N_23534,N_13162,N_13703);
nor U23535 (N_23535,N_13175,N_13250);
nand U23536 (N_23536,N_13575,N_15884);
nand U23537 (N_23537,N_12495,N_15468);
or U23538 (N_23538,N_16527,N_15045);
nand U23539 (N_23539,N_17906,N_17291);
nand U23540 (N_23540,N_13164,N_12016);
and U23541 (N_23541,N_14864,N_13645);
nand U23542 (N_23542,N_17067,N_13224);
nor U23543 (N_23543,N_13517,N_17948);
nor U23544 (N_23544,N_17577,N_14453);
nor U23545 (N_23545,N_12922,N_14774);
or U23546 (N_23546,N_15504,N_12849);
nand U23547 (N_23547,N_12015,N_13164);
nand U23548 (N_23548,N_12529,N_17235);
xor U23549 (N_23549,N_15230,N_15778);
nor U23550 (N_23550,N_13208,N_16299);
xor U23551 (N_23551,N_17972,N_16973);
or U23552 (N_23552,N_12033,N_16895);
nand U23553 (N_23553,N_13219,N_14140);
and U23554 (N_23554,N_13804,N_17360);
nand U23555 (N_23555,N_12754,N_12303);
nor U23556 (N_23556,N_13800,N_12087);
xor U23557 (N_23557,N_12924,N_12070);
nor U23558 (N_23558,N_17866,N_13942);
or U23559 (N_23559,N_16086,N_17615);
or U23560 (N_23560,N_16142,N_17106);
and U23561 (N_23561,N_17877,N_16062);
or U23562 (N_23562,N_13062,N_16925);
and U23563 (N_23563,N_14605,N_13127);
nor U23564 (N_23564,N_14477,N_13438);
nor U23565 (N_23565,N_16455,N_15968);
and U23566 (N_23566,N_16851,N_15818);
nand U23567 (N_23567,N_17949,N_12875);
or U23568 (N_23568,N_17740,N_17436);
or U23569 (N_23569,N_12030,N_12823);
nor U23570 (N_23570,N_12809,N_12375);
or U23571 (N_23571,N_15344,N_17859);
nor U23572 (N_23572,N_15281,N_17426);
or U23573 (N_23573,N_17404,N_12335);
xnor U23574 (N_23574,N_17615,N_17630);
nand U23575 (N_23575,N_17413,N_17511);
or U23576 (N_23576,N_16452,N_15058);
and U23577 (N_23577,N_13492,N_12937);
and U23578 (N_23578,N_14446,N_15046);
or U23579 (N_23579,N_15530,N_14844);
or U23580 (N_23580,N_13867,N_13118);
or U23581 (N_23581,N_17593,N_16439);
or U23582 (N_23582,N_17947,N_12009);
and U23583 (N_23583,N_13408,N_15517);
nor U23584 (N_23584,N_14026,N_16947);
or U23585 (N_23585,N_13599,N_14823);
nor U23586 (N_23586,N_15454,N_12706);
or U23587 (N_23587,N_14791,N_14664);
nand U23588 (N_23588,N_15391,N_13286);
xnor U23589 (N_23589,N_13001,N_17606);
and U23590 (N_23590,N_15978,N_13143);
xnor U23591 (N_23591,N_12004,N_12889);
and U23592 (N_23592,N_15259,N_13257);
nand U23593 (N_23593,N_17154,N_12297);
or U23594 (N_23594,N_16596,N_12693);
or U23595 (N_23595,N_12289,N_17226);
and U23596 (N_23596,N_14155,N_15566);
nand U23597 (N_23597,N_17743,N_14216);
and U23598 (N_23598,N_12999,N_12174);
nor U23599 (N_23599,N_13956,N_17318);
nor U23600 (N_23600,N_13216,N_13713);
xnor U23601 (N_23601,N_14471,N_15113);
nor U23602 (N_23602,N_15655,N_14432);
nor U23603 (N_23603,N_14050,N_17498);
nand U23604 (N_23604,N_13516,N_14261);
or U23605 (N_23605,N_15286,N_16366);
and U23606 (N_23606,N_15326,N_15625);
and U23607 (N_23607,N_15616,N_12595);
and U23608 (N_23608,N_16489,N_15865);
or U23609 (N_23609,N_15390,N_13543);
nand U23610 (N_23610,N_17832,N_13021);
or U23611 (N_23611,N_16876,N_16853);
and U23612 (N_23612,N_17374,N_15585);
nand U23613 (N_23613,N_17819,N_17273);
nand U23614 (N_23614,N_13686,N_13750);
and U23615 (N_23615,N_17445,N_12199);
nor U23616 (N_23616,N_15929,N_16030);
or U23617 (N_23617,N_13206,N_12681);
nand U23618 (N_23618,N_14333,N_13888);
or U23619 (N_23619,N_16585,N_15954);
nand U23620 (N_23620,N_12880,N_15496);
and U23621 (N_23621,N_13072,N_14811);
nand U23622 (N_23622,N_15647,N_16254);
and U23623 (N_23623,N_12833,N_16777);
nand U23624 (N_23624,N_15951,N_13175);
or U23625 (N_23625,N_17739,N_17218);
nor U23626 (N_23626,N_15189,N_16736);
or U23627 (N_23627,N_14676,N_17286);
nor U23628 (N_23628,N_14060,N_16238);
and U23629 (N_23629,N_13651,N_12709);
nor U23630 (N_23630,N_16010,N_13731);
xnor U23631 (N_23631,N_17589,N_15291);
nand U23632 (N_23632,N_17939,N_17759);
nor U23633 (N_23633,N_15106,N_12720);
and U23634 (N_23634,N_17280,N_16936);
nor U23635 (N_23635,N_12048,N_16076);
xor U23636 (N_23636,N_13160,N_13300);
nor U23637 (N_23637,N_16966,N_16330);
and U23638 (N_23638,N_16750,N_15405);
nand U23639 (N_23639,N_16749,N_17013);
and U23640 (N_23640,N_16472,N_16684);
and U23641 (N_23641,N_17270,N_13396);
and U23642 (N_23642,N_12399,N_14740);
nor U23643 (N_23643,N_16472,N_17254);
nand U23644 (N_23644,N_12611,N_14633);
or U23645 (N_23645,N_13400,N_16505);
nand U23646 (N_23646,N_14167,N_14716);
nor U23647 (N_23647,N_14123,N_14074);
or U23648 (N_23648,N_17874,N_13686);
nor U23649 (N_23649,N_13336,N_15122);
nand U23650 (N_23650,N_15312,N_13382);
nor U23651 (N_23651,N_14119,N_12484);
or U23652 (N_23652,N_16971,N_17254);
or U23653 (N_23653,N_15891,N_17448);
or U23654 (N_23654,N_12163,N_16730);
nor U23655 (N_23655,N_17447,N_16330);
xor U23656 (N_23656,N_13497,N_17490);
nand U23657 (N_23657,N_12107,N_14529);
nor U23658 (N_23658,N_12358,N_17118);
and U23659 (N_23659,N_12126,N_14407);
nor U23660 (N_23660,N_14220,N_14279);
nor U23661 (N_23661,N_16704,N_12953);
and U23662 (N_23662,N_17232,N_14940);
nand U23663 (N_23663,N_17147,N_13803);
xnor U23664 (N_23664,N_13584,N_14786);
or U23665 (N_23665,N_17651,N_12417);
nand U23666 (N_23666,N_12575,N_12353);
or U23667 (N_23667,N_16654,N_16252);
nand U23668 (N_23668,N_14594,N_17407);
and U23669 (N_23669,N_13502,N_15059);
and U23670 (N_23670,N_12676,N_16556);
and U23671 (N_23671,N_14286,N_14559);
and U23672 (N_23672,N_15672,N_15894);
or U23673 (N_23673,N_16942,N_13114);
xnor U23674 (N_23674,N_14436,N_13249);
xnor U23675 (N_23675,N_15099,N_13390);
xnor U23676 (N_23676,N_13677,N_16738);
nand U23677 (N_23677,N_12734,N_13559);
or U23678 (N_23678,N_15271,N_17800);
nand U23679 (N_23679,N_13494,N_16076);
nor U23680 (N_23680,N_14206,N_15187);
nor U23681 (N_23681,N_12310,N_15373);
xor U23682 (N_23682,N_17045,N_15071);
or U23683 (N_23683,N_17512,N_15705);
xor U23684 (N_23684,N_16726,N_13134);
or U23685 (N_23685,N_14414,N_16030);
or U23686 (N_23686,N_17976,N_17107);
nand U23687 (N_23687,N_13089,N_13408);
and U23688 (N_23688,N_15915,N_14423);
nor U23689 (N_23689,N_16296,N_16190);
or U23690 (N_23690,N_12474,N_16059);
or U23691 (N_23691,N_15408,N_13261);
and U23692 (N_23692,N_15943,N_15541);
xnor U23693 (N_23693,N_12346,N_17051);
or U23694 (N_23694,N_13431,N_13222);
nor U23695 (N_23695,N_17983,N_12171);
nand U23696 (N_23696,N_13988,N_17032);
nand U23697 (N_23697,N_17073,N_16347);
nand U23698 (N_23698,N_15115,N_16020);
or U23699 (N_23699,N_12303,N_17244);
and U23700 (N_23700,N_13536,N_16793);
nor U23701 (N_23701,N_13824,N_16362);
or U23702 (N_23702,N_13526,N_16963);
xor U23703 (N_23703,N_15750,N_16200);
or U23704 (N_23704,N_15090,N_12384);
nor U23705 (N_23705,N_17721,N_14671);
nand U23706 (N_23706,N_15057,N_15407);
and U23707 (N_23707,N_14933,N_14509);
nor U23708 (N_23708,N_13400,N_15149);
nand U23709 (N_23709,N_13677,N_15061);
and U23710 (N_23710,N_16092,N_17715);
nor U23711 (N_23711,N_16951,N_14305);
or U23712 (N_23712,N_15177,N_15990);
nand U23713 (N_23713,N_12998,N_17498);
nor U23714 (N_23714,N_15062,N_15522);
nand U23715 (N_23715,N_15650,N_16762);
nor U23716 (N_23716,N_14962,N_14583);
nand U23717 (N_23717,N_12192,N_15484);
or U23718 (N_23718,N_13258,N_16514);
or U23719 (N_23719,N_13289,N_15090);
nor U23720 (N_23720,N_15708,N_13856);
xnor U23721 (N_23721,N_16709,N_17098);
nor U23722 (N_23722,N_15490,N_13738);
xor U23723 (N_23723,N_14742,N_13555);
or U23724 (N_23724,N_17650,N_12124);
xnor U23725 (N_23725,N_14819,N_15575);
xor U23726 (N_23726,N_12926,N_14174);
or U23727 (N_23727,N_12964,N_15810);
and U23728 (N_23728,N_14665,N_17635);
nor U23729 (N_23729,N_15117,N_17152);
nor U23730 (N_23730,N_15368,N_14106);
or U23731 (N_23731,N_17845,N_13912);
or U23732 (N_23732,N_14448,N_17713);
or U23733 (N_23733,N_15451,N_14911);
and U23734 (N_23734,N_17208,N_17907);
and U23735 (N_23735,N_14218,N_15333);
xnor U23736 (N_23736,N_16211,N_12159);
and U23737 (N_23737,N_12055,N_13590);
nor U23738 (N_23738,N_12305,N_14848);
and U23739 (N_23739,N_12165,N_17880);
nand U23740 (N_23740,N_13897,N_14992);
and U23741 (N_23741,N_12296,N_17819);
nand U23742 (N_23742,N_15581,N_17738);
nand U23743 (N_23743,N_13002,N_12571);
nand U23744 (N_23744,N_13105,N_16377);
nand U23745 (N_23745,N_13167,N_17200);
nand U23746 (N_23746,N_16032,N_17169);
nor U23747 (N_23747,N_15726,N_16626);
xor U23748 (N_23748,N_15271,N_12855);
nor U23749 (N_23749,N_12115,N_15187);
nor U23750 (N_23750,N_16541,N_12810);
and U23751 (N_23751,N_16187,N_13259);
xnor U23752 (N_23752,N_17690,N_16892);
and U23753 (N_23753,N_16535,N_14744);
nor U23754 (N_23754,N_15349,N_14243);
or U23755 (N_23755,N_15706,N_15923);
nor U23756 (N_23756,N_16750,N_15882);
xnor U23757 (N_23757,N_17582,N_16141);
nand U23758 (N_23758,N_12033,N_15564);
nand U23759 (N_23759,N_16286,N_13354);
nor U23760 (N_23760,N_16337,N_17269);
nand U23761 (N_23761,N_13353,N_12833);
and U23762 (N_23762,N_13256,N_16437);
and U23763 (N_23763,N_13360,N_15762);
xor U23764 (N_23764,N_16623,N_14223);
nor U23765 (N_23765,N_17312,N_12967);
nor U23766 (N_23766,N_16609,N_13688);
xnor U23767 (N_23767,N_12516,N_16474);
or U23768 (N_23768,N_12996,N_15703);
and U23769 (N_23769,N_17779,N_12501);
xnor U23770 (N_23770,N_17753,N_15950);
and U23771 (N_23771,N_15942,N_12440);
nor U23772 (N_23772,N_14631,N_13832);
or U23773 (N_23773,N_13892,N_14557);
and U23774 (N_23774,N_15965,N_13052);
and U23775 (N_23775,N_13311,N_14782);
xor U23776 (N_23776,N_13946,N_15975);
and U23777 (N_23777,N_12662,N_15628);
or U23778 (N_23778,N_12108,N_12663);
nor U23779 (N_23779,N_13968,N_16433);
nand U23780 (N_23780,N_16238,N_12443);
or U23781 (N_23781,N_17299,N_14303);
and U23782 (N_23782,N_13202,N_17067);
xnor U23783 (N_23783,N_15183,N_14359);
nor U23784 (N_23784,N_13991,N_16729);
and U23785 (N_23785,N_17233,N_17540);
nor U23786 (N_23786,N_14621,N_12590);
nor U23787 (N_23787,N_15348,N_12182);
xnor U23788 (N_23788,N_13422,N_12291);
nor U23789 (N_23789,N_13344,N_17109);
nand U23790 (N_23790,N_14683,N_16117);
xor U23791 (N_23791,N_14069,N_17541);
and U23792 (N_23792,N_14209,N_16544);
nand U23793 (N_23793,N_13880,N_17806);
xor U23794 (N_23794,N_16035,N_12829);
nand U23795 (N_23795,N_13551,N_14220);
nor U23796 (N_23796,N_14601,N_17966);
nand U23797 (N_23797,N_17404,N_13663);
and U23798 (N_23798,N_15089,N_15015);
nor U23799 (N_23799,N_13689,N_17383);
nand U23800 (N_23800,N_12361,N_17679);
nor U23801 (N_23801,N_16544,N_16188);
nor U23802 (N_23802,N_17106,N_17559);
xnor U23803 (N_23803,N_13781,N_15214);
and U23804 (N_23804,N_12610,N_17847);
nand U23805 (N_23805,N_17782,N_15599);
and U23806 (N_23806,N_14087,N_16644);
or U23807 (N_23807,N_13602,N_17683);
nor U23808 (N_23808,N_15794,N_13610);
nand U23809 (N_23809,N_12840,N_12230);
xnor U23810 (N_23810,N_14854,N_14299);
and U23811 (N_23811,N_14911,N_13606);
and U23812 (N_23812,N_13227,N_15408);
nand U23813 (N_23813,N_16708,N_13771);
nand U23814 (N_23814,N_17648,N_13487);
nor U23815 (N_23815,N_15854,N_17814);
or U23816 (N_23816,N_12900,N_14816);
and U23817 (N_23817,N_15991,N_17070);
or U23818 (N_23818,N_13740,N_14591);
and U23819 (N_23819,N_12277,N_15614);
nor U23820 (N_23820,N_14930,N_17916);
nand U23821 (N_23821,N_14774,N_15669);
and U23822 (N_23822,N_14121,N_14320);
nand U23823 (N_23823,N_17256,N_12745);
and U23824 (N_23824,N_15858,N_14039);
xor U23825 (N_23825,N_16782,N_12900);
nor U23826 (N_23826,N_15581,N_14143);
or U23827 (N_23827,N_12092,N_15486);
nand U23828 (N_23828,N_13594,N_12254);
xor U23829 (N_23829,N_12351,N_17052);
and U23830 (N_23830,N_16787,N_13589);
xnor U23831 (N_23831,N_14747,N_14770);
nor U23832 (N_23832,N_13111,N_13959);
or U23833 (N_23833,N_14007,N_12226);
or U23834 (N_23834,N_15024,N_13948);
or U23835 (N_23835,N_12485,N_15696);
and U23836 (N_23836,N_15612,N_16847);
or U23837 (N_23837,N_17286,N_17180);
nor U23838 (N_23838,N_17782,N_17334);
or U23839 (N_23839,N_16087,N_15232);
xor U23840 (N_23840,N_17515,N_16571);
and U23841 (N_23841,N_14998,N_17577);
nand U23842 (N_23842,N_14508,N_12371);
or U23843 (N_23843,N_16663,N_13160);
nor U23844 (N_23844,N_16872,N_12073);
and U23845 (N_23845,N_12598,N_16637);
and U23846 (N_23846,N_14583,N_13977);
xor U23847 (N_23847,N_15494,N_12865);
nand U23848 (N_23848,N_12698,N_16205);
nand U23849 (N_23849,N_14170,N_15962);
nor U23850 (N_23850,N_16659,N_16336);
nor U23851 (N_23851,N_17970,N_17246);
nor U23852 (N_23852,N_17997,N_15308);
or U23853 (N_23853,N_16450,N_12358);
and U23854 (N_23854,N_16346,N_15183);
nor U23855 (N_23855,N_16625,N_17933);
and U23856 (N_23856,N_13812,N_16166);
nand U23857 (N_23857,N_17164,N_15139);
nor U23858 (N_23858,N_17108,N_17350);
nand U23859 (N_23859,N_14840,N_16631);
xor U23860 (N_23860,N_12662,N_12961);
nand U23861 (N_23861,N_13282,N_16693);
and U23862 (N_23862,N_15380,N_12140);
nor U23863 (N_23863,N_17412,N_16550);
or U23864 (N_23864,N_13808,N_13958);
or U23865 (N_23865,N_15936,N_14794);
or U23866 (N_23866,N_13643,N_15074);
and U23867 (N_23867,N_14516,N_14002);
nand U23868 (N_23868,N_17496,N_14070);
nor U23869 (N_23869,N_15767,N_17285);
nor U23870 (N_23870,N_14487,N_16772);
nor U23871 (N_23871,N_12295,N_16737);
and U23872 (N_23872,N_12965,N_15175);
and U23873 (N_23873,N_16943,N_13906);
and U23874 (N_23874,N_12069,N_17466);
nor U23875 (N_23875,N_17390,N_15000);
nand U23876 (N_23876,N_15842,N_14126);
or U23877 (N_23877,N_14815,N_17100);
nand U23878 (N_23878,N_17473,N_12852);
xnor U23879 (N_23879,N_12390,N_17698);
and U23880 (N_23880,N_16428,N_13246);
nor U23881 (N_23881,N_17495,N_15827);
or U23882 (N_23882,N_15253,N_16511);
nand U23883 (N_23883,N_16659,N_14089);
nand U23884 (N_23884,N_12156,N_17316);
nor U23885 (N_23885,N_16063,N_12616);
nor U23886 (N_23886,N_14392,N_17142);
or U23887 (N_23887,N_13788,N_17924);
or U23888 (N_23888,N_13683,N_15082);
xnor U23889 (N_23889,N_14262,N_12936);
nand U23890 (N_23890,N_17129,N_12816);
or U23891 (N_23891,N_16998,N_16612);
or U23892 (N_23892,N_15244,N_14034);
nand U23893 (N_23893,N_16632,N_17060);
or U23894 (N_23894,N_15726,N_13485);
or U23895 (N_23895,N_13192,N_14278);
nand U23896 (N_23896,N_13740,N_17068);
xor U23897 (N_23897,N_12970,N_13122);
nand U23898 (N_23898,N_16330,N_17225);
nand U23899 (N_23899,N_17033,N_16960);
xor U23900 (N_23900,N_14646,N_17494);
nand U23901 (N_23901,N_13223,N_16510);
and U23902 (N_23902,N_17791,N_16894);
or U23903 (N_23903,N_14711,N_17145);
nor U23904 (N_23904,N_13667,N_14768);
and U23905 (N_23905,N_17050,N_15581);
and U23906 (N_23906,N_12754,N_14149);
nor U23907 (N_23907,N_15160,N_15847);
and U23908 (N_23908,N_16692,N_17809);
or U23909 (N_23909,N_14689,N_15267);
nor U23910 (N_23910,N_14268,N_12175);
xor U23911 (N_23911,N_14477,N_17049);
xor U23912 (N_23912,N_15887,N_13831);
xor U23913 (N_23913,N_16334,N_12237);
nand U23914 (N_23914,N_13024,N_16815);
or U23915 (N_23915,N_14167,N_13551);
xor U23916 (N_23916,N_15130,N_15855);
or U23917 (N_23917,N_14777,N_12689);
and U23918 (N_23918,N_14621,N_17593);
or U23919 (N_23919,N_14767,N_15434);
nor U23920 (N_23920,N_12357,N_13424);
and U23921 (N_23921,N_15234,N_17508);
nor U23922 (N_23922,N_16655,N_14166);
nor U23923 (N_23923,N_16570,N_14884);
nor U23924 (N_23924,N_13136,N_16633);
or U23925 (N_23925,N_15515,N_13042);
or U23926 (N_23926,N_17523,N_15294);
nand U23927 (N_23927,N_16149,N_17914);
nor U23928 (N_23928,N_16719,N_13366);
or U23929 (N_23929,N_13405,N_17475);
nand U23930 (N_23930,N_15487,N_16829);
nand U23931 (N_23931,N_16601,N_16123);
and U23932 (N_23932,N_13017,N_17610);
nor U23933 (N_23933,N_17889,N_14311);
nand U23934 (N_23934,N_16305,N_13543);
and U23935 (N_23935,N_14667,N_13376);
and U23936 (N_23936,N_12234,N_16895);
or U23937 (N_23937,N_15313,N_14049);
nand U23938 (N_23938,N_17961,N_14330);
and U23939 (N_23939,N_13897,N_17900);
nand U23940 (N_23940,N_16758,N_12148);
or U23941 (N_23941,N_14741,N_15688);
nand U23942 (N_23942,N_12026,N_14478);
or U23943 (N_23943,N_15518,N_14358);
or U23944 (N_23944,N_17987,N_14348);
and U23945 (N_23945,N_15322,N_13744);
or U23946 (N_23946,N_17656,N_17216);
nor U23947 (N_23947,N_13405,N_13864);
and U23948 (N_23948,N_13188,N_17667);
nor U23949 (N_23949,N_14328,N_14449);
nand U23950 (N_23950,N_13379,N_13786);
nand U23951 (N_23951,N_12618,N_13361);
or U23952 (N_23952,N_12441,N_12126);
nor U23953 (N_23953,N_17501,N_16970);
or U23954 (N_23954,N_13246,N_17163);
and U23955 (N_23955,N_16531,N_17627);
nor U23956 (N_23956,N_15907,N_14480);
or U23957 (N_23957,N_13561,N_13357);
or U23958 (N_23958,N_15333,N_17697);
nand U23959 (N_23959,N_16542,N_14579);
nand U23960 (N_23960,N_14715,N_17373);
nor U23961 (N_23961,N_13963,N_13419);
and U23962 (N_23962,N_16103,N_14625);
nor U23963 (N_23963,N_17136,N_13777);
nand U23964 (N_23964,N_12884,N_17762);
nor U23965 (N_23965,N_12930,N_13755);
and U23966 (N_23966,N_12758,N_17594);
nor U23967 (N_23967,N_12788,N_14623);
nor U23968 (N_23968,N_14667,N_15465);
nand U23969 (N_23969,N_16893,N_17577);
and U23970 (N_23970,N_13908,N_13963);
nor U23971 (N_23971,N_15347,N_12245);
and U23972 (N_23972,N_12871,N_12248);
or U23973 (N_23973,N_16254,N_14080);
or U23974 (N_23974,N_15325,N_14284);
nand U23975 (N_23975,N_13223,N_16183);
xor U23976 (N_23976,N_13496,N_14179);
nor U23977 (N_23977,N_13466,N_16117);
or U23978 (N_23978,N_14806,N_12532);
and U23979 (N_23979,N_13241,N_16738);
and U23980 (N_23980,N_16779,N_13000);
nor U23981 (N_23981,N_13652,N_15776);
or U23982 (N_23982,N_14563,N_12485);
xnor U23983 (N_23983,N_12026,N_14970);
or U23984 (N_23984,N_14791,N_15451);
and U23985 (N_23985,N_12356,N_12669);
nand U23986 (N_23986,N_13893,N_13725);
nand U23987 (N_23987,N_13481,N_12512);
and U23988 (N_23988,N_12595,N_12496);
and U23989 (N_23989,N_16417,N_15445);
and U23990 (N_23990,N_14261,N_14778);
xnor U23991 (N_23991,N_13832,N_17047);
nor U23992 (N_23992,N_16826,N_14725);
nand U23993 (N_23993,N_16992,N_17944);
or U23994 (N_23994,N_16692,N_12450);
and U23995 (N_23995,N_14793,N_17761);
and U23996 (N_23996,N_17760,N_13121);
xnor U23997 (N_23997,N_12545,N_14860);
xnor U23998 (N_23998,N_17985,N_16032);
or U23999 (N_23999,N_14861,N_15926);
nand U24000 (N_24000,N_22143,N_20040);
nand U24001 (N_24001,N_23651,N_21505);
nor U24002 (N_24002,N_20163,N_18699);
or U24003 (N_24003,N_22200,N_23359);
xor U24004 (N_24004,N_18718,N_18552);
or U24005 (N_24005,N_21020,N_18369);
nor U24006 (N_24006,N_23284,N_22584);
nand U24007 (N_24007,N_21573,N_20593);
or U24008 (N_24008,N_22253,N_18687);
and U24009 (N_24009,N_23518,N_22046);
and U24010 (N_24010,N_18980,N_20223);
nor U24011 (N_24011,N_22088,N_18550);
xnor U24012 (N_24012,N_19322,N_21280);
or U24013 (N_24013,N_18525,N_20601);
and U24014 (N_24014,N_21862,N_20075);
nand U24015 (N_24015,N_20893,N_23537);
nor U24016 (N_24016,N_22328,N_20897);
and U24017 (N_24017,N_19227,N_21756);
or U24018 (N_24018,N_18493,N_19191);
xnor U24019 (N_24019,N_19194,N_21844);
and U24020 (N_24020,N_21256,N_20221);
nor U24021 (N_24021,N_23876,N_18356);
and U24022 (N_24022,N_20395,N_18491);
and U24023 (N_24023,N_19656,N_19504);
nand U24024 (N_24024,N_20311,N_23026);
or U24025 (N_24025,N_22426,N_18436);
nor U24026 (N_24026,N_19458,N_21690);
or U24027 (N_24027,N_21611,N_23423);
and U24028 (N_24028,N_18033,N_21547);
xor U24029 (N_24029,N_22134,N_23633);
nand U24030 (N_24030,N_18285,N_23113);
nor U24031 (N_24031,N_21343,N_18109);
or U24032 (N_24032,N_18524,N_20646);
and U24033 (N_24033,N_20306,N_18795);
or U24034 (N_24034,N_22066,N_21358);
nand U24035 (N_24035,N_21563,N_21203);
nor U24036 (N_24036,N_23390,N_18751);
nor U24037 (N_24037,N_22577,N_20572);
nand U24038 (N_24038,N_20145,N_18926);
nand U24039 (N_24039,N_22551,N_23144);
nor U24040 (N_24040,N_20070,N_23103);
nor U24041 (N_24041,N_22843,N_20976);
nand U24042 (N_24042,N_19556,N_20415);
xor U24043 (N_24043,N_19747,N_21523);
nor U24044 (N_24044,N_22827,N_23279);
or U24045 (N_24045,N_21999,N_20804);
nand U24046 (N_24046,N_20850,N_18603);
nand U24047 (N_24047,N_18511,N_19988);
and U24048 (N_24048,N_20488,N_21994);
nand U24049 (N_24049,N_23757,N_18092);
nand U24050 (N_24050,N_22456,N_21717);
nor U24051 (N_24051,N_21222,N_21646);
nand U24052 (N_24052,N_21527,N_18851);
and U24053 (N_24053,N_23458,N_19996);
and U24054 (N_24054,N_19925,N_18015);
nor U24055 (N_24055,N_20541,N_23678);
nand U24056 (N_24056,N_23072,N_21710);
and U24057 (N_24057,N_20104,N_19992);
and U24058 (N_24058,N_23524,N_18424);
nor U24059 (N_24059,N_22202,N_18238);
nand U24060 (N_24060,N_21040,N_21009);
nand U24061 (N_24061,N_19123,N_18147);
nor U24062 (N_24062,N_22000,N_21148);
nor U24063 (N_24063,N_18024,N_21115);
and U24064 (N_24064,N_23308,N_23219);
nor U24065 (N_24065,N_18573,N_19786);
and U24066 (N_24066,N_23469,N_20180);
nor U24067 (N_24067,N_23092,N_21725);
and U24068 (N_24068,N_22756,N_19290);
or U24069 (N_24069,N_22594,N_21917);
or U24070 (N_24070,N_22842,N_21186);
xor U24071 (N_24071,N_20573,N_19735);
nor U24072 (N_24072,N_22530,N_21403);
and U24073 (N_24073,N_18653,N_18696);
nand U24074 (N_24074,N_19120,N_19644);
nor U24075 (N_24075,N_20041,N_18957);
nand U24076 (N_24076,N_23237,N_21997);
nor U24077 (N_24077,N_21491,N_21220);
nand U24078 (N_24078,N_23886,N_20817);
and U24079 (N_24079,N_18669,N_18518);
nor U24080 (N_24080,N_19528,N_21544);
xnor U24081 (N_24081,N_18277,N_19128);
or U24082 (N_24082,N_22948,N_19985);
nand U24083 (N_24083,N_21194,N_22719);
or U24084 (N_24084,N_18005,N_21159);
nor U24085 (N_24085,N_22888,N_21441);
and U24086 (N_24086,N_18786,N_22159);
nor U24087 (N_24087,N_20014,N_23100);
nand U24088 (N_24088,N_22383,N_21951);
nor U24089 (N_24089,N_18106,N_22668);
and U24090 (N_24090,N_22778,N_19443);
nand U24091 (N_24091,N_21421,N_23869);
nor U24092 (N_24092,N_21883,N_22515);
and U24093 (N_24093,N_23706,N_21109);
nand U24094 (N_24094,N_22512,N_23354);
xnor U24095 (N_24095,N_18812,N_20858);
nand U24096 (N_24096,N_19508,N_19479);
nor U24097 (N_24097,N_23595,N_19400);
nor U24098 (N_24098,N_22701,N_21129);
nor U24099 (N_24099,N_23874,N_21735);
nor U24100 (N_24100,N_23168,N_23720);
and U24101 (N_24101,N_22273,N_18568);
and U24102 (N_24102,N_21977,N_18296);
and U24103 (N_24103,N_22798,N_22228);
nor U24104 (N_24104,N_18040,N_20176);
and U24105 (N_24105,N_21496,N_21528);
nor U24106 (N_24106,N_22607,N_22508);
nor U24107 (N_24107,N_18672,N_22745);
or U24108 (N_24108,N_23663,N_23615);
nor U24109 (N_24109,N_22525,N_19439);
nand U24110 (N_24110,N_21647,N_22186);
nor U24111 (N_24111,N_21378,N_20590);
xor U24112 (N_24112,N_20362,N_19696);
nor U24113 (N_24113,N_22762,N_19608);
or U24114 (N_24114,N_23752,N_19484);
nor U24115 (N_24115,N_22978,N_22680);
and U24116 (N_24116,N_23282,N_19205);
nor U24117 (N_24117,N_21818,N_18788);
nand U24118 (N_24118,N_19064,N_22513);
xnor U24119 (N_24119,N_18947,N_21393);
or U24120 (N_24120,N_22149,N_18304);
or U24121 (N_24121,N_20371,N_23783);
or U24122 (N_24122,N_20607,N_19200);
and U24123 (N_24123,N_19981,N_21036);
nand U24124 (N_24124,N_18251,N_21435);
or U24125 (N_24125,N_20473,N_19975);
and U24126 (N_24126,N_23968,N_22444);
and U24127 (N_24127,N_22960,N_20275);
nand U24128 (N_24128,N_22748,N_23089);
nand U24129 (N_24129,N_23955,N_18260);
or U24130 (N_24130,N_22212,N_19033);
nor U24131 (N_24131,N_19351,N_19095);
nor U24132 (N_24132,N_21352,N_22992);
and U24133 (N_24133,N_23197,N_22464);
nand U24134 (N_24134,N_23393,N_20309);
nor U24135 (N_24135,N_18688,N_21433);
xor U24136 (N_24136,N_18737,N_18708);
and U24137 (N_24137,N_18218,N_19107);
nor U24138 (N_24138,N_22891,N_20592);
and U24139 (N_24139,N_18314,N_22340);
or U24140 (N_24140,N_21254,N_21790);
xor U24141 (N_24141,N_23829,N_19580);
or U24142 (N_24142,N_19715,N_20403);
or U24143 (N_24143,N_22550,N_22575);
nor U24144 (N_24144,N_21512,N_21169);
and U24145 (N_24145,N_23491,N_18281);
or U24146 (N_24146,N_18240,N_23281);
nand U24147 (N_24147,N_23837,N_21426);
xnor U24148 (N_24148,N_22192,N_23149);
nor U24149 (N_24149,N_19264,N_22310);
xnor U24150 (N_24150,N_23713,N_19456);
nand U24151 (N_24151,N_22004,N_20004);
xnor U24152 (N_24152,N_21049,N_20516);
or U24153 (N_24153,N_23966,N_21929);
or U24154 (N_24154,N_20924,N_19089);
nor U24155 (N_24155,N_23351,N_20615);
and U24156 (N_24156,N_19461,N_22103);
nor U24157 (N_24157,N_22029,N_22071);
nand U24158 (N_24158,N_19012,N_22145);
nor U24159 (N_24159,N_19904,N_23724);
nand U24160 (N_24160,N_20860,N_20227);
or U24161 (N_24161,N_19415,N_19815);
nor U24162 (N_24162,N_23055,N_20894);
xor U24163 (N_24163,N_20660,N_21584);
nand U24164 (N_24164,N_18702,N_18585);
and U24165 (N_24165,N_18089,N_22583);
nand U24166 (N_24166,N_22437,N_18482);
nand U24167 (N_24167,N_20661,N_21150);
or U24168 (N_24168,N_23374,N_18685);
nor U24169 (N_24169,N_22611,N_19794);
nand U24170 (N_24170,N_18862,N_18073);
or U24171 (N_24171,N_19687,N_21926);
or U24172 (N_24172,N_22742,N_18198);
and U24173 (N_24173,N_19592,N_19550);
nor U24174 (N_24174,N_23224,N_21861);
and U24175 (N_24175,N_19278,N_19062);
xor U24176 (N_24176,N_19116,N_23930);
nor U24177 (N_24177,N_20792,N_20820);
xnor U24178 (N_24178,N_22276,N_22929);
and U24179 (N_24179,N_18834,N_21726);
xnor U24180 (N_24180,N_23647,N_23261);
or U24181 (N_24181,N_18257,N_20353);
and U24182 (N_24182,N_20768,N_22234);
xnor U24183 (N_24183,N_18084,N_20654);
nor U24184 (N_24184,N_20251,N_21945);
nor U24185 (N_24185,N_23610,N_19811);
nor U24186 (N_24186,N_22334,N_22527);
or U24187 (N_24187,N_19980,N_20803);
xor U24188 (N_24188,N_19006,N_20274);
and U24189 (N_24189,N_23635,N_20891);
or U24190 (N_24190,N_21916,N_21987);
or U24191 (N_24191,N_22519,N_20290);
nand U24192 (N_24192,N_23076,N_20335);
or U24193 (N_24193,N_23420,N_22120);
and U24194 (N_24194,N_20262,N_19094);
or U24195 (N_24195,N_20356,N_22647);
xnor U24196 (N_24196,N_22917,N_23865);
nor U24197 (N_24197,N_19146,N_18102);
nand U24198 (N_24198,N_21503,N_18818);
nand U24199 (N_24199,N_20647,N_22593);
nand U24200 (N_24200,N_18527,N_21759);
nor U24201 (N_24201,N_23022,N_18767);
nand U24202 (N_24202,N_19075,N_18284);
and U24203 (N_24203,N_20605,N_23870);
or U24204 (N_24204,N_18079,N_20732);
nor U24205 (N_24205,N_22191,N_19282);
nor U24206 (N_24206,N_23499,N_20819);
nand U24207 (N_24207,N_20788,N_21811);
or U24208 (N_24208,N_23705,N_22060);
nand U24209 (N_24209,N_22419,N_19713);
and U24210 (N_24210,N_20568,N_21661);
or U24211 (N_24211,N_22546,N_21405);
nor U24212 (N_24212,N_18389,N_20297);
nand U24213 (N_24213,N_23848,N_23441);
or U24214 (N_24214,N_18744,N_21154);
and U24215 (N_24215,N_21117,N_20440);
nand U24216 (N_24216,N_22499,N_22567);
nor U24217 (N_24217,N_18039,N_23943);
nor U24218 (N_24218,N_19192,N_19764);
and U24219 (N_24219,N_18167,N_20463);
xnor U24220 (N_24220,N_18857,N_23685);
nand U24221 (N_24221,N_23266,N_22876);
and U24222 (N_24222,N_20148,N_22396);
or U24223 (N_24223,N_22574,N_18395);
or U24224 (N_24224,N_20324,N_21139);
xnor U24225 (N_24225,N_19664,N_19912);
and U24226 (N_24226,N_23523,N_20310);
nor U24227 (N_24227,N_19701,N_22187);
and U24228 (N_24228,N_23174,N_21940);
nand U24229 (N_24229,N_18557,N_20373);
and U24230 (N_24230,N_18316,N_20898);
or U24231 (N_24231,N_21388,N_22984);
nand U24232 (N_24232,N_22589,N_21114);
and U24233 (N_24233,N_19809,N_20688);
and U24234 (N_24234,N_23856,N_19438);
and U24235 (N_24235,N_19999,N_23327);
or U24236 (N_24236,N_20168,N_21755);
and U24237 (N_24237,N_23127,N_19011);
and U24238 (N_24238,N_21390,N_21263);
nand U24239 (N_24239,N_18155,N_20754);
and U24240 (N_24240,N_23547,N_23937);
and U24241 (N_24241,N_22037,N_21796);
nor U24242 (N_24242,N_19335,N_22799);
nand U24243 (N_24243,N_22372,N_23249);
nor U24244 (N_24244,N_20873,N_22211);
or U24245 (N_24245,N_21011,N_23987);
xor U24246 (N_24246,N_22836,N_20518);
nor U24247 (N_24247,N_18878,N_21093);
nand U24248 (N_24248,N_23861,N_18589);
and U24249 (N_24249,N_19712,N_23689);
nand U24250 (N_24250,N_18308,N_23932);
xnor U24251 (N_24251,N_22613,N_22818);
nor U24252 (N_24252,N_21073,N_21734);
xor U24253 (N_24253,N_22223,N_20971);
and U24254 (N_24254,N_23305,N_22473);
xor U24255 (N_24255,N_18430,N_20825);
nand U24256 (N_24256,N_19787,N_22106);
xnor U24257 (N_24257,N_20095,N_23388);
and U24258 (N_24258,N_20706,N_22664);
nor U24259 (N_24259,N_22727,N_19650);
nor U24260 (N_24260,N_18833,N_23244);
and U24261 (N_24261,N_22774,N_18605);
or U24262 (N_24262,N_22180,N_22715);
and U24263 (N_24263,N_20624,N_21067);
nand U24264 (N_24264,N_19963,N_22353);
nand U24265 (N_24265,N_22216,N_20312);
or U24266 (N_24266,N_19683,N_22706);
or U24267 (N_24267,N_18738,N_20512);
and U24268 (N_24268,N_18866,N_22246);
nor U24269 (N_24269,N_19417,N_18139);
nand U24270 (N_24270,N_22309,N_20442);
nand U24271 (N_24271,N_20955,N_23669);
or U24272 (N_24272,N_18160,N_21655);
nand U24273 (N_24273,N_20332,N_20899);
nor U24274 (N_24274,N_21134,N_23431);
nand U24275 (N_24275,N_22481,N_23812);
or U24276 (N_24276,N_20669,N_22315);
or U24277 (N_24277,N_22123,N_23257);
and U24278 (N_24278,N_22986,N_23295);
and U24279 (N_24279,N_19299,N_23522);
and U24280 (N_24280,N_20038,N_18062);
and U24281 (N_24281,N_19250,N_21122);
nor U24282 (N_24282,N_23950,N_19537);
nand U24283 (N_24283,N_20808,N_18419);
and U24284 (N_24284,N_23508,N_22557);
and U24285 (N_24285,N_21550,N_21166);
nand U24286 (N_24286,N_20695,N_21246);
nor U24287 (N_24287,N_21092,N_20935);
xor U24288 (N_24288,N_23478,N_21449);
or U24289 (N_24289,N_19621,N_20886);
or U24290 (N_24290,N_21319,N_18793);
and U24291 (N_24291,N_22213,N_20492);
or U24292 (N_24292,N_21000,N_20462);
and U24293 (N_24293,N_20635,N_20954);
nand U24294 (N_24294,N_18918,N_19379);
and U24295 (N_24295,N_23403,N_18875);
nand U24296 (N_24296,N_23167,N_20197);
nand U24297 (N_24297,N_21659,N_23915);
nand U24298 (N_24298,N_19475,N_21443);
and U24299 (N_24299,N_21698,N_22003);
and U24300 (N_24300,N_20979,N_20417);
and U24301 (N_24301,N_23065,N_20547);
or U24302 (N_24302,N_19587,N_18533);
or U24303 (N_24303,N_21805,N_23572);
nand U24304 (N_24304,N_21781,N_20677);
nor U24305 (N_24305,N_23992,N_18376);
and U24306 (N_24306,N_22943,N_22666);
xor U24307 (N_24307,N_22453,N_18666);
xor U24308 (N_24308,N_22539,N_18768);
nor U24309 (N_24309,N_23977,N_22327);
nand U24310 (N_24310,N_23655,N_20295);
or U24311 (N_24311,N_21737,N_18811);
nor U24312 (N_24312,N_23083,N_19164);
xnor U24313 (N_24313,N_22823,N_20600);
nor U24314 (N_24314,N_20116,N_18072);
or U24315 (N_24315,N_18655,N_21630);
xor U24316 (N_24316,N_23109,N_22934);
and U24317 (N_24317,N_19202,N_19665);
or U24318 (N_24318,N_20464,N_18633);
nor U24319 (N_24319,N_20617,N_19884);
or U24320 (N_24320,N_23419,N_18108);
nand U24321 (N_24321,N_22829,N_20425);
nand U24322 (N_24322,N_19394,N_19455);
nor U24323 (N_24323,N_21307,N_19406);
nor U24324 (N_24324,N_22402,N_21170);
nor U24325 (N_24325,N_23933,N_21021);
or U24326 (N_24326,N_22714,N_18231);
nor U24327 (N_24327,N_20733,N_21250);
and U24328 (N_24328,N_21185,N_19420);
nor U24329 (N_24329,N_20544,N_19134);
nand U24330 (N_24330,N_21401,N_19676);
or U24331 (N_24331,N_23225,N_20638);
and U24332 (N_24332,N_23521,N_21138);
and U24333 (N_24333,N_18836,N_18402);
or U24334 (N_24334,N_20103,N_22695);
and U24335 (N_24335,N_21764,N_19964);
nor U24336 (N_24336,N_21045,N_22395);
xor U24337 (N_24337,N_23708,N_21869);
nor U24338 (N_24338,N_21809,N_22681);
or U24339 (N_24339,N_20009,N_21095);
and U24340 (N_24340,N_21793,N_21302);
or U24341 (N_24341,N_21498,N_23820);
nor U24342 (N_24342,N_19293,N_21601);
and U24343 (N_24343,N_20080,N_20991);
nand U24344 (N_24344,N_22973,N_20548);
nor U24345 (N_24345,N_20006,N_19234);
nand U24346 (N_24346,N_19396,N_19059);
nand U24347 (N_24347,N_23289,N_22693);
or U24348 (N_24348,N_23033,N_21858);
xor U24349 (N_24349,N_21415,N_18674);
or U24350 (N_24350,N_20459,N_18275);
or U24351 (N_24351,N_20537,N_20652);
or U24352 (N_24352,N_18428,N_22653);
and U24353 (N_24353,N_20880,N_21085);
nor U24354 (N_24354,N_19339,N_21062);
nand U24355 (N_24355,N_22198,N_23749);
nor U24356 (N_24356,N_19101,N_23736);
xnor U24357 (N_24357,N_21489,N_18839);
and U24358 (N_24358,N_19097,N_18606);
or U24359 (N_24359,N_23658,N_20257);
nand U24360 (N_24360,N_18288,N_18394);
or U24361 (N_24361,N_20182,N_22981);
nor U24362 (N_24362,N_22218,N_22835);
and U24363 (N_24363,N_23392,N_19639);
or U24364 (N_24364,N_19703,N_21618);
and U24365 (N_24365,N_23287,N_22313);
or U24366 (N_24366,N_18255,N_19541);
and U24367 (N_24367,N_21189,N_18574);
xor U24368 (N_24368,N_18597,N_18224);
or U24369 (N_24369,N_22887,N_22392);
and U24370 (N_24370,N_21599,N_20179);
and U24371 (N_24371,N_21675,N_19355);
and U24372 (N_24372,N_22980,N_19637);
and U24373 (N_24373,N_18272,N_21003);
nor U24374 (N_24374,N_20158,N_18380);
nor U24375 (N_24375,N_20618,N_20948);
xnor U24376 (N_24376,N_22330,N_23555);
nor U24377 (N_24377,N_21897,N_18298);
nor U24378 (N_24378,N_20937,N_21305);
nor U24379 (N_24379,N_23339,N_19300);
nor U24380 (N_24380,N_21622,N_21824);
nor U24381 (N_24381,N_23074,N_21836);
and U24382 (N_24382,N_20837,N_21943);
and U24383 (N_24383,N_21931,N_19432);
or U24384 (N_24384,N_18270,N_23031);
and U24385 (N_24385,N_22119,N_20591);
nand U24386 (N_24386,N_23021,N_23621);
nor U24387 (N_24387,N_18104,N_21613);
nand U24388 (N_24388,N_19209,N_23200);
and U24389 (N_24389,N_21939,N_23700);
and U24390 (N_24390,N_19180,N_18779);
nor U24391 (N_24391,N_20294,N_18956);
nand U24392 (N_24392,N_19441,N_21668);
or U24393 (N_24393,N_19737,N_22105);
nand U24394 (N_24394,N_20187,N_21090);
nor U24395 (N_24395,N_18991,N_20961);
nand U24396 (N_24396,N_20121,N_21652);
or U24397 (N_24397,N_18127,N_19152);
or U24398 (N_24398,N_21412,N_23426);
nand U24399 (N_24399,N_18888,N_21876);
or U24400 (N_24400,N_23468,N_20322);
nor U24401 (N_24401,N_23411,N_20039);
and U24402 (N_24402,N_18210,N_18520);
nand U24403 (N_24403,N_18826,N_21703);
nand U24404 (N_24404,N_18332,N_18549);
and U24405 (N_24405,N_18010,N_23422);
nand U24406 (N_24406,N_19170,N_23529);
or U24407 (N_24407,N_22840,N_23810);
xor U24408 (N_24408,N_23068,N_18382);
or U24409 (N_24409,N_19700,N_20761);
or U24410 (N_24410,N_23862,N_20444);
and U24411 (N_24411,N_22898,N_19969);
nor U24412 (N_24412,N_23798,N_22906);
nor U24413 (N_24413,N_22744,N_23296);
and U24414 (N_24414,N_19800,N_23479);
nor U24415 (N_24415,N_21476,N_19270);
and U24416 (N_24416,N_20515,N_20623);
nand U24417 (N_24417,N_21979,N_22081);
and U24418 (N_24418,N_22563,N_23911);
or U24419 (N_24419,N_19920,N_18649);
nand U24420 (N_24420,N_21502,N_20017);
nand U24421 (N_24421,N_22290,N_23493);
and U24422 (N_24422,N_18831,N_18982);
and U24423 (N_24423,N_22239,N_22969);
nand U24424 (N_24424,N_22413,N_23527);
nor U24425 (N_24425,N_23201,N_19052);
nand U24426 (N_24426,N_21454,N_22480);
and U24427 (N_24427,N_23541,N_21304);
xnor U24428 (N_24428,N_21721,N_21758);
nor U24429 (N_24429,N_22296,N_21827);
or U24430 (N_24430,N_21413,N_23054);
or U24431 (N_24431,N_21429,N_19524);
nor U24432 (N_24432,N_21656,N_18264);
nand U24433 (N_24433,N_18841,N_18949);
or U24434 (N_24434,N_19574,N_22016);
nor U24435 (N_24435,N_23677,N_20319);
nor U24436 (N_24436,N_22294,N_23385);
nand U24437 (N_24437,N_19416,N_22698);
xnor U24438 (N_24438,N_23583,N_22291);
nor U24439 (N_24439,N_18697,N_18996);
xor U24440 (N_24440,N_22414,N_19341);
and U24441 (N_24441,N_19098,N_18090);
and U24442 (N_24442,N_23566,N_20409);
nor U24443 (N_24443,N_23847,N_20760);
nor U24444 (N_24444,N_21740,N_20926);
nor U24445 (N_24445,N_21341,N_18145);
xor U24446 (N_24446,N_18323,N_20285);
xor U24447 (N_24447,N_19765,N_23676);
nand U24448 (N_24448,N_21484,N_21205);
xor U24449 (N_24449,N_22006,N_18720);
and U24450 (N_24450,N_19544,N_23410);
and U24451 (N_24451,N_21658,N_20633);
xnor U24452 (N_24452,N_18924,N_20222);
or U24453 (N_24453,N_21075,N_22616);
nand U24454 (N_24454,N_22796,N_19359);
nand U24455 (N_24455,N_20670,N_18973);
or U24456 (N_24456,N_21325,N_20918);
nor U24457 (N_24457,N_23459,N_18873);
xor U24458 (N_24458,N_21494,N_22924);
or U24459 (N_24459,N_18769,N_23141);
or U24460 (N_24460,N_19796,N_20149);
and U24461 (N_24461,N_23516,N_19802);
nand U24462 (N_24462,N_19410,N_23640);
nor U24463 (N_24463,N_18785,N_19719);
or U24464 (N_24464,N_22777,N_22788);
xor U24465 (N_24465,N_18704,N_18753);
or U24466 (N_24466,N_19569,N_20342);
or U24467 (N_24467,N_23742,N_21101);
and U24468 (N_24468,N_20922,N_18935);
xor U24469 (N_24469,N_23101,N_18403);
nand U24470 (N_24470,N_21992,N_22516);
nor U24471 (N_24471,N_18012,N_22122);
xnor U24472 (N_24472,N_20479,N_18870);
nand U24473 (N_24473,N_18623,N_20582);
and U24474 (N_24474,N_23412,N_18920);
nand U24475 (N_24475,N_18908,N_23693);
nor U24476 (N_24476,N_18128,N_19869);
xor U24477 (N_24477,N_22990,N_22225);
xor U24478 (N_24478,N_21024,N_21752);
nand U24479 (N_24479,N_22286,N_21568);
nand U24480 (N_24480,N_21142,N_18842);
nor U24481 (N_24481,N_19933,N_23851);
xor U24482 (N_24482,N_19133,N_18679);
nor U24483 (N_24483,N_23438,N_19135);
or U24484 (N_24484,N_20522,N_19588);
xor U24485 (N_24485,N_21176,N_20265);
or U24486 (N_24486,N_20739,N_22832);
nor U24487 (N_24487,N_19636,N_19780);
xnor U24488 (N_24488,N_22112,N_20308);
nor U24489 (N_24489,N_19620,N_18215);
and U24490 (N_24490,N_19433,N_23665);
or U24491 (N_24491,N_19031,N_22250);
and U24492 (N_24492,N_21680,N_23041);
nor U24493 (N_24493,N_23088,N_18684);
xnor U24494 (N_24494,N_22504,N_22966);
nand U24495 (N_24495,N_23975,N_19125);
or U24496 (N_24496,N_21981,N_18921);
nor U24497 (N_24497,N_19077,N_18975);
or U24498 (N_24498,N_22826,N_23983);
xnor U24499 (N_24499,N_19091,N_19552);
or U24500 (N_24500,N_19321,N_23051);
or U24501 (N_24501,N_19598,N_23671);
nand U24502 (N_24502,N_22498,N_20904);
nor U24503 (N_24503,N_22627,N_20982);
nor U24504 (N_24504,N_22749,N_21400);
nand U24505 (N_24505,N_18905,N_21666);
nor U24506 (N_24506,N_19576,N_19855);
nor U24507 (N_24507,N_19888,N_18351);
or U24508 (N_24508,N_22961,N_21697);
or U24509 (N_24509,N_19890,N_19808);
nor U24510 (N_24510,N_19830,N_21389);
xor U24511 (N_24511,N_23451,N_22947);
nor U24512 (N_24512,N_18563,N_21379);
and U24513 (N_24513,N_23883,N_23292);
and U24514 (N_24514,N_20852,N_21417);
and U24515 (N_24515,N_22683,N_21168);
nand U24516 (N_24516,N_18489,N_20244);
nor U24517 (N_24517,N_19944,N_20359);
nand U24518 (N_24518,N_19162,N_18437);
nor U24519 (N_24519,N_21837,N_23242);
and U24520 (N_24520,N_23286,N_19797);
and U24521 (N_24521,N_20723,N_19442);
nand U24522 (N_24522,N_21462,N_18116);
or U24523 (N_24523,N_21113,N_18821);
and U24524 (N_24524,N_18286,N_23122);
and U24525 (N_24525,N_22254,N_23310);
and U24526 (N_24526,N_22388,N_23750);
nor U24527 (N_24527,N_19466,N_21175);
nand U24528 (N_24528,N_20069,N_22758);
and U24529 (N_24529,N_20089,N_21081);
or U24530 (N_24530,N_22457,N_20962);
or U24531 (N_24531,N_23425,N_18388);
nand U24532 (N_24532,N_20186,N_23260);
and U24533 (N_24533,N_19280,N_21806);
and U24534 (N_24534,N_19099,N_22654);
and U24535 (N_24535,N_20558,N_22989);
xnor U24536 (N_24536,N_21171,N_22522);
and U24537 (N_24537,N_18820,N_18750);
and U24538 (N_24538,N_22765,N_22020);
and U24539 (N_24539,N_21161,N_21466);
nor U24540 (N_24540,N_20436,N_23816);
nand U24541 (N_24541,N_23938,N_18640);
and U24542 (N_24542,N_23071,N_22764);
nor U24543 (N_24543,N_20538,N_19088);
nor U24544 (N_24544,N_21475,N_19629);
and U24545 (N_24545,N_20703,N_19363);
nand U24546 (N_24546,N_22013,N_21334);
nor U24547 (N_24547,N_20057,N_22559);
nor U24548 (N_24548,N_22995,N_20764);
or U24549 (N_24549,N_18107,N_20657);
xor U24550 (N_24550,N_19114,N_18060);
nor U24551 (N_24551,N_18301,N_21187);
or U24552 (N_24552,N_18941,N_19225);
nor U24553 (N_24553,N_21718,N_22167);
xnor U24554 (N_24554,N_23680,N_20906);
nand U24555 (N_24555,N_22158,N_18118);
and U24556 (N_24556,N_19345,N_18483);
and U24557 (N_24557,N_23731,N_23220);
or U24558 (N_24558,N_22630,N_20725);
and U24559 (N_24559,N_18006,N_21097);
or U24560 (N_24560,N_18852,N_19886);
or U24561 (N_24561,N_23995,N_19304);
xor U24562 (N_24562,N_19954,N_22824);
xnor U24563 (N_24563,N_19440,N_21603);
nand U24564 (N_24564,N_20200,N_19003);
or U24565 (N_24565,N_22482,N_19388);
nand U24566 (N_24566,N_19242,N_18962);
nor U24567 (N_24567,N_22637,N_22323);
nor U24568 (N_24568,N_22152,N_20491);
and U24569 (N_24569,N_18799,N_18995);
nor U24570 (N_24570,N_20448,N_22976);
xnor U24571 (N_24571,N_22178,N_19983);
nor U24572 (N_24572,N_19269,N_21270);
and U24573 (N_24573,N_22983,N_21266);
xnor U24574 (N_24574,N_18481,N_21531);
xnor U24575 (N_24575,N_20184,N_23118);
xnor U24576 (N_24576,N_19930,N_19942);
nand U24577 (N_24577,N_20468,N_19896);
or U24578 (N_24578,N_23389,N_21792);
or U24579 (N_24579,N_18477,N_19850);
or U24580 (N_24580,N_18173,N_23205);
or U24581 (N_24581,N_19543,N_19389);
or U24582 (N_24582,N_22168,N_21448);
or U24583 (N_24583,N_21530,N_20779);
nand U24584 (N_24584,N_22270,N_20799);
and U24585 (N_24585,N_19086,N_18840);
nand U24586 (N_24586,N_20471,N_19470);
nand U24587 (N_24587,N_19469,N_21165);
nand U24588 (N_24588,N_19903,N_23085);
nor U24589 (N_24589,N_19326,N_20508);
xnor U24590 (N_24590,N_21849,N_20164);
or U24591 (N_24591,N_20741,N_22407);
nand U24592 (N_24592,N_23195,N_19902);
nand U24593 (N_24593,N_19693,N_20445);
nor U24594 (N_24594,N_23276,N_21229);
or U24595 (N_24595,N_23790,N_21933);
nand U24596 (N_24596,N_23391,N_23058);
nor U24597 (N_24597,N_23871,N_19691);
nor U24598 (N_24598,N_18249,N_22580);
or U24599 (N_24599,N_20721,N_22118);
nand U24600 (N_24600,N_20305,N_20950);
nor U24601 (N_24601,N_19295,N_23312);
nand U24602 (N_24602,N_22502,N_21200);
and U24603 (N_24603,N_22677,N_19739);
nand U24604 (N_24604,N_20875,N_22204);
nand U24605 (N_24605,N_22136,N_18410);
nor U24606 (N_24606,N_23002,N_22855);
nor U24607 (N_24607,N_18582,N_20698);
and U24608 (N_24608,N_18783,N_21089);
or U24609 (N_24609,N_18627,N_19292);
nor U24610 (N_24610,N_18338,N_18321);
or U24611 (N_24611,N_21609,N_20361);
nand U24612 (N_24612,N_23573,N_20636);
and U24613 (N_24613,N_23698,N_21451);
nand U24614 (N_24614,N_23802,N_23780);
xnor U24615 (N_24615,N_20055,N_18282);
nand U24616 (N_24616,N_18578,N_22977);
nor U24617 (N_24617,N_19881,N_23519);
nor U24618 (N_24618,N_19667,N_18148);
nand U24619 (N_24619,N_22345,N_20389);
or U24620 (N_24620,N_20869,N_23035);
nor U24621 (N_24621,N_21214,N_21387);
or U24622 (N_24622,N_22874,N_21514);
xnor U24623 (N_24623,N_21960,N_20836);
nor U24624 (N_24624,N_21991,N_18567);
nor U24625 (N_24625,N_23733,N_18576);
or U24626 (N_24626,N_19061,N_19229);
and U24627 (N_24627,N_18273,N_21007);
and U24628 (N_24628,N_19478,N_21553);
nand U24629 (N_24629,N_22586,N_22130);
and U24630 (N_24630,N_21794,N_23512);
and U24631 (N_24631,N_23809,N_21495);
or U24632 (N_24632,N_18522,N_18928);
nor U24633 (N_24633,N_20071,N_18103);
xnor U24634 (N_24634,N_22387,N_18446);
or U24635 (N_24635,N_22803,N_20242);
nand U24636 (N_24636,N_18584,N_23878);
and U24637 (N_24637,N_19889,N_21232);
xnor U24638 (N_24638,N_20120,N_20499);
nor U24639 (N_24639,N_22189,N_18223);
nor U24640 (N_24640,N_19601,N_19661);
or U24641 (N_24641,N_19414,N_19217);
and U24642 (N_24642,N_22148,N_19392);
or U24643 (N_24643,N_23639,N_20790);
nor U24644 (N_24644,N_21900,N_20431);
or U24645 (N_24645,N_18137,N_19894);
nand U24646 (N_24646,N_19685,N_19378);
nand U24647 (N_24647,N_23817,N_22779);
or U24648 (N_24648,N_18521,N_23513);
nor U24649 (N_24649,N_19327,N_23526);
or U24650 (N_24650,N_20801,N_21969);
xor U24651 (N_24651,N_21966,N_22236);
or U24652 (N_24652,N_22787,N_19843);
or U24653 (N_24653,N_21754,N_21519);
nor U24654 (N_24654,N_23177,N_20390);
or U24655 (N_24655,N_21446,N_19273);
nand U24656 (N_24656,N_20291,N_18004);
and U24657 (N_24657,N_21303,N_22650);
nand U24658 (N_24658,N_21286,N_18462);
or U24659 (N_24659,N_21577,N_18721);
xor U24660 (N_24660,N_19418,N_19235);
or U24661 (N_24661,N_21155,N_20901);
nand U24662 (N_24662,N_18199,N_22051);
nand U24663 (N_24663,N_21641,N_18650);
nor U24664 (N_24664,N_22126,N_23716);
xnor U24665 (N_24665,N_19010,N_23417);
nand U24666 (N_24666,N_22679,N_23234);
or U24667 (N_24667,N_19181,N_20997);
nor U24668 (N_24668,N_21582,N_18994);
or U24669 (N_24669,N_21571,N_21911);
nand U24670 (N_24670,N_23066,N_23472);
or U24671 (N_24671,N_21469,N_20671);
or U24672 (N_24672,N_23466,N_22467);
nand U24673 (N_24673,N_18064,N_21207);
and U24674 (N_24674,N_21932,N_20815);
nand U24675 (N_24675,N_18624,N_18115);
and U24676 (N_24676,N_19934,N_23563);
or U24677 (N_24677,N_18318,N_18987);
xor U24678 (N_24678,N_19434,N_18228);
nand U24679 (N_24679,N_19605,N_21340);
nand U24680 (N_24680,N_23495,N_21416);
nand U24681 (N_24681,N_18887,N_18754);
and U24682 (N_24682,N_19305,N_19654);
nand U24683 (N_24683,N_18731,N_18313);
nand U24684 (N_24684,N_21082,N_20236);
or U24685 (N_24685,N_20169,N_18536);
nand U24686 (N_24686,N_18871,N_20493);
nand U24687 (N_24687,N_20243,N_23578);
and U24688 (N_24688,N_23165,N_20778);
nand U24689 (N_24689,N_19195,N_19251);
nand U24690 (N_24690,N_19361,N_18423);
or U24691 (N_24691,N_18561,N_19510);
nand U24692 (N_24692,N_21749,N_18890);
and U24693 (N_24693,N_21673,N_19928);
nor U24694 (N_24694,N_18844,N_23487);
xor U24695 (N_24695,N_18401,N_18637);
or U24696 (N_24696,N_21453,N_20855);
or U24697 (N_24697,N_22114,N_21423);
nor U24698 (N_24698,N_19677,N_18805);
nor U24699 (N_24699,N_20822,N_22640);
nor U24700 (N_24700,N_23363,N_21606);
and U24701 (N_24701,N_18989,N_21975);
or U24702 (N_24702,N_20005,N_18448);
nand U24703 (N_24703,N_21654,N_22510);
or U24704 (N_24704,N_18174,N_22865);
or U24705 (N_24705,N_22099,N_21288);
or U24706 (N_24706,N_23971,N_19130);
or U24707 (N_24707,N_23903,N_20456);
nor U24708 (N_24708,N_22012,N_19854);
or U24709 (N_24709,N_18706,N_19558);
or U24710 (N_24710,N_21110,N_20810);
nor U24711 (N_24711,N_18938,N_18782);
and U24712 (N_24712,N_20367,N_23046);
or U24713 (N_24713,N_22802,N_19773);
nand U24714 (N_24714,N_22951,N_18752);
nor U24715 (N_24715,N_23936,N_18464);
xnor U24716 (N_24716,N_19401,N_19518);
and U24717 (N_24717,N_19697,N_21136);
xor U24718 (N_24718,N_23835,N_22955);
nor U24719 (N_24719,N_23759,N_21241);
nor U24720 (N_24720,N_20846,N_20694);
and U24721 (N_24721,N_21671,N_21013);
nand U24722 (N_24722,N_23213,N_19371);
or U24723 (N_24723,N_22602,N_22804);
nor U24724 (N_24724,N_18345,N_23766);
or U24725 (N_24725,N_22825,N_23806);
nand U24726 (N_24726,N_20051,N_22182);
xor U24727 (N_24727,N_19680,N_22565);
nor U24728 (N_24728,N_22019,N_20237);
nand U24729 (N_24729,N_21464,N_18003);
and U24730 (N_24730,N_18170,N_18189);
nand U24731 (N_24731,N_21619,N_23474);
or U24732 (N_24732,N_20890,N_19505);
nand U24733 (N_24733,N_22878,N_22370);
xor U24734 (N_24734,N_19806,N_21026);
nand U24735 (N_24735,N_23427,N_18848);
nor U24736 (N_24736,N_18580,N_20263);
and U24737 (N_24737,N_21258,N_19210);
or U24738 (N_24738,N_23991,N_21330);
and U24739 (N_24739,N_23607,N_23970);
nor U24740 (N_24740,N_22335,N_18735);
or U24741 (N_24741,N_18474,N_22449);
and U24742 (N_24742,N_18670,N_18440);
nand U24743 (N_24743,N_21889,N_20159);
xnor U24744 (N_24744,N_23357,N_21653);
or U24745 (N_24745,N_20749,N_23553);
and U24746 (N_24746,N_20108,N_22177);
xnor U24747 (N_24747,N_19253,N_23447);
and U24748 (N_24748,N_23320,N_23381);
xor U24749 (N_24749,N_22311,N_18449);
nor U24750 (N_24750,N_20313,N_18097);
nand U24751 (N_24751,N_23232,N_22085);
nand U24752 (N_24752,N_19173,N_23247);
nor U24753 (N_24753,N_18059,N_21976);
and U24754 (N_24754,N_21868,N_21834);
or U24755 (N_24755,N_18607,N_20967);
nand U24756 (N_24756,N_18384,N_23931);
and U24757 (N_24757,N_23134,N_20928);
and U24758 (N_24758,N_22684,N_21875);
or U24759 (N_24759,N_23015,N_18562);
nand U24760 (N_24760,N_20876,N_21339);
nor U24761 (N_24761,N_23335,N_21585);
nor U24762 (N_24762,N_22107,N_21284);
xor U24763 (N_24763,N_23845,N_20023);
xnor U24764 (N_24764,N_22044,N_19138);
nor U24765 (N_24765,N_22900,N_23044);
xor U24766 (N_24766,N_19147,N_22588);
and U24767 (N_24767,N_23952,N_23446);
or U24768 (N_24768,N_18029,N_19947);
and U24769 (N_24769,N_21276,N_23227);
and U24770 (N_24770,N_20958,N_21799);
xor U24771 (N_24771,N_22700,N_21409);
and U24772 (N_24772,N_19435,N_23407);
nor U24773 (N_24773,N_19198,N_22027);
or U24774 (N_24774,N_21457,N_20727);
or U24775 (N_24775,N_23908,N_21572);
nand U24776 (N_24776,N_22894,N_18558);
and U24777 (N_24777,N_23329,N_19929);
nand U24778 (N_24778,N_21111,N_20433);
nand U24779 (N_24779,N_21785,N_22185);
nand U24780 (N_24780,N_23979,N_23603);
and U24781 (N_24781,N_20963,N_22406);
and U24782 (N_24782,N_20514,N_19953);
and U24783 (N_24783,N_23138,N_19990);
and U24784 (N_24784,N_20224,N_21615);
nand U24785 (N_24785,N_19641,N_20198);
or U24786 (N_24786,N_23444,N_19021);
and U24787 (N_24787,N_21455,N_20859);
nand U24788 (N_24788,N_19041,N_23501);
nor U24789 (N_24789,N_18480,N_21950);
or U24790 (N_24790,N_18807,N_18796);
or U24791 (N_24791,N_23365,N_20386);
nand U24792 (N_24792,N_22780,N_20765);
or U24793 (N_24793,N_23557,N_20602);
or U24794 (N_24794,N_19474,N_21346);
or U24795 (N_24795,N_22624,N_18343);
xor U24796 (N_24796,N_21775,N_19705);
and U24797 (N_24797,N_19237,N_21391);
nor U24798 (N_24798,N_19143,N_18978);
and U24799 (N_24799,N_23852,N_20135);
or U24800 (N_24800,N_22753,N_20715);
or U24801 (N_24801,N_21076,N_18478);
nand U24802 (N_24802,N_22558,N_19267);
or U24803 (N_24803,N_18268,N_21716);
nand U24804 (N_24804,N_21487,N_23695);
nand U24805 (N_24805,N_22572,N_21102);
and U24806 (N_24806,N_18140,N_23872);
nor U24807 (N_24807,N_19065,N_19666);
nand U24808 (N_24808,N_21182,N_22466);
nor U24809 (N_24809,N_23670,N_19437);
xor U24810 (N_24810,N_20049,N_22768);
and U24811 (N_24811,N_18011,N_23818);
nand U24812 (N_24812,N_23299,N_22321);
and U24813 (N_24813,N_21427,N_22626);
and U24814 (N_24814,N_20497,N_22628);
or U24815 (N_24815,N_21993,N_22389);
nand U24816 (N_24816,N_22484,N_19917);
nand U24817 (N_24817,N_22600,N_23973);
nand U24818 (N_24818,N_20970,N_21878);
or U24819 (N_24819,N_19916,N_20533);
nor U24820 (N_24820,N_23214,N_18049);
or U24821 (N_24821,N_19426,N_23293);
nor U24822 (N_24822,N_18432,N_19531);
or U24823 (N_24823,N_21551,N_20844);
or U24824 (N_24824,N_23542,N_19613);
and U24825 (N_24825,N_18258,N_20466);
and U24826 (N_24826,N_19647,N_22262);
or U24827 (N_24827,N_20323,N_21414);
nand U24828 (N_24828,N_23823,N_19575);
nand U24829 (N_24829,N_19709,N_18013);
or U24830 (N_24830,N_18066,N_20011);
nand U24831 (N_24831,N_20532,N_23888);
or U24832 (N_24832,N_18484,N_23785);
nand U24833 (N_24833,N_22493,N_19213);
or U24834 (N_24834,N_20705,N_21404);
nor U24835 (N_24835,N_21635,N_23687);
and U24836 (N_24836,N_19004,N_23875);
nor U24837 (N_24837,N_21974,N_23306);
and U24838 (N_24838,N_18772,N_21816);
nand U24839 (N_24839,N_22921,N_20136);
nand U24840 (N_24840,N_18916,N_22377);
nand U24841 (N_24841,N_23409,N_19841);
nand U24842 (N_24842,N_23330,N_23940);
nor U24843 (N_24843,N_19684,N_21468);
nor U24844 (N_24844,N_20578,N_22828);
nor U24845 (N_24845,N_20566,N_22304);
or U24846 (N_24846,N_23707,N_18457);
nand U24847 (N_24847,N_23012,N_18069);
or U24848 (N_24848,N_19892,N_19239);
and U24849 (N_24849,N_23342,N_22895);
and U24850 (N_24850,N_22362,N_23755);
nor U24851 (N_24851,N_19759,N_22424);
nor U24852 (N_24852,N_18931,N_21251);
or U24853 (N_24853,N_19989,N_22521);
and U24854 (N_24854,N_22023,N_22735);
or U24855 (N_24855,N_18512,N_20597);
nand U24856 (N_24856,N_21516,N_18329);
nor U24857 (N_24857,N_22722,N_19412);
xnor U24858 (N_24858,N_21804,N_22500);
nor U24859 (N_24859,N_23577,N_20854);
and U24860 (N_24860,N_23400,N_19131);
xor U24861 (N_24861,N_22873,N_22659);
nand U24862 (N_24862,N_23456,N_22523);
or U24863 (N_24863,N_22761,N_23275);
nor U24864 (N_24864,N_18233,N_18705);
or U24865 (N_24865,N_18466,N_23246);
nand U24866 (N_24866,N_19945,N_21172);
nand U24867 (N_24867,N_21912,N_19877);
nand U24868 (N_24868,N_20299,N_20383);
nor U24869 (N_24869,N_19717,N_18306);
or U24870 (N_24870,N_18933,N_23187);
and U24871 (N_24871,N_21839,N_23965);
or U24872 (N_24872,N_21482,N_22360);
nor U24873 (N_24873,N_19395,N_23540);
xor U24874 (N_24874,N_20964,N_20394);
or U24875 (N_24875,N_18761,N_18770);
xnor U24876 (N_24876,N_21437,N_23063);
nand U24877 (N_24877,N_20861,N_19571);
xnor U24878 (N_24878,N_21771,N_22479);
and U24879 (N_24879,N_22035,N_18701);
nor U24880 (N_24880,N_20230,N_19660);
nand U24881 (N_24881,N_22303,N_21879);
xor U24882 (N_24882,N_23059,N_19568);
nand U24883 (N_24883,N_19362,N_19967);
nor U24884 (N_24884,N_20503,N_22077);
and U24885 (N_24885,N_19971,N_21623);
nand U24886 (N_24886,N_23154,N_22342);
and U24887 (N_24887,N_21407,N_18739);
xnor U24888 (N_24888,N_18386,N_20419);
and U24889 (N_24889,N_19652,N_23988);
and U24890 (N_24890,N_21990,N_22096);
nand U24891 (N_24891,N_23811,N_22931);
or U24892 (N_24892,N_18677,N_22083);
or U24893 (N_24893,N_20782,N_22274);
nor U24894 (N_24894,N_20915,N_23199);
or U24895 (N_24895,N_21526,N_20021);
or U24896 (N_24896,N_23481,N_19402);
or U24897 (N_24897,N_21100,N_23864);
and U24898 (N_24898,N_18164,N_21888);
and U24899 (N_24899,N_18954,N_18801);
or U24900 (N_24900,N_23019,N_18125);
and U24901 (N_24901,N_23398,N_19847);
nand U24902 (N_24902,N_23771,N_19103);
xnor U24903 (N_24903,N_19307,N_21285);
xnor U24904 (N_24904,N_20162,N_23539);
xnor U24905 (N_24905,N_22226,N_23860);
or U24906 (N_24906,N_19596,N_22501);
nor U24907 (N_24907,N_20905,N_19630);
nand U24908 (N_24908,N_20840,N_23832);
nor U24909 (N_24909,N_19853,N_19081);
nand U24910 (N_24910,N_18455,N_19728);
nand U24911 (N_24911,N_20973,N_21347);
nor U24912 (N_24912,N_21855,N_22231);
or U24913 (N_24913,N_22224,N_21640);
or U24914 (N_24914,N_19102,N_22993);
or U24915 (N_24915,N_22068,N_18209);
xor U24916 (N_24916,N_19905,N_23598);
and U24917 (N_24917,N_22863,N_18379);
and U24918 (N_24918,N_20511,N_19411);
nor U24919 (N_24919,N_19901,N_23014);
and U24920 (N_24920,N_19584,N_23683);
xor U24921 (N_24921,N_23107,N_23384);
and U24922 (N_24922,N_20596,N_22890);
and U24923 (N_24923,N_21143,N_21370);
and U24924 (N_24924,N_21520,N_21252);
nor U24925 (N_24925,N_20209,N_23782);
xnor U24926 (N_24926,N_23753,N_19167);
and U24927 (N_24927,N_18469,N_21277);
nor U24928 (N_24928,N_19519,N_23280);
xor U24929 (N_24929,N_20107,N_23914);
nand U24930 (N_24930,N_20351,N_23815);
nand U24931 (N_24931,N_21517,N_21087);
nor U24932 (N_24932,N_20033,N_23891);
nand U24933 (N_24933,N_21317,N_23311);
nand U24934 (N_24934,N_20526,N_22378);
nor U24935 (N_24935,N_20577,N_20560);
or U24936 (N_24936,N_19082,N_20517);
and U24937 (N_24937,N_18874,N_20037);
nor U24938 (N_24938,N_21206,N_19344);
xnor U24939 (N_24939,N_21492,N_20229);
or U24940 (N_24940,N_21434,N_21638);
and U24941 (N_24941,N_19994,N_20172);
nor U24942 (N_24942,N_23129,N_23561);
and U24943 (N_24943,N_22181,N_23125);
or U24944 (N_24944,N_22674,N_21774);
or U24945 (N_24945,N_18736,N_20079);
or U24946 (N_24946,N_22398,N_22731);
nand U24947 (N_24947,N_18682,N_20284);
or U24948 (N_24948,N_22988,N_21894);
nor U24949 (N_24949,N_22691,N_19215);
or U24950 (N_24950,N_23840,N_19822);
or U24951 (N_24951,N_19035,N_23505);
xor U24952 (N_24952,N_21050,N_20719);
nand U24953 (N_24953,N_18244,N_21264);
nand U24954 (N_24954,N_19956,N_19922);
xor U24955 (N_24955,N_19866,N_21255);
and U24956 (N_24956,N_23944,N_21846);
and U24957 (N_24957,N_21281,N_19334);
and U24958 (N_24958,N_19523,N_21942);
nor U24959 (N_24959,N_22220,N_18378);
nor U24960 (N_24960,N_19725,N_21569);
nand U24961 (N_24961,N_22656,N_20052);
nor U24962 (N_24962,N_23490,N_21204);
and U24963 (N_24963,N_19813,N_20907);
and U24964 (N_24964,N_23255,N_19489);
nor U24965 (N_24965,N_20772,N_20432);
nand U24966 (N_24966,N_19895,N_23387);
and U24967 (N_24967,N_18569,N_18044);
or U24968 (N_24968,N_22316,N_18433);
xor U24969 (N_24969,N_22707,N_18832);
nor U24970 (N_24970,N_22686,N_23614);
or U24971 (N_24971,N_22201,N_19044);
nor U24972 (N_24972,N_22307,N_22945);
xnor U24973 (N_24973,N_23946,N_20382);
nor U24974 (N_24974,N_18902,N_22548);
nor U24975 (N_24975,N_23416,N_19150);
nor U24976 (N_24976,N_23509,N_22411);
and U24977 (N_24977,N_18747,N_23684);
and U24978 (N_24978,N_18259,N_22690);
or U24979 (N_24979,N_23906,N_23696);
nor U24980 (N_24980,N_23788,N_20449);
xnor U24981 (N_24981,N_19405,N_18180);
nor U24982 (N_24982,N_18397,N_19695);
and U24983 (N_24983,N_22601,N_18219);
nor U24984 (N_24984,N_18710,N_22944);
and U24985 (N_24985,N_23673,N_21738);
nand U24986 (N_24986,N_19530,N_23686);
or U24987 (N_24987,N_22959,N_22067);
xor U24988 (N_24988,N_21359,N_23098);
nand U24989 (N_24989,N_19393,N_18291);
nor U24990 (N_24990,N_23792,N_20889);
or U24991 (N_24991,N_18427,N_20490);
and U24992 (N_24992,N_22562,N_21230);
or U24993 (N_24993,N_22688,N_23568);
nand U24994 (N_24994,N_22171,N_18201);
or U24995 (N_24995,N_20384,N_19001);
nand U24996 (N_24996,N_21565,N_18577);
nand U24997 (N_24997,N_21273,N_19893);
nand U24998 (N_24998,N_20966,N_18965);
or U24999 (N_24999,N_19882,N_20087);
or U25000 (N_25000,N_22422,N_22111);
and U25001 (N_25001,N_18534,N_23006);
and U25002 (N_25002,N_21335,N_23024);
nor U25003 (N_25003,N_23000,N_18979);
nor U25004 (N_25004,N_20947,N_18778);
and U25005 (N_25005,N_20909,N_19224);
or U25006 (N_25006,N_20150,N_20649);
nand U25007 (N_25007,N_20157,N_18968);
nor U25008 (N_25008,N_23025,N_22497);
and U25009 (N_25009,N_22667,N_19669);
nand U25010 (N_25010,N_20282,N_22047);
nand U25011 (N_25011,N_23954,N_22195);
or U25012 (N_25012,N_22709,N_20144);
xor U25013 (N_25013,N_20783,N_19761);
nor U25014 (N_25014,N_19419,N_23239);
and U25015 (N_25015,N_18925,N_23776);
nand U25016 (N_25016,N_20430,N_21620);
and U25017 (N_25017,N_23978,N_22259);
nand U25018 (N_25018,N_22232,N_21614);
or U25019 (N_25019,N_22244,N_21376);
nor U25020 (N_25020,N_19337,N_22769);
and U25021 (N_25021,N_20379,N_23132);
xnor U25022 (N_25022,N_23316,N_19632);
nand U25023 (N_25023,N_20457,N_23489);
nand U25024 (N_25024,N_18354,N_22431);
nand U25025 (N_25025,N_20101,N_22346);
or U25026 (N_25026,N_21729,N_22401);
nand U25027 (N_25027,N_20206,N_20644);
nor U25028 (N_25028,N_21373,N_19104);
nor U25029 (N_25029,N_23061,N_18447);
nor U25030 (N_25030,N_22063,N_19754);
xor U25031 (N_25031,N_20561,N_18548);
nor U25032 (N_25032,N_20085,N_21539);
and U25033 (N_25033,N_23023,N_18050);
or U25034 (N_25034,N_22483,N_20631);
nor U25035 (N_25035,N_22032,N_19607);
nand U25036 (N_25036,N_21644,N_19635);
nand U25037 (N_25037,N_20348,N_21628);
nor U25038 (N_25038,N_23920,N_22257);
nand U25039 (N_25039,N_21705,N_19681);
or U25040 (N_25040,N_18910,N_20304);
nor U25041 (N_25041,N_23483,N_23898);
nor U25042 (N_25042,N_19463,N_23355);
nand U25043 (N_25043,N_20881,N_22905);
and U25044 (N_25044,N_23953,N_20266);
or U25045 (N_25045,N_21015,N_19865);
and U25046 (N_25046,N_21240,N_23745);
xor U25047 (N_25047,N_23842,N_22812);
or U25048 (N_25048,N_22366,N_19063);
and U25049 (N_25049,N_19330,N_18038);
or U25050 (N_25050,N_18153,N_23345);
or U25051 (N_25051,N_22582,N_18227);
nor U25052 (N_25052,N_18048,N_22297);
nand U25053 (N_25053,N_20470,N_19978);
nor U25054 (N_25054,N_18628,N_21874);
nor U25055 (N_25055,N_23831,N_22946);
xor U25056 (N_25056,N_22462,N_21221);
xor U25057 (N_25057,N_23530,N_20567);
or U25058 (N_25058,N_23361,N_21261);
and U25059 (N_25059,N_22117,N_22069);
nor U25060 (N_25060,N_20769,N_22822);
nand U25061 (N_25061,N_21177,N_19555);
nor U25062 (N_25062,N_19085,N_23048);
nor U25063 (N_25063,N_21054,N_20298);
and U25064 (N_25064,N_23604,N_19499);
nor U25065 (N_25065,N_22755,N_23942);
or U25066 (N_25066,N_19346,N_20340);
nor U25067 (N_25067,N_21301,N_22518);
nor U25068 (N_25068,N_22903,N_22433);
nor U25069 (N_25069,N_23256,N_20030);
nor U25070 (N_25070,N_20476,N_19015);
nand U25071 (N_25071,N_22104,N_22184);
nor U25072 (N_25072,N_22048,N_22496);
nand U25073 (N_25073,N_19494,N_23660);
nand U25074 (N_25074,N_20068,N_23272);
and U25075 (N_25075,N_22288,N_23629);
nand U25076 (N_25076,N_18713,N_18668);
and U25077 (N_25077,N_21444,N_21126);
nor U25078 (N_25078,N_18396,N_20542);
or U25079 (N_25079,N_20003,N_18454);
and U25080 (N_25080,N_23738,N_21515);
nand U25081 (N_25081,N_21913,N_20751);
or U25082 (N_25082,N_21770,N_18399);
or U25083 (N_25083,N_22110,N_23801);
or U25084 (N_25084,N_18490,N_20933);
or U25085 (N_25085,N_20557,N_19491);
and U25086 (N_25086,N_23586,N_21299);
or U25087 (N_25087,N_23143,N_22663);
xor U25088 (N_25088,N_18547,N_19973);
nand U25089 (N_25089,N_20167,N_21866);
xor U25090 (N_25090,N_20662,N_21728);
nor U25091 (N_25091,N_21744,N_20634);
and U25092 (N_25092,N_18884,N_21228);
nor U25093 (N_25093,N_22347,N_18998);
nor U25094 (N_25094,N_20334,N_18780);
xor U25095 (N_25095,N_18468,N_19373);
nor U25096 (N_25096,N_22229,N_18195);
nand U25097 (N_25097,N_22754,N_21891);
or U25098 (N_25098,N_23248,N_20314);
and U25099 (N_25099,N_23727,N_20192);
nor U25100 (N_25100,N_18813,N_22045);
or U25101 (N_25101,N_22260,N_19106);
and U25102 (N_25102,N_20461,N_22264);
and U25103 (N_25103,N_21438,N_20925);
or U25104 (N_25104,N_20126,N_19885);
nand U25105 (N_25105,N_21248,N_21127);
or U25106 (N_25106,N_18893,N_19161);
or U25107 (N_25107,N_22124,N_22357);
and U25108 (N_25108,N_21762,N_22914);
and U25109 (N_25109,N_20195,N_20388);
nand U25110 (N_25110,N_20024,N_20273);
and U25111 (N_25111,N_23001,N_20994);
nor U25112 (N_25112,N_19554,N_20056);
nor U25113 (N_25113,N_19748,N_21174);
nor U25114 (N_25114,N_19577,N_22400);
and U25115 (N_25115,N_19668,N_23866);
nand U25116 (N_25116,N_21027,N_18418);
and U25117 (N_25117,N_19906,N_23994);
or U25118 (N_25118,N_22856,N_19240);
or U25119 (N_25119,N_22547,N_19216);
nor U25120 (N_25120,N_23297,N_22792);
and U25121 (N_25121,N_23517,N_19525);
or U25122 (N_25122,N_20398,N_22718);
and U25123 (N_25123,N_21103,N_20921);
xnor U25124 (N_25124,N_23981,N_22997);
nand U25125 (N_25125,N_19774,N_23719);
or U25126 (N_25126,N_20699,N_22949);
nand U25127 (N_25127,N_20289,N_19640);
nand U25128 (N_25128,N_20360,N_20396);
nor U25129 (N_25129,N_21354,N_20743);
and U25130 (N_25130,N_18634,N_23135);
nand U25131 (N_25131,N_21125,N_21972);
nor U25132 (N_25132,N_18373,N_21119);
nand U25133 (N_25133,N_20500,N_21202);
and U25134 (N_25134,N_21481,N_21840);
nor U25135 (N_25135,N_23747,N_22834);
and U25136 (N_25136,N_22846,N_22573);
nor U25137 (N_25137,N_19776,N_20032);
nand U25138 (N_25138,N_19384,N_18143);
nand U25139 (N_25139,N_22880,N_18342);
or U25140 (N_25140,N_18026,N_21902);
nand U25141 (N_25141,N_20099,N_18620);
nand U25142 (N_25142,N_22821,N_21549);
or U25143 (N_25143,N_22174,N_21300);
nor U25144 (N_25144,N_19178,N_18934);
or U25145 (N_25145,N_18337,N_20202);
nor U25146 (N_25146,N_21669,N_18017);
xor U25147 (N_25147,N_18294,N_20146);
and U25148 (N_25148,N_18861,N_20293);
and U25149 (N_25149,N_20211,N_20076);
nand U25150 (N_25150,N_23927,N_18479);
and U25151 (N_25151,N_20555,N_19272);
nor U25152 (N_25152,N_21848,N_21915);
nor U25153 (N_25153,N_22368,N_23654);
nor U25154 (N_25154,N_21898,N_18317);
or U25155 (N_25155,N_22710,N_18763);
nand U25156 (N_25156,N_20917,N_21105);
nand U25157 (N_25157,N_20272,N_21356);
nor U25158 (N_25158,N_22549,N_20530);
or U25159 (N_25159,N_22397,N_21432);
nand U25160 (N_25160,N_19448,N_22716);
nand U25161 (N_25161,N_20728,N_18798);
or U25162 (N_25162,N_21779,N_21763);
or U25163 (N_25163,N_23413,N_21372);
or U25164 (N_25164,N_22221,N_20152);
nand U25165 (N_25165,N_22404,N_22833);
and U25166 (N_25166,N_21327,N_20827);
nor U25167 (N_25167,N_20632,N_22859);
and U25168 (N_25168,N_20196,N_20064);
nand U25169 (N_25169,N_21022,N_23997);
and U25170 (N_25170,N_23910,N_20036);
nand U25171 (N_25171,N_18923,N_22618);
nand U25172 (N_25172,N_19604,N_20402);
or U25173 (N_25173,N_18865,N_22086);
and U25174 (N_25174,N_20945,N_19805);
xnor U25175 (N_25175,N_22994,N_18271);
and U25176 (N_25176,N_20151,N_18901);
nand U25177 (N_25177,N_21597,N_21575);
and U25178 (N_25178,N_20115,N_20520);
and U25179 (N_25179,N_23096,N_18760);
or U25180 (N_25180,N_23596,N_18088);
nand U25181 (N_25181,N_19368,N_23030);
nor U25182 (N_25182,N_19507,N_18184);
or U25183 (N_25183,N_21425,N_20640);
nand U25184 (N_25184,N_22494,N_19651);
or U25185 (N_25185,N_23515,N_18971);
nand U25186 (N_25186,N_22420,N_18639);
nand U25187 (N_25187,N_19560,N_19066);
or U25188 (N_25188,N_19222,N_23902);
or U25189 (N_25189,N_23148,N_19935);
or U25190 (N_25190,N_20949,N_20443);
nand U25191 (N_25191,N_19232,N_22736);
nor U25192 (N_25192,N_21439,N_18644);
and U25193 (N_25193,N_22214,N_20234);
or U25194 (N_25194,N_21593,N_20426);
and U25195 (N_25195,N_19959,N_20341);
nor U25196 (N_25196,N_20042,N_21162);
nand U25197 (N_25197,N_19289,N_23039);
and U25198 (N_25198,N_21497,N_18471);
nor U25199 (N_25199,N_23056,N_18732);
nor U25200 (N_25200,N_21504,N_19151);
nor U25201 (N_25201,N_19014,N_19960);
or U25202 (N_25202,N_22447,N_21329);
nand U25203 (N_25203,N_23887,N_23160);
and U25204 (N_25204,N_22040,N_23949);
or U25205 (N_25205,N_18953,N_20350);
nand U25206 (N_25206,N_19506,N_23222);
and U25207 (N_25207,N_18651,N_22365);
or U25208 (N_25208,N_21472,N_20862);
nand U25209 (N_25209,N_21820,N_20240);
or U25210 (N_25210,N_19817,N_18787);
and U25211 (N_25211,N_21814,N_21747);
and U25212 (N_25212,N_20753,N_22738);
xnor U25213 (N_25213,N_23198,N_22807);
nand U25214 (N_25214,N_19803,N_22416);
nor U25215 (N_25215,N_19034,N_21616);
nand U25216 (N_25216,N_20951,N_20002);
nor U25217 (N_25217,N_21949,N_22703);
nor U25218 (N_25218,N_22967,N_21431);
xnor U25219 (N_25219,N_22794,N_20460);
nand U25220 (N_25220,N_23352,N_23549);
nor U25221 (N_25221,N_23619,N_19155);
nor U25222 (N_25222,N_21326,N_22429);
or U25223 (N_25223,N_23638,N_20865);
or U25224 (N_25224,N_23418,N_23880);
xor U25225 (N_25225,N_21424,N_23146);
nor U25226 (N_25226,N_23395,N_23584);
xnor U25227 (N_25227,N_18232,N_22737);
nand U25228 (N_25228,N_20378,N_20513);
or U25229 (N_25229,N_18331,N_19408);
and U25230 (N_25230,N_19768,N_20536);
nand U25231 (N_25231,N_22405,N_23648);
or U25232 (N_25232,N_21419,N_19376);
nand U25233 (N_25233,N_19111,N_19188);
nor U25234 (N_25234,N_18324,N_22733);
nor U25235 (N_25235,N_23590,N_18940);
nand U25236 (N_25236,N_23796,N_19875);
nor U25237 (N_25237,N_21769,N_20791);
nand U25238 (N_25238,N_18037,N_20483);
or U25239 (N_25239,N_21402,N_23661);
nand U25240 (N_25240,N_23912,N_20992);
nor U25241 (N_25241,N_20139,N_19431);
xor U25242 (N_25242,N_21822,N_18588);
nand U25243 (N_25243,N_23258,N_20684);
nand U25244 (N_25244,N_23961,N_18408);
nand U25245 (N_25245,N_21164,N_19835);
or U25246 (N_25246,N_22289,N_20216);
and U25247 (N_25247,N_19409,N_19746);
or U25248 (N_25248,N_20278,N_23094);
or U25249 (N_25249,N_19177,N_23675);
nor U25250 (N_25250,N_21060,N_22478);
nor U25251 (N_25251,N_23585,N_23114);
and U25252 (N_25252,N_21670,N_18969);
nor U25253 (N_25253,N_22612,N_23034);
nand U25254 (N_25254,N_20013,N_21219);
xnor U25255 (N_25255,N_18146,N_19493);
xnor U25256 (N_25256,N_22161,N_23120);
nor U25257 (N_25257,N_23534,N_18543);
nand U25258 (N_25258,N_22625,N_21688);
nand U25259 (N_25259,N_23659,N_21063);
nand U25260 (N_25260,N_21687,N_18283);
and U25261 (N_25261,N_21802,N_23121);
nor U25262 (N_25262,N_22617,N_22904);
nor U25263 (N_25263,N_18742,N_19671);
or U25264 (N_25264,N_18952,N_20943);
xnor U25265 (N_25265,N_18709,N_18906);
nor U25266 (N_25266,N_20784,N_23959);
or U25267 (N_25267,N_23923,N_23465);
or U25268 (N_25268,N_22154,N_20411);
nor U25269 (N_25269,N_22272,N_19732);
and U25270 (N_25270,N_22520,N_21178);
and U25271 (N_25271,N_22868,N_18693);
nand U25272 (N_25272,N_20710,N_18823);
nand U25273 (N_25273,N_23070,N_18110);
nor U25274 (N_25274,N_21295,N_22095);
nor U25275 (N_25275,N_20109,N_18335);
nor U25276 (N_25276,N_20016,N_19924);
nor U25277 (N_25277,N_21323,N_20065);
xor U25278 (N_25278,N_18997,N_21039);
and U25279 (N_25279,N_18810,N_20495);
and U25280 (N_25280,N_21783,N_20789);
nor U25281 (N_25281,N_20025,N_18014);
nor U25282 (N_25282,N_20454,N_18554);
nor U25283 (N_25283,N_20629,N_23078);
nor U25284 (N_25284,N_22881,N_23503);
nor U25285 (N_25285,N_20770,N_20354);
or U25286 (N_25286,N_21038,N_18800);
nand U25287 (N_25287,N_18364,N_20856);
nor U25288 (N_25288,N_19755,N_18055);
or U25289 (N_25289,N_23037,N_22685);
nand U25290 (N_25290,N_23075,N_22875);
and U25291 (N_25291,N_18312,N_23704);
and U25292 (N_25292,N_22100,N_23723);
nor U25293 (N_25293,N_23926,N_20847);
xor U25294 (N_25294,N_18598,N_19076);
and U25295 (N_25295,N_18041,N_19160);
nor U25296 (N_25296,N_18877,N_19793);
xnor U25297 (N_25297,N_21094,N_20609);
nor U25298 (N_25298,N_21239,N_20043);
xnor U25299 (N_25299,N_21290,N_19212);
or U25300 (N_25300,N_20911,N_20730);
nor U25301 (N_25301,N_23106,N_19857);
nor U25302 (N_25302,N_23544,N_21901);
nand U25303 (N_25303,N_22423,N_19868);
nand U25304 (N_25304,N_23740,N_19047);
nand U25305 (N_25305,N_21722,N_22043);
nand U25306 (N_25306,N_23370,N_23839);
nor U25307 (N_25307,N_19936,N_23605);
nand U25308 (N_25308,N_18305,N_21461);
nor U25309 (N_25309,N_21364,N_19074);
or U25310 (N_25310,N_20685,N_23464);
or U25311 (N_25311,N_22348,N_18629);
or U25312 (N_25312,N_19864,N_22775);
or U25313 (N_25313,N_23834,N_19294);
or U25314 (N_25314,N_23460,N_21914);
nand U25315 (N_25315,N_18057,N_21580);
and U25316 (N_25316,N_21973,N_20201);
nor U25317 (N_25317,N_18056,N_19731);
nand U25318 (N_25318,N_18892,N_21518);
nor U25319 (N_25319,N_19899,N_19628);
and U25320 (N_25320,N_21395,N_18564);
or U25321 (N_25321,N_19118,N_21541);
and U25322 (N_25322,N_19939,N_20809);
nor U25323 (N_25323,N_20047,N_19287);
and U25324 (N_25324,N_21946,N_22197);
or U25325 (N_25325,N_21545,N_19002);
or U25326 (N_25326,N_22252,N_22062);
xor U25327 (N_25327,N_23963,N_23005);
xnor U25328 (N_25328,N_20527,N_23445);
xor U25329 (N_25329,N_21546,N_23185);
xnor U25330 (N_25330,N_22230,N_22534);
and U25331 (N_25331,N_23245,N_20027);
and U25332 (N_25332,N_22705,N_20724);
nand U25333 (N_25333,N_23535,N_21921);
and U25334 (N_25334,N_21574,N_21279);
or U25335 (N_25335,N_22460,N_19228);
nand U25336 (N_25336,N_23032,N_20228);
or U25337 (N_25337,N_18964,N_19055);
nor U25338 (N_25338,N_19199,N_22789);
and U25339 (N_25339,N_22344,N_18671);
nor U25340 (N_25340,N_21944,N_18112);
nand U25341 (N_25341,N_18353,N_22415);
xor U25342 (N_25342,N_18434,N_19812);
or U25343 (N_25343,N_22925,N_20748);
nand U25344 (N_25344,N_20983,N_23470);
nand U25345 (N_25345,N_20154,N_21662);
and U25346 (N_25346,N_21587,N_21034);
and U25347 (N_25347,N_18516,N_22810);
nor U25348 (N_25348,N_23084,N_19718);
xor U25349 (N_25349,N_20375,N_19238);
nand U25350 (N_25350,N_20161,N_23328);
and U25351 (N_25351,N_21694,N_20942);
nor U25352 (N_25352,N_22643,N_23725);
and U25353 (N_25353,N_18599,N_19870);
and U25354 (N_25354,N_18352,N_18133);
or U25355 (N_25355,N_19814,N_18404);
nor U25356 (N_25356,N_19233,N_23767);
nor U25357 (N_25357,N_19686,N_22882);
nand U25358 (N_25358,N_18643,N_22317);
or U25359 (N_25359,N_20358,N_18771);
nor U25360 (N_25360,N_21146,N_22844);
nor U25361 (N_25361,N_21488,N_18504);
or U25362 (N_25362,N_22970,N_18156);
nor U25363 (N_25363,N_22795,N_18441);
and U25364 (N_25364,N_21123,N_20521);
or U25365 (N_25365,N_22319,N_22421);
nand U25366 (N_25366,N_21683,N_21483);
or U25367 (N_25367,N_22222,N_19986);
or U25368 (N_25368,N_21895,N_23408);
nor U25369 (N_25369,N_22670,N_19473);
xor U25370 (N_25370,N_21033,N_21084);
xnor U25371 (N_25371,N_23069,N_23728);
nor U25372 (N_25372,N_22352,N_23600);
or U25373 (N_25373,N_19744,N_18983);
or U25374 (N_25374,N_22109,N_18121);
and U25375 (N_25375,N_18171,N_18129);
nor U25376 (N_25376,N_21436,N_19391);
or U25377 (N_25377,N_19255,N_19775);
nand U25378 (N_25378,N_18722,N_22373);
nor U25379 (N_25379,N_21768,N_23825);
and U25380 (N_25380,N_23343,N_21777);
and U25381 (N_25381,N_22528,N_23376);
and U25382 (N_25382,N_20738,N_19136);
and U25383 (N_25383,N_18854,N_19129);
xnor U25384 (N_25384,N_18377,N_22441);
nor U25385 (N_25385,N_22269,N_18766);
nor U25386 (N_25386,N_20814,N_23921);
or U25387 (N_25387,N_19919,N_19148);
and U25388 (N_25388,N_22702,N_22791);
and U25389 (N_25389,N_19009,N_23830);
and U25390 (N_25390,N_21336,N_18027);
and U25391 (N_25391,N_18762,N_20811);
nand U25392 (N_25392,N_22058,N_20931);
nand U25393 (N_25393,N_20549,N_20325);
nor U25394 (N_25394,N_20932,N_22968);
xor U25395 (N_25395,N_18175,N_18370);
xor U25396 (N_25396,N_20125,N_19429);
xnor U25397 (N_25397,N_22010,N_23366);
and U25398 (N_25398,N_22266,N_22172);
or U25399 (N_25399,N_19423,N_22432);
nor U25400 (N_25400,N_20477,N_19459);
or U25401 (N_25401,N_19663,N_18409);
nand U25402 (N_25402,N_20884,N_18042);
nand U25403 (N_25403,N_18864,N_20913);
and U25404 (N_25404,N_23203,N_19675);
or U25405 (N_25405,N_18581,N_21017);
and U25406 (N_25406,N_21954,N_22569);
nand U25407 (N_25407,N_22538,N_22541);
and U25408 (N_25408,N_23091,N_23781);
nand U25409 (N_25409,N_22786,N_18456);
and U25410 (N_25410,N_20137,N_21018);
and U25411 (N_25411,N_23443,N_20793);
or U25412 (N_25412,N_21314,N_20581);
nor U25413 (N_25413,N_20007,N_21522);
or U25414 (N_25414,N_20486,N_20773);
or U25415 (N_25415,N_21988,N_19425);
nand U25416 (N_25416,N_19230,N_20614);
nor U25417 (N_25417,N_21321,N_20902);
nand U25418 (N_25418,N_20336,N_18642);
nand U25419 (N_25419,N_21598,N_21002);
xnor U25420 (N_25420,N_23833,N_18149);
xnor U25421 (N_25421,N_23497,N_23027);
xor U25422 (N_25422,N_19252,N_19471);
or U25423 (N_25423,N_19451,N_18724);
xnor U25424 (N_25424,N_18619,N_22082);
nand U25425 (N_25425,N_21612,N_19827);
nand U25426 (N_25426,N_18570,N_23574);
and U25427 (N_25427,N_22241,N_19352);
or U25428 (N_25428,N_20528,N_19297);
nand U25429 (N_25429,N_19481,N_18183);
nor U25430 (N_25430,N_20132,N_23029);
nor U25431 (N_25431,N_19625,N_23147);
xnor U25432 (N_25432,N_19900,N_20929);
or U25433 (N_25433,N_22375,N_22061);
nand U25434 (N_25434,N_18507,N_22450);
or U25435 (N_25435,N_19548,N_19185);
nand U25436 (N_25436,N_20084,N_21397);
nor U25437 (N_25437,N_20028,N_20757);
nor U25438 (N_25438,N_19038,N_23016);
nor U25439 (N_25439,N_20119,N_19027);
nand U25440 (N_25440,N_19403,N_23849);
nand U25441 (N_25441,N_20212,N_19594);
nor U25442 (N_25442,N_21743,N_22322);
or U25443 (N_25443,N_23819,N_18016);
or U25444 (N_25444,N_23636,N_18895);
or U25445 (N_25445,N_23709,N_18859);
nor U25446 (N_25446,N_23156,N_20090);
or U25447 (N_25447,N_19171,N_22235);
nand U25448 (N_25448,N_19848,N_19751);
xor U25449 (N_25449,N_19856,N_21223);
and U25450 (N_25450,N_20637,N_22007);
or U25451 (N_25451,N_23193,N_21179);
xor U25452 (N_25452,N_18667,N_21467);
nand U25453 (N_25453,N_21736,N_19268);
nand U25454 (N_25454,N_23439,N_21621);
nor U25455 (N_25455,N_22193,N_22721);
or U25456 (N_25456,N_23184,N_21310);
and U25457 (N_25457,N_18505,N_23710);
nor U25458 (N_25458,N_22492,N_19156);
and U25459 (N_25459,N_22418,N_20446);
nand U25460 (N_25460,N_18075,N_19444);
and U25461 (N_25461,N_18136,N_22800);
and U25462 (N_25462,N_19950,N_19862);
nand U25463 (N_25463,N_21543,N_19879);
or U25464 (N_25464,N_18302,N_20034);
nand U25465 (N_25465,N_20588,N_19343);
nand U25466 (N_25466,N_20975,N_22320);
nor U25467 (N_25467,N_23332,N_19166);
and U25468 (N_25468,N_22850,N_23786);
nand U25469 (N_25469,N_20653,N_20774);
nand U25470 (N_25470,N_22639,N_23769);
nand U25471 (N_25471,N_22784,N_19716);
nor U25472 (N_25472,N_23457,N_23536);
nand U25473 (N_25473,N_20318,N_22285);
or U25474 (N_25474,N_20794,N_23627);
nand U25475 (N_25475,N_23804,N_20000);
nand U25476 (N_25476,N_18608,N_21086);
or U25477 (N_25477,N_20220,N_21506);
and U25478 (N_25478,N_20406,N_23744);
nor U25479 (N_25479,N_19846,N_19487);
or U25480 (N_25480,N_21447,N_20543);
nand U25481 (N_25481,N_18135,N_21218);
and U25482 (N_25482,N_20665,N_22723);
or U25483 (N_25483,N_23916,N_22902);
nand U25484 (N_25484,N_22490,N_21333);
nor U25485 (N_25485,N_20619,N_23212);
nor U25486 (N_25486,N_19141,N_21810);
and U25487 (N_25487,N_22115,N_23102);
nor U25488 (N_25488,N_19586,N_21714);
and U25489 (N_25489,N_23440,N_18185);
nor U25490 (N_25490,N_18822,N_22278);
or U25491 (N_25491,N_23947,N_21235);
and U25492 (N_25492,N_19132,N_19823);
nand U25493 (N_25493,N_22560,N_19674);
nor U25494 (N_25494,N_23179,N_19279);
or U25495 (N_25495,N_20974,N_23449);
nand U25496 (N_25496,N_23004,N_18625);
or U25497 (N_25497,N_23188,N_19096);
and U25498 (N_25498,N_22644,N_22926);
and U25499 (N_25499,N_18119,N_18086);
nand U25500 (N_25500,N_21685,N_23646);
or U25501 (N_25501,N_23485,N_21210);
or U25502 (N_25502,N_19005,N_20648);
nand U25503 (N_25503,N_19387,N_18429);
nand U25504 (N_25504,N_22240,N_18287);
nand U25505 (N_25505,N_18486,N_21452);
and U25506 (N_25506,N_22393,N_20178);
nand U25507 (N_25507,N_20936,N_23007);
or U25508 (N_25508,N_20664,N_20797);
nor U25509 (N_25509,N_23777,N_23349);
or U25510 (N_25510,N_20447,N_20366);
nand U25511 (N_25511,N_19539,N_18290);
and U25512 (N_25512,N_22790,N_20381);
nor U25513 (N_25513,N_22566,N_19570);
nor U25514 (N_25514,N_20401,N_23473);
and U25515 (N_25515,N_22603,N_19154);
or U25516 (N_25516,N_23433,N_23528);
nor U25517 (N_25517,N_19777,N_18727);
or U25518 (N_25518,N_23892,N_18579);
and U25519 (N_25519,N_20365,N_23371);
nor U25520 (N_25520,N_18365,N_20142);
nor U25521 (N_25521,N_19124,N_23119);
or U25522 (N_25522,N_21061,N_18729);
nor U25523 (N_25523,N_21739,N_20110);
or U25524 (N_25524,N_23093,N_20117);
nor U25525 (N_25525,N_20716,N_19609);
nor U25526 (N_25526,N_20029,N_18087);
or U25527 (N_25527,N_20128,N_20245);
or U25528 (N_25528,N_19698,N_19923);
xnor U25529 (N_25529,N_19053,N_19873);
nand U25530 (N_25530,N_18764,N_21184);
nor U25531 (N_25531,N_21242,N_20878);
or U25532 (N_25532,N_19563,N_23741);
nor U25533 (N_25533,N_22064,N_19108);
or U25534 (N_25534,N_22129,N_23104);
nand U25535 (N_25535,N_18246,N_22646);
or U25536 (N_25536,N_19374,N_19126);
or U25537 (N_25537,N_22299,N_22408);
or U25538 (N_25538,N_18254,N_18172);
nor U25539 (N_25539,N_20235,N_19979);
xor U25540 (N_25540,N_22203,N_18372);
nor U25541 (N_25541,N_22438,N_23382);
and U25542 (N_25542,N_21850,N_20097);
and U25543 (N_25543,N_19722,N_23452);
or U25544 (N_25544,N_19054,N_23650);
and U25545 (N_25545,N_19955,N_20867);
nor U25546 (N_25546,N_19582,N_18792);
or U25547 (N_25547,N_21099,N_18618);
nor U25548 (N_25548,N_19265,N_18556);
and U25549 (N_25549,N_20140,N_20094);
or U25550 (N_25550,N_20659,N_21361);
and U25551 (N_25551,N_20868,N_23592);
nor U25552 (N_25552,N_19839,N_18202);
nand U25553 (N_25553,N_18809,N_20166);
and U25554 (N_25554,N_20231,N_23151);
nand U25555 (N_25555,N_20562,N_18829);
nand U25556 (N_25556,N_22517,N_19281);
nor U25557 (N_25557,N_20428,N_19602);
xnor U25558 (N_25558,N_22446,N_23701);
nand U25559 (N_25559,N_20331,N_21430);
or U25560 (N_25560,N_18200,N_19040);
and U25561 (N_25561,N_21069,N_23064);
nor U25562 (N_25562,N_19310,N_19315);
and U25563 (N_25563,N_21919,N_21311);
nor U25564 (N_25564,N_20296,N_18817);
or U25565 (N_25565,N_22175,N_20704);
or U25566 (N_25566,N_23052,N_22165);
or U25567 (N_25567,N_19536,N_21348);
nand U25568 (N_25568,N_20063,N_20993);
xor U25569 (N_25569,N_19799,N_19562);
nor U25570 (N_25570,N_20673,N_21507);
nor U25571 (N_25571,N_18659,N_23672);
or U25572 (N_25572,N_18723,N_20816);
xor U25573 (N_25573,N_21751,N_22312);
nor U25574 (N_25574,N_21925,N_23575);
or U25575 (N_25575,N_22782,N_18126);
and U25576 (N_25576,N_21887,N_22751);
nand U25577 (N_25577,N_20392,N_20747);
and U25578 (N_25578,N_23929,N_19730);
nand U25579 (N_25579,N_18452,N_20627);
nand U25580 (N_25580,N_21392,N_21141);
nor U25581 (N_25581,N_18993,N_18058);
nor U25582 (N_25582,N_22675,N_18593);
nand U25583 (N_25583,N_22609,N_20374);
nor U25584 (N_25584,N_21923,N_22869);
and U25585 (N_25585,N_23732,N_22938);
or U25586 (N_25586,N_18930,N_18960);
nand U25587 (N_25587,N_20939,N_18827);
or U25588 (N_25588,N_22942,N_19056);
or U25589 (N_25589,N_19860,N_18292);
nor U25590 (N_25590,N_21537,N_21029);
nor U25591 (N_25591,N_21056,N_21450);
and U25592 (N_25592,N_22367,N_20213);
or U25593 (N_25593,N_23303,N_19829);
or U25594 (N_25594,N_20960,N_21529);
nor U25595 (N_25595,N_23045,N_18676);
and U25596 (N_25596,N_21967,N_18385);
and U25597 (N_25597,N_21344,N_19826);
and U25598 (N_25598,N_21098,N_19206);
and U25599 (N_25599,N_19517,N_18680);
nand U25600 (N_25600,N_23551,N_23889);
and U25601 (N_25601,N_18740,N_22556);
nor U25602 (N_25602,N_20941,N_19336);
xor U25603 (N_25603,N_22939,N_18344);
nand U25604 (N_25604,N_21996,N_19328);
xor U25605 (N_25605,N_22631,N_20124);
nor U25606 (N_25606,N_23397,N_20977);
nand U25607 (N_25607,N_21349,N_21208);
or U25608 (N_25608,N_20238,N_22940);
and U25609 (N_25609,N_21964,N_20579);
nand U25610 (N_25610,N_22741,N_19624);
nand U25611 (N_25611,N_21382,N_23925);
or U25612 (N_25612,N_21051,N_19365);
or U25613 (N_25613,N_18211,N_18881);
nor U25614 (N_25614,N_20736,N_21624);
nand U25615 (N_25615,N_21842,N_19642);
and U25616 (N_25616,N_18743,N_21645);
nor U25617 (N_25617,N_21188,N_18194);
and U25618 (N_25618,N_18944,N_19527);
or U25619 (N_25619,N_18638,N_23770);
nand U25620 (N_25620,N_21890,N_18806);
nand U25621 (N_25621,N_21637,N_19176);
nand U25622 (N_25622,N_23697,N_22660);
and U25623 (N_25623,N_20564,N_19883);
nor U25624 (N_25624,N_22958,N_19546);
and U25625 (N_25625,N_18804,N_23087);
or U25626 (N_25626,N_19974,N_19612);
and U25627 (N_25627,N_23867,N_23360);
nand U25628 (N_25628,N_20551,N_20697);
nand U25629 (N_25629,N_22374,N_23899);
nor U25630 (N_25630,N_19521,N_20498);
xnor U25631 (N_25631,N_22199,N_20327);
or U25632 (N_25632,N_18970,N_21513);
nor U25633 (N_25633,N_19201,N_18346);
nor U25634 (N_25634,N_20616,N_22760);
nor U25635 (N_25635,N_20226,N_21561);
or U25636 (N_25636,N_23808,N_22475);
nor U25637 (N_25637,N_22708,N_21980);
and U25638 (N_25638,N_22632,N_22852);
and U25639 (N_25639,N_19302,N_19318);
or U25640 (N_25640,N_18797,N_22329);
xnor U25641 (N_25641,N_22156,N_23794);
nor U25642 (N_25642,N_19533,N_20965);
and U25643 (N_25643,N_19673,N_21843);
or U25644 (N_25644,N_18239,N_20189);
nor U25645 (N_25645,N_20435,N_19704);
nor U25646 (N_25646,N_18340,N_18021);
or U25647 (N_25647,N_20264,N_21440);
nor U25648 (N_25648,N_19301,N_22985);
nor U25649 (N_25649,N_19734,N_21293);
nor U25650 (N_25650,N_21877,N_22079);
nor U25651 (N_25651,N_20766,N_21905);
and U25652 (N_25652,N_20529,N_21629);
nand U25653 (N_25653,N_20346,N_23877);
and U25654 (N_25654,N_22633,N_22747);
or U25655 (N_25655,N_19790,N_20062);
xnor U25656 (N_25656,N_21723,N_19246);
nor U25657 (N_25657,N_18411,N_19020);
nor U25658 (N_25658,N_18391,N_20307);
nand U25659 (N_25659,N_19589,N_23570);
nor U25660 (N_25660,N_18999,N_23945);
nor U25661 (N_25661,N_19043,N_18885);
xnor U25662 (N_25662,N_19296,N_18539);
nor U25663 (N_25663,N_19943,N_19898);
nor U25664 (N_25664,N_19071,N_19729);
xor U25665 (N_25665,N_18100,N_21761);
nand U25666 (N_25666,N_21957,N_22920);
and U25667 (N_25667,N_21350,N_19175);
nor U25668 (N_25668,N_23183,N_20494);
nand U25669 (N_25669,N_18756,N_22503);
nor U25670 (N_25670,N_19998,N_20174);
or U25671 (N_25671,N_18775,N_21262);
or U25672 (N_25672,N_19204,N_18879);
or U25673 (N_25673,N_18883,N_19165);
nand U25674 (N_25674,N_23532,N_20074);
or U25675 (N_25675,N_21365,N_20208);
nor U25676 (N_25676,N_21867,N_18032);
nand U25677 (N_25677,N_18094,N_19785);
and U25678 (N_25678,N_23463,N_22219);
or U25679 (N_25679,N_18336,N_23136);
and U25680 (N_25680,N_21604,N_18867);
or U25681 (N_25681,N_20478,N_18571);
and U25682 (N_25682,N_20689,N_22636);
and U25683 (N_25683,N_21120,N_19468);
and U25684 (N_25684,N_19742,N_19342);
or U25685 (N_25685,N_19000,N_18863);
nor U25686 (N_25686,N_19984,N_22098);
or U25687 (N_25687,N_21041,N_22635);
xnor U25688 (N_25688,N_20073,N_23905);
nand U25689 (N_25689,N_20507,N_22242);
nor U25690 (N_25690,N_21552,N_22814);
or U25691 (N_25691,N_18141,N_22194);
and U25692 (N_25692,N_23191,N_18689);
xor U25693 (N_25693,N_20177,N_19196);
nand U25694 (N_25694,N_19277,N_21953);
nand U25695 (N_25695,N_20259,N_19819);
and U25696 (N_25696,N_22205,N_20740);
nor U25697 (N_25697,N_19643,N_18675);
nand U25698 (N_25698,N_22544,N_23890);
nand U25699 (N_25699,N_18101,N_18444);
nand U25700 (N_25700,N_20553,N_21362);
and U25701 (N_25701,N_18280,N_21149);
nor U25702 (N_25702,N_22363,N_18193);
or U25703 (N_25703,N_21681,N_20475);
and U25704 (N_25704,N_23215,N_20496);
or U25705 (N_25705,N_20438,N_22176);
and U25706 (N_25706,N_23543,N_21287);
nor U25707 (N_25707,N_23624,N_23207);
or U25708 (N_25708,N_18008,N_21137);
or U25709 (N_25709,N_19338,N_21077);
nand U25710 (N_25710,N_22896,N_19977);
or U25711 (N_25711,N_19721,N_18501);
nor U25712 (N_25712,N_18467,N_21536);
nor U25713 (N_25713,N_18341,N_22127);
nand U25714 (N_25714,N_22915,N_19760);
xnor U25715 (N_25715,N_22897,N_22463);
and U25716 (N_25716,N_21477,N_19026);
nand U25717 (N_25717,N_19369,N_20050);
or U25718 (N_25718,N_22293,N_19645);
and U25719 (N_25719,N_22465,N_19340);
and U25720 (N_25720,N_21854,N_20487);
or U25721 (N_25721,N_19672,N_22793);
or U25722 (N_25722,N_18662,N_18252);
or U25723 (N_25723,N_20919,N_20812);
and U25724 (N_25724,N_23897,N_19553);
nor U25725 (N_25725,N_23112,N_23313);
nand U25726 (N_25726,N_18077,N_23231);
nor U25727 (N_25727,N_21375,N_18439);
or U25728 (N_25728,N_20397,N_20469);
nor U25729 (N_25729,N_22819,N_21042);
or U25730 (N_25730,N_20750,N_21590);
nand U25731 (N_25731,N_23326,N_23726);
and U25732 (N_25732,N_20286,N_21947);
nor U25733 (N_25733,N_19492,N_22907);
or U25734 (N_25734,N_19070,N_20368);
or U25735 (N_25735,N_20241,N_20376);
nand U25736 (N_25736,N_20709,N_18398);
nor U25737 (N_25737,N_20611,N_23462);
or U25738 (N_25738,N_19303,N_23318);
nor U25739 (N_25739,N_19581,N_23294);
nand U25740 (N_25740,N_19836,N_18942);
or U25741 (N_25741,N_20300,N_22813);
and U25742 (N_25742,N_20546,N_23394);
xor U25743 (N_25743,N_19243,N_20427);
or U25744 (N_25744,N_23611,N_20540);
xor U25745 (N_25745,N_21357,N_18612);
and U25746 (N_25746,N_18113,N_22923);
nand U25747 (N_25747,N_18683,N_20835);
and U25748 (N_25748,N_23904,N_19149);
or U25749 (N_25749,N_20787,N_22916);
and U25750 (N_25750,N_19678,N_22054);
and U25751 (N_25751,N_20509,N_22854);
or U25752 (N_25752,N_21247,N_21046);
or U25753 (N_25753,N_18765,N_18886);
nor U25754 (N_25754,N_20828,N_18746);
nor U25755 (N_25755,N_18431,N_19025);
nand U25756 (N_25756,N_18748,N_19214);
nand U25757 (N_25757,N_21579,N_18082);
xor U25758 (N_25758,N_21773,N_23990);
and U25759 (N_25759,N_23511,N_21428);
nor U25760 (N_25760,N_19631,N_22477);
nor U25761 (N_25761,N_19648,N_20357);
nand U25762 (N_25762,N_22757,N_22536);
xor U25763 (N_25763,N_18182,N_22694);
and U25764 (N_25764,N_19821,N_18664);
nand U25765 (N_25765,N_23763,N_20676);
nand U25766 (N_25766,N_22359,N_18134);
nand U25767 (N_25767,N_23105,N_21216);
and U25768 (N_25768,N_23934,N_23569);
xnor U25769 (N_25769,N_18350,N_18781);
nor U25770 (N_25770,N_20877,N_23192);
or U25771 (N_25771,N_23238,N_18465);
xnor U25772 (N_25772,N_21699,N_18907);
nand U25773 (N_25773,N_19961,N_18755);
or U25774 (N_25774,N_19223,N_21871);
or U25775 (N_25775,N_21961,N_20019);
and U25776 (N_25776,N_23901,N_20914);
and U25777 (N_25777,N_18192,N_18245);
nand U25778 (N_25778,N_21930,N_20834);
xor U25779 (N_25779,N_18621,N_22243);
or U25780 (N_25780,N_23754,N_23879);
xnor U25781 (N_25781,N_20701,N_23379);
nor U25782 (N_25782,N_23003,N_21377);
or U25783 (N_25783,N_19465,N_22078);
and U25784 (N_25784,N_23919,N_18610);
or U25785 (N_25785,N_20292,N_21984);
or U25786 (N_25786,N_23868,N_19258);
and U25787 (N_25787,N_18663,N_19007);
nand U25788 (N_25788,N_23841,N_18445);
or U25789 (N_25789,N_19457,N_21152);
or U25790 (N_25790,N_23455,N_21534);
or U25791 (N_25791,N_23209,N_18330);
or U25792 (N_25792,N_22596,N_23502);
or U25793 (N_25793,N_21478,N_20655);
nand U25794 (N_25794,N_23336,N_23805);
and U25795 (N_25795,N_21408,N_22514);
and U25796 (N_25796,N_18035,N_18407);
nor U25797 (N_25797,N_18759,N_22255);
and U25798 (N_25798,N_21558,N_22196);
or U25799 (N_25799,N_18816,N_19311);
xor U25800 (N_25800,N_20058,N_18734);
and U25801 (N_25801,N_20088,N_22207);
and U25802 (N_25802,N_19157,N_20096);
nand U25803 (N_25803,N_18635,N_22084);
nand U25804 (N_25804,N_19706,N_19467);
nand U25805 (N_25805,N_23013,N_19208);
and U25806 (N_25806,N_23153,N_22655);
nand U25807 (N_25807,N_21808,N_20260);
xor U25808 (N_25808,N_22649,N_21499);
nor U25809 (N_25809,N_23475,N_23081);
and U25810 (N_25810,N_18207,N_18151);
and U25811 (N_25811,N_19284,N_18665);
nor U25812 (N_25812,N_18869,N_20333);
xnor U25813 (N_25813,N_23180,N_19042);
nand U25814 (N_25814,N_21509,N_19019);
nand U25815 (N_25815,N_20267,N_18498);
nand U25816 (N_25816,N_19172,N_20130);
nand U25817 (N_25817,N_20081,N_22306);
nor U25818 (N_25818,N_18707,N_18078);
and U25819 (N_25819,N_19397,N_20729);
nor U25820 (N_25820,N_21044,N_22469);
nand U25821 (N_25821,N_20363,N_20434);
or U25822 (N_25822,N_20400,N_18984);
nand U25823 (N_25823,N_20957,N_18830);
nand U25824 (N_25824,N_19430,N_21825);
and U25825 (N_25825,N_23404,N_19614);
nor U25826 (N_25826,N_20105,N_22505);
nor U25827 (N_25827,N_20952,N_20679);
and U25828 (N_25828,N_21116,N_18566);
nand U25829 (N_25829,N_22030,N_22005);
nand U25830 (N_25830,N_22911,N_20545);
nor U25831 (N_25831,N_18528,N_22386);
xor U25832 (N_25832,N_19515,N_18976);
xnor U25833 (N_25833,N_23972,N_19313);
xor U25834 (N_25834,N_23718,N_23240);
or U25835 (N_25835,N_22991,N_18165);
nand U25836 (N_25836,N_20247,N_19909);
and U25837 (N_25837,N_21118,N_21511);
and U25838 (N_25838,N_21418,N_20826);
xor U25839 (N_25839,N_23267,N_18459);
nand U25840 (N_25840,N_22726,N_23131);
nor U25841 (N_25841,N_18912,N_19183);
or U25842 (N_25842,N_19937,N_18297);
nor U25843 (N_25843,N_18927,N_20287);
and U25844 (N_25844,N_19512,N_23863);
or U25845 (N_25845,N_21091,N_23028);
nor U25846 (N_25846,N_23662,N_21600);
xnor U25847 (N_25847,N_20642,N_19018);
and U25848 (N_25848,N_23178,N_21243);
nand U25849 (N_25849,N_19067,N_23625);
or U25850 (N_25850,N_22591,N_21269);
or U25851 (N_25851,N_22864,N_19182);
or U25852 (N_25852,N_19633,N_21096);
nand U25853 (N_25853,N_23507,N_19262);
nand U25854 (N_25854,N_18319,N_23807);
and U25855 (N_25855,N_23217,N_20691);
nor U25856 (N_25856,N_21952,N_23428);
and U25857 (N_25857,N_22507,N_22623);
nor U25858 (N_25858,N_20277,N_23784);
xnor U25859 (N_25859,N_20574,N_22210);
and U25860 (N_25860,N_22661,N_23768);
and U25861 (N_25861,N_22476,N_23594);
or U25862 (N_25862,N_22849,N_22385);
and U25863 (N_25863,N_21275,N_21660);
nor U25864 (N_25864,N_18144,N_21935);
or U25865 (N_25865,N_18414,N_18320);
or U25866 (N_25866,N_19453,N_20414);
or U25867 (N_25867,N_22314,N_20258);
and U25868 (N_25868,N_19559,N_22615);
xor U25869 (N_25869,N_22399,N_23009);
and U25870 (N_25870,N_22021,N_22281);
xnor U25871 (N_25871,N_21211,N_23998);
or U25872 (N_25872,N_20114,N_20091);
and U25873 (N_25873,N_21265,N_18698);
nand U25874 (N_25874,N_20315,N_23642);
xnor U25875 (N_25875,N_18716,N_20010);
nor U25876 (N_25876,N_18267,N_23694);
and U25877 (N_25877,N_19845,N_19997);
or U25878 (N_25878,N_20352,N_18658);
and U25879 (N_25879,N_21217,N_22361);
nor U25880 (N_25880,N_20625,N_19965);
nor U25881 (N_25881,N_20687,N_19211);
nor U25882 (N_25882,N_19325,N_23356);
or U25883 (N_25883,N_18575,N_23735);
nor U25884 (N_25884,N_18472,N_18334);
and U25885 (N_25885,N_23520,N_18470);
nor U25886 (N_25886,N_18315,N_20839);
nand U25887 (N_25887,N_21893,N_19179);
and U25888 (N_25888,N_18532,N_20405);
nor U25889 (N_25889,N_22472,N_21617);
and U25890 (N_25890,N_18660,N_23873);
nor U25891 (N_25891,N_20989,N_18714);
and U25892 (N_25892,N_23435,N_21535);
nor U25893 (N_25893,N_21970,N_19516);
nor U25894 (N_25894,N_21005,N_19139);
xnor U25895 (N_25895,N_21420,N_23484);
and U25896 (N_25896,N_19688,N_23270);
nand U25897 (N_25897,N_18741,N_19740);
xor U25898 (N_25898,N_19372,N_22725);
or U25899 (N_25899,N_20083,N_21500);
and U25900 (N_25900,N_21282,N_21485);
or U25901 (N_25901,N_18105,N_20420);
or U25902 (N_25902,N_19949,N_23471);
and U25903 (N_25903,N_22073,N_23353);
nand U25904 (N_25904,N_21986,N_22665);
nor U25905 (N_25905,N_22128,N_20986);
xnor U25906 (N_25906,N_21742,N_21962);
and U25907 (N_25907,N_20474,N_22188);
or U25908 (N_25908,N_22443,N_19068);
nor U25909 (N_25909,N_20253,N_20502);
nor U25910 (N_25910,N_23226,N_19495);
or U25911 (N_25911,N_18868,N_20681);
nand U25912 (N_25912,N_20194,N_21322);
and U25913 (N_25913,N_20594,N_19115);
nor U25914 (N_25914,N_21267,N_22409);
nand U25915 (N_25915,N_19972,N_21648);
nor U25916 (N_25916,N_23743,N_22356);
or U25917 (N_25917,N_22564,N_20608);
nor U25918 (N_25918,N_23116,N_22209);
nor U25919 (N_25919,N_18416,N_22830);
or U25920 (N_25920,N_21766,N_23506);
and U25921 (N_25921,N_22350,N_23779);
nand U25922 (N_25922,N_18540,N_22933);
nand U25923 (N_25923,N_21745,N_20054);
nor U25924 (N_25924,N_21132,N_19163);
nor U25925 (N_25925,N_18690,N_22816);
or U25926 (N_25926,N_19750,N_19995);
nor U25927 (N_25927,N_22910,N_20510);
or U25928 (N_25928,N_19332,N_18776);
xor U25929 (N_25929,N_20726,N_21852);
nor U25930 (N_25930,N_21566,N_18208);
nor U25931 (N_25931,N_20421,N_23322);
xor U25932 (N_25932,N_23315,N_19878);
nand U25933 (N_25933,N_23274,N_22390);
or U25934 (N_25934,N_23974,N_21257);
or U25935 (N_25935,N_23644,N_18712);
nand U25936 (N_25936,N_20481,N_22179);
nand U25937 (N_25937,N_20191,N_18914);
nor U25938 (N_25938,N_20343,N_20505);
or U25939 (N_25939,N_22732,N_18531);
nand U25940 (N_25940,N_20848,N_19367);
and U25941 (N_25941,N_18051,N_22645);
or U25942 (N_25942,N_18673,N_19013);
xor U25943 (N_25943,N_21047,N_21832);
or U25944 (N_25944,N_18152,N_23340);
or U25945 (N_25945,N_21679,N_21813);
and U25946 (N_25946,N_19991,N_23190);
and U25947 (N_25947,N_23882,N_19825);
nand U25948 (N_25948,N_19770,N_19078);
xor U25949 (N_25949,N_22162,N_19699);
nand U25950 (N_25950,N_23894,N_22908);
and U25951 (N_25951,N_19271,N_22430);
nor U25952 (N_25952,N_22776,N_18325);
nand U25953 (N_25953,N_20001,N_23241);
nor U25954 (N_25954,N_18492,N_22999);
nand U25955 (N_25955,N_18122,N_22009);
xor U25956 (N_25956,N_20552,N_19585);
or U25957 (N_25957,N_18711,N_21695);
or U25958 (N_25958,N_20147,N_22928);
and U25959 (N_25959,N_21209,N_18846);
or U25960 (N_25960,N_22936,N_21198);
or U25961 (N_25961,N_20276,N_20824);
and U25962 (N_25962,N_22090,N_18413);
nor U25963 (N_25963,N_23645,N_18876);
nor U25964 (N_25964,N_22267,N_23250);
and U25965 (N_25965,N_21442,N_19858);
nor U25966 (N_25966,N_18600,N_18359);
and U25967 (N_25967,N_21784,N_19274);
nand U25968 (N_25968,N_19424,N_22971);
nor U25969 (N_25969,N_22739,N_21748);
and U25970 (N_25970,N_22853,N_21578);
nor U25971 (N_25971,N_23364,N_19247);
or U25972 (N_25972,N_20956,N_19520);
and U25973 (N_25973,N_21886,N_18691);
xnor U25974 (N_25974,N_23323,N_22208);
or U25975 (N_25975,N_20524,N_18421);
nor U25976 (N_25976,N_18604,N_19597);
or U25977 (N_25977,N_18733,N_18899);
or U25978 (N_25978,N_19591,N_23711);
nand U25979 (N_25979,N_23243,N_19189);
or U25980 (N_25980,N_21570,N_23567);
or U25981 (N_25981,N_23836,N_19941);
and U25982 (N_25982,N_18406,N_23288);
nand U25983 (N_25983,N_18535,N_19317);
nor U25984 (N_25984,N_23317,N_18880);
or U25985 (N_25985,N_22972,N_18719);
or U25986 (N_25986,N_22131,N_22634);
nor U25987 (N_25987,N_18163,N_23278);
nand U25988 (N_25988,N_21342,N_20199);
and U25989 (N_25989,N_19256,N_23760);
xnor U25990 (N_25990,N_22858,N_22841);
nor U25991 (N_25991,N_18387,N_18333);
xor U25992 (N_25992,N_21133,N_20045);
and U25993 (N_25993,N_20380,N_20190);
xnor U25994 (N_25994,N_19557,N_20281);
nand U25995 (N_25995,N_20329,N_19741);
nor U25996 (N_25996,N_20853,N_19144);
nand U25997 (N_25997,N_18274,N_18496);
nor U25998 (N_25998,N_19957,N_20345);
nor U25999 (N_25999,N_22140,N_22692);
and U26000 (N_26000,N_18917,N_21899);
nor U26001 (N_26001,N_23467,N_20980);
or U26002 (N_26002,N_19762,N_19333);
nand U26003 (N_26003,N_19532,N_21639);
and U26004 (N_26004,N_19048,N_22542);
nand U26005 (N_26005,N_22251,N_20534);
nor U26006 (N_26006,N_18241,N_18263);
or U26007 (N_26007,N_20678,N_20539);
nand U26008 (N_26008,N_20864,N_23703);
xor U26009 (N_26009,N_19485,N_18790);
xnor U26010 (N_26010,N_23751,N_20138);
or U26011 (N_26011,N_20857,N_20450);
xnor U26012 (N_26012,N_18415,N_18196);
and U26013 (N_26013,N_20141,N_20621);
or U26014 (N_26014,N_21072,N_21025);
nand U26015 (N_26015,N_19259,N_22033);
nand U26016 (N_26016,N_23591,N_19658);
nand U26017 (N_26017,N_23576,N_22190);
and U26018 (N_26018,N_20482,N_22553);
nand U26019 (N_26019,N_19789,N_19220);
or U26020 (N_26020,N_20734,N_20467);
xnor U26021 (N_26021,N_23533,N_19051);
or U26022 (N_26022,N_23714,N_23290);
or U26023 (N_26023,N_21065,N_18262);
nand U26024 (N_26024,N_21035,N_20896);
nand U26025 (N_26025,N_23924,N_23748);
nand U26026 (N_26026,N_19818,N_23166);
and U26027 (N_26027,N_19758,N_19874);
and U26028 (N_26028,N_20531,N_21004);
or U26029 (N_26029,N_22474,N_20953);
nor U26030 (N_26030,N_18460,N_22717);
nand U26031 (N_26031,N_21971,N_23011);
or U26032 (N_26032,N_22820,N_19590);
nand U26033 (N_26033,N_20805,N_20595);
and U26034 (N_26034,N_20317,N_21351);
xor U26035 (N_26035,N_23597,N_19502);
and U26036 (N_26036,N_22435,N_23415);
and U26037 (N_26037,N_18269,N_20246);
nand U26038 (N_26038,N_23010,N_19540);
or U26039 (N_26039,N_23559,N_18046);
and U26040 (N_26040,N_19820,N_22922);
and U26041 (N_26041,N_21521,N_22712);
nand U26042 (N_26042,N_22535,N_20692);
nand U26043 (N_26043,N_23298,N_18458);
xnor U26044 (N_26044,N_22277,N_20271);
and U26045 (N_26045,N_22862,N_21835);
nor U26046 (N_26046,N_23488,N_21108);
nor U26047 (N_26047,N_18889,N_21829);
and U26048 (N_26048,N_22785,N_22998);
and U26049 (N_26049,N_18476,N_23510);
nor U26050 (N_26050,N_22773,N_20626);
nor U26051 (N_26051,N_20046,N_19381);
and U26052 (N_26052,N_23170,N_18553);
and U26053 (N_26053,N_22783,N_19193);
nor U26054 (N_26054,N_23552,N_21274);
nand U26055 (N_26055,N_23140,N_23414);
and U26056 (N_26056,N_19708,N_19714);
or U26057 (N_26057,N_23699,N_19257);
and U26058 (N_26058,N_21306,N_18295);
or U26059 (N_26059,N_20802,N_23176);
and U26060 (N_26060,N_23789,N_23210);
or U26061 (N_26061,N_23049,N_22713);
or U26062 (N_26062,N_23681,N_20066);
nand U26063 (N_26063,N_22417,N_23893);
and U26064 (N_26064,N_20672,N_18541);
xnor U26065 (N_26065,N_18717,N_19653);
nor U26066 (N_26066,N_18860,N_21470);
nand U26067 (N_26067,N_22509,N_19447);
nor U26068 (N_26068,N_18124,N_18853);
nor U26069 (N_26069,N_21057,N_18177);
or U26070 (N_26070,N_18645,N_19788);
and U26071 (N_26071,N_18648,N_20523);
or U26072 (N_26072,N_20988,N_20061);
nand U26073 (N_26073,N_22470,N_18572);
nand U26074 (N_26074,N_19140,N_21733);
nand U26075 (N_26075,N_23620,N_19030);
and U26076 (N_26076,N_18587,N_23613);
or U26077 (N_26077,N_18559,N_22604);
nor U26078 (N_26078,N_22838,N_19807);
nor U26079 (N_26079,N_21819,N_19231);
nand U26080 (N_26080,N_23623,N_19599);
and U26081 (N_26081,N_18131,N_18043);
nand U26082 (N_26082,N_19050,N_22157);
nor U26083 (N_26083,N_21831,N_20959);
nor U26084 (N_26084,N_19724,N_20569);
or U26085 (N_26085,N_19918,N_23909);
nor U26086 (N_26086,N_19500,N_18896);
and U26087 (N_26087,N_21702,N_19350);
nand U26088 (N_26088,N_18632,N_21731);
nand U26089 (N_26089,N_20885,N_19711);
nand U26090 (N_26090,N_19073,N_23172);
nor U26091 (N_26091,N_21676,N_21066);
nand U26092 (N_26092,N_20078,N_22962);
nand U26093 (N_26093,N_22002,N_18858);
nor U26094 (N_26094,N_22279,N_20031);
or U26095 (N_26095,N_22343,N_18891);
nand U26096 (N_26096,N_21157,N_20969);
nor U26097 (N_26097,N_20018,N_21225);
or U26098 (N_26098,N_21190,N_20193);
or U26099 (N_26099,N_19772,N_18034);
or U26100 (N_26100,N_20720,N_20984);
nand U26101 (N_26101,N_20369,N_21833);
or U26102 (N_26102,N_22070,N_21213);
and U26103 (N_26103,N_21782,N_19831);
or U26104 (N_26104,N_23230,N_21938);
and U26105 (N_26105,N_21626,N_22872);
xnor U26106 (N_26106,N_22265,N_22052);
nand U26107 (N_26107,N_22302,N_19377);
nor U26108 (N_26108,N_23765,N_20756);
xnor U26109 (N_26109,N_18181,N_23208);
and U26110 (N_26110,N_20232,N_18383);
nand U26111 (N_26111,N_23599,N_22382);
and U26112 (N_26112,N_19261,N_23406);
and U26113 (N_26113,N_19323,N_20895);
or U26114 (N_26114,N_19927,N_23602);
nor U26115 (N_26115,N_20599,N_20843);
or U26116 (N_26116,N_20338,N_19851);
or U26117 (N_26117,N_21383,N_19039);
and U26118 (N_26118,N_20303,N_21224);
nor U26119 (N_26119,N_19932,N_23843);
xnor U26120 (N_26120,N_23157,N_20718);
nor U26121 (N_26121,N_22015,N_18235);
nor U26122 (N_26122,N_21857,N_20613);
nand U26123 (N_26123,N_20035,N_21167);
or U26124 (N_26124,N_21696,N_19859);
nand U26125 (N_26125,N_18617,N_18815);
or U26126 (N_26126,N_20439,N_21384);
and U26127 (N_26127,N_19298,N_22953);
or U26128 (N_26128,N_21374,N_21078);
nand U26129 (N_26129,N_20735,N_22585);
and U26130 (N_26130,N_23436,N_19121);
nor U26131 (N_26131,N_19174,N_23601);
nor U26132 (N_26132,N_20344,N_22284);
and U26133 (N_26133,N_23589,N_23111);
nor U26134 (N_26134,N_21107,N_18913);
or U26135 (N_26135,N_20712,N_22217);
nand U26136 (N_26136,N_21924,N_21965);
nor U26137 (N_26137,N_19616,N_22455);
nor U26138 (N_26138,N_21595,N_18091);
and U26139 (N_26139,N_18031,N_19399);
or U26140 (N_26140,N_21767,N_22237);
nand U26141 (N_26141,N_18791,N_19314);
or U26142 (N_26142,N_21147,N_21856);
or U26143 (N_26143,N_21456,N_21360);
nor U26144 (N_26144,N_22815,N_19488);
nor U26145 (N_26145,N_18794,N_20219);
and U26146 (N_26146,N_20269,N_18161);
xnor U26147 (N_26147,N_18808,N_21128);
nor U26148 (N_26148,N_23739,N_18250);
nor U26149 (N_26149,N_23737,N_19951);
or U26150 (N_26150,N_22116,N_22049);
or U26151 (N_26151,N_23900,N_21253);
xnor U26152 (N_26152,N_18206,N_19682);
nand U26153 (N_26153,N_20188,N_23494);
and U26154 (N_26154,N_23053,N_22442);
nor U26155 (N_26155,N_19309,N_21934);
nand U26156 (N_26156,N_23634,N_19655);
nor U26157 (N_26157,N_23989,N_18545);
nand U26158 (N_26158,N_20833,N_21088);
nor U26159 (N_26159,N_21682,N_21791);
and U26160 (N_26160,N_22094,N_22597);
xnor U26161 (N_26161,N_18030,N_23372);
and U26162 (N_26162,N_22380,N_18837);
nor U26163 (N_26163,N_19940,N_18613);
and U26164 (N_26164,N_21367,N_22275);
nand U26165 (N_26165,N_21135,N_18849);
xor U26166 (N_26166,N_20916,N_18068);
or U26167 (N_26167,N_18349,N_18692);
and U26168 (N_26168,N_18609,N_22901);
nor U26169 (N_26169,N_21363,N_21490);
and U26170 (N_26170,N_18630,N_18647);
and U26171 (N_26171,N_18560,N_19260);
nor U26172 (N_26172,N_23341,N_20452);
and U26173 (N_26173,N_19617,N_22974);
nand U26174 (N_26174,N_23692,N_23907);
or U26175 (N_26175,N_20370,N_18123);
nor U26176 (N_26176,N_18120,N_20416);
nand U26177 (N_26177,N_21998,N_19358);
nor U26178 (N_26178,N_20217,N_21704);
and U26179 (N_26179,N_22132,N_21328);
or U26180 (N_26180,N_20781,N_21231);
nor U26181 (N_26181,N_23969,N_22866);
xor U26182 (N_26182,N_19824,N_21757);
nand U26183 (N_26183,N_22305,N_18197);
or U26184 (N_26184,N_18098,N_23558);
nor U26185 (N_26185,N_19275,N_21234);
nor U26186 (N_26186,N_21458,N_21927);
and U26187 (N_26187,N_21564,N_22324);
nand U26188 (N_26188,N_20583,N_19908);
and U26189 (N_26189,N_22300,N_22287);
nand U26190 (N_26190,N_21008,N_22730);
nor U26191 (N_26191,N_19871,N_21803);
or U26192 (N_26192,N_20207,N_21153);
nand U26193 (N_26193,N_20092,N_22379);
and U26194 (N_26194,N_19757,N_23047);
and U26195 (N_26195,N_22540,N_18695);
and U26196 (N_26196,N_19486,N_18897);
and U26197 (N_26197,N_18360,N_23158);
nor U26198 (N_26198,N_18222,N_21215);
nor U26199 (N_26199,N_19203,N_23562);
nor U26200 (N_26200,N_20175,N_19689);
and U26201 (N_26201,N_20930,N_23858);
and U26202 (N_26202,N_23884,N_22489);
nand U26203 (N_26203,N_22183,N_19833);
or U26204 (N_26204,N_19349,N_22461);
and U26205 (N_26205,N_20872,N_23486);
nand U26206 (N_26206,N_22488,N_19036);
or U26207 (N_26207,N_18071,N_20610);
and U26208 (N_26208,N_22554,N_21480);
and U26209 (N_26209,N_23896,N_20996);
and U26210 (N_26210,N_21865,N_20717);
xor U26211 (N_26211,N_23333,N_21633);
nand U26212 (N_26212,N_23609,N_23531);
nor U26213 (N_26213,N_20026,N_23314);
and U26214 (N_26214,N_18715,N_19952);
and U26215 (N_26215,N_20667,N_22927);
nand U26216 (N_26216,N_21642,N_22337);
nor U26217 (N_26217,N_18725,N_21473);
and U26218 (N_26218,N_21882,N_21236);
nand U26219 (N_26219,N_21037,N_18279);
nor U26220 (N_26220,N_20280,N_22391);
nor U26221 (N_26221,N_22121,N_19060);
nand U26222 (N_26222,N_18363,N_20806);
or U26223 (N_26223,N_23653,N_20628);
or U26224 (N_26224,N_21181,N_23525);
or U26225 (N_26225,N_19707,N_18242);
or U26226 (N_26226,N_18157,N_21196);
nand U26227 (N_26227,N_23453,N_22952);
nor U26228 (N_26228,N_23854,N_18546);
or U26229 (N_26229,N_22412,N_23229);
or U26230 (N_26230,N_19383,N_18850);
or U26231 (N_26231,N_23254,N_19501);
xor U26232 (N_26232,N_22139,N_23331);
xnor U26233 (N_26233,N_23211,N_22018);
or U26234 (N_26234,N_23885,N_19286);
nand U26235 (N_26235,N_21068,N_21283);
or U26236 (N_26236,N_23855,N_20215);
nor U26237 (N_26237,N_18611,N_22651);
xor U26238 (N_26238,N_18749,N_18309);
or U26239 (N_26239,N_23715,N_22954);
xnor U26240 (N_26240,N_20696,N_20571);
nor U26241 (N_26241,N_19627,N_21581);
and U26242 (N_26242,N_21873,N_19583);
or U26243 (N_26243,N_19634,N_23273);
xor U26244 (N_26244,N_21591,N_22102);
nor U26245 (N_26245,N_21510,N_22552);
and U26246 (N_26246,N_20339,N_20882);
xnor U26247 (N_26247,N_20680,N_23062);
nand U26248 (N_26248,N_23309,N_19353);
nor U26249 (N_26249,N_23712,N_22672);
xor U26250 (N_26250,N_22886,N_21385);
and U26251 (N_26251,N_18500,N_22371);
and U26252 (N_26252,N_23588,N_20938);
nand U26253 (N_26253,N_21006,N_22965);
nor U26254 (N_26254,N_20674,N_20330);
nand U26255 (N_26255,N_22772,N_22268);
or U26256 (N_26256,N_18220,N_21948);
nor U26257 (N_26257,N_21227,N_23913);
nor U26258 (N_26258,N_18132,N_20077);
and U26259 (N_26259,N_23380,N_18176);
nand U26260 (N_26260,N_18903,N_19982);
and U26261 (N_26261,N_20410,N_21016);
and U26262 (N_26262,N_21903,N_19490);
nand U26263 (N_26263,N_23277,N_18654);
and U26264 (N_26264,N_23050,N_18237);
xor U26265 (N_26265,N_19375,N_18236);
nor U26266 (N_26266,N_23962,N_19763);
and U26267 (N_26267,N_23773,N_20328);
nor U26268 (N_26268,N_21750,N_20713);
nand U26269 (N_26269,N_20700,N_19572);
or U26270 (N_26270,N_19159,N_22355);
nand U26271 (N_26271,N_18187,N_19837);
and U26272 (N_26272,N_19834,N_20892);
and U26273 (N_26273,N_20316,N_23690);
nand U26274 (N_26274,N_18614,N_22014);
nand U26275 (N_26275,N_22436,N_18328);
nand U26276 (N_26276,N_23038,N_22024);
xor U26277 (N_26277,N_22682,N_22740);
nor U26278 (N_26278,N_18990,N_21807);
nand U26279 (N_26279,N_23514,N_20556);
and U26280 (N_26280,N_19913,N_23181);
and U26281 (N_26281,N_19319,N_23235);
or U26282 (N_26282,N_18070,N_23664);
nand U26283 (N_26283,N_19117,N_18299);
nor U26284 (N_26284,N_22759,N_23682);
or U26285 (N_26285,N_22642,N_23301);
nand U26286 (N_26286,N_22831,N_22641);
nor U26287 (N_26287,N_21712,N_18368);
nor U26288 (N_26288,N_18307,N_18367);
and U26289 (N_26289,N_22097,N_21772);
nand U26290 (N_26290,N_18234,N_20767);
or U26291 (N_26291,N_19567,N_19449);
and U26292 (N_26292,N_22039,N_23173);
nor U26293 (N_26293,N_23377,N_23941);
nand U26294 (N_26294,N_18519,N_23189);
nand U26295 (N_26295,N_21019,N_22657);
or U26296 (N_26296,N_19464,N_23632);
nor U26297 (N_26297,N_18595,N_19069);
or U26298 (N_26298,N_20160,N_21643);
or U26299 (N_26299,N_20437,N_18510);
or U26300 (N_26300,N_20838,N_22325);
nand U26301 (N_26301,N_19606,N_18067);
and U26302 (N_26302,N_20525,N_21366);
and U26303 (N_26303,N_22141,N_18838);
nor U26304 (N_26304,N_20866,N_20489);
xnor U26305 (N_26305,N_18355,N_18339);
nand U26306 (N_26306,N_18204,N_18542);
and U26307 (N_26307,N_23795,N_18289);
and U26308 (N_26308,N_23251,N_19962);
nor U26309 (N_26309,N_22238,N_20422);
nor U26310 (N_26310,N_22770,N_22025);
nor U26311 (N_26311,N_20480,N_20580);
nor U26312 (N_26312,N_21798,N_18565);
nand U26313 (N_26313,N_23442,N_19622);
nand U26314 (N_26314,N_19080,N_19849);
or U26315 (N_26315,N_18977,N_18159);
nand U26316 (N_26316,N_21318,N_23204);
nand U26317 (N_26317,N_21028,N_22595);
or U26318 (N_26318,N_23302,N_21826);
and U26319 (N_26319,N_19386,N_20218);
xnor U26320 (N_26320,N_19771,N_23667);
nand U26321 (N_26321,N_20465,N_23228);
and U26322 (N_26322,N_22590,N_19407);
and U26323 (N_26323,N_18190,N_18169);
nand U26324 (N_26324,N_23086,N_18261);
nor U26325 (N_26325,N_22771,N_22537);
nand U26326 (N_26326,N_18602,N_23814);
nor U26327 (N_26327,N_23587,N_20210);
or U26328 (N_26328,N_22629,N_21634);
or U26329 (N_26329,N_20879,N_21272);
nand U26330 (N_26330,N_19810,N_18229);
nor U26331 (N_26331,N_20519,N_21244);
and U26332 (N_26332,N_23996,N_23008);
and U26333 (N_26333,N_22877,N_20347);
and U26334 (N_26334,N_21124,N_20391);
or U26335 (N_26335,N_19385,N_18596);
nand U26336 (N_26336,N_20981,N_18636);
and U26337 (N_26337,N_23082,N_19245);
nand U26338 (N_26338,N_19891,N_19276);
or U26339 (N_26339,N_18488,N_18497);
nand U26340 (N_26340,N_18036,N_23186);
and U26341 (N_26341,N_21910,N_22282);
and U26342 (N_26342,N_20288,N_18392);
xor U26343 (N_26343,N_20722,N_19460);
and U26344 (N_26344,N_20106,N_22913);
nor U26345 (N_26345,N_21776,N_18443);
xnor U26346 (N_26346,N_20887,N_19462);
nor U26347 (N_26347,N_20780,N_18188);
or U26348 (N_26348,N_23133,N_23067);
nand U26349 (N_26349,N_20821,N_21501);
or U26350 (N_26350,N_18080,N_22036);
nor U26351 (N_26351,N_18592,N_18955);
or U26352 (N_26352,N_21586,N_20453);
xnor U26353 (N_26353,N_21237,N_19348);
and U26354 (N_26354,N_19710,N_20455);
nand U26355 (N_26355,N_22608,N_22851);
or U26356 (N_26356,N_21158,N_22860);
nor U26357 (N_26357,N_22150,N_20261);
nand U26358 (N_26358,N_23976,N_22979);
or U26359 (N_26359,N_22261,N_23721);
and U26360 (N_26360,N_23137,N_23162);
xnor U26361 (N_26361,N_19784,N_21608);
xor U26362 (N_26362,N_18828,N_22138);
nand U26363 (N_26363,N_21131,N_20641);
and U26364 (N_26364,N_20870,N_20059);
or U26365 (N_26365,N_21337,N_22318);
and U26366 (N_26366,N_21880,N_21080);
and U26367 (N_26367,N_20205,N_23378);
or U26368 (N_26368,N_21567,N_20603);
and U26369 (N_26369,N_22458,N_23827);
and U26370 (N_26370,N_21278,N_23917);
nand U26371 (N_26371,N_23772,N_22248);
nand U26372 (N_26372,N_18946,N_23437);
nor U26373 (N_26373,N_21338,N_23964);
xor U26374 (N_26374,N_21588,N_23152);
or U26375 (N_26375,N_22621,N_21386);
xor U26376 (N_26376,N_22673,N_18366);
nand U26377 (N_26377,N_22511,N_21560);
nor U26378 (N_26378,N_19404,N_19112);
and U26379 (N_26379,N_23347,N_23263);
xor U26380 (N_26380,N_21576,N_22950);
or U26381 (N_26381,N_21296,N_22797);
nor U26382 (N_26382,N_21556,N_23935);
and U26383 (N_26383,N_19938,N_19626);
and U26384 (N_26384,N_23175,N_21870);
or U26385 (N_26385,N_23080,N_21355);
and U26386 (N_26386,N_22652,N_23560);
nor U26387 (N_26387,N_22746,N_20372);
nand U26388 (N_26388,N_23496,N_23334);
nor U26389 (N_26389,N_20451,N_23828);
xor U26390 (N_26390,N_19720,N_21083);
nor U26391 (N_26391,N_22704,N_22892);
nor U26392 (N_26392,N_23729,N_19316);
and U26393 (N_26393,N_21711,N_19320);
and U26394 (N_26394,N_20181,N_21471);
xnor U26395 (N_26395,N_18463,N_20999);
nor U26396 (N_26396,N_18371,N_23821);
and U26397 (N_26397,N_22957,N_22448);
nor U26398 (N_26398,N_18063,N_18138);
nand U26399 (N_26399,N_20321,N_19670);
or U26400 (N_26400,N_19547,N_23824);
and U26401 (N_26401,N_21956,N_21371);
and U26402 (N_26402,N_20612,N_19694);
or U26403 (N_26403,N_23612,N_19023);
nand U26404 (N_26404,N_22301,N_19263);
nor U26405 (N_26405,N_20565,N_23985);
xnor U26406 (N_26406,N_19887,N_20183);
nand U26407 (N_26407,N_18803,N_21885);
and U26408 (N_26408,N_20060,N_23124);
or U26409 (N_26409,N_18915,N_21048);
nand U26410 (N_26410,N_23608,N_19249);
or U26411 (N_26411,N_20385,N_20874);
xor U26412 (N_26412,N_21649,N_21160);
nor U26413 (N_26413,N_21765,N_21592);
and U26414 (N_26414,N_19756,N_22333);
or U26415 (N_26415,N_21853,N_23957);
or U26416 (N_26416,N_23182,N_19513);
or U26417 (N_26417,N_20584,N_18678);
or U26418 (N_26418,N_20249,N_18311);
or U26419 (N_26419,N_19119,N_22941);
xor U26420 (N_26420,N_23268,N_19084);
and U26421 (N_26421,N_19024,N_19619);
xnor U26422 (N_26422,N_21043,N_23482);
or U26423 (N_26423,N_23171,N_19221);
and U26424 (N_26424,N_22937,N_22233);
or U26425 (N_26425,N_19733,N_18937);
and U26426 (N_26426,N_18646,N_21823);
nor U26427 (N_26427,N_22571,N_23939);
nand U26428 (N_26428,N_20086,N_23161);
nand U26429 (N_26429,N_20484,N_22845);
nor U26430 (N_26430,N_23077,N_22263);
xnor U26431 (N_26431,N_21315,N_21693);
or U26432 (N_26432,N_23628,N_23756);
or U26433 (N_26433,N_18111,N_19649);
nand U26434 (N_26434,N_21760,N_18855);
and U26435 (N_26435,N_19832,N_18936);
and U26436 (N_26436,N_19542,N_23956);
nor U26437 (N_26437,N_21524,N_22459);
nor U26438 (N_26438,N_21151,N_22428);
or U26439 (N_26439,N_21817,N_22669);
or U26440 (N_26440,N_22879,N_21238);
and U26441 (N_26441,N_19816,N_22918);
and U26442 (N_26442,N_21851,N_20711);
and U26443 (N_26443,N_20559,N_22605);
nor U26444 (N_26444,N_23498,N_21199);
nand U26445 (N_26445,N_23126,N_21106);
or U26446 (N_26446,N_20093,N_21650);
and U26447 (N_26447,N_23618,N_22351);
and U26448 (N_26448,N_18963,N_21678);
nor U26449 (N_26449,N_23846,N_21937);
nor U26450 (N_26450,N_19057,N_20946);
xor U26451 (N_26451,N_20563,N_21074);
nand U26452 (N_26452,N_19058,N_21320);
or U26453 (N_26453,N_18583,N_23649);
nor U26454 (N_26454,N_19593,N_22728);
and U26455 (N_26455,N_21922,N_22133);
nand U26456 (N_26456,N_21289,N_23060);
nand U26457 (N_26457,N_23476,N_18616);
or U26458 (N_26458,N_21058,N_21055);
and U26459 (N_26459,N_18214,N_22364);
nand U26460 (N_26460,N_18438,N_21881);
xnor U26461 (N_26461,N_21691,N_21052);
nand U26462 (N_26462,N_22055,N_18939);
nor U26463 (N_26463,N_19186,N_21381);
xor U26464 (N_26464,N_22720,N_19312);
or U26465 (N_26465,N_21801,N_21298);
and U26466 (N_26466,N_21053,N_23216);
and U26467 (N_26467,N_21312,N_19187);
and U26468 (N_26468,N_18327,N_20123);
nand U26469 (N_26469,N_22543,N_21445);
nand U26470 (N_26470,N_21023,N_19472);
nor U26471 (N_26471,N_19197,N_20413);
and U26472 (N_26472,N_22147,N_23373);
and U26473 (N_26473,N_21830,N_21847);
nor U26474 (N_26474,N_18130,N_23764);
nand U26475 (N_26475,N_21692,N_19079);
or U26476 (N_26476,N_19926,N_23202);
or U26477 (N_26477,N_20252,N_20883);
xor U26478 (N_26478,N_19840,N_18774);
and U26479 (N_26479,N_20418,N_19966);
and U26480 (N_26480,N_20845,N_21720);
and U26481 (N_26481,N_18326,N_21059);
and U26482 (N_26482,N_18216,N_22292);
and U26483 (N_26483,N_18142,N_21192);
nor U26484 (N_26484,N_23504,N_19766);
nand U26485 (N_26485,N_20504,N_19910);
nand U26486 (N_26486,N_18009,N_20832);
or U26487 (N_26487,N_21828,N_22087);
nand U26488 (N_26488,N_20998,N_19779);
nor U26489 (N_26489,N_23159,N_19987);
xor U26490 (N_26490,N_21465,N_23402);
nor U26491 (N_26491,N_23117,N_23221);
or U26492 (N_26492,N_21410,N_21309);
and U26493 (N_26493,N_19308,N_19029);
nand U26494 (N_26494,N_22376,N_21838);
or U26495 (N_26495,N_18900,N_22326);
nand U26496 (N_26496,N_22533,N_19110);
nand U26497 (N_26497,N_21493,N_22687);
and U26498 (N_26498,N_19782,N_18538);
nand U26499 (N_26499,N_20777,N_23556);
or U26500 (N_26500,N_21636,N_22341);
nor U26501 (N_26501,N_21163,N_19692);
and U26502 (N_26502,N_19329,N_23079);
or U26503 (N_26503,N_20127,N_23252);
or U26504 (N_26504,N_23564,N_20714);
nor U26505 (N_26505,N_18217,N_20171);
nand U26506 (N_26506,N_22581,N_20785);
and U26507 (N_26507,N_19921,N_21778);
and U26508 (N_26508,N_18420,N_23545);
nor U26509 (N_26509,N_22041,N_20283);
nand U26510 (N_26510,N_20233,N_23565);
or U26511 (N_26511,N_19657,N_19324);
or U26512 (N_26512,N_21982,N_23169);
and U26513 (N_26513,N_20100,N_21197);
or U26514 (N_26514,N_21399,N_18300);
and U26515 (N_26515,N_20908,N_22620);
nor U26516 (N_26516,N_22805,N_18374);
or U26517 (N_26517,N_18348,N_18266);
and U26518 (N_26518,N_22781,N_23691);
xor U26519 (N_26519,N_19867,N_20934);
nand U26520 (N_26520,N_20643,N_18487);
and U26521 (N_26521,N_19566,N_21010);
nand U26522 (N_26522,N_21508,N_23073);
xor U26523 (N_26523,N_22369,N_21707);
and U26524 (N_26524,N_20762,N_20131);
and U26525 (N_26525,N_20841,N_19145);
or U26526 (N_26526,N_20048,N_22648);
nor U26527 (N_26527,N_19767,N_19285);
xor U26528 (N_26528,N_22101,N_18375);
or U26529 (N_26529,N_21030,N_22057);
nor U26530 (N_26530,N_20775,N_19615);
or U26531 (N_26531,N_22671,N_18451);
nand U26532 (N_26532,N_20441,N_19783);
or U26533 (N_26533,N_20842,N_20587);
and U26534 (N_26534,N_20658,N_23358);
or U26535 (N_26535,N_18293,N_19347);
or U26536 (N_26536,N_20807,N_19113);
or U26537 (N_26537,N_18494,N_21896);
and U26538 (N_26538,N_23369,N_22996);
and U26539 (N_26539,N_18065,N_23430);
nor U26540 (N_26540,N_23734,N_23657);
and U26541 (N_26541,N_22871,N_20987);
nand U26542 (N_26542,N_23960,N_21918);
or U26543 (N_26543,N_19738,N_22975);
nor U26544 (N_26544,N_20248,N_18961);
nor U26545 (N_26545,N_21941,N_21012);
nand U26546 (N_26546,N_18212,N_23538);
or U26547 (N_26547,N_22164,N_18225);
and U26548 (N_26548,N_21316,N_19610);
and U26549 (N_26549,N_23325,N_18622);
nand U26550 (N_26550,N_23958,N_21294);
nand U26551 (N_26551,N_19522,N_23826);
and U26552 (N_26552,N_22080,N_23838);
nand U26553 (N_26553,N_19623,N_22258);
or U26554 (N_26554,N_22750,N_22956);
nor U26555 (N_26555,N_23853,N_22614);
nand U26556 (N_26556,N_20072,N_22861);
nand U26557 (N_26557,N_20408,N_22963);
xnor U26558 (N_26558,N_21212,N_22169);
xnor U26559 (N_26559,N_21474,N_19477);
nor U26560 (N_26560,N_18226,N_21486);
nand U26561 (N_26561,N_23922,N_21538);
nand U26562 (N_26562,N_21398,N_20268);
nor U26563 (N_26563,N_18694,N_19861);
and U26564 (N_26564,N_21928,N_19370);
nor U26565 (N_26565,N_18347,N_19356);
and U26566 (N_26566,N_19288,N_18773);
nor U26567 (N_26567,N_20985,N_23787);
xor U26568 (N_26568,N_22381,N_18357);
xor U26569 (N_26569,N_22495,N_19842);
nand U26570 (N_26570,N_20786,N_20320);
nand U26571 (N_26571,N_19791,N_18422);
xnor U26572 (N_26572,N_22982,N_19611);
nor U26573 (N_26573,N_20737,N_22930);
or U26574 (N_26574,N_23480,N_19993);
or U26575 (N_26575,N_20995,N_22008);
nand U26576 (N_26576,N_22336,N_20752);
or U26577 (N_26577,N_22151,N_20798);
or U26578 (N_26578,N_22256,N_18529);
xnor U26579 (N_26579,N_22471,N_21700);
and U26580 (N_26580,N_22487,N_23643);
nor U26581 (N_26581,N_18114,N_22271);
nor U26582 (N_26582,N_19072,N_18358);
nor U26583 (N_26583,N_19497,N_19595);
and U26584 (N_26584,N_20133,N_23793);
nand U26585 (N_26585,N_19137,N_20067);
nand U26586 (N_26586,N_21746,N_19545);
and U26587 (N_26587,N_22163,N_22034);
and U26588 (N_26588,N_18381,N_22729);
or U26589 (N_26589,N_20731,N_20302);
or U26590 (N_26590,N_21787,N_19032);
or U26591 (N_26591,N_22987,N_22022);
nor U26592 (N_26592,N_21963,N_19122);
and U26593 (N_26593,N_20472,N_19798);
nor U26594 (N_26594,N_22227,N_23778);
or U26595 (N_26595,N_19509,N_21554);
and U26596 (N_26596,N_18023,N_23020);
nand U26597 (N_26597,N_21532,N_22394);
nand U26598 (N_26598,N_19413,N_18154);
or U26599 (N_26599,N_18473,N_18085);
xor U26600 (N_26600,N_22622,N_18179);
or U26601 (N_26601,N_21291,N_23844);
and U26602 (N_26602,N_22142,N_19781);
xnor U26603 (N_26603,N_19291,N_18514);
nand U26604 (N_26604,N_21892,N_20683);
nor U26605 (N_26605,N_20755,N_18758);
nand U26606 (N_26606,N_20429,N_19421);
nor U26607 (N_26607,N_22445,N_22485);
or U26608 (N_26608,N_19801,N_21140);
xor U26609 (N_26609,N_22662,N_21605);
xnor U26610 (N_26610,N_19022,N_21797);
or U26611 (N_26611,N_21201,N_22439);
nor U26612 (N_26612,N_21479,N_18757);
and U26613 (N_26613,N_21627,N_23099);
and U26614 (N_26614,N_19422,N_23641);
and U26615 (N_26615,N_18045,N_19795);
xnor U26616 (N_26616,N_23401,N_22349);
nor U26617 (N_26617,N_18278,N_19872);
nand U26618 (N_26618,N_18205,N_18203);
and U26619 (N_26619,N_22108,N_21292);
nand U26620 (N_26620,N_23368,N_18390);
nor U26621 (N_26621,N_23454,N_22883);
xnor U26622 (N_26622,N_19236,N_19127);
nor U26623 (N_26623,N_18002,N_20250);
nor U26624 (N_26624,N_21463,N_23399);
or U26625 (N_26625,N_21724,N_23461);
nand U26626 (N_26626,N_20301,N_19390);
nand U26627 (N_26627,N_22678,N_23580);
nand U26628 (N_26628,N_23616,N_18789);
nor U26629 (N_26629,N_19428,N_19100);
nand U26630 (N_26630,N_18904,N_18843);
and U26631 (N_26631,N_23477,N_18594);
nand U26632 (N_26632,N_21396,N_22338);
or U26633 (N_26633,N_20682,N_18909);
nor U26634 (N_26634,N_22091,N_18453);
xnor U26635 (N_26635,N_20851,N_21664);
and U26636 (N_26636,N_20920,N_22899);
or U26637 (N_26637,N_20763,N_20118);
nand U26638 (N_26638,N_20053,N_23042);
nor U26639 (N_26639,N_19876,N_19357);
nand U26640 (N_26640,N_18117,N_18019);
nand U26641 (N_26641,N_18819,N_20153);
or U26642 (N_26642,N_20412,N_18243);
and U26643 (N_26643,N_22076,N_22964);
nand U26644 (N_26644,N_18922,N_18499);
and U26645 (N_26645,N_23405,N_19743);
and U26646 (N_26646,N_19573,N_22410);
nand U26647 (N_26647,N_21741,N_19538);
and U26648 (N_26648,N_18485,N_18631);
nand U26649 (N_26649,N_23758,N_21665);
nand U26650 (N_26650,N_19207,N_19450);
nand U26651 (N_26651,N_22599,N_22857);
nor U26652 (N_26652,N_21884,N_23548);
nor U26653 (N_26653,N_20143,N_19254);
nand U26654 (N_26654,N_18700,N_18985);
nor U26655 (N_26655,N_23582,N_22308);
and U26656 (N_26656,N_18615,N_22561);
nor U26657 (N_26657,N_23652,N_22113);
xnor U26658 (N_26658,N_20185,N_18322);
or U26659 (N_26659,N_18814,N_22042);
xnor U26660 (N_26660,N_22696,N_18442);
and U26661 (N_26661,N_22354,N_20606);
and U26662 (N_26662,N_19037,N_21180);
nor U26663 (N_26663,N_22817,N_20585);
nor U26664 (N_26664,N_20458,N_21860);
nand U26665 (N_26665,N_21812,N_19907);
nand U26666 (N_26666,N_21719,N_19690);
xnor U26667 (N_26667,N_21651,N_21032);
and U26668 (N_26668,N_21706,N_21583);
nand U26669 (N_26669,N_18526,N_20393);
xnor U26670 (N_26670,N_20554,N_23223);
and U26671 (N_26671,N_23450,N_19331);
and U26672 (N_26672,N_19749,N_21121);
and U26673 (N_26673,N_20111,N_18047);
nor U26674 (N_26674,N_23375,N_20645);
nand U26675 (N_26675,N_21245,N_21859);
nor U26676 (N_26676,N_19931,N_22332);
nor U26677 (N_26677,N_23948,N_21632);
and U26678 (N_26678,N_23637,N_21233);
and U26679 (N_26679,N_18972,N_23656);
nor U26680 (N_26680,N_19105,N_22249);
nand U26681 (N_26681,N_18303,N_22870);
and U26682 (N_26682,N_19360,N_21014);
and U26683 (N_26683,N_21249,N_21674);
nand U26684 (N_26684,N_18728,N_19970);
and U26685 (N_26685,N_23115,N_23951);
xnor U26686 (N_26686,N_20823,N_19723);
nor U26687 (N_26687,N_20746,N_19745);
and U26688 (N_26688,N_19679,N_18361);
nand U26689 (N_26689,N_23206,N_18186);
nand U26690 (N_26690,N_22811,N_22053);
or U26691 (N_26691,N_23606,N_21786);
nor U26692 (N_26692,N_22531,N_21800);
nor U26693 (N_26693,N_19093,N_23291);
or U26694 (N_26694,N_19503,N_21906);
or U26695 (N_26695,N_22215,N_18551);
or U26696 (N_26696,N_19452,N_18530);
and U26697 (N_26697,N_21525,N_18061);
nand U26698 (N_26698,N_23421,N_23928);
and U26699 (N_26699,N_18513,N_19662);
or U26700 (N_26700,N_18400,N_23679);
and U26701 (N_26701,N_23774,N_20404);
and U26702 (N_26702,N_23362,N_23367);
and U26703 (N_26703,N_22576,N_19852);
nand U26704 (N_26704,N_21324,N_23881);
and U26705 (N_26705,N_22031,N_23253);
or U26706 (N_26706,N_23304,N_23617);
and U26707 (N_26707,N_22766,N_23017);
or U26708 (N_26708,N_19158,N_20663);
nor U26709 (N_26709,N_18802,N_21555);
and U26710 (N_26710,N_23194,N_19008);
or U26711 (N_26711,N_22570,N_20622);
and U26712 (N_26712,N_20968,N_19638);
nand U26713 (N_26713,N_18845,N_23571);
and U26714 (N_26714,N_22919,N_23674);
and U26715 (N_26715,N_18590,N_19092);
nand U26716 (N_26716,N_20589,N_23043);
or U26717 (N_26717,N_21332,N_23622);
nor U26718 (N_26718,N_21226,N_22767);
nor U26719 (N_26719,N_22153,N_23319);
nand U26720 (N_26720,N_18929,N_19454);
nor U26721 (N_26721,N_21713,N_21841);
or U26722 (N_26722,N_20829,N_20849);
or U26723 (N_26723,N_20424,N_21271);
nor U26724 (N_26724,N_23337,N_21907);
xor U26725 (N_26725,N_22001,N_18882);
or U26726 (N_26726,N_18076,N_19109);
or U26727 (N_26727,N_18221,N_20758);
nand U26728 (N_26728,N_23057,N_20759);
nand U26729 (N_26729,N_20708,N_19483);
xor U26730 (N_26730,N_21959,N_21789);
xor U26731 (N_26731,N_23386,N_22427);
or U26732 (N_26732,N_19702,N_18099);
or U26733 (N_26733,N_23145,N_19659);
xnor U26734 (N_26734,N_23982,N_20364);
and U26735 (N_26735,N_18052,N_22072);
nor U26736 (N_26736,N_21663,N_22884);
or U26737 (N_26737,N_20818,N_19445);
and U26738 (N_26738,N_19549,N_23150);
and U26739 (N_26739,N_22555,N_22135);
xnor U26740 (N_26740,N_21958,N_19184);
and U26741 (N_26741,N_22801,N_20831);
nand U26742 (N_26742,N_23859,N_19769);
nand U26743 (N_26743,N_22598,N_18426);
xnor U26744 (N_26744,N_20156,N_19579);
nand U26745 (N_26745,N_20506,N_20122);
or U26746 (N_26746,N_19090,N_22932);
nand U26747 (N_26747,N_22606,N_21308);
or U26748 (N_26748,N_21031,N_18555);
or U26749 (N_26749,N_20800,N_22170);
nor U26750 (N_26750,N_21672,N_21411);
xnor U26751 (N_26751,N_20707,N_18475);
nor U26752 (N_26752,N_18405,N_22532);
nand U26753 (N_26753,N_21422,N_23688);
nand U26754 (N_26754,N_18523,N_18824);
or U26755 (N_26755,N_23321,N_20377);
or U26756 (N_26756,N_18966,N_18641);
nand U26757 (N_26757,N_22529,N_20813);
or U26758 (N_26758,N_20485,N_18726);
or U26759 (N_26759,N_22017,N_23123);
or U26760 (N_26760,N_22206,N_21730);
nor U26761 (N_26761,N_23986,N_23097);
nand U26762 (N_26762,N_19561,N_22074);
and U26763 (N_26763,N_18018,N_19436);
nand U26764 (N_26764,N_22434,N_20423);
nor U26765 (N_26765,N_20990,N_21394);
nor U26766 (N_26766,N_23429,N_20203);
and U26767 (N_26767,N_20978,N_23492);
or U26768 (N_26768,N_21909,N_18515);
xor U26769 (N_26769,N_21701,N_20165);
nor U26770 (N_26770,N_20903,N_19153);
nor U26771 (N_26771,N_18362,N_21983);
nor U26772 (N_26772,N_23813,N_19427);
nand U26773 (N_26773,N_23196,N_18053);
nor U26774 (N_26774,N_22734,N_20940);
and U26775 (N_26775,N_22689,N_23761);
nor U26776 (N_26776,N_18959,N_18856);
and U26777 (N_26777,N_23550,N_20675);
xor U26778 (N_26778,N_22056,N_23630);
and U26779 (N_26779,N_22038,N_19976);
or U26780 (N_26780,N_21540,N_19914);
and U26781 (N_26781,N_18586,N_19600);
or U26782 (N_26782,N_18988,N_19752);
nand U26783 (N_26783,N_20012,N_18495);
or U26784 (N_26784,N_19526,N_22075);
nor U26785 (N_26785,N_22848,N_21260);
nor U26786 (N_26786,N_23259,N_19219);
or U26787 (N_26787,N_21845,N_19915);
nor U26788 (N_26788,N_20214,N_18967);
nand U26789 (N_26789,N_19169,N_20098);
and U26790 (N_26790,N_18393,N_21985);
and U26791 (N_26791,N_23850,N_19241);
nand U26792 (N_26792,N_21144,N_21259);
nand U26793 (N_26793,N_21594,N_21406);
or U26794 (N_26794,N_23999,N_22486);
or U26795 (N_26795,N_23350,N_21345);
nand U26796 (N_26796,N_21070,N_20771);
and U26797 (N_26797,N_23344,N_23271);
nand U26798 (N_26798,N_22280,N_18745);
nand U26799 (N_26799,N_18310,N_19565);
and U26800 (N_26800,N_19863,N_21596);
or U26801 (N_26801,N_19804,N_19792);
nand U26802 (N_26802,N_21156,N_18461);
or U26803 (N_26803,N_21079,N_22839);
or U26804 (N_26804,N_21727,N_20225);
nor U26805 (N_26805,N_21631,N_23631);
nand U26806 (N_26806,N_23803,N_20337);
nor U26807 (N_26807,N_22468,N_21920);
or U26808 (N_26808,N_20204,N_22893);
nor U26809 (N_26809,N_18425,N_21709);
and U26810 (N_26810,N_23984,N_21112);
nand U26811 (N_26811,N_22160,N_18000);
or U26812 (N_26812,N_22452,N_20702);
nor U26813 (N_26813,N_23300,N_21313);
or U26814 (N_26814,N_18835,N_23895);
nor U26815 (N_26815,N_22867,N_23090);
nor U26816 (N_26816,N_22146,N_22837);
nand U26817 (N_26817,N_18919,N_20923);
or U26818 (N_26818,N_21297,N_23163);
nor U26819 (N_26819,N_19578,N_19087);
or U26820 (N_26820,N_19535,N_23348);
and U26821 (N_26821,N_23285,N_18591);
nor U26822 (N_26822,N_18626,N_22592);
and U26823 (N_26823,N_21533,N_23108);
nor U26824 (N_26824,N_23918,N_20639);
and U26825 (N_26825,N_19016,N_22699);
or U26826 (N_26826,N_22587,N_21978);
and U26827 (N_26827,N_22173,N_23791);
or U26828 (N_26828,N_21815,N_20575);
or U26829 (N_26829,N_22011,N_19482);
and U26830 (N_26830,N_20598,N_20326);
nor U26831 (N_26831,N_23799,N_23128);
and U26832 (N_26832,N_20134,N_19618);
or U26833 (N_26833,N_23036,N_21380);
and U26834 (N_26834,N_23546,N_22295);
xnor U26835 (N_26835,N_22638,N_23500);
or U26836 (N_26836,N_20279,N_19382);
nor U26837 (N_26837,N_19496,N_20745);
or U26838 (N_26838,N_22809,N_23746);
and U26839 (N_26839,N_20630,N_20686);
or U26840 (N_26840,N_22724,N_19446);
nand U26841 (N_26841,N_22579,N_18213);
or U26842 (N_26842,N_18435,N_20022);
and U26843 (N_26843,N_23110,N_21064);
or U26844 (N_26844,N_22743,N_18950);
nor U26845 (N_26845,N_20239,N_18509);
or U26846 (N_26846,N_23262,N_19226);
and U26847 (N_26847,N_18025,N_20693);
and U26848 (N_26848,N_18898,N_19283);
or U26849 (N_26849,N_19366,N_22610);
xnor U26850 (N_26850,N_18911,N_18095);
nand U26851 (N_26851,N_20407,N_19534);
or U26852 (N_26852,N_21195,N_20586);
or U26853 (N_26853,N_22676,N_22545);
nor U26854 (N_26854,N_21677,N_20501);
and U26855 (N_26855,N_20550,N_21708);
nor U26856 (N_26856,N_20155,N_19480);
nor U26857 (N_26857,N_19564,N_22144);
or U26858 (N_26858,N_22092,N_20650);
and U26859 (N_26859,N_22425,N_18074);
or U26860 (N_26860,N_22711,N_19083);
nand U26861 (N_26861,N_18894,N_19646);
nor U26862 (N_26862,N_23857,N_20255);
nand U26863 (N_26863,N_18096,N_23702);
and U26864 (N_26864,N_21625,N_20656);
and U26865 (N_26865,N_18992,N_18503);
and U26866 (N_26866,N_21753,N_22358);
nor U26867 (N_26867,N_18256,N_18230);
nand U26868 (N_26868,N_20112,N_20690);
nor U26869 (N_26869,N_18652,N_22050);
or U26870 (N_26870,N_19168,N_20651);
or U26871 (N_26871,N_19244,N_21542);
and U26872 (N_26872,N_19948,N_20349);
nand U26873 (N_26873,N_22808,N_21353);
nand U26874 (N_26874,N_20020,N_19364);
and U26875 (N_26875,N_22026,N_20113);
nor U26876 (N_26876,N_21460,N_19603);
nand U26877 (N_26877,N_19778,N_18020);
nor U26878 (N_26878,N_20270,N_21559);
and U26879 (N_26879,N_21908,N_21684);
or U26880 (N_26880,N_18191,N_22298);
and U26881 (N_26881,N_21715,N_19511);
xor U26882 (N_26882,N_19218,N_18508);
nor U26883 (N_26883,N_18158,N_20972);
nand U26884 (N_26884,N_18847,N_21369);
and U26885 (N_26885,N_23265,N_22125);
or U26886 (N_26886,N_20863,N_18502);
or U26887 (N_26887,N_22847,N_18948);
nor U26888 (N_26888,N_23581,N_18784);
and U26889 (N_26889,N_19828,N_20015);
nor U26890 (N_26890,N_18974,N_21955);
and U26891 (N_26891,N_23993,N_21864);
or U26892 (N_26892,N_20830,N_22155);
nor U26893 (N_26893,N_20173,N_22331);
nor U26894 (N_26894,N_18981,N_21145);
and U26895 (N_26895,N_23626,N_20102);
nor U26896 (N_26896,N_21368,N_21548);
or U26897 (N_26897,N_21686,N_20927);
nor U26898 (N_26898,N_18657,N_22093);
and U26899 (N_26899,N_21995,N_22440);
xor U26900 (N_26900,N_18178,N_18412);
xor U26901 (N_26901,N_21183,N_19968);
or U26902 (N_26902,N_18730,N_19266);
nor U26903 (N_26903,N_20576,N_22912);
nand U26904 (N_26904,N_21331,N_21863);
nand U26905 (N_26905,N_21557,N_18943);
nor U26906 (N_26906,N_22885,N_22245);
or U26907 (N_26907,N_22065,N_23233);
or U26908 (N_26908,N_20776,N_20044);
and U26909 (N_26909,N_18417,N_23383);
or U26910 (N_26910,N_19028,N_23730);
or U26911 (N_26911,N_19498,N_21459);
and U26912 (N_26912,N_23432,N_22697);
nor U26913 (N_26913,N_18945,N_21193);
nor U26914 (N_26914,N_21657,N_18168);
nand U26915 (N_26915,N_18001,N_19248);
and U26916 (N_26916,N_18986,N_22384);
xor U26917 (N_26917,N_18054,N_20744);
xnor U26918 (N_26918,N_22909,N_22166);
nand U26919 (N_26919,N_22451,N_18007);
and U26920 (N_26920,N_23155,N_22403);
and U26921 (N_26921,N_23762,N_19514);
and U26922 (N_26922,N_19736,N_20795);
nor U26923 (N_26923,N_22454,N_19551);
nand U26924 (N_26924,N_23338,N_23269);
nor U26925 (N_26925,N_18656,N_23593);
nor U26926 (N_26926,N_19726,N_23722);
or U26927 (N_26927,N_23980,N_20082);
and U26928 (N_26928,N_18544,N_18681);
xnor U26929 (N_26929,N_20796,N_19753);
nand U26930 (N_26930,N_21104,N_22619);
xnor U26931 (N_26931,N_18265,N_18276);
nor U26932 (N_26932,N_22339,N_18601);
and U26933 (N_26933,N_21795,N_21732);
or U26934 (N_26934,N_20888,N_19958);
and U26935 (N_26935,N_18162,N_21788);
xnor U26936 (N_26936,N_20871,N_21904);
nand U26937 (N_26937,N_22524,N_20008);
xnor U26938 (N_26938,N_23424,N_23095);
nor U26939 (N_26939,N_21191,N_22658);
nand U26940 (N_26940,N_20387,N_18150);
and U26941 (N_26941,N_18537,N_19017);
or U26942 (N_26942,N_20570,N_22283);
nand U26943 (N_26943,N_23396,N_21562);
or U26944 (N_26944,N_19306,N_23018);
nor U26945 (N_26945,N_20129,N_23040);
and U26946 (N_26946,N_22247,N_21872);
and U26947 (N_26947,N_23967,N_23800);
and U26948 (N_26948,N_20668,N_23666);
nand U26949 (N_26949,N_23434,N_21001);
and U26950 (N_26950,N_20254,N_18825);
or U26951 (N_26951,N_18777,N_22506);
xnor U26952 (N_26952,N_21667,N_23283);
and U26953 (N_26953,N_22089,N_21780);
nand U26954 (N_26954,N_18081,N_22028);
and U26955 (N_26955,N_21173,N_21968);
and U26956 (N_26956,N_19529,N_18028);
or U26957 (N_26957,N_19946,N_23448);
xnor U26958 (N_26958,N_19838,N_18093);
and U26959 (N_26959,N_18247,N_18703);
nand U26960 (N_26960,N_22806,N_18083);
and U26961 (N_26961,N_23218,N_23579);
and U26962 (N_26962,N_22889,N_23264);
xor U26963 (N_26963,N_19049,N_19190);
nor U26964 (N_26964,N_18450,N_23164);
nor U26965 (N_26965,N_20912,N_20170);
nand U26966 (N_26966,N_21989,N_21130);
nor U26967 (N_26967,N_20256,N_19142);
nand U26968 (N_26968,N_22491,N_20355);
or U26969 (N_26969,N_22578,N_23142);
nor U26970 (N_26970,N_22752,N_23139);
or U26971 (N_26971,N_20535,N_18517);
and U26972 (N_26972,N_22059,N_18661);
and U26973 (N_26973,N_19045,N_19046);
or U26974 (N_26974,N_19897,N_20604);
nand U26975 (N_26975,N_20910,N_19398);
nand U26976 (N_26976,N_19911,N_23775);
nand U26977 (N_26977,N_22763,N_22137);
or U26978 (N_26978,N_21602,N_23236);
nor U26979 (N_26979,N_23797,N_19727);
and U26980 (N_26980,N_19380,N_18022);
nor U26981 (N_26981,N_20944,N_21589);
nand U26982 (N_26982,N_22568,N_19476);
and U26983 (N_26983,N_23324,N_19844);
and U26984 (N_26984,N_23822,N_21936);
and U26985 (N_26985,N_20399,N_18506);
or U26986 (N_26986,N_21071,N_21821);
or U26987 (N_26987,N_23717,N_20620);
nand U26988 (N_26988,N_18248,N_18253);
nand U26989 (N_26989,N_23554,N_20666);
nand U26990 (N_26990,N_18166,N_23307);
nand U26991 (N_26991,N_23346,N_18686);
and U26992 (N_26992,N_18958,N_21268);
nand U26993 (N_26993,N_19354,N_20900);
nor U26994 (N_26994,N_18872,N_21610);
nor U26995 (N_26995,N_19880,N_23130);
or U26996 (N_26996,N_22526,N_23668);
nor U26997 (N_26997,N_22935,N_21689);
nor U26998 (N_26998,N_21607,N_18951);
nor U26999 (N_26999,N_18932,N_20742);
or U27000 (N_27000,N_18076,N_23981);
or U27001 (N_27001,N_22038,N_21801);
or U27002 (N_27002,N_21736,N_23268);
nand U27003 (N_27003,N_18947,N_23365);
and U27004 (N_27004,N_22328,N_20694);
xor U27005 (N_27005,N_21674,N_22731);
or U27006 (N_27006,N_23414,N_18779);
nor U27007 (N_27007,N_20670,N_19921);
nor U27008 (N_27008,N_22009,N_18780);
nor U27009 (N_27009,N_21798,N_22241);
and U27010 (N_27010,N_20367,N_22500);
and U27011 (N_27011,N_23712,N_18826);
and U27012 (N_27012,N_23182,N_21016);
nand U27013 (N_27013,N_22921,N_23406);
xor U27014 (N_27014,N_23555,N_20959);
xnor U27015 (N_27015,N_20759,N_18016);
nor U27016 (N_27016,N_23152,N_19656);
and U27017 (N_27017,N_22010,N_21462);
xor U27018 (N_27018,N_23012,N_22460);
and U27019 (N_27019,N_19642,N_18123);
nor U27020 (N_27020,N_18127,N_19379);
nor U27021 (N_27021,N_18923,N_19510);
nor U27022 (N_27022,N_20301,N_22967);
and U27023 (N_27023,N_20314,N_21793);
nor U27024 (N_27024,N_23014,N_19684);
nor U27025 (N_27025,N_21064,N_23448);
nand U27026 (N_27026,N_18555,N_19910);
nand U27027 (N_27027,N_23898,N_22806);
nand U27028 (N_27028,N_23008,N_23695);
or U27029 (N_27029,N_20360,N_20373);
or U27030 (N_27030,N_23914,N_21516);
or U27031 (N_27031,N_21043,N_21978);
xnor U27032 (N_27032,N_20110,N_22138);
and U27033 (N_27033,N_18500,N_20683);
xor U27034 (N_27034,N_22767,N_22165);
and U27035 (N_27035,N_21723,N_21405);
nand U27036 (N_27036,N_21959,N_20465);
xor U27037 (N_27037,N_21979,N_19422);
and U27038 (N_27038,N_19318,N_21269);
nand U27039 (N_27039,N_18874,N_22015);
and U27040 (N_27040,N_21913,N_18716);
nor U27041 (N_27041,N_23468,N_19799);
nor U27042 (N_27042,N_18045,N_18328);
and U27043 (N_27043,N_20939,N_18822);
or U27044 (N_27044,N_18133,N_21398);
xnor U27045 (N_27045,N_23559,N_20566);
or U27046 (N_27046,N_21673,N_22388);
nand U27047 (N_27047,N_21966,N_19075);
or U27048 (N_27048,N_20641,N_20998);
and U27049 (N_27049,N_22182,N_18624);
nor U27050 (N_27050,N_20744,N_20802);
or U27051 (N_27051,N_22690,N_22617);
nand U27052 (N_27052,N_19405,N_22195);
and U27053 (N_27053,N_19482,N_20479);
or U27054 (N_27054,N_20148,N_21178);
xor U27055 (N_27055,N_19332,N_20003);
nand U27056 (N_27056,N_21010,N_21709);
or U27057 (N_27057,N_19431,N_18958);
nor U27058 (N_27058,N_18222,N_20872);
nand U27059 (N_27059,N_20808,N_23141);
or U27060 (N_27060,N_23519,N_22153);
nor U27061 (N_27061,N_20098,N_20861);
nand U27062 (N_27062,N_21782,N_22083);
or U27063 (N_27063,N_22046,N_19685);
nand U27064 (N_27064,N_23557,N_19592);
nand U27065 (N_27065,N_23865,N_21050);
nor U27066 (N_27066,N_19214,N_21470);
or U27067 (N_27067,N_20469,N_21045);
and U27068 (N_27068,N_18851,N_19633);
or U27069 (N_27069,N_23333,N_20594);
nand U27070 (N_27070,N_21886,N_18800);
nor U27071 (N_27071,N_20875,N_21356);
nand U27072 (N_27072,N_20519,N_19323);
and U27073 (N_27073,N_20325,N_21090);
nor U27074 (N_27074,N_22046,N_19849);
xor U27075 (N_27075,N_18372,N_21687);
xnor U27076 (N_27076,N_23485,N_23950);
or U27077 (N_27077,N_22966,N_22125);
nor U27078 (N_27078,N_20245,N_22315);
or U27079 (N_27079,N_19197,N_21042);
or U27080 (N_27080,N_20578,N_23047);
and U27081 (N_27081,N_22836,N_23681);
nand U27082 (N_27082,N_18754,N_23271);
nor U27083 (N_27083,N_21737,N_21127);
or U27084 (N_27084,N_22731,N_20493);
nand U27085 (N_27085,N_19113,N_23479);
and U27086 (N_27086,N_18671,N_18184);
or U27087 (N_27087,N_21948,N_18270);
or U27088 (N_27088,N_21279,N_22662);
xor U27089 (N_27089,N_20398,N_19976);
and U27090 (N_27090,N_18641,N_22132);
nand U27091 (N_27091,N_23149,N_18234);
nor U27092 (N_27092,N_23220,N_23188);
nand U27093 (N_27093,N_20093,N_19781);
nand U27094 (N_27094,N_20789,N_19254);
xor U27095 (N_27095,N_22264,N_23351);
or U27096 (N_27096,N_22659,N_18080);
nor U27097 (N_27097,N_23384,N_19464);
xor U27098 (N_27098,N_22379,N_21788);
nand U27099 (N_27099,N_19386,N_21566);
or U27100 (N_27100,N_23521,N_18846);
nor U27101 (N_27101,N_23092,N_19592);
nand U27102 (N_27102,N_21939,N_21862);
and U27103 (N_27103,N_20106,N_19122);
or U27104 (N_27104,N_23566,N_23962);
nor U27105 (N_27105,N_19437,N_21870);
and U27106 (N_27106,N_18627,N_19951);
and U27107 (N_27107,N_19120,N_19856);
nor U27108 (N_27108,N_22186,N_20763);
xnor U27109 (N_27109,N_21289,N_18483);
nand U27110 (N_27110,N_23032,N_20630);
nand U27111 (N_27111,N_21156,N_22372);
nand U27112 (N_27112,N_19660,N_19549);
nor U27113 (N_27113,N_22103,N_18426);
nor U27114 (N_27114,N_23350,N_20255);
and U27115 (N_27115,N_23387,N_18752);
and U27116 (N_27116,N_22205,N_20046);
nor U27117 (N_27117,N_23959,N_22319);
or U27118 (N_27118,N_20134,N_22154);
nor U27119 (N_27119,N_18535,N_18961);
xnor U27120 (N_27120,N_21788,N_21900);
and U27121 (N_27121,N_21159,N_19342);
nand U27122 (N_27122,N_21935,N_21337);
or U27123 (N_27123,N_20182,N_18059);
nand U27124 (N_27124,N_23275,N_19494);
nor U27125 (N_27125,N_23798,N_23220);
or U27126 (N_27126,N_20212,N_18815);
nand U27127 (N_27127,N_22182,N_22993);
xnor U27128 (N_27128,N_21513,N_21855);
xor U27129 (N_27129,N_18956,N_18253);
or U27130 (N_27130,N_23007,N_19896);
xor U27131 (N_27131,N_19515,N_19959);
or U27132 (N_27132,N_19746,N_18524);
or U27133 (N_27133,N_18330,N_18788);
nand U27134 (N_27134,N_20760,N_23109);
nand U27135 (N_27135,N_22459,N_18605);
nand U27136 (N_27136,N_23137,N_23638);
or U27137 (N_27137,N_18591,N_23122);
nor U27138 (N_27138,N_21682,N_22900);
nor U27139 (N_27139,N_22873,N_23454);
xnor U27140 (N_27140,N_18160,N_19149);
or U27141 (N_27141,N_20819,N_23155);
nor U27142 (N_27142,N_18501,N_20892);
and U27143 (N_27143,N_23796,N_21164);
or U27144 (N_27144,N_22985,N_20504);
nand U27145 (N_27145,N_21253,N_20458);
nor U27146 (N_27146,N_23493,N_20461);
and U27147 (N_27147,N_23790,N_20664);
and U27148 (N_27148,N_23303,N_22626);
and U27149 (N_27149,N_19323,N_22940);
xor U27150 (N_27150,N_23996,N_21038);
nand U27151 (N_27151,N_23185,N_22656);
nor U27152 (N_27152,N_23920,N_19771);
nor U27153 (N_27153,N_21281,N_23122);
and U27154 (N_27154,N_22000,N_19186);
nand U27155 (N_27155,N_22177,N_20575);
xor U27156 (N_27156,N_21473,N_18424);
nor U27157 (N_27157,N_18298,N_19916);
nand U27158 (N_27158,N_19596,N_23089);
nand U27159 (N_27159,N_22069,N_22012);
or U27160 (N_27160,N_18297,N_23220);
nand U27161 (N_27161,N_19126,N_19646);
and U27162 (N_27162,N_21962,N_21638);
nor U27163 (N_27163,N_23081,N_18910);
and U27164 (N_27164,N_21459,N_19177);
and U27165 (N_27165,N_18973,N_20251);
and U27166 (N_27166,N_22029,N_20120);
nor U27167 (N_27167,N_23246,N_21605);
nor U27168 (N_27168,N_21145,N_21132);
nor U27169 (N_27169,N_19134,N_19775);
xnor U27170 (N_27170,N_23772,N_19501);
nand U27171 (N_27171,N_23999,N_22589);
xor U27172 (N_27172,N_21025,N_18406);
or U27173 (N_27173,N_23775,N_18689);
nand U27174 (N_27174,N_23880,N_22961);
or U27175 (N_27175,N_19697,N_23649);
or U27176 (N_27176,N_23825,N_21406);
or U27177 (N_27177,N_19061,N_23698);
nand U27178 (N_27178,N_19575,N_21392);
and U27179 (N_27179,N_23679,N_18968);
nand U27180 (N_27180,N_22165,N_22138);
nand U27181 (N_27181,N_18656,N_20229);
xor U27182 (N_27182,N_23420,N_23892);
nand U27183 (N_27183,N_23988,N_23128);
or U27184 (N_27184,N_23804,N_21282);
nand U27185 (N_27185,N_20939,N_22963);
nor U27186 (N_27186,N_21744,N_19164);
and U27187 (N_27187,N_18228,N_20938);
nor U27188 (N_27188,N_19734,N_22347);
nor U27189 (N_27189,N_18169,N_19295);
and U27190 (N_27190,N_20671,N_20728);
or U27191 (N_27191,N_21025,N_20513);
nor U27192 (N_27192,N_22855,N_18126);
nor U27193 (N_27193,N_19788,N_20835);
nor U27194 (N_27194,N_23392,N_21222);
or U27195 (N_27195,N_23467,N_18116);
xor U27196 (N_27196,N_20788,N_19433);
nor U27197 (N_27197,N_22246,N_23054);
xor U27198 (N_27198,N_18041,N_22152);
or U27199 (N_27199,N_20704,N_20563);
nor U27200 (N_27200,N_20513,N_22928);
or U27201 (N_27201,N_23887,N_20259);
and U27202 (N_27202,N_20626,N_18858);
or U27203 (N_27203,N_23635,N_20511);
or U27204 (N_27204,N_18050,N_18906);
or U27205 (N_27205,N_19356,N_23387);
and U27206 (N_27206,N_21778,N_20671);
xnor U27207 (N_27207,N_18354,N_21532);
or U27208 (N_27208,N_21565,N_21989);
or U27209 (N_27209,N_18543,N_22356);
or U27210 (N_27210,N_20748,N_23180);
and U27211 (N_27211,N_20116,N_22551);
nor U27212 (N_27212,N_20278,N_20107);
nand U27213 (N_27213,N_18291,N_20083);
nor U27214 (N_27214,N_22689,N_23798);
and U27215 (N_27215,N_18184,N_19154);
nor U27216 (N_27216,N_19980,N_23941);
and U27217 (N_27217,N_20718,N_20146);
nor U27218 (N_27218,N_18353,N_19600);
or U27219 (N_27219,N_22210,N_23947);
nand U27220 (N_27220,N_19336,N_21308);
nor U27221 (N_27221,N_23910,N_20822);
and U27222 (N_27222,N_19819,N_18114);
or U27223 (N_27223,N_18486,N_20968);
or U27224 (N_27224,N_18699,N_23553);
nand U27225 (N_27225,N_23432,N_22083);
xor U27226 (N_27226,N_20827,N_19964);
nand U27227 (N_27227,N_19794,N_23549);
or U27228 (N_27228,N_21041,N_19873);
xnor U27229 (N_27229,N_18586,N_20433);
nand U27230 (N_27230,N_21925,N_21622);
nand U27231 (N_27231,N_19458,N_20756);
and U27232 (N_27232,N_18895,N_23206);
nand U27233 (N_27233,N_20902,N_18207);
and U27234 (N_27234,N_23693,N_23653);
and U27235 (N_27235,N_20776,N_18869);
xnor U27236 (N_27236,N_20949,N_19836);
nand U27237 (N_27237,N_23616,N_20788);
nor U27238 (N_27238,N_21837,N_18148);
or U27239 (N_27239,N_20419,N_23074);
xor U27240 (N_27240,N_20864,N_21181);
xnor U27241 (N_27241,N_19528,N_19161);
and U27242 (N_27242,N_23283,N_23316);
nor U27243 (N_27243,N_23495,N_22588);
nand U27244 (N_27244,N_22087,N_19273);
nand U27245 (N_27245,N_21140,N_19803);
or U27246 (N_27246,N_19399,N_19772);
and U27247 (N_27247,N_20704,N_22669);
nor U27248 (N_27248,N_23310,N_21741);
and U27249 (N_27249,N_23322,N_23617);
nand U27250 (N_27250,N_20717,N_22522);
nor U27251 (N_27251,N_23843,N_22432);
or U27252 (N_27252,N_23449,N_18380);
nand U27253 (N_27253,N_23394,N_20547);
and U27254 (N_27254,N_22822,N_23057);
and U27255 (N_27255,N_18421,N_23651);
and U27256 (N_27256,N_23095,N_23758);
or U27257 (N_27257,N_22258,N_21478);
and U27258 (N_27258,N_21687,N_20506);
nor U27259 (N_27259,N_20266,N_21707);
nand U27260 (N_27260,N_20985,N_19612);
xor U27261 (N_27261,N_21747,N_19246);
and U27262 (N_27262,N_23977,N_22892);
nor U27263 (N_27263,N_19415,N_18610);
or U27264 (N_27264,N_22064,N_20925);
or U27265 (N_27265,N_20363,N_18025);
nor U27266 (N_27266,N_19491,N_21436);
or U27267 (N_27267,N_19129,N_19366);
xor U27268 (N_27268,N_20872,N_22207);
nand U27269 (N_27269,N_21805,N_18991);
or U27270 (N_27270,N_20388,N_19497);
or U27271 (N_27271,N_18005,N_18410);
nand U27272 (N_27272,N_18612,N_22940);
and U27273 (N_27273,N_21658,N_19978);
and U27274 (N_27274,N_18484,N_21117);
and U27275 (N_27275,N_23463,N_22524);
xnor U27276 (N_27276,N_19339,N_23970);
nor U27277 (N_27277,N_21429,N_21691);
and U27278 (N_27278,N_19884,N_19307);
or U27279 (N_27279,N_18221,N_23024);
and U27280 (N_27280,N_21170,N_20294);
nand U27281 (N_27281,N_23098,N_22639);
and U27282 (N_27282,N_18084,N_23472);
nor U27283 (N_27283,N_20401,N_20967);
nand U27284 (N_27284,N_21014,N_18354);
nand U27285 (N_27285,N_22442,N_18166);
nor U27286 (N_27286,N_20450,N_20604);
and U27287 (N_27287,N_20596,N_18682);
nand U27288 (N_27288,N_18330,N_20788);
or U27289 (N_27289,N_19515,N_22907);
nand U27290 (N_27290,N_23504,N_18343);
and U27291 (N_27291,N_22586,N_18908);
nand U27292 (N_27292,N_23605,N_19952);
xnor U27293 (N_27293,N_23891,N_21367);
or U27294 (N_27294,N_22106,N_23164);
nor U27295 (N_27295,N_22141,N_20823);
nor U27296 (N_27296,N_20755,N_20311);
nor U27297 (N_27297,N_19098,N_20929);
and U27298 (N_27298,N_20026,N_23078);
and U27299 (N_27299,N_23707,N_23279);
nand U27300 (N_27300,N_19992,N_23021);
nor U27301 (N_27301,N_18878,N_21722);
and U27302 (N_27302,N_23853,N_23368);
and U27303 (N_27303,N_20739,N_23098);
nor U27304 (N_27304,N_23321,N_23942);
and U27305 (N_27305,N_19047,N_21063);
or U27306 (N_27306,N_23805,N_20745);
nand U27307 (N_27307,N_22501,N_22416);
or U27308 (N_27308,N_20260,N_23446);
xnor U27309 (N_27309,N_23570,N_18643);
or U27310 (N_27310,N_22529,N_20169);
nor U27311 (N_27311,N_18694,N_18184);
xnor U27312 (N_27312,N_19607,N_19429);
nand U27313 (N_27313,N_19605,N_23473);
xnor U27314 (N_27314,N_22808,N_21825);
or U27315 (N_27315,N_21893,N_23288);
nor U27316 (N_27316,N_20071,N_19621);
and U27317 (N_27317,N_20517,N_23006);
nor U27318 (N_27318,N_23691,N_22063);
and U27319 (N_27319,N_19464,N_18614);
or U27320 (N_27320,N_21277,N_19128);
xor U27321 (N_27321,N_20674,N_21223);
nor U27322 (N_27322,N_18392,N_22895);
and U27323 (N_27323,N_18801,N_23400);
and U27324 (N_27324,N_21772,N_22813);
nand U27325 (N_27325,N_18318,N_21181);
and U27326 (N_27326,N_22789,N_19620);
and U27327 (N_27327,N_21751,N_18112);
xor U27328 (N_27328,N_19813,N_18338);
nor U27329 (N_27329,N_22776,N_20404);
and U27330 (N_27330,N_18583,N_18513);
nand U27331 (N_27331,N_21466,N_20757);
xnor U27332 (N_27332,N_23374,N_19340);
nand U27333 (N_27333,N_21826,N_19449);
xor U27334 (N_27334,N_22953,N_18454);
xnor U27335 (N_27335,N_23693,N_18163);
or U27336 (N_27336,N_19023,N_23391);
or U27337 (N_27337,N_23931,N_19809);
and U27338 (N_27338,N_21750,N_21267);
or U27339 (N_27339,N_20902,N_18615);
nand U27340 (N_27340,N_22278,N_21769);
xnor U27341 (N_27341,N_20766,N_22961);
nand U27342 (N_27342,N_22353,N_18631);
and U27343 (N_27343,N_19114,N_19161);
nor U27344 (N_27344,N_19624,N_21198);
nand U27345 (N_27345,N_18867,N_23676);
nor U27346 (N_27346,N_22469,N_19987);
nor U27347 (N_27347,N_18542,N_20282);
nand U27348 (N_27348,N_20114,N_22533);
nor U27349 (N_27349,N_21135,N_22031);
xnor U27350 (N_27350,N_18093,N_18478);
nor U27351 (N_27351,N_19925,N_20564);
and U27352 (N_27352,N_19718,N_19627);
nand U27353 (N_27353,N_22965,N_22646);
nor U27354 (N_27354,N_19419,N_23606);
nor U27355 (N_27355,N_18777,N_19774);
or U27356 (N_27356,N_21544,N_20900);
or U27357 (N_27357,N_20936,N_22505);
or U27358 (N_27358,N_19213,N_23393);
xnor U27359 (N_27359,N_18464,N_20790);
nor U27360 (N_27360,N_21903,N_23523);
and U27361 (N_27361,N_21924,N_22334);
or U27362 (N_27362,N_20385,N_21600);
nor U27363 (N_27363,N_23119,N_23494);
xnor U27364 (N_27364,N_21542,N_20998);
nand U27365 (N_27365,N_19283,N_18706);
or U27366 (N_27366,N_20694,N_19933);
nand U27367 (N_27367,N_19344,N_18717);
xor U27368 (N_27368,N_20506,N_18277);
nor U27369 (N_27369,N_23061,N_19913);
nand U27370 (N_27370,N_23778,N_21575);
nor U27371 (N_27371,N_20137,N_21801);
or U27372 (N_27372,N_20130,N_23614);
or U27373 (N_27373,N_20505,N_18480);
nand U27374 (N_27374,N_22489,N_23156);
nor U27375 (N_27375,N_21808,N_22242);
or U27376 (N_27376,N_21280,N_18809);
and U27377 (N_27377,N_18913,N_18938);
and U27378 (N_27378,N_23302,N_22175);
or U27379 (N_27379,N_23522,N_18120);
and U27380 (N_27380,N_18529,N_21382);
nor U27381 (N_27381,N_19432,N_18897);
or U27382 (N_27382,N_18171,N_20365);
nor U27383 (N_27383,N_23159,N_19156);
nor U27384 (N_27384,N_23588,N_23434);
nand U27385 (N_27385,N_22781,N_23477);
nand U27386 (N_27386,N_21531,N_20649);
nor U27387 (N_27387,N_21587,N_23148);
and U27388 (N_27388,N_20428,N_23598);
nor U27389 (N_27389,N_23227,N_22596);
and U27390 (N_27390,N_21879,N_18555);
or U27391 (N_27391,N_22397,N_23700);
nor U27392 (N_27392,N_22641,N_23094);
xnor U27393 (N_27393,N_20972,N_19548);
or U27394 (N_27394,N_18151,N_18895);
nor U27395 (N_27395,N_20927,N_23619);
nand U27396 (N_27396,N_22684,N_23624);
nor U27397 (N_27397,N_20175,N_19962);
or U27398 (N_27398,N_22952,N_19022);
or U27399 (N_27399,N_20840,N_23289);
nor U27400 (N_27400,N_19306,N_20855);
nand U27401 (N_27401,N_22706,N_21399);
nor U27402 (N_27402,N_20314,N_21323);
and U27403 (N_27403,N_20280,N_23537);
xnor U27404 (N_27404,N_21861,N_22013);
nor U27405 (N_27405,N_21992,N_21410);
and U27406 (N_27406,N_22666,N_20842);
nor U27407 (N_27407,N_19129,N_20619);
and U27408 (N_27408,N_18371,N_20317);
and U27409 (N_27409,N_22959,N_20367);
or U27410 (N_27410,N_21324,N_19965);
xnor U27411 (N_27411,N_23741,N_20621);
nand U27412 (N_27412,N_20760,N_20702);
nand U27413 (N_27413,N_19487,N_18310);
or U27414 (N_27414,N_23875,N_23125);
nor U27415 (N_27415,N_20456,N_20759);
or U27416 (N_27416,N_23116,N_18925);
or U27417 (N_27417,N_23187,N_22158);
nand U27418 (N_27418,N_18045,N_23467);
and U27419 (N_27419,N_21234,N_19719);
and U27420 (N_27420,N_22412,N_23380);
nand U27421 (N_27421,N_21729,N_22642);
xnor U27422 (N_27422,N_21233,N_21953);
nand U27423 (N_27423,N_22229,N_20856);
or U27424 (N_27424,N_22940,N_20026);
nand U27425 (N_27425,N_19564,N_23439);
nand U27426 (N_27426,N_23153,N_18384);
nor U27427 (N_27427,N_23512,N_22028);
nor U27428 (N_27428,N_19863,N_23234);
nor U27429 (N_27429,N_20433,N_19857);
nor U27430 (N_27430,N_20775,N_23000);
xnor U27431 (N_27431,N_19134,N_22019);
or U27432 (N_27432,N_23717,N_20904);
nand U27433 (N_27433,N_22351,N_18967);
nor U27434 (N_27434,N_21954,N_20699);
or U27435 (N_27435,N_21742,N_20150);
and U27436 (N_27436,N_22925,N_18608);
and U27437 (N_27437,N_23288,N_20449);
nor U27438 (N_27438,N_18442,N_21978);
and U27439 (N_27439,N_22998,N_20187);
or U27440 (N_27440,N_22952,N_21430);
or U27441 (N_27441,N_20349,N_22236);
nor U27442 (N_27442,N_19126,N_18910);
and U27443 (N_27443,N_20992,N_22793);
or U27444 (N_27444,N_21141,N_19469);
nand U27445 (N_27445,N_20720,N_22518);
or U27446 (N_27446,N_21937,N_18475);
nor U27447 (N_27447,N_22722,N_18312);
nand U27448 (N_27448,N_18036,N_19478);
and U27449 (N_27449,N_21340,N_23661);
nand U27450 (N_27450,N_18307,N_22216);
or U27451 (N_27451,N_19944,N_22577);
nand U27452 (N_27452,N_18587,N_23627);
nor U27453 (N_27453,N_20035,N_22659);
nand U27454 (N_27454,N_19027,N_19558);
nand U27455 (N_27455,N_23157,N_18392);
nand U27456 (N_27456,N_18209,N_21470);
nor U27457 (N_27457,N_18161,N_19452);
or U27458 (N_27458,N_22485,N_23107);
or U27459 (N_27459,N_19936,N_18122);
xor U27460 (N_27460,N_22414,N_19628);
or U27461 (N_27461,N_23029,N_21385);
and U27462 (N_27462,N_18687,N_22254);
nor U27463 (N_27463,N_18297,N_18786);
and U27464 (N_27464,N_20713,N_18767);
or U27465 (N_27465,N_23678,N_21969);
nor U27466 (N_27466,N_19615,N_18792);
or U27467 (N_27467,N_18202,N_22891);
nor U27468 (N_27468,N_22112,N_22166);
and U27469 (N_27469,N_22225,N_21373);
nor U27470 (N_27470,N_21388,N_19059);
or U27471 (N_27471,N_22272,N_19871);
nor U27472 (N_27472,N_22762,N_23899);
and U27473 (N_27473,N_23478,N_19625);
nor U27474 (N_27474,N_19351,N_23579);
nor U27475 (N_27475,N_18199,N_20126);
xnor U27476 (N_27476,N_19862,N_20069);
nand U27477 (N_27477,N_18987,N_19720);
or U27478 (N_27478,N_20170,N_21073);
nand U27479 (N_27479,N_23619,N_18193);
nand U27480 (N_27480,N_20147,N_22848);
nor U27481 (N_27481,N_22369,N_21264);
and U27482 (N_27482,N_22963,N_19041);
or U27483 (N_27483,N_23749,N_19287);
nand U27484 (N_27484,N_20969,N_18096);
nand U27485 (N_27485,N_18553,N_18124);
or U27486 (N_27486,N_20729,N_19119);
or U27487 (N_27487,N_21591,N_21133);
or U27488 (N_27488,N_19486,N_19750);
and U27489 (N_27489,N_21328,N_21280);
and U27490 (N_27490,N_18537,N_22322);
and U27491 (N_27491,N_22653,N_18801);
nor U27492 (N_27492,N_22392,N_22127);
nor U27493 (N_27493,N_22542,N_23645);
and U27494 (N_27494,N_19671,N_19128);
xnor U27495 (N_27495,N_22526,N_21347);
nor U27496 (N_27496,N_23704,N_23722);
and U27497 (N_27497,N_18793,N_22496);
or U27498 (N_27498,N_23547,N_19896);
xor U27499 (N_27499,N_21258,N_22411);
nand U27500 (N_27500,N_20316,N_23222);
or U27501 (N_27501,N_20988,N_23225);
nor U27502 (N_27502,N_19814,N_19035);
or U27503 (N_27503,N_20990,N_18091);
nor U27504 (N_27504,N_20496,N_21985);
or U27505 (N_27505,N_23821,N_18544);
and U27506 (N_27506,N_20158,N_19539);
nor U27507 (N_27507,N_22285,N_18024);
and U27508 (N_27508,N_19685,N_22463);
nor U27509 (N_27509,N_23428,N_19263);
xnor U27510 (N_27510,N_18930,N_23709);
nor U27511 (N_27511,N_18536,N_23641);
nand U27512 (N_27512,N_21260,N_20243);
or U27513 (N_27513,N_18825,N_18706);
or U27514 (N_27514,N_23897,N_19271);
and U27515 (N_27515,N_19433,N_18764);
or U27516 (N_27516,N_19905,N_21888);
nor U27517 (N_27517,N_20435,N_22025);
nand U27518 (N_27518,N_18952,N_20030);
nand U27519 (N_27519,N_18699,N_18529);
and U27520 (N_27520,N_23982,N_22854);
xor U27521 (N_27521,N_23950,N_19863);
nand U27522 (N_27522,N_22280,N_20638);
or U27523 (N_27523,N_20397,N_21174);
nor U27524 (N_27524,N_18700,N_19610);
nand U27525 (N_27525,N_19123,N_18698);
nor U27526 (N_27526,N_19933,N_20683);
or U27527 (N_27527,N_18661,N_23913);
nor U27528 (N_27528,N_19999,N_20457);
and U27529 (N_27529,N_23702,N_20806);
nor U27530 (N_27530,N_23948,N_22548);
nor U27531 (N_27531,N_18130,N_21050);
nand U27532 (N_27532,N_19723,N_20893);
and U27533 (N_27533,N_20656,N_18270);
and U27534 (N_27534,N_20343,N_23170);
and U27535 (N_27535,N_18903,N_20220);
or U27536 (N_27536,N_21258,N_23170);
or U27537 (N_27537,N_20685,N_20469);
and U27538 (N_27538,N_19593,N_19341);
and U27539 (N_27539,N_23455,N_20757);
xor U27540 (N_27540,N_21047,N_21594);
nor U27541 (N_27541,N_19308,N_20315);
xnor U27542 (N_27542,N_22195,N_20964);
nor U27543 (N_27543,N_19454,N_18229);
nor U27544 (N_27544,N_22471,N_21010);
nor U27545 (N_27545,N_21307,N_21989);
nand U27546 (N_27546,N_19062,N_23460);
nand U27547 (N_27547,N_22301,N_20226);
nand U27548 (N_27548,N_21277,N_18351);
nand U27549 (N_27549,N_20399,N_23322);
or U27550 (N_27550,N_22865,N_19944);
nand U27551 (N_27551,N_22828,N_19919);
and U27552 (N_27552,N_21845,N_22806);
or U27553 (N_27553,N_20305,N_22817);
nor U27554 (N_27554,N_21526,N_18612);
nand U27555 (N_27555,N_23414,N_22546);
and U27556 (N_27556,N_21359,N_19811);
nor U27557 (N_27557,N_18214,N_22331);
nor U27558 (N_27558,N_21524,N_23377);
and U27559 (N_27559,N_20978,N_22178);
or U27560 (N_27560,N_18487,N_22563);
nor U27561 (N_27561,N_22287,N_18135);
nor U27562 (N_27562,N_20241,N_22512);
nor U27563 (N_27563,N_19981,N_18206);
nor U27564 (N_27564,N_20412,N_21542);
nor U27565 (N_27565,N_22669,N_21821);
and U27566 (N_27566,N_22746,N_21595);
nand U27567 (N_27567,N_21089,N_19057);
nor U27568 (N_27568,N_20588,N_22987);
or U27569 (N_27569,N_18280,N_22676);
nand U27570 (N_27570,N_20940,N_21311);
nand U27571 (N_27571,N_18782,N_18596);
nand U27572 (N_27572,N_19471,N_22980);
or U27573 (N_27573,N_23184,N_23314);
or U27574 (N_27574,N_21497,N_21670);
nor U27575 (N_27575,N_18592,N_18741);
or U27576 (N_27576,N_20668,N_20780);
or U27577 (N_27577,N_23660,N_18970);
nor U27578 (N_27578,N_19290,N_20287);
nand U27579 (N_27579,N_22622,N_18395);
and U27580 (N_27580,N_19281,N_22922);
nand U27581 (N_27581,N_19417,N_23490);
xnor U27582 (N_27582,N_22043,N_19807);
nand U27583 (N_27583,N_21500,N_19578);
or U27584 (N_27584,N_22149,N_19057);
or U27585 (N_27585,N_22824,N_21335);
or U27586 (N_27586,N_18923,N_23783);
or U27587 (N_27587,N_20378,N_21628);
and U27588 (N_27588,N_23373,N_21257);
and U27589 (N_27589,N_21144,N_22896);
and U27590 (N_27590,N_20617,N_21524);
or U27591 (N_27591,N_22920,N_22396);
nand U27592 (N_27592,N_18747,N_22755);
and U27593 (N_27593,N_19444,N_22858);
nor U27594 (N_27594,N_19357,N_22979);
nor U27595 (N_27595,N_19202,N_22936);
nor U27596 (N_27596,N_22524,N_18422);
or U27597 (N_27597,N_19775,N_23802);
nor U27598 (N_27598,N_20158,N_21481);
and U27599 (N_27599,N_22435,N_23437);
and U27600 (N_27600,N_18667,N_22698);
or U27601 (N_27601,N_22343,N_18150);
or U27602 (N_27602,N_20168,N_22843);
or U27603 (N_27603,N_19510,N_19572);
and U27604 (N_27604,N_19131,N_19486);
and U27605 (N_27605,N_20547,N_20920);
nor U27606 (N_27606,N_18279,N_19984);
or U27607 (N_27607,N_18191,N_22492);
nor U27608 (N_27608,N_21583,N_23275);
nand U27609 (N_27609,N_20670,N_23585);
or U27610 (N_27610,N_21725,N_20176);
nor U27611 (N_27611,N_23644,N_18055);
or U27612 (N_27612,N_18929,N_23232);
and U27613 (N_27613,N_19681,N_23498);
nor U27614 (N_27614,N_22025,N_21571);
nor U27615 (N_27615,N_20146,N_18658);
nand U27616 (N_27616,N_20592,N_22906);
and U27617 (N_27617,N_20795,N_18736);
nor U27618 (N_27618,N_21038,N_22426);
or U27619 (N_27619,N_20202,N_21441);
nor U27620 (N_27620,N_22653,N_21714);
and U27621 (N_27621,N_18338,N_22908);
nor U27622 (N_27622,N_18684,N_21022);
nor U27623 (N_27623,N_23899,N_18875);
nor U27624 (N_27624,N_18200,N_19618);
or U27625 (N_27625,N_21033,N_23873);
nor U27626 (N_27626,N_21764,N_22784);
nand U27627 (N_27627,N_20628,N_20192);
and U27628 (N_27628,N_21142,N_20597);
or U27629 (N_27629,N_20345,N_23562);
or U27630 (N_27630,N_19322,N_23311);
nand U27631 (N_27631,N_19901,N_18924);
or U27632 (N_27632,N_22165,N_21813);
or U27633 (N_27633,N_22333,N_22112);
xor U27634 (N_27634,N_22271,N_20507);
or U27635 (N_27635,N_22350,N_20163);
and U27636 (N_27636,N_18523,N_21609);
nand U27637 (N_27637,N_20803,N_23806);
or U27638 (N_27638,N_20354,N_23171);
and U27639 (N_27639,N_21983,N_18016);
nor U27640 (N_27640,N_20577,N_18248);
and U27641 (N_27641,N_18962,N_21527);
nand U27642 (N_27642,N_21117,N_21346);
nor U27643 (N_27643,N_23305,N_18909);
and U27644 (N_27644,N_21868,N_18754);
nand U27645 (N_27645,N_22023,N_23954);
nor U27646 (N_27646,N_23483,N_23884);
and U27647 (N_27647,N_22604,N_20711);
or U27648 (N_27648,N_19190,N_19034);
nor U27649 (N_27649,N_22071,N_19216);
or U27650 (N_27650,N_18431,N_23722);
nor U27651 (N_27651,N_19891,N_21227);
nor U27652 (N_27652,N_21105,N_22472);
or U27653 (N_27653,N_21149,N_19248);
or U27654 (N_27654,N_23304,N_19149);
and U27655 (N_27655,N_23416,N_22707);
and U27656 (N_27656,N_20757,N_19660);
and U27657 (N_27657,N_20084,N_22434);
and U27658 (N_27658,N_20166,N_18894);
nand U27659 (N_27659,N_19593,N_23524);
or U27660 (N_27660,N_18265,N_19478);
nand U27661 (N_27661,N_20651,N_22184);
and U27662 (N_27662,N_20661,N_20084);
and U27663 (N_27663,N_20335,N_22039);
nor U27664 (N_27664,N_22729,N_20572);
and U27665 (N_27665,N_18761,N_19919);
nand U27666 (N_27666,N_19573,N_21942);
nor U27667 (N_27667,N_20287,N_18804);
or U27668 (N_27668,N_23082,N_18121);
or U27669 (N_27669,N_19681,N_21738);
xnor U27670 (N_27670,N_19329,N_22814);
or U27671 (N_27671,N_20637,N_18558);
nand U27672 (N_27672,N_18642,N_19433);
and U27673 (N_27673,N_20622,N_20916);
or U27674 (N_27674,N_23639,N_20480);
nand U27675 (N_27675,N_18887,N_18546);
xor U27676 (N_27676,N_22738,N_19444);
or U27677 (N_27677,N_19141,N_21367);
or U27678 (N_27678,N_21690,N_21021);
nor U27679 (N_27679,N_20894,N_21625);
nor U27680 (N_27680,N_23671,N_19392);
nor U27681 (N_27681,N_20940,N_20886);
nand U27682 (N_27682,N_22260,N_22727);
nand U27683 (N_27683,N_19005,N_19649);
nand U27684 (N_27684,N_21791,N_21627);
nor U27685 (N_27685,N_18236,N_23719);
and U27686 (N_27686,N_21853,N_20174);
and U27687 (N_27687,N_22830,N_20476);
or U27688 (N_27688,N_19383,N_20039);
and U27689 (N_27689,N_22685,N_23002);
and U27690 (N_27690,N_20224,N_21837);
nand U27691 (N_27691,N_18311,N_20343);
xor U27692 (N_27692,N_22877,N_18902);
and U27693 (N_27693,N_18536,N_20714);
xnor U27694 (N_27694,N_21480,N_21906);
and U27695 (N_27695,N_22887,N_23283);
and U27696 (N_27696,N_20947,N_21880);
nor U27697 (N_27697,N_20568,N_18068);
and U27698 (N_27698,N_21418,N_21495);
nor U27699 (N_27699,N_19816,N_18409);
nand U27700 (N_27700,N_18792,N_21064);
and U27701 (N_27701,N_22065,N_19433);
nand U27702 (N_27702,N_19085,N_20142);
or U27703 (N_27703,N_18240,N_18058);
or U27704 (N_27704,N_23283,N_22376);
and U27705 (N_27705,N_18085,N_21764);
and U27706 (N_27706,N_23615,N_18681);
and U27707 (N_27707,N_21422,N_21845);
nor U27708 (N_27708,N_18242,N_21269);
nand U27709 (N_27709,N_22289,N_21183);
or U27710 (N_27710,N_22743,N_18447);
nand U27711 (N_27711,N_19603,N_20124);
and U27712 (N_27712,N_23711,N_19207);
or U27713 (N_27713,N_21340,N_18694);
or U27714 (N_27714,N_19661,N_18996);
nor U27715 (N_27715,N_20238,N_21288);
or U27716 (N_27716,N_22472,N_20057);
nor U27717 (N_27717,N_19397,N_21717);
xnor U27718 (N_27718,N_20669,N_22425);
nor U27719 (N_27719,N_18669,N_21807);
or U27720 (N_27720,N_23349,N_18958);
and U27721 (N_27721,N_23953,N_23805);
or U27722 (N_27722,N_18418,N_19904);
and U27723 (N_27723,N_22732,N_21433);
or U27724 (N_27724,N_18668,N_21127);
or U27725 (N_27725,N_19816,N_21520);
xnor U27726 (N_27726,N_19854,N_19043);
xor U27727 (N_27727,N_21798,N_20224);
nor U27728 (N_27728,N_22591,N_18457);
and U27729 (N_27729,N_22448,N_19349);
nor U27730 (N_27730,N_22500,N_23285);
and U27731 (N_27731,N_23319,N_19471);
or U27732 (N_27732,N_19380,N_22853);
or U27733 (N_27733,N_19870,N_20761);
nand U27734 (N_27734,N_23971,N_23979);
nor U27735 (N_27735,N_21229,N_19812);
nor U27736 (N_27736,N_22372,N_18405);
nor U27737 (N_27737,N_19989,N_23893);
nand U27738 (N_27738,N_20099,N_21455);
and U27739 (N_27739,N_23392,N_19738);
nor U27740 (N_27740,N_20542,N_21946);
or U27741 (N_27741,N_23665,N_22378);
and U27742 (N_27742,N_19280,N_23974);
nand U27743 (N_27743,N_21606,N_21582);
nand U27744 (N_27744,N_22347,N_21278);
nor U27745 (N_27745,N_21809,N_21417);
nor U27746 (N_27746,N_22169,N_23904);
and U27747 (N_27747,N_20191,N_19405);
or U27748 (N_27748,N_21628,N_23767);
and U27749 (N_27749,N_18658,N_22113);
nand U27750 (N_27750,N_19542,N_23476);
and U27751 (N_27751,N_21080,N_23566);
nor U27752 (N_27752,N_18255,N_18936);
nand U27753 (N_27753,N_22983,N_20021);
nor U27754 (N_27754,N_23125,N_21145);
xor U27755 (N_27755,N_19892,N_18445);
xnor U27756 (N_27756,N_20988,N_20458);
nor U27757 (N_27757,N_20888,N_20919);
or U27758 (N_27758,N_21144,N_22719);
nor U27759 (N_27759,N_21223,N_22323);
and U27760 (N_27760,N_20139,N_19683);
and U27761 (N_27761,N_23444,N_22487);
and U27762 (N_27762,N_20155,N_20975);
and U27763 (N_27763,N_19467,N_23553);
nand U27764 (N_27764,N_22696,N_22398);
xor U27765 (N_27765,N_18667,N_22741);
or U27766 (N_27766,N_22500,N_19154);
or U27767 (N_27767,N_18145,N_21431);
or U27768 (N_27768,N_18770,N_18334);
nor U27769 (N_27769,N_20204,N_20788);
xnor U27770 (N_27770,N_21840,N_22068);
nor U27771 (N_27771,N_19865,N_20783);
xnor U27772 (N_27772,N_21251,N_20089);
xor U27773 (N_27773,N_18879,N_23625);
nand U27774 (N_27774,N_20245,N_23259);
or U27775 (N_27775,N_19476,N_20753);
or U27776 (N_27776,N_21796,N_20461);
xnor U27777 (N_27777,N_22755,N_18654);
xnor U27778 (N_27778,N_23082,N_22449);
nor U27779 (N_27779,N_20623,N_19547);
nor U27780 (N_27780,N_20392,N_21254);
nand U27781 (N_27781,N_18320,N_23173);
or U27782 (N_27782,N_23039,N_18150);
and U27783 (N_27783,N_22296,N_21625);
xnor U27784 (N_27784,N_22644,N_22416);
or U27785 (N_27785,N_18887,N_19255);
or U27786 (N_27786,N_22486,N_20337);
nand U27787 (N_27787,N_20965,N_19324);
or U27788 (N_27788,N_20358,N_22269);
or U27789 (N_27789,N_20237,N_19936);
and U27790 (N_27790,N_19607,N_22426);
nand U27791 (N_27791,N_21895,N_20631);
or U27792 (N_27792,N_23721,N_20982);
and U27793 (N_27793,N_22021,N_18034);
and U27794 (N_27794,N_21071,N_21022);
and U27795 (N_27795,N_19780,N_19144);
and U27796 (N_27796,N_20312,N_18462);
nor U27797 (N_27797,N_20952,N_22028);
or U27798 (N_27798,N_20336,N_22756);
and U27799 (N_27799,N_20658,N_21665);
or U27800 (N_27800,N_20552,N_21120);
xor U27801 (N_27801,N_18869,N_23128);
nand U27802 (N_27802,N_18609,N_23911);
nor U27803 (N_27803,N_20561,N_21717);
nor U27804 (N_27804,N_18085,N_18048);
nor U27805 (N_27805,N_19988,N_19031);
and U27806 (N_27806,N_22601,N_20445);
nor U27807 (N_27807,N_21152,N_19541);
nand U27808 (N_27808,N_18255,N_21991);
and U27809 (N_27809,N_21896,N_23961);
nand U27810 (N_27810,N_20433,N_18833);
or U27811 (N_27811,N_21299,N_19163);
and U27812 (N_27812,N_19470,N_19602);
nand U27813 (N_27813,N_22784,N_20729);
or U27814 (N_27814,N_20629,N_18993);
xor U27815 (N_27815,N_22932,N_18780);
nor U27816 (N_27816,N_19318,N_23999);
nor U27817 (N_27817,N_20422,N_18677);
or U27818 (N_27818,N_19464,N_20806);
nand U27819 (N_27819,N_19828,N_23022);
and U27820 (N_27820,N_22773,N_22734);
nand U27821 (N_27821,N_22606,N_20831);
nor U27822 (N_27822,N_21072,N_22225);
nor U27823 (N_27823,N_20857,N_20101);
nand U27824 (N_27824,N_23886,N_23419);
xor U27825 (N_27825,N_19513,N_18527);
and U27826 (N_27826,N_19374,N_19948);
nand U27827 (N_27827,N_20570,N_21995);
nor U27828 (N_27828,N_22548,N_18516);
or U27829 (N_27829,N_20380,N_21160);
xor U27830 (N_27830,N_21673,N_18491);
or U27831 (N_27831,N_22961,N_23030);
and U27832 (N_27832,N_23180,N_23702);
or U27833 (N_27833,N_19522,N_19035);
nor U27834 (N_27834,N_18182,N_20402);
or U27835 (N_27835,N_22173,N_20233);
and U27836 (N_27836,N_21929,N_18268);
xnor U27837 (N_27837,N_21323,N_22767);
or U27838 (N_27838,N_20923,N_19861);
nor U27839 (N_27839,N_19646,N_19989);
xnor U27840 (N_27840,N_18713,N_21329);
or U27841 (N_27841,N_23553,N_22454);
nor U27842 (N_27842,N_18370,N_19962);
and U27843 (N_27843,N_21371,N_19954);
or U27844 (N_27844,N_22208,N_23803);
nor U27845 (N_27845,N_22829,N_20324);
xor U27846 (N_27846,N_21335,N_18516);
and U27847 (N_27847,N_18896,N_22867);
and U27848 (N_27848,N_20038,N_18029);
nor U27849 (N_27849,N_22259,N_20671);
or U27850 (N_27850,N_20729,N_18322);
and U27851 (N_27851,N_19342,N_21576);
or U27852 (N_27852,N_23693,N_21722);
xnor U27853 (N_27853,N_18109,N_18250);
nor U27854 (N_27854,N_19611,N_18776);
or U27855 (N_27855,N_23556,N_22734);
xnor U27856 (N_27856,N_18884,N_22892);
nand U27857 (N_27857,N_19255,N_23686);
nand U27858 (N_27858,N_19024,N_21910);
or U27859 (N_27859,N_23795,N_23903);
and U27860 (N_27860,N_23097,N_18532);
and U27861 (N_27861,N_21592,N_18708);
or U27862 (N_27862,N_20970,N_23917);
nand U27863 (N_27863,N_20044,N_20623);
and U27864 (N_27864,N_22276,N_22745);
nor U27865 (N_27865,N_20584,N_23401);
and U27866 (N_27866,N_20808,N_20017);
and U27867 (N_27867,N_19230,N_20715);
nor U27868 (N_27868,N_22834,N_21100);
or U27869 (N_27869,N_19319,N_21065);
and U27870 (N_27870,N_18443,N_21890);
xnor U27871 (N_27871,N_20173,N_22760);
or U27872 (N_27872,N_20588,N_20448);
nor U27873 (N_27873,N_22417,N_18500);
and U27874 (N_27874,N_22211,N_22261);
or U27875 (N_27875,N_20138,N_23154);
nor U27876 (N_27876,N_22794,N_22712);
nor U27877 (N_27877,N_23971,N_22532);
nand U27878 (N_27878,N_22127,N_23440);
or U27879 (N_27879,N_22409,N_23874);
nor U27880 (N_27880,N_21436,N_20314);
or U27881 (N_27881,N_20393,N_22274);
nor U27882 (N_27882,N_23252,N_21326);
nor U27883 (N_27883,N_21677,N_23716);
and U27884 (N_27884,N_19289,N_23157);
nor U27885 (N_27885,N_20281,N_23188);
or U27886 (N_27886,N_21067,N_19963);
nand U27887 (N_27887,N_18830,N_18201);
nand U27888 (N_27888,N_21004,N_20860);
nand U27889 (N_27889,N_21528,N_22975);
and U27890 (N_27890,N_21050,N_22055);
nor U27891 (N_27891,N_21112,N_19424);
and U27892 (N_27892,N_22800,N_19525);
and U27893 (N_27893,N_20942,N_20626);
and U27894 (N_27894,N_22299,N_21943);
nand U27895 (N_27895,N_20199,N_18208);
or U27896 (N_27896,N_19425,N_19247);
or U27897 (N_27897,N_20806,N_23596);
nand U27898 (N_27898,N_20810,N_18336);
nor U27899 (N_27899,N_21912,N_19525);
nor U27900 (N_27900,N_23995,N_22866);
nor U27901 (N_27901,N_18978,N_19930);
nor U27902 (N_27902,N_20745,N_21121);
nor U27903 (N_27903,N_20512,N_22722);
nand U27904 (N_27904,N_19358,N_19173);
nand U27905 (N_27905,N_23521,N_18924);
nor U27906 (N_27906,N_21317,N_23840);
or U27907 (N_27907,N_23484,N_21027);
nand U27908 (N_27908,N_23242,N_18628);
or U27909 (N_27909,N_22071,N_21948);
or U27910 (N_27910,N_21686,N_19702);
or U27911 (N_27911,N_18983,N_23196);
xnor U27912 (N_27912,N_22517,N_20654);
or U27913 (N_27913,N_22339,N_20805);
xor U27914 (N_27914,N_21376,N_21660);
and U27915 (N_27915,N_19529,N_20547);
or U27916 (N_27916,N_22267,N_18245);
and U27917 (N_27917,N_23336,N_19864);
nand U27918 (N_27918,N_22683,N_20910);
nand U27919 (N_27919,N_18481,N_22043);
nor U27920 (N_27920,N_19572,N_20444);
nor U27921 (N_27921,N_18439,N_18837);
or U27922 (N_27922,N_18824,N_18765);
nor U27923 (N_27923,N_20317,N_21356);
and U27924 (N_27924,N_18501,N_23525);
xor U27925 (N_27925,N_19433,N_18857);
and U27926 (N_27926,N_18886,N_23176);
and U27927 (N_27927,N_20441,N_22280);
nand U27928 (N_27928,N_18949,N_23973);
and U27929 (N_27929,N_21029,N_20276);
nand U27930 (N_27930,N_20224,N_21648);
nor U27931 (N_27931,N_20872,N_20634);
nand U27932 (N_27932,N_19058,N_20053);
nand U27933 (N_27933,N_23248,N_21616);
nor U27934 (N_27934,N_23112,N_21818);
or U27935 (N_27935,N_19202,N_21930);
or U27936 (N_27936,N_19983,N_23410);
and U27937 (N_27937,N_18245,N_18579);
xnor U27938 (N_27938,N_19456,N_18809);
and U27939 (N_27939,N_18210,N_18544);
nor U27940 (N_27940,N_22537,N_23437);
and U27941 (N_27941,N_19654,N_18002);
nor U27942 (N_27942,N_19962,N_20605);
or U27943 (N_27943,N_18100,N_18857);
and U27944 (N_27944,N_20417,N_20307);
and U27945 (N_27945,N_19987,N_21489);
xnor U27946 (N_27946,N_20822,N_21716);
or U27947 (N_27947,N_20374,N_23179);
and U27948 (N_27948,N_21594,N_18785);
nor U27949 (N_27949,N_22567,N_19319);
or U27950 (N_27950,N_21158,N_18138);
xor U27951 (N_27951,N_19607,N_21108);
and U27952 (N_27952,N_21314,N_22262);
nor U27953 (N_27953,N_22242,N_19969);
nand U27954 (N_27954,N_19609,N_20531);
or U27955 (N_27955,N_23783,N_21910);
and U27956 (N_27956,N_18830,N_21246);
or U27957 (N_27957,N_18412,N_19512);
xnor U27958 (N_27958,N_21902,N_23851);
nand U27959 (N_27959,N_19630,N_20759);
and U27960 (N_27960,N_19273,N_22430);
nand U27961 (N_27961,N_19379,N_19445);
nor U27962 (N_27962,N_18008,N_19081);
nor U27963 (N_27963,N_20110,N_19403);
or U27964 (N_27964,N_21428,N_18656);
nand U27965 (N_27965,N_22073,N_23451);
xor U27966 (N_27966,N_20098,N_23163);
or U27967 (N_27967,N_18624,N_23546);
or U27968 (N_27968,N_20146,N_22830);
nand U27969 (N_27969,N_19254,N_23148);
or U27970 (N_27970,N_19338,N_18042);
nand U27971 (N_27971,N_23157,N_20414);
or U27972 (N_27972,N_18275,N_22220);
nor U27973 (N_27973,N_19177,N_20671);
or U27974 (N_27974,N_18494,N_22999);
nand U27975 (N_27975,N_18418,N_18869);
nand U27976 (N_27976,N_20509,N_21573);
nand U27977 (N_27977,N_23408,N_22029);
or U27978 (N_27978,N_22147,N_19779);
or U27979 (N_27979,N_22071,N_20929);
nor U27980 (N_27980,N_20738,N_22132);
and U27981 (N_27981,N_22117,N_18764);
nand U27982 (N_27982,N_23618,N_22867);
nand U27983 (N_27983,N_19845,N_22576);
or U27984 (N_27984,N_23949,N_22029);
and U27985 (N_27985,N_18200,N_20321);
nor U27986 (N_27986,N_21234,N_18447);
and U27987 (N_27987,N_18458,N_22250);
and U27988 (N_27988,N_19420,N_20136);
xnor U27989 (N_27989,N_19775,N_20556);
or U27990 (N_27990,N_23772,N_22423);
nor U27991 (N_27991,N_18572,N_18082);
or U27992 (N_27992,N_19982,N_18010);
nand U27993 (N_27993,N_20202,N_20142);
and U27994 (N_27994,N_22491,N_20078);
and U27995 (N_27995,N_23092,N_18080);
nand U27996 (N_27996,N_21710,N_22691);
or U27997 (N_27997,N_23374,N_21924);
nor U27998 (N_27998,N_19381,N_23368);
or U27999 (N_27999,N_22268,N_19699);
xnor U28000 (N_28000,N_19564,N_21782);
or U28001 (N_28001,N_23693,N_19227);
nand U28002 (N_28002,N_19453,N_20955);
nor U28003 (N_28003,N_21183,N_20210);
xor U28004 (N_28004,N_23364,N_20522);
xnor U28005 (N_28005,N_20696,N_19307);
and U28006 (N_28006,N_21399,N_23874);
and U28007 (N_28007,N_18427,N_19912);
and U28008 (N_28008,N_22103,N_23709);
and U28009 (N_28009,N_21456,N_23450);
xnor U28010 (N_28010,N_23573,N_19961);
xnor U28011 (N_28011,N_22182,N_20313);
and U28012 (N_28012,N_19021,N_20296);
nand U28013 (N_28013,N_22821,N_21414);
nand U28014 (N_28014,N_19150,N_20756);
nor U28015 (N_28015,N_21202,N_18477);
nor U28016 (N_28016,N_20446,N_23318);
nor U28017 (N_28017,N_23483,N_18991);
nand U28018 (N_28018,N_19327,N_23330);
nor U28019 (N_28019,N_21250,N_21824);
or U28020 (N_28020,N_18907,N_23658);
and U28021 (N_28021,N_19328,N_18730);
and U28022 (N_28022,N_22993,N_22190);
or U28023 (N_28023,N_20374,N_21044);
xor U28024 (N_28024,N_19149,N_21917);
or U28025 (N_28025,N_19399,N_23970);
or U28026 (N_28026,N_18655,N_22365);
nor U28027 (N_28027,N_22442,N_20607);
nand U28028 (N_28028,N_23401,N_22062);
nand U28029 (N_28029,N_21832,N_23821);
and U28030 (N_28030,N_18491,N_19740);
and U28031 (N_28031,N_22282,N_22137);
and U28032 (N_28032,N_21920,N_22837);
or U28033 (N_28033,N_20126,N_23361);
and U28034 (N_28034,N_18262,N_18825);
nand U28035 (N_28035,N_21267,N_23773);
nand U28036 (N_28036,N_18039,N_20856);
or U28037 (N_28037,N_21201,N_18295);
or U28038 (N_28038,N_19155,N_19606);
nand U28039 (N_28039,N_19705,N_21805);
xnor U28040 (N_28040,N_22955,N_18368);
and U28041 (N_28041,N_20675,N_21837);
or U28042 (N_28042,N_20860,N_20212);
nand U28043 (N_28043,N_19020,N_23940);
and U28044 (N_28044,N_22950,N_19300);
nor U28045 (N_28045,N_21128,N_21554);
or U28046 (N_28046,N_20178,N_21484);
nand U28047 (N_28047,N_18264,N_20783);
nor U28048 (N_28048,N_22277,N_20518);
and U28049 (N_28049,N_23963,N_23763);
or U28050 (N_28050,N_23272,N_23323);
or U28051 (N_28051,N_23592,N_19704);
xnor U28052 (N_28052,N_22880,N_21572);
xor U28053 (N_28053,N_22472,N_20184);
xnor U28054 (N_28054,N_23544,N_18444);
or U28055 (N_28055,N_20880,N_22007);
xor U28056 (N_28056,N_23209,N_22852);
and U28057 (N_28057,N_23884,N_19716);
xor U28058 (N_28058,N_20219,N_18591);
nand U28059 (N_28059,N_18267,N_18354);
xnor U28060 (N_28060,N_22380,N_19976);
nand U28061 (N_28061,N_19029,N_19109);
nand U28062 (N_28062,N_23938,N_19452);
xnor U28063 (N_28063,N_22780,N_21567);
and U28064 (N_28064,N_21500,N_21561);
xor U28065 (N_28065,N_18753,N_19354);
or U28066 (N_28066,N_18081,N_22978);
nand U28067 (N_28067,N_21129,N_20535);
or U28068 (N_28068,N_23147,N_18967);
nand U28069 (N_28069,N_19225,N_23548);
and U28070 (N_28070,N_21401,N_19746);
and U28071 (N_28071,N_23023,N_20081);
and U28072 (N_28072,N_22344,N_19626);
nand U28073 (N_28073,N_18423,N_23567);
xnor U28074 (N_28074,N_20158,N_20562);
nor U28075 (N_28075,N_20958,N_20406);
or U28076 (N_28076,N_18771,N_23808);
nor U28077 (N_28077,N_19945,N_22963);
nor U28078 (N_28078,N_18073,N_19409);
nand U28079 (N_28079,N_19484,N_18272);
nand U28080 (N_28080,N_19776,N_19725);
or U28081 (N_28081,N_19167,N_18191);
nor U28082 (N_28082,N_23514,N_23117);
and U28083 (N_28083,N_21530,N_19977);
nor U28084 (N_28084,N_19834,N_21110);
nand U28085 (N_28085,N_18069,N_23414);
nor U28086 (N_28086,N_19178,N_23723);
nand U28087 (N_28087,N_18403,N_22266);
nand U28088 (N_28088,N_21709,N_18502);
nand U28089 (N_28089,N_21225,N_22261);
xnor U28090 (N_28090,N_18004,N_22313);
nor U28091 (N_28091,N_23189,N_20795);
or U28092 (N_28092,N_22574,N_23187);
and U28093 (N_28093,N_18880,N_23313);
and U28094 (N_28094,N_19308,N_21495);
nand U28095 (N_28095,N_19737,N_21481);
or U28096 (N_28096,N_19985,N_20433);
or U28097 (N_28097,N_22209,N_19619);
and U28098 (N_28098,N_21681,N_23152);
nor U28099 (N_28099,N_21037,N_21347);
or U28100 (N_28100,N_22124,N_21863);
nand U28101 (N_28101,N_21211,N_20719);
and U28102 (N_28102,N_21152,N_21339);
nand U28103 (N_28103,N_20648,N_20845);
and U28104 (N_28104,N_19215,N_20559);
and U28105 (N_28105,N_20639,N_19757);
nor U28106 (N_28106,N_22417,N_22059);
nand U28107 (N_28107,N_21413,N_21879);
or U28108 (N_28108,N_19674,N_23137);
and U28109 (N_28109,N_21811,N_23790);
nor U28110 (N_28110,N_19208,N_21330);
nor U28111 (N_28111,N_20581,N_22935);
nand U28112 (N_28112,N_23782,N_18729);
and U28113 (N_28113,N_19328,N_21658);
nor U28114 (N_28114,N_23945,N_20257);
nor U28115 (N_28115,N_23715,N_23230);
and U28116 (N_28116,N_19533,N_23578);
nor U28117 (N_28117,N_22011,N_22490);
and U28118 (N_28118,N_22044,N_21307);
nor U28119 (N_28119,N_21388,N_21656);
and U28120 (N_28120,N_23454,N_22582);
xor U28121 (N_28121,N_22868,N_21892);
nor U28122 (N_28122,N_18230,N_22483);
nor U28123 (N_28123,N_19018,N_22388);
and U28124 (N_28124,N_19597,N_21311);
or U28125 (N_28125,N_23841,N_18497);
or U28126 (N_28126,N_18823,N_21608);
nand U28127 (N_28127,N_22209,N_19744);
nand U28128 (N_28128,N_20330,N_20589);
and U28129 (N_28129,N_18154,N_22004);
nor U28130 (N_28130,N_22840,N_21402);
and U28131 (N_28131,N_18854,N_18472);
nand U28132 (N_28132,N_18402,N_20317);
nand U28133 (N_28133,N_23402,N_19894);
nor U28134 (N_28134,N_22474,N_19183);
and U28135 (N_28135,N_18868,N_20293);
or U28136 (N_28136,N_19334,N_20327);
or U28137 (N_28137,N_18029,N_18037);
or U28138 (N_28138,N_21626,N_23003);
or U28139 (N_28139,N_23965,N_19109);
nor U28140 (N_28140,N_23365,N_22673);
or U28141 (N_28141,N_22684,N_19366);
or U28142 (N_28142,N_19548,N_19871);
nor U28143 (N_28143,N_18215,N_22545);
nor U28144 (N_28144,N_20666,N_23578);
and U28145 (N_28145,N_22625,N_21696);
or U28146 (N_28146,N_19908,N_18025);
or U28147 (N_28147,N_18295,N_21401);
and U28148 (N_28148,N_22424,N_19485);
or U28149 (N_28149,N_19407,N_19840);
nor U28150 (N_28150,N_22957,N_23934);
or U28151 (N_28151,N_21006,N_23087);
xnor U28152 (N_28152,N_22317,N_22016);
nand U28153 (N_28153,N_23226,N_22604);
or U28154 (N_28154,N_18845,N_21327);
nand U28155 (N_28155,N_21837,N_18954);
and U28156 (N_28156,N_23306,N_19592);
or U28157 (N_28157,N_21025,N_18069);
nand U28158 (N_28158,N_23339,N_22180);
xor U28159 (N_28159,N_23838,N_22517);
nor U28160 (N_28160,N_20617,N_21041);
nand U28161 (N_28161,N_23619,N_21013);
and U28162 (N_28162,N_18972,N_22433);
nand U28163 (N_28163,N_20132,N_21528);
or U28164 (N_28164,N_21200,N_18934);
or U28165 (N_28165,N_22862,N_22749);
nor U28166 (N_28166,N_23539,N_18748);
and U28167 (N_28167,N_22667,N_19283);
nor U28168 (N_28168,N_22840,N_23825);
nand U28169 (N_28169,N_19601,N_18003);
nand U28170 (N_28170,N_19585,N_22659);
nor U28171 (N_28171,N_19992,N_18655);
and U28172 (N_28172,N_21548,N_20293);
or U28173 (N_28173,N_19406,N_18348);
and U28174 (N_28174,N_20585,N_20229);
or U28175 (N_28175,N_19723,N_22192);
nor U28176 (N_28176,N_19284,N_23886);
and U28177 (N_28177,N_22102,N_21176);
and U28178 (N_28178,N_22287,N_20481);
nand U28179 (N_28179,N_22879,N_19911);
nor U28180 (N_28180,N_21434,N_20380);
xor U28181 (N_28181,N_21777,N_20299);
nor U28182 (N_28182,N_23666,N_22548);
and U28183 (N_28183,N_20087,N_18694);
xnor U28184 (N_28184,N_18768,N_23798);
nor U28185 (N_28185,N_20014,N_19503);
nand U28186 (N_28186,N_19276,N_22393);
and U28187 (N_28187,N_20904,N_22048);
or U28188 (N_28188,N_23087,N_20055);
nor U28189 (N_28189,N_18936,N_19534);
xor U28190 (N_28190,N_21248,N_21792);
xnor U28191 (N_28191,N_18081,N_22472);
or U28192 (N_28192,N_20070,N_18172);
nor U28193 (N_28193,N_21153,N_21902);
and U28194 (N_28194,N_18160,N_20624);
and U28195 (N_28195,N_20882,N_18716);
nand U28196 (N_28196,N_18602,N_19888);
nand U28197 (N_28197,N_18620,N_20490);
and U28198 (N_28198,N_18435,N_21378);
xnor U28199 (N_28199,N_18942,N_19871);
nand U28200 (N_28200,N_19764,N_19655);
xor U28201 (N_28201,N_19025,N_21376);
or U28202 (N_28202,N_22845,N_18183);
and U28203 (N_28203,N_23829,N_19923);
or U28204 (N_28204,N_18651,N_22668);
or U28205 (N_28205,N_18148,N_18217);
or U28206 (N_28206,N_20189,N_19535);
nor U28207 (N_28207,N_18979,N_22658);
nand U28208 (N_28208,N_23974,N_22110);
and U28209 (N_28209,N_18898,N_23197);
xnor U28210 (N_28210,N_21019,N_20273);
or U28211 (N_28211,N_18180,N_18057);
nor U28212 (N_28212,N_23350,N_23297);
nand U28213 (N_28213,N_22975,N_23772);
xor U28214 (N_28214,N_19595,N_20739);
nor U28215 (N_28215,N_21348,N_22313);
or U28216 (N_28216,N_18220,N_21567);
or U28217 (N_28217,N_20530,N_19130);
xnor U28218 (N_28218,N_18066,N_22912);
nor U28219 (N_28219,N_21232,N_22172);
nand U28220 (N_28220,N_20364,N_22456);
xor U28221 (N_28221,N_23742,N_20393);
nand U28222 (N_28222,N_21222,N_23099);
nand U28223 (N_28223,N_21364,N_20020);
and U28224 (N_28224,N_22894,N_21534);
and U28225 (N_28225,N_22999,N_22918);
or U28226 (N_28226,N_21189,N_23888);
or U28227 (N_28227,N_19063,N_21201);
xor U28228 (N_28228,N_20086,N_22466);
or U28229 (N_28229,N_23601,N_21044);
xnor U28230 (N_28230,N_22470,N_19084);
nor U28231 (N_28231,N_21956,N_23219);
or U28232 (N_28232,N_22936,N_20228);
nor U28233 (N_28233,N_22680,N_23848);
nor U28234 (N_28234,N_18757,N_23759);
nand U28235 (N_28235,N_20584,N_23954);
and U28236 (N_28236,N_21551,N_20216);
nand U28237 (N_28237,N_18142,N_22322);
or U28238 (N_28238,N_23910,N_18302);
or U28239 (N_28239,N_18779,N_19502);
nand U28240 (N_28240,N_18439,N_19339);
nor U28241 (N_28241,N_18473,N_18728);
nand U28242 (N_28242,N_20655,N_20904);
or U28243 (N_28243,N_20656,N_21502);
or U28244 (N_28244,N_20169,N_20058);
xnor U28245 (N_28245,N_18646,N_23527);
or U28246 (N_28246,N_21220,N_20845);
xor U28247 (N_28247,N_20660,N_23939);
nor U28248 (N_28248,N_19431,N_21524);
or U28249 (N_28249,N_21145,N_18000);
xnor U28250 (N_28250,N_21355,N_22798);
nor U28251 (N_28251,N_22354,N_23067);
and U28252 (N_28252,N_20420,N_23436);
nand U28253 (N_28253,N_19083,N_23502);
nor U28254 (N_28254,N_19435,N_23028);
and U28255 (N_28255,N_20690,N_19321);
nand U28256 (N_28256,N_23968,N_18906);
xnor U28257 (N_28257,N_22613,N_20938);
nand U28258 (N_28258,N_18706,N_19896);
nand U28259 (N_28259,N_23937,N_18495);
nor U28260 (N_28260,N_23477,N_18524);
nand U28261 (N_28261,N_22955,N_18184);
nand U28262 (N_28262,N_18057,N_18898);
or U28263 (N_28263,N_23860,N_23160);
or U28264 (N_28264,N_21136,N_23648);
nor U28265 (N_28265,N_22409,N_20429);
nor U28266 (N_28266,N_22904,N_22976);
or U28267 (N_28267,N_18539,N_22498);
and U28268 (N_28268,N_23033,N_19055);
nor U28269 (N_28269,N_23462,N_23977);
xnor U28270 (N_28270,N_20799,N_23377);
and U28271 (N_28271,N_23850,N_20353);
nand U28272 (N_28272,N_19615,N_20466);
and U28273 (N_28273,N_22759,N_21218);
and U28274 (N_28274,N_19049,N_20000);
nor U28275 (N_28275,N_19017,N_23784);
nor U28276 (N_28276,N_18052,N_20395);
and U28277 (N_28277,N_20494,N_21862);
nor U28278 (N_28278,N_21402,N_22591);
nor U28279 (N_28279,N_22042,N_22280);
nor U28280 (N_28280,N_21796,N_20447);
nor U28281 (N_28281,N_19224,N_22815);
and U28282 (N_28282,N_23934,N_20632);
or U28283 (N_28283,N_23364,N_23976);
nand U28284 (N_28284,N_21938,N_18005);
nand U28285 (N_28285,N_20866,N_22857);
and U28286 (N_28286,N_21802,N_23986);
or U28287 (N_28287,N_22421,N_23266);
xnor U28288 (N_28288,N_19563,N_23300);
nand U28289 (N_28289,N_18987,N_22773);
and U28290 (N_28290,N_22977,N_18548);
or U28291 (N_28291,N_22864,N_20663);
or U28292 (N_28292,N_20109,N_18299);
and U28293 (N_28293,N_18594,N_21704);
or U28294 (N_28294,N_20686,N_18372);
and U28295 (N_28295,N_19376,N_23654);
nand U28296 (N_28296,N_23233,N_18906);
nor U28297 (N_28297,N_21834,N_19937);
nand U28298 (N_28298,N_19439,N_19959);
or U28299 (N_28299,N_22415,N_18602);
or U28300 (N_28300,N_20612,N_19256);
nand U28301 (N_28301,N_20662,N_18540);
and U28302 (N_28302,N_19771,N_23103);
nand U28303 (N_28303,N_22096,N_21111);
or U28304 (N_28304,N_22094,N_18580);
and U28305 (N_28305,N_23660,N_22200);
and U28306 (N_28306,N_23552,N_19776);
or U28307 (N_28307,N_18818,N_22628);
and U28308 (N_28308,N_21301,N_23887);
nor U28309 (N_28309,N_21642,N_19622);
nand U28310 (N_28310,N_18414,N_19275);
xnor U28311 (N_28311,N_21607,N_23886);
nor U28312 (N_28312,N_18166,N_20207);
or U28313 (N_28313,N_23540,N_23890);
nand U28314 (N_28314,N_23675,N_22733);
and U28315 (N_28315,N_19888,N_22820);
and U28316 (N_28316,N_23736,N_21314);
nand U28317 (N_28317,N_23004,N_19596);
and U28318 (N_28318,N_23275,N_21298);
nor U28319 (N_28319,N_18755,N_18795);
nor U28320 (N_28320,N_21407,N_21895);
xnor U28321 (N_28321,N_21898,N_18448);
nand U28322 (N_28322,N_21429,N_20349);
or U28323 (N_28323,N_18291,N_21446);
xnor U28324 (N_28324,N_23467,N_20712);
and U28325 (N_28325,N_23732,N_20278);
nor U28326 (N_28326,N_19229,N_22175);
and U28327 (N_28327,N_23075,N_19440);
and U28328 (N_28328,N_18019,N_20254);
and U28329 (N_28329,N_18141,N_18620);
and U28330 (N_28330,N_19331,N_18073);
nor U28331 (N_28331,N_23961,N_18198);
nor U28332 (N_28332,N_23739,N_19804);
and U28333 (N_28333,N_20916,N_23140);
and U28334 (N_28334,N_19641,N_23018);
nor U28335 (N_28335,N_20508,N_20970);
xor U28336 (N_28336,N_22273,N_20964);
nor U28337 (N_28337,N_19517,N_22643);
and U28338 (N_28338,N_23756,N_18219);
or U28339 (N_28339,N_22260,N_20103);
and U28340 (N_28340,N_19348,N_23076);
and U28341 (N_28341,N_23032,N_22717);
and U28342 (N_28342,N_22106,N_22643);
and U28343 (N_28343,N_20440,N_21128);
or U28344 (N_28344,N_22909,N_20046);
xor U28345 (N_28345,N_18692,N_23433);
nand U28346 (N_28346,N_18447,N_22183);
and U28347 (N_28347,N_18861,N_21203);
nor U28348 (N_28348,N_18811,N_23701);
nor U28349 (N_28349,N_18200,N_20599);
nor U28350 (N_28350,N_19907,N_22375);
or U28351 (N_28351,N_22405,N_19508);
nor U28352 (N_28352,N_18503,N_19813);
and U28353 (N_28353,N_21995,N_18923);
nand U28354 (N_28354,N_20037,N_21666);
xor U28355 (N_28355,N_23092,N_19022);
or U28356 (N_28356,N_23639,N_19729);
nor U28357 (N_28357,N_21026,N_20695);
nor U28358 (N_28358,N_20825,N_18537);
or U28359 (N_28359,N_19165,N_19496);
nand U28360 (N_28360,N_21799,N_18872);
and U28361 (N_28361,N_23978,N_23020);
nor U28362 (N_28362,N_21236,N_22283);
nor U28363 (N_28363,N_20699,N_21028);
nor U28364 (N_28364,N_19184,N_23507);
or U28365 (N_28365,N_19650,N_19915);
and U28366 (N_28366,N_18430,N_20255);
or U28367 (N_28367,N_23352,N_18754);
and U28368 (N_28368,N_18566,N_19064);
nor U28369 (N_28369,N_20387,N_23188);
nor U28370 (N_28370,N_22524,N_22728);
nand U28371 (N_28371,N_21958,N_19538);
nor U28372 (N_28372,N_19553,N_23954);
or U28373 (N_28373,N_20835,N_22002);
nor U28374 (N_28374,N_20837,N_20614);
nor U28375 (N_28375,N_21036,N_20343);
and U28376 (N_28376,N_20727,N_19856);
or U28377 (N_28377,N_18715,N_23721);
and U28378 (N_28378,N_20496,N_20132);
or U28379 (N_28379,N_21964,N_23723);
nor U28380 (N_28380,N_20902,N_22397);
or U28381 (N_28381,N_18681,N_22062);
and U28382 (N_28382,N_21214,N_18156);
nand U28383 (N_28383,N_18191,N_21145);
and U28384 (N_28384,N_20091,N_18466);
xnor U28385 (N_28385,N_23683,N_23041);
or U28386 (N_28386,N_23015,N_18387);
nor U28387 (N_28387,N_20520,N_23380);
nand U28388 (N_28388,N_23946,N_21947);
nor U28389 (N_28389,N_23704,N_22604);
nor U28390 (N_28390,N_22137,N_18738);
or U28391 (N_28391,N_19586,N_18876);
nor U28392 (N_28392,N_20243,N_19288);
and U28393 (N_28393,N_18900,N_20990);
xnor U28394 (N_28394,N_23273,N_20063);
xnor U28395 (N_28395,N_19384,N_20633);
xnor U28396 (N_28396,N_18383,N_20819);
xnor U28397 (N_28397,N_22823,N_21917);
nand U28398 (N_28398,N_22928,N_21079);
nor U28399 (N_28399,N_21851,N_18409);
or U28400 (N_28400,N_18335,N_20837);
nand U28401 (N_28401,N_18419,N_21499);
nor U28402 (N_28402,N_20633,N_23307);
and U28403 (N_28403,N_23262,N_18045);
nor U28404 (N_28404,N_23625,N_19210);
nand U28405 (N_28405,N_21863,N_19462);
nand U28406 (N_28406,N_22486,N_20565);
or U28407 (N_28407,N_19717,N_22147);
and U28408 (N_28408,N_21678,N_21571);
or U28409 (N_28409,N_18340,N_20174);
or U28410 (N_28410,N_19635,N_23389);
xor U28411 (N_28411,N_18626,N_23366);
nor U28412 (N_28412,N_18548,N_22935);
and U28413 (N_28413,N_22935,N_20728);
and U28414 (N_28414,N_23328,N_18542);
and U28415 (N_28415,N_20223,N_22593);
or U28416 (N_28416,N_18437,N_23460);
nor U28417 (N_28417,N_21484,N_20604);
nand U28418 (N_28418,N_20917,N_21648);
nand U28419 (N_28419,N_23371,N_20437);
nand U28420 (N_28420,N_18084,N_22273);
or U28421 (N_28421,N_21411,N_19787);
nor U28422 (N_28422,N_23994,N_18158);
and U28423 (N_28423,N_18654,N_20569);
and U28424 (N_28424,N_20113,N_22326);
and U28425 (N_28425,N_19516,N_23771);
nand U28426 (N_28426,N_18236,N_21836);
and U28427 (N_28427,N_23425,N_22307);
and U28428 (N_28428,N_19407,N_23730);
nor U28429 (N_28429,N_18353,N_18627);
or U28430 (N_28430,N_20537,N_19446);
nand U28431 (N_28431,N_19147,N_18524);
nor U28432 (N_28432,N_22374,N_23985);
and U28433 (N_28433,N_19029,N_22461);
or U28434 (N_28434,N_23341,N_20397);
or U28435 (N_28435,N_22155,N_23599);
nand U28436 (N_28436,N_23583,N_18899);
and U28437 (N_28437,N_22545,N_18478);
nor U28438 (N_28438,N_18834,N_19899);
or U28439 (N_28439,N_20478,N_21528);
and U28440 (N_28440,N_18369,N_23118);
nand U28441 (N_28441,N_18072,N_19530);
and U28442 (N_28442,N_21851,N_22885);
nor U28443 (N_28443,N_19771,N_23269);
or U28444 (N_28444,N_23644,N_18601);
xor U28445 (N_28445,N_21498,N_22732);
and U28446 (N_28446,N_23310,N_23950);
or U28447 (N_28447,N_21110,N_18010);
and U28448 (N_28448,N_20787,N_18255);
nand U28449 (N_28449,N_23986,N_18979);
nor U28450 (N_28450,N_22785,N_18966);
and U28451 (N_28451,N_19503,N_19324);
nand U28452 (N_28452,N_23281,N_18696);
nand U28453 (N_28453,N_18617,N_23983);
nand U28454 (N_28454,N_23835,N_23251);
nand U28455 (N_28455,N_18004,N_19640);
and U28456 (N_28456,N_18563,N_20523);
and U28457 (N_28457,N_23502,N_23410);
nor U28458 (N_28458,N_18200,N_19185);
and U28459 (N_28459,N_19706,N_23217);
nor U28460 (N_28460,N_18957,N_23871);
and U28461 (N_28461,N_18574,N_19089);
or U28462 (N_28462,N_20172,N_21149);
and U28463 (N_28463,N_22422,N_22806);
and U28464 (N_28464,N_18868,N_20649);
nor U28465 (N_28465,N_22256,N_21176);
nor U28466 (N_28466,N_20697,N_19672);
or U28467 (N_28467,N_21976,N_20452);
and U28468 (N_28468,N_18375,N_18436);
nand U28469 (N_28469,N_20440,N_18672);
nand U28470 (N_28470,N_22633,N_22523);
nor U28471 (N_28471,N_19148,N_21788);
nor U28472 (N_28472,N_21274,N_20367);
and U28473 (N_28473,N_22579,N_21116);
xnor U28474 (N_28474,N_19635,N_20751);
nand U28475 (N_28475,N_18565,N_21100);
nor U28476 (N_28476,N_19107,N_20807);
xor U28477 (N_28477,N_21830,N_18467);
nand U28478 (N_28478,N_20849,N_23190);
nor U28479 (N_28479,N_23308,N_19229);
nor U28480 (N_28480,N_18602,N_18106);
and U28481 (N_28481,N_18970,N_18202);
nand U28482 (N_28482,N_21311,N_21163);
nor U28483 (N_28483,N_18073,N_22118);
xor U28484 (N_28484,N_20219,N_19884);
nand U28485 (N_28485,N_20376,N_19657);
nand U28486 (N_28486,N_23470,N_18930);
nor U28487 (N_28487,N_18469,N_19592);
and U28488 (N_28488,N_22318,N_20902);
or U28489 (N_28489,N_22589,N_20388);
xnor U28490 (N_28490,N_18834,N_21140);
xor U28491 (N_28491,N_19962,N_19469);
nor U28492 (N_28492,N_22649,N_18156);
nand U28493 (N_28493,N_22414,N_20918);
nand U28494 (N_28494,N_20543,N_19115);
xor U28495 (N_28495,N_22890,N_23043);
nand U28496 (N_28496,N_18928,N_18686);
or U28497 (N_28497,N_21467,N_18179);
or U28498 (N_28498,N_22217,N_18289);
nor U28499 (N_28499,N_18481,N_19118);
or U28500 (N_28500,N_20439,N_21788);
or U28501 (N_28501,N_19775,N_20394);
nand U28502 (N_28502,N_19141,N_23034);
nor U28503 (N_28503,N_21522,N_22716);
nor U28504 (N_28504,N_23958,N_18208);
and U28505 (N_28505,N_20753,N_18483);
nand U28506 (N_28506,N_20414,N_18866);
nor U28507 (N_28507,N_22987,N_22424);
nor U28508 (N_28508,N_18598,N_23592);
nand U28509 (N_28509,N_23304,N_23554);
nor U28510 (N_28510,N_19117,N_20792);
xnor U28511 (N_28511,N_18277,N_21294);
nor U28512 (N_28512,N_19850,N_22295);
and U28513 (N_28513,N_20059,N_19933);
nor U28514 (N_28514,N_20853,N_21898);
or U28515 (N_28515,N_20255,N_22941);
or U28516 (N_28516,N_21181,N_21656);
and U28517 (N_28517,N_22165,N_22495);
or U28518 (N_28518,N_23289,N_19617);
nor U28519 (N_28519,N_18903,N_21348);
or U28520 (N_28520,N_21497,N_21003);
and U28521 (N_28521,N_18051,N_23928);
nor U28522 (N_28522,N_20015,N_22598);
nor U28523 (N_28523,N_23337,N_21157);
xnor U28524 (N_28524,N_23894,N_20332);
xor U28525 (N_28525,N_21837,N_22928);
or U28526 (N_28526,N_19373,N_22110);
and U28527 (N_28527,N_18819,N_20576);
nor U28528 (N_28528,N_22216,N_18693);
nor U28529 (N_28529,N_22399,N_23067);
and U28530 (N_28530,N_23474,N_21064);
nor U28531 (N_28531,N_20961,N_21379);
and U28532 (N_28532,N_23302,N_22444);
nor U28533 (N_28533,N_21155,N_18665);
nor U28534 (N_28534,N_18124,N_23990);
nand U28535 (N_28535,N_23372,N_18148);
or U28536 (N_28536,N_19402,N_20278);
nor U28537 (N_28537,N_19135,N_20296);
or U28538 (N_28538,N_19002,N_18082);
nor U28539 (N_28539,N_22275,N_18301);
nor U28540 (N_28540,N_21621,N_22041);
nor U28541 (N_28541,N_18770,N_23251);
and U28542 (N_28542,N_19514,N_20086);
xnor U28543 (N_28543,N_21910,N_19325);
nand U28544 (N_28544,N_22074,N_23605);
nand U28545 (N_28545,N_21046,N_19134);
and U28546 (N_28546,N_18007,N_23978);
or U28547 (N_28547,N_23255,N_18100);
or U28548 (N_28548,N_18629,N_18075);
or U28549 (N_28549,N_22296,N_21281);
or U28550 (N_28550,N_19792,N_23131);
xor U28551 (N_28551,N_18786,N_18229);
and U28552 (N_28552,N_20933,N_22882);
nand U28553 (N_28553,N_19225,N_22289);
and U28554 (N_28554,N_20536,N_19169);
or U28555 (N_28555,N_21583,N_22625);
and U28556 (N_28556,N_23759,N_20506);
or U28557 (N_28557,N_22530,N_22037);
nor U28558 (N_28558,N_21658,N_23068);
and U28559 (N_28559,N_22363,N_20909);
nand U28560 (N_28560,N_22690,N_23357);
nor U28561 (N_28561,N_20773,N_21668);
nor U28562 (N_28562,N_20851,N_18445);
and U28563 (N_28563,N_21197,N_23035);
or U28564 (N_28564,N_20707,N_19430);
nand U28565 (N_28565,N_22834,N_19865);
nand U28566 (N_28566,N_18086,N_21973);
nor U28567 (N_28567,N_19986,N_20311);
xor U28568 (N_28568,N_20664,N_19014);
nor U28569 (N_28569,N_18350,N_19572);
nand U28570 (N_28570,N_20597,N_22541);
and U28571 (N_28571,N_19768,N_19562);
nand U28572 (N_28572,N_19349,N_23458);
xnor U28573 (N_28573,N_18092,N_20755);
or U28574 (N_28574,N_18537,N_22142);
and U28575 (N_28575,N_20457,N_23737);
and U28576 (N_28576,N_20395,N_22219);
nor U28577 (N_28577,N_20124,N_20352);
nand U28578 (N_28578,N_21195,N_18299);
or U28579 (N_28579,N_18892,N_19642);
nand U28580 (N_28580,N_18124,N_20418);
nand U28581 (N_28581,N_23399,N_23218);
nor U28582 (N_28582,N_19617,N_21297);
or U28583 (N_28583,N_23270,N_21578);
nand U28584 (N_28584,N_23524,N_19512);
nor U28585 (N_28585,N_21437,N_20378);
nand U28586 (N_28586,N_18832,N_20975);
or U28587 (N_28587,N_22603,N_21539);
or U28588 (N_28588,N_19857,N_23710);
nor U28589 (N_28589,N_19127,N_22064);
or U28590 (N_28590,N_23225,N_21129);
and U28591 (N_28591,N_19343,N_22182);
nor U28592 (N_28592,N_18240,N_23822);
xor U28593 (N_28593,N_20744,N_23683);
or U28594 (N_28594,N_19870,N_19347);
nor U28595 (N_28595,N_20229,N_22763);
nand U28596 (N_28596,N_21261,N_21656);
nand U28597 (N_28597,N_19736,N_22034);
nand U28598 (N_28598,N_18282,N_22702);
and U28599 (N_28599,N_18385,N_22668);
xnor U28600 (N_28600,N_22602,N_18471);
and U28601 (N_28601,N_20939,N_20135);
nor U28602 (N_28602,N_18702,N_23744);
and U28603 (N_28603,N_19436,N_23697);
and U28604 (N_28604,N_19764,N_19165);
and U28605 (N_28605,N_22805,N_23082);
and U28606 (N_28606,N_23099,N_19226);
or U28607 (N_28607,N_23705,N_18813);
nor U28608 (N_28608,N_22250,N_18508);
and U28609 (N_28609,N_19547,N_19385);
or U28610 (N_28610,N_23194,N_23285);
or U28611 (N_28611,N_21138,N_19541);
xor U28612 (N_28612,N_18013,N_19580);
or U28613 (N_28613,N_18522,N_20707);
and U28614 (N_28614,N_23393,N_23532);
or U28615 (N_28615,N_23885,N_21232);
or U28616 (N_28616,N_18133,N_20153);
nor U28617 (N_28617,N_20650,N_19229);
nor U28618 (N_28618,N_21654,N_22346);
or U28619 (N_28619,N_22202,N_21585);
nand U28620 (N_28620,N_19984,N_21389);
or U28621 (N_28621,N_21842,N_19557);
or U28622 (N_28622,N_20639,N_20354);
nor U28623 (N_28623,N_19732,N_22950);
nand U28624 (N_28624,N_22836,N_19043);
and U28625 (N_28625,N_19249,N_19999);
and U28626 (N_28626,N_20663,N_23230);
nor U28627 (N_28627,N_23198,N_18011);
nand U28628 (N_28628,N_22951,N_23258);
or U28629 (N_28629,N_23506,N_20164);
and U28630 (N_28630,N_20762,N_21902);
nor U28631 (N_28631,N_23218,N_18582);
nand U28632 (N_28632,N_18116,N_22373);
xor U28633 (N_28633,N_18201,N_22275);
nor U28634 (N_28634,N_18191,N_21214);
or U28635 (N_28635,N_22506,N_20227);
nand U28636 (N_28636,N_21783,N_19146);
and U28637 (N_28637,N_22924,N_20549);
and U28638 (N_28638,N_18527,N_22639);
or U28639 (N_28639,N_22755,N_18714);
nor U28640 (N_28640,N_23153,N_19889);
nor U28641 (N_28641,N_18553,N_18489);
nor U28642 (N_28642,N_18963,N_19526);
nor U28643 (N_28643,N_18026,N_18427);
and U28644 (N_28644,N_23532,N_23251);
nor U28645 (N_28645,N_19144,N_23404);
nor U28646 (N_28646,N_22011,N_18168);
nand U28647 (N_28647,N_23634,N_22716);
or U28648 (N_28648,N_21255,N_21682);
nand U28649 (N_28649,N_18849,N_20295);
nor U28650 (N_28650,N_18669,N_21251);
and U28651 (N_28651,N_18234,N_23305);
nand U28652 (N_28652,N_22515,N_22461);
nand U28653 (N_28653,N_19015,N_19778);
and U28654 (N_28654,N_23401,N_18442);
and U28655 (N_28655,N_19884,N_19511);
nor U28656 (N_28656,N_20764,N_20630);
or U28657 (N_28657,N_18623,N_20339);
or U28658 (N_28658,N_22656,N_22286);
nand U28659 (N_28659,N_23501,N_20791);
nand U28660 (N_28660,N_22261,N_20883);
nand U28661 (N_28661,N_21485,N_21897);
nand U28662 (N_28662,N_18934,N_20327);
xnor U28663 (N_28663,N_20709,N_18058);
and U28664 (N_28664,N_18237,N_22654);
or U28665 (N_28665,N_23234,N_21476);
and U28666 (N_28666,N_18767,N_22251);
nor U28667 (N_28667,N_23995,N_22444);
or U28668 (N_28668,N_18464,N_18181);
or U28669 (N_28669,N_22199,N_20403);
nand U28670 (N_28670,N_22332,N_18982);
and U28671 (N_28671,N_21405,N_22570);
nor U28672 (N_28672,N_22836,N_21689);
xor U28673 (N_28673,N_20411,N_23892);
and U28674 (N_28674,N_18065,N_18111);
nor U28675 (N_28675,N_22075,N_19193);
nor U28676 (N_28676,N_23331,N_21695);
or U28677 (N_28677,N_21232,N_19763);
nand U28678 (N_28678,N_20200,N_19100);
and U28679 (N_28679,N_22758,N_21156);
or U28680 (N_28680,N_18222,N_21822);
and U28681 (N_28681,N_23590,N_19591);
and U28682 (N_28682,N_21099,N_23889);
xnor U28683 (N_28683,N_20891,N_22611);
or U28684 (N_28684,N_18913,N_19532);
nor U28685 (N_28685,N_19470,N_18460);
nand U28686 (N_28686,N_22278,N_21646);
and U28687 (N_28687,N_22267,N_23145);
nand U28688 (N_28688,N_21404,N_23279);
or U28689 (N_28689,N_18883,N_22847);
nor U28690 (N_28690,N_21658,N_23094);
or U28691 (N_28691,N_22459,N_19451);
and U28692 (N_28692,N_23167,N_19885);
and U28693 (N_28693,N_18620,N_22987);
nor U28694 (N_28694,N_19798,N_20384);
nor U28695 (N_28695,N_22177,N_22692);
nand U28696 (N_28696,N_19566,N_23807);
or U28697 (N_28697,N_22788,N_20740);
or U28698 (N_28698,N_22709,N_18886);
nor U28699 (N_28699,N_19323,N_18223);
nor U28700 (N_28700,N_18780,N_19264);
xor U28701 (N_28701,N_22875,N_21963);
and U28702 (N_28702,N_23534,N_21075);
nor U28703 (N_28703,N_20231,N_20391);
and U28704 (N_28704,N_18293,N_20050);
xor U28705 (N_28705,N_22707,N_23999);
nand U28706 (N_28706,N_18083,N_23306);
nand U28707 (N_28707,N_21445,N_20254);
and U28708 (N_28708,N_22261,N_23821);
nor U28709 (N_28709,N_21635,N_18758);
nor U28710 (N_28710,N_22780,N_20327);
and U28711 (N_28711,N_18453,N_19929);
and U28712 (N_28712,N_20695,N_23937);
nor U28713 (N_28713,N_23721,N_21813);
nand U28714 (N_28714,N_19886,N_19222);
nand U28715 (N_28715,N_21834,N_23862);
or U28716 (N_28716,N_22403,N_23978);
nand U28717 (N_28717,N_20017,N_23088);
xor U28718 (N_28718,N_22048,N_22860);
nand U28719 (N_28719,N_19651,N_18417);
nand U28720 (N_28720,N_21442,N_19722);
and U28721 (N_28721,N_21266,N_18635);
nor U28722 (N_28722,N_23067,N_23825);
nor U28723 (N_28723,N_20809,N_19803);
or U28724 (N_28724,N_20356,N_20040);
xor U28725 (N_28725,N_23198,N_18303);
nand U28726 (N_28726,N_23868,N_22068);
nand U28727 (N_28727,N_21652,N_20566);
and U28728 (N_28728,N_18803,N_20303);
nor U28729 (N_28729,N_21283,N_23470);
nand U28730 (N_28730,N_22640,N_23612);
nand U28731 (N_28731,N_19633,N_21994);
nor U28732 (N_28732,N_18886,N_20743);
nand U28733 (N_28733,N_23137,N_18865);
and U28734 (N_28734,N_20615,N_20738);
nor U28735 (N_28735,N_21144,N_21639);
xnor U28736 (N_28736,N_19252,N_21870);
nor U28737 (N_28737,N_22638,N_21405);
and U28738 (N_28738,N_19928,N_22580);
nor U28739 (N_28739,N_20305,N_19760);
or U28740 (N_28740,N_22594,N_19700);
nand U28741 (N_28741,N_21259,N_21878);
xnor U28742 (N_28742,N_19343,N_23073);
xor U28743 (N_28743,N_18588,N_19391);
and U28744 (N_28744,N_18574,N_20460);
and U28745 (N_28745,N_19923,N_19715);
nor U28746 (N_28746,N_18459,N_22221);
and U28747 (N_28747,N_18129,N_20371);
and U28748 (N_28748,N_18396,N_22987);
and U28749 (N_28749,N_21148,N_20192);
nor U28750 (N_28750,N_19094,N_19720);
and U28751 (N_28751,N_19485,N_19291);
and U28752 (N_28752,N_18611,N_22374);
nand U28753 (N_28753,N_20228,N_23189);
or U28754 (N_28754,N_21735,N_19897);
nor U28755 (N_28755,N_20666,N_23212);
nor U28756 (N_28756,N_19561,N_21221);
or U28757 (N_28757,N_22761,N_18784);
nand U28758 (N_28758,N_22795,N_19814);
or U28759 (N_28759,N_22891,N_18859);
nor U28760 (N_28760,N_18317,N_18415);
nor U28761 (N_28761,N_19652,N_23122);
nand U28762 (N_28762,N_20425,N_18793);
nor U28763 (N_28763,N_23719,N_21126);
nand U28764 (N_28764,N_20460,N_21798);
nand U28765 (N_28765,N_21063,N_23230);
nand U28766 (N_28766,N_20173,N_18870);
or U28767 (N_28767,N_18664,N_19064);
nor U28768 (N_28768,N_22498,N_22262);
nor U28769 (N_28769,N_19541,N_19770);
or U28770 (N_28770,N_23468,N_18765);
xor U28771 (N_28771,N_18079,N_22471);
nor U28772 (N_28772,N_21124,N_23439);
and U28773 (N_28773,N_19184,N_23945);
or U28774 (N_28774,N_23900,N_22692);
nand U28775 (N_28775,N_18423,N_22236);
xnor U28776 (N_28776,N_22638,N_19367);
and U28777 (N_28777,N_19500,N_23157);
nor U28778 (N_28778,N_22186,N_18409);
or U28779 (N_28779,N_21988,N_23633);
and U28780 (N_28780,N_18224,N_21681);
nand U28781 (N_28781,N_21539,N_19425);
or U28782 (N_28782,N_20375,N_19860);
nor U28783 (N_28783,N_20685,N_23291);
nor U28784 (N_28784,N_22635,N_21347);
nor U28785 (N_28785,N_18777,N_20093);
or U28786 (N_28786,N_22559,N_23591);
nand U28787 (N_28787,N_20782,N_18733);
nand U28788 (N_28788,N_19136,N_18792);
nor U28789 (N_28789,N_18908,N_22533);
or U28790 (N_28790,N_23053,N_22954);
or U28791 (N_28791,N_20310,N_20297);
nand U28792 (N_28792,N_22916,N_19614);
or U28793 (N_28793,N_23832,N_22271);
and U28794 (N_28794,N_22825,N_18001);
xor U28795 (N_28795,N_21767,N_23933);
xor U28796 (N_28796,N_19195,N_20548);
xnor U28797 (N_28797,N_21187,N_18564);
or U28798 (N_28798,N_20939,N_19291);
and U28799 (N_28799,N_19202,N_18636);
or U28800 (N_28800,N_20632,N_19278);
nor U28801 (N_28801,N_22441,N_18886);
nor U28802 (N_28802,N_21756,N_22022);
and U28803 (N_28803,N_21095,N_21132);
and U28804 (N_28804,N_20105,N_20887);
nand U28805 (N_28805,N_18111,N_22567);
or U28806 (N_28806,N_18102,N_23787);
or U28807 (N_28807,N_21868,N_19953);
xnor U28808 (N_28808,N_21523,N_19116);
xor U28809 (N_28809,N_22719,N_22295);
nor U28810 (N_28810,N_23382,N_23855);
or U28811 (N_28811,N_21322,N_20413);
nor U28812 (N_28812,N_21493,N_22795);
nand U28813 (N_28813,N_18957,N_21801);
or U28814 (N_28814,N_22855,N_22582);
or U28815 (N_28815,N_22402,N_23107);
nor U28816 (N_28816,N_22814,N_21589);
nand U28817 (N_28817,N_19344,N_20831);
xnor U28818 (N_28818,N_21858,N_22842);
and U28819 (N_28819,N_18559,N_20413);
nand U28820 (N_28820,N_21857,N_19825);
nand U28821 (N_28821,N_20164,N_18954);
and U28822 (N_28822,N_23482,N_19093);
or U28823 (N_28823,N_23608,N_21175);
and U28824 (N_28824,N_19321,N_21575);
nor U28825 (N_28825,N_19945,N_22514);
or U28826 (N_28826,N_21338,N_18405);
and U28827 (N_28827,N_19322,N_18224);
nor U28828 (N_28828,N_18179,N_21434);
or U28829 (N_28829,N_19329,N_23808);
nand U28830 (N_28830,N_21419,N_20833);
xor U28831 (N_28831,N_19986,N_18475);
and U28832 (N_28832,N_18163,N_22127);
xnor U28833 (N_28833,N_19932,N_20714);
nand U28834 (N_28834,N_23885,N_18537);
nand U28835 (N_28835,N_22312,N_22903);
nand U28836 (N_28836,N_23395,N_18047);
nand U28837 (N_28837,N_21976,N_19111);
nand U28838 (N_28838,N_23694,N_20696);
or U28839 (N_28839,N_22866,N_18194);
nand U28840 (N_28840,N_19914,N_22997);
nand U28841 (N_28841,N_23282,N_19308);
or U28842 (N_28842,N_22088,N_20827);
nor U28843 (N_28843,N_22822,N_18767);
nor U28844 (N_28844,N_20130,N_19574);
nor U28845 (N_28845,N_21724,N_22256);
or U28846 (N_28846,N_21974,N_22802);
or U28847 (N_28847,N_22398,N_21125);
nor U28848 (N_28848,N_20507,N_22705);
nor U28849 (N_28849,N_21924,N_23756);
nand U28850 (N_28850,N_22635,N_23892);
nand U28851 (N_28851,N_23255,N_21835);
or U28852 (N_28852,N_21222,N_19411);
xor U28853 (N_28853,N_22499,N_23249);
nor U28854 (N_28854,N_19909,N_18013);
and U28855 (N_28855,N_21695,N_18683);
nor U28856 (N_28856,N_23531,N_18425);
xor U28857 (N_28857,N_22744,N_18388);
and U28858 (N_28858,N_18154,N_19438);
and U28859 (N_28859,N_18774,N_18931);
and U28860 (N_28860,N_21284,N_19311);
nor U28861 (N_28861,N_19326,N_23623);
and U28862 (N_28862,N_20885,N_22780);
nor U28863 (N_28863,N_18634,N_22186);
nor U28864 (N_28864,N_20352,N_19493);
or U28865 (N_28865,N_20606,N_19691);
nand U28866 (N_28866,N_19512,N_18743);
nor U28867 (N_28867,N_22666,N_20426);
nor U28868 (N_28868,N_22482,N_18785);
xnor U28869 (N_28869,N_21995,N_23665);
and U28870 (N_28870,N_18800,N_19359);
nor U28871 (N_28871,N_21401,N_21132);
or U28872 (N_28872,N_20947,N_20167);
nand U28873 (N_28873,N_21870,N_19673);
and U28874 (N_28874,N_23921,N_22581);
nor U28875 (N_28875,N_20241,N_22183);
and U28876 (N_28876,N_22916,N_20594);
and U28877 (N_28877,N_22219,N_18844);
nand U28878 (N_28878,N_22777,N_20266);
nor U28879 (N_28879,N_18236,N_22977);
or U28880 (N_28880,N_23555,N_19463);
or U28881 (N_28881,N_23658,N_21025);
nor U28882 (N_28882,N_21136,N_22416);
nor U28883 (N_28883,N_20416,N_18395);
nand U28884 (N_28884,N_20869,N_23064);
or U28885 (N_28885,N_19844,N_20575);
nor U28886 (N_28886,N_19971,N_20006);
nand U28887 (N_28887,N_21184,N_21929);
nor U28888 (N_28888,N_20947,N_19478);
and U28889 (N_28889,N_20829,N_20039);
or U28890 (N_28890,N_22963,N_23523);
xor U28891 (N_28891,N_19812,N_19610);
xnor U28892 (N_28892,N_20727,N_21928);
or U28893 (N_28893,N_22385,N_22641);
and U28894 (N_28894,N_21124,N_18974);
nor U28895 (N_28895,N_23550,N_20306);
or U28896 (N_28896,N_22598,N_23116);
or U28897 (N_28897,N_21370,N_18896);
and U28898 (N_28898,N_21349,N_21435);
nor U28899 (N_28899,N_20117,N_23707);
nor U28900 (N_28900,N_18319,N_21018);
nand U28901 (N_28901,N_20780,N_19486);
or U28902 (N_28902,N_19181,N_20944);
and U28903 (N_28903,N_19241,N_18352);
and U28904 (N_28904,N_21349,N_19551);
nor U28905 (N_28905,N_23191,N_19730);
and U28906 (N_28906,N_22578,N_20457);
and U28907 (N_28907,N_19780,N_20685);
or U28908 (N_28908,N_18796,N_20440);
nand U28909 (N_28909,N_22730,N_22194);
nand U28910 (N_28910,N_20355,N_19264);
xor U28911 (N_28911,N_21402,N_19174);
nand U28912 (N_28912,N_21224,N_21229);
nor U28913 (N_28913,N_19810,N_23103);
xnor U28914 (N_28914,N_20684,N_20552);
nor U28915 (N_28915,N_21271,N_20031);
nor U28916 (N_28916,N_21059,N_20304);
and U28917 (N_28917,N_22873,N_22707);
or U28918 (N_28918,N_23824,N_18208);
or U28919 (N_28919,N_18999,N_21683);
or U28920 (N_28920,N_19524,N_18861);
nor U28921 (N_28921,N_20149,N_18145);
xnor U28922 (N_28922,N_22739,N_19757);
and U28923 (N_28923,N_23492,N_19580);
nor U28924 (N_28924,N_23797,N_23619);
and U28925 (N_28925,N_20420,N_22828);
or U28926 (N_28926,N_19924,N_23150);
and U28927 (N_28927,N_19232,N_21377);
or U28928 (N_28928,N_23763,N_20058);
and U28929 (N_28929,N_18460,N_21196);
nand U28930 (N_28930,N_21731,N_20046);
nand U28931 (N_28931,N_21789,N_18307);
or U28932 (N_28932,N_18108,N_21079);
or U28933 (N_28933,N_23470,N_21483);
nor U28934 (N_28934,N_23899,N_22131);
nand U28935 (N_28935,N_23028,N_19944);
xor U28936 (N_28936,N_22624,N_23270);
or U28937 (N_28937,N_22335,N_18163);
or U28938 (N_28938,N_19494,N_21225);
nor U28939 (N_28939,N_22451,N_23407);
or U28940 (N_28940,N_23697,N_19795);
xor U28941 (N_28941,N_19356,N_23608);
or U28942 (N_28942,N_19760,N_22741);
nor U28943 (N_28943,N_19032,N_19684);
or U28944 (N_28944,N_20391,N_18672);
nand U28945 (N_28945,N_19611,N_22383);
or U28946 (N_28946,N_20061,N_23854);
xor U28947 (N_28947,N_21157,N_22690);
nor U28948 (N_28948,N_19174,N_21556);
or U28949 (N_28949,N_23536,N_18505);
nand U28950 (N_28950,N_18779,N_22259);
nor U28951 (N_28951,N_18307,N_21586);
or U28952 (N_28952,N_21335,N_22099);
nand U28953 (N_28953,N_18338,N_19147);
or U28954 (N_28954,N_19328,N_21120);
nand U28955 (N_28955,N_18190,N_22708);
nand U28956 (N_28956,N_22655,N_20733);
and U28957 (N_28957,N_20945,N_20059);
and U28958 (N_28958,N_22856,N_22810);
or U28959 (N_28959,N_21107,N_23596);
and U28960 (N_28960,N_22441,N_23937);
nor U28961 (N_28961,N_19263,N_23648);
or U28962 (N_28962,N_23969,N_19443);
or U28963 (N_28963,N_20902,N_20173);
nor U28964 (N_28964,N_18926,N_23023);
or U28965 (N_28965,N_20152,N_19695);
or U28966 (N_28966,N_23530,N_19004);
or U28967 (N_28967,N_20239,N_18900);
nor U28968 (N_28968,N_22438,N_19424);
nor U28969 (N_28969,N_20861,N_18151);
nand U28970 (N_28970,N_21531,N_21827);
and U28971 (N_28971,N_20211,N_19068);
nand U28972 (N_28972,N_22590,N_19715);
or U28973 (N_28973,N_23652,N_19996);
nand U28974 (N_28974,N_21579,N_19552);
and U28975 (N_28975,N_19661,N_23798);
xnor U28976 (N_28976,N_23852,N_22643);
or U28977 (N_28977,N_19474,N_21024);
nor U28978 (N_28978,N_18459,N_21148);
and U28979 (N_28979,N_21827,N_22652);
nor U28980 (N_28980,N_18755,N_23260);
nor U28981 (N_28981,N_19022,N_18220);
or U28982 (N_28982,N_23629,N_21033);
or U28983 (N_28983,N_22967,N_23234);
and U28984 (N_28984,N_21213,N_18156);
nor U28985 (N_28985,N_21726,N_18342);
and U28986 (N_28986,N_18732,N_21503);
nand U28987 (N_28987,N_19339,N_20217);
nand U28988 (N_28988,N_23072,N_19344);
nor U28989 (N_28989,N_18520,N_20902);
and U28990 (N_28990,N_19395,N_19349);
or U28991 (N_28991,N_22399,N_20578);
or U28992 (N_28992,N_18421,N_20892);
nand U28993 (N_28993,N_21805,N_20529);
or U28994 (N_28994,N_20200,N_20283);
and U28995 (N_28995,N_19151,N_18565);
nor U28996 (N_28996,N_23568,N_20684);
nand U28997 (N_28997,N_19863,N_18903);
nand U28998 (N_28998,N_21618,N_19256);
or U28999 (N_28999,N_22572,N_21142);
nand U29000 (N_29000,N_19939,N_21892);
and U29001 (N_29001,N_21625,N_23206);
or U29002 (N_29002,N_20823,N_20765);
nor U29003 (N_29003,N_19436,N_19193);
xnor U29004 (N_29004,N_22944,N_18803);
nand U29005 (N_29005,N_22536,N_22307);
and U29006 (N_29006,N_23879,N_18859);
and U29007 (N_29007,N_19196,N_22530);
or U29008 (N_29008,N_22357,N_18195);
nor U29009 (N_29009,N_20808,N_18199);
and U29010 (N_29010,N_20417,N_20867);
and U29011 (N_29011,N_18698,N_21384);
nor U29012 (N_29012,N_20916,N_22665);
and U29013 (N_29013,N_22256,N_19261);
nand U29014 (N_29014,N_23501,N_20137);
nor U29015 (N_29015,N_22794,N_18321);
or U29016 (N_29016,N_21470,N_23782);
nand U29017 (N_29017,N_21085,N_21566);
and U29018 (N_29018,N_21565,N_22153);
nand U29019 (N_29019,N_19294,N_19529);
nor U29020 (N_29020,N_18400,N_23637);
or U29021 (N_29021,N_23293,N_19182);
nor U29022 (N_29022,N_18452,N_21431);
nor U29023 (N_29023,N_21124,N_20224);
or U29024 (N_29024,N_18295,N_18133);
or U29025 (N_29025,N_21396,N_20227);
xor U29026 (N_29026,N_21498,N_23440);
nor U29027 (N_29027,N_18127,N_20469);
and U29028 (N_29028,N_23187,N_18402);
nand U29029 (N_29029,N_20141,N_20003);
nand U29030 (N_29030,N_23130,N_20859);
nor U29031 (N_29031,N_18244,N_21852);
or U29032 (N_29032,N_23104,N_20592);
and U29033 (N_29033,N_22342,N_18543);
nor U29034 (N_29034,N_21019,N_19935);
xor U29035 (N_29035,N_22180,N_19212);
nand U29036 (N_29036,N_20748,N_22987);
xnor U29037 (N_29037,N_19526,N_22359);
xor U29038 (N_29038,N_19143,N_21079);
nor U29039 (N_29039,N_21050,N_20460);
xnor U29040 (N_29040,N_23256,N_22235);
xor U29041 (N_29041,N_18504,N_21381);
xnor U29042 (N_29042,N_23382,N_23250);
and U29043 (N_29043,N_22597,N_23971);
nor U29044 (N_29044,N_21748,N_19227);
nand U29045 (N_29045,N_23150,N_21601);
and U29046 (N_29046,N_22613,N_22806);
nand U29047 (N_29047,N_20507,N_21169);
and U29048 (N_29048,N_20558,N_20794);
nand U29049 (N_29049,N_23499,N_19062);
xor U29050 (N_29050,N_21478,N_19657);
nand U29051 (N_29051,N_21287,N_20461);
and U29052 (N_29052,N_18895,N_23093);
nand U29053 (N_29053,N_21440,N_22199);
nand U29054 (N_29054,N_21133,N_20648);
or U29055 (N_29055,N_23580,N_21142);
nor U29056 (N_29056,N_20837,N_20252);
nor U29057 (N_29057,N_19394,N_23046);
nor U29058 (N_29058,N_23689,N_18459);
nor U29059 (N_29059,N_21201,N_23584);
or U29060 (N_29060,N_22093,N_22316);
or U29061 (N_29061,N_21022,N_20469);
or U29062 (N_29062,N_22333,N_20520);
and U29063 (N_29063,N_19487,N_21077);
and U29064 (N_29064,N_21235,N_23982);
nor U29065 (N_29065,N_21232,N_18551);
or U29066 (N_29066,N_20560,N_20682);
and U29067 (N_29067,N_20104,N_21572);
xnor U29068 (N_29068,N_19218,N_23525);
nand U29069 (N_29069,N_19472,N_21207);
and U29070 (N_29070,N_18053,N_20830);
and U29071 (N_29071,N_20419,N_21734);
xnor U29072 (N_29072,N_22275,N_23758);
or U29073 (N_29073,N_19545,N_21963);
nand U29074 (N_29074,N_19470,N_22406);
nand U29075 (N_29075,N_21983,N_19015);
or U29076 (N_29076,N_23508,N_19955);
and U29077 (N_29077,N_21685,N_22120);
nor U29078 (N_29078,N_18073,N_22083);
or U29079 (N_29079,N_19183,N_18450);
or U29080 (N_29080,N_18325,N_23721);
nor U29081 (N_29081,N_20295,N_21168);
or U29082 (N_29082,N_22109,N_20229);
or U29083 (N_29083,N_23126,N_21450);
or U29084 (N_29084,N_23207,N_19122);
or U29085 (N_29085,N_18226,N_22015);
nand U29086 (N_29086,N_19293,N_21891);
and U29087 (N_29087,N_21826,N_18038);
and U29088 (N_29088,N_23804,N_21608);
and U29089 (N_29089,N_22024,N_23024);
or U29090 (N_29090,N_19368,N_18570);
and U29091 (N_29091,N_18072,N_22640);
nor U29092 (N_29092,N_23247,N_19034);
xnor U29093 (N_29093,N_18143,N_23095);
or U29094 (N_29094,N_18038,N_22955);
or U29095 (N_29095,N_18344,N_23177);
nand U29096 (N_29096,N_20613,N_18033);
nor U29097 (N_29097,N_23460,N_23033);
nand U29098 (N_29098,N_21702,N_23457);
xor U29099 (N_29099,N_22659,N_22769);
xnor U29100 (N_29100,N_18858,N_21467);
nor U29101 (N_29101,N_19080,N_18858);
or U29102 (N_29102,N_22869,N_23196);
nand U29103 (N_29103,N_20086,N_23505);
or U29104 (N_29104,N_20102,N_22907);
xor U29105 (N_29105,N_23808,N_23562);
and U29106 (N_29106,N_19365,N_19734);
and U29107 (N_29107,N_18963,N_23387);
and U29108 (N_29108,N_23845,N_18494);
nand U29109 (N_29109,N_23418,N_18523);
or U29110 (N_29110,N_18249,N_21542);
nand U29111 (N_29111,N_23651,N_19492);
nor U29112 (N_29112,N_18867,N_22506);
xnor U29113 (N_29113,N_18193,N_22099);
or U29114 (N_29114,N_20855,N_21053);
nand U29115 (N_29115,N_19897,N_20361);
nand U29116 (N_29116,N_18509,N_23703);
nor U29117 (N_29117,N_20973,N_22731);
and U29118 (N_29118,N_19714,N_23533);
xnor U29119 (N_29119,N_21687,N_19455);
and U29120 (N_29120,N_23833,N_20442);
or U29121 (N_29121,N_21864,N_20462);
nor U29122 (N_29122,N_23822,N_21925);
or U29123 (N_29123,N_18365,N_22635);
and U29124 (N_29124,N_21248,N_19676);
or U29125 (N_29125,N_19808,N_22021);
and U29126 (N_29126,N_21182,N_20480);
and U29127 (N_29127,N_19908,N_20999);
xnor U29128 (N_29128,N_22757,N_22107);
or U29129 (N_29129,N_22345,N_21634);
nand U29130 (N_29130,N_21616,N_19274);
or U29131 (N_29131,N_21475,N_20120);
nand U29132 (N_29132,N_23599,N_21857);
or U29133 (N_29133,N_19058,N_21342);
or U29134 (N_29134,N_19311,N_19129);
or U29135 (N_29135,N_19804,N_20220);
nor U29136 (N_29136,N_23646,N_19055);
nand U29137 (N_29137,N_21040,N_22887);
and U29138 (N_29138,N_22829,N_20878);
nor U29139 (N_29139,N_18758,N_22126);
xnor U29140 (N_29140,N_22088,N_22501);
xnor U29141 (N_29141,N_22106,N_22827);
nor U29142 (N_29142,N_20218,N_20855);
nand U29143 (N_29143,N_21308,N_23604);
and U29144 (N_29144,N_23608,N_19902);
and U29145 (N_29145,N_23007,N_19895);
xnor U29146 (N_29146,N_23205,N_21336);
or U29147 (N_29147,N_22594,N_18861);
nor U29148 (N_29148,N_19325,N_22676);
nand U29149 (N_29149,N_22414,N_19608);
xor U29150 (N_29150,N_21701,N_18280);
or U29151 (N_29151,N_18817,N_21324);
and U29152 (N_29152,N_20807,N_21546);
xor U29153 (N_29153,N_20714,N_19822);
nand U29154 (N_29154,N_18555,N_21224);
nand U29155 (N_29155,N_20316,N_19942);
xnor U29156 (N_29156,N_22037,N_20074);
and U29157 (N_29157,N_18047,N_23791);
or U29158 (N_29158,N_19246,N_18027);
nand U29159 (N_29159,N_22826,N_18248);
nor U29160 (N_29160,N_18624,N_23593);
xor U29161 (N_29161,N_20207,N_21703);
nor U29162 (N_29162,N_21869,N_20612);
nor U29163 (N_29163,N_18981,N_20713);
nor U29164 (N_29164,N_23984,N_20600);
and U29165 (N_29165,N_22119,N_20473);
and U29166 (N_29166,N_18556,N_20775);
nor U29167 (N_29167,N_20583,N_18747);
or U29168 (N_29168,N_19989,N_18354);
nor U29169 (N_29169,N_21137,N_21258);
nand U29170 (N_29170,N_18061,N_22555);
or U29171 (N_29171,N_23368,N_23416);
nor U29172 (N_29172,N_22881,N_19636);
nor U29173 (N_29173,N_22183,N_23226);
and U29174 (N_29174,N_22096,N_19773);
nand U29175 (N_29175,N_21512,N_20804);
or U29176 (N_29176,N_21109,N_19069);
nand U29177 (N_29177,N_18935,N_18794);
and U29178 (N_29178,N_21392,N_19098);
nand U29179 (N_29179,N_18421,N_20973);
or U29180 (N_29180,N_22883,N_21282);
nor U29181 (N_29181,N_20381,N_20900);
and U29182 (N_29182,N_23135,N_20946);
or U29183 (N_29183,N_23335,N_21961);
nand U29184 (N_29184,N_18465,N_22278);
xor U29185 (N_29185,N_21879,N_21631);
nor U29186 (N_29186,N_20028,N_22970);
nand U29187 (N_29187,N_19604,N_18772);
or U29188 (N_29188,N_20471,N_22897);
xor U29189 (N_29189,N_23287,N_22583);
xor U29190 (N_29190,N_22413,N_23213);
nor U29191 (N_29191,N_21731,N_23053);
nand U29192 (N_29192,N_23021,N_21969);
or U29193 (N_29193,N_19776,N_22058);
nor U29194 (N_29194,N_22409,N_21540);
xor U29195 (N_29195,N_19703,N_23218);
nand U29196 (N_29196,N_19402,N_19685);
nand U29197 (N_29197,N_20626,N_23445);
nor U29198 (N_29198,N_18415,N_20920);
nand U29199 (N_29199,N_21235,N_19935);
nor U29200 (N_29200,N_18991,N_23082);
and U29201 (N_29201,N_21483,N_22293);
nor U29202 (N_29202,N_22276,N_18420);
or U29203 (N_29203,N_18455,N_20317);
nor U29204 (N_29204,N_18893,N_22048);
nand U29205 (N_29205,N_19029,N_18264);
nand U29206 (N_29206,N_20926,N_23064);
or U29207 (N_29207,N_22515,N_23240);
nor U29208 (N_29208,N_19961,N_23043);
and U29209 (N_29209,N_21865,N_23814);
and U29210 (N_29210,N_20115,N_22670);
nand U29211 (N_29211,N_23241,N_22438);
or U29212 (N_29212,N_19995,N_19167);
or U29213 (N_29213,N_21546,N_23977);
nand U29214 (N_29214,N_19953,N_20136);
nor U29215 (N_29215,N_23092,N_23459);
nor U29216 (N_29216,N_23474,N_19740);
and U29217 (N_29217,N_18302,N_20167);
nand U29218 (N_29218,N_22227,N_23421);
nor U29219 (N_29219,N_23092,N_20506);
nand U29220 (N_29220,N_19989,N_19320);
nor U29221 (N_29221,N_22212,N_19532);
or U29222 (N_29222,N_22437,N_18803);
nand U29223 (N_29223,N_21774,N_22743);
xnor U29224 (N_29224,N_18701,N_22603);
and U29225 (N_29225,N_22258,N_22828);
nand U29226 (N_29226,N_23398,N_20541);
and U29227 (N_29227,N_23319,N_23594);
and U29228 (N_29228,N_21550,N_20836);
or U29229 (N_29229,N_22446,N_23635);
or U29230 (N_29230,N_19309,N_19041);
or U29231 (N_29231,N_21211,N_21683);
nand U29232 (N_29232,N_18238,N_20882);
and U29233 (N_29233,N_21798,N_19834);
nor U29234 (N_29234,N_21788,N_22969);
nor U29235 (N_29235,N_19830,N_18966);
or U29236 (N_29236,N_21341,N_20304);
nor U29237 (N_29237,N_23286,N_20370);
and U29238 (N_29238,N_18170,N_20402);
nand U29239 (N_29239,N_22347,N_19186);
nand U29240 (N_29240,N_20289,N_21912);
nor U29241 (N_29241,N_19369,N_21992);
and U29242 (N_29242,N_18163,N_20039);
nor U29243 (N_29243,N_19190,N_19351);
and U29244 (N_29244,N_23896,N_23224);
nor U29245 (N_29245,N_18200,N_20769);
and U29246 (N_29246,N_22240,N_19921);
nand U29247 (N_29247,N_22266,N_20572);
and U29248 (N_29248,N_22937,N_19848);
and U29249 (N_29249,N_20461,N_19132);
nand U29250 (N_29250,N_20197,N_23496);
and U29251 (N_29251,N_19215,N_22533);
and U29252 (N_29252,N_22522,N_19641);
nor U29253 (N_29253,N_19834,N_20802);
and U29254 (N_29254,N_21026,N_20360);
xor U29255 (N_29255,N_23835,N_21460);
or U29256 (N_29256,N_19653,N_19690);
and U29257 (N_29257,N_19068,N_21934);
nand U29258 (N_29258,N_23552,N_20923);
nor U29259 (N_29259,N_23388,N_18808);
or U29260 (N_29260,N_21885,N_23325);
and U29261 (N_29261,N_21968,N_18960);
nor U29262 (N_29262,N_18695,N_23256);
nor U29263 (N_29263,N_19129,N_23109);
and U29264 (N_29264,N_21488,N_23741);
or U29265 (N_29265,N_20986,N_18943);
and U29266 (N_29266,N_22238,N_20944);
or U29267 (N_29267,N_23749,N_23439);
or U29268 (N_29268,N_20266,N_20772);
or U29269 (N_29269,N_18652,N_20595);
and U29270 (N_29270,N_23829,N_20952);
and U29271 (N_29271,N_23580,N_20178);
nand U29272 (N_29272,N_19127,N_23595);
nor U29273 (N_29273,N_19912,N_22125);
nor U29274 (N_29274,N_23807,N_22072);
xnor U29275 (N_29275,N_22513,N_18806);
or U29276 (N_29276,N_18549,N_19799);
or U29277 (N_29277,N_20152,N_22090);
and U29278 (N_29278,N_20412,N_20369);
nor U29279 (N_29279,N_19435,N_23184);
nor U29280 (N_29280,N_19735,N_21228);
nor U29281 (N_29281,N_22691,N_22933);
nand U29282 (N_29282,N_21538,N_20293);
or U29283 (N_29283,N_20507,N_18278);
xnor U29284 (N_29284,N_23503,N_19512);
nor U29285 (N_29285,N_19381,N_19007);
and U29286 (N_29286,N_21901,N_21608);
and U29287 (N_29287,N_20238,N_20096);
or U29288 (N_29288,N_18252,N_19420);
nand U29289 (N_29289,N_20510,N_22496);
and U29290 (N_29290,N_22921,N_19892);
and U29291 (N_29291,N_18147,N_19649);
or U29292 (N_29292,N_22101,N_19202);
or U29293 (N_29293,N_21980,N_23673);
nor U29294 (N_29294,N_20103,N_22671);
or U29295 (N_29295,N_23032,N_21263);
or U29296 (N_29296,N_20606,N_19807);
nand U29297 (N_29297,N_18436,N_18953);
and U29298 (N_29298,N_20941,N_23207);
nor U29299 (N_29299,N_23113,N_20851);
or U29300 (N_29300,N_22393,N_22356);
nand U29301 (N_29301,N_18906,N_20281);
nor U29302 (N_29302,N_20414,N_21042);
nor U29303 (N_29303,N_18539,N_19551);
nor U29304 (N_29304,N_20277,N_23642);
and U29305 (N_29305,N_22983,N_23891);
nand U29306 (N_29306,N_18465,N_22350);
or U29307 (N_29307,N_20711,N_19828);
xnor U29308 (N_29308,N_20861,N_21581);
nor U29309 (N_29309,N_20346,N_21942);
and U29310 (N_29310,N_19275,N_19657);
and U29311 (N_29311,N_23762,N_19840);
or U29312 (N_29312,N_18610,N_19254);
and U29313 (N_29313,N_20627,N_19604);
or U29314 (N_29314,N_22139,N_18973);
nand U29315 (N_29315,N_18418,N_22203);
and U29316 (N_29316,N_23881,N_18146);
nor U29317 (N_29317,N_23584,N_21309);
or U29318 (N_29318,N_18825,N_19109);
or U29319 (N_29319,N_19077,N_23374);
nor U29320 (N_29320,N_18835,N_22947);
nor U29321 (N_29321,N_23223,N_19662);
nand U29322 (N_29322,N_23931,N_22105);
nand U29323 (N_29323,N_23323,N_21949);
xor U29324 (N_29324,N_19434,N_18440);
nand U29325 (N_29325,N_18834,N_19190);
nor U29326 (N_29326,N_18524,N_22407);
or U29327 (N_29327,N_19533,N_18795);
nor U29328 (N_29328,N_19435,N_19833);
nand U29329 (N_29329,N_22676,N_18480);
nand U29330 (N_29330,N_23820,N_18286);
xnor U29331 (N_29331,N_19473,N_22701);
or U29332 (N_29332,N_18261,N_18883);
nand U29333 (N_29333,N_18887,N_22688);
nor U29334 (N_29334,N_19786,N_23155);
nor U29335 (N_29335,N_23832,N_18939);
or U29336 (N_29336,N_20791,N_20291);
or U29337 (N_29337,N_20824,N_23221);
nor U29338 (N_29338,N_22443,N_22305);
nand U29339 (N_29339,N_22580,N_19099);
and U29340 (N_29340,N_20621,N_18029);
or U29341 (N_29341,N_22532,N_18728);
nor U29342 (N_29342,N_22673,N_20393);
nand U29343 (N_29343,N_20504,N_21493);
nand U29344 (N_29344,N_22886,N_21328);
or U29345 (N_29345,N_21431,N_20812);
or U29346 (N_29346,N_19520,N_23622);
xor U29347 (N_29347,N_23297,N_19280);
and U29348 (N_29348,N_21883,N_23148);
nand U29349 (N_29349,N_21363,N_18289);
or U29350 (N_29350,N_18357,N_18263);
and U29351 (N_29351,N_19737,N_23742);
nor U29352 (N_29352,N_23907,N_21677);
nor U29353 (N_29353,N_22549,N_22845);
nor U29354 (N_29354,N_23139,N_19604);
nand U29355 (N_29355,N_23622,N_21795);
nor U29356 (N_29356,N_18601,N_20280);
nor U29357 (N_29357,N_22102,N_22476);
nand U29358 (N_29358,N_18957,N_19120);
or U29359 (N_29359,N_22602,N_22696);
and U29360 (N_29360,N_20355,N_19614);
nand U29361 (N_29361,N_21309,N_19653);
or U29362 (N_29362,N_21980,N_19478);
nor U29363 (N_29363,N_21033,N_18064);
or U29364 (N_29364,N_23794,N_21848);
xor U29365 (N_29365,N_23389,N_22530);
or U29366 (N_29366,N_21705,N_23879);
or U29367 (N_29367,N_18354,N_20831);
nand U29368 (N_29368,N_21231,N_20569);
nor U29369 (N_29369,N_19465,N_19323);
xor U29370 (N_29370,N_20748,N_21554);
nor U29371 (N_29371,N_18447,N_21304);
nor U29372 (N_29372,N_21292,N_22578);
nand U29373 (N_29373,N_18362,N_19380);
nand U29374 (N_29374,N_19275,N_19173);
nand U29375 (N_29375,N_19451,N_23000);
nand U29376 (N_29376,N_21244,N_21879);
nor U29377 (N_29377,N_20789,N_20575);
or U29378 (N_29378,N_19404,N_19565);
or U29379 (N_29379,N_19574,N_18528);
nand U29380 (N_29380,N_21622,N_23204);
nand U29381 (N_29381,N_21057,N_21155);
and U29382 (N_29382,N_23553,N_20370);
nor U29383 (N_29383,N_18763,N_23786);
nor U29384 (N_29384,N_20935,N_20338);
or U29385 (N_29385,N_20230,N_21114);
and U29386 (N_29386,N_21698,N_18946);
nand U29387 (N_29387,N_19932,N_19397);
and U29388 (N_29388,N_18863,N_20217);
and U29389 (N_29389,N_18460,N_19315);
or U29390 (N_29390,N_19392,N_19064);
and U29391 (N_29391,N_21791,N_21010);
or U29392 (N_29392,N_21271,N_18371);
and U29393 (N_29393,N_21118,N_18161);
nor U29394 (N_29394,N_20967,N_22666);
nand U29395 (N_29395,N_23852,N_20423);
nand U29396 (N_29396,N_21988,N_20214);
nand U29397 (N_29397,N_18385,N_22795);
nor U29398 (N_29398,N_18236,N_18826);
nand U29399 (N_29399,N_22479,N_20780);
and U29400 (N_29400,N_21853,N_19332);
nor U29401 (N_29401,N_18504,N_18726);
or U29402 (N_29402,N_21992,N_19336);
xor U29403 (N_29403,N_21934,N_20624);
and U29404 (N_29404,N_19115,N_23876);
and U29405 (N_29405,N_19899,N_22520);
xnor U29406 (N_29406,N_22200,N_20950);
or U29407 (N_29407,N_23714,N_21992);
nor U29408 (N_29408,N_19582,N_22896);
and U29409 (N_29409,N_19462,N_18421);
and U29410 (N_29410,N_21787,N_23912);
or U29411 (N_29411,N_22732,N_18539);
xor U29412 (N_29412,N_21591,N_23861);
xor U29413 (N_29413,N_19581,N_22323);
xnor U29414 (N_29414,N_19021,N_19606);
nor U29415 (N_29415,N_20144,N_23011);
nor U29416 (N_29416,N_19166,N_19499);
nor U29417 (N_29417,N_20266,N_22218);
or U29418 (N_29418,N_18201,N_22727);
nor U29419 (N_29419,N_20645,N_19038);
and U29420 (N_29420,N_23521,N_23858);
or U29421 (N_29421,N_21574,N_18529);
nand U29422 (N_29422,N_21912,N_21167);
and U29423 (N_29423,N_23817,N_23057);
and U29424 (N_29424,N_22163,N_20709);
nand U29425 (N_29425,N_21703,N_23991);
and U29426 (N_29426,N_18023,N_19900);
and U29427 (N_29427,N_23973,N_22782);
and U29428 (N_29428,N_22732,N_19253);
nor U29429 (N_29429,N_21007,N_23723);
nor U29430 (N_29430,N_20258,N_18841);
or U29431 (N_29431,N_23912,N_20412);
or U29432 (N_29432,N_18766,N_23036);
nand U29433 (N_29433,N_21185,N_20617);
nand U29434 (N_29434,N_23878,N_22279);
nor U29435 (N_29435,N_23004,N_23710);
nor U29436 (N_29436,N_18582,N_22131);
nand U29437 (N_29437,N_22494,N_18008);
or U29438 (N_29438,N_20231,N_19324);
and U29439 (N_29439,N_21772,N_23445);
nand U29440 (N_29440,N_23413,N_18170);
and U29441 (N_29441,N_23707,N_19247);
or U29442 (N_29442,N_22916,N_21314);
and U29443 (N_29443,N_22055,N_18654);
nor U29444 (N_29444,N_20268,N_18766);
or U29445 (N_29445,N_20541,N_22572);
or U29446 (N_29446,N_21003,N_20135);
and U29447 (N_29447,N_23274,N_22065);
nor U29448 (N_29448,N_22315,N_22523);
and U29449 (N_29449,N_19587,N_19213);
or U29450 (N_29450,N_18482,N_22307);
nor U29451 (N_29451,N_22433,N_20438);
nor U29452 (N_29452,N_20345,N_23054);
or U29453 (N_29453,N_20182,N_23385);
or U29454 (N_29454,N_22940,N_20544);
nor U29455 (N_29455,N_22605,N_23981);
and U29456 (N_29456,N_22634,N_21275);
and U29457 (N_29457,N_20574,N_20546);
and U29458 (N_29458,N_21882,N_19049);
nor U29459 (N_29459,N_18586,N_21039);
or U29460 (N_29460,N_23522,N_22461);
and U29461 (N_29461,N_23692,N_20623);
or U29462 (N_29462,N_20078,N_20417);
and U29463 (N_29463,N_23269,N_22460);
or U29464 (N_29464,N_18952,N_23790);
and U29465 (N_29465,N_19919,N_22975);
nor U29466 (N_29466,N_18822,N_20832);
or U29467 (N_29467,N_19362,N_18766);
nand U29468 (N_29468,N_18251,N_23147);
nand U29469 (N_29469,N_18681,N_21467);
nand U29470 (N_29470,N_20309,N_20279);
nand U29471 (N_29471,N_21274,N_22033);
or U29472 (N_29472,N_20321,N_21758);
nand U29473 (N_29473,N_19441,N_23026);
xor U29474 (N_29474,N_20488,N_20512);
nor U29475 (N_29475,N_21791,N_18745);
nor U29476 (N_29476,N_23169,N_21605);
nand U29477 (N_29477,N_19833,N_23304);
or U29478 (N_29478,N_23008,N_18380);
and U29479 (N_29479,N_19212,N_19957);
nor U29480 (N_29480,N_22661,N_21641);
nor U29481 (N_29481,N_21311,N_23116);
nand U29482 (N_29482,N_20338,N_22584);
xor U29483 (N_29483,N_19709,N_21712);
nor U29484 (N_29484,N_20687,N_23377);
nand U29485 (N_29485,N_21044,N_22484);
xnor U29486 (N_29486,N_21165,N_20315);
nor U29487 (N_29487,N_23053,N_21752);
or U29488 (N_29488,N_19062,N_22231);
and U29489 (N_29489,N_23952,N_21046);
nor U29490 (N_29490,N_20351,N_19890);
nor U29491 (N_29491,N_22276,N_22076);
nand U29492 (N_29492,N_20343,N_23917);
nand U29493 (N_29493,N_22020,N_18246);
nand U29494 (N_29494,N_19478,N_23056);
nor U29495 (N_29495,N_22655,N_23171);
nand U29496 (N_29496,N_19965,N_18728);
nand U29497 (N_29497,N_23114,N_22022);
and U29498 (N_29498,N_22209,N_20341);
or U29499 (N_29499,N_23979,N_20204);
nor U29500 (N_29500,N_23005,N_20402);
nor U29501 (N_29501,N_18990,N_18744);
or U29502 (N_29502,N_18227,N_21637);
or U29503 (N_29503,N_23941,N_18074);
and U29504 (N_29504,N_23982,N_22174);
nor U29505 (N_29505,N_18382,N_22887);
or U29506 (N_29506,N_20784,N_21591);
nor U29507 (N_29507,N_18447,N_18874);
nor U29508 (N_29508,N_18765,N_19393);
or U29509 (N_29509,N_20165,N_21736);
and U29510 (N_29510,N_19992,N_21132);
nor U29511 (N_29511,N_18650,N_18720);
nand U29512 (N_29512,N_19979,N_20697);
nor U29513 (N_29513,N_23211,N_23380);
nor U29514 (N_29514,N_21373,N_19325);
xnor U29515 (N_29515,N_23473,N_22366);
nand U29516 (N_29516,N_22150,N_21775);
nor U29517 (N_29517,N_20323,N_22341);
or U29518 (N_29518,N_22068,N_22382);
nand U29519 (N_29519,N_23196,N_19320);
or U29520 (N_29520,N_20279,N_20708);
and U29521 (N_29521,N_22943,N_23111);
xnor U29522 (N_29522,N_18912,N_22177);
nand U29523 (N_29523,N_18753,N_18101);
or U29524 (N_29524,N_19603,N_22592);
and U29525 (N_29525,N_23048,N_20774);
and U29526 (N_29526,N_22959,N_19495);
and U29527 (N_29527,N_23888,N_22679);
and U29528 (N_29528,N_23396,N_20779);
nor U29529 (N_29529,N_21378,N_21452);
nor U29530 (N_29530,N_21494,N_22675);
and U29531 (N_29531,N_23155,N_19996);
nand U29532 (N_29532,N_23876,N_22078);
and U29533 (N_29533,N_19195,N_22581);
and U29534 (N_29534,N_18841,N_19117);
nand U29535 (N_29535,N_23714,N_22882);
nand U29536 (N_29536,N_20042,N_23220);
or U29537 (N_29537,N_21627,N_19045);
xor U29538 (N_29538,N_23702,N_21961);
and U29539 (N_29539,N_23935,N_18882);
nand U29540 (N_29540,N_18530,N_18825);
and U29541 (N_29541,N_20755,N_21849);
and U29542 (N_29542,N_21677,N_20321);
nor U29543 (N_29543,N_22155,N_21256);
nor U29544 (N_29544,N_18852,N_22606);
nor U29545 (N_29545,N_21743,N_21678);
nand U29546 (N_29546,N_21437,N_23273);
and U29547 (N_29547,N_19924,N_20112);
nor U29548 (N_29548,N_18591,N_23185);
and U29549 (N_29549,N_23416,N_18048);
and U29550 (N_29550,N_21319,N_20484);
nand U29551 (N_29551,N_21345,N_20502);
or U29552 (N_29552,N_23442,N_21624);
nand U29553 (N_29553,N_23922,N_22175);
nand U29554 (N_29554,N_23587,N_22814);
or U29555 (N_29555,N_20247,N_18242);
xnor U29556 (N_29556,N_19086,N_21047);
xnor U29557 (N_29557,N_23430,N_21981);
or U29558 (N_29558,N_22795,N_20752);
nand U29559 (N_29559,N_23440,N_20252);
nand U29560 (N_29560,N_20016,N_21176);
xnor U29561 (N_29561,N_18376,N_20263);
or U29562 (N_29562,N_18198,N_20819);
and U29563 (N_29563,N_23789,N_20607);
nor U29564 (N_29564,N_21985,N_19151);
nand U29565 (N_29565,N_23250,N_20065);
and U29566 (N_29566,N_18802,N_21045);
nor U29567 (N_29567,N_19697,N_20671);
or U29568 (N_29568,N_18935,N_23449);
nor U29569 (N_29569,N_22409,N_23397);
and U29570 (N_29570,N_19193,N_21116);
xor U29571 (N_29571,N_18393,N_23761);
or U29572 (N_29572,N_22107,N_22911);
and U29573 (N_29573,N_23237,N_18215);
nand U29574 (N_29574,N_21141,N_23920);
or U29575 (N_29575,N_19165,N_18000);
xor U29576 (N_29576,N_23514,N_22820);
and U29577 (N_29577,N_21784,N_23306);
nand U29578 (N_29578,N_18908,N_20174);
nand U29579 (N_29579,N_21107,N_20308);
and U29580 (N_29580,N_18154,N_20156);
or U29581 (N_29581,N_19080,N_19611);
nor U29582 (N_29582,N_19724,N_21205);
nor U29583 (N_29583,N_20542,N_20213);
or U29584 (N_29584,N_21540,N_21061);
nor U29585 (N_29585,N_23714,N_18703);
and U29586 (N_29586,N_21484,N_22878);
nand U29587 (N_29587,N_20927,N_22817);
nor U29588 (N_29588,N_23414,N_19534);
nand U29589 (N_29589,N_23856,N_22118);
xnor U29590 (N_29590,N_19499,N_22960);
and U29591 (N_29591,N_19815,N_20118);
nand U29592 (N_29592,N_23316,N_19558);
or U29593 (N_29593,N_22749,N_20988);
nand U29594 (N_29594,N_19137,N_21493);
or U29595 (N_29595,N_22507,N_19366);
and U29596 (N_29596,N_18106,N_20837);
or U29597 (N_29597,N_19491,N_22469);
xnor U29598 (N_29598,N_23179,N_21768);
nand U29599 (N_29599,N_19168,N_21506);
xor U29600 (N_29600,N_22904,N_22190);
or U29601 (N_29601,N_21571,N_22502);
nand U29602 (N_29602,N_22043,N_22917);
nand U29603 (N_29603,N_19490,N_21923);
nand U29604 (N_29604,N_22510,N_19510);
nand U29605 (N_29605,N_21929,N_20642);
nand U29606 (N_29606,N_21256,N_18405);
and U29607 (N_29607,N_21839,N_22981);
or U29608 (N_29608,N_18856,N_22312);
or U29609 (N_29609,N_21502,N_21223);
and U29610 (N_29610,N_23253,N_23275);
and U29611 (N_29611,N_21002,N_19603);
and U29612 (N_29612,N_18211,N_19255);
nor U29613 (N_29613,N_19827,N_20950);
nand U29614 (N_29614,N_23562,N_22241);
xnor U29615 (N_29615,N_20104,N_19491);
nor U29616 (N_29616,N_20895,N_18330);
and U29617 (N_29617,N_20610,N_22310);
and U29618 (N_29618,N_21509,N_22998);
and U29619 (N_29619,N_22998,N_21470);
nand U29620 (N_29620,N_21849,N_23468);
nand U29621 (N_29621,N_19850,N_23009);
nand U29622 (N_29622,N_22655,N_21864);
nand U29623 (N_29623,N_21938,N_22208);
nor U29624 (N_29624,N_22173,N_22639);
or U29625 (N_29625,N_23550,N_22214);
nand U29626 (N_29626,N_18173,N_18167);
nor U29627 (N_29627,N_19392,N_21803);
nor U29628 (N_29628,N_23479,N_21971);
xnor U29629 (N_29629,N_18996,N_23158);
and U29630 (N_29630,N_19679,N_18452);
nand U29631 (N_29631,N_19330,N_19482);
or U29632 (N_29632,N_23295,N_18375);
nor U29633 (N_29633,N_23601,N_18433);
nand U29634 (N_29634,N_19141,N_22091);
nor U29635 (N_29635,N_23883,N_21257);
nand U29636 (N_29636,N_23110,N_21485);
nor U29637 (N_29637,N_21835,N_21470);
nor U29638 (N_29638,N_23237,N_22136);
nor U29639 (N_29639,N_21589,N_20117);
nand U29640 (N_29640,N_21952,N_19690);
and U29641 (N_29641,N_20004,N_18843);
or U29642 (N_29642,N_23845,N_18386);
nand U29643 (N_29643,N_21581,N_21107);
nand U29644 (N_29644,N_23961,N_20813);
nor U29645 (N_29645,N_18414,N_18891);
and U29646 (N_29646,N_19215,N_21206);
or U29647 (N_29647,N_21353,N_22305);
xor U29648 (N_29648,N_19124,N_22931);
nor U29649 (N_29649,N_22482,N_21672);
xor U29650 (N_29650,N_18091,N_22808);
nor U29651 (N_29651,N_23550,N_23061);
and U29652 (N_29652,N_21203,N_22187);
and U29653 (N_29653,N_23687,N_18003);
nor U29654 (N_29654,N_21542,N_22774);
or U29655 (N_29655,N_22861,N_18357);
nand U29656 (N_29656,N_18643,N_19591);
and U29657 (N_29657,N_23701,N_20352);
xor U29658 (N_29658,N_22526,N_23639);
nand U29659 (N_29659,N_18174,N_23860);
or U29660 (N_29660,N_22490,N_21736);
or U29661 (N_29661,N_18315,N_23187);
nand U29662 (N_29662,N_18115,N_18732);
nand U29663 (N_29663,N_21405,N_20608);
or U29664 (N_29664,N_23778,N_23707);
nor U29665 (N_29665,N_18553,N_18965);
nor U29666 (N_29666,N_21136,N_23473);
nor U29667 (N_29667,N_23343,N_18240);
nor U29668 (N_29668,N_20598,N_22562);
nor U29669 (N_29669,N_18837,N_19206);
or U29670 (N_29670,N_20959,N_20504);
or U29671 (N_29671,N_18163,N_20092);
nor U29672 (N_29672,N_18592,N_22788);
or U29673 (N_29673,N_23679,N_21421);
and U29674 (N_29674,N_20569,N_20402);
and U29675 (N_29675,N_23293,N_19055);
or U29676 (N_29676,N_21714,N_18874);
and U29677 (N_29677,N_21304,N_18042);
nor U29678 (N_29678,N_21043,N_19085);
nor U29679 (N_29679,N_20266,N_21062);
nand U29680 (N_29680,N_19766,N_18124);
xor U29681 (N_29681,N_23645,N_23464);
nand U29682 (N_29682,N_18862,N_23526);
or U29683 (N_29683,N_18266,N_20593);
and U29684 (N_29684,N_19105,N_22278);
or U29685 (N_29685,N_20405,N_21010);
and U29686 (N_29686,N_20096,N_21958);
and U29687 (N_29687,N_19216,N_19059);
nand U29688 (N_29688,N_22453,N_19167);
xnor U29689 (N_29689,N_23851,N_20211);
and U29690 (N_29690,N_19058,N_21755);
nor U29691 (N_29691,N_23096,N_22295);
and U29692 (N_29692,N_18680,N_19898);
or U29693 (N_29693,N_23139,N_23565);
or U29694 (N_29694,N_23943,N_19807);
nand U29695 (N_29695,N_19110,N_19855);
or U29696 (N_29696,N_23690,N_19629);
nand U29697 (N_29697,N_23705,N_22539);
nor U29698 (N_29698,N_19257,N_19353);
or U29699 (N_29699,N_21469,N_22099);
nand U29700 (N_29700,N_19851,N_19211);
or U29701 (N_29701,N_23993,N_21447);
nor U29702 (N_29702,N_23976,N_22235);
nand U29703 (N_29703,N_19475,N_22463);
nor U29704 (N_29704,N_20240,N_19071);
nor U29705 (N_29705,N_22243,N_20353);
and U29706 (N_29706,N_23914,N_22042);
nand U29707 (N_29707,N_18417,N_21898);
nor U29708 (N_29708,N_19713,N_19497);
or U29709 (N_29709,N_18172,N_19155);
nor U29710 (N_29710,N_21774,N_18663);
and U29711 (N_29711,N_21334,N_20587);
or U29712 (N_29712,N_23185,N_18674);
nor U29713 (N_29713,N_23389,N_21498);
nor U29714 (N_29714,N_22049,N_19349);
nand U29715 (N_29715,N_21297,N_22916);
or U29716 (N_29716,N_22830,N_23849);
and U29717 (N_29717,N_22676,N_18185);
nor U29718 (N_29718,N_18171,N_21002);
xor U29719 (N_29719,N_23149,N_21114);
nand U29720 (N_29720,N_20261,N_19329);
and U29721 (N_29721,N_22028,N_21337);
nor U29722 (N_29722,N_18716,N_19880);
and U29723 (N_29723,N_22085,N_21734);
or U29724 (N_29724,N_18365,N_22357);
nor U29725 (N_29725,N_20044,N_20556);
or U29726 (N_29726,N_18622,N_21751);
and U29727 (N_29727,N_22119,N_22288);
or U29728 (N_29728,N_18381,N_19908);
nor U29729 (N_29729,N_22839,N_21057);
or U29730 (N_29730,N_21510,N_22671);
or U29731 (N_29731,N_23845,N_21529);
or U29732 (N_29732,N_21616,N_23719);
xnor U29733 (N_29733,N_20959,N_18760);
or U29734 (N_29734,N_19359,N_22867);
xnor U29735 (N_29735,N_19401,N_21039);
xor U29736 (N_29736,N_20564,N_18783);
and U29737 (N_29737,N_20622,N_22758);
or U29738 (N_29738,N_18205,N_23484);
nand U29739 (N_29739,N_23901,N_20013);
nand U29740 (N_29740,N_18005,N_21822);
or U29741 (N_29741,N_21005,N_18018);
xor U29742 (N_29742,N_18502,N_20053);
nor U29743 (N_29743,N_18674,N_20773);
or U29744 (N_29744,N_20142,N_19090);
or U29745 (N_29745,N_23311,N_19570);
nand U29746 (N_29746,N_23791,N_22124);
or U29747 (N_29747,N_21484,N_19551);
nand U29748 (N_29748,N_21942,N_21230);
xor U29749 (N_29749,N_20875,N_23270);
and U29750 (N_29750,N_20742,N_19959);
nand U29751 (N_29751,N_20227,N_18439);
nand U29752 (N_29752,N_19783,N_20536);
or U29753 (N_29753,N_18223,N_19568);
nand U29754 (N_29754,N_23004,N_23992);
or U29755 (N_29755,N_21004,N_22306);
nor U29756 (N_29756,N_22667,N_21866);
and U29757 (N_29757,N_18810,N_23870);
or U29758 (N_29758,N_18990,N_19412);
xnor U29759 (N_29759,N_20616,N_21324);
xor U29760 (N_29760,N_19863,N_19128);
xor U29761 (N_29761,N_21771,N_21071);
and U29762 (N_29762,N_19758,N_20723);
nand U29763 (N_29763,N_18185,N_22666);
or U29764 (N_29764,N_18712,N_21504);
and U29765 (N_29765,N_23654,N_18214);
and U29766 (N_29766,N_21186,N_21475);
nand U29767 (N_29767,N_23215,N_19664);
and U29768 (N_29768,N_21591,N_20249);
or U29769 (N_29769,N_23795,N_23948);
or U29770 (N_29770,N_20313,N_19834);
and U29771 (N_29771,N_22071,N_21797);
nor U29772 (N_29772,N_18567,N_22880);
nor U29773 (N_29773,N_21469,N_19778);
nor U29774 (N_29774,N_19086,N_21937);
nor U29775 (N_29775,N_23701,N_22182);
and U29776 (N_29776,N_23521,N_23457);
nor U29777 (N_29777,N_22777,N_22078);
or U29778 (N_29778,N_23015,N_22070);
and U29779 (N_29779,N_21754,N_20340);
xor U29780 (N_29780,N_23074,N_21851);
nor U29781 (N_29781,N_21122,N_21773);
nand U29782 (N_29782,N_18243,N_22805);
nor U29783 (N_29783,N_20280,N_19919);
or U29784 (N_29784,N_22018,N_22334);
or U29785 (N_29785,N_21584,N_21842);
xor U29786 (N_29786,N_19107,N_21661);
and U29787 (N_29787,N_23802,N_22741);
nand U29788 (N_29788,N_23513,N_18107);
or U29789 (N_29789,N_18449,N_23144);
nand U29790 (N_29790,N_20895,N_19071);
nor U29791 (N_29791,N_21752,N_23251);
and U29792 (N_29792,N_23530,N_22430);
nand U29793 (N_29793,N_22475,N_18991);
or U29794 (N_29794,N_22313,N_20643);
nor U29795 (N_29795,N_22353,N_23978);
or U29796 (N_29796,N_22274,N_23256);
nor U29797 (N_29797,N_20957,N_22467);
or U29798 (N_29798,N_21494,N_19228);
nand U29799 (N_29799,N_21320,N_22460);
nor U29800 (N_29800,N_22745,N_20257);
nand U29801 (N_29801,N_22715,N_20606);
xnor U29802 (N_29802,N_23426,N_18664);
or U29803 (N_29803,N_22723,N_23728);
nand U29804 (N_29804,N_21313,N_19942);
nor U29805 (N_29805,N_20435,N_19445);
xnor U29806 (N_29806,N_19930,N_21429);
and U29807 (N_29807,N_19644,N_22656);
or U29808 (N_29808,N_23396,N_21522);
xor U29809 (N_29809,N_20618,N_19380);
or U29810 (N_29810,N_20349,N_21712);
nand U29811 (N_29811,N_18393,N_23507);
and U29812 (N_29812,N_23740,N_23552);
and U29813 (N_29813,N_21541,N_20795);
or U29814 (N_29814,N_21538,N_23043);
or U29815 (N_29815,N_18668,N_23926);
or U29816 (N_29816,N_21596,N_21058);
nand U29817 (N_29817,N_18335,N_19495);
nor U29818 (N_29818,N_20143,N_23878);
and U29819 (N_29819,N_20989,N_23974);
xor U29820 (N_29820,N_20809,N_23495);
nand U29821 (N_29821,N_20056,N_19239);
and U29822 (N_29822,N_19105,N_21712);
nand U29823 (N_29823,N_20728,N_22408);
nor U29824 (N_29824,N_22362,N_22909);
or U29825 (N_29825,N_23149,N_19049);
nand U29826 (N_29826,N_23807,N_19597);
or U29827 (N_29827,N_23541,N_20055);
nor U29828 (N_29828,N_18978,N_18448);
and U29829 (N_29829,N_23200,N_20142);
or U29830 (N_29830,N_20857,N_22780);
or U29831 (N_29831,N_20602,N_23017);
xor U29832 (N_29832,N_19662,N_23960);
or U29833 (N_29833,N_20007,N_23178);
or U29834 (N_29834,N_19779,N_21999);
and U29835 (N_29835,N_19087,N_19237);
nand U29836 (N_29836,N_20811,N_18613);
or U29837 (N_29837,N_23945,N_18620);
nor U29838 (N_29838,N_20365,N_19178);
or U29839 (N_29839,N_23846,N_22850);
nor U29840 (N_29840,N_21680,N_21177);
or U29841 (N_29841,N_22634,N_22881);
nor U29842 (N_29842,N_22541,N_20309);
nor U29843 (N_29843,N_21411,N_20779);
nand U29844 (N_29844,N_20134,N_22406);
nand U29845 (N_29845,N_23511,N_19523);
or U29846 (N_29846,N_19823,N_20138);
nand U29847 (N_29847,N_19508,N_19955);
nand U29848 (N_29848,N_19273,N_21284);
nand U29849 (N_29849,N_19004,N_20170);
nor U29850 (N_29850,N_23764,N_23448);
nor U29851 (N_29851,N_21159,N_23398);
nor U29852 (N_29852,N_20377,N_19732);
nor U29853 (N_29853,N_20504,N_21688);
xor U29854 (N_29854,N_22583,N_22609);
xnor U29855 (N_29855,N_20669,N_21108);
nand U29856 (N_29856,N_20804,N_18427);
nor U29857 (N_29857,N_21509,N_18214);
or U29858 (N_29858,N_23775,N_21061);
and U29859 (N_29859,N_20092,N_20848);
nand U29860 (N_29860,N_20684,N_18317);
nor U29861 (N_29861,N_18005,N_18519);
xnor U29862 (N_29862,N_21804,N_18351);
nor U29863 (N_29863,N_21009,N_22660);
and U29864 (N_29864,N_21583,N_22189);
and U29865 (N_29865,N_22268,N_18589);
nor U29866 (N_29866,N_22911,N_19174);
nand U29867 (N_29867,N_18590,N_19814);
nand U29868 (N_29868,N_23107,N_22265);
nand U29869 (N_29869,N_18191,N_18888);
and U29870 (N_29870,N_19716,N_18021);
or U29871 (N_29871,N_21171,N_21665);
nor U29872 (N_29872,N_18382,N_21552);
nor U29873 (N_29873,N_21232,N_23970);
nand U29874 (N_29874,N_21296,N_18450);
or U29875 (N_29875,N_22587,N_20067);
xor U29876 (N_29876,N_20530,N_19454);
or U29877 (N_29877,N_18101,N_18324);
nor U29878 (N_29878,N_19128,N_23498);
or U29879 (N_29879,N_19652,N_19038);
nand U29880 (N_29880,N_18252,N_21216);
xnor U29881 (N_29881,N_22997,N_20803);
and U29882 (N_29882,N_18013,N_20069);
or U29883 (N_29883,N_21758,N_21050);
nor U29884 (N_29884,N_20951,N_22719);
or U29885 (N_29885,N_22574,N_18676);
nor U29886 (N_29886,N_19647,N_21744);
and U29887 (N_29887,N_18490,N_23985);
or U29888 (N_29888,N_19336,N_20576);
nand U29889 (N_29889,N_23250,N_20229);
nand U29890 (N_29890,N_21271,N_22092);
and U29891 (N_29891,N_23888,N_18296);
and U29892 (N_29892,N_18295,N_23923);
or U29893 (N_29893,N_22849,N_21352);
and U29894 (N_29894,N_22262,N_19832);
and U29895 (N_29895,N_19540,N_19339);
or U29896 (N_29896,N_21154,N_18721);
nand U29897 (N_29897,N_19992,N_20261);
nor U29898 (N_29898,N_18115,N_21141);
nor U29899 (N_29899,N_18723,N_22625);
or U29900 (N_29900,N_18845,N_18882);
nand U29901 (N_29901,N_20823,N_19667);
nor U29902 (N_29902,N_18522,N_22685);
and U29903 (N_29903,N_21437,N_19736);
nand U29904 (N_29904,N_21839,N_22657);
nand U29905 (N_29905,N_21089,N_19362);
and U29906 (N_29906,N_20255,N_18155);
nor U29907 (N_29907,N_20992,N_18798);
nand U29908 (N_29908,N_18177,N_21939);
or U29909 (N_29909,N_20194,N_21204);
nor U29910 (N_29910,N_23779,N_22105);
nor U29911 (N_29911,N_20803,N_23493);
nor U29912 (N_29912,N_22031,N_22532);
or U29913 (N_29913,N_21366,N_19300);
and U29914 (N_29914,N_21739,N_23976);
nor U29915 (N_29915,N_23395,N_21711);
or U29916 (N_29916,N_19515,N_23226);
and U29917 (N_29917,N_22826,N_22503);
and U29918 (N_29918,N_21363,N_20803);
nor U29919 (N_29919,N_19307,N_23096);
nand U29920 (N_29920,N_23666,N_20024);
nand U29921 (N_29921,N_20176,N_22600);
nand U29922 (N_29922,N_23407,N_18147);
and U29923 (N_29923,N_21911,N_21565);
nand U29924 (N_29924,N_18402,N_23005);
nand U29925 (N_29925,N_23139,N_18087);
and U29926 (N_29926,N_23310,N_18232);
nor U29927 (N_29927,N_19445,N_21777);
xnor U29928 (N_29928,N_21255,N_22053);
and U29929 (N_29929,N_18198,N_19810);
nor U29930 (N_29930,N_18672,N_19644);
nand U29931 (N_29931,N_23537,N_23853);
or U29932 (N_29932,N_23801,N_19744);
nor U29933 (N_29933,N_19677,N_23824);
nor U29934 (N_29934,N_20490,N_22326);
nand U29935 (N_29935,N_22087,N_22478);
xor U29936 (N_29936,N_23676,N_19566);
nand U29937 (N_29937,N_21249,N_21279);
or U29938 (N_29938,N_18883,N_23136);
xnor U29939 (N_29939,N_21134,N_19863);
and U29940 (N_29940,N_18186,N_18129);
and U29941 (N_29941,N_19329,N_20337);
or U29942 (N_29942,N_19126,N_22527);
and U29943 (N_29943,N_18047,N_20632);
and U29944 (N_29944,N_18100,N_19550);
and U29945 (N_29945,N_23774,N_18848);
nand U29946 (N_29946,N_21197,N_19577);
or U29947 (N_29947,N_23601,N_22279);
nand U29948 (N_29948,N_22444,N_20562);
and U29949 (N_29949,N_20727,N_22285);
nand U29950 (N_29950,N_23931,N_22595);
nor U29951 (N_29951,N_23172,N_20121);
and U29952 (N_29952,N_22943,N_19123);
or U29953 (N_29953,N_23906,N_18632);
and U29954 (N_29954,N_20638,N_19507);
and U29955 (N_29955,N_21392,N_19813);
xnor U29956 (N_29956,N_23636,N_20058);
nand U29957 (N_29957,N_18225,N_22433);
nor U29958 (N_29958,N_20847,N_20284);
and U29959 (N_29959,N_23192,N_20542);
nand U29960 (N_29960,N_23185,N_20730);
or U29961 (N_29961,N_20107,N_20162);
nor U29962 (N_29962,N_22319,N_21128);
nor U29963 (N_29963,N_21049,N_18236);
nand U29964 (N_29964,N_18546,N_23279);
nor U29965 (N_29965,N_19683,N_19007);
or U29966 (N_29966,N_18328,N_20333);
nor U29967 (N_29967,N_21175,N_20565);
and U29968 (N_29968,N_21638,N_21944);
xnor U29969 (N_29969,N_18590,N_20250);
nand U29970 (N_29970,N_22488,N_22805);
and U29971 (N_29971,N_18339,N_19351);
nor U29972 (N_29972,N_23193,N_23895);
and U29973 (N_29973,N_21436,N_19591);
or U29974 (N_29974,N_18435,N_23658);
and U29975 (N_29975,N_18266,N_21227);
nor U29976 (N_29976,N_20828,N_19674);
nor U29977 (N_29977,N_20237,N_20401);
nor U29978 (N_29978,N_22530,N_22593);
or U29979 (N_29979,N_22838,N_19593);
nor U29980 (N_29980,N_23883,N_23191);
nand U29981 (N_29981,N_18030,N_18286);
nor U29982 (N_29982,N_19104,N_18241);
xor U29983 (N_29983,N_22047,N_18401);
nor U29984 (N_29984,N_22853,N_20448);
and U29985 (N_29985,N_20682,N_23610);
nand U29986 (N_29986,N_19995,N_23286);
or U29987 (N_29987,N_18279,N_20953);
nor U29988 (N_29988,N_23096,N_23444);
or U29989 (N_29989,N_19594,N_23305);
nand U29990 (N_29990,N_23018,N_20169);
and U29991 (N_29991,N_19411,N_20187);
or U29992 (N_29992,N_18767,N_21849);
or U29993 (N_29993,N_18505,N_23067);
nor U29994 (N_29994,N_20134,N_20216);
nor U29995 (N_29995,N_19098,N_23802);
nand U29996 (N_29996,N_18541,N_20116);
xnor U29997 (N_29997,N_23352,N_19211);
nor U29998 (N_29998,N_22378,N_18063);
nor U29999 (N_29999,N_19976,N_21817);
or UO_0 (O_0,N_29760,N_29551);
and UO_1 (O_1,N_25446,N_27227);
or UO_2 (O_2,N_24304,N_25063);
nor UO_3 (O_3,N_26813,N_28600);
xor UO_4 (O_4,N_27692,N_28151);
and UO_5 (O_5,N_27526,N_28014);
and UO_6 (O_6,N_24280,N_27414);
and UO_7 (O_7,N_24481,N_28290);
xor UO_8 (O_8,N_24373,N_26806);
nor UO_9 (O_9,N_26491,N_26354);
and UO_10 (O_10,N_29106,N_28410);
and UO_11 (O_11,N_28509,N_28325);
and UO_12 (O_12,N_25046,N_27049);
and UO_13 (O_13,N_29416,N_25923);
or UO_14 (O_14,N_24581,N_26614);
nand UO_15 (O_15,N_27774,N_27258);
nor UO_16 (O_16,N_29914,N_24763);
nand UO_17 (O_17,N_28741,N_28982);
nand UO_18 (O_18,N_26812,N_29816);
or UO_19 (O_19,N_25317,N_25837);
and UO_20 (O_20,N_26244,N_25381);
nand UO_21 (O_21,N_29011,N_25251);
nand UO_22 (O_22,N_24276,N_29877);
xor UO_23 (O_23,N_25474,N_26419);
nand UO_24 (O_24,N_28739,N_26867);
or UO_25 (O_25,N_27303,N_26370);
or UO_26 (O_26,N_27013,N_26821);
nand UO_27 (O_27,N_24410,N_27617);
or UO_28 (O_28,N_29888,N_26360);
xnor UO_29 (O_29,N_24720,N_26390);
nand UO_30 (O_30,N_26189,N_28830);
nand UO_31 (O_31,N_27741,N_28770);
nor UO_32 (O_32,N_27708,N_29792);
nand UO_33 (O_33,N_24774,N_26226);
nor UO_34 (O_34,N_26619,N_25127);
nor UO_35 (O_35,N_24629,N_25714);
nand UO_36 (O_36,N_24782,N_27084);
nor UO_37 (O_37,N_24744,N_27018);
and UO_38 (O_38,N_29402,N_28404);
nand UO_39 (O_39,N_24022,N_25948);
or UO_40 (O_40,N_27546,N_28440);
and UO_41 (O_41,N_27942,N_24787);
or UO_42 (O_42,N_24094,N_26225);
and UO_43 (O_43,N_26047,N_29084);
and UO_44 (O_44,N_24290,N_27566);
xor UO_45 (O_45,N_27914,N_25229);
nand UO_46 (O_46,N_27534,N_27957);
and UO_47 (O_47,N_28894,N_29170);
nor UO_48 (O_48,N_26259,N_29297);
nand UO_49 (O_49,N_24722,N_27365);
nand UO_50 (O_50,N_29775,N_27464);
nand UO_51 (O_51,N_28213,N_29182);
nor UO_52 (O_52,N_29615,N_27346);
xor UO_53 (O_53,N_27614,N_26532);
nor UO_54 (O_54,N_28783,N_24854);
and UO_55 (O_55,N_26470,N_28993);
nand UO_56 (O_56,N_26086,N_26411);
or UO_57 (O_57,N_24256,N_24267);
and UO_58 (O_58,N_27480,N_25295);
and UO_59 (O_59,N_28375,N_25760);
nand UO_60 (O_60,N_29504,N_29431);
xor UO_61 (O_61,N_26272,N_29249);
nor UO_62 (O_62,N_26495,N_25783);
or UO_63 (O_63,N_24622,N_26228);
nand UO_64 (O_64,N_25458,N_27832);
nand UO_65 (O_65,N_29741,N_26933);
or UO_66 (O_66,N_27153,N_24526);
or UO_67 (O_67,N_24610,N_29190);
or UO_68 (O_68,N_26547,N_27055);
nand UO_69 (O_69,N_27073,N_25161);
and UO_70 (O_70,N_29440,N_24509);
or UO_71 (O_71,N_29569,N_24014);
and UO_72 (O_72,N_25542,N_27670);
and UO_73 (O_73,N_26981,N_27148);
or UO_74 (O_74,N_27651,N_29452);
and UO_75 (O_75,N_26582,N_27511);
or UO_76 (O_76,N_26635,N_25489);
nor UO_77 (O_77,N_27770,N_24514);
nor UO_78 (O_78,N_24490,N_26801);
and UO_79 (O_79,N_26923,N_25374);
nor UO_80 (O_80,N_29386,N_29141);
or UO_81 (O_81,N_24510,N_28769);
xor UO_82 (O_82,N_26171,N_29938);
and UO_83 (O_83,N_25723,N_27856);
nor UO_84 (O_84,N_25033,N_28652);
nor UO_85 (O_85,N_24092,N_26580);
nand UO_86 (O_86,N_27739,N_26456);
or UO_87 (O_87,N_25601,N_29359);
or UO_88 (O_88,N_24487,N_25766);
or UO_89 (O_89,N_28117,N_25029);
or UO_90 (O_90,N_25720,N_27560);
xor UO_91 (O_91,N_26686,N_27290);
nand UO_92 (O_92,N_28210,N_25071);
or UO_93 (O_93,N_24077,N_25176);
nor UO_94 (O_94,N_29063,N_25757);
and UO_95 (O_95,N_29673,N_27982);
xnor UO_96 (O_96,N_29663,N_26040);
nor UO_97 (O_97,N_28198,N_26604);
nand UO_98 (O_98,N_24516,N_25701);
and UO_99 (O_99,N_25526,N_27890);
nor UO_100 (O_100,N_27090,N_24137);
nor UO_101 (O_101,N_24289,N_27568);
nor UO_102 (O_102,N_28633,N_24456);
and UO_103 (O_103,N_25985,N_29468);
or UO_104 (O_104,N_24306,N_27452);
nand UO_105 (O_105,N_28272,N_27396);
nor UO_106 (O_106,N_25461,N_24495);
and UO_107 (O_107,N_26583,N_29171);
xor UO_108 (O_108,N_29574,N_25727);
and UO_109 (O_109,N_29890,N_24529);
nor UO_110 (O_110,N_28716,N_29484);
and UO_111 (O_111,N_28271,N_29969);
or UO_112 (O_112,N_28348,N_25619);
and UO_113 (O_113,N_25730,N_25551);
nor UO_114 (O_114,N_29116,N_27214);
nor UO_115 (O_115,N_28631,N_29318);
and UO_116 (O_116,N_28753,N_27537);
nand UO_117 (O_117,N_26964,N_24450);
nand UO_118 (O_118,N_24590,N_27091);
nand UO_119 (O_119,N_24036,N_29537);
and UO_120 (O_120,N_26528,N_28461);
nand UO_121 (O_121,N_25379,N_25777);
nor UO_122 (O_122,N_24753,N_25280);
xor UO_123 (O_123,N_28368,N_25561);
or UO_124 (O_124,N_26022,N_29566);
nand UO_125 (O_125,N_28657,N_24929);
or UO_126 (O_126,N_24649,N_29616);
nand UO_127 (O_127,N_25967,N_27118);
nor UO_128 (O_128,N_27187,N_26865);
and UO_129 (O_129,N_26416,N_24217);
and UO_130 (O_130,N_25538,N_29902);
nand UO_131 (O_131,N_27151,N_25175);
and UO_132 (O_132,N_29438,N_25368);
and UO_133 (O_133,N_28275,N_27740);
nand UO_134 (O_134,N_26277,N_27017);
nand UO_135 (O_135,N_24931,N_25205);
or UO_136 (O_136,N_27532,N_26036);
nand UO_137 (O_137,N_28081,N_25825);
nor UO_138 (O_138,N_29721,N_27970);
and UO_139 (O_139,N_27494,N_28629);
nand UO_140 (O_140,N_29686,N_26027);
or UO_141 (O_141,N_29373,N_26151);
xnor UO_142 (O_142,N_29062,N_29494);
nand UO_143 (O_143,N_28510,N_25607);
nor UO_144 (O_144,N_25569,N_29202);
or UO_145 (O_145,N_29517,N_25740);
nor UO_146 (O_146,N_29633,N_27001);
nor UO_147 (O_147,N_26765,N_25143);
nor UO_148 (O_148,N_28417,N_25077);
nand UO_149 (O_149,N_25259,N_26957);
nor UO_150 (O_150,N_29611,N_24947);
nor UO_151 (O_151,N_28330,N_26887);
nor UO_152 (O_152,N_29844,N_28845);
nand UO_153 (O_153,N_24012,N_26335);
or UO_154 (O_154,N_24983,N_29681);
nand UO_155 (O_155,N_29174,N_25291);
nor UO_156 (O_156,N_27007,N_29164);
or UO_157 (O_157,N_26164,N_25741);
nand UO_158 (O_158,N_27045,N_27766);
or UO_159 (O_159,N_27887,N_27893);
nand UO_160 (O_160,N_24329,N_27563);
xor UO_161 (O_161,N_28972,N_28393);
or UO_162 (O_162,N_24240,N_26632);
or UO_163 (O_163,N_29530,N_26123);
nand UO_164 (O_164,N_26165,N_29898);
nand UO_165 (O_165,N_27334,N_26915);
xor UO_166 (O_166,N_27570,N_28152);
nor UO_167 (O_167,N_25832,N_27158);
nand UO_168 (O_168,N_27004,N_28082);
and UO_169 (O_169,N_28777,N_24806);
and UO_170 (O_170,N_26548,N_26644);
nand UO_171 (O_171,N_28345,N_28350);
and UO_172 (O_172,N_25342,N_24169);
nor UO_173 (O_173,N_25166,N_29463);
nand UO_174 (O_174,N_24299,N_24684);
and UO_175 (O_175,N_27831,N_25906);
nor UO_176 (O_176,N_28609,N_24551);
and UO_177 (O_177,N_29756,N_24208);
nor UO_178 (O_178,N_27975,N_28215);
and UO_179 (O_179,N_28146,N_28954);
or UO_180 (O_180,N_29052,N_25540);
nor UO_181 (O_181,N_25828,N_27427);
nand UO_182 (O_182,N_25674,N_25678);
and UO_183 (O_183,N_24016,N_28487);
and UO_184 (O_184,N_27724,N_27213);
nand UO_185 (O_185,N_28431,N_27763);
nor UO_186 (O_186,N_29997,N_29753);
and UO_187 (O_187,N_28551,N_28898);
and UO_188 (O_188,N_29090,N_28274);
nand UO_189 (O_189,N_26121,N_28385);
xnor UO_190 (O_190,N_27329,N_29475);
nand UO_191 (O_191,N_27256,N_25450);
and UO_192 (O_192,N_24350,N_28493);
and UO_193 (O_193,N_28425,N_25931);
nand UO_194 (O_194,N_25628,N_26706);
xor UO_195 (O_195,N_25328,N_27752);
nor UO_196 (O_196,N_28495,N_29820);
and UO_197 (O_197,N_27907,N_28423);
and UO_198 (O_198,N_25979,N_28411);
and UO_199 (O_199,N_29549,N_24205);
xor UO_200 (O_200,N_28126,N_28683);
or UO_201 (O_201,N_25774,N_24407);
or UO_202 (O_202,N_24628,N_27133);
and UO_203 (O_203,N_26603,N_27143);
and UO_204 (O_204,N_28344,N_25498);
xnor UO_205 (O_205,N_27330,N_24078);
nor UO_206 (O_206,N_27418,N_27218);
and UO_207 (O_207,N_29958,N_24991);
nand UO_208 (O_208,N_27631,N_28907);
nor UO_209 (O_209,N_24583,N_26024);
nand UO_210 (O_210,N_29007,N_27124);
nor UO_211 (O_211,N_25758,N_27152);
or UO_212 (O_212,N_25057,N_26602);
nor UO_213 (O_213,N_29845,N_25467);
nand UO_214 (O_214,N_26886,N_24275);
xnor UO_215 (O_215,N_27367,N_26820);
or UO_216 (O_216,N_25167,N_25662);
nand UO_217 (O_217,N_29409,N_28719);
nor UO_218 (O_218,N_29300,N_27040);
nor UO_219 (O_219,N_29237,N_24598);
nor UO_220 (O_220,N_27591,N_28457);
or UO_221 (O_221,N_26477,N_26270);
and UO_222 (O_222,N_28178,N_26714);
xnor UO_223 (O_223,N_25594,N_25506);
xor UO_224 (O_224,N_24406,N_27729);
and UO_225 (O_225,N_28278,N_25853);
nor UO_226 (O_226,N_25657,N_26336);
nand UO_227 (O_227,N_29602,N_28458);
or UO_228 (O_228,N_27405,N_28538);
and UO_229 (O_229,N_25611,N_26633);
and UO_230 (O_230,N_28462,N_28966);
and UO_231 (O_231,N_29331,N_28060);
and UO_232 (O_232,N_27082,N_24172);
and UO_233 (O_233,N_25862,N_29443);
nand UO_234 (O_234,N_29789,N_27483);
or UO_235 (O_235,N_24361,N_29570);
nor UO_236 (O_236,N_27521,N_25924);
nor UO_237 (O_237,N_28134,N_26381);
nor UO_238 (O_238,N_27713,N_29461);
and UO_239 (O_239,N_24918,N_27478);
nand UO_240 (O_240,N_29637,N_29307);
or UO_241 (O_241,N_28402,N_29508);
xnor UO_242 (O_242,N_27261,N_27446);
and UO_243 (O_243,N_26041,N_27720);
nand UO_244 (O_244,N_24059,N_25243);
or UO_245 (O_245,N_27941,N_27497);
and UO_246 (O_246,N_24285,N_29632);
nand UO_247 (O_247,N_27829,N_29874);
nor UO_248 (O_248,N_24040,N_25350);
or UO_249 (O_249,N_24080,N_27398);
nor UO_250 (O_250,N_27658,N_24884);
nand UO_251 (O_251,N_27307,N_29675);
and UO_252 (O_252,N_24367,N_27275);
or UO_253 (O_253,N_29030,N_28920);
xnor UO_254 (O_254,N_25391,N_25797);
nor UO_255 (O_255,N_26681,N_28670);
xor UO_256 (O_256,N_27571,N_26288);
and UO_257 (O_257,N_25492,N_25304);
or UO_258 (O_258,N_28756,N_24126);
nor UO_259 (O_259,N_27698,N_28960);
nand UO_260 (O_260,N_24477,N_28908);
and UO_261 (O_261,N_28465,N_25729);
nor UO_262 (O_262,N_27798,N_27431);
or UO_263 (O_263,N_29626,N_26345);
nor UO_264 (O_264,N_28361,N_29762);
or UO_265 (O_265,N_28842,N_28099);
and UO_266 (O_266,N_29897,N_24681);
and UO_267 (O_267,N_26972,N_27401);
and UO_268 (O_268,N_27963,N_27613);
or UO_269 (O_269,N_26304,N_24967);
and UO_270 (O_270,N_26715,N_27604);
nand UO_271 (O_271,N_27687,N_24885);
xor UO_272 (O_272,N_27181,N_25749);
or UO_273 (O_273,N_26422,N_28566);
nand UO_274 (O_274,N_24143,N_27313);
nor UO_275 (O_275,N_25670,N_25691);
xor UO_276 (O_276,N_24969,N_26233);
nand UO_277 (O_277,N_29708,N_26624);
or UO_278 (O_278,N_29638,N_26408);
or UO_279 (O_279,N_29892,N_27689);
or UO_280 (O_280,N_27634,N_24480);
xor UO_281 (O_281,N_26671,N_29781);
nand UO_282 (O_282,N_26800,N_24250);
xnor UO_283 (O_283,N_26198,N_28531);
or UO_284 (O_284,N_25253,N_29613);
xnor UO_285 (O_285,N_28890,N_28723);
nor UO_286 (O_286,N_26462,N_26137);
nand UO_287 (O_287,N_25095,N_28424);
and UO_288 (O_288,N_24537,N_28659);
or UO_289 (O_289,N_29885,N_25930);
or UO_290 (O_290,N_29793,N_25372);
nor UO_291 (O_291,N_25703,N_27823);
nor UO_292 (O_292,N_27594,N_27482);
xor UO_293 (O_293,N_24976,N_26471);
xor UO_294 (O_294,N_29516,N_28292);
or UO_295 (O_295,N_24687,N_28694);
and UO_296 (O_296,N_24951,N_29867);
xor UO_297 (O_297,N_26677,N_24411);
or UO_298 (O_298,N_24536,N_28252);
nand UO_299 (O_299,N_27704,N_28833);
xor UO_300 (O_300,N_28790,N_28264);
or UO_301 (O_301,N_25278,N_27026);
xor UO_302 (O_302,N_26122,N_29479);
nand UO_303 (O_303,N_29072,N_27977);
or UO_304 (O_304,N_24438,N_29244);
nor UO_305 (O_305,N_25738,N_24385);
nor UO_306 (O_306,N_24245,N_24916);
nand UO_307 (O_307,N_27850,N_28864);
or UO_308 (O_308,N_25026,N_26852);
xnor UO_309 (O_309,N_24404,N_25643);
or UO_310 (O_310,N_24990,N_29654);
nand UO_311 (O_311,N_27157,N_26026);
and UO_312 (O_312,N_27293,N_25110);
nor UO_313 (O_313,N_24502,N_24336);
nand UO_314 (O_314,N_27419,N_25710);
or UO_315 (O_315,N_24165,N_28862);
or UO_316 (O_316,N_28572,N_28595);
nor UO_317 (O_317,N_25871,N_28637);
nand UO_318 (O_318,N_26911,N_27519);
and UO_319 (O_319,N_29911,N_27297);
or UO_320 (O_320,N_28500,N_26754);
and UO_321 (O_321,N_26746,N_27363);
nor UO_322 (O_322,N_26163,N_29230);
nor UO_323 (O_323,N_29866,N_26530);
nand UO_324 (O_324,N_29028,N_29413);
nor UO_325 (O_325,N_26088,N_28042);
and UO_326 (O_326,N_29543,N_29374);
or UO_327 (O_327,N_24207,N_25106);
nor UO_328 (O_328,N_29150,N_25994);
and UO_329 (O_329,N_29937,N_28009);
nand UO_330 (O_330,N_25524,N_27128);
and UO_331 (O_331,N_26145,N_29082);
nor UO_332 (O_332,N_28693,N_28162);
and UO_333 (O_333,N_29662,N_29565);
and UO_334 (O_334,N_29357,N_26147);
and UO_335 (O_335,N_25505,N_28205);
and UO_336 (O_336,N_28517,N_24387);
nor UO_337 (O_337,N_24911,N_25991);
nor UO_338 (O_338,N_26083,N_27059);
nand UO_339 (O_339,N_28123,N_25936);
xor UO_340 (O_340,N_27621,N_28055);
nand UO_341 (O_341,N_27439,N_27107);
or UO_342 (O_342,N_29050,N_26312);
and UO_343 (O_343,N_29776,N_26104);
nand UO_344 (O_344,N_24009,N_29159);
nand UO_345 (O_345,N_27701,N_27402);
nand UO_346 (O_346,N_29783,N_24769);
nor UO_347 (O_347,N_29056,N_28771);
nor UO_348 (O_348,N_27973,N_27068);
nor UO_349 (O_349,N_27006,N_28218);
xor UO_350 (O_350,N_29077,N_28552);
nor UO_351 (O_351,N_27197,N_29184);
nor UO_352 (O_352,N_24935,N_24879);
nand UO_353 (O_353,N_28445,N_26777);
or UO_354 (O_354,N_27088,N_28876);
or UO_355 (O_355,N_25215,N_29059);
and UO_356 (O_356,N_28248,N_24142);
or UO_357 (O_357,N_24791,N_24982);
nor UO_358 (O_358,N_26357,N_24847);
nor UO_359 (O_359,N_29629,N_27529);
nand UO_360 (O_360,N_26237,N_28610);
nor UO_361 (O_361,N_28114,N_27686);
or UO_362 (O_362,N_24826,N_26114);
xnor UO_363 (O_363,N_28435,N_24321);
and UO_364 (O_364,N_27474,N_28010);
nor UO_365 (O_365,N_27747,N_28748);
nor UO_366 (O_366,N_28524,N_24718);
nand UO_367 (O_367,N_28561,N_24269);
nor UO_368 (O_368,N_29608,N_24444);
nor UO_369 (O_369,N_28223,N_27678);
nand UO_370 (O_370,N_25355,N_27504);
nand UO_371 (O_371,N_24039,N_27036);
nor UO_372 (O_372,N_28708,N_24534);
nand UO_373 (O_373,N_29136,N_25145);
nand UO_374 (O_374,N_28639,N_25116);
and UO_375 (O_375,N_27841,N_28563);
nor UO_376 (O_376,N_24155,N_28412);
and UO_377 (O_377,N_29278,N_28396);
or UO_378 (O_378,N_27284,N_28291);
nor UO_379 (O_379,N_24591,N_28388);
nor UO_380 (O_380,N_27865,N_28718);
nand UO_381 (O_381,N_28138,N_28983);
nor UO_382 (O_382,N_28220,N_25541);
and UO_383 (O_383,N_27415,N_29218);
or UO_384 (O_384,N_28879,N_27456);
or UO_385 (O_385,N_25584,N_24372);
nor UO_386 (O_386,N_27250,N_25692);
xnor UO_387 (O_387,N_28003,N_24202);
nor UO_388 (O_388,N_24797,N_29540);
nand UO_389 (O_389,N_25773,N_24291);
or UO_390 (O_390,N_25510,N_25273);
nand UO_391 (O_391,N_27345,N_24749);
nor UO_392 (O_392,N_25576,N_25297);
xor UO_393 (O_393,N_28280,N_24596);
or UO_394 (O_394,N_26590,N_28745);
xnor UO_395 (O_395,N_28934,N_29149);
nor UO_396 (O_396,N_25312,N_26728);
nand UO_397 (O_397,N_25868,N_26692);
or UO_398 (O_398,N_26436,N_28505);
nor UO_399 (O_399,N_28488,N_28807);
or UO_400 (O_400,N_28946,N_27775);
nand UO_401 (O_401,N_28587,N_24027);
or UO_402 (O_402,N_27985,N_25512);
nor UO_403 (O_403,N_27586,N_25362);
nor UO_404 (O_404,N_27799,N_27074);
nand UO_405 (O_405,N_28324,N_29575);
and UO_406 (O_406,N_27886,N_24279);
or UO_407 (O_407,N_25423,N_24355);
or UO_408 (O_408,N_26606,N_28621);
or UO_409 (O_409,N_25789,N_24882);
nand UO_410 (O_410,N_29197,N_25174);
nor UO_411 (O_411,N_25990,N_27325);
nand UO_412 (O_412,N_26492,N_25784);
nor UO_413 (O_413,N_28506,N_25976);
nand UO_414 (O_414,N_29073,N_27790);
nand UO_415 (O_415,N_27503,N_26653);
or UO_416 (O_416,N_24630,N_25150);
or UO_417 (O_417,N_29919,N_24613);
and UO_418 (O_418,N_27792,N_28596);
nor UO_419 (O_419,N_27233,N_25098);
xor UO_420 (O_420,N_24535,N_24433);
nand UO_421 (O_421,N_27622,N_29485);
xnor UO_422 (O_422,N_24825,N_25842);
nor UO_423 (O_423,N_24013,N_27241);
nand UO_424 (O_424,N_29970,N_27936);
or UO_425 (O_425,N_28507,N_28101);
nor UO_426 (O_426,N_26660,N_26937);
nor UO_427 (O_427,N_24286,N_24010);
nor UO_428 (O_428,N_24875,N_24021);
xnor UO_429 (O_429,N_28747,N_24159);
nor UO_430 (O_430,N_27911,N_29837);
or UO_431 (O_431,N_29907,N_24726);
and UO_432 (O_432,N_27409,N_27216);
nand UO_433 (O_433,N_24398,N_25866);
nand UO_434 (O_434,N_28405,N_27811);
nor UO_435 (O_435,N_27318,N_27995);
nor UO_436 (O_436,N_25397,N_29419);
nor UO_437 (O_437,N_26386,N_29734);
nand UO_438 (O_438,N_26103,N_27206);
or UO_439 (O_439,N_25831,N_24869);
or UO_440 (O_440,N_28931,N_28937);
nor UO_441 (O_441,N_26181,N_25005);
or UO_442 (O_442,N_27468,N_25290);
nor UO_443 (O_443,N_29018,N_27457);
and UO_444 (O_444,N_24553,N_24166);
and UO_445 (O_445,N_26250,N_28371);
nand UO_446 (O_446,N_28654,N_24562);
nor UO_447 (O_447,N_25241,N_26879);
nand UO_448 (O_448,N_24656,N_25160);
nor UO_449 (O_449,N_29000,N_28688);
and UO_450 (O_450,N_25800,N_28376);
xor UO_451 (O_451,N_29710,N_29643);
and UO_452 (O_452,N_29634,N_27208);
or UO_453 (O_453,N_24272,N_24149);
and UO_454 (O_454,N_27145,N_27654);
xnor UO_455 (O_455,N_27642,N_28407);
or UO_456 (O_456,N_28779,N_25438);
or UO_457 (O_457,N_28449,N_29024);
and UO_458 (O_458,N_28562,N_27885);
nand UO_459 (O_459,N_26142,N_24895);
nand UO_460 (O_460,N_25261,N_25861);
nor UO_461 (O_461,N_27500,N_25457);
nand UO_462 (O_462,N_24531,N_29241);
or UO_463 (O_463,N_26720,N_27210);
and UO_464 (O_464,N_27971,N_27810);
nor UO_465 (O_465,N_26420,N_25435);
or UO_466 (O_466,N_27354,N_24539);
and UO_467 (O_467,N_28037,N_27357);
nand UO_468 (O_468,N_25886,N_27417);
and UO_469 (O_469,N_27039,N_29458);
nor UO_470 (O_470,N_29497,N_25724);
nand UO_471 (O_471,N_29194,N_29521);
nand UO_472 (O_472,N_27510,N_28140);
nor UO_473 (O_473,N_28203,N_28415);
xnor UO_474 (O_474,N_25052,N_29811);
nor UO_475 (O_475,N_28464,N_29689);
and UO_476 (O_476,N_27020,N_29260);
and UO_477 (O_477,N_28814,N_27660);
or UO_478 (O_478,N_27430,N_27242);
and UO_479 (O_479,N_27754,N_26703);
xnor UO_480 (O_480,N_29142,N_27295);
and UO_481 (O_481,N_27437,N_24823);
xnor UO_482 (O_482,N_26516,N_28869);
xor UO_483 (O_483,N_24334,N_24742);
nor UO_484 (O_484,N_28139,N_29875);
or UO_485 (O_485,N_25238,N_26907);
and UO_486 (O_486,N_27322,N_27127);
xor UO_487 (O_487,N_27805,N_28991);
nand UO_488 (O_488,N_28367,N_29916);
nand UO_489 (O_489,N_25378,N_24625);
xor UO_490 (O_490,N_28143,N_29819);
or UO_491 (O_491,N_29074,N_27795);
nand UO_492 (O_492,N_28355,N_25747);
xor UO_493 (O_493,N_25182,N_29381);
nand UO_494 (O_494,N_25283,N_27635);
and UO_495 (O_495,N_27087,N_26804);
and UO_496 (O_496,N_28917,N_24917);
or UO_497 (O_497,N_24631,N_26741);
and UO_498 (O_498,N_24443,N_24429);
nand UO_499 (O_499,N_28172,N_26870);
and UO_500 (O_500,N_24263,N_27783);
nand UO_501 (O_501,N_28840,N_28296);
nor UO_502 (O_502,N_25780,N_25928);
and UO_503 (O_503,N_26751,N_26910);
nor UO_504 (O_504,N_28671,N_24643);
nor UO_505 (O_505,N_27897,N_25860);
or UO_506 (O_506,N_24765,N_29042);
xor UO_507 (O_507,N_24697,N_25237);
nor UO_508 (O_508,N_27582,N_27493);
nand UO_509 (O_509,N_26740,N_28459);
nor UO_510 (O_510,N_28992,N_25211);
nor UO_511 (O_511,N_29262,N_26874);
nand UO_512 (O_512,N_27327,N_27714);
and UO_513 (O_513,N_25660,N_25055);
nor UO_514 (O_514,N_25959,N_24563);
or UO_515 (O_515,N_28408,N_25580);
or UO_516 (O_516,N_26249,N_26756);
xnor UO_517 (O_517,N_25059,N_25549);
nor UO_518 (O_518,N_26192,N_29581);
nand UO_519 (O_519,N_29546,N_28984);
xor UO_520 (O_520,N_25014,N_27667);
nand UO_521 (O_521,N_24352,N_25523);
nor UO_522 (O_522,N_24281,N_25909);
nor UO_523 (O_523,N_27423,N_25228);
nor UO_524 (O_524,N_28384,N_29720);
nand UO_525 (O_525,N_27541,N_26329);
or UO_526 (O_526,N_24366,N_26880);
nor UO_527 (O_527,N_24015,N_26534);
nor UO_528 (O_528,N_28682,N_25840);
nand UO_529 (O_529,N_25798,N_27772);
or UO_530 (O_530,N_29255,N_28791);
and UO_531 (O_531,N_29451,N_24978);
and UO_532 (O_532,N_25889,N_26055);
xnor UO_533 (O_533,N_26747,N_25341);
nand UO_534 (O_534,N_26939,N_27688);
or UO_535 (O_535,N_29325,N_27903);
and UO_536 (O_536,N_27673,N_29707);
or UO_537 (O_537,N_25126,N_28317);
xnor UO_538 (O_538,N_26166,N_29423);
xnor UO_539 (O_539,N_26125,N_26004);
nand UO_540 (O_540,N_27523,N_26019);
xnor UO_541 (O_541,N_25699,N_29617);
nand UO_542 (O_542,N_25180,N_28059);
or UO_543 (O_543,N_27845,N_24396);
nand UO_544 (O_544,N_27425,N_28301);
or UO_545 (O_545,N_28576,N_29940);
nor UO_546 (O_546,N_26628,N_27615);
or UO_547 (O_547,N_26906,N_27544);
nand UO_548 (O_548,N_25882,N_25499);
and UO_549 (O_549,N_26139,N_26905);
and UO_550 (O_550,N_29766,N_28980);
xor UO_551 (O_551,N_28892,N_28822);
nand UO_552 (O_552,N_28363,N_26182);
and UO_553 (O_553,N_26480,N_27837);
nand UO_554 (O_554,N_27411,N_28260);
or UO_555 (O_555,N_27922,N_27876);
and UO_556 (O_556,N_28701,N_27513);
nand UO_557 (O_557,N_27364,N_29147);
nor UO_558 (O_558,N_27436,N_26504);
nor UO_559 (O_559,N_28288,N_28251);
nand UO_560 (O_560,N_25249,N_29157);
and UO_561 (O_561,N_27709,N_24754);
nor UO_562 (O_562,N_28228,N_27574);
xnor UO_563 (O_563,N_27454,N_26639);
and UO_564 (O_564,N_25354,N_24347);
nor UO_565 (O_565,N_25626,N_27685);
or UO_566 (O_566,N_29071,N_29718);
xnor UO_567 (O_567,N_24545,N_28340);
nand UO_568 (O_568,N_29245,N_29651);
nand UO_569 (O_569,N_24528,N_24345);
and UO_570 (O_570,N_28062,N_27530);
or UO_571 (O_571,N_27175,N_27761);
and UO_572 (O_572,N_29833,N_29646);
and UO_573 (O_573,N_29338,N_24136);
and UO_574 (O_574,N_25926,N_28884);
xnor UO_575 (O_575,N_28821,N_27352);
xor UO_576 (O_576,N_25776,N_27818);
nor UO_577 (O_577,N_24793,N_29367);
or UO_578 (O_578,N_25856,N_24233);
or UO_579 (O_579,N_28996,N_25247);
nand UO_580 (O_580,N_27579,N_27916);
or UO_581 (O_581,N_28035,N_28430);
xor UO_582 (O_582,N_27520,N_24652);
xnor UO_583 (O_583,N_25813,N_27035);
nand UO_584 (O_584,N_29918,N_29972);
nor UO_585 (O_585,N_28782,N_29435);
and UO_586 (O_586,N_26843,N_24828);
or UO_587 (O_587,N_24795,N_25987);
and UO_588 (O_588,N_26161,N_29005);
and UO_589 (O_589,N_26824,N_28369);
and UO_590 (O_590,N_28331,N_24700);
and UO_591 (O_591,N_29354,N_26509);
nor UO_592 (O_592,N_28047,N_26097);
nand UO_593 (O_593,N_29559,N_24655);
and UO_594 (O_594,N_29578,N_26982);
and UO_595 (O_595,N_24550,N_26263);
nand UO_596 (O_596,N_28548,N_27255);
or UO_597 (O_597,N_25129,N_24930);
or UO_598 (O_598,N_29183,N_27676);
nand UO_599 (O_599,N_24151,N_25102);
nor UO_600 (O_600,N_27735,N_25490);
or UO_601 (O_601,N_25793,N_29387);
and UO_602 (O_602,N_24944,N_25320);
and UO_603 (O_603,N_24686,N_29850);
or UO_604 (O_604,N_29787,N_24147);
nand UO_605 (O_605,N_25433,N_24454);
nand UO_606 (O_606,N_24780,N_25340);
or UO_607 (O_607,N_29812,N_24678);
or UO_608 (O_608,N_28391,N_24724);
xnor UO_609 (O_609,N_25881,N_26216);
or UO_610 (O_610,N_24871,N_28005);
nand UO_611 (O_611,N_29547,N_24170);
or UO_612 (O_612,N_29983,N_24028);
or UO_613 (O_613,N_28863,N_29723);
nand UO_614 (O_614,N_29027,N_24738);
or UO_615 (O_615,N_24762,N_27159);
nand UO_616 (O_616,N_27778,N_26111);
xor UO_617 (O_617,N_28474,N_24565);
and UO_618 (O_618,N_26434,N_28705);
or UO_619 (O_619,N_27142,N_26115);
and UO_620 (O_620,N_24287,N_27736);
nand UO_621 (O_621,N_29282,N_25203);
nor UO_622 (O_622,N_28043,N_29679);
or UO_623 (O_623,N_24893,N_29296);
or UO_624 (O_624,N_27949,N_27956);
or UO_625 (O_625,N_29098,N_26501);
and UO_626 (O_626,N_24556,N_25517);
or UO_627 (O_627,N_28526,N_26752);
or UO_628 (O_628,N_24402,N_28760);
xor UO_629 (O_629,N_24601,N_25302);
nand UO_630 (O_630,N_26900,N_27680);
nor UO_631 (O_631,N_24062,N_29587);
and UO_632 (O_632,N_28370,N_24032);
and UO_633 (O_633,N_29625,N_29921);
or UO_634 (O_634,N_27177,N_28021);
xor UO_635 (O_635,N_24451,N_24064);
or UO_636 (O_636,N_27116,N_26048);
or UO_637 (O_637,N_26002,N_24986);
and UO_638 (O_638,N_24705,N_26455);
or UO_639 (O_639,N_27077,N_28575);
and UO_640 (O_640,N_29751,N_29589);
and UO_641 (O_641,N_25545,N_26524);
and UO_642 (O_642,N_25184,N_25191);
or UO_643 (O_643,N_29899,N_24530);
and UO_644 (O_644,N_24173,N_26096);
nand UO_645 (O_645,N_29456,N_24734);
and UO_646 (O_646,N_26372,N_29148);
nand UO_647 (O_647,N_27308,N_29065);
and UO_648 (O_648,N_27502,N_29100);
nand UO_649 (O_649,N_29614,N_24418);
nor UO_650 (O_650,N_29731,N_26224);
xor UO_651 (O_651,N_26872,N_26584);
and UO_652 (O_652,N_24437,N_28004);
and UO_653 (O_653,N_28788,N_24856);
nor UO_654 (O_654,N_25912,N_27199);
xnor UO_655 (O_655,N_28520,N_24266);
and UO_656 (O_656,N_26935,N_27536);
nand UO_657 (O_657,N_28832,N_27838);
and UO_658 (O_658,N_25650,N_25637);
or UO_659 (O_659,N_25478,N_26735);
nor UO_660 (O_660,N_24056,N_27803);
nand UO_661 (O_661,N_27601,N_27027);
or UO_662 (O_662,N_28473,N_28429);
nand UO_663 (O_663,N_24431,N_27655);
or UO_664 (O_664,N_26625,N_28560);
nor UO_665 (O_665,N_24727,N_25009);
nor UO_666 (O_666,N_29685,N_25535);
nor UO_667 (O_667,N_27378,N_25493);
nor UO_668 (O_668,N_28028,N_26368);
nor UO_669 (O_669,N_27784,N_26637);
or UO_670 (O_670,N_28534,N_26831);
or UO_671 (O_671,N_29422,N_28818);
and UO_672 (O_672,N_28079,N_24082);
nand UO_673 (O_673,N_27420,N_24511);
and UO_674 (O_674,N_24735,N_24097);
or UO_675 (O_675,N_26341,N_27122);
nand UO_676 (O_676,N_26814,N_27809);
nand UO_677 (O_677,N_27121,N_27375);
nor UO_678 (O_678,N_24206,N_27535);
nand UO_679 (O_679,N_28503,N_25024);
or UO_680 (O_680,N_25164,N_29441);
or UO_681 (O_681,N_24855,N_29519);
or UO_682 (O_682,N_25755,N_26257);
and UO_683 (O_683,N_27244,N_28281);
nor UO_684 (O_684,N_26229,N_26367);
or UO_685 (O_685,N_24393,N_25646);
xor UO_686 (O_686,N_28689,N_27926);
nor UO_687 (O_687,N_28630,N_27451);
nand UO_688 (O_688,N_26724,N_29499);
or UO_689 (O_689,N_24099,N_27254);
and UO_690 (O_690,N_29693,N_24045);
or UO_691 (O_691,N_24838,N_28592);
xnor UO_692 (O_692,N_27930,N_28486);
and UO_693 (O_693,N_24925,N_25330);
nor UO_694 (O_694,N_24308,N_25659);
nand UO_695 (O_695,N_27125,N_24818);
nand UO_696 (O_696,N_29501,N_25622);
nor UO_697 (O_697,N_25880,N_26134);
nor UO_698 (O_698,N_26993,N_26043);
xor UO_699 (O_699,N_26427,N_25468);
xnor UO_700 (O_700,N_28456,N_26621);
and UO_701 (O_701,N_27966,N_27003);
and UO_702 (O_702,N_27131,N_29267);
nor UO_703 (O_703,N_24047,N_29936);
or UO_704 (O_704,N_25661,N_29410);
or UO_705 (O_705,N_27839,N_29904);
nor UO_706 (O_706,N_26319,N_28071);
and UO_707 (O_707,N_28988,N_27705);
and UO_708 (O_708,N_26930,N_28605);
xor UO_709 (O_709,N_24288,N_26718);
nor UO_710 (O_710,N_26818,N_25079);
or UO_711 (O_711,N_29732,N_26207);
and UO_712 (O_712,N_29355,N_25155);
nand UO_713 (O_713,N_25763,N_28646);
or UO_714 (O_714,N_25254,N_29298);
and UO_715 (O_715,N_27076,N_25412);
and UO_716 (O_716,N_26894,N_28116);
nor UO_717 (O_717,N_27304,N_29988);
or UO_718 (O_718,N_26902,N_24111);
or UO_719 (O_719,N_24446,N_26325);
xnor UO_720 (O_720,N_28949,N_27034);
nand UO_721 (O_721,N_26811,N_28279);
nor UO_722 (O_722,N_26442,N_26396);
nand UO_723 (O_723,N_28607,N_25685);
and UO_724 (O_724,N_25230,N_25146);
nand UO_725 (O_725,N_27465,N_26196);
and UO_726 (O_726,N_24690,N_24073);
or UO_727 (O_727,N_27577,N_27955);
or UO_728 (O_728,N_26385,N_25984);
and UO_729 (O_729,N_29603,N_27797);
nand UO_730 (O_730,N_25263,N_27872);
or UO_731 (O_731,N_28641,N_26519);
and UO_732 (O_732,N_25553,N_28968);
and UO_733 (O_733,N_29683,N_25313);
or UO_734 (O_734,N_27165,N_28467);
and UO_735 (O_735,N_24184,N_29697);
or UO_736 (O_736,N_25074,N_29838);
nand UO_737 (O_737,N_25613,N_27170);
nor UO_738 (O_738,N_29544,N_28513);
or UO_739 (O_739,N_26068,N_27215);
nor UO_740 (O_740,N_24403,N_29290);
nand UO_741 (O_741,N_29327,N_24428);
or UO_742 (O_742,N_29449,N_26709);
and UO_743 (O_743,N_29401,N_28843);
or UO_744 (O_744,N_26209,N_28967);
and UO_745 (O_745,N_26438,N_25756);
nor UO_746 (O_746,N_28820,N_28707);
nor UO_747 (O_747,N_24498,N_24558);
nor UO_748 (O_748,N_27992,N_28692);
and UO_749 (O_749,N_29061,N_26545);
and UO_750 (O_750,N_29214,N_26485);
and UO_751 (O_751,N_28033,N_27057);
and UO_752 (O_752,N_29466,N_25196);
nand UO_753 (O_753,N_29601,N_26551);
nor UO_754 (O_754,N_28602,N_29160);
and UO_755 (O_755,N_28297,N_29524);
xor UO_756 (O_756,N_25399,N_26494);
and UO_757 (O_757,N_27948,N_26075);
or UO_758 (O_758,N_27768,N_29865);
or UO_759 (O_759,N_28667,N_26000);
and UO_760 (O_760,N_25639,N_28649);
nand UO_761 (O_761,N_28307,N_24989);
nand UO_762 (O_762,N_27937,N_24277);
and UO_763 (O_763,N_25801,N_29120);
and UO_764 (O_764,N_25431,N_27848);
and UO_765 (O_765,N_28466,N_25904);
nand UO_766 (O_766,N_26726,N_25799);
and UO_767 (O_767,N_26931,N_26987);
and UO_768 (O_768,N_24070,N_26556);
and UO_769 (O_769,N_29019,N_29004);
nand UO_770 (O_770,N_24731,N_28880);
nand UO_771 (O_771,N_29800,N_25501);
and UO_772 (O_772,N_28365,N_28925);
or UO_773 (O_773,N_27416,N_25792);
and UO_774 (O_774,N_25668,N_24654);
and UO_775 (O_775,N_28118,N_25025);
and UO_776 (O_776,N_29406,N_29563);
nand UO_777 (O_777,N_26687,N_27996);
nor UO_778 (O_778,N_24463,N_27952);
nor UO_779 (O_779,N_29848,N_24641);
xnor UO_780 (O_780,N_27287,N_26654);
and UO_781 (O_781,N_27791,N_29102);
nand UO_782 (O_782,N_25497,N_26702);
or UO_783 (O_783,N_29586,N_29991);
and UO_784 (O_784,N_29226,N_27989);
nand UO_785 (O_785,N_29652,N_29870);
nor UO_786 (O_786,N_25193,N_26755);
nor UO_787 (O_787,N_29849,N_26331);
and UO_788 (O_788,N_27368,N_28354);
or UO_789 (O_789,N_26269,N_26180);
or UO_790 (O_790,N_29920,N_26489);
and UO_791 (O_791,N_24075,N_29444);
nand UO_792 (O_792,N_24333,N_29464);
xor UO_793 (O_793,N_27864,N_26693);
nand UO_794 (O_794,N_28874,N_28940);
nor UO_795 (O_795,N_27249,N_25296);
nand UO_796 (O_796,N_29067,N_24824);
or UO_797 (O_797,N_25989,N_26960);
nand UO_798 (O_798,N_26690,N_24846);
or UO_799 (O_799,N_27093,N_27866);
xor UO_800 (O_800,N_29115,N_28665);
or UO_801 (O_801,N_24751,N_26862);
xor UO_802 (O_802,N_27796,N_26618);
or UO_803 (O_803,N_28938,N_26955);
nand UO_804 (O_804,N_29645,N_29259);
nor UO_805 (O_805,N_26559,N_24561);
nand UO_806 (O_806,N_25504,N_29326);
xor UO_807 (O_807,N_25768,N_24185);
or UO_808 (O_808,N_24804,N_27969);
nand UO_809 (O_809,N_24802,N_28030);
nor UO_810 (O_810,N_26733,N_25870);
nor UO_811 (O_811,N_26260,N_29754);
and UO_812 (O_812,N_24758,N_27350);
or UO_813 (O_813,N_28104,N_28776);
and UO_814 (O_814,N_24689,N_29252);
nand UO_815 (O_815,N_29688,N_29852);
nor UO_816 (O_816,N_29799,N_28900);
nand UO_817 (O_817,N_28569,N_28087);
and UO_818 (O_818,N_27361,N_26600);
or UO_819 (O_819,N_29526,N_26734);
or UO_820 (O_820,N_25424,N_28176);
nor UO_821 (O_821,N_25616,N_26555);
or UO_822 (O_822,N_29994,N_24132);
nand UO_823 (O_823,N_25144,N_28761);
nand UO_824 (O_824,N_26346,N_24506);
or UO_825 (O_825,N_25343,N_24167);
and UO_826 (O_826,N_24704,N_28944);
or UO_827 (O_827,N_28684,N_25686);
nor UO_828 (O_828,N_27716,N_29801);
or UO_829 (O_829,N_25068,N_29949);
xnor UO_830 (O_830,N_27373,N_28537);
or UO_831 (O_831,N_25236,N_29332);
nor UO_832 (O_832,N_24907,N_24029);
or UO_833 (O_833,N_27212,N_29627);
nor UO_834 (O_834,N_29717,N_25963);
nand UO_835 (O_835,N_29105,N_24546);
and UO_836 (O_836,N_29719,N_24813);
nor UO_837 (O_837,N_26965,N_29089);
nor UO_838 (O_838,N_24896,N_24771);
and UO_839 (O_839,N_29749,N_25208);
nor UO_840 (O_840,N_26352,N_26661);
xor UO_841 (O_841,N_27557,N_28803);
xnor UO_842 (O_842,N_28026,N_27292);
or UO_843 (O_843,N_24274,N_25265);
nor UO_844 (O_844,N_26415,N_28819);
nor UO_845 (O_845,N_29680,N_27332);
nand UO_846 (O_846,N_24035,N_29043);
or UO_847 (O_847,N_27032,N_24442);
nand UO_848 (O_848,N_29510,N_26376);
and UO_849 (O_849,N_26279,N_27440);
nand UO_850 (O_850,N_28478,N_26028);
xnor UO_851 (O_851,N_26840,N_24434);
or UO_852 (O_852,N_28226,N_28672);
or UO_853 (O_853,N_28808,N_28357);
or UO_854 (O_854,N_26452,N_29698);
nor UO_855 (O_855,N_24887,N_27163);
nor UO_856 (O_856,N_26120,N_24303);
and UO_857 (O_857,N_25746,N_29154);
xor UO_858 (O_858,N_25560,N_24644);
and UO_859 (O_859,N_26766,N_25154);
nand UO_860 (O_860,N_25728,N_24921);
nand UO_861 (O_861,N_26947,N_26146);
and UO_862 (O_862,N_27458,N_28650);
nand UO_863 (O_863,N_27819,N_28627);
nand UO_864 (O_864,N_24400,N_25310);
and UO_865 (O_865,N_26593,N_26406);
and UO_866 (O_866,N_28935,N_27755);
nand UO_867 (O_867,N_27934,N_25010);
and UO_868 (O_868,N_24380,N_26634);
nand UO_869 (O_869,N_26711,N_29054);
or UO_870 (O_870,N_26949,N_28170);
nor UO_871 (O_871,N_25219,N_25765);
nor UO_872 (O_872,N_27382,N_26183);
and UO_873 (O_873,N_25069,N_29655);
or UO_874 (O_874,N_27644,N_28454);
nand UO_875 (O_875,N_29960,N_25969);
and UO_876 (O_876,N_25632,N_24815);
nand UO_877 (O_877,N_27023,N_25531);
or UO_878 (O_878,N_27920,N_29025);
or UO_879 (O_879,N_29500,N_28011);
and UO_880 (O_880,N_26951,N_25970);
nor UO_881 (O_881,N_24088,N_25076);
or UO_882 (O_882,N_29097,N_26184);
xnor UO_883 (O_883,N_25752,N_25496);
and UO_884 (O_884,N_28799,N_25019);
or UO_885 (O_885,N_25597,N_27224);
or UO_886 (O_886,N_26255,N_24360);
or UO_887 (O_887,N_29671,N_25878);
nor UO_888 (O_888,N_26236,N_26557);
and UO_889 (O_889,N_27561,N_25272);
or UO_890 (O_890,N_29424,N_29630);
and UO_891 (O_891,N_25258,N_26529);
nand UO_892 (O_892,N_27815,N_29247);
or UO_893 (O_893,N_25008,N_26869);
nor UO_894 (O_894,N_27648,N_26505);
nor UO_895 (O_895,N_28829,N_27429);
and UO_896 (O_896,N_29631,N_26280);
nor UO_897 (O_897,N_28190,N_28635);
nand UO_898 (O_898,N_25631,N_27612);
xor UO_899 (O_899,N_27098,N_27780);
and UO_900 (O_900,N_26310,N_29933);
nand UO_901 (O_901,N_25748,N_24914);
nand UO_902 (O_902,N_25181,N_28400);
or UO_903 (O_903,N_28795,N_24262);
and UO_904 (O_904,N_26875,N_26179);
nand UO_905 (O_905,N_24532,N_25839);
or UO_906 (O_906,N_28921,N_29281);
nor UO_907 (O_907,N_29814,N_26684);
or UO_908 (O_908,N_29058,N_25092);
or UO_909 (O_909,N_26053,N_28432);
or UO_910 (O_910,N_27869,N_24066);
nor UO_911 (O_911,N_28212,N_24636);
nand UO_912 (O_912,N_27154,N_28801);
xnor UO_913 (O_913,N_29453,N_25084);
and UO_914 (O_914,N_24048,N_25791);
or UO_915 (O_915,N_24264,N_27251);
and UO_916 (O_916,N_27089,N_24603);
and UO_917 (O_917,N_24669,N_27852);
and UO_918 (O_918,N_29477,N_27964);
or UO_919 (O_919,N_24365,N_25679);
and UO_920 (O_920,N_29187,N_27645);
or UO_921 (O_921,N_24378,N_24740);
nand UO_922 (O_922,N_27348,N_25402);
or UO_923 (O_923,N_27598,N_29376);
nand UO_924 (O_924,N_25292,N_26992);
nor UO_925 (O_925,N_25118,N_25833);
and UO_926 (O_926,N_26503,N_27400);
nor UO_927 (O_927,N_24179,N_25598);
nand UO_928 (O_928,N_29378,N_29828);
or UO_929 (O_929,N_27403,N_29140);
or UO_930 (O_930,N_28120,N_29308);
xnor UO_931 (O_931,N_28549,N_28962);
and UO_932 (O_932,N_26753,N_29322);
nand UO_933 (O_933,N_28924,N_28455);
nand UO_934 (O_934,N_26285,N_25786);
nand UO_935 (O_935,N_25572,N_28221);
nor UO_936 (O_936,N_24523,N_27750);
or UO_937 (O_937,N_26135,N_29474);
nand UO_938 (O_938,N_27954,N_29977);
and UO_939 (O_939,N_24777,N_24866);
or UO_940 (O_940,N_29724,N_24948);
or UO_941 (O_941,N_27022,N_28865);
xor UO_942 (O_942,N_28525,N_26531);
nand UO_943 (O_943,N_28374,N_25767);
nand UO_944 (O_944,N_29235,N_29349);
and UO_945 (O_945,N_28269,N_24843);
or UO_946 (O_946,N_29807,N_24125);
and UO_947 (O_947,N_24216,N_26332);
and UO_948 (O_948,N_24131,N_29974);
nand UO_949 (O_949,N_24965,N_27661);
and UO_950 (O_950,N_27610,N_26441);
and UO_951 (O_951,N_24187,N_25992);
nand UO_952 (O_952,N_25218,N_26344);
nor UO_953 (O_953,N_27868,N_29429);
nand UO_954 (O_954,N_25602,N_24790);
nor UO_955 (O_955,N_25835,N_27961);
xnor UO_956 (O_956,N_25621,N_25314);
or UO_957 (O_957,N_26849,N_28824);
nand UO_958 (O_958,N_24394,N_25306);
or UO_959 (O_959,N_24330,N_26805);
and UO_960 (O_960,N_25554,N_27789);
nand UO_961 (O_961,N_25183,N_28480);
or UO_962 (O_962,N_28054,N_28891);
and UO_963 (O_963,N_24096,N_24960);
nand UO_964 (O_964,N_24215,N_28722);
nor UO_965 (O_965,N_28183,N_29730);
or UO_966 (O_966,N_25892,N_28644);
nand UO_967 (O_967,N_26425,N_26031);
and UO_968 (O_968,N_25877,N_27289);
nand UO_969 (O_969,N_29736,N_26340);
nand UO_970 (O_970,N_26328,N_28608);
or UO_971 (O_971,N_29273,N_28337);
or UO_972 (O_972,N_28318,N_25618);
xnor UO_973 (O_973,N_27515,N_24515);
or UO_974 (O_974,N_29292,N_28219);
and UO_975 (O_975,N_25380,N_24421);
or UO_976 (O_976,N_25999,N_24189);
nor UO_977 (O_977,N_24470,N_25591);
or UO_978 (O_978,N_24113,N_26085);
nand UO_979 (O_979,N_28057,N_29996);
or UO_980 (O_980,N_25371,N_27399);
xor UO_981 (O_981,N_27569,N_28620);
nand UO_982 (O_982,N_26908,N_24640);
nor UO_983 (O_983,N_24086,N_24491);
and UO_984 (O_984,N_26167,N_25473);
xnor UO_985 (O_985,N_24091,N_25062);
nor UO_986 (O_986,N_25232,N_27106);
nor UO_987 (O_987,N_24023,N_26116);
and UO_988 (O_988,N_25782,N_26459);
and UO_989 (O_989,N_26057,N_26514);
or UO_990 (O_990,N_25702,N_28591);
or UO_991 (O_991,N_25406,N_27857);
nor UO_992 (O_992,N_28346,N_25287);
nand UO_993 (O_993,N_25859,N_27587);
nand UO_994 (O_994,N_29999,N_25899);
nand UO_995 (O_995,N_29470,N_29993);
and UO_996 (O_996,N_27609,N_28157);
nor UO_997 (O_997,N_25546,N_25135);
or UO_998 (O_998,N_25325,N_29945);
or UO_999 (O_999,N_25893,N_28072);
and UO_1000 (O_1000,N_26566,N_25627);
and UO_1001 (O_1001,N_24063,N_26643);
nor UO_1002 (O_1002,N_26883,N_28153);
xnor UO_1003 (O_1003,N_25539,N_28119);
or UO_1004 (O_1004,N_28625,N_28381);
nand UO_1005 (O_1005,N_25567,N_25642);
nor UO_1006 (O_1006,N_28678,N_24759);
nor UO_1007 (O_1007,N_28848,N_24209);
nor UO_1008 (O_1008,N_25030,N_26994);
and UO_1009 (O_1009,N_24486,N_26066);
or UO_1010 (O_1010,N_25222,N_27979);
or UO_1011 (O_1011,N_28909,N_28556);
or UO_1012 (O_1012,N_24344,N_29196);
nor UO_1013 (O_1013,N_29702,N_25246);
nor UO_1014 (O_1014,N_25884,N_27272);
nand UO_1015 (O_1015,N_27816,N_24371);
nor UO_1016 (O_1016,N_27788,N_24133);
nor UO_1017 (O_1017,N_27573,N_28485);
nor UO_1018 (O_1018,N_24923,N_26571);
nand UO_1019 (O_1019,N_28573,N_26118);
and UO_1020 (O_1020,N_25101,N_24607);
and UO_1021 (O_1021,N_29363,N_28339);
nand UO_1022 (O_1022,N_26796,N_25943);
or UO_1023 (O_1023,N_25413,N_25204);
or UO_1024 (O_1024,N_28077,N_27619);
nand UO_1025 (O_1025,N_27737,N_29761);
and UO_1026 (O_1026,N_28173,N_24157);
or UO_1027 (O_1027,N_27826,N_29505);
or UO_1028 (O_1028,N_26950,N_26678);
and UO_1029 (O_1029,N_28581,N_25038);
nor UO_1030 (O_1030,N_25089,N_27912);
nor UO_1031 (O_1031,N_27883,N_24874);
nor UO_1032 (O_1032,N_29175,N_24322);
nor UO_1033 (O_1033,N_26791,N_26717);
nand UO_1034 (O_1034,N_26848,N_29432);
nand UO_1035 (O_1035,N_24507,N_26963);
nand UO_1036 (O_1036,N_27487,N_25142);
or UO_1037 (O_1037,N_26305,N_27461);
nor UO_1038 (O_1038,N_29156,N_26478);
nand UO_1039 (O_1039,N_26770,N_26889);
or UO_1040 (O_1040,N_29460,N_24750);
nor UO_1041 (O_1041,N_28243,N_24177);
nand UO_1042 (O_1042,N_29927,N_25103);
xnor UO_1043 (O_1043,N_28362,N_27879);
or UO_1044 (O_1044,N_26157,N_24364);
nor UO_1045 (O_1045,N_25898,N_25981);
nand UO_1046 (O_1046,N_28019,N_24693);
and UO_1047 (O_1047,N_29358,N_24316);
or UO_1048 (O_1048,N_29590,N_29478);
and UO_1049 (O_1049,N_26084,N_26102);
nor UO_1050 (O_1050,N_26369,N_27044);
nand UO_1051 (O_1051,N_28977,N_27728);
xor UO_1052 (O_1052,N_24268,N_24183);
nor UO_1053 (O_1053,N_27953,N_29582);
and UO_1054 (O_1054,N_26483,N_27862);
nor UO_1055 (O_1055,N_25398,N_26978);
xor UO_1056 (O_1056,N_25826,N_24295);
nor UO_1057 (O_1057,N_26691,N_26927);
nor UO_1058 (O_1058,N_27744,N_25226);
nand UO_1059 (O_1059,N_27267,N_24633);
and UO_1060 (O_1060,N_26130,N_25907);
nor UO_1061 (O_1061,N_25897,N_24374);
nor UO_1062 (O_1062,N_29572,N_28078);
and UO_1063 (O_1063,N_29795,N_27522);
and UO_1064 (O_1064,N_29271,N_24608);
nor UO_1065 (O_1065,N_27620,N_25787);
and UO_1066 (O_1066,N_29483,N_26803);
xor UO_1067 (O_1067,N_26926,N_29293);
and UO_1068 (O_1068,N_27962,N_24508);
and UO_1069 (O_1069,N_29139,N_27769);
nor UO_1070 (O_1070,N_29434,N_25407);
nor UO_1071 (O_1071,N_24447,N_29369);
nand UO_1072 (O_1072,N_25107,N_26845);
and UO_1073 (O_1073,N_28867,N_26676);
and UO_1074 (O_1074,N_28978,N_28326);
or UO_1075 (O_1075,N_27484,N_24766);
and UO_1076 (O_1076,N_25443,N_24679);
nor UO_1077 (O_1077,N_28232,N_28854);
xor UO_1078 (O_1078,N_25709,N_24176);
and UO_1079 (O_1079,N_25396,N_27700);
xor UO_1080 (O_1080,N_29989,N_28558);
nand UO_1081 (O_1081,N_24822,N_26668);
nand UO_1082 (O_1082,N_28188,N_28923);
xor UO_1083 (O_1083,N_25652,N_29947);
or UO_1084 (O_1084,N_25288,N_28746);
nand UO_1085 (O_1085,N_28726,N_26858);
and UO_1086 (O_1086,N_25522,N_25891);
nand UO_1087 (O_1087,N_28191,N_26178);
nand UO_1088 (O_1088,N_26835,N_26251);
and UO_1089 (O_1089,N_27097,N_28928);
or UO_1090 (O_1090,N_24309,N_24060);
nor UO_1091 (O_1091,N_27311,N_28837);
or UO_1092 (O_1092,N_26383,N_28490);
and UO_1093 (O_1093,N_26670,N_27746);
and UO_1094 (O_1094,N_29138,N_27756);
and UO_1095 (O_1095,N_24741,N_26620);
and UO_1096 (O_1096,N_25806,N_28137);
or UO_1097 (O_1097,N_27820,N_25239);
and UO_1098 (O_1098,N_29403,N_27901);
nor UO_1099 (O_1099,N_29407,N_26318);
nand UO_1100 (O_1100,N_29015,N_25547);
and UO_1101 (O_1101,N_24980,N_27384);
nor UO_1102 (O_1102,N_29324,N_26798);
or UO_1103 (O_1103,N_26888,N_24144);
or UO_1104 (O_1104,N_24538,N_26153);
nand UO_1105 (O_1105,N_28696,N_25937);
nor UO_1106 (O_1106,N_24003,N_24619);
nand UO_1107 (O_1107,N_26464,N_24368);
nand UO_1108 (O_1108,N_25442,N_26458);
and UO_1109 (O_1109,N_29995,N_29316);
xnor UO_1110 (O_1110,N_28319,N_25114);
nor UO_1111 (O_1111,N_25697,N_26890);
or UO_1112 (O_1112,N_27139,N_27663);
nand UO_1113 (O_1113,N_25484,N_25242);
nand UO_1114 (O_1114,N_29053,N_25331);
or UO_1115 (O_1115,N_29436,N_28167);
and UO_1116 (O_1116,N_29782,N_28311);
nor UO_1117 (O_1117,N_29619,N_28952);
or UO_1118 (O_1118,N_26934,N_29674);
nor UO_1119 (O_1119,N_26710,N_28781);
nor UO_1120 (O_1120,N_24701,N_29179);
or UO_1121 (O_1121,N_24124,N_25051);
xnor UO_1122 (O_1122,N_24721,N_24800);
nor UO_1123 (O_1123,N_27608,N_27722);
xnor UO_1124 (O_1124,N_26866,N_24415);
and UO_1125 (O_1125,N_28395,N_29250);
and UO_1126 (O_1126,N_25153,N_25188);
or UO_1127 (O_1127,N_27908,N_24593);
or UO_1128 (O_1128,N_28796,N_24587);
nand UO_1129 (O_1129,N_25574,N_25067);
xor UO_1130 (O_1130,N_27102,N_29057);
nor UO_1131 (O_1131,N_27983,N_29623);
nand UO_1132 (O_1132,N_26289,N_29313);
nand UO_1133 (O_1133,N_29503,N_26107);
nor UO_1134 (O_1134,N_24615,N_28765);
nor UO_1135 (O_1135,N_26234,N_24313);
or UO_1136 (O_1136,N_25293,N_26044);
or UO_1137 (O_1137,N_27219,N_27633);
and UO_1138 (O_1138,N_26262,N_27141);
nand UO_1139 (O_1139,N_26912,N_26645);
nor UO_1140 (O_1140,N_25935,N_29036);
and UO_1141 (O_1141,N_27498,N_26607);
nand UO_1142 (O_1142,N_24945,N_24203);
nor UO_1143 (O_1143,N_26705,N_24821);
and UO_1144 (O_1144,N_26759,N_29498);
xor UO_1145 (O_1145,N_26299,N_27366);
nand UO_1146 (O_1146,N_27277,N_29490);
or UO_1147 (O_1147,N_24861,N_28258);
nand UO_1148 (O_1148,N_29968,N_29329);
nand UO_1149 (O_1149,N_27777,N_24339);
nor UO_1150 (O_1150,N_25346,N_28744);
nand UO_1151 (O_1151,N_28144,N_27426);
and UO_1152 (O_1152,N_24943,N_29869);
and UO_1153 (O_1153,N_27328,N_28080);
or UO_1154 (O_1154,N_28380,N_28446);
nor UO_1155 (O_1155,N_25808,N_29101);
nor UO_1156 (O_1156,N_28614,N_25426);
or UO_1157 (O_1157,N_25735,N_25386);
xnor UO_1158 (O_1158,N_28397,N_25586);
nand UO_1159 (O_1159,N_24671,N_28567);
and UO_1160 (O_1160,N_29333,N_24222);
nor UO_1161 (O_1161,N_24030,N_29690);
nand UO_1162 (O_1162,N_29123,N_26856);
or UO_1163 (O_1163,N_26646,N_25945);
and UO_1164 (O_1164,N_25289,N_28899);
nor UO_1165 (O_1165,N_29206,N_28976);
nor UO_1166 (O_1166,N_25073,N_26961);
and UO_1167 (O_1167,N_29393,N_28073);
nand UO_1168 (O_1168,N_29729,N_28893);
and UO_1169 (O_1169,N_28870,N_28702);
nor UO_1170 (O_1170,N_27386,N_24729);
nor UO_1171 (O_1171,N_24101,N_26424);
or UO_1172 (O_1172,N_24711,N_24932);
nand UO_1173 (O_1173,N_24572,N_24876);
and UO_1174 (O_1174,N_25439,N_24079);
or UO_1175 (O_1175,N_25736,N_27771);
or UO_1176 (O_1176,N_25690,N_24441);
nand UO_1177 (O_1177,N_25704,N_29284);
and UO_1178 (O_1178,N_27800,N_28048);
nand UO_1179 (O_1179,N_25952,N_28245);
nand UO_1180 (O_1180,N_27269,N_27718);
nor UO_1181 (O_1181,N_25123,N_29201);
nor UO_1182 (O_1182,N_28277,N_29108);
or UO_1183 (O_1183,N_25179,N_26286);
or UO_1184 (O_1184,N_28479,N_29114);
or UO_1185 (O_1185,N_24878,N_28554);
nor UO_1186 (O_1186,N_28642,N_28700);
xnor UO_1187 (O_1187,N_24061,N_24436);
nor UO_1188 (O_1188,N_29356,N_25361);
nand UO_1189 (O_1189,N_29467,N_27188);
nand UO_1190 (O_1190,N_28024,N_27909);
and UO_1191 (O_1191,N_29258,N_25344);
nor UO_1192 (O_1192,N_26760,N_26988);
and UO_1193 (O_1193,N_24053,N_26651);
and UO_1194 (O_1194,N_29345,N_29181);
nand UO_1195 (O_1195,N_27234,N_26268);
nor UO_1196 (O_1196,N_24662,N_29901);
xnor UO_1197 (O_1197,N_27730,N_27424);
nor UO_1198 (O_1198,N_29660,N_29351);
and UO_1199 (O_1199,N_28979,N_25390);
or UO_1200 (O_1200,N_29152,N_27176);
and UO_1201 (O_1201,N_26439,N_27564);
nor UO_1202 (O_1202,N_26612,N_24474);
and UO_1203 (O_1203,N_24559,N_25844);
and UO_1204 (O_1204,N_25257,N_25971);
nor UO_1205 (O_1205,N_26786,N_25422);
and UO_1206 (O_1206,N_24747,N_28882);
or UO_1207 (O_1207,N_24231,N_28855);
and UO_1208 (O_1208,N_24829,N_27703);
nand UO_1209 (O_1209,N_27203,N_24959);
or UO_1210 (O_1210,N_27450,N_26141);
nor UO_1211 (O_1211,N_24717,N_26080);
and UO_1212 (O_1212,N_26642,N_28570);
xor UO_1213 (O_1213,N_25120,N_26149);
nor UO_1214 (O_1214,N_24614,N_25887);
or UO_1215 (O_1215,N_29930,N_28112);
nor UO_1216 (O_1216,N_26597,N_25525);
and UO_1217 (O_1217,N_28872,N_25441);
nor UO_1218 (O_1218,N_24164,N_28358);
or UO_1219 (O_1219,N_27524,N_29522);
or UO_1220 (O_1220,N_28989,N_26205);
or UO_1221 (O_1221,N_29925,N_24044);
nor UO_1222 (O_1222,N_29853,N_28904);
xnor UO_1223 (O_1223,N_28847,N_29856);
or UO_1224 (O_1224,N_29527,N_24121);
and UO_1225 (O_1225,N_24152,N_26117);
nand UO_1226 (O_1226,N_25564,N_26893);
xor UO_1227 (O_1227,N_24401,N_27508);
nand UO_1228 (O_1228,N_26986,N_28294);
nand UO_1229 (O_1229,N_29010,N_29854);
nor UO_1230 (O_1230,N_28174,N_27475);
nor UO_1231 (O_1231,N_24100,N_28859);
and UO_1232 (O_1232,N_27453,N_28974);
nor UO_1233 (O_1233,N_27021,N_24540);
and UO_1234 (O_1234,N_29975,N_25130);
and UO_1235 (O_1235,N_27071,N_28398);
and UO_1236 (O_1236,N_28343,N_29254);
nand UO_1237 (O_1237,N_24382,N_26238);
xor UO_1238 (O_1238,N_28161,N_24904);
or UO_1239 (O_1239,N_24695,N_26359);
or UO_1240 (O_1240,N_24542,N_27355);
or UO_1241 (O_1241,N_27144,N_29561);
and UO_1242 (O_1242,N_29980,N_27531);
and UO_1243 (O_1243,N_28023,N_25849);
or UO_1244 (O_1244,N_27824,N_24997);
xnor UO_1245 (O_1245,N_29562,N_24192);
nand UO_1246 (O_1246,N_25305,N_29408);
nand UO_1247 (O_1247,N_26525,N_27050);
and UO_1248 (O_1248,N_28124,N_25315);
nor UO_1249 (O_1249,N_27349,N_29773);
and UO_1250 (O_1250,N_25585,N_26499);
nor UO_1251 (O_1251,N_26578,N_29037);
nand UO_1252 (O_1252,N_27980,N_25248);
xor UO_1253 (O_1253,N_25128,N_24549);
nand UO_1254 (O_1254,N_28749,N_29597);
and UO_1255 (O_1255,N_28130,N_27968);
nor UO_1256 (O_1256,N_26330,N_28135);
nand UO_1257 (O_1257,N_25453,N_25028);
xnor UO_1258 (O_1258,N_24518,N_24888);
or UO_1259 (O_1259,N_29668,N_25841);
and UO_1260 (O_1260,N_26248,N_29203);
and UO_1261 (O_1261,N_25281,N_26361);
or UO_1262 (O_1262,N_25483,N_24479);
nand UO_1263 (O_1263,N_26732,N_26523);
and UO_1264 (O_1264,N_29768,N_28242);
nand UO_1265 (O_1265,N_27434,N_24586);
xor UO_1266 (O_1266,N_26431,N_28100);
nand UO_1267 (O_1267,N_24314,N_25001);
xor UO_1268 (O_1268,N_29714,N_27987);
or UO_1269 (O_1269,N_28685,N_24489);
nor UO_1270 (O_1270,N_25775,N_27408);
nand UO_1271 (O_1271,N_24253,N_27605);
nand UO_1272 (O_1272,N_29389,N_26780);
nor UO_1273 (O_1273,N_24899,N_26769);
nor UO_1274 (O_1274,N_26898,N_25778);
and UO_1275 (O_1275,N_29309,N_25845);
nor UO_1276 (O_1276,N_28168,N_29863);
or UO_1277 (O_1277,N_25929,N_26020);
nand UO_1278 (O_1278,N_24775,N_29842);
nor UO_1279 (O_1279,N_28711,N_24999);
and UO_1280 (O_1280,N_29802,N_28040);
nor UO_1281 (O_1281,N_25901,N_29131);
and UO_1282 (O_1282,N_24328,N_27965);
or UO_1283 (O_1283,N_26402,N_28295);
and UO_1284 (O_1284,N_26037,N_24568);
or UO_1285 (O_1285,N_29492,N_24973);
or UO_1286 (O_1286,N_27785,N_27932);
nand UO_1287 (O_1287,N_27137,N_29847);
and UO_1288 (O_1288,N_28470,N_25138);
xor UO_1289 (O_1289,N_25980,N_29287);
and UO_1290 (O_1290,N_27470,N_25240);
or UO_1291 (O_1291,N_27878,N_28313);
nand UO_1292 (O_1292,N_27479,N_24600);
and UO_1293 (O_1293,N_26672,N_24778);
or UO_1294 (O_1294,N_25725,N_26410);
nand UO_1295 (O_1295,N_26089,N_26010);
nand UO_1296 (O_1296,N_29512,N_25087);
or UO_1297 (O_1297,N_29857,N_28496);
nor UO_1298 (O_1298,N_25448,N_29476);
or UO_1299 (O_1299,N_26347,N_27509);
nand UO_1300 (O_1300,N_27913,N_25099);
xor UO_1301 (O_1301,N_28585,N_26334);
nor UO_1302 (O_1302,N_25227,N_29026);
or UO_1303 (O_1303,N_27173,N_26261);
nor UO_1304 (O_1304,N_24284,N_29133);
and UO_1305 (O_1305,N_26520,N_29711);
nor UO_1306 (O_1306,N_24657,N_27252);
nand UO_1307 (O_1307,N_26126,N_25223);
and UO_1308 (O_1308,N_26897,N_25949);
and UO_1309 (O_1309,N_27274,N_26351);
or UO_1310 (O_1310,N_25172,N_26035);
xnor UO_1311 (O_1311,N_28911,N_26552);
xor UO_1312 (O_1312,N_28312,N_26536);
or UO_1313 (O_1313,N_24840,N_24890);
nor UO_1314 (O_1314,N_25978,N_28482);
and UO_1315 (O_1315,N_29959,N_26533);
nand UO_1316 (O_1316,N_25604,N_24448);
nor UO_1317 (O_1317,N_29017,N_24220);
nor UO_1318 (O_1318,N_24666,N_24533);
or UO_1319 (O_1319,N_27028,N_27441);
nor UO_1320 (O_1320,N_24492,N_28255);
and UO_1321 (O_1321,N_29104,N_24258);
and UO_1322 (O_1322,N_28961,N_24377);
or UO_1323 (O_1323,N_29347,N_27449);
nand UO_1324 (O_1324,N_25475,N_27488);
or UO_1325 (O_1325,N_24419,N_28656);
or UO_1326 (O_1326,N_24604,N_25097);
xnor UO_1327 (O_1327,N_27174,N_27527);
nor UO_1328 (O_1328,N_29088,N_24420);
nand UO_1329 (O_1329,N_29716,N_28053);
and UO_1330 (O_1330,N_26538,N_27518);
nand UO_1331 (O_1331,N_27075,N_27632);
and UO_1332 (O_1332,N_25169,N_26850);
nor UO_1333 (O_1333,N_27745,N_27340);
nand UO_1334 (O_1334,N_24235,N_26997);
or UO_1335 (O_1335,N_29135,N_27553);
nor UO_1336 (O_1336,N_26953,N_25836);
and UO_1337 (O_1337,N_28626,N_24494);
and UO_1338 (O_1338,N_24055,N_26664);
xor UO_1339 (O_1339,N_29111,N_26321);
or UO_1340 (O_1340,N_24193,N_24025);
or UO_1341 (O_1341,N_28437,N_24244);
or UO_1342 (O_1342,N_25508,N_24933);
or UO_1343 (O_1343,N_26658,N_29319);
or UO_1344 (O_1344,N_26487,N_28755);
and UO_1345 (O_1345,N_27472,N_26941);
and UO_1346 (O_1346,N_25610,N_29827);
or UO_1347 (O_1347,N_29554,N_26045);
and UO_1348 (O_1348,N_29585,N_25054);
nand UO_1349 (O_1349,N_29012,N_29533);
and UO_1350 (O_1350,N_25321,N_29618);
nor UO_1351 (O_1351,N_26110,N_24915);
nor UO_1352 (O_1352,N_28655,N_29173);
nor UO_1353 (O_1353,N_27933,N_26968);
and UO_1354 (O_1354,N_28536,N_26191);
and UO_1355 (O_1355,N_26374,N_27851);
xor UO_1356 (O_1356,N_25338,N_25817);
nand UO_1357 (O_1357,N_28158,N_24462);
and UO_1358 (O_1358,N_28481,N_28261);
nor UO_1359 (O_1359,N_29112,N_26223);
and UO_1360 (O_1360,N_26543,N_29794);
xnor UO_1361 (O_1361,N_28521,N_27732);
and UO_1362 (O_1362,N_24210,N_25299);
nand UO_1363 (O_1363,N_29656,N_27679);
xor UO_1364 (O_1364,N_28839,N_24831);
nor UO_1365 (O_1365,N_27094,N_28492);
or UO_1366 (O_1366,N_28186,N_28031);
and UO_1367 (O_1367,N_29709,N_24694);
and UO_1368 (O_1368,N_28956,N_25807);
nand UO_1369 (O_1369,N_27239,N_25220);
nor UO_1370 (O_1370,N_27664,N_24348);
and UO_1371 (O_1371,N_24796,N_24188);
nor UO_1372 (O_1372,N_28329,N_25638);
nand UO_1373 (O_1373,N_24621,N_29006);
or UO_1374 (O_1374,N_29964,N_25595);
and UO_1375 (O_1375,N_29473,N_24471);
nand UO_1376 (O_1376,N_26586,N_27636);
nand UO_1377 (O_1377,N_29188,N_25307);
and UO_1378 (O_1378,N_25011,N_25571);
and UO_1379 (O_1379,N_25664,N_28075);
or UO_1380 (O_1380,N_28617,N_27205);
and UO_1381 (O_1381,N_26173,N_27200);
nand UO_1382 (O_1382,N_28338,N_27606);
nor UO_1383 (O_1383,N_29635,N_24660);
nor UO_1384 (O_1384,N_26046,N_24154);
and UO_1385 (O_1385,N_27247,N_29191);
and UO_1386 (O_1386,N_29846,N_28679);
xor UO_1387 (O_1387,N_24238,N_27389);
nand UO_1388 (O_1388,N_27047,N_28225);
or UO_1389 (O_1389,N_25848,N_27786);
nor UO_1390 (O_1390,N_24389,N_29185);
and UO_1391 (O_1391,N_27525,N_28599);
xor UO_1392 (O_1392,N_24198,N_28612);
xnor UO_1393 (O_1393,N_26235,N_26984);
or UO_1394 (O_1394,N_29404,N_29198);
nor UO_1395 (O_1395,N_29430,N_26323);
or UO_1396 (O_1396,N_25045,N_24026);
nand UO_1397 (O_1397,N_28785,N_24788);
and UO_1398 (O_1398,N_25731,N_26364);
or UO_1399 (O_1399,N_28706,N_28309);
xor UO_1400 (O_1400,N_28555,N_24141);
nor UO_1401 (O_1401,N_28164,N_27759);
or UO_1402 (O_1402,N_24469,N_29815);
and UO_1403 (O_1403,N_27902,N_29311);
nor UO_1404 (O_1404,N_26663,N_24792);
nand UO_1405 (O_1405,N_28266,N_26338);
and UO_1406 (O_1406,N_25528,N_27010);
and UO_1407 (O_1407,N_29390,N_27240);
nor UO_1408 (O_1408,N_27166,N_24234);
xnor UO_1409 (O_1409,N_29288,N_24067);
nor UO_1410 (O_1410,N_28175,N_28058);
and UO_1411 (O_1411,N_24650,N_24212);
and UO_1412 (O_1412,N_28953,N_27855);
nand UO_1413 (O_1413,N_26011,N_29143);
nand UO_1414 (O_1414,N_26952,N_27337);
or UO_1415 (O_1415,N_26970,N_26061);
and UO_1416 (O_1416,N_26453,N_26091);
nand UO_1417 (O_1417,N_27695,N_26573);
nand UO_1418 (O_1418,N_25168,N_24435);
nor UO_1419 (O_1419,N_29310,N_27666);
nor UO_1420 (O_1420,N_24756,N_28827);
nand UO_1421 (O_1421,N_25056,N_24358);
nor UO_1422 (O_1422,N_26003,N_29124);
nand UO_1423 (O_1423,N_26208,N_24970);
or UO_1424 (O_1424,N_25579,N_26472);
nor UO_1425 (O_1425,N_24938,N_24430);
or UO_1426 (O_1426,N_28421,N_27370);
or UO_1427 (O_1427,N_24872,N_26842);
and UO_1428 (O_1428,N_28873,N_26188);
xnor UO_1429 (O_1429,N_25698,N_26544);
nand UO_1430 (O_1430,N_29536,N_28352);
nor UO_1431 (O_1431,N_24521,N_27921);
xor UO_1432 (O_1432,N_25189,N_29205);
xnor UO_1433 (O_1433,N_24706,N_26362);
nor UO_1434 (O_1434,N_27888,N_25916);
and UO_1435 (O_1435,N_25485,N_25908);
nor UO_1436 (O_1436,N_29151,N_29405);
xnor UO_1437 (O_1437,N_26349,N_24342);
or UO_1438 (O_1438,N_29064,N_29525);
xor UO_1439 (O_1439,N_26976,N_27994);
nor UO_1440 (O_1440,N_25869,N_27991);
nor UO_1441 (O_1441,N_29591,N_24648);
nand UO_1442 (O_1442,N_29903,N_27814);
nand UO_1443 (O_1443,N_27031,N_26355);
nand UO_1444 (O_1444,N_24952,N_28142);
or UO_1445 (O_1445,N_25078,N_28841);
and UO_1446 (O_1446,N_25064,N_25482);
xnor UO_1447 (O_1447,N_27998,N_26194);
and UO_1448 (O_1448,N_25666,N_29055);
or UO_1449 (O_1449,N_25946,N_24645);
xnor UO_1450 (O_1450,N_24140,N_27138);
and UO_1451 (O_1451,N_24624,N_24555);
or UO_1452 (O_1452,N_28386,N_26392);
nor UO_1453 (O_1453,N_24071,N_25364);
and UO_1454 (O_1454,N_24730,N_29664);
xor UO_1455 (O_1455,N_25617,N_28254);
nor UO_1456 (O_1456,N_25708,N_29669);
nand UO_1457 (O_1457,N_29976,N_25408);
or UO_1458 (O_1458,N_26159,N_25552);
xor UO_1459 (O_1459,N_29336,N_24034);
xor UO_1460 (O_1460,N_26847,N_26176);
xnor UO_1461 (O_1461,N_24922,N_28308);
xnor UO_1462 (O_1462,N_25577,N_28710);
and UO_1463 (O_1463,N_28107,N_25814);
and UO_1464 (O_1464,N_25932,N_25521);
or UO_1465 (O_1465,N_25334,N_25986);
and UO_1466 (O_1466,N_29137,N_29167);
or UO_1467 (O_1467,N_25185,N_27581);
and UO_1468 (O_1468,N_28532,N_24122);
or UO_1469 (O_1469,N_27331,N_28293);
nand UO_1470 (O_1470,N_26857,N_24934);
nor UO_1471 (O_1471,N_25905,N_25165);
and UO_1472 (O_1472,N_27891,N_29177);
and UO_1473 (O_1473,N_26358,N_24292);
or UO_1474 (O_1474,N_29400,N_25683);
nand UO_1475 (O_1475,N_29091,N_25920);
nand UO_1476 (O_1476,N_29628,N_27565);
nor UO_1477 (O_1477,N_24642,N_25608);
and UO_1478 (O_1478,N_27668,N_26219);
xor UO_1479 (O_1479,N_25600,N_25514);
nor UO_1480 (O_1480,N_25234,N_27584);
or UO_1481 (O_1481,N_24104,N_29087);
nand UO_1482 (O_1482,N_25404,N_27376);
nor UO_1483 (O_1483,N_27029,N_26222);
or UO_1484 (O_1484,N_28074,N_29248);
or UO_1485 (O_1485,N_24570,N_24237);
or UO_1486 (O_1486,N_27195,N_28322);
nor UO_1487 (O_1487,N_29895,N_25058);
nor UO_1488 (O_1488,N_26220,N_27505);
nand UO_1489 (O_1489,N_29385,N_29531);
or UO_1490 (O_1490,N_25718,N_27993);
nand UO_1491 (O_1491,N_29841,N_27650);
and UO_1492 (O_1492,N_27575,N_25915);
and UO_1493 (O_1493,N_28093,N_28129);
nor UO_1494 (O_1494,N_26899,N_25843);
or UO_1495 (O_1495,N_25339,N_29195);
and UO_1496 (O_1496,N_24954,N_25519);
nand UO_1497 (O_1497,N_26301,N_28502);
nand UO_1498 (O_1498,N_26554,N_26510);
nor UO_1499 (O_1499,N_24050,N_26785);
nand UO_1500 (O_1500,N_26570,N_28267);
nand UO_1501 (O_1501,N_25300,N_24354);
and UO_1502 (O_1502,N_26481,N_27665);
nor UO_1503 (O_1503,N_28184,N_29340);
nor UO_1504 (O_1504,N_27939,N_28334);
nor UO_1505 (O_1505,N_27607,N_25104);
nand UO_1506 (O_1506,N_25141,N_25075);
xor UO_1507 (O_1507,N_24211,N_27822);
and UO_1508 (O_1508,N_27134,N_28875);
nor UO_1509 (O_1509,N_24488,N_24632);
nand UO_1510 (O_1510,N_29417,N_26860);
nand UO_1511 (O_1511,N_28499,N_28150);
or UO_1512 (O_1512,N_26892,N_29256);
nand UO_1513 (O_1513,N_28154,N_26895);
nand UO_1514 (O_1514,N_26700,N_28713);
nand UO_1515 (O_1515,N_25609,N_26966);
and UO_1516 (O_1516,N_24908,N_28758);
nor UO_1517 (O_1517,N_27374,N_28310);
nor UO_1518 (O_1518,N_24910,N_27599);
nor UO_1519 (O_1519,N_25277,N_27643);
nor UO_1520 (O_1520,N_29604,N_25375);
or UO_1521 (O_1521,N_26716,N_26928);
and UO_1522 (O_1522,N_25013,N_24466);
nor UO_1523 (O_1523,N_28438,N_29532);
nor UO_1524 (O_1524,N_29395,N_27404);
nand UO_1525 (O_1525,N_25515,N_24500);
nor UO_1526 (O_1526,N_24665,N_26204);
xor UO_1527 (O_1527,N_24008,N_27058);
or UO_1528 (O_1528,N_28106,N_29599);
nor UO_1529 (O_1529,N_26885,N_28964);
and UO_1530 (O_1530,N_29986,N_24852);
nor UO_1531 (O_1531,N_25163,N_28995);
or UO_1532 (O_1532,N_27656,N_25158);
nand UO_1533 (O_1533,N_27600,N_28553);
or UO_1534 (O_1534,N_28888,N_25434);
xnor UO_1535 (O_1535,N_28426,N_28522);
nand UO_1536 (O_1536,N_24331,N_27385);
nor UO_1537 (O_1537,N_29641,N_25085);
nand UO_1538 (O_1538,N_25518,N_24504);
or UO_1539 (O_1539,N_26596,N_27012);
nand UO_1540 (O_1540,N_29973,N_27014);
xnor UO_1541 (O_1541,N_28239,N_27997);
nor UO_1542 (O_1542,N_29824,N_27111);
or UO_1543 (O_1543,N_26124,N_25680);
or UO_1544 (O_1544,N_25960,N_27164);
nor UO_1545 (O_1545,N_26513,N_24041);
or UO_1546 (O_1546,N_24108,N_27333);
nor UO_1547 (O_1547,N_25855,N_27435);
nand UO_1548 (O_1548,N_27288,N_28922);
nand UO_1549 (O_1549,N_25113,N_24709);
nand UO_1550 (O_1550,N_28237,N_25301);
and UO_1551 (O_1551,N_28877,N_24961);
xor UO_1552 (O_1552,N_25454,N_29855);
nor UO_1553 (O_1553,N_26435,N_27981);
and UO_1554 (O_1554,N_28802,N_26138);
xnor UO_1555 (O_1555,N_27136,N_26418);
nand UO_1556 (O_1556,N_29075,N_28039);
or UO_1557 (O_1557,N_24482,N_28105);
xor UO_1558 (O_1558,N_25982,N_25327);
and UO_1559 (O_1559,N_28712,N_24112);
or UO_1560 (O_1560,N_25156,N_28918);
or UO_1561 (O_1561,N_25544,N_26776);
nor UO_1562 (O_1562,N_25387,N_25954);
or UO_1563 (O_1563,N_24781,N_26802);
and UO_1564 (O_1564,N_27825,N_27041);
nand UO_1565 (O_1565,N_28497,N_24809);
nor UO_1566 (O_1566,N_29242,N_29961);
and UO_1567 (O_1567,N_25309,N_25463);
or UO_1568 (O_1568,N_26460,N_24962);
and UO_1569 (O_1569,N_26009,N_29595);
or UO_1570 (O_1570,N_27538,N_28103);
or UO_1571 (O_1571,N_26924,N_28256);
nand UO_1572 (O_1572,N_26221,N_26844);
or UO_1573 (O_1573,N_24255,N_26649);
and UO_1574 (O_1574,N_26736,N_27757);
or UO_1575 (O_1575,N_26211,N_29117);
or UO_1576 (O_1576,N_25534,N_26511);
or UO_1577 (O_1577,N_25815,N_26808);
and UO_1578 (O_1578,N_29513,N_28740);
and UO_1579 (O_1579,N_29621,N_28113);
and UO_1580 (O_1580,N_25491,N_29778);
xnor UO_1581 (O_1581,N_29555,N_25507);
and UO_1582 (O_1582,N_25712,N_26278);
or UO_1583 (O_1583,N_27207,N_25563);
nor UO_1584 (O_1584,N_28209,N_25953);
or UO_1585 (O_1585,N_25065,N_24799);
nor UO_1586 (O_1586,N_26382,N_26326);
or UO_1587 (O_1587,N_27342,N_25357);
and UO_1588 (O_1588,N_24180,N_25605);
nor UO_1589 (O_1589,N_28927,N_25027);
and UO_1590 (O_1590,N_25367,N_25271);
and UO_1591 (O_1591,N_29593,N_28109);
nand UO_1592 (O_1592,N_27360,N_28851);
nor UO_1593 (O_1593,N_28111,N_28632);
nor UO_1594 (O_1594,N_28017,N_27918);
or UO_1595 (O_1595,N_26884,N_24182);
xnor UO_1596 (O_1596,N_28985,N_24807);
xor UO_1597 (O_1597,N_24668,N_26393);
and UO_1598 (O_1598,N_29132,N_28715);
nor UO_1599 (O_1599,N_25040,N_26871);
nor UO_1600 (O_1600,N_26727,N_29836);
nand UO_1601 (O_1601,N_26830,N_27377);
and UO_1602 (O_1602,N_24369,N_25867);
or UO_1603 (O_1603,N_27283,N_28601);
xor UO_1604 (O_1604,N_28813,N_27639);
and UO_1605 (O_1605,N_27265,N_29851);
nand UO_1606 (O_1606,N_29769,N_24319);
or UO_1607 (O_1607,N_24936,N_29328);
nand UO_1608 (O_1608,N_29253,N_29777);
or UO_1609 (O_1609,N_25311,N_26377);
nor UO_1610 (O_1610,N_28283,N_27019);
xnor UO_1611 (O_1611,N_28342,N_27444);
or UO_1612 (O_1612,N_28955,N_28673);
nand UO_1613 (O_1613,N_27974,N_29556);
nor UO_1614 (O_1614,N_26508,N_27410);
nand UO_1615 (O_1615,N_27884,N_28622);
nor UO_1616 (O_1616,N_29998,N_26767);
nor UO_1617 (O_1617,N_25148,N_25088);
nor UO_1618 (O_1618,N_29909,N_24712);
and UO_1619 (O_1619,N_25788,N_26868);
and UO_1620 (O_1620,N_28051,N_29805);
nor UO_1621 (O_1621,N_24626,N_28002);
nand UO_1622 (O_1622,N_28618,N_25694);
nand UO_1623 (O_1623,N_25159,N_26876);
nand UO_1624 (O_1624,N_29511,N_27543);
nand UO_1625 (O_1625,N_24957,N_24842);
or UO_1626 (O_1626,N_26913,N_25322);
or UO_1627 (O_1627,N_29040,N_26675);
or UO_1628 (O_1628,N_28825,N_25091);
nand UO_1629 (O_1629,N_26921,N_26779);
or UO_1630 (O_1630,N_28441,N_24218);
nor UO_1631 (O_1631,N_24699,N_28528);
nand UO_1632 (O_1632,N_29362,N_25214);
xnor UO_1633 (O_1633,N_26750,N_29277);
and UO_1634 (O_1634,N_27764,N_26863);
nand UO_1635 (O_1635,N_29060,N_26465);
or UO_1636 (O_1636,N_24000,N_28565);
and UO_1637 (O_1637,N_25037,N_29128);
nand UO_1638 (O_1638,N_25734,N_28403);
nand UO_1639 (O_1639,N_29955,N_29509);
and UO_1640 (O_1640,N_25432,N_25875);
nand UO_1641 (O_1641,N_29304,N_29118);
nor UO_1642 (O_1642,N_27638,N_28686);
and UO_1643 (O_1643,N_25653,N_28450);
nand UO_1644 (O_1644,N_28638,N_24623);
and UO_1645 (O_1645,N_25122,N_24340);
nor UO_1646 (O_1646,N_26995,N_28378);
and UO_1647 (O_1647,N_28419,N_25516);
nand UO_1648 (O_1648,N_26293,N_24658);
nor UO_1649 (O_1649,N_25436,N_29981);
nand UO_1650 (O_1650,N_28943,N_28038);
nor UO_1651 (O_1651,N_25565,N_28483);
nor UO_1652 (O_1652,N_29785,N_28356);
or UO_1653 (O_1653,N_24580,N_25279);
xnor UO_1654 (O_1654,N_29653,N_24478);
nand UO_1655 (O_1655,N_24178,N_29963);
or UO_1656 (O_1656,N_28453,N_29238);
nand UO_1657 (O_1657,N_26498,N_26265);
nand UO_1658 (O_1658,N_27126,N_26609);
or UO_1659 (O_1659,N_28751,N_28155);
nor UO_1660 (O_1660,N_25353,N_28268);
nand UO_1661 (O_1661,N_29790,N_29079);
nor UO_1662 (O_1662,N_27467,N_27103);
or UO_1663 (O_1663,N_26659,N_29687);
nor UO_1664 (O_1664,N_29219,N_24670);
and UO_1665 (O_1665,N_29840,N_26445);
nand UO_1666 (O_1666,N_24278,N_28885);
nor UO_1667 (O_1667,N_25401,N_29950);
nor UO_1668 (O_1668,N_26034,N_29233);
xnor UO_1669 (O_1669,N_28606,N_29829);
nor UO_1670 (O_1670,N_24249,N_26630);
nand UO_1671 (O_1671,N_29883,N_27310);
nor UO_1672 (O_1672,N_25658,N_25636);
nand UO_1673 (O_1673,N_29303,N_28550);
xor UO_1674 (O_1674,N_29830,N_28947);
nand UO_1675 (O_1675,N_25556,N_29648);
or UO_1676 (O_1676,N_27990,N_26281);
or UO_1677 (O_1677,N_25136,N_27549);
or UO_1678 (O_1678,N_29394,N_29571);
or UO_1679 (O_1679,N_25112,N_24850);
or UO_1680 (O_1680,N_29003,N_25500);
nand UO_1681 (O_1681,N_25589,N_26996);
and UO_1682 (O_1682,N_25444,N_24453);
or UO_1683 (O_1683,N_28303,N_24228);
nand UO_1684 (O_1684,N_26579,N_26615);
or UO_1685 (O_1685,N_25962,N_27830);
or UO_1686 (O_1686,N_25911,N_27115);
or UO_1687 (O_1687,N_25590,N_24602);
or UO_1688 (O_1688,N_27341,N_25416);
nor UO_1689 (O_1689,N_27495,N_25269);
nor UO_1690 (O_1690,N_26017,N_29125);
nor UO_1691 (O_1691,N_26429,N_26148);
and UO_1692 (O_1692,N_26712,N_29144);
or UO_1693 (O_1693,N_26404,N_29935);
or UO_1694 (O_1694,N_24001,N_24186);
nand UO_1695 (O_1695,N_27555,N_24107);
or UO_1696 (O_1696,N_24803,N_25751);
or UO_1697 (O_1697,N_27924,N_24145);
nand UO_1698 (O_1698,N_27945,N_27262);
nor UO_1699 (O_1699,N_28416,N_24270);
or UO_1700 (O_1700,N_29552,N_26227);
nor UO_1701 (O_1701,N_28418,N_25693);
nand UO_1702 (O_1702,N_25732,N_25093);
nor UO_1703 (O_1703,N_24892,N_24472);
nor UO_1704 (O_1704,N_29725,N_28328);
nor UO_1705 (O_1705,N_24175,N_25366);
xor UO_1706 (O_1706,N_28392,N_24351);
and UO_1707 (O_1707,N_29520,N_24163);
nand UO_1708 (O_1708,N_24862,N_29414);
nor UO_1709 (O_1709,N_24293,N_29168);
and UO_1710 (O_1710,N_25365,N_24832);
or UO_1711 (O_1711,N_26838,N_28469);
xor UO_1712 (O_1712,N_24757,N_29747);
and UO_1713 (O_1713,N_29798,N_27711);
or UO_1714 (O_1714,N_27641,N_25647);
nand UO_1715 (O_1715,N_25629,N_26698);
and UO_1716 (O_1716,N_25829,N_26025);
or UO_1717 (O_1717,N_27767,N_29305);
or UO_1718 (O_1718,N_24522,N_29825);
nor UO_1719 (O_1719,N_27940,N_24301);
nor UO_1720 (O_1720,N_27392,N_27171);
and UO_1721 (O_1721,N_27066,N_29457);
nor UO_1722 (O_1722,N_29350,N_24977);
nand UO_1723 (O_1723,N_24748,N_24994);
nand UO_1724 (O_1724,N_27691,N_24716);
and UO_1725 (O_1725,N_29535,N_29227);
nor UO_1726 (O_1726,N_28768,N_26467);
xnor UO_1727 (O_1727,N_29606,N_29272);
and UO_1728 (O_1728,N_29487,N_26030);
and UO_1729 (O_1729,N_24808,N_26792);
nor UO_1730 (O_1730,N_25879,N_29486);
nor UO_1731 (O_1731,N_26039,N_28588);
and UO_1732 (O_1732,N_27353,N_27222);
nor UO_1733 (O_1733,N_28809,N_28881);
nand UO_1734 (O_1734,N_29039,N_29165);
nor UO_1735 (O_1735,N_24860,N_28941);
and UO_1736 (O_1736,N_29178,N_24617);
nand UO_1737 (O_1737,N_29642,N_24953);
nor UO_1738 (O_1738,N_24296,N_29217);
and UO_1739 (O_1739,N_27951,N_27383);
xor UO_1740 (O_1740,N_26423,N_25958);
nor UO_1741 (O_1741,N_27455,N_24006);
nand UO_1742 (O_1742,N_29312,N_26731);
nor UO_1743 (O_1743,N_28778,N_24226);
nor UO_1744 (O_1744,N_24664,N_25082);
nor UO_1745 (O_1745,N_25804,N_28511);
or UO_1746 (O_1746,N_29335,N_26773);
nor UO_1747 (O_1747,N_25385,N_27381);
nand UO_1748 (O_1748,N_28128,N_26144);
nor UO_1749 (O_1749,N_25988,N_28422);
and UO_1750 (O_1750,N_27005,N_27616);
xor UO_1751 (O_1751,N_28196,N_24639);
or UO_1752 (O_1752,N_24674,N_24343);
nand UO_1753 (O_1753,N_26989,N_27640);
and UO_1754 (O_1754,N_24682,N_28583);
nand UO_1755 (O_1755,N_26108,N_28156);
nor UO_1756 (O_1756,N_24051,N_27109);
nor UO_1757 (O_1757,N_24698,N_28805);
nor UO_1758 (O_1758,N_25996,N_28333);
nor UO_1759 (O_1759,N_28729,N_27875);
nand UO_1760 (O_1760,N_26679,N_25888);
xor UO_1761 (O_1761,N_25190,N_26093);
nand UO_1762 (O_1762,N_24956,N_26721);
nor UO_1763 (O_1763,N_25857,N_29022);
xor UO_1764 (O_1764,N_25252,N_26685);
and UO_1765 (O_1765,N_26680,N_27085);
or UO_1766 (O_1766,N_26823,N_25624);
nor UO_1767 (O_1767,N_24294,N_26861);
or UO_1768 (O_1768,N_27929,N_28774);
nand UO_1769 (O_1769,N_28543,N_25850);
nand UO_1770 (O_1770,N_27733,N_29366);
nand UO_1771 (O_1771,N_25221,N_24496);
nand UO_1772 (O_1772,N_27202,N_27552);
xor UO_1773 (O_1773,N_27950,N_28052);
or UO_1774 (O_1774,N_29861,N_26610);
and UO_1775 (O_1775,N_26611,N_28076);
nand UO_1776 (O_1776,N_28016,N_27276);
and UO_1777 (O_1777,N_27273,N_29045);
nand UO_1778 (O_1778,N_29694,N_28564);
or UO_1779 (O_1779,N_29647,N_28068);
or UO_1780 (O_1780,N_26245,N_25745);
nor UO_1781 (O_1781,N_27813,N_25447);
or UO_1782 (O_1782,N_24541,N_24683);
and UO_1783 (O_1783,N_25480,N_27236);
and UO_1784 (O_1784,N_27237,N_29392);
nor UO_1785 (O_1785,N_26232,N_24786);
or UO_1786 (O_1786,N_25117,N_24224);
nand UO_1787 (O_1787,N_29942,N_25041);
and UO_1788 (O_1788,N_24002,N_27870);
nand UO_1789 (O_1789,N_27706,N_26296);
nor UO_1790 (O_1790,N_29713,N_27314);
nand UO_1791 (O_1791,N_29910,N_28594);
and UO_1792 (O_1792,N_26247,N_27081);
and UO_1793 (O_1793,N_26819,N_25061);
nor UO_1794 (O_1794,N_29705,N_27445);
xor UO_1795 (O_1795,N_29371,N_24031);
or UO_1796 (O_1796,N_26168,N_26241);
nand UO_1797 (O_1797,N_26468,N_26591);
nand UO_1798 (O_1798,N_28828,N_27282);
and UO_1799 (O_1799,N_26737,N_25559);
nand UO_1800 (O_1800,N_25048,N_25675);
nand UO_1801 (O_1801,N_25794,N_25477);
or UO_1802 (O_1802,N_26457,N_27853);
nor UO_1803 (O_1803,N_27742,N_29127);
or UO_1804 (O_1804,N_24547,N_27836);
or UO_1805 (O_1805,N_28148,N_24527);
and UO_1806 (O_1806,N_27743,N_24467);
nand UO_1807 (O_1807,N_24440,N_27182);
nor UO_1808 (O_1808,N_27873,N_24905);
nor UO_1809 (O_1809,N_28582,N_25503);
nand UO_1810 (O_1810,N_26585,N_27466);
nor UO_1811 (O_1811,N_25418,N_27300);
nor UO_1812 (O_1812,N_24552,N_27749);
and UO_1813 (O_1813,N_27180,N_26787);
and UO_1814 (O_1814,N_27597,N_27356);
nand UO_1815 (O_1815,N_29797,N_24119);
or UO_1816 (O_1816,N_24046,N_24005);
nor UO_1817 (O_1817,N_24924,N_29155);
nor UO_1818 (O_1818,N_28628,N_29126);
and UO_1819 (O_1819,N_25805,N_24297);
nand UO_1820 (O_1820,N_27753,N_25596);
nand UO_1821 (O_1821,N_28936,N_29739);
xnor UO_1822 (O_1822,N_27037,N_26160);
or UO_1823 (O_1823,N_27156,N_26512);
and UO_1824 (O_1824,N_28149,N_28094);
and UO_1825 (O_1825,N_26050,N_26757);
nand UO_1826 (O_1826,N_26440,N_25902);
nand UO_1827 (O_1827,N_26598,N_24505);
xnor UO_1828 (O_1828,N_26991,N_28732);
nand UO_1829 (O_1829,N_29649,N_25606);
and UO_1830 (O_1830,N_27072,N_27306);
nand UO_1831 (O_1831,N_25032,N_29507);
nor UO_1832 (O_1832,N_26032,N_28020);
and UO_1833 (O_1833,N_24937,N_25481);
nor UO_1834 (O_1834,N_29992,N_27721);
nand UO_1835 (O_1835,N_24219,N_28122);
or UO_1836 (O_1836,N_24767,N_26187);
nand UO_1837 (O_1837,N_26764,N_29929);
and UO_1838 (O_1838,N_26696,N_26729);
or UO_1839 (O_1839,N_28676,N_24635);
nor UO_1840 (O_1840,N_26738,N_26565);
or UO_1841 (O_1841,N_28414,N_24337);
or UO_1842 (O_1842,N_26657,N_25360);
nand UO_1843 (O_1843,N_29372,N_26444);
nor UO_1844 (O_1844,N_29692,N_24543);
nor UO_1845 (O_1845,N_26074,N_26854);
or UO_1846 (O_1846,N_28579,N_29579);
nand UO_1847 (O_1847,N_25268,N_26212);
and UO_1848 (O_1848,N_27662,N_27393);
nand UO_1849 (O_1849,N_28315,N_27551);
or UO_1850 (O_1850,N_27162,N_25873);
nand UO_1851 (O_1851,N_29482,N_26292);
or UO_1852 (O_1852,N_25044,N_29068);
nor UO_1853 (O_1853,N_25885,N_27477);
nand UO_1854 (O_1854,N_24381,N_26315);
or UO_1855 (O_1855,N_29270,N_29377);
and UO_1856 (O_1856,N_25821,N_26079);
and UO_1857 (O_1857,N_29580,N_24229);
and UO_1858 (O_1858,N_27682,N_28448);
nor UO_1859 (O_1859,N_28728,N_27776);
nand UO_1860 (O_1860,N_27590,N_29691);
nand UO_1861 (O_1861,N_29696,N_27183);
nor UO_1862 (O_1862,N_24903,N_28235);
nor UO_1863 (O_1863,N_28651,N_26694);
nand UO_1864 (O_1864,N_25667,N_24900);
or UO_1865 (O_1865,N_24708,N_27067);
nor UO_1866 (O_1866,N_26891,N_24359);
nand UO_1867 (O_1867,N_27580,N_28508);
nand UO_1868 (O_1868,N_29134,N_24102);
and UO_1869 (O_1869,N_28817,N_26076);
nor UO_1870 (O_1870,N_28069,N_25352);
nand UO_1871 (O_1871,N_26665,N_28523);
or UO_1872 (O_1872,N_27960,N_24848);
and UO_1873 (O_1873,N_26563,N_24038);
or UO_1874 (O_1874,N_25020,N_29542);
and UO_1875 (O_1875,N_28443,N_26042);
or UO_1876 (O_1876,N_24920,N_24265);
nor UO_1877 (O_1877,N_25109,N_24578);
xor UO_1878 (O_1878,N_24426,N_24736);
nand UO_1879 (O_1879,N_24975,N_25739);
or UO_1880 (O_1880,N_25303,N_29415);
nand UO_1881 (O_1881,N_29953,N_26303);
and UO_1882 (O_1882,N_28975,N_24940);
or UO_1883 (O_1883,N_24408,N_27802);
or UO_1884 (O_1884,N_24849,N_24835);
or UO_1885 (O_1885,N_28793,N_29266);
or UO_1886 (O_1886,N_27105,N_24409);
nand UO_1887 (O_1887,N_24672,N_26008);
nand UO_1888 (O_1888,N_26081,N_26697);
nand UO_1889 (O_1889,N_28179,N_24376);
nor UO_1890 (O_1890,N_28766,N_27683);
xor UO_1891 (O_1891,N_27827,N_24311);
nand UO_1892 (O_1892,N_24326,N_29418);
nand UO_1893 (O_1893,N_25810,N_25178);
and UO_1894 (O_1894,N_26599,N_27150);
and UO_1895 (O_1895,N_26807,N_29099);
and UO_1896 (O_1896,N_29086,N_24190);
nor UO_1897 (O_1897,N_29186,N_25972);
nor UO_1898 (O_1898,N_27030,N_27562);
and UO_1899 (O_1899,N_28662,N_26095);
nor UO_1900 (O_1900,N_27046,N_27086);
and UO_1901 (O_1901,N_26550,N_28349);
xor UO_1902 (O_1902,N_28738,N_27507);
nand UO_1903 (O_1903,N_27078,N_25023);
nor UO_1904 (O_1904,N_24913,N_24955);
and UO_1905 (O_1905,N_27009,N_25060);
and UO_1906 (O_1906,N_26400,N_27583);
or UO_1907 (O_1907,N_27702,N_24427);
xnor UO_1908 (O_1908,N_25140,N_29523);
and UO_1909 (O_1909,N_26105,N_29821);
or UO_1910 (O_1910,N_25086,N_28262);
nor UO_1911 (O_1911,N_26380,N_25645);
nand UO_1912 (O_1912,N_26650,N_28912);
nand UO_1913 (O_1913,N_24575,N_27280);
and UO_1914 (O_1914,N_29199,N_25570);
nor UO_1915 (O_1915,N_27988,N_27715);
and UO_1916 (O_1916,N_28083,N_28095);
and UO_1917 (O_1917,N_24723,N_27025);
nand UO_1918 (O_1918,N_26517,N_28494);
nor UO_1919 (O_1919,N_26388,N_24349);
xor UO_1920 (O_1920,N_26540,N_25934);
or UO_1921 (O_1921,N_29640,N_27860);
or UO_1922 (O_1922,N_28568,N_29979);
and UO_1923 (O_1923,N_28372,N_27369);
nand UO_1924 (O_1924,N_27849,N_29954);
nand UO_1925 (O_1925,N_24197,N_25460);
and UO_1926 (O_1926,N_26072,N_29491);
and UO_1927 (O_1927,N_26172,N_26652);
or UO_1928 (O_1928,N_27279,N_29450);
and UO_1929 (O_1929,N_29014,N_27184);
nand UO_1930 (O_1930,N_27731,N_27978);
nor UO_1931 (O_1931,N_29858,N_28838);
or UO_1932 (O_1932,N_26549,N_27925);
nor UO_1933 (O_1933,N_28049,N_24606);
nand UO_1934 (O_1934,N_27944,N_24357);
and UO_1935 (O_1935,N_25042,N_27448);
xnor UO_1936 (O_1936,N_28849,N_25137);
nand UO_1937 (O_1937,N_27629,N_29433);
xor UO_1938 (O_1938,N_27840,N_28653);
nor UO_1939 (O_1939,N_26589,N_25332);
nand UO_1940 (O_1940,N_25706,N_29596);
nor UO_1941 (O_1941,N_28025,N_27486);
xor UO_1942 (O_1942,N_25895,N_28535);
nand UO_1943 (O_1943,N_29094,N_24588);
or UO_1944 (O_1944,N_28085,N_25383);
or UO_1945 (O_1945,N_26560,N_24573);
nor UO_1946 (O_1946,N_26938,N_24120);
nor UO_1947 (O_1947,N_24085,N_26940);
xnor UO_1948 (O_1948,N_26140,N_25640);
nor UO_1949 (O_1949,N_24156,N_28533);
or UO_1950 (O_1950,N_28289,N_26302);
nand UO_1951 (O_1951,N_26391,N_28950);
nand UO_1952 (O_1952,N_24020,N_24049);
nor UO_1953 (O_1953,N_28577,N_25411);
or UO_1954 (O_1954,N_26925,N_28858);
and UO_1955 (O_1955,N_29764,N_25919);
xnor UO_1956 (O_1956,N_27051,N_24733);
nand UO_1957 (O_1957,N_29121,N_24995);
nand UO_1958 (O_1958,N_25750,N_28108);
xor UO_1959 (O_1959,N_26294,N_25941);
nor UO_1960 (O_1960,N_28913,N_26291);
nand UO_1961 (O_1961,N_24725,N_25864);
nand UO_1962 (O_1962,N_25419,N_29667);
nor UO_1963 (O_1963,N_24065,N_25707);
and UO_1964 (O_1964,N_28468,N_24127);
nand UO_1965 (O_1965,N_27130,N_27305);
and UO_1966 (O_1966,N_26240,N_25575);
nand UO_1967 (O_1967,N_26778,N_28208);
and UO_1968 (O_1968,N_24320,N_29439);
nand UO_1969 (O_1969,N_24353,N_27438);
nand UO_1970 (O_1970,N_27707,N_27407);
nand UO_1971 (O_1971,N_29695,N_25363);
nand UO_1972 (O_1972,N_26021,N_26366);
nor UO_1973 (O_1973,N_25285,N_27821);
nand UO_1974 (O_1974,N_26131,N_25715);
and UO_1975 (O_1975,N_24567,N_28044);
or UO_1976 (O_1976,N_29346,N_29454);
and UO_1977 (O_1977,N_24637,N_26060);
nor UO_1978 (O_1978,N_27723,N_29737);
nor UO_1979 (O_1979,N_24423,N_29445);
nor UO_1980 (O_1980,N_24405,N_24386);
or UO_1981 (O_1981,N_27052,N_24902);
and UO_1982 (O_1982,N_28231,N_26082);
nor UO_1983 (O_1983,N_24128,N_25726);
and UO_1984 (O_1984,N_27877,N_29289);
and UO_1985 (O_1985,N_26394,N_25213);
nand UO_1986 (O_1986,N_28823,N_27828);
or UO_1987 (O_1987,N_27033,N_28091);
xor UO_1988 (O_1988,N_26699,N_28382);
or UO_1989 (O_1989,N_25235,N_29539);
nand UO_1990 (O_1990,N_27625,N_27725);
nand UO_1991 (O_1991,N_26851,N_24392);
nor UO_1992 (O_1992,N_26809,N_29661);
nor UO_1993 (O_1993,N_28615,N_27413);
nand UO_1994 (O_1994,N_27324,N_26414);
nand UO_1995 (O_1995,N_29261,N_24195);
and UO_1996 (O_1996,N_27185,N_28754);
nor UO_1997 (O_1997,N_24199,N_26999);
nand UO_1998 (O_1998,N_25039,N_24271);
nor UO_1999 (O_1999,N_24576,N_29588);
nand UO_2000 (O_2000,N_27782,N_24667);
nor UO_2001 (O_2001,N_29163,N_28265);
and UO_2002 (O_2002,N_25803,N_24798);
and UO_2003 (O_2003,N_27492,N_24677);
or UO_2004 (O_2004,N_25004,N_24889);
nand UO_2005 (O_2005,N_27080,N_26451);
or UO_2006 (O_2006,N_28504,N_28022);
nor UO_2007 (O_2007,N_27652,N_24685);
or UO_2008 (O_2008,N_25066,N_25527);
or UO_2009 (O_2009,N_25818,N_25834);
nor UO_2010 (O_2010,N_29035,N_28165);
nand UO_2011 (O_2011,N_27999,N_29020);
nand UO_2012 (O_2012,N_28514,N_27002);
nand UO_2013 (O_2013,N_27043,N_25581);
and UO_2014 (O_2014,N_27694,N_27123);
or UO_2015 (O_2015,N_29502,N_25743);
nor UO_2016 (O_2016,N_26588,N_29383);
nor UO_2017 (O_2017,N_27958,N_29752);
xnor UO_2018 (O_2018,N_24675,N_24196);
nand UO_2019 (O_2019,N_26795,N_24483);
nor UO_2020 (O_2020,N_27917,N_28420);
or UO_2021 (O_2021,N_28578,N_27833);
nor UO_2022 (O_2022,N_25903,N_27647);
or UO_2023 (O_2023,N_26825,N_25105);
or UO_2024 (O_2024,N_26450,N_27611);
or UO_2025 (O_2025,N_24390,N_24988);
nor UO_2026 (O_2026,N_26197,N_28282);
xor UO_2027 (O_2027,N_26816,N_25072);
or UO_2028 (O_2028,N_26463,N_24457);
nor UO_2029 (O_2029,N_24998,N_27104);
nor UO_2030 (O_2030,N_29420,N_24362);
nor UO_2031 (O_2031,N_28399,N_26822);
or UO_2032 (O_2032,N_29038,N_26613);
or UO_2033 (O_2033,N_29210,N_25231);
and UO_2034 (O_2034,N_26826,N_28351);
nand UO_2035 (O_2035,N_25070,N_25472);
and UO_2036 (O_2036,N_29598,N_28163);
or UO_2037 (O_2037,N_24115,N_25115);
or UO_2038 (O_2038,N_24307,N_27447);
or UO_2039 (O_2039,N_29906,N_25764);
and UO_2040 (O_2040,N_29636,N_27286);
or UO_2041 (O_2041,N_26150,N_25007);
nand UO_2042 (O_2042,N_27846,N_29380);
nand UO_2043 (O_2043,N_25388,N_24663);
nand UO_2044 (O_2044,N_26474,N_26317);
nor UO_2045 (O_2045,N_26846,N_29541);
xor UO_2046 (O_2046,N_29745,N_25599);
and UO_2047 (O_2047,N_24715,N_27927);
nand UO_2048 (O_2048,N_26094,N_26077);
nor UO_2049 (O_2049,N_28428,N_26655);
nand UO_2050 (O_2050,N_26956,N_24412);
or UO_2051 (O_2051,N_28542,N_24375);
nand UO_2052 (O_2052,N_24906,N_26437);
or UO_2053 (O_2053,N_26253,N_29774);
nor UO_2054 (O_2054,N_27245,N_26561);
or UO_2055 (O_2055,N_24123,N_29220);
or UO_2056 (O_2056,N_26507,N_25000);
or UO_2057 (O_2057,N_25162,N_28804);
or UO_2058 (O_2058,N_26389,N_28593);
and UO_2059 (O_2059,N_24117,N_24909);
or UO_2060 (O_2060,N_27896,N_28703);
or UO_2061 (O_2061,N_27858,N_27462);
xnor UO_2062 (O_2062,N_29213,N_24242);
nand UO_2063 (O_2063,N_25006,N_27011);
and UO_2064 (O_2064,N_29275,N_29315);
xor UO_2065 (O_2065,N_25612,N_28323);
or UO_2066 (O_2066,N_25876,N_27390);
nand UO_2067 (O_2067,N_26948,N_26316);
nor UO_2068 (O_2068,N_24200,N_26572);
or UO_2069 (O_2069,N_24676,N_29224);
or UO_2070 (O_2070,N_26479,N_29908);
or UO_2071 (O_2071,N_25358,N_26012);
nand UO_2072 (O_2072,N_28206,N_24465);
nor UO_2073 (O_2073,N_28246,N_26100);
or UO_2074 (O_2074,N_25471,N_25681);
nor UO_2075 (O_2075,N_26169,N_29657);
or UO_2076 (O_2076,N_26943,N_27946);
nand UO_2077 (O_2077,N_29146,N_28866);
nor UO_2078 (O_2078,N_25822,N_29893);
nor UO_2079 (O_2079,N_24755,N_27817);
nor UO_2080 (O_2080,N_26276,N_28767);
or UO_2081 (O_2081,N_27899,N_24571);
nand UO_2082 (O_2082,N_29917,N_27473);
nor UO_2083 (O_2083,N_28834,N_28018);
nand UO_2084 (O_2084,N_27882,N_24476);
nand UO_2085 (O_2085,N_29364,N_29299);
or UO_2086 (O_2086,N_27490,N_26832);
nor UO_2087 (O_2087,N_26493,N_28733);
nand UO_2088 (O_2088,N_25614,N_29557);
and UO_2089 (O_2089,N_28236,N_25682);
xor UO_2090 (O_2090,N_28133,N_27285);
xnor UO_2091 (O_2091,N_28519,N_28597);
xor UO_2092 (O_2092,N_27943,N_26283);
and UO_2093 (O_2093,N_27684,N_28675);
nor UO_2094 (O_2094,N_26337,N_27630);
and UO_2095 (O_2095,N_25687,N_29735);
or UO_2096 (O_2096,N_24103,N_27335);
and UO_2097 (O_2097,N_29317,N_24772);
nand UO_2098 (O_2098,N_26307,N_26143);
xor UO_2099 (O_2099,N_27959,N_25633);
xor UO_2100 (O_2100,N_28195,N_26308);
nand UO_2101 (O_2101,N_29779,N_28166);
xor UO_2102 (O_2102,N_26322,N_27751);
nand UO_2103 (O_2103,N_27863,N_29122);
or UO_2104 (O_2104,N_26413,N_29209);
xor UO_2105 (O_2105,N_29952,N_24130);
and UO_2106 (O_2106,N_24585,N_24499);
nand UO_2107 (O_2107,N_29926,N_26213);
and UO_2108 (O_2108,N_29670,N_29085);
or UO_2109 (O_2109,N_28211,N_28910);
and UO_2110 (O_2110,N_27690,N_28559);
nor UO_2111 (O_2111,N_26306,N_28406);
and UO_2112 (O_2112,N_27391,N_27765);
and UO_2113 (O_2113,N_28546,N_29558);
nand UO_2114 (O_2114,N_25872,N_25896);
nand UO_2115 (O_2115,N_29314,N_28604);
and UO_2116 (O_2116,N_29427,N_26006);
nand UO_2117 (O_2117,N_25754,N_24638);
and UO_2118 (O_2118,N_28238,N_24341);
nor UO_2119 (O_2119,N_24422,N_29728);
nor UO_2120 (O_2120,N_27514,N_25615);
or UO_2121 (O_2121,N_25015,N_29677);
nor UO_2122 (O_2122,N_29034,N_27986);
and UO_2123 (O_2123,N_24302,N_24171);
nand UO_2124 (O_2124,N_25284,N_25914);
nor UO_2125 (O_2125,N_29703,N_28674);
or UO_2126 (O_2126,N_29379,N_27972);
nand UO_2127 (O_2127,N_26371,N_25587);
nand UO_2128 (O_2128,N_29748,N_26298);
nor UO_2129 (O_2129,N_28895,N_27079);
and UO_2130 (O_2130,N_29882,N_27738);
nor UO_2131 (O_2131,N_28247,N_29583);
and UO_2132 (O_2132,N_26071,N_28798);
and UO_2133 (O_2133,N_29321,N_26016);
or UO_2134 (O_2134,N_28939,N_29391);
nand UO_2135 (O_2135,N_25459,N_26195);
or UO_2136 (O_2136,N_24805,N_29251);
and UO_2137 (O_2137,N_28856,N_25950);
xnor UO_2138 (O_2138,N_25890,N_27264);
or UO_2139 (O_2139,N_27923,N_29881);
nor UO_2140 (O_2140,N_25319,N_24519);
or UO_2141 (O_2141,N_25157,N_27773);
or UO_2142 (O_2142,N_27696,N_26231);
nand UO_2143 (O_2143,N_26397,N_29831);
nor UO_2144 (O_2144,N_26106,N_24985);
nand UO_2145 (O_2145,N_25417,N_24616);
nand UO_2146 (O_2146,N_27301,N_24383);
nand UO_2147 (O_2147,N_29832,N_28366);
nand UO_2148 (O_2148,N_29279,N_28811);
and UO_2149 (O_2149,N_26177,N_27270);
or UO_2150 (O_2150,N_28177,N_27338);
nor UO_2151 (O_2151,N_29342,N_26014);
and UO_2152 (O_2152,N_25939,N_25260);
or UO_2153 (O_2153,N_26587,N_25649);
or UO_2154 (O_2154,N_25286,N_24544);
and UO_2155 (O_2155,N_26617,N_27193);
and UO_2156 (O_2156,N_29567,N_29932);
and UO_2157 (O_2157,N_26309,N_28012);
nor UO_2158 (O_2158,N_28868,N_28187);
nor UO_2159 (O_2159,N_26056,N_26641);
and UO_2160 (O_2160,N_29080,N_24459);
nor UO_2161 (O_2161,N_29110,N_28623);
and UO_2162 (O_2162,N_26629,N_27379);
or UO_2163 (O_2163,N_25753,N_27657);
or UO_2164 (O_2164,N_28204,N_26287);
nor UO_2165 (O_2165,N_28660,N_27693);
nand UO_2166 (O_2166,N_27915,N_25002);
or UO_2167 (O_2167,N_24174,N_25555);
nor UO_2168 (O_2168,N_24004,N_25210);
xor UO_2169 (O_2169,N_25194,N_27558);
or UO_2170 (O_2170,N_28491,N_28413);
and UO_2171 (O_2171,N_26873,N_27428);
and UO_2172 (O_2172,N_28452,N_26258);
nor UO_2173 (O_2173,N_25017,N_24068);
and UO_2174 (O_2174,N_24760,N_24248);
and UO_2175 (O_2175,N_25684,N_24611);
nand UO_2176 (O_2176,N_26342,N_24864);
and UO_2177 (O_2177,N_25771,N_28951);
or UO_2178 (O_2178,N_28598,N_25369);
nand UO_2179 (O_2179,N_29755,N_25207);
and UO_2180 (O_2180,N_27919,N_25922);
or UO_2181 (O_2181,N_26616,N_26794);
and UO_2182 (O_2182,N_29032,N_24129);
nor UO_2183 (O_2183,N_26300,N_27895);
and UO_2184 (O_2184,N_24972,N_27119);
and UO_2185 (O_2185,N_29109,N_25420);
nor UO_2186 (O_2186,N_28759,N_26881);
nor UO_2187 (O_2187,N_28216,N_28061);
nand UO_2188 (O_2188,N_26412,N_28948);
nand UO_2189 (O_2189,N_25995,N_29894);
or UO_2190 (O_2190,N_25673,N_26215);
and UO_2191 (O_2191,N_28965,N_25838);
or UO_2192 (O_2192,N_29361,N_26449);
nand UO_2193 (O_2193,N_28515,N_25377);
or UO_2194 (O_2194,N_29382,N_24841);
or UO_2195 (O_2195,N_29446,N_24618);
nand UO_2196 (O_2196,N_28300,N_25333);
nor UO_2197 (O_2197,N_25918,N_27319);
nor UO_2198 (O_2198,N_25425,N_26558);
nand UO_2199 (O_2199,N_25451,N_24743);
nand UO_2200 (O_2200,N_29323,N_24703);
nand UO_2201 (O_2201,N_28327,N_26174);
nand UO_2202 (O_2202,N_26486,N_27517);
nand UO_2203 (O_2203,N_29207,N_24898);
nand UO_2204 (O_2204,N_25250,N_27299);
xnor UO_2205 (O_2205,N_25671,N_27762);
nor UO_2206 (O_2206,N_28724,N_25487);
and UO_2207 (O_2207,N_26763,N_25761);
nor UO_2208 (O_2208,N_29934,N_26567);
and UO_2209 (O_2209,N_29239,N_25947);
nor UO_2210 (O_2210,N_28886,N_27096);
nand UO_2211 (O_2211,N_29818,N_26522);
nand UO_2212 (O_2212,N_26200,N_28590);
or UO_2213 (O_2213,N_24417,N_25266);
or UO_2214 (O_2214,N_26527,N_25536);
nor UO_2215 (O_2215,N_26742,N_26674);
or UO_2216 (O_2216,N_29806,N_29341);
and UO_2217 (O_2217,N_25816,N_27100);
nor UO_2218 (O_2218,N_26909,N_27146);
nor UO_2219 (O_2219,N_29868,N_26070);
or UO_2220 (O_2220,N_28359,N_25348);
and UO_2221 (O_2221,N_26749,N_29119);
or UO_2222 (O_2222,N_28387,N_28697);
nor UO_2223 (O_2223,N_28200,N_27576);
and UO_2224 (O_2224,N_24912,N_24019);
or UO_2225 (O_2225,N_29228,N_24927);
and UO_2226 (O_2226,N_24752,N_24283);
and UO_2227 (O_2227,N_27844,N_25533);
nand UO_2228 (O_2228,N_27516,N_29553);
and UO_2229 (O_2229,N_28762,N_24707);
nor UO_2230 (O_2230,N_26275,N_24414);
nor UO_2231 (O_2231,N_29078,N_25274);
nand UO_2232 (O_2232,N_28987,N_26243);
nor UO_2233 (O_2233,N_27271,N_28285);
and UO_2234 (O_2234,N_25711,N_27257);
nand UO_2235 (O_2235,N_24069,N_25654);
nand UO_2236 (O_2236,N_25393,N_29757);
or UO_2237 (O_2237,N_29330,N_27967);
nor UO_2238 (O_2238,N_29915,N_25329);
or UO_2239 (O_2239,N_29771,N_28008);
nor UO_2240 (O_2240,N_26348,N_27190);
nand UO_2241 (O_2241,N_29462,N_28734);
nor UO_2242 (O_2242,N_24058,N_29984);
nand UO_2243 (O_2243,N_24356,N_25644);
nor UO_2244 (O_2244,N_25983,N_28227);
nand UO_2245 (O_2245,N_27108,N_25449);
and UO_2246 (O_2246,N_29758,N_24627);
nor UO_2247 (O_2247,N_29600,N_24949);
xor UO_2248 (O_2248,N_26797,N_25811);
nand UO_2249 (O_2249,N_27618,N_24963);
and UO_2250 (O_2250,N_27259,N_25035);
nand UO_2251 (O_2251,N_27070,N_26959);
and UO_2252 (O_2252,N_25043,N_29889);
or UO_2253 (O_2253,N_24323,N_26049);
and UO_2254 (O_2254,N_27064,N_27659);
xor UO_2255 (O_2255,N_26152,N_25392);
and UO_2256 (O_2256,N_28257,N_29095);
xor UO_2257 (O_2257,N_29211,N_25031);
and UO_2258 (O_2258,N_27315,N_25139);
nand UO_2259 (O_2259,N_25421,N_24560);
nor UO_2260 (O_2260,N_28439,N_26719);
nand UO_2261 (O_2261,N_24857,N_24620);
nor UO_2262 (O_2262,N_26363,N_29886);
or UO_2263 (O_2263,N_29948,N_24084);
xor UO_2264 (O_2264,N_25427,N_28580);
and UO_2265 (O_2265,N_28240,N_25998);
and UO_2266 (O_2266,N_26569,N_26623);
nand UO_2267 (O_2267,N_26932,N_26761);
xnor UO_2268 (O_2268,N_27422,N_25964);
and UO_2269 (O_2269,N_27653,N_26136);
nor UO_2270 (O_2270,N_28958,N_27063);
nand UO_2271 (O_2271,N_26666,N_26005);
nand UO_2272 (O_2272,N_24971,N_25620);
nand UO_2273 (O_2273,N_27649,N_29528);
or UO_2274 (O_2274,N_24397,N_24834);
nor UO_2275 (O_2275,N_25452,N_26790);
nand UO_2276 (O_2276,N_24713,N_28250);
or UO_2277 (O_2277,N_28463,N_29967);
nor UO_2278 (O_2278,N_28015,N_26922);
or UO_2279 (O_2279,N_28360,N_28263);
nand UO_2280 (O_2280,N_24310,N_25669);
and UO_2281 (O_2281,N_26473,N_24968);
or UO_2282 (O_2282,N_29878,N_25440);
or UO_2283 (O_2283,N_25713,N_25648);
and UO_2284 (O_2284,N_24868,N_26067);
nand UO_2285 (O_2285,N_24745,N_28185);
xor UO_2286 (O_2286,N_26339,N_25874);
nor UO_2287 (O_2287,N_29448,N_29876);
and UO_2288 (O_2288,N_29518,N_26707);
and UO_2289 (O_2289,N_27793,N_28731);
xnor UO_2290 (O_2290,N_27092,N_25400);
xnor UO_2291 (O_2291,N_26052,N_28390);
or UO_2292 (O_2292,N_26695,N_28194);
or UO_2293 (O_2293,N_28098,N_25742);
and UO_2294 (O_2294,N_29971,N_25455);
or UO_2295 (O_2295,N_24714,N_29665);
nand UO_2296 (O_2296,N_27672,N_25566);
nor UO_2297 (O_2297,N_26920,N_28244);
and UO_2298 (O_2298,N_26379,N_24332);
xnor UO_2299 (O_2299,N_27231,N_29584);
xnor UO_2300 (O_2300,N_25152,N_24520);
nand UO_2301 (O_2301,N_28092,N_25997);
nor UO_2302 (O_2302,N_28981,N_24493);
xnor UO_2303 (O_2303,N_29609,N_28063);
nand UO_2304 (O_2304,N_26133,N_26730);
xnor UO_2305 (O_2305,N_28027,N_24728);
nand UO_2306 (O_2306,N_25625,N_29337);
nand UO_2307 (O_2307,N_29076,N_27550);
xor UO_2308 (O_2308,N_25486,N_26788);
nand UO_2309 (O_2309,N_28699,N_26793);
nand UO_2310 (O_2310,N_27559,N_29568);
or UO_2311 (O_2311,N_28241,N_26395);
nor UO_2312 (O_2312,N_28332,N_28460);
nor UO_2313 (O_2313,N_24497,N_29860);
nor UO_2314 (O_2314,N_27726,N_28645);
nand UO_2315 (O_2315,N_28727,N_26430);
or UO_2316 (O_2316,N_28472,N_25047);
or UO_2317 (O_2317,N_29425,N_29044);
nand UO_2318 (O_2318,N_28763,N_29538);
nor UO_2319 (O_2319,N_25655,N_29941);
or UO_2320 (O_2320,N_26373,N_29700);
xnor UO_2321 (O_2321,N_26098,N_28132);
nor UO_2322 (O_2322,N_29650,N_25716);
nand UO_2323 (O_2323,N_29437,N_26673);
or UO_2324 (O_2324,N_26446,N_28036);
nor UO_2325 (O_2325,N_24042,N_27871);
and UO_2326 (O_2326,N_26799,N_27278);
nor UO_2327 (O_2327,N_25795,N_29283);
nor UO_2328 (O_2328,N_25973,N_26901);
and UO_2329 (O_2329,N_27238,N_24996);
nand UO_2330 (O_2330,N_24719,N_25147);
or UO_2331 (O_2331,N_26217,N_27861);
xor UO_2332 (O_2332,N_28029,N_24259);
nand UO_2333 (O_2333,N_29564,N_26980);
xor UO_2334 (O_2334,N_28202,N_25456);
or UO_2335 (O_2335,N_24883,N_25977);
nand UO_2336 (O_2336,N_25022,N_29887);
nand UO_2337 (O_2337,N_28127,N_25410);
and UO_2338 (O_2338,N_25927,N_25298);
nor UO_2339 (O_2339,N_25294,N_24243);
or UO_2340 (O_2340,N_25405,N_27794);
xor UO_2341 (O_2341,N_27083,N_24072);
nor UO_2342 (O_2342,N_28447,N_24820);
or UO_2343 (O_2343,N_29592,N_25630);
nand UO_2344 (O_2344,N_29506,N_24513);
nor UO_2345 (O_2345,N_29659,N_25282);
or UO_2346 (O_2346,N_25537,N_24926);
nand UO_2347 (O_2347,N_27372,N_29455);
and UO_2348 (O_2348,N_27015,N_28284);
and UO_2349 (O_2349,N_27699,N_27246);
or UO_2350 (O_2350,N_24118,N_28471);
nor UO_2351 (O_2351,N_25224,N_25894);
nor UO_2352 (O_2352,N_29624,N_27779);
nand UO_2353 (O_2353,N_25373,N_26320);
and UO_2354 (O_2354,N_24773,N_27395);
or UO_2355 (O_2355,N_27412,N_24252);
or UO_2356 (O_2356,N_29295,N_24564);
or UO_2357 (O_2357,N_28730,N_29740);
and UO_2358 (O_2358,N_25933,N_27351);
nand UO_2359 (O_2359,N_29166,N_27221);
nand UO_2360 (O_2360,N_29859,N_28915);
or UO_2361 (O_2361,N_25199,N_25488);
nand UO_2362 (O_2362,N_24247,N_27854);
or UO_2363 (O_2363,N_25623,N_28110);
xnor UO_2364 (O_2364,N_24696,N_29607);
and UO_2365 (O_2365,N_25414,N_29236);
or UO_2366 (O_2366,N_28557,N_27801);
nor UO_2367 (O_2367,N_26018,N_27388);
nand UO_2368 (O_2368,N_24992,N_28273);
or UO_2369 (O_2369,N_27061,N_26789);
nor UO_2370 (O_2370,N_28180,N_29672);
nand UO_2371 (O_2371,N_29192,N_27499);
nor UO_2372 (O_2372,N_24273,N_28489);
and UO_2373 (O_2373,N_25762,N_26708);
or UO_2374 (O_2374,N_27585,N_24827);
and UO_2375 (O_2375,N_29348,N_29286);
or UO_2376 (O_2376,N_24810,N_25347);
nor UO_2377 (O_2377,N_24214,N_28957);
nor UO_2378 (O_2378,N_27501,N_27397);
or UO_2379 (O_2379,N_29922,N_29880);
nor UO_2380 (O_2380,N_28032,N_26461);
nor UO_2381 (O_2381,N_24801,N_27572);
or UO_2382 (O_2382,N_26762,N_24811);
nand UO_2383 (O_2383,N_26537,N_26113);
or UO_2384 (O_2384,N_26448,N_29770);
or UO_2385 (O_2385,N_24083,N_24844);
nor UO_2386 (O_2386,N_26916,N_28287);
and UO_2387 (O_2387,N_27220,N_29873);
and UO_2388 (O_2388,N_27343,N_29047);
or UO_2389 (O_2389,N_24605,N_28787);
nor UO_2390 (O_2390,N_24958,N_24794);
nor UO_2391 (O_2391,N_25464,N_28045);
and UO_2392 (O_2392,N_24692,N_27593);
nand UO_2393 (O_2393,N_29360,N_25852);
or UO_2394 (O_2394,N_24865,N_28007);
nand UO_2395 (O_2395,N_25149,N_24691);
and UO_2396 (O_2396,N_24318,N_28335);
and UO_2397 (O_2397,N_24251,N_25469);
nand UO_2398 (O_2398,N_27229,N_24784);
or UO_2399 (O_2399,N_27596,N_25053);
or UO_2400 (O_2400,N_24399,N_24300);
or UO_2401 (O_2401,N_28249,N_26433);
nand UO_2402 (O_2402,N_27060,N_25900);
or UO_2403 (O_2403,N_29987,N_28512);
nand UO_2404 (O_2404,N_28160,N_24939);
or UO_2405 (O_2405,N_27191,N_28433);
nor UO_2406 (O_2406,N_27235,N_25466);
nor UO_2407 (O_2407,N_27906,N_25968);
and UO_2408 (O_2408,N_28887,N_24090);
or UO_2409 (O_2409,N_26682,N_29204);
nand UO_2410 (O_2410,N_29016,N_25275);
or UO_2411 (O_2411,N_24011,N_27485);
or UO_2412 (O_2412,N_25131,N_26568);
nand UO_2413 (O_2413,N_29180,N_27232);
or UO_2414 (O_2414,N_25173,N_28305);
or UO_2415 (O_2415,N_27463,N_27095);
or UO_2416 (O_2416,N_28945,N_26185);
nor UO_2417 (O_2417,N_28089,N_24870);
or UO_2418 (O_2418,N_25796,N_26246);
or UO_2419 (O_2419,N_27178,N_27253);
nand UO_2420 (O_2420,N_27263,N_26622);
and UO_2421 (O_2421,N_29990,N_29823);
nand UO_2422 (O_2422,N_29722,N_25470);
xnor UO_2423 (O_2423,N_25975,N_29469);
nor UO_2424 (O_2424,N_25656,N_27432);
and UO_2425 (O_2425,N_24468,N_27135);
nor UO_2426 (O_2426,N_27904,N_29759);
nand UO_2427 (O_2427,N_26033,N_27406);
nand UO_2428 (O_2428,N_25462,N_26099);
nor UO_2429 (O_2429,N_25700,N_25790);
nor UO_2430 (O_2430,N_28498,N_25827);
and UO_2431 (O_2431,N_24881,N_26758);
xnor UO_2432 (O_2432,N_25021,N_28736);
nand UO_2433 (O_2433,N_28141,N_24388);
and UO_2434 (O_2434,N_24974,N_28013);
xor UO_2435 (O_2435,N_24139,N_26202);
nor UO_2436 (O_2436,N_26155,N_29276);
nor UO_2437 (O_2437,N_25588,N_25910);
xor UO_2438 (O_2438,N_26775,N_29481);
xnor UO_2439 (O_2439,N_25267,N_25382);
or UO_2440 (O_2440,N_27588,N_29240);
nand UO_2441 (O_2441,N_26154,N_24223);
nor UO_2442 (O_2442,N_24146,N_24460);
nand UO_2443 (O_2443,N_25316,N_29496);
and UO_2444 (O_2444,N_29678,N_28159);
or UO_2445 (O_2445,N_28214,N_29545);
nand UO_2446 (O_2446,N_29048,N_24732);
nor UO_2447 (O_2447,N_28896,N_28389);
or UO_2448 (O_2448,N_27443,N_27460);
and UO_2449 (O_2449,N_25415,N_25151);
and UO_2450 (O_2450,N_26267,N_28658);
nand UO_2451 (O_2451,N_26810,N_26745);
or UO_2452 (O_2452,N_29113,N_26781);
or UO_2453 (O_2453,N_28056,N_26626);
and UO_2454 (O_2454,N_28484,N_27787);
or UO_2455 (O_2455,N_28298,N_24439);
nand UO_2456 (O_2456,N_26428,N_29879);
and UO_2457 (O_2457,N_28698,N_26535);
or UO_2458 (O_2458,N_26230,N_25543);
nor UO_2459 (O_2459,N_28844,N_24789);
nand UO_2460 (O_2460,N_29421,N_27371);
and UO_2461 (O_2461,N_29092,N_26063);
nand UO_2462 (O_2462,N_28436,N_26918);
or UO_2463 (O_2463,N_29577,N_29306);
and UO_2464 (O_2464,N_29550,N_24257);
nor UO_2465 (O_2465,N_26954,N_26496);
nor UO_2466 (O_2466,N_29397,N_27101);
and UO_2467 (O_2467,N_28929,N_24830);
and UO_2468 (O_2468,N_27316,N_29130);
and UO_2469 (O_2469,N_29002,N_27326);
nor UO_2470 (O_2470,N_29772,N_29375);
xnor UO_2471 (O_2471,N_27248,N_26608);
or UO_2472 (O_2472,N_28752,N_26946);
or UO_2473 (O_2473,N_25938,N_27359);
nand UO_2474 (O_2474,N_26264,N_28871);
nand UO_2475 (O_2475,N_26162,N_26023);
nor UO_2476 (O_2476,N_25318,N_25349);
and UO_2477 (O_2477,N_24584,N_25819);
xor UO_2478 (O_2478,N_25171,N_27347);
and UO_2479 (O_2479,N_27344,N_26713);
nand UO_2480 (O_2480,N_27807,N_26384);
or UO_2481 (O_2481,N_24837,N_27748);
and UO_2482 (O_2482,N_28664,N_27491);
nor UO_2483 (O_2483,N_25925,N_28611);
nand UO_2484 (O_2484,N_24981,N_25080);
or UO_2485 (O_2485,N_25993,N_29514);
xor UO_2486 (O_2486,N_26919,N_25264);
or UO_2487 (O_2487,N_25663,N_27808);
and UO_2488 (O_2488,N_24816,N_26314);
and UO_2489 (O_2489,N_28197,N_28640);
xor UO_2490 (O_2490,N_24007,N_28998);
nand UO_2491 (O_2491,N_25942,N_29172);
nor UO_2492 (O_2492,N_28171,N_25854);
or UO_2493 (O_2493,N_25785,N_26203);
nor UO_2494 (O_2494,N_25705,N_24680);
nor UO_2495 (O_2495,N_29765,N_27938);
nor UO_2496 (O_2496,N_25677,N_28541);
nor UO_2497 (O_2497,N_24325,N_28794);
or UO_2498 (O_2498,N_25955,N_28709);
or UO_2499 (O_2499,N_29924,N_26375);
nor UO_2500 (O_2500,N_26199,N_27421);
xnor UO_2501 (O_2501,N_24191,N_25376);
nor UO_2502 (O_2502,N_25529,N_29682);
and UO_2503 (O_2503,N_26667,N_26029);
nand UO_2504 (O_2504,N_27323,N_24609);
and UO_2505 (O_2505,N_25772,N_24942);
nand UO_2506 (O_2506,N_24461,N_29676);
nor UO_2507 (O_2507,N_28902,N_28812);
and UO_2508 (O_2508,N_25494,N_28914);
nand UO_2509 (O_2509,N_26836,N_25744);
and UO_2510 (O_2510,N_29701,N_25201);
and UO_2511 (O_2511,N_25359,N_25944);
nor UO_2512 (O_2512,N_28687,N_26521);
nor UO_2513 (O_2513,N_25125,N_26242);
and UO_2514 (O_2514,N_29398,N_29231);
or UO_2515 (O_2515,N_29368,N_24105);
xor UO_2516 (O_2516,N_24201,N_24646);
or UO_2517 (O_2517,N_25197,N_26917);
nand UO_2518 (O_2518,N_29145,N_24599);
and UO_2519 (O_2519,N_27317,N_26454);
nand UO_2520 (O_2520,N_24746,N_26193);
or UO_2521 (O_2521,N_29639,N_24946);
xor UO_2522 (O_2522,N_24737,N_25593);
or UO_2523 (O_2523,N_27626,N_28259);
nor UO_2524 (O_2524,N_24054,N_24093);
or UO_2525 (O_2525,N_24204,N_29939);
nand UO_2526 (O_2526,N_29726,N_24168);
xor UO_2527 (O_2527,N_28616,N_29746);
and UO_2528 (O_2528,N_25177,N_29495);
nand UO_2529 (O_2529,N_25100,N_25851);
nor UO_2530 (O_2530,N_24317,N_29229);
or UO_2531 (O_2531,N_27198,N_27160);
nor UO_2532 (O_2532,N_26942,N_25170);
nor UO_2533 (O_2533,N_24391,N_28681);
nor UO_2534 (O_2534,N_24432,N_26914);
and UO_2535 (O_2535,N_29612,N_26827);
nand UO_2536 (O_2536,N_28786,N_29031);
nor UO_2537 (O_2537,N_27172,N_25558);
and UO_2538 (O_2538,N_29066,N_27309);
xor UO_2539 (O_2539,N_28475,N_26969);
or UO_2540 (O_2540,N_24653,N_27042);
or UO_2541 (O_2541,N_29225,N_28743);
and UO_2542 (O_2542,N_28619,N_29023);
and UO_2543 (O_2543,N_27189,N_24739);
or UO_2544 (O_2544,N_26882,N_26432);
nor UO_2545 (O_2545,N_29843,N_24395);
nand UO_2546 (O_2546,N_24225,N_29706);
or UO_2547 (O_2547,N_27016,N_27433);
nand UO_2548 (O_2548,N_24779,N_28304);
nor UO_2549 (O_2549,N_25389,N_29750);
nand UO_2550 (O_2550,N_28680,N_25403);
or UO_2551 (O_2551,N_24582,N_26201);
xnor UO_2552 (O_2552,N_26647,N_29041);
xnor UO_2553 (O_2553,N_25090,N_28634);
and UO_2554 (O_2554,N_27471,N_24647);
and UO_2555 (O_2555,N_27834,N_26343);
or UO_2556 (O_2556,N_29742,N_29103);
nand UO_2557 (O_2557,N_24702,N_26069);
xnor UO_2558 (O_2558,N_26013,N_28725);
or UO_2559 (O_2559,N_29353,N_28906);
nand UO_2560 (O_2560,N_24305,N_25276);
nand UO_2561 (O_2561,N_25966,N_25409);
nand UO_2562 (O_2562,N_29715,N_26575);
nor UO_2563 (O_2563,N_25012,N_28364);
or UO_2564 (O_2564,N_26945,N_28695);
xnor UO_2565 (O_2565,N_28810,N_29912);
and UO_2566 (O_2566,N_26774,N_26975);
xor UO_2567 (O_2567,N_26290,N_25430);
xnor UO_2568 (O_2568,N_24138,N_24579);
nor UO_2569 (O_2569,N_27358,N_27260);
and UO_2570 (O_2570,N_25465,N_28336);
or UO_2571 (O_2571,N_28253,N_26974);
nand UO_2572 (O_2572,N_29265,N_29232);
nand UO_2573 (O_2573,N_27489,N_28773);
and UO_2574 (O_2574,N_28217,N_28530);
and UO_2575 (O_2575,N_25384,N_24109);
nand UO_2576 (O_2576,N_26190,N_24298);
xor UO_2577 (O_2577,N_26282,N_26206);
and UO_2578 (O_2578,N_27056,N_26725);
nor UO_2579 (O_2579,N_29804,N_25913);
nor UO_2580 (O_2580,N_29834,N_27266);
and UO_2581 (O_2581,N_29070,N_26601);
nor UO_2582 (O_2582,N_28571,N_28136);
xor UO_2583 (O_2583,N_25770,N_29269);
and UO_2584 (O_2584,N_27069,N_24458);
nand UO_2585 (O_2585,N_29872,N_28383);
or UO_2586 (O_2586,N_26398,N_25356);
nor UO_2587 (O_2587,N_27223,N_25820);
nor UO_2588 (O_2588,N_24894,N_24589);
or UO_2589 (O_2589,N_29966,N_24873);
nand UO_2590 (O_2590,N_24524,N_29234);
and UO_2591 (O_2591,N_27889,N_25119);
or UO_2592 (O_2592,N_28181,N_28853);
xnor UO_2593 (O_2593,N_28321,N_29803);
or UO_2594 (O_2594,N_26090,N_28926);
nor UO_2595 (O_2595,N_24853,N_25520);
or UO_2596 (O_2596,N_29243,N_25689);
xnor UO_2597 (O_2597,N_26506,N_25111);
nor UO_2598 (O_2598,N_28169,N_29370);
nor UO_2599 (O_2599,N_27496,N_26638);
xnor UO_2600 (O_2600,N_28857,N_28066);
or UO_2601 (O_2601,N_27935,N_26132);
or UO_2602 (O_2602,N_29788,N_25225);
nand UO_2603 (O_2603,N_27843,N_24057);
or UO_2604 (O_2604,N_25592,N_25961);
nor UO_2605 (O_2605,N_29738,N_27149);
and UO_2606 (O_2606,N_29862,N_28930);
nand UO_2607 (O_2607,N_26903,N_28603);
nor UO_2608 (O_2608,N_29334,N_26904);
and UO_2609 (O_2609,N_29280,N_26783);
or UO_2610 (O_2610,N_25094,N_26062);
nor UO_2611 (O_2611,N_28270,N_26853);
and UO_2612 (O_2612,N_29957,N_24501);
or UO_2613 (O_2613,N_28224,N_29576);
nand UO_2614 (O_2614,N_28088,N_28540);
and UO_2615 (O_2615,N_27186,N_29021);
or UO_2616 (O_2616,N_29780,N_29489);
and UO_2617 (O_2617,N_28201,N_27595);
or UO_2618 (O_2618,N_25548,N_28000);
nand UO_2619 (O_2619,N_27226,N_28086);
and UO_2620 (O_2620,N_25018,N_24979);
and UO_2621 (O_2621,N_25370,N_29274);
nand UO_2622 (O_2622,N_25351,N_24768);
nand UO_2623 (O_2623,N_24181,N_27038);
nor UO_2624 (O_2624,N_27320,N_28831);
nand UO_2625 (O_2625,N_25212,N_25812);
nor UO_2626 (O_2626,N_24659,N_24836);
or UO_2627 (O_2627,N_29158,N_27984);
nor UO_2628 (O_2628,N_24098,N_27681);
or UO_2629 (O_2629,N_27847,N_28353);
nor UO_2630 (O_2630,N_26546,N_29169);
nand UO_2631 (O_2631,N_24863,N_27054);
and UO_2632 (O_2632,N_26256,N_29294);
and UO_2633 (O_2633,N_26421,N_26266);
nand UO_2634 (O_2634,N_26284,N_28973);
or UO_2635 (O_2635,N_29684,N_26744);
nor UO_2636 (O_2636,N_27898,N_26502);
and UO_2637 (O_2637,N_29339,N_25187);
nor UO_2638 (O_2638,N_27321,N_29428);
and UO_2639 (O_2639,N_27760,N_24194);
nor UO_2640 (O_2640,N_24557,N_27129);
nor UO_2641 (O_2641,N_24919,N_28427);
and UO_2642 (O_2642,N_27545,N_28434);
or UO_2643 (O_2643,N_25323,N_26967);
xor UO_2644 (O_2644,N_27835,N_28772);
and UO_2645 (O_2645,N_26399,N_27155);
nor UO_2646 (O_2646,N_26979,N_27442);
nor UO_2647 (O_2647,N_25308,N_28316);
or UO_2648 (O_2648,N_27000,N_26553);
and UO_2649 (O_2649,N_28084,N_24817);
and UO_2650 (O_2650,N_29871,N_25206);
or UO_2651 (O_2651,N_29302,N_24452);
or UO_2652 (O_2652,N_27147,N_25428);
nand UO_2653 (O_2653,N_28704,N_25345);
or UO_2654 (O_2654,N_29049,N_26689);
nor UO_2655 (O_2655,N_29712,N_25096);
and UO_2656 (O_2656,N_26627,N_27394);
and UO_2657 (O_2657,N_29666,N_27110);
and UO_2658 (O_2658,N_26350,N_27734);
nand UO_2659 (O_2659,N_27910,N_26704);
nor UO_2660 (O_2660,N_26640,N_24783);
or UO_2661 (O_2661,N_25769,N_26101);
nor UO_2662 (O_2662,N_26859,N_27481);
nor UO_2663 (O_2663,N_28518,N_24845);
or UO_2664 (O_2664,N_28102,N_28994);
nand UO_2665 (O_2665,N_27548,N_29009);
nand UO_2666 (O_2666,N_28971,N_29200);
nor UO_2667 (O_2667,N_27167,N_28544);
nor UO_2668 (O_2668,N_26864,N_25476);
and UO_2669 (O_2669,N_29744,N_27296);
xnor UO_2670 (O_2670,N_29268,N_26594);
nor UO_2671 (O_2671,N_29784,N_25108);
xor UO_2672 (O_2672,N_28784,N_29605);
nor UO_2673 (O_2673,N_26186,N_24851);
nand UO_2674 (O_2674,N_24485,N_29013);
nor UO_2675 (O_2675,N_26353,N_27697);
nor UO_2676 (O_2676,N_29285,N_28826);
nand UO_2677 (O_2677,N_25255,N_24554);
or UO_2678 (O_2678,N_24464,N_26990);
xnor UO_2679 (O_2679,N_28970,N_25722);
nand UO_2680 (O_2680,N_29534,N_25573);
nor UO_2681 (O_2681,N_27362,N_26156);
or UO_2682 (O_2682,N_24941,N_27528);
nor UO_2683 (O_2683,N_25395,N_25216);
nand UO_2684 (O_2684,N_29743,N_24153);
nor UO_2685 (O_2685,N_24984,N_26855);
or UO_2686 (O_2686,N_28800,N_28050);
or UO_2687 (O_2687,N_26295,N_29189);
nor UO_2688 (O_2688,N_28286,N_28878);
or UO_2689 (O_2689,N_29365,N_26015);
or UO_2690 (O_2690,N_25957,N_24886);
xnor UO_2691 (O_2691,N_24950,N_27758);
or UO_2692 (O_2692,N_29083,N_25696);
and UO_2693 (O_2693,N_26092,N_27931);
and UO_2694 (O_2694,N_28815,N_25394);
and UO_2695 (O_2695,N_29216,N_27540);
xnor UO_2696 (O_2696,N_24867,N_29956);
and UO_2697 (O_2697,N_27380,N_28663);
nand UO_2698 (O_2698,N_25511,N_28852);
and UO_2699 (O_2699,N_25324,N_26841);
nand UO_2700 (O_2700,N_29161,N_25940);
and UO_2701 (O_2701,N_28229,N_27099);
nand UO_2702 (O_2702,N_29388,N_29985);
xor UO_2703 (O_2703,N_26768,N_29426);
or UO_2704 (O_2704,N_25688,N_28373);
and UO_2705 (O_2705,N_26417,N_24595);
nor UO_2706 (O_2706,N_26701,N_25133);
nand UO_2707 (O_2707,N_28690,N_26839);
or UO_2708 (O_2708,N_25186,N_27712);
nor UO_2709 (O_2709,N_28199,N_26576);
nand UO_2710 (O_2710,N_25921,N_27387);
xnor UO_2711 (O_2711,N_24282,N_26688);
or UO_2712 (O_2712,N_24597,N_28742);
nor UO_2713 (O_2713,N_27291,N_26815);
and UO_2714 (O_2714,N_28669,N_28041);
xnor UO_2715 (O_2715,N_27161,N_27674);
or UO_2716 (O_2716,N_28299,N_28182);
xnor UO_2717 (O_2717,N_25823,N_25337);
nand UO_2718 (O_2718,N_25192,N_29786);
and UO_2719 (O_2719,N_29658,N_28806);
nor UO_2720 (O_2720,N_27459,N_25568);
xnor UO_2721 (O_2721,N_28691,N_27859);
nor UO_2722 (O_2722,N_26127,N_26722);
nand UO_2723 (O_2723,N_28648,N_25121);
and UO_2724 (O_2724,N_26669,N_24236);
or UO_2725 (O_2725,N_24052,N_26001);
nor UO_2726 (O_2726,N_26828,N_28501);
or UO_2727 (O_2727,N_26985,N_26877);
nor UO_2728 (O_2728,N_25081,N_26356);
nand UO_2729 (O_2729,N_27669,N_26490);
or UO_2730 (O_2730,N_29951,N_27053);
nor UO_2731 (O_2731,N_28624,N_29033);
or UO_2732 (O_2732,N_25830,N_24413);
or UO_2733 (O_2733,N_28070,N_28379);
or UO_2734 (O_2734,N_25583,N_24241);
nand UO_2735 (O_2735,N_26539,N_29808);
nor UO_2736 (O_2736,N_24363,N_28720);
or UO_2737 (O_2737,N_28192,N_24346);
nor UO_2738 (O_2738,N_24148,N_29864);
or UO_2739 (O_2739,N_26944,N_28046);
nor UO_2740 (O_2740,N_27781,N_24517);
nand UO_2741 (O_2741,N_25951,N_28750);
or UO_2742 (O_2742,N_25195,N_29835);
nand UO_2743 (O_2743,N_26387,N_24651);
and UO_2744 (O_2744,N_27592,N_28775);
or UO_2745 (O_2745,N_27312,N_24484);
nor UO_2746 (O_2746,N_24338,N_26401);
nor UO_2747 (O_2747,N_26058,N_24134);
xnor UO_2748 (O_2748,N_25217,N_26409);
xor UO_2749 (O_2749,N_29215,N_26656);
and UO_2750 (O_2750,N_28302,N_29529);
nand UO_2751 (O_2751,N_25124,N_27062);
nor UO_2752 (O_2752,N_28222,N_26447);
and UO_2753 (O_2753,N_29488,N_26407);
xor UO_2754 (O_2754,N_27627,N_26834);
nor UO_2755 (O_2755,N_25557,N_29839);
and UO_2756 (O_2756,N_26648,N_27120);
and UO_2757 (O_2757,N_24877,N_25665);
or UO_2758 (O_2758,N_28714,N_26896);
nor UO_2759 (O_2759,N_26064,N_28883);
xor UO_2760 (O_2760,N_24770,N_29320);
and UO_2761 (O_2761,N_26109,N_24612);
and UO_2762 (O_2762,N_26723,N_25603);
and UO_2763 (O_2763,N_26748,N_24839);
nand UO_2764 (O_2764,N_24966,N_26239);
and UO_2765 (O_2765,N_26378,N_26254);
and UO_2766 (O_2766,N_24246,N_28643);
nor UO_2767 (O_2767,N_28897,N_25865);
or UO_2768 (O_2768,N_28347,N_25737);
nand UO_2769 (O_2769,N_25651,N_29399);
or UO_2770 (O_2770,N_27302,N_29069);
xor UO_2771 (O_2771,N_28539,N_27533);
nand UO_2772 (O_2772,N_27228,N_27547);
and UO_2773 (O_2773,N_27900,N_29891);
xor UO_2774 (O_2774,N_29396,N_24227);
and UO_2775 (O_2775,N_26574,N_24569);
or UO_2776 (O_2776,N_28789,N_26327);
nor UO_2777 (O_2777,N_28668,N_27225);
and UO_2778 (O_2778,N_24445,N_28477);
or UO_2779 (O_2779,N_24135,N_24819);
or UO_2780 (O_2780,N_24548,N_29493);
nand UO_2781 (O_2781,N_27947,N_26087);
nor UO_2782 (O_2782,N_25134,N_29176);
or UO_2783 (O_2783,N_28997,N_28861);
nand UO_2784 (O_2784,N_26476,N_27217);
nor UO_2785 (O_2785,N_27294,N_25676);
and UO_2786 (O_2786,N_25050,N_28444);
or UO_2787 (O_2787,N_28527,N_24370);
nand UO_2788 (O_2788,N_27717,N_25495);
nand UO_2789 (O_2789,N_28306,N_24449);
or UO_2790 (O_2790,N_28451,N_29573);
xnor UO_2791 (O_2791,N_25445,N_26324);
nand UO_2792 (O_2792,N_28115,N_29965);
nor UO_2793 (O_2793,N_29733,N_29153);
nor UO_2794 (O_2794,N_26564,N_25429);
or UO_2795 (O_2795,N_27867,N_28147);
xor UO_2796 (O_2796,N_25479,N_25802);
or UO_2797 (O_2797,N_25016,N_28764);
or UO_2798 (O_2798,N_26515,N_26469);
and UO_2799 (O_2799,N_28547,N_28529);
nor UO_2800 (O_2800,N_24089,N_28933);
or UO_2801 (O_2801,N_26214,N_26175);
nand UO_2802 (O_2802,N_28586,N_27928);
nand UO_2803 (O_2803,N_26577,N_29264);
nor UO_2804 (O_2804,N_27476,N_28320);
and UO_2805 (O_2805,N_24081,N_25036);
nand UO_2806 (O_2806,N_26526,N_24993);
and UO_2807 (O_2807,N_28189,N_25530);
and UO_2808 (O_2808,N_24761,N_29620);
nand UO_2809 (O_2809,N_27204,N_26581);
and UO_2810 (O_2810,N_24764,N_26112);
xnor UO_2811 (O_2811,N_28193,N_25883);
xnor UO_2812 (O_2812,N_28990,N_24116);
nand UO_2813 (O_2813,N_28792,N_25262);
nand UO_2814 (O_2814,N_27602,N_27140);
nand UO_2815 (O_2815,N_28314,N_29622);
or UO_2816 (O_2816,N_24315,N_24230);
or UO_2817 (O_2817,N_24928,N_29447);
nor UO_2818 (O_2818,N_26743,N_28889);
or UO_2819 (O_2819,N_28276,N_26313);
or UO_2820 (O_2820,N_28377,N_29344);
xnor UO_2821 (O_2821,N_29896,N_24416);
and UO_2822 (O_2822,N_29001,N_27905);
xnor UO_2823 (O_2823,N_29096,N_25974);
or UO_2824 (O_2824,N_26488,N_29472);
or UO_2825 (O_2825,N_27008,N_25721);
nor UO_2826 (O_2826,N_24673,N_25502);
nor UO_2827 (O_2827,N_26365,N_29699);
and UO_2828 (O_2828,N_27671,N_25509);
and UO_2829 (O_2829,N_27114,N_24076);
nor UO_2830 (O_2830,N_29051,N_26038);
or UO_2831 (O_2831,N_27169,N_27065);
nand UO_2832 (O_2832,N_27874,N_28835);
xnor UO_2833 (O_2833,N_26739,N_25672);
nand UO_2834 (O_2834,N_26878,N_29343);
or UO_2835 (O_2835,N_25256,N_29962);
xnor UO_2836 (O_2836,N_29193,N_24833);
nand UO_2837 (O_2837,N_27339,N_29471);
nor UO_2838 (O_2838,N_24891,N_26170);
or UO_2839 (O_2839,N_26426,N_28959);
xor UO_2840 (O_2840,N_27192,N_29884);
nand UO_2841 (O_2841,N_27894,N_25132);
or UO_2842 (O_2842,N_25634,N_27637);
or UO_2843 (O_2843,N_26782,N_27243);
or UO_2844 (O_2844,N_28034,N_25847);
or UO_2845 (O_2845,N_28516,N_28735);
and UO_2846 (O_2846,N_28442,N_24475);
or UO_2847 (O_2847,N_24880,N_26929);
nor UO_2848 (O_2848,N_28131,N_29560);
nor UO_2849 (O_2849,N_26962,N_28666);
nand UO_2850 (O_2850,N_27024,N_24095);
and UO_2851 (O_2851,N_26158,N_28121);
xnor UO_2852 (O_2852,N_28932,N_25245);
nand UO_2853 (O_2853,N_28717,N_27201);
or UO_2854 (O_2854,N_25003,N_29905);
and UO_2855 (O_2855,N_29301,N_28574);
nor UO_2856 (O_2856,N_28233,N_28090);
xor UO_2857 (O_2857,N_28097,N_27132);
nand UO_2858 (O_2858,N_25513,N_28816);
nand UO_2859 (O_2859,N_29727,N_26595);
nand UO_2860 (O_2860,N_27512,N_27719);
and UO_2861 (O_2861,N_24043,N_26129);
and UO_2862 (O_2862,N_29791,N_24566);
and UO_2863 (O_2863,N_28901,N_26817);
or UO_2864 (O_2864,N_29208,N_29246);
and UO_2865 (O_2865,N_28797,N_28916);
nand UO_2866 (O_2866,N_27539,N_26542);
nor UO_2867 (O_2867,N_29515,N_26059);
nand UO_2868 (O_2868,N_24261,N_24785);
and UO_2869 (O_2869,N_29594,N_27211);
nand UO_2870 (O_2870,N_25034,N_25717);
nor UO_2871 (O_2871,N_27727,N_29913);
nor UO_2872 (O_2872,N_26562,N_24473);
or UO_2873 (O_2873,N_27881,N_24710);
nor UO_2874 (O_2874,N_29223,N_27196);
and UO_2875 (O_2875,N_26683,N_24335);
nor UO_2876 (O_2876,N_29946,N_24424);
nor UO_2877 (O_2877,N_29817,N_25779);
or UO_2878 (O_2878,N_27578,N_24260);
nand UO_2879 (O_2879,N_28647,N_25233);
xor UO_2880 (O_2880,N_28903,N_27842);
or UO_2881 (O_2881,N_24158,N_24577);
nand UO_2882 (O_2882,N_29257,N_27117);
and UO_2883 (O_2883,N_29943,N_27675);
or UO_2884 (O_2884,N_28234,N_25326);
nand UO_2885 (O_2885,N_27710,N_29767);
nand UO_2886 (O_2886,N_26443,N_27336);
or UO_2887 (O_2887,N_28125,N_29944);
xnor UO_2888 (O_2888,N_25846,N_25719);
or UO_2889 (O_2889,N_25781,N_27268);
nor UO_2890 (O_2890,N_26119,N_24024);
nor UO_2891 (O_2891,N_26073,N_28986);
nand UO_2892 (O_2892,N_24254,N_28589);
or UO_2893 (O_2893,N_29107,N_25209);
nand UO_2894 (O_2894,N_24221,N_28230);
and UO_2895 (O_2895,N_24232,N_26475);
nor UO_2896 (O_2896,N_26631,N_26936);
and UO_2897 (O_2897,N_24525,N_25336);
xnor UO_2898 (O_2898,N_24661,N_24017);
xnor UO_2899 (O_2899,N_26500,N_25733);
or UO_2900 (O_2900,N_27589,N_24033);
nand UO_2901 (O_2901,N_24160,N_24384);
or UO_2902 (O_2902,N_24162,N_28409);
nand UO_2903 (O_2903,N_29162,N_27542);
nor UO_2904 (O_2904,N_27179,N_26078);
or UO_2905 (O_2905,N_29809,N_29411);
nor UO_2906 (O_2906,N_24503,N_26833);
or UO_2907 (O_2907,N_25965,N_29810);
and UO_2908 (O_2908,N_29826,N_28919);
or UO_2909 (O_2909,N_25202,N_24964);
and UO_2910 (O_2910,N_28145,N_29548);
or UO_2911 (O_2911,N_28905,N_26252);
or UO_2912 (O_2912,N_29978,N_29222);
and UO_2913 (O_2913,N_25809,N_26958);
or UO_2914 (O_2914,N_28661,N_24312);
and UO_2915 (O_2915,N_28096,N_29352);
nor UO_2916 (O_2916,N_28757,N_28846);
nor UO_2917 (O_2917,N_24018,N_25437);
nand UO_2918 (O_2918,N_28860,N_24897);
nand UO_2919 (O_2919,N_29822,N_26592);
and UO_2920 (O_2920,N_29129,N_28584);
xnor UO_2921 (O_2921,N_28001,N_27554);
and UO_2922 (O_2922,N_28401,N_25582);
xor UO_2923 (O_2923,N_24239,N_28963);
xor UO_2924 (O_2924,N_29813,N_25200);
nand UO_2925 (O_2925,N_26973,N_26497);
nand UO_2926 (O_2926,N_25956,N_26403);
or UO_2927 (O_2927,N_26998,N_28942);
and UO_2928 (O_2928,N_28780,N_25270);
or UO_2929 (O_2929,N_29442,N_24812);
or UO_2930 (O_2930,N_28545,N_24161);
or UO_2931 (O_2931,N_27880,N_29081);
xor UO_2932 (O_2932,N_26636,N_29459);
nand UO_2933 (O_2933,N_29046,N_24106);
and UO_2934 (O_2934,N_29093,N_29480);
nand UO_2935 (O_2935,N_24324,N_26333);
or UO_2936 (O_2936,N_24037,N_28969);
or UO_2937 (O_2937,N_25695,N_29465);
and UO_2938 (O_2938,N_27506,N_29982);
nor UO_2939 (O_2939,N_28476,N_24594);
and UO_2940 (O_2940,N_24634,N_25641);
or UO_2941 (O_2941,N_28999,N_24150);
or UO_2942 (O_2942,N_29610,N_27556);
or UO_2943 (O_2943,N_27976,N_27623);
or UO_2944 (O_2944,N_24114,N_26541);
and UO_2945 (O_2945,N_27624,N_28613);
or UO_2946 (O_2946,N_24110,N_25083);
and UO_2947 (O_2947,N_25198,N_24213);
or UO_2948 (O_2948,N_26605,N_24425);
and UO_2949 (O_2949,N_25858,N_27892);
nor UO_2950 (O_2950,N_29212,N_27646);
or UO_2951 (O_2951,N_27806,N_29796);
nor UO_2952 (O_2952,N_27230,N_28677);
or UO_2953 (O_2953,N_26271,N_29928);
or UO_2954 (O_2954,N_26051,N_26837);
or UO_2955 (O_2955,N_26829,N_24455);
or UO_2956 (O_2956,N_25550,N_24512);
and UO_2957 (O_2957,N_24574,N_28065);
nor UO_2958 (O_2958,N_29291,N_26210);
nand UO_2959 (O_2959,N_25049,N_26218);
nor UO_2960 (O_2960,N_26405,N_28850);
nor UO_2961 (O_2961,N_29412,N_25917);
nor UO_2962 (O_2962,N_26662,N_25635);
nor UO_2963 (O_2963,N_24327,N_28207);
xnor UO_2964 (O_2964,N_27812,N_28737);
nor UO_2965 (O_2965,N_26484,N_26297);
nand UO_2966 (O_2966,N_28341,N_28636);
and UO_2967 (O_2967,N_29644,N_26784);
nand UO_2968 (O_2968,N_25335,N_29763);
nor UO_2969 (O_2969,N_24814,N_27628);
and UO_2970 (O_2970,N_25578,N_25244);
nand UO_2971 (O_2971,N_29931,N_26482);
xnor UO_2972 (O_2972,N_28006,N_24379);
and UO_2973 (O_2973,N_27567,N_27209);
and UO_2974 (O_2974,N_25562,N_29384);
xnor UO_2975 (O_2975,N_27603,N_26772);
nor UO_2976 (O_2976,N_26466,N_26983);
nand UO_2977 (O_2977,N_25532,N_25824);
or UO_2978 (O_2978,N_26054,N_27113);
nor UO_2979 (O_2979,N_29900,N_26065);
nor UO_2980 (O_2980,N_27194,N_26977);
nor UO_2981 (O_2981,N_24087,N_27112);
nor UO_2982 (O_2982,N_27804,N_29263);
nand UO_2983 (O_2983,N_27469,N_24901);
or UO_2984 (O_2984,N_29221,N_26518);
or UO_2985 (O_2985,N_28836,N_27168);
and UO_2986 (O_2986,N_24858,N_29704);
nand UO_2987 (O_2987,N_29923,N_29029);
or UO_2988 (O_2988,N_26128,N_28067);
nand UO_2989 (O_2989,N_27677,N_28064);
nor UO_2990 (O_2990,N_24987,N_28394);
or UO_2991 (O_2991,N_24074,N_24859);
xnor UO_2992 (O_2992,N_25863,N_24592);
xnor UO_2993 (O_2993,N_25759,N_27048);
and UO_2994 (O_2994,N_24688,N_27298);
and UO_2995 (O_2995,N_29008,N_26311);
nand UO_2996 (O_2996,N_26274,N_26771);
nor UO_2997 (O_2997,N_24776,N_26007);
nand UO_2998 (O_2998,N_27281,N_26971);
or UO_2999 (O_2999,N_26273,N_28721);
nand UO_3000 (O_3000,N_25422,N_24886);
nand UO_3001 (O_3001,N_26872,N_25789);
nand UO_3002 (O_3002,N_28233,N_29322);
nor UO_3003 (O_3003,N_24033,N_28984);
or UO_3004 (O_3004,N_26428,N_28322);
nor UO_3005 (O_3005,N_25188,N_27570);
and UO_3006 (O_3006,N_26376,N_27373);
or UO_3007 (O_3007,N_26661,N_24051);
and UO_3008 (O_3008,N_27075,N_27230);
or UO_3009 (O_3009,N_26888,N_27830);
or UO_3010 (O_3010,N_25607,N_28251);
xor UO_3011 (O_3011,N_28007,N_28939);
and UO_3012 (O_3012,N_25605,N_29424);
nor UO_3013 (O_3013,N_29170,N_27976);
nor UO_3014 (O_3014,N_24899,N_25506);
nand UO_3015 (O_3015,N_24422,N_29829);
xnor UO_3016 (O_3016,N_24167,N_24859);
nand UO_3017 (O_3017,N_26409,N_29111);
and UO_3018 (O_3018,N_24043,N_27320);
and UO_3019 (O_3019,N_25759,N_27040);
and UO_3020 (O_3020,N_28852,N_28046);
and UO_3021 (O_3021,N_29300,N_24533);
nand UO_3022 (O_3022,N_29843,N_29315);
nor UO_3023 (O_3023,N_27226,N_25911);
nand UO_3024 (O_3024,N_25174,N_28910);
or UO_3025 (O_3025,N_26306,N_26986);
nand UO_3026 (O_3026,N_25444,N_29165);
nor UO_3027 (O_3027,N_26992,N_29160);
nor UO_3028 (O_3028,N_27597,N_26427);
nand UO_3029 (O_3029,N_26085,N_28877);
nor UO_3030 (O_3030,N_25204,N_25818);
and UO_3031 (O_3031,N_28081,N_29958);
nand UO_3032 (O_3032,N_28852,N_29296);
nand UO_3033 (O_3033,N_24373,N_28913);
nand UO_3034 (O_3034,N_29584,N_29066);
nand UO_3035 (O_3035,N_27472,N_29982);
xnor UO_3036 (O_3036,N_27264,N_24195);
nand UO_3037 (O_3037,N_25107,N_24500);
and UO_3038 (O_3038,N_25965,N_25460);
or UO_3039 (O_3039,N_25586,N_28822);
nor UO_3040 (O_3040,N_25257,N_28229);
and UO_3041 (O_3041,N_28937,N_24003);
and UO_3042 (O_3042,N_25408,N_29868);
or UO_3043 (O_3043,N_25732,N_28999);
or UO_3044 (O_3044,N_24005,N_26372);
or UO_3045 (O_3045,N_24404,N_25204);
nand UO_3046 (O_3046,N_28768,N_28388);
or UO_3047 (O_3047,N_26694,N_27809);
xor UO_3048 (O_3048,N_29134,N_24937);
nand UO_3049 (O_3049,N_28822,N_28978);
or UO_3050 (O_3050,N_26867,N_25094);
nand UO_3051 (O_3051,N_28486,N_26728);
and UO_3052 (O_3052,N_26499,N_24307);
or UO_3053 (O_3053,N_28132,N_26139);
nand UO_3054 (O_3054,N_25241,N_28178);
or UO_3055 (O_3055,N_26088,N_29331);
and UO_3056 (O_3056,N_28846,N_24793);
nor UO_3057 (O_3057,N_26712,N_24479);
xnor UO_3058 (O_3058,N_26563,N_29959);
and UO_3059 (O_3059,N_25420,N_29361);
and UO_3060 (O_3060,N_29970,N_29829);
nand UO_3061 (O_3061,N_25313,N_24547);
nand UO_3062 (O_3062,N_26891,N_27621);
and UO_3063 (O_3063,N_26487,N_24423);
and UO_3064 (O_3064,N_28813,N_29906);
and UO_3065 (O_3065,N_24532,N_27781);
or UO_3066 (O_3066,N_24197,N_26223);
nor UO_3067 (O_3067,N_25659,N_24104);
or UO_3068 (O_3068,N_29737,N_28511);
nand UO_3069 (O_3069,N_28628,N_27150);
or UO_3070 (O_3070,N_27571,N_29440);
or UO_3071 (O_3071,N_27421,N_26588);
xnor UO_3072 (O_3072,N_27050,N_28742);
and UO_3073 (O_3073,N_25144,N_29494);
or UO_3074 (O_3074,N_25512,N_25558);
nor UO_3075 (O_3075,N_25746,N_26950);
and UO_3076 (O_3076,N_26174,N_29400);
and UO_3077 (O_3077,N_27929,N_27491);
or UO_3078 (O_3078,N_25198,N_29133);
nor UO_3079 (O_3079,N_26892,N_24202);
xnor UO_3080 (O_3080,N_24271,N_29818);
or UO_3081 (O_3081,N_27658,N_28878);
nor UO_3082 (O_3082,N_28790,N_24442);
nand UO_3083 (O_3083,N_24529,N_28257);
nor UO_3084 (O_3084,N_27079,N_25715);
nor UO_3085 (O_3085,N_29087,N_29816);
and UO_3086 (O_3086,N_26780,N_26608);
or UO_3087 (O_3087,N_27811,N_27695);
or UO_3088 (O_3088,N_26873,N_24233);
nand UO_3089 (O_3089,N_25710,N_26093);
nor UO_3090 (O_3090,N_24556,N_29877);
nor UO_3091 (O_3091,N_27387,N_24616);
nor UO_3092 (O_3092,N_28803,N_27856);
nor UO_3093 (O_3093,N_24394,N_25443);
and UO_3094 (O_3094,N_26695,N_25551);
nor UO_3095 (O_3095,N_29202,N_24302);
and UO_3096 (O_3096,N_26654,N_24328);
or UO_3097 (O_3097,N_29300,N_25205);
and UO_3098 (O_3098,N_26761,N_25188);
and UO_3099 (O_3099,N_25708,N_24873);
nor UO_3100 (O_3100,N_26564,N_27464);
xor UO_3101 (O_3101,N_25318,N_29368);
or UO_3102 (O_3102,N_27993,N_26669);
nor UO_3103 (O_3103,N_25220,N_25941);
or UO_3104 (O_3104,N_28699,N_29106);
or UO_3105 (O_3105,N_28574,N_24169);
and UO_3106 (O_3106,N_25459,N_29564);
or UO_3107 (O_3107,N_27205,N_26325);
or UO_3108 (O_3108,N_28852,N_28461);
xnor UO_3109 (O_3109,N_29504,N_29105);
nand UO_3110 (O_3110,N_28191,N_24703);
nor UO_3111 (O_3111,N_24466,N_27605);
nand UO_3112 (O_3112,N_26747,N_26924);
or UO_3113 (O_3113,N_24465,N_24621);
nand UO_3114 (O_3114,N_26881,N_28545);
nor UO_3115 (O_3115,N_25098,N_24909);
or UO_3116 (O_3116,N_25099,N_28109);
and UO_3117 (O_3117,N_28499,N_28617);
xnor UO_3118 (O_3118,N_28141,N_27324);
or UO_3119 (O_3119,N_29336,N_26862);
nor UO_3120 (O_3120,N_26013,N_29678);
or UO_3121 (O_3121,N_28460,N_24596);
nand UO_3122 (O_3122,N_28879,N_28100);
and UO_3123 (O_3123,N_24883,N_29946);
nor UO_3124 (O_3124,N_28135,N_28170);
and UO_3125 (O_3125,N_28838,N_28706);
nor UO_3126 (O_3126,N_26056,N_25269);
nand UO_3127 (O_3127,N_29502,N_27395);
nor UO_3128 (O_3128,N_24049,N_29804);
or UO_3129 (O_3129,N_29144,N_25390);
and UO_3130 (O_3130,N_29720,N_24342);
nor UO_3131 (O_3131,N_29966,N_28811);
and UO_3132 (O_3132,N_27711,N_25195);
nor UO_3133 (O_3133,N_24181,N_28007);
or UO_3134 (O_3134,N_24175,N_25141);
or UO_3135 (O_3135,N_29255,N_24249);
nand UO_3136 (O_3136,N_29001,N_24753);
and UO_3137 (O_3137,N_25557,N_28765);
nand UO_3138 (O_3138,N_24966,N_27035);
and UO_3139 (O_3139,N_24399,N_26742);
nor UO_3140 (O_3140,N_29918,N_27011);
nor UO_3141 (O_3141,N_29003,N_27538);
nand UO_3142 (O_3142,N_27821,N_28299);
nand UO_3143 (O_3143,N_28969,N_27368);
nor UO_3144 (O_3144,N_26740,N_28602);
and UO_3145 (O_3145,N_26242,N_24468);
nand UO_3146 (O_3146,N_29782,N_27043);
or UO_3147 (O_3147,N_24363,N_24525);
or UO_3148 (O_3148,N_28167,N_26005);
or UO_3149 (O_3149,N_26590,N_24689);
or UO_3150 (O_3150,N_29481,N_29523);
nor UO_3151 (O_3151,N_24927,N_29131);
and UO_3152 (O_3152,N_25684,N_25064);
nor UO_3153 (O_3153,N_28343,N_29150);
and UO_3154 (O_3154,N_26158,N_29854);
and UO_3155 (O_3155,N_29524,N_26675);
and UO_3156 (O_3156,N_28192,N_26647);
and UO_3157 (O_3157,N_26146,N_26335);
xor UO_3158 (O_3158,N_25395,N_27216);
or UO_3159 (O_3159,N_27599,N_29028);
and UO_3160 (O_3160,N_26401,N_29387);
and UO_3161 (O_3161,N_27160,N_28328);
or UO_3162 (O_3162,N_28049,N_28034);
nor UO_3163 (O_3163,N_26895,N_26828);
nor UO_3164 (O_3164,N_27031,N_27058);
and UO_3165 (O_3165,N_27132,N_24372);
xor UO_3166 (O_3166,N_24797,N_27351);
nand UO_3167 (O_3167,N_28623,N_27627);
or UO_3168 (O_3168,N_29244,N_25780);
or UO_3169 (O_3169,N_28898,N_24213);
xor UO_3170 (O_3170,N_28842,N_24222);
nor UO_3171 (O_3171,N_24105,N_27244);
or UO_3172 (O_3172,N_26556,N_26878);
or UO_3173 (O_3173,N_26069,N_28522);
nand UO_3174 (O_3174,N_25608,N_24313);
nand UO_3175 (O_3175,N_27581,N_25860);
and UO_3176 (O_3176,N_26947,N_27419);
nand UO_3177 (O_3177,N_27236,N_24024);
nand UO_3178 (O_3178,N_27806,N_26363);
or UO_3179 (O_3179,N_29565,N_26348);
and UO_3180 (O_3180,N_24143,N_26814);
or UO_3181 (O_3181,N_25633,N_27809);
nand UO_3182 (O_3182,N_29561,N_27240);
nand UO_3183 (O_3183,N_27505,N_28324);
and UO_3184 (O_3184,N_26404,N_25993);
nand UO_3185 (O_3185,N_24563,N_26988);
nor UO_3186 (O_3186,N_25318,N_24867);
nand UO_3187 (O_3187,N_27049,N_28338);
xnor UO_3188 (O_3188,N_29050,N_27106);
and UO_3189 (O_3189,N_25544,N_28555);
and UO_3190 (O_3190,N_27175,N_28841);
or UO_3191 (O_3191,N_29595,N_26165);
nand UO_3192 (O_3192,N_29612,N_28333);
or UO_3193 (O_3193,N_24883,N_28600);
nand UO_3194 (O_3194,N_27948,N_25006);
and UO_3195 (O_3195,N_26538,N_26939);
and UO_3196 (O_3196,N_24559,N_24849);
xnor UO_3197 (O_3197,N_27846,N_24124);
and UO_3198 (O_3198,N_27163,N_28753);
or UO_3199 (O_3199,N_25695,N_27911);
nor UO_3200 (O_3200,N_25060,N_25279);
nand UO_3201 (O_3201,N_27263,N_24387);
or UO_3202 (O_3202,N_27074,N_27493);
nor UO_3203 (O_3203,N_25130,N_25466);
or UO_3204 (O_3204,N_29816,N_24224);
nand UO_3205 (O_3205,N_29392,N_27497);
or UO_3206 (O_3206,N_27926,N_26931);
and UO_3207 (O_3207,N_24910,N_24652);
or UO_3208 (O_3208,N_29678,N_28667);
or UO_3209 (O_3209,N_27449,N_28018);
xnor UO_3210 (O_3210,N_26781,N_27443);
and UO_3211 (O_3211,N_28203,N_25960);
and UO_3212 (O_3212,N_27914,N_25378);
nand UO_3213 (O_3213,N_24835,N_24295);
nor UO_3214 (O_3214,N_25102,N_26322);
or UO_3215 (O_3215,N_27092,N_25681);
nand UO_3216 (O_3216,N_25586,N_29190);
and UO_3217 (O_3217,N_25637,N_24036);
nor UO_3218 (O_3218,N_24309,N_25071);
and UO_3219 (O_3219,N_27338,N_26643);
or UO_3220 (O_3220,N_26595,N_24837);
nor UO_3221 (O_3221,N_25807,N_24542);
and UO_3222 (O_3222,N_25376,N_29153);
or UO_3223 (O_3223,N_25862,N_29751);
or UO_3224 (O_3224,N_27643,N_28819);
and UO_3225 (O_3225,N_26833,N_26505);
nand UO_3226 (O_3226,N_27063,N_28082);
or UO_3227 (O_3227,N_26568,N_29266);
nor UO_3228 (O_3228,N_25458,N_27225);
nor UO_3229 (O_3229,N_25290,N_29441);
nand UO_3230 (O_3230,N_26269,N_25236);
nor UO_3231 (O_3231,N_27353,N_27356);
or UO_3232 (O_3232,N_29228,N_25511);
or UO_3233 (O_3233,N_26739,N_24072);
and UO_3234 (O_3234,N_26729,N_29971);
nand UO_3235 (O_3235,N_27113,N_28547);
or UO_3236 (O_3236,N_26830,N_27932);
xor UO_3237 (O_3237,N_27190,N_29363);
nor UO_3238 (O_3238,N_26951,N_26956);
nand UO_3239 (O_3239,N_27514,N_25133);
nor UO_3240 (O_3240,N_26236,N_26805);
xor UO_3241 (O_3241,N_28964,N_24760);
and UO_3242 (O_3242,N_25802,N_24589);
or UO_3243 (O_3243,N_28264,N_29459);
xor UO_3244 (O_3244,N_29846,N_29197);
or UO_3245 (O_3245,N_24578,N_29771);
or UO_3246 (O_3246,N_29528,N_29876);
or UO_3247 (O_3247,N_25174,N_26589);
or UO_3248 (O_3248,N_29766,N_28546);
and UO_3249 (O_3249,N_28479,N_25993);
or UO_3250 (O_3250,N_24704,N_29846);
nand UO_3251 (O_3251,N_25109,N_26467);
or UO_3252 (O_3252,N_24080,N_24192);
and UO_3253 (O_3253,N_24101,N_28059);
nand UO_3254 (O_3254,N_27003,N_25834);
or UO_3255 (O_3255,N_29704,N_27750);
and UO_3256 (O_3256,N_24336,N_26982);
or UO_3257 (O_3257,N_27539,N_26722);
nand UO_3258 (O_3258,N_25613,N_28377);
nand UO_3259 (O_3259,N_28108,N_28665);
nor UO_3260 (O_3260,N_25503,N_25104);
nand UO_3261 (O_3261,N_28576,N_25508);
or UO_3262 (O_3262,N_26229,N_29226);
nor UO_3263 (O_3263,N_25733,N_28260);
or UO_3264 (O_3264,N_28471,N_24727);
nand UO_3265 (O_3265,N_27895,N_28639);
nor UO_3266 (O_3266,N_29883,N_27336);
nor UO_3267 (O_3267,N_29275,N_25111);
and UO_3268 (O_3268,N_24117,N_28925);
xnor UO_3269 (O_3269,N_28084,N_28017);
nor UO_3270 (O_3270,N_27403,N_27555);
and UO_3271 (O_3271,N_27197,N_25551);
and UO_3272 (O_3272,N_27835,N_29940);
nand UO_3273 (O_3273,N_28499,N_28207);
or UO_3274 (O_3274,N_26864,N_29654);
and UO_3275 (O_3275,N_29952,N_27207);
nor UO_3276 (O_3276,N_26199,N_29660);
nand UO_3277 (O_3277,N_25557,N_26608);
and UO_3278 (O_3278,N_25948,N_27609);
nor UO_3279 (O_3279,N_24987,N_25831);
nand UO_3280 (O_3280,N_29605,N_24656);
nand UO_3281 (O_3281,N_24917,N_25212);
or UO_3282 (O_3282,N_28708,N_29536);
nor UO_3283 (O_3283,N_25875,N_29808);
or UO_3284 (O_3284,N_29254,N_27003);
and UO_3285 (O_3285,N_25274,N_28849);
and UO_3286 (O_3286,N_28378,N_27377);
nand UO_3287 (O_3287,N_24266,N_28892);
and UO_3288 (O_3288,N_28128,N_27528);
and UO_3289 (O_3289,N_26613,N_28458);
nand UO_3290 (O_3290,N_28042,N_24240);
nor UO_3291 (O_3291,N_24294,N_26278);
nor UO_3292 (O_3292,N_26427,N_28151);
and UO_3293 (O_3293,N_24420,N_25591);
and UO_3294 (O_3294,N_26519,N_27485);
nor UO_3295 (O_3295,N_26473,N_27046);
and UO_3296 (O_3296,N_28536,N_25363);
xnor UO_3297 (O_3297,N_28287,N_28260);
nand UO_3298 (O_3298,N_25290,N_24602);
and UO_3299 (O_3299,N_28183,N_25422);
nor UO_3300 (O_3300,N_28303,N_24436);
or UO_3301 (O_3301,N_26422,N_26785);
nor UO_3302 (O_3302,N_24031,N_28446);
nor UO_3303 (O_3303,N_24199,N_29056);
and UO_3304 (O_3304,N_25226,N_25758);
and UO_3305 (O_3305,N_29514,N_29862);
or UO_3306 (O_3306,N_28466,N_28034);
nor UO_3307 (O_3307,N_25907,N_28288);
or UO_3308 (O_3308,N_24491,N_25493);
nand UO_3309 (O_3309,N_28783,N_28026);
nor UO_3310 (O_3310,N_27670,N_27641);
and UO_3311 (O_3311,N_29369,N_25595);
nor UO_3312 (O_3312,N_27340,N_25540);
or UO_3313 (O_3313,N_29940,N_24829);
or UO_3314 (O_3314,N_29481,N_24826);
nor UO_3315 (O_3315,N_29853,N_26200);
xor UO_3316 (O_3316,N_24821,N_26031);
or UO_3317 (O_3317,N_27539,N_27345);
nand UO_3318 (O_3318,N_29411,N_29163);
or UO_3319 (O_3319,N_28273,N_29477);
nand UO_3320 (O_3320,N_28247,N_27182);
or UO_3321 (O_3321,N_27751,N_24481);
nand UO_3322 (O_3322,N_25096,N_24550);
or UO_3323 (O_3323,N_29539,N_29567);
and UO_3324 (O_3324,N_25950,N_27205);
nor UO_3325 (O_3325,N_24112,N_26144);
xor UO_3326 (O_3326,N_25636,N_29671);
xor UO_3327 (O_3327,N_26370,N_24734);
or UO_3328 (O_3328,N_27953,N_28122);
or UO_3329 (O_3329,N_25243,N_25971);
nand UO_3330 (O_3330,N_29925,N_25928);
or UO_3331 (O_3331,N_29620,N_29044);
nor UO_3332 (O_3332,N_26196,N_28312);
and UO_3333 (O_3333,N_24487,N_24095);
and UO_3334 (O_3334,N_28361,N_24590);
or UO_3335 (O_3335,N_26319,N_26098);
xnor UO_3336 (O_3336,N_27471,N_24612);
nor UO_3337 (O_3337,N_24858,N_29370);
nor UO_3338 (O_3338,N_24105,N_27238);
nor UO_3339 (O_3339,N_24214,N_29882);
and UO_3340 (O_3340,N_28008,N_24005);
nand UO_3341 (O_3341,N_27624,N_25107);
or UO_3342 (O_3342,N_24469,N_25687);
and UO_3343 (O_3343,N_29331,N_25225);
and UO_3344 (O_3344,N_24455,N_26383);
nor UO_3345 (O_3345,N_27237,N_24467);
and UO_3346 (O_3346,N_24821,N_25497);
and UO_3347 (O_3347,N_25823,N_25553);
xor UO_3348 (O_3348,N_25623,N_28714);
nand UO_3349 (O_3349,N_28261,N_24979);
nor UO_3350 (O_3350,N_24577,N_28048);
nand UO_3351 (O_3351,N_27498,N_24367);
nor UO_3352 (O_3352,N_25638,N_26405);
nand UO_3353 (O_3353,N_28599,N_26628);
nor UO_3354 (O_3354,N_26544,N_24991);
nand UO_3355 (O_3355,N_28149,N_29082);
or UO_3356 (O_3356,N_28603,N_24716);
xor UO_3357 (O_3357,N_24303,N_28986);
or UO_3358 (O_3358,N_26171,N_27812);
and UO_3359 (O_3359,N_25665,N_27571);
nand UO_3360 (O_3360,N_25241,N_28732);
and UO_3361 (O_3361,N_24068,N_29623);
and UO_3362 (O_3362,N_25273,N_27277);
xnor UO_3363 (O_3363,N_27745,N_29405);
xnor UO_3364 (O_3364,N_25574,N_29402);
nor UO_3365 (O_3365,N_24549,N_29676);
nand UO_3366 (O_3366,N_29239,N_25898);
nand UO_3367 (O_3367,N_28429,N_25326);
and UO_3368 (O_3368,N_24705,N_28117);
or UO_3369 (O_3369,N_26789,N_26077);
or UO_3370 (O_3370,N_26354,N_28848);
xor UO_3371 (O_3371,N_24097,N_27708);
nand UO_3372 (O_3372,N_26781,N_27120);
and UO_3373 (O_3373,N_26635,N_26887);
nand UO_3374 (O_3374,N_24443,N_24575);
xnor UO_3375 (O_3375,N_29163,N_29057);
and UO_3376 (O_3376,N_24214,N_25264);
nand UO_3377 (O_3377,N_24899,N_26924);
or UO_3378 (O_3378,N_29956,N_29314);
nor UO_3379 (O_3379,N_28521,N_25153);
nand UO_3380 (O_3380,N_26500,N_24129);
or UO_3381 (O_3381,N_25063,N_27531);
xor UO_3382 (O_3382,N_25382,N_27509);
xnor UO_3383 (O_3383,N_25912,N_24852);
and UO_3384 (O_3384,N_26501,N_24480);
and UO_3385 (O_3385,N_26120,N_27127);
nand UO_3386 (O_3386,N_26965,N_25529);
and UO_3387 (O_3387,N_28556,N_28675);
nand UO_3388 (O_3388,N_29016,N_25202);
xor UO_3389 (O_3389,N_29651,N_27495);
or UO_3390 (O_3390,N_28837,N_24080);
or UO_3391 (O_3391,N_25395,N_28671);
nand UO_3392 (O_3392,N_26100,N_27695);
nand UO_3393 (O_3393,N_28552,N_28635);
nor UO_3394 (O_3394,N_28055,N_27781);
or UO_3395 (O_3395,N_25517,N_29134);
and UO_3396 (O_3396,N_26074,N_24487);
nand UO_3397 (O_3397,N_27937,N_25037);
or UO_3398 (O_3398,N_25577,N_26101);
nand UO_3399 (O_3399,N_29647,N_28078);
or UO_3400 (O_3400,N_25331,N_27581);
and UO_3401 (O_3401,N_27290,N_24395);
xor UO_3402 (O_3402,N_24783,N_27765);
xor UO_3403 (O_3403,N_28375,N_27041);
and UO_3404 (O_3404,N_29881,N_24352);
nor UO_3405 (O_3405,N_28692,N_24943);
nand UO_3406 (O_3406,N_25187,N_27953);
and UO_3407 (O_3407,N_25354,N_29838);
and UO_3408 (O_3408,N_26888,N_25561);
nand UO_3409 (O_3409,N_26734,N_26135);
nand UO_3410 (O_3410,N_26197,N_29534);
or UO_3411 (O_3411,N_24707,N_26444);
or UO_3412 (O_3412,N_27249,N_29096);
nand UO_3413 (O_3413,N_29412,N_29609);
nand UO_3414 (O_3414,N_28740,N_27527);
or UO_3415 (O_3415,N_27068,N_25724);
nand UO_3416 (O_3416,N_29466,N_29646);
and UO_3417 (O_3417,N_26211,N_25168);
and UO_3418 (O_3418,N_28763,N_25114);
or UO_3419 (O_3419,N_24396,N_24563);
xnor UO_3420 (O_3420,N_28700,N_28998);
nor UO_3421 (O_3421,N_24874,N_29132);
xor UO_3422 (O_3422,N_29358,N_24016);
and UO_3423 (O_3423,N_28405,N_25746);
nor UO_3424 (O_3424,N_28416,N_24649);
nand UO_3425 (O_3425,N_26683,N_29450);
nor UO_3426 (O_3426,N_28351,N_29139);
nor UO_3427 (O_3427,N_24958,N_25334);
or UO_3428 (O_3428,N_24258,N_26691);
and UO_3429 (O_3429,N_24847,N_25038);
nor UO_3430 (O_3430,N_24391,N_29870);
and UO_3431 (O_3431,N_25971,N_29426);
nor UO_3432 (O_3432,N_27767,N_26588);
nand UO_3433 (O_3433,N_25316,N_28695);
or UO_3434 (O_3434,N_24060,N_28990);
or UO_3435 (O_3435,N_28038,N_28266);
nand UO_3436 (O_3436,N_25307,N_29816);
and UO_3437 (O_3437,N_24389,N_29664);
nand UO_3438 (O_3438,N_27566,N_27178);
or UO_3439 (O_3439,N_24975,N_27618);
nor UO_3440 (O_3440,N_25056,N_27717);
nand UO_3441 (O_3441,N_27722,N_27519);
nor UO_3442 (O_3442,N_26386,N_25620);
nor UO_3443 (O_3443,N_29428,N_25440);
nand UO_3444 (O_3444,N_29727,N_24249);
xnor UO_3445 (O_3445,N_27167,N_29691);
nor UO_3446 (O_3446,N_24648,N_24381);
nor UO_3447 (O_3447,N_27845,N_27572);
or UO_3448 (O_3448,N_26726,N_28125);
and UO_3449 (O_3449,N_25436,N_29517);
nor UO_3450 (O_3450,N_27606,N_25757);
and UO_3451 (O_3451,N_28376,N_25694);
or UO_3452 (O_3452,N_27197,N_28896);
nor UO_3453 (O_3453,N_24727,N_25164);
or UO_3454 (O_3454,N_27677,N_28347);
and UO_3455 (O_3455,N_25637,N_25728);
nor UO_3456 (O_3456,N_25615,N_24505);
and UO_3457 (O_3457,N_24536,N_27005);
and UO_3458 (O_3458,N_28383,N_27430);
nor UO_3459 (O_3459,N_27546,N_28802);
nand UO_3460 (O_3460,N_24798,N_28335);
xnor UO_3461 (O_3461,N_29188,N_27171);
or UO_3462 (O_3462,N_29535,N_29323);
nand UO_3463 (O_3463,N_28718,N_29666);
and UO_3464 (O_3464,N_26972,N_25284);
xnor UO_3465 (O_3465,N_25022,N_24613);
nand UO_3466 (O_3466,N_28953,N_29401);
or UO_3467 (O_3467,N_27470,N_27854);
and UO_3468 (O_3468,N_29832,N_25605);
or UO_3469 (O_3469,N_29544,N_26775);
and UO_3470 (O_3470,N_25038,N_24698);
nand UO_3471 (O_3471,N_29093,N_29365);
nand UO_3472 (O_3472,N_27937,N_28760);
nand UO_3473 (O_3473,N_28248,N_25576);
and UO_3474 (O_3474,N_28124,N_25718);
or UO_3475 (O_3475,N_24268,N_26053);
and UO_3476 (O_3476,N_25839,N_29711);
nand UO_3477 (O_3477,N_27514,N_27060);
nor UO_3478 (O_3478,N_29995,N_29438);
nor UO_3479 (O_3479,N_27270,N_29644);
nor UO_3480 (O_3480,N_29126,N_28911);
and UO_3481 (O_3481,N_28143,N_28916);
nor UO_3482 (O_3482,N_29127,N_26081);
nand UO_3483 (O_3483,N_26829,N_28274);
and UO_3484 (O_3484,N_28759,N_25679);
nor UO_3485 (O_3485,N_26117,N_28322);
and UO_3486 (O_3486,N_27488,N_26057);
nor UO_3487 (O_3487,N_27536,N_27585);
nand UO_3488 (O_3488,N_25834,N_26164);
xor UO_3489 (O_3489,N_27017,N_26225);
or UO_3490 (O_3490,N_28461,N_26962);
or UO_3491 (O_3491,N_24189,N_25197);
nand UO_3492 (O_3492,N_29083,N_24677);
nor UO_3493 (O_3493,N_26982,N_29918);
or UO_3494 (O_3494,N_27714,N_29216);
xnor UO_3495 (O_3495,N_25808,N_24448);
nand UO_3496 (O_3496,N_29501,N_24635);
and UO_3497 (O_3497,N_24376,N_27617);
or UO_3498 (O_3498,N_24334,N_24738);
or UO_3499 (O_3499,N_25042,N_25811);
endmodule