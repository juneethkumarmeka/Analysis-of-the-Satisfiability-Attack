module basic_750_5000_1000_2_levels_1xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2511,N_2513,N_2514,N_2515,N_2517,N_2519,N_2520,N_2521,N_2522,N_2524,N_2525,N_2526,N_2527,N_2529,N_2530,N_2531,N_2532,N_2533,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2545,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2569,N_2570,N_2572,N_2573,N_2574,N_2575,N_2577,N_2578,N_2579,N_2581,N_2582,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2612,N_2613,N_2614,N_2615,N_2616,N_2620,N_2621,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2643,N_2645,N_2648,N_2649,N_2650,N_2651,N_2653,N_2654,N_2655,N_2656,N_2659,N_2660,N_2662,N_2664,N_2665,N_2666,N_2667,N_2670,N_2672,N_2673,N_2674,N_2675,N_2678,N_2680,N_2681,N_2682,N_2683,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2692,N_2693,N_2694,N_2695,N_2697,N_2698,N_2699,N_2700,N_2701,N_2703,N_2704,N_2705,N_2706,N_2707,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2748,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2766,N_2768,N_2770,N_2771,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2788,N_2789,N_2790,N_2791,N_2792,N_2794,N_2795,N_2796,N_2797,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2841,N_2842,N_2843,N_2845,N_2846,N_2848,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2862,N_2863,N_2864,N_2866,N_2867,N_2868,N_2869,N_2871,N_2872,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2882,N_2883,N_2884,N_2885,N_2887,N_2888,N_2889,N_2891,N_2892,N_2893,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2904,N_2906,N_2908,N_2910,N_2911,N_2912,N_2913,N_2915,N_2916,N_2917,N_2919,N_2920,N_2921,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2931,N_2932,N_2933,N_2935,N_2936,N_2939,N_2940,N_2941,N_2944,N_2945,N_2946,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2960,N_2961,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2974,N_2975,N_2977,N_2978,N_2979,N_2980,N_2981,N_2983,N_2984,N_2985,N_2987,N_2988,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3006,N_3008,N_3009,N_3010,N_3011,N_3014,N_3015,N_3016,N_3017,N_3018,N_3020,N_3021,N_3022,N_3023,N_3024,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3043,N_3044,N_3045,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3066,N_3067,N_3068,N_3069,N_3071,N_3072,N_3074,N_3076,N_3077,N_3078,N_3079,N_3080,N_3082,N_3083,N_3085,N_3087,N_3088,N_3089,N_3091,N_3093,N_3094,N_3095,N_3096,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3105,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3124,N_3125,N_3126,N_3127,N_3128,N_3131,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3142,N_3143,N_3144,N_3146,N_3148,N_3149,N_3150,N_3151,N_3152,N_3154,N_3155,N_3157,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3196,N_3197,N_3198,N_3199,N_3201,N_3202,N_3203,N_3205,N_3206,N_3208,N_3209,N_3212,N_3213,N_3214,N_3215,N_3216,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3225,N_3226,N_3227,N_3228,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3255,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3292,N_3293,N_3294,N_3295,N_3298,N_3299,N_3301,N_3302,N_3303,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3324,N_3325,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3337,N_3339,N_3340,N_3341,N_3342,N_3347,N_3348,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3360,N_3361,N_3362,N_3363,N_3364,N_3366,N_3367,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3386,N_3387,N_3388,N_3389,N_3390,N_3393,N_3395,N_3398,N_3399,N_3400,N_3401,N_3405,N_3406,N_3407,N_3408,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3448,N_3449,N_3450,N_3451,N_3452,N_3454,N_3455,N_3457,N_3458,N_3460,N_3463,N_3464,N_3465,N_3466,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3481,N_3482,N_3485,N_3486,N_3487,N_3489,N_3490,N_3491,N_3493,N_3494,N_3495,N_3497,N_3498,N_3499,N_3500,N_3501,N_3503,N_3504,N_3505,N_3506,N_3507,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3541,N_3542,N_3545,N_3546,N_3547,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3569,N_3573,N_3576,N_3577,N_3578,N_3580,N_3582,N_3583,N_3586,N_3587,N_3588,N_3589,N_3590,N_3592,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3603,N_3605,N_3606,N_3607,N_3608,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3617,N_3618,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3629,N_3630,N_3631,N_3634,N_3635,N_3636,N_3639,N_3640,N_3641,N_3644,N_3645,N_3646,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3658,N_3659,N_3661,N_3662,N_3663,N_3665,N_3666,N_3667,N_3669,N_3670,N_3673,N_3674,N_3675,N_3676,N_3678,N_3679,N_3680,N_3682,N_3683,N_3684,N_3685,N_3686,N_3688,N_3689,N_3690,N_3691,N_3692,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3709,N_3710,N_3711,N_3712,N_3713,N_3715,N_3717,N_3718,N_3719,N_3720,N_3721,N_3723,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3742,N_3744,N_3745,N_3746,N_3747,N_3748,N_3750,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3767,N_3769,N_3770,N_3772,N_3773,N_3775,N_3776,N_3778,N_3779,N_3780,N_3781,N_3783,N_3785,N_3786,N_3789,N_3790,N_3791,N_3792,N_3794,N_3795,N_3796,N_3797,N_3799,N_3800,N_3801,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3845,N_3846,N_3847,N_3848,N_3850,N_3851,N_3852,N_3853,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3875,N_3876,N_3878,N_3879,N_3880,N_3881,N_3882,N_3884,N_3885,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3905,N_3906,N_3907,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3925,N_3928,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3940,N_3942,N_3943,N_3947,N_3949,N_3950,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3960,N_3962,N_3963,N_3965,N_3966,N_3968,N_3969,N_3970,N_3971,N_3973,N_3974,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3985,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4007,N_4009,N_4010,N_4011,N_4012,N_4014,N_4016,N_4017,N_4018,N_4019,N_4020,N_4022,N_4024,N_4025,N_4026,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4039,N_4040,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4055,N_4056,N_4058,N_4059,N_4060,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4083,N_4084,N_4085,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4094,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4103,N_4104,N_4105,N_4106,N_4107,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4120,N_4122,N_4124,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4137,N_4138,N_4140,N_4141,N_4143,N_4145,N_4146,N_4148,N_4149,N_4150,N_4151,N_4153,N_4154,N_4155,N_4156,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4167,N_4168,N_4170,N_4171,N_4173,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4187,N_4188,N_4190,N_4191,N_4192,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4214,N_4215,N_4216,N_4217,N_4218,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4251,N_4252,N_4253,N_4254,N_4256,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4287,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4301,N_4302,N_4303,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4314,N_4317,N_4318,N_4319,N_4320,N_4322,N_4323,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4356,N_4357,N_4359,N_4360,N_4361,N_4362,N_4364,N_4365,N_4367,N_4368,N_4369,N_4371,N_4372,N_4373,N_4374,N_4375,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4385,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4400,N_4401,N_4402,N_4403,N_4405,N_4406,N_4407,N_4408,N_4409,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4425,N_4426,N_4427,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4443,N_4444,N_4445,N_4446,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4458,N_4459,N_4460,N_4461,N_4462,N_4464,N_4466,N_4467,N_4468,N_4472,N_4474,N_4475,N_4476,N_4478,N_4479,N_4480,N_4481,N_4483,N_4484,N_4485,N_4489,N_4491,N_4492,N_4493,N_4494,N_4495,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4507,N_4508,N_4509,N_4512,N_4513,N_4515,N_4516,N_4519,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4536,N_4537,N_4538,N_4540,N_4541,N_4544,N_4545,N_4546,N_4547,N_4549,N_4550,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4566,N_4567,N_4568,N_4570,N_4572,N_4574,N_4575,N_4576,N_4577,N_4578,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4588,N_4590,N_4592,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4602,N_4603,N_4605,N_4606,N_4607,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4620,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4650,N_4651,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4660,N_4661,N_4663,N_4664,N_4665,N_4666,N_4668,N_4669,N_4670,N_4671,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4681,N_4682,N_4683,N_4685,N_4686,N_4688,N_4690,N_4692,N_4693,N_4694,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4717,N_4718,N_4720,N_4721,N_4724,N_4726,N_4728,N_4729,N_4730,N_4731,N_4733,N_4734,N_4736,N_4737,N_4738,N_4739,N_4740,N_4742,N_4744,N_4746,N_4747,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4756,N_4757,N_4759,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4788,N_4789,N_4790,N_4791,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4801,N_4804,N_4805,N_4806,N_4807,N_4808,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4821,N_4822,N_4824,N_4826,N_4827,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4841,N_4842,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4851,N_4852,N_4853,N_4855,N_4856,N_4857,N_4858,N_4860,N_4863,N_4864,N_4865,N_4866,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4883,N_4884,N_4886,N_4888,N_4889,N_4890,N_4891,N_4893,N_4894,N_4895,N_4897,N_4898,N_4899,N_4900,N_4901,N_4903,N_4904,N_4906,N_4907,N_4910,N_4911,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4922,N_4924,N_4925,N_4926,N_4927,N_4928,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4988,N_4991,N_4995,N_4997,N_4998,N_4999;
nand U0 (N_0,In_418,In_227);
and U1 (N_1,In_16,In_595);
or U2 (N_2,In_170,In_317);
nor U3 (N_3,In_698,In_38);
nor U4 (N_4,In_279,In_191);
or U5 (N_5,In_402,In_129);
nand U6 (N_6,In_510,In_79);
or U7 (N_7,In_328,In_161);
and U8 (N_8,In_245,In_122);
or U9 (N_9,In_333,In_326);
nor U10 (N_10,In_253,In_638);
nand U11 (N_11,In_549,In_186);
nand U12 (N_12,In_351,In_662);
or U13 (N_13,In_426,In_81);
nand U14 (N_14,In_578,In_360);
nor U15 (N_15,In_98,In_142);
nor U16 (N_16,In_444,In_18);
or U17 (N_17,In_659,In_195);
nor U18 (N_18,In_221,In_41);
nor U19 (N_19,In_667,In_190);
and U20 (N_20,In_302,In_180);
or U21 (N_21,In_384,In_475);
nor U22 (N_22,In_162,In_622);
nor U23 (N_23,In_387,In_263);
or U24 (N_24,In_434,In_584);
or U25 (N_25,In_17,In_347);
nor U26 (N_26,In_681,In_348);
xor U27 (N_27,In_218,In_108);
and U28 (N_28,In_518,In_0);
and U29 (N_29,In_59,In_255);
and U30 (N_30,In_741,In_281);
nor U31 (N_31,In_72,In_600);
and U32 (N_32,In_345,In_690);
nand U33 (N_33,In_587,In_254);
nor U34 (N_34,In_494,In_504);
nor U35 (N_35,In_153,In_496);
or U36 (N_36,In_528,In_313);
and U37 (N_37,In_67,In_433);
nor U38 (N_38,In_643,In_749);
or U39 (N_39,In_216,In_175);
nor U40 (N_40,In_316,In_231);
nand U41 (N_41,In_329,In_113);
and U42 (N_42,In_439,In_624);
nor U43 (N_43,In_453,In_267);
nor U44 (N_44,In_93,In_53);
and U45 (N_45,In_295,In_286);
nand U46 (N_46,In_337,In_451);
nand U47 (N_47,In_620,In_582);
or U48 (N_48,In_469,In_487);
nand U49 (N_49,In_722,In_382);
and U50 (N_50,In_45,In_590);
nor U51 (N_51,In_48,In_725);
nand U52 (N_52,In_399,In_557);
and U53 (N_53,In_711,In_696);
xnor U54 (N_54,In_233,In_131);
nand U55 (N_55,In_378,In_686);
nand U56 (N_56,In_523,In_211);
and U57 (N_57,In_520,In_393);
or U58 (N_58,In_85,In_394);
or U59 (N_59,In_219,In_648);
and U60 (N_60,In_572,In_693);
nand U61 (N_61,In_728,In_168);
or U62 (N_62,In_82,In_630);
nand U63 (N_63,In_558,In_71);
and U64 (N_64,In_178,In_63);
and U65 (N_65,In_465,In_127);
nor U66 (N_66,In_410,In_181);
or U67 (N_67,In_604,In_565);
or U68 (N_68,In_193,In_401);
nand U69 (N_69,In_720,In_466);
or U70 (N_70,In_117,In_336);
or U71 (N_71,In_99,In_357);
nor U72 (N_72,In_602,In_265);
or U73 (N_73,In_610,In_513);
nand U74 (N_74,In_42,In_737);
nor U75 (N_75,In_629,In_704);
or U76 (N_76,In_516,In_432);
nor U77 (N_77,In_14,In_101);
nor U78 (N_78,In_311,In_152);
and U79 (N_79,In_588,In_207);
or U80 (N_80,In_301,In_293);
nor U81 (N_81,In_519,In_413);
nor U82 (N_82,In_577,In_96);
and U83 (N_83,In_146,In_362);
nor U84 (N_84,In_47,In_442);
and U85 (N_85,In_187,In_546);
nand U86 (N_86,In_566,In_223);
nor U87 (N_87,In_296,In_213);
nand U88 (N_88,In_372,In_273);
and U89 (N_89,In_331,In_228);
nand U90 (N_90,In_585,In_349);
and U91 (N_91,In_11,In_60);
nor U92 (N_92,In_226,In_3);
nand U93 (N_93,In_116,In_506);
nor U94 (N_94,In_593,In_389);
xnor U95 (N_95,In_613,In_661);
and U96 (N_96,In_441,In_208);
nand U97 (N_97,In_135,In_94);
or U98 (N_98,In_555,In_647);
or U99 (N_99,In_673,In_31);
nor U100 (N_100,In_144,In_561);
nor U101 (N_101,In_498,In_283);
or U102 (N_102,In_395,In_609);
nor U103 (N_103,In_714,In_700);
and U104 (N_104,In_318,In_633);
and U105 (N_105,In_635,In_199);
nand U106 (N_106,In_710,In_30);
or U107 (N_107,In_49,In_644);
nor U108 (N_108,In_458,In_437);
nor U109 (N_109,In_392,In_627);
or U110 (N_110,In_192,In_503);
or U111 (N_111,In_292,In_145);
or U112 (N_112,In_352,In_545);
nor U113 (N_113,In_478,In_482);
nor U114 (N_114,In_535,In_87);
or U115 (N_115,In_637,In_525);
and U116 (N_116,In_636,In_137);
and U117 (N_117,In_297,In_385);
nor U118 (N_118,In_745,In_205);
and U119 (N_119,In_568,In_452);
or U120 (N_120,In_134,In_438);
and U121 (N_121,In_576,In_65);
and U122 (N_122,In_697,In_685);
and U123 (N_123,In_88,In_386);
nand U124 (N_124,In_90,In_376);
nand U125 (N_125,In_684,In_550);
nand U126 (N_126,In_455,In_705);
nand U127 (N_127,In_78,In_111);
nand U128 (N_128,In_562,In_107);
or U129 (N_129,In_381,In_414);
or U130 (N_130,In_32,In_702);
or U131 (N_131,In_532,In_20);
nand U132 (N_132,In_325,In_259);
and U133 (N_133,In_327,In_43);
or U134 (N_134,In_95,In_574);
and U135 (N_135,In_533,In_304);
xor U136 (N_136,In_420,In_21);
or U137 (N_137,In_375,In_54);
or U138 (N_138,In_201,In_105);
and U139 (N_139,In_654,In_726);
nor U140 (N_140,In_133,In_173);
or U141 (N_141,In_524,In_28);
or U142 (N_142,In_341,In_448);
and U143 (N_143,In_1,In_614);
and U144 (N_144,In_27,In_499);
and U145 (N_145,In_666,In_118);
nand U146 (N_146,In_365,In_39);
or U147 (N_147,In_37,In_421);
or U148 (N_148,In_548,In_46);
nand U149 (N_149,In_575,In_148);
xnor U150 (N_150,In_224,In_723);
nand U151 (N_151,In_154,In_282);
nand U152 (N_152,In_670,In_493);
nor U153 (N_153,In_51,In_55);
or U154 (N_154,In_564,In_605);
or U155 (N_155,In_40,In_547);
nand U156 (N_156,In_159,In_290);
nor U157 (N_157,In_121,In_650);
nand U158 (N_158,In_529,In_669);
nor U159 (N_159,In_731,In_677);
nor U160 (N_160,In_174,In_517);
and U161 (N_161,In_459,In_657);
nor U162 (N_162,In_663,In_243);
nor U163 (N_163,In_109,In_242);
nor U164 (N_164,In_371,In_474);
or U165 (N_165,In_664,In_230);
and U166 (N_166,In_483,In_713);
nor U167 (N_167,In_244,In_573);
or U168 (N_168,In_124,In_406);
and U169 (N_169,In_692,In_257);
or U170 (N_170,In_652,In_138);
nor U171 (N_171,In_68,In_640);
and U172 (N_172,In_8,In_342);
and U173 (N_173,In_521,In_511);
nor U174 (N_174,In_495,In_250);
nor U175 (N_175,In_457,In_143);
nand U176 (N_176,In_727,In_552);
nor U177 (N_177,In_730,In_425);
nor U178 (N_178,In_431,In_102);
nand U179 (N_179,In_215,In_294);
or U180 (N_180,In_559,In_123);
or U181 (N_181,In_625,In_678);
and U182 (N_182,In_140,In_403);
nand U183 (N_183,In_355,In_268);
and U184 (N_184,In_736,In_707);
or U185 (N_185,In_165,In_262);
and U186 (N_186,In_125,In_26);
and U187 (N_187,In_739,In_260);
nor U188 (N_188,In_343,In_130);
nand U189 (N_189,In_299,In_75);
nand U190 (N_190,In_668,In_194);
and U191 (N_191,In_471,In_701);
and U192 (N_192,In_50,In_449);
nand U193 (N_193,In_497,In_734);
nor U194 (N_194,In_412,In_157);
nand U195 (N_195,In_653,In_200);
and U196 (N_196,In_411,In_570);
and U197 (N_197,In_490,In_370);
or U198 (N_198,In_571,In_592);
or U199 (N_199,In_359,In_354);
and U200 (N_200,In_247,In_672);
and U201 (N_201,In_225,In_719);
and U202 (N_202,In_703,In_276);
or U203 (N_203,In_665,In_373);
or U204 (N_204,In_679,In_631);
nor U205 (N_205,In_2,In_248);
xnor U206 (N_206,In_177,In_197);
nand U207 (N_207,In_275,In_405);
or U208 (N_208,In_708,In_540);
or U209 (N_209,In_34,In_450);
and U210 (N_210,In_324,In_618);
nor U211 (N_211,In_86,In_440);
and U212 (N_212,In_256,In_500);
or U213 (N_213,In_278,In_84);
or U214 (N_214,In_699,In_512);
or U215 (N_215,In_522,In_641);
and U216 (N_216,In_4,In_423);
or U217 (N_217,In_132,In_361);
nor U218 (N_218,In_612,In_464);
or U219 (N_219,In_589,In_408);
or U220 (N_220,In_407,In_400);
xor U221 (N_221,In_310,In_473);
nand U222 (N_222,In_556,In_676);
and U223 (N_223,In_445,In_551);
and U224 (N_224,In_718,In_476);
nor U225 (N_225,In_66,In_307);
and U226 (N_226,In_150,In_155);
nand U227 (N_227,In_743,In_646);
nand U228 (N_228,In_601,In_485);
nor U229 (N_229,In_52,In_339);
and U230 (N_230,In_484,In_7);
or U231 (N_231,In_314,In_312);
nand U232 (N_232,In_323,In_356);
and U233 (N_233,In_176,In_369);
and U234 (N_234,In_70,In_716);
or U235 (N_235,In_306,In_607);
or U236 (N_236,In_580,In_206);
nand U237 (N_237,In_460,In_747);
and U238 (N_238,In_235,In_319);
nand U239 (N_239,In_683,In_56);
nor U240 (N_240,In_688,In_196);
nor U241 (N_241,In_489,In_687);
and U242 (N_242,In_100,In_91);
and U243 (N_243,In_332,In_682);
and U244 (N_244,In_15,In_80);
nor U245 (N_245,In_163,In_237);
nor U246 (N_246,In_379,In_468);
nand U247 (N_247,In_591,In_239);
nor U248 (N_248,In_183,In_322);
and U249 (N_249,In_274,In_151);
nand U250 (N_250,In_172,In_106);
or U251 (N_251,In_409,In_526);
nand U252 (N_252,In_606,In_220);
and U253 (N_253,In_706,In_287);
nand U254 (N_254,In_309,In_338);
and U255 (N_255,In_655,In_210);
nand U256 (N_256,In_232,In_158);
or U257 (N_257,In_581,In_492);
and U258 (N_258,In_443,In_350);
nor U259 (N_259,In_44,In_530);
nand U260 (N_260,In_436,In_502);
nor U261 (N_261,In_507,In_628);
nand U262 (N_262,In_746,In_479);
nand U263 (N_263,In_6,In_611);
or U264 (N_264,In_5,In_430);
nand U265 (N_265,In_583,In_742);
and U266 (N_266,In_112,In_553);
nor U267 (N_267,In_315,In_505);
nand U268 (N_268,In_488,In_89);
nand U269 (N_269,In_398,In_73);
or U270 (N_270,In_481,In_599);
nor U271 (N_271,In_639,In_461);
or U272 (N_272,In_623,In_320);
nand U273 (N_273,In_115,In_415);
or U274 (N_274,In_266,In_390);
and U275 (N_275,In_380,In_22);
or U276 (N_276,In_9,In_169);
nand U277 (N_277,In_212,In_462);
and U278 (N_278,In_188,In_184);
nand U279 (N_279,In_642,In_527);
and U280 (N_280,In_217,In_674);
or U281 (N_281,In_164,In_76);
or U282 (N_282,In_57,In_391);
or U283 (N_283,In_141,In_691);
or U284 (N_284,In_374,In_74);
or U285 (N_285,In_694,In_486);
nor U286 (N_286,In_744,In_396);
and U287 (N_287,In_501,In_596);
nand U288 (N_288,In_61,In_156);
and U289 (N_289,In_598,In_649);
nor U290 (N_290,In_23,In_542);
and U291 (N_291,In_616,In_104);
and U292 (N_292,In_185,In_543);
and U293 (N_293,In_238,In_285);
and U294 (N_294,In_363,In_480);
and U295 (N_295,In_36,In_536);
and U296 (N_296,In_563,In_554);
nor U297 (N_297,In_416,In_579);
nor U298 (N_298,In_660,In_586);
and U299 (N_299,In_58,In_29);
nor U300 (N_300,In_229,In_249);
nor U301 (N_301,In_308,In_748);
nor U302 (N_302,In_209,In_368);
nand U303 (N_303,In_198,In_732);
nor U304 (N_304,In_695,In_64);
nand U305 (N_305,In_77,In_321);
or U306 (N_306,In_422,In_615);
or U307 (N_307,In_671,In_621);
and U308 (N_308,In_291,In_364);
nand U309 (N_309,In_538,In_358);
or U310 (N_310,In_179,In_298);
xnor U311 (N_311,In_251,In_597);
and U312 (N_312,In_632,In_246);
and U313 (N_313,In_634,In_160);
or U314 (N_314,In_424,In_234);
nor U315 (N_315,In_417,In_35);
nand U316 (N_316,In_626,In_569);
nand U317 (N_317,In_709,In_12);
nor U318 (N_318,In_62,In_258);
nand U319 (N_319,In_272,In_446);
and U320 (N_320,In_594,In_271);
or U321 (N_321,In_388,In_537);
or U322 (N_322,In_689,In_608);
or U323 (N_323,In_284,In_539);
nor U324 (N_324,In_203,In_472);
nand U325 (N_325,In_477,In_264);
and U326 (N_326,In_738,In_658);
or U327 (N_327,In_340,In_427);
nand U328 (N_328,In_435,In_167);
nand U329 (N_329,In_136,In_97);
and U330 (N_330,In_366,In_344);
nor U331 (N_331,In_397,In_675);
nand U332 (N_332,In_288,In_335);
or U333 (N_333,In_114,In_25);
nand U334 (N_334,In_724,In_269);
nand U335 (N_335,In_383,In_603);
or U336 (N_336,In_712,In_470);
nor U337 (N_337,In_300,In_353);
and U338 (N_338,In_456,In_24);
nor U339 (N_339,In_567,In_305);
and U340 (N_340,In_139,In_346);
and U341 (N_341,In_447,In_110);
or U342 (N_342,In_651,In_252);
nand U343 (N_343,In_182,In_166);
or U344 (N_344,In_656,In_147);
nor U345 (N_345,In_544,In_419);
or U346 (N_346,In_270,In_289);
nor U347 (N_347,In_204,In_240);
and U348 (N_348,In_241,In_729);
and U349 (N_349,In_171,In_280);
and U350 (N_350,In_721,In_189);
nor U351 (N_351,In_645,In_508);
nand U352 (N_352,In_428,In_541);
nand U353 (N_353,In_128,In_83);
nand U354 (N_354,In_236,In_715);
or U355 (N_355,In_491,In_120);
and U356 (N_356,In_531,In_149);
and U357 (N_357,In_733,In_534);
nor U358 (N_358,In_202,In_334);
nor U359 (N_359,In_467,In_126);
nand U360 (N_360,In_740,In_367);
nor U361 (N_361,In_69,In_509);
nor U362 (N_362,In_330,In_377);
and U363 (N_363,In_222,In_735);
or U364 (N_364,In_680,In_10);
nor U365 (N_365,In_617,In_463);
nand U366 (N_366,In_515,In_454);
nor U367 (N_367,In_33,In_619);
or U368 (N_368,In_429,In_717);
nor U369 (N_369,In_261,In_103);
and U370 (N_370,In_119,In_13);
nor U371 (N_371,In_560,In_19);
nor U372 (N_372,In_404,In_514);
nand U373 (N_373,In_214,In_303);
or U374 (N_374,In_277,In_92);
nand U375 (N_375,In_62,In_588);
nand U376 (N_376,In_437,In_734);
and U377 (N_377,In_177,In_140);
nand U378 (N_378,In_48,In_353);
or U379 (N_379,In_223,In_490);
and U380 (N_380,In_335,In_341);
nor U381 (N_381,In_301,In_514);
or U382 (N_382,In_605,In_369);
or U383 (N_383,In_454,In_598);
and U384 (N_384,In_122,In_92);
and U385 (N_385,In_730,In_542);
nand U386 (N_386,In_603,In_636);
and U387 (N_387,In_236,In_345);
and U388 (N_388,In_285,In_310);
or U389 (N_389,In_167,In_367);
nor U390 (N_390,In_37,In_287);
nor U391 (N_391,In_557,In_142);
nor U392 (N_392,In_460,In_447);
nor U393 (N_393,In_269,In_427);
or U394 (N_394,In_413,In_697);
nor U395 (N_395,In_508,In_373);
nor U396 (N_396,In_417,In_464);
nand U397 (N_397,In_731,In_88);
and U398 (N_398,In_151,In_413);
nand U399 (N_399,In_112,In_728);
nor U400 (N_400,In_97,In_482);
and U401 (N_401,In_439,In_286);
and U402 (N_402,In_607,In_359);
and U403 (N_403,In_260,In_628);
and U404 (N_404,In_143,In_490);
and U405 (N_405,In_486,In_372);
and U406 (N_406,In_719,In_657);
nand U407 (N_407,In_325,In_112);
nor U408 (N_408,In_406,In_73);
or U409 (N_409,In_674,In_704);
and U410 (N_410,In_540,In_236);
or U411 (N_411,In_553,In_215);
and U412 (N_412,In_535,In_64);
and U413 (N_413,In_302,In_58);
or U414 (N_414,In_260,In_63);
nand U415 (N_415,In_33,In_542);
nand U416 (N_416,In_487,In_523);
nand U417 (N_417,In_263,In_115);
or U418 (N_418,In_478,In_396);
or U419 (N_419,In_400,In_89);
and U420 (N_420,In_214,In_713);
and U421 (N_421,In_704,In_247);
and U422 (N_422,In_307,In_120);
or U423 (N_423,In_12,In_428);
nand U424 (N_424,In_631,In_609);
nand U425 (N_425,In_1,In_472);
or U426 (N_426,In_127,In_88);
or U427 (N_427,In_200,In_571);
or U428 (N_428,In_30,In_148);
or U429 (N_429,In_621,In_730);
nand U430 (N_430,In_445,In_186);
nand U431 (N_431,In_675,In_585);
or U432 (N_432,In_74,In_400);
nand U433 (N_433,In_223,In_659);
nand U434 (N_434,In_729,In_92);
or U435 (N_435,In_282,In_42);
nand U436 (N_436,In_325,In_436);
and U437 (N_437,In_239,In_498);
or U438 (N_438,In_214,In_564);
xnor U439 (N_439,In_601,In_495);
and U440 (N_440,In_625,In_536);
and U441 (N_441,In_237,In_105);
nor U442 (N_442,In_705,In_647);
and U443 (N_443,In_494,In_642);
nor U444 (N_444,In_660,In_602);
nand U445 (N_445,In_374,In_326);
xnor U446 (N_446,In_624,In_659);
nand U447 (N_447,In_113,In_579);
xnor U448 (N_448,In_123,In_175);
or U449 (N_449,In_251,In_620);
nor U450 (N_450,In_63,In_745);
or U451 (N_451,In_147,In_631);
or U452 (N_452,In_292,In_604);
nand U453 (N_453,In_99,In_596);
nand U454 (N_454,In_52,In_105);
nand U455 (N_455,In_471,In_359);
or U456 (N_456,In_509,In_514);
or U457 (N_457,In_396,In_414);
nor U458 (N_458,In_482,In_466);
or U459 (N_459,In_699,In_674);
or U460 (N_460,In_175,In_127);
and U461 (N_461,In_594,In_153);
and U462 (N_462,In_164,In_484);
nand U463 (N_463,In_488,In_671);
nand U464 (N_464,In_684,In_486);
and U465 (N_465,In_16,In_573);
and U466 (N_466,In_442,In_670);
or U467 (N_467,In_111,In_360);
and U468 (N_468,In_606,In_189);
and U469 (N_469,In_616,In_591);
and U470 (N_470,In_549,In_310);
or U471 (N_471,In_47,In_379);
or U472 (N_472,In_726,In_187);
nor U473 (N_473,In_717,In_593);
nor U474 (N_474,In_240,In_446);
nor U475 (N_475,In_539,In_443);
or U476 (N_476,In_580,In_266);
nand U477 (N_477,In_721,In_114);
nand U478 (N_478,In_58,In_269);
or U479 (N_479,In_268,In_318);
or U480 (N_480,In_558,In_512);
nand U481 (N_481,In_222,In_599);
or U482 (N_482,In_454,In_131);
or U483 (N_483,In_454,In_501);
nor U484 (N_484,In_187,In_286);
nor U485 (N_485,In_321,In_511);
or U486 (N_486,In_367,In_43);
or U487 (N_487,In_335,In_692);
nor U488 (N_488,In_269,In_334);
or U489 (N_489,In_606,In_730);
nor U490 (N_490,In_53,In_60);
nor U491 (N_491,In_614,In_272);
and U492 (N_492,In_494,In_255);
and U493 (N_493,In_336,In_644);
or U494 (N_494,In_629,In_531);
nor U495 (N_495,In_254,In_235);
nor U496 (N_496,In_567,In_749);
nor U497 (N_497,In_710,In_467);
and U498 (N_498,In_481,In_730);
xnor U499 (N_499,In_747,In_246);
nand U500 (N_500,In_544,In_660);
or U501 (N_501,In_701,In_104);
or U502 (N_502,In_24,In_579);
nor U503 (N_503,In_491,In_456);
nand U504 (N_504,In_27,In_128);
or U505 (N_505,In_576,In_230);
nor U506 (N_506,In_554,In_82);
xor U507 (N_507,In_487,In_334);
or U508 (N_508,In_425,In_86);
nor U509 (N_509,In_446,In_363);
or U510 (N_510,In_13,In_556);
nand U511 (N_511,In_394,In_162);
or U512 (N_512,In_431,In_79);
and U513 (N_513,In_504,In_295);
nand U514 (N_514,In_703,In_205);
or U515 (N_515,In_188,In_150);
nor U516 (N_516,In_715,In_217);
nor U517 (N_517,In_363,In_189);
and U518 (N_518,In_507,In_365);
nand U519 (N_519,In_576,In_245);
or U520 (N_520,In_86,In_19);
and U521 (N_521,In_332,In_563);
nor U522 (N_522,In_636,In_196);
and U523 (N_523,In_409,In_24);
nor U524 (N_524,In_555,In_474);
nor U525 (N_525,In_209,In_454);
nor U526 (N_526,In_596,In_646);
nand U527 (N_527,In_283,In_698);
or U528 (N_528,In_209,In_283);
or U529 (N_529,In_312,In_707);
or U530 (N_530,In_153,In_578);
and U531 (N_531,In_403,In_332);
nand U532 (N_532,In_112,In_42);
or U533 (N_533,In_729,In_240);
or U534 (N_534,In_502,In_181);
and U535 (N_535,In_672,In_747);
nand U536 (N_536,In_257,In_736);
nand U537 (N_537,In_402,In_332);
nand U538 (N_538,In_452,In_42);
or U539 (N_539,In_317,In_223);
and U540 (N_540,In_522,In_402);
and U541 (N_541,In_327,In_203);
nor U542 (N_542,In_208,In_547);
and U543 (N_543,In_423,In_223);
and U544 (N_544,In_576,In_673);
nor U545 (N_545,In_203,In_130);
or U546 (N_546,In_160,In_537);
xor U547 (N_547,In_479,In_653);
and U548 (N_548,In_28,In_272);
and U549 (N_549,In_159,In_691);
or U550 (N_550,In_484,In_720);
nor U551 (N_551,In_534,In_685);
and U552 (N_552,In_631,In_550);
or U553 (N_553,In_461,In_706);
and U554 (N_554,In_195,In_260);
nor U555 (N_555,In_9,In_550);
nor U556 (N_556,In_396,In_19);
nor U557 (N_557,In_541,In_670);
nand U558 (N_558,In_137,In_598);
nand U559 (N_559,In_704,In_123);
nand U560 (N_560,In_290,In_349);
nand U561 (N_561,In_145,In_559);
and U562 (N_562,In_258,In_643);
nor U563 (N_563,In_307,In_9);
nor U564 (N_564,In_379,In_664);
nor U565 (N_565,In_523,In_608);
nor U566 (N_566,In_442,In_187);
nor U567 (N_567,In_411,In_504);
or U568 (N_568,In_311,In_453);
and U569 (N_569,In_559,In_84);
nand U570 (N_570,In_55,In_421);
nand U571 (N_571,In_259,In_623);
or U572 (N_572,In_733,In_503);
and U573 (N_573,In_536,In_721);
and U574 (N_574,In_523,In_558);
and U575 (N_575,In_473,In_383);
and U576 (N_576,In_46,In_326);
or U577 (N_577,In_526,In_19);
and U578 (N_578,In_329,In_388);
nand U579 (N_579,In_311,In_230);
and U580 (N_580,In_516,In_110);
nor U581 (N_581,In_662,In_476);
nand U582 (N_582,In_505,In_35);
and U583 (N_583,In_372,In_496);
nor U584 (N_584,In_380,In_264);
nand U585 (N_585,In_269,In_147);
or U586 (N_586,In_655,In_667);
xor U587 (N_587,In_387,In_676);
nor U588 (N_588,In_8,In_242);
and U589 (N_589,In_602,In_342);
and U590 (N_590,In_405,In_244);
or U591 (N_591,In_371,In_173);
nand U592 (N_592,In_392,In_702);
nand U593 (N_593,In_295,In_719);
nand U594 (N_594,In_131,In_87);
nor U595 (N_595,In_477,In_522);
nand U596 (N_596,In_526,In_254);
and U597 (N_597,In_343,In_293);
nor U598 (N_598,In_192,In_69);
or U599 (N_599,In_247,In_719);
nor U600 (N_600,In_532,In_324);
nand U601 (N_601,In_495,In_695);
and U602 (N_602,In_436,In_407);
nand U603 (N_603,In_352,In_179);
nand U604 (N_604,In_108,In_263);
or U605 (N_605,In_177,In_52);
nor U606 (N_606,In_44,In_260);
and U607 (N_607,In_103,In_722);
nor U608 (N_608,In_362,In_425);
nand U609 (N_609,In_204,In_586);
and U610 (N_610,In_582,In_247);
and U611 (N_611,In_332,In_736);
and U612 (N_612,In_564,In_560);
or U613 (N_613,In_602,In_81);
nand U614 (N_614,In_430,In_670);
and U615 (N_615,In_255,In_556);
or U616 (N_616,In_735,In_554);
nor U617 (N_617,In_318,In_92);
or U618 (N_618,In_588,In_15);
nor U619 (N_619,In_19,In_172);
xnor U620 (N_620,In_652,In_392);
and U621 (N_621,In_357,In_180);
nor U622 (N_622,In_683,In_681);
and U623 (N_623,In_195,In_270);
or U624 (N_624,In_473,In_152);
nand U625 (N_625,In_690,In_150);
and U626 (N_626,In_447,In_720);
nand U627 (N_627,In_569,In_253);
nor U628 (N_628,In_50,In_73);
nand U629 (N_629,In_328,In_437);
nor U630 (N_630,In_316,In_291);
nor U631 (N_631,In_20,In_137);
or U632 (N_632,In_452,In_378);
or U633 (N_633,In_277,In_224);
or U634 (N_634,In_270,In_425);
nand U635 (N_635,In_261,In_530);
nor U636 (N_636,In_658,In_741);
nand U637 (N_637,In_573,In_569);
nand U638 (N_638,In_281,In_190);
and U639 (N_639,In_544,In_33);
nand U640 (N_640,In_255,In_428);
nand U641 (N_641,In_137,In_684);
and U642 (N_642,In_116,In_695);
nand U643 (N_643,In_218,In_334);
nand U644 (N_644,In_10,In_448);
nor U645 (N_645,In_545,In_315);
nor U646 (N_646,In_575,In_432);
nand U647 (N_647,In_220,In_613);
or U648 (N_648,In_253,In_648);
and U649 (N_649,In_57,In_196);
nor U650 (N_650,In_653,In_545);
and U651 (N_651,In_379,In_410);
and U652 (N_652,In_465,In_392);
or U653 (N_653,In_613,In_718);
nand U654 (N_654,In_189,In_529);
nand U655 (N_655,In_669,In_4);
and U656 (N_656,In_669,In_551);
nand U657 (N_657,In_252,In_332);
or U658 (N_658,In_374,In_161);
xnor U659 (N_659,In_68,In_104);
or U660 (N_660,In_592,In_373);
and U661 (N_661,In_239,In_253);
nor U662 (N_662,In_348,In_282);
and U663 (N_663,In_99,In_329);
nor U664 (N_664,In_384,In_345);
and U665 (N_665,In_396,In_273);
or U666 (N_666,In_740,In_624);
or U667 (N_667,In_2,In_176);
or U668 (N_668,In_311,In_246);
nor U669 (N_669,In_541,In_38);
nor U670 (N_670,In_300,In_544);
or U671 (N_671,In_88,In_312);
nor U672 (N_672,In_597,In_549);
and U673 (N_673,In_146,In_57);
nand U674 (N_674,In_275,In_628);
and U675 (N_675,In_47,In_343);
or U676 (N_676,In_361,In_625);
nand U677 (N_677,In_736,In_604);
nand U678 (N_678,In_644,In_593);
or U679 (N_679,In_137,In_563);
nand U680 (N_680,In_582,In_302);
nor U681 (N_681,In_577,In_475);
and U682 (N_682,In_96,In_40);
nor U683 (N_683,In_147,In_260);
nand U684 (N_684,In_384,In_403);
and U685 (N_685,In_521,In_403);
nor U686 (N_686,In_469,In_23);
and U687 (N_687,In_726,In_628);
nor U688 (N_688,In_471,In_421);
nand U689 (N_689,In_48,In_157);
nor U690 (N_690,In_646,In_303);
nand U691 (N_691,In_6,In_494);
or U692 (N_692,In_567,In_172);
nor U693 (N_693,In_81,In_707);
or U694 (N_694,In_352,In_142);
and U695 (N_695,In_294,In_124);
or U696 (N_696,In_699,In_23);
nand U697 (N_697,In_407,In_590);
and U698 (N_698,In_570,In_155);
or U699 (N_699,In_663,In_638);
nor U700 (N_700,In_267,In_672);
nor U701 (N_701,In_688,In_159);
or U702 (N_702,In_531,In_64);
or U703 (N_703,In_131,In_353);
nor U704 (N_704,In_562,In_33);
or U705 (N_705,In_426,In_309);
nand U706 (N_706,In_578,In_1);
or U707 (N_707,In_371,In_200);
and U708 (N_708,In_131,In_376);
nor U709 (N_709,In_384,In_649);
xnor U710 (N_710,In_383,In_737);
nand U711 (N_711,In_605,In_748);
nor U712 (N_712,In_415,In_653);
nor U713 (N_713,In_741,In_335);
and U714 (N_714,In_519,In_601);
or U715 (N_715,In_712,In_643);
nand U716 (N_716,In_179,In_202);
and U717 (N_717,In_288,In_600);
or U718 (N_718,In_671,In_117);
nand U719 (N_719,In_684,In_17);
and U720 (N_720,In_315,In_639);
or U721 (N_721,In_374,In_357);
or U722 (N_722,In_745,In_140);
nand U723 (N_723,In_64,In_604);
nand U724 (N_724,In_538,In_688);
nand U725 (N_725,In_639,In_436);
and U726 (N_726,In_298,In_557);
nand U727 (N_727,In_259,In_98);
nor U728 (N_728,In_383,In_49);
nor U729 (N_729,In_121,In_273);
nor U730 (N_730,In_1,In_358);
and U731 (N_731,In_354,In_360);
or U732 (N_732,In_621,In_182);
and U733 (N_733,In_184,In_47);
nor U734 (N_734,In_178,In_736);
nand U735 (N_735,In_407,In_634);
or U736 (N_736,In_227,In_148);
and U737 (N_737,In_352,In_365);
and U738 (N_738,In_557,In_32);
nor U739 (N_739,In_571,In_208);
nor U740 (N_740,In_729,In_527);
or U741 (N_741,In_361,In_615);
nor U742 (N_742,In_120,In_612);
or U743 (N_743,In_687,In_209);
nand U744 (N_744,In_686,In_440);
nor U745 (N_745,In_514,In_435);
and U746 (N_746,In_698,In_210);
and U747 (N_747,In_686,In_401);
or U748 (N_748,In_413,In_146);
nor U749 (N_749,In_453,In_739);
nand U750 (N_750,In_719,In_406);
and U751 (N_751,In_511,In_694);
or U752 (N_752,In_276,In_678);
nand U753 (N_753,In_46,In_579);
xor U754 (N_754,In_736,In_493);
nand U755 (N_755,In_381,In_216);
nor U756 (N_756,In_208,In_654);
and U757 (N_757,In_624,In_735);
nor U758 (N_758,In_46,In_55);
nand U759 (N_759,In_737,In_483);
or U760 (N_760,In_241,In_64);
or U761 (N_761,In_450,In_466);
nand U762 (N_762,In_428,In_625);
or U763 (N_763,In_401,In_405);
nand U764 (N_764,In_722,In_99);
nand U765 (N_765,In_542,In_415);
nand U766 (N_766,In_403,In_285);
or U767 (N_767,In_52,In_585);
and U768 (N_768,In_284,In_584);
and U769 (N_769,In_701,In_43);
nor U770 (N_770,In_523,In_355);
or U771 (N_771,In_442,In_487);
and U772 (N_772,In_230,In_569);
or U773 (N_773,In_250,In_85);
nor U774 (N_774,In_634,In_415);
or U775 (N_775,In_166,In_360);
nor U776 (N_776,In_408,In_141);
nor U777 (N_777,In_90,In_643);
or U778 (N_778,In_424,In_589);
and U779 (N_779,In_365,In_748);
nor U780 (N_780,In_260,In_649);
nand U781 (N_781,In_53,In_444);
nand U782 (N_782,In_208,In_356);
or U783 (N_783,In_426,In_370);
or U784 (N_784,In_456,In_201);
and U785 (N_785,In_68,In_202);
or U786 (N_786,In_132,In_7);
or U787 (N_787,In_46,In_138);
and U788 (N_788,In_4,In_413);
nand U789 (N_789,In_97,In_293);
and U790 (N_790,In_41,In_609);
or U791 (N_791,In_105,In_361);
and U792 (N_792,In_738,In_666);
and U793 (N_793,In_290,In_749);
nor U794 (N_794,In_742,In_108);
or U795 (N_795,In_390,In_382);
and U796 (N_796,In_370,In_522);
or U797 (N_797,In_515,In_313);
nand U798 (N_798,In_284,In_182);
and U799 (N_799,In_19,In_653);
nor U800 (N_800,In_232,In_634);
or U801 (N_801,In_569,In_214);
nor U802 (N_802,In_359,In_22);
nor U803 (N_803,In_128,In_9);
nand U804 (N_804,In_23,In_166);
nand U805 (N_805,In_2,In_373);
nor U806 (N_806,In_120,In_739);
xnor U807 (N_807,In_194,In_365);
nor U808 (N_808,In_604,In_634);
nand U809 (N_809,In_440,In_688);
nor U810 (N_810,In_576,In_144);
nand U811 (N_811,In_329,In_493);
nor U812 (N_812,In_709,In_337);
nand U813 (N_813,In_663,In_569);
or U814 (N_814,In_365,In_279);
nor U815 (N_815,In_476,In_671);
nor U816 (N_816,In_274,In_569);
nand U817 (N_817,In_123,In_147);
and U818 (N_818,In_156,In_408);
nor U819 (N_819,In_638,In_312);
xor U820 (N_820,In_472,In_566);
nand U821 (N_821,In_375,In_74);
nor U822 (N_822,In_385,In_649);
and U823 (N_823,In_431,In_5);
or U824 (N_824,In_490,In_12);
and U825 (N_825,In_63,In_46);
and U826 (N_826,In_640,In_678);
and U827 (N_827,In_437,In_700);
nand U828 (N_828,In_294,In_164);
and U829 (N_829,In_538,In_653);
or U830 (N_830,In_538,In_80);
and U831 (N_831,In_708,In_570);
and U832 (N_832,In_171,In_707);
nor U833 (N_833,In_108,In_505);
or U834 (N_834,In_265,In_132);
nor U835 (N_835,In_743,In_228);
nor U836 (N_836,In_340,In_628);
and U837 (N_837,In_596,In_257);
nand U838 (N_838,In_83,In_2);
and U839 (N_839,In_353,In_590);
nand U840 (N_840,In_198,In_378);
nor U841 (N_841,In_464,In_620);
nor U842 (N_842,In_568,In_289);
nor U843 (N_843,In_468,In_312);
or U844 (N_844,In_221,In_540);
nand U845 (N_845,In_707,In_121);
or U846 (N_846,In_315,In_478);
nor U847 (N_847,In_712,In_260);
or U848 (N_848,In_77,In_99);
nand U849 (N_849,In_147,In_454);
and U850 (N_850,In_55,In_627);
or U851 (N_851,In_110,In_83);
and U852 (N_852,In_236,In_502);
or U853 (N_853,In_728,In_258);
nand U854 (N_854,In_279,In_295);
nor U855 (N_855,In_324,In_302);
nor U856 (N_856,In_237,In_716);
or U857 (N_857,In_469,In_106);
or U858 (N_858,In_178,In_505);
and U859 (N_859,In_596,In_290);
and U860 (N_860,In_552,In_391);
nor U861 (N_861,In_577,In_617);
or U862 (N_862,In_34,In_257);
nor U863 (N_863,In_104,In_552);
nand U864 (N_864,In_239,In_74);
nor U865 (N_865,In_374,In_486);
and U866 (N_866,In_232,In_92);
nor U867 (N_867,In_124,In_565);
and U868 (N_868,In_434,In_87);
nor U869 (N_869,In_608,In_403);
or U870 (N_870,In_323,In_372);
nor U871 (N_871,In_464,In_633);
nor U872 (N_872,In_334,In_591);
and U873 (N_873,In_736,In_168);
or U874 (N_874,In_523,In_405);
or U875 (N_875,In_298,In_169);
nor U876 (N_876,In_656,In_570);
nand U877 (N_877,In_435,In_724);
nor U878 (N_878,In_519,In_388);
nand U879 (N_879,In_467,In_196);
or U880 (N_880,In_378,In_453);
nor U881 (N_881,In_490,In_567);
nor U882 (N_882,In_445,In_41);
or U883 (N_883,In_710,In_425);
nor U884 (N_884,In_618,In_201);
nand U885 (N_885,In_293,In_26);
and U886 (N_886,In_672,In_76);
nor U887 (N_887,In_43,In_587);
or U888 (N_888,In_318,In_574);
or U889 (N_889,In_448,In_460);
or U890 (N_890,In_265,In_502);
nor U891 (N_891,In_279,In_15);
or U892 (N_892,In_55,In_429);
or U893 (N_893,In_421,In_732);
nor U894 (N_894,In_590,In_701);
or U895 (N_895,In_137,In_348);
and U896 (N_896,In_656,In_125);
and U897 (N_897,In_180,In_342);
nand U898 (N_898,In_184,In_544);
or U899 (N_899,In_79,In_256);
nor U900 (N_900,In_696,In_199);
and U901 (N_901,In_386,In_484);
and U902 (N_902,In_488,In_118);
or U903 (N_903,In_49,In_355);
or U904 (N_904,In_482,In_463);
or U905 (N_905,In_136,In_25);
or U906 (N_906,In_227,In_413);
nor U907 (N_907,In_464,In_262);
and U908 (N_908,In_306,In_573);
nand U909 (N_909,In_290,In_464);
nand U910 (N_910,In_702,In_57);
nand U911 (N_911,In_438,In_53);
nand U912 (N_912,In_504,In_355);
nand U913 (N_913,In_1,In_79);
and U914 (N_914,In_277,In_61);
nor U915 (N_915,In_364,In_102);
nor U916 (N_916,In_157,In_279);
nor U917 (N_917,In_128,In_437);
nor U918 (N_918,In_686,In_600);
nor U919 (N_919,In_27,In_646);
nor U920 (N_920,In_378,In_627);
nor U921 (N_921,In_152,In_314);
nand U922 (N_922,In_584,In_612);
nand U923 (N_923,In_416,In_622);
and U924 (N_924,In_614,In_20);
nor U925 (N_925,In_295,In_711);
and U926 (N_926,In_634,In_159);
nand U927 (N_927,In_62,In_107);
nand U928 (N_928,In_75,In_214);
or U929 (N_929,In_70,In_656);
nor U930 (N_930,In_363,In_22);
nand U931 (N_931,In_364,In_590);
nor U932 (N_932,In_732,In_673);
and U933 (N_933,In_243,In_17);
nand U934 (N_934,In_563,In_631);
and U935 (N_935,In_254,In_452);
or U936 (N_936,In_726,In_405);
nor U937 (N_937,In_230,In_644);
nand U938 (N_938,In_689,In_198);
and U939 (N_939,In_491,In_160);
nor U940 (N_940,In_156,In_682);
nor U941 (N_941,In_364,In_551);
nand U942 (N_942,In_694,In_709);
nand U943 (N_943,In_741,In_272);
xor U944 (N_944,In_91,In_130);
and U945 (N_945,In_451,In_296);
and U946 (N_946,In_680,In_145);
nor U947 (N_947,In_481,In_3);
and U948 (N_948,In_198,In_34);
nand U949 (N_949,In_181,In_687);
and U950 (N_950,In_2,In_296);
nand U951 (N_951,In_736,In_517);
and U952 (N_952,In_198,In_384);
and U953 (N_953,In_55,In_576);
or U954 (N_954,In_303,In_178);
nor U955 (N_955,In_564,In_515);
or U956 (N_956,In_26,In_452);
nand U957 (N_957,In_53,In_439);
nand U958 (N_958,In_482,In_181);
and U959 (N_959,In_522,In_520);
or U960 (N_960,In_726,In_329);
or U961 (N_961,In_166,In_3);
or U962 (N_962,In_156,In_448);
nor U963 (N_963,In_536,In_10);
or U964 (N_964,In_732,In_213);
and U965 (N_965,In_33,In_524);
and U966 (N_966,In_320,In_51);
and U967 (N_967,In_348,In_645);
and U968 (N_968,In_721,In_458);
nand U969 (N_969,In_488,In_691);
nand U970 (N_970,In_691,In_350);
and U971 (N_971,In_105,In_711);
nor U972 (N_972,In_163,In_528);
and U973 (N_973,In_337,In_347);
nor U974 (N_974,In_525,In_318);
or U975 (N_975,In_357,In_402);
nor U976 (N_976,In_286,In_679);
and U977 (N_977,In_726,In_326);
and U978 (N_978,In_264,In_580);
or U979 (N_979,In_739,In_413);
nand U980 (N_980,In_185,In_263);
nand U981 (N_981,In_362,In_279);
nand U982 (N_982,In_501,In_203);
xnor U983 (N_983,In_321,In_194);
nor U984 (N_984,In_228,In_370);
nand U985 (N_985,In_407,In_408);
nor U986 (N_986,In_629,In_650);
nor U987 (N_987,In_439,In_496);
and U988 (N_988,In_88,In_511);
or U989 (N_989,In_536,In_583);
and U990 (N_990,In_443,In_63);
or U991 (N_991,In_722,In_97);
nor U992 (N_992,In_227,In_209);
nor U993 (N_993,In_178,In_493);
nor U994 (N_994,In_156,In_338);
nand U995 (N_995,In_676,In_62);
nand U996 (N_996,In_169,In_1);
nand U997 (N_997,In_99,In_462);
and U998 (N_998,In_174,In_172);
or U999 (N_999,In_388,In_638);
nor U1000 (N_1000,In_40,In_292);
or U1001 (N_1001,In_247,In_170);
and U1002 (N_1002,In_489,In_54);
nor U1003 (N_1003,In_173,In_246);
or U1004 (N_1004,In_103,In_383);
and U1005 (N_1005,In_716,In_229);
or U1006 (N_1006,In_28,In_581);
or U1007 (N_1007,In_131,In_443);
nand U1008 (N_1008,In_562,In_80);
or U1009 (N_1009,In_336,In_327);
nor U1010 (N_1010,In_303,In_122);
nor U1011 (N_1011,In_383,In_57);
nand U1012 (N_1012,In_367,In_749);
or U1013 (N_1013,In_749,In_31);
nor U1014 (N_1014,In_700,In_653);
nor U1015 (N_1015,In_204,In_651);
nor U1016 (N_1016,In_423,In_411);
or U1017 (N_1017,In_97,In_740);
and U1018 (N_1018,In_148,In_425);
or U1019 (N_1019,In_241,In_664);
or U1020 (N_1020,In_699,In_413);
or U1021 (N_1021,In_87,In_385);
or U1022 (N_1022,In_81,In_455);
and U1023 (N_1023,In_574,In_229);
and U1024 (N_1024,In_88,In_275);
nor U1025 (N_1025,In_499,In_68);
nand U1026 (N_1026,In_620,In_693);
nor U1027 (N_1027,In_507,In_174);
nor U1028 (N_1028,In_249,In_578);
nand U1029 (N_1029,In_582,In_434);
nor U1030 (N_1030,In_619,In_654);
nand U1031 (N_1031,In_207,In_665);
nand U1032 (N_1032,In_213,In_123);
nand U1033 (N_1033,In_613,In_617);
or U1034 (N_1034,In_347,In_598);
and U1035 (N_1035,In_320,In_358);
nor U1036 (N_1036,In_84,In_172);
and U1037 (N_1037,In_458,In_631);
or U1038 (N_1038,In_526,In_186);
or U1039 (N_1039,In_69,In_396);
nand U1040 (N_1040,In_480,In_589);
nand U1041 (N_1041,In_244,In_563);
or U1042 (N_1042,In_182,In_513);
and U1043 (N_1043,In_681,In_288);
and U1044 (N_1044,In_676,In_65);
nand U1045 (N_1045,In_301,In_512);
nor U1046 (N_1046,In_35,In_740);
nor U1047 (N_1047,In_641,In_352);
nor U1048 (N_1048,In_228,In_514);
or U1049 (N_1049,In_151,In_262);
and U1050 (N_1050,In_481,In_139);
nor U1051 (N_1051,In_749,In_165);
or U1052 (N_1052,In_666,In_28);
and U1053 (N_1053,In_731,In_570);
nand U1054 (N_1054,In_249,In_184);
nand U1055 (N_1055,In_82,In_258);
and U1056 (N_1056,In_487,In_176);
and U1057 (N_1057,In_416,In_395);
and U1058 (N_1058,In_328,In_462);
nor U1059 (N_1059,In_443,In_96);
and U1060 (N_1060,In_514,In_483);
nand U1061 (N_1061,In_456,In_192);
and U1062 (N_1062,In_208,In_98);
nand U1063 (N_1063,In_45,In_471);
and U1064 (N_1064,In_352,In_328);
and U1065 (N_1065,In_721,In_733);
and U1066 (N_1066,In_713,In_158);
or U1067 (N_1067,In_197,In_376);
nand U1068 (N_1068,In_428,In_275);
nand U1069 (N_1069,In_427,In_663);
nor U1070 (N_1070,In_392,In_525);
and U1071 (N_1071,In_54,In_346);
nand U1072 (N_1072,In_231,In_439);
nor U1073 (N_1073,In_321,In_375);
nor U1074 (N_1074,In_597,In_28);
or U1075 (N_1075,In_602,In_442);
and U1076 (N_1076,In_338,In_626);
and U1077 (N_1077,In_621,In_205);
nand U1078 (N_1078,In_320,In_409);
nand U1079 (N_1079,In_154,In_87);
or U1080 (N_1080,In_693,In_583);
or U1081 (N_1081,In_212,In_737);
nand U1082 (N_1082,In_155,In_113);
nor U1083 (N_1083,In_288,In_505);
and U1084 (N_1084,In_662,In_730);
nand U1085 (N_1085,In_162,In_708);
nor U1086 (N_1086,In_222,In_186);
nand U1087 (N_1087,In_341,In_281);
nor U1088 (N_1088,In_536,In_627);
and U1089 (N_1089,In_231,In_334);
nand U1090 (N_1090,In_43,In_289);
nand U1091 (N_1091,In_94,In_149);
and U1092 (N_1092,In_565,In_211);
nand U1093 (N_1093,In_215,In_287);
and U1094 (N_1094,In_512,In_698);
nand U1095 (N_1095,In_221,In_704);
nor U1096 (N_1096,In_701,In_406);
nor U1097 (N_1097,In_511,In_512);
and U1098 (N_1098,In_500,In_667);
nand U1099 (N_1099,In_665,In_282);
nor U1100 (N_1100,In_209,In_300);
nor U1101 (N_1101,In_604,In_76);
nor U1102 (N_1102,In_96,In_494);
nor U1103 (N_1103,In_630,In_615);
or U1104 (N_1104,In_749,In_735);
nor U1105 (N_1105,In_173,In_474);
or U1106 (N_1106,In_289,In_302);
xnor U1107 (N_1107,In_642,In_688);
or U1108 (N_1108,In_644,In_218);
nand U1109 (N_1109,In_417,In_538);
or U1110 (N_1110,In_87,In_279);
nor U1111 (N_1111,In_266,In_21);
nand U1112 (N_1112,In_734,In_325);
nand U1113 (N_1113,In_194,In_323);
or U1114 (N_1114,In_560,In_109);
or U1115 (N_1115,In_322,In_235);
and U1116 (N_1116,In_58,In_401);
or U1117 (N_1117,In_258,In_93);
nor U1118 (N_1118,In_358,In_5);
or U1119 (N_1119,In_661,In_621);
and U1120 (N_1120,In_707,In_230);
and U1121 (N_1121,In_671,In_324);
and U1122 (N_1122,In_571,In_691);
or U1123 (N_1123,In_191,In_246);
and U1124 (N_1124,In_633,In_29);
and U1125 (N_1125,In_620,In_294);
or U1126 (N_1126,In_593,In_253);
xor U1127 (N_1127,In_604,In_135);
nor U1128 (N_1128,In_361,In_121);
xnor U1129 (N_1129,In_64,In_19);
nor U1130 (N_1130,In_18,In_728);
nor U1131 (N_1131,In_595,In_647);
and U1132 (N_1132,In_292,In_160);
or U1133 (N_1133,In_383,In_172);
nand U1134 (N_1134,In_382,In_45);
and U1135 (N_1135,In_299,In_536);
or U1136 (N_1136,In_413,In_140);
and U1137 (N_1137,In_311,In_160);
nand U1138 (N_1138,In_428,In_453);
or U1139 (N_1139,In_175,In_121);
nand U1140 (N_1140,In_473,In_409);
and U1141 (N_1141,In_723,In_40);
or U1142 (N_1142,In_46,In_246);
nand U1143 (N_1143,In_318,In_192);
nor U1144 (N_1144,In_515,In_309);
and U1145 (N_1145,In_705,In_83);
nand U1146 (N_1146,In_690,In_78);
and U1147 (N_1147,In_61,In_570);
and U1148 (N_1148,In_347,In_429);
or U1149 (N_1149,In_548,In_27);
nor U1150 (N_1150,In_383,In_705);
nor U1151 (N_1151,In_374,In_730);
nand U1152 (N_1152,In_557,In_725);
nor U1153 (N_1153,In_370,In_587);
and U1154 (N_1154,In_439,In_264);
nor U1155 (N_1155,In_533,In_421);
nand U1156 (N_1156,In_151,In_253);
nand U1157 (N_1157,In_615,In_367);
and U1158 (N_1158,In_337,In_193);
nor U1159 (N_1159,In_461,In_419);
or U1160 (N_1160,In_253,In_495);
or U1161 (N_1161,In_210,In_518);
nor U1162 (N_1162,In_330,In_60);
or U1163 (N_1163,In_568,In_78);
and U1164 (N_1164,In_549,In_592);
or U1165 (N_1165,In_649,In_36);
or U1166 (N_1166,In_560,In_725);
nand U1167 (N_1167,In_670,In_55);
nor U1168 (N_1168,In_25,In_13);
and U1169 (N_1169,In_319,In_672);
or U1170 (N_1170,In_529,In_349);
or U1171 (N_1171,In_638,In_465);
and U1172 (N_1172,In_680,In_218);
nor U1173 (N_1173,In_71,In_520);
nor U1174 (N_1174,In_575,In_258);
nand U1175 (N_1175,In_196,In_35);
and U1176 (N_1176,In_688,In_383);
nand U1177 (N_1177,In_393,In_216);
nor U1178 (N_1178,In_526,In_502);
or U1179 (N_1179,In_466,In_571);
and U1180 (N_1180,In_236,In_53);
nor U1181 (N_1181,In_95,In_609);
nor U1182 (N_1182,In_715,In_314);
or U1183 (N_1183,In_513,In_711);
nand U1184 (N_1184,In_665,In_96);
and U1185 (N_1185,In_36,In_332);
nor U1186 (N_1186,In_672,In_277);
or U1187 (N_1187,In_555,In_239);
nor U1188 (N_1188,In_685,In_259);
nor U1189 (N_1189,In_629,In_745);
nand U1190 (N_1190,In_305,In_367);
nand U1191 (N_1191,In_115,In_223);
xnor U1192 (N_1192,In_366,In_421);
and U1193 (N_1193,In_148,In_716);
nand U1194 (N_1194,In_238,In_128);
and U1195 (N_1195,In_543,In_59);
and U1196 (N_1196,In_380,In_590);
nand U1197 (N_1197,In_587,In_58);
nor U1198 (N_1198,In_737,In_295);
nand U1199 (N_1199,In_600,In_171);
and U1200 (N_1200,In_581,In_395);
nor U1201 (N_1201,In_545,In_283);
nor U1202 (N_1202,In_703,In_115);
nand U1203 (N_1203,In_607,In_219);
nand U1204 (N_1204,In_495,In_21);
or U1205 (N_1205,In_212,In_717);
and U1206 (N_1206,In_392,In_123);
or U1207 (N_1207,In_634,In_595);
or U1208 (N_1208,In_495,In_288);
nor U1209 (N_1209,In_209,In_10);
and U1210 (N_1210,In_514,In_701);
or U1211 (N_1211,In_661,In_591);
and U1212 (N_1212,In_565,In_451);
or U1213 (N_1213,In_364,In_336);
nand U1214 (N_1214,In_73,In_491);
nor U1215 (N_1215,In_108,In_377);
nand U1216 (N_1216,In_689,In_598);
nor U1217 (N_1217,In_658,In_227);
and U1218 (N_1218,In_286,In_597);
nand U1219 (N_1219,In_644,In_725);
nand U1220 (N_1220,In_728,In_69);
or U1221 (N_1221,In_572,In_178);
and U1222 (N_1222,In_11,In_584);
and U1223 (N_1223,In_619,In_328);
and U1224 (N_1224,In_372,In_330);
or U1225 (N_1225,In_161,In_116);
or U1226 (N_1226,In_342,In_200);
nor U1227 (N_1227,In_202,In_295);
nor U1228 (N_1228,In_683,In_257);
or U1229 (N_1229,In_5,In_474);
and U1230 (N_1230,In_612,In_407);
or U1231 (N_1231,In_304,In_395);
and U1232 (N_1232,In_44,In_701);
and U1233 (N_1233,In_623,In_294);
and U1234 (N_1234,In_19,In_439);
nor U1235 (N_1235,In_78,In_134);
xor U1236 (N_1236,In_44,In_363);
or U1237 (N_1237,In_467,In_351);
nand U1238 (N_1238,In_79,In_388);
or U1239 (N_1239,In_432,In_271);
nor U1240 (N_1240,In_13,In_19);
or U1241 (N_1241,In_203,In_641);
nor U1242 (N_1242,In_589,In_429);
nand U1243 (N_1243,In_488,In_683);
nor U1244 (N_1244,In_144,In_6);
and U1245 (N_1245,In_182,In_509);
or U1246 (N_1246,In_703,In_340);
nand U1247 (N_1247,In_308,In_196);
nor U1248 (N_1248,In_367,In_218);
nor U1249 (N_1249,In_151,In_650);
or U1250 (N_1250,In_339,In_576);
nand U1251 (N_1251,In_452,In_364);
or U1252 (N_1252,In_565,In_77);
nor U1253 (N_1253,In_194,In_45);
nand U1254 (N_1254,In_501,In_547);
and U1255 (N_1255,In_221,In_588);
and U1256 (N_1256,In_437,In_301);
nor U1257 (N_1257,In_712,In_102);
or U1258 (N_1258,In_39,In_717);
or U1259 (N_1259,In_226,In_522);
or U1260 (N_1260,In_174,In_561);
nor U1261 (N_1261,In_589,In_679);
and U1262 (N_1262,In_736,In_569);
or U1263 (N_1263,In_62,In_311);
or U1264 (N_1264,In_688,In_467);
nand U1265 (N_1265,In_87,In_49);
nand U1266 (N_1266,In_353,In_745);
and U1267 (N_1267,In_662,In_350);
and U1268 (N_1268,In_435,In_14);
or U1269 (N_1269,In_668,In_256);
nand U1270 (N_1270,In_464,In_663);
nor U1271 (N_1271,In_647,In_67);
or U1272 (N_1272,In_259,In_36);
nor U1273 (N_1273,In_625,In_698);
or U1274 (N_1274,In_748,In_190);
nor U1275 (N_1275,In_235,In_393);
and U1276 (N_1276,In_110,In_628);
nand U1277 (N_1277,In_635,In_269);
nor U1278 (N_1278,In_229,In_696);
nor U1279 (N_1279,In_278,In_374);
nand U1280 (N_1280,In_395,In_689);
or U1281 (N_1281,In_613,In_647);
nor U1282 (N_1282,In_243,In_385);
nor U1283 (N_1283,In_342,In_701);
and U1284 (N_1284,In_641,In_703);
nor U1285 (N_1285,In_676,In_637);
nor U1286 (N_1286,In_616,In_252);
nor U1287 (N_1287,In_133,In_400);
and U1288 (N_1288,In_709,In_599);
nor U1289 (N_1289,In_741,In_255);
nor U1290 (N_1290,In_143,In_96);
or U1291 (N_1291,In_157,In_128);
or U1292 (N_1292,In_113,In_81);
or U1293 (N_1293,In_708,In_139);
nor U1294 (N_1294,In_345,In_548);
nand U1295 (N_1295,In_563,In_131);
and U1296 (N_1296,In_522,In_559);
nand U1297 (N_1297,In_119,In_622);
nor U1298 (N_1298,In_312,In_343);
or U1299 (N_1299,In_478,In_62);
and U1300 (N_1300,In_249,In_525);
nand U1301 (N_1301,In_423,In_286);
or U1302 (N_1302,In_159,In_676);
nand U1303 (N_1303,In_452,In_613);
nand U1304 (N_1304,In_22,In_406);
nor U1305 (N_1305,In_21,In_330);
and U1306 (N_1306,In_113,In_236);
nor U1307 (N_1307,In_500,In_338);
and U1308 (N_1308,In_214,In_322);
nand U1309 (N_1309,In_624,In_368);
nor U1310 (N_1310,In_417,In_191);
or U1311 (N_1311,In_53,In_517);
nor U1312 (N_1312,In_263,In_132);
nor U1313 (N_1313,In_382,In_617);
or U1314 (N_1314,In_151,In_556);
nor U1315 (N_1315,In_122,In_669);
nor U1316 (N_1316,In_210,In_17);
and U1317 (N_1317,In_257,In_319);
and U1318 (N_1318,In_350,In_274);
nor U1319 (N_1319,In_173,In_383);
nor U1320 (N_1320,In_315,In_404);
or U1321 (N_1321,In_234,In_197);
and U1322 (N_1322,In_422,In_623);
nor U1323 (N_1323,In_275,In_35);
and U1324 (N_1324,In_193,In_651);
and U1325 (N_1325,In_380,In_79);
and U1326 (N_1326,In_396,In_307);
nand U1327 (N_1327,In_75,In_376);
and U1328 (N_1328,In_100,In_652);
or U1329 (N_1329,In_313,In_520);
nor U1330 (N_1330,In_713,In_478);
nand U1331 (N_1331,In_189,In_95);
or U1332 (N_1332,In_243,In_92);
or U1333 (N_1333,In_11,In_372);
nand U1334 (N_1334,In_138,In_310);
nand U1335 (N_1335,In_733,In_681);
or U1336 (N_1336,In_505,In_455);
nor U1337 (N_1337,In_394,In_210);
nand U1338 (N_1338,In_189,In_84);
nand U1339 (N_1339,In_168,In_737);
nor U1340 (N_1340,In_361,In_464);
and U1341 (N_1341,In_553,In_435);
and U1342 (N_1342,In_542,In_247);
nor U1343 (N_1343,In_74,In_500);
or U1344 (N_1344,In_563,In_351);
nor U1345 (N_1345,In_650,In_171);
and U1346 (N_1346,In_527,In_204);
nand U1347 (N_1347,In_184,In_322);
and U1348 (N_1348,In_196,In_445);
nor U1349 (N_1349,In_91,In_625);
nand U1350 (N_1350,In_583,In_214);
nor U1351 (N_1351,In_155,In_529);
nor U1352 (N_1352,In_496,In_557);
nor U1353 (N_1353,In_552,In_226);
and U1354 (N_1354,In_59,In_508);
nand U1355 (N_1355,In_302,In_238);
or U1356 (N_1356,In_106,In_447);
or U1357 (N_1357,In_447,In_442);
or U1358 (N_1358,In_482,In_332);
nand U1359 (N_1359,In_218,In_328);
nor U1360 (N_1360,In_29,In_553);
and U1361 (N_1361,In_168,In_606);
nor U1362 (N_1362,In_644,In_434);
nor U1363 (N_1363,In_745,In_464);
nand U1364 (N_1364,In_622,In_324);
nand U1365 (N_1365,In_592,In_8);
nor U1366 (N_1366,In_718,In_594);
and U1367 (N_1367,In_394,In_431);
nand U1368 (N_1368,In_501,In_516);
nand U1369 (N_1369,In_688,In_362);
xor U1370 (N_1370,In_146,In_440);
and U1371 (N_1371,In_12,In_547);
nor U1372 (N_1372,In_672,In_450);
and U1373 (N_1373,In_423,In_734);
nor U1374 (N_1374,In_526,In_306);
xor U1375 (N_1375,In_355,In_416);
and U1376 (N_1376,In_687,In_646);
or U1377 (N_1377,In_358,In_127);
nand U1378 (N_1378,In_21,In_614);
xnor U1379 (N_1379,In_483,In_169);
nand U1380 (N_1380,In_620,In_250);
and U1381 (N_1381,In_459,In_734);
nor U1382 (N_1382,In_255,In_69);
nor U1383 (N_1383,In_439,In_36);
nor U1384 (N_1384,In_357,In_606);
and U1385 (N_1385,In_55,In_714);
nor U1386 (N_1386,In_75,In_293);
and U1387 (N_1387,In_423,In_303);
xnor U1388 (N_1388,In_649,In_539);
nand U1389 (N_1389,In_421,In_745);
and U1390 (N_1390,In_207,In_215);
nand U1391 (N_1391,In_562,In_331);
nor U1392 (N_1392,In_290,In_556);
nor U1393 (N_1393,In_352,In_236);
or U1394 (N_1394,In_27,In_397);
and U1395 (N_1395,In_33,In_396);
and U1396 (N_1396,In_706,In_380);
or U1397 (N_1397,In_139,In_698);
nand U1398 (N_1398,In_445,In_703);
nand U1399 (N_1399,In_248,In_115);
and U1400 (N_1400,In_516,In_1);
and U1401 (N_1401,In_186,In_664);
nand U1402 (N_1402,In_218,In_350);
or U1403 (N_1403,In_61,In_123);
nand U1404 (N_1404,In_6,In_315);
nand U1405 (N_1405,In_597,In_424);
nand U1406 (N_1406,In_567,In_121);
or U1407 (N_1407,In_524,In_459);
or U1408 (N_1408,In_433,In_574);
nor U1409 (N_1409,In_302,In_622);
nor U1410 (N_1410,In_585,In_673);
and U1411 (N_1411,In_633,In_606);
nand U1412 (N_1412,In_523,In_60);
or U1413 (N_1413,In_516,In_688);
nand U1414 (N_1414,In_380,In_296);
or U1415 (N_1415,In_656,In_328);
or U1416 (N_1416,In_259,In_682);
nor U1417 (N_1417,In_157,In_319);
nor U1418 (N_1418,In_271,In_549);
and U1419 (N_1419,In_602,In_200);
or U1420 (N_1420,In_386,In_613);
nor U1421 (N_1421,In_64,In_2);
nand U1422 (N_1422,In_460,In_395);
or U1423 (N_1423,In_125,In_733);
nand U1424 (N_1424,In_405,In_340);
or U1425 (N_1425,In_516,In_723);
or U1426 (N_1426,In_250,In_170);
nand U1427 (N_1427,In_739,In_553);
nand U1428 (N_1428,In_377,In_569);
or U1429 (N_1429,In_381,In_687);
or U1430 (N_1430,In_693,In_15);
nor U1431 (N_1431,In_504,In_125);
and U1432 (N_1432,In_294,In_349);
nor U1433 (N_1433,In_397,In_195);
or U1434 (N_1434,In_38,In_34);
nand U1435 (N_1435,In_177,In_118);
nor U1436 (N_1436,In_711,In_188);
or U1437 (N_1437,In_284,In_504);
or U1438 (N_1438,In_16,In_242);
or U1439 (N_1439,In_342,In_451);
nand U1440 (N_1440,In_629,In_561);
or U1441 (N_1441,In_270,In_207);
and U1442 (N_1442,In_659,In_561);
nor U1443 (N_1443,In_117,In_647);
nor U1444 (N_1444,In_406,In_547);
nand U1445 (N_1445,In_484,In_653);
nor U1446 (N_1446,In_164,In_641);
nor U1447 (N_1447,In_399,In_46);
or U1448 (N_1448,In_560,In_80);
nand U1449 (N_1449,In_256,In_61);
nand U1450 (N_1450,In_602,In_189);
or U1451 (N_1451,In_732,In_415);
nand U1452 (N_1452,In_627,In_27);
nand U1453 (N_1453,In_62,In_727);
or U1454 (N_1454,In_264,In_226);
nor U1455 (N_1455,In_258,In_248);
or U1456 (N_1456,In_172,In_551);
nor U1457 (N_1457,In_343,In_120);
nand U1458 (N_1458,In_591,In_78);
and U1459 (N_1459,In_113,In_542);
and U1460 (N_1460,In_11,In_309);
or U1461 (N_1461,In_382,In_37);
or U1462 (N_1462,In_399,In_405);
nand U1463 (N_1463,In_413,In_280);
and U1464 (N_1464,In_599,In_642);
nor U1465 (N_1465,In_491,In_545);
or U1466 (N_1466,In_131,In_397);
or U1467 (N_1467,In_339,In_647);
nand U1468 (N_1468,In_102,In_670);
nand U1469 (N_1469,In_619,In_484);
or U1470 (N_1470,In_72,In_608);
nor U1471 (N_1471,In_441,In_614);
or U1472 (N_1472,In_617,In_618);
and U1473 (N_1473,In_715,In_263);
and U1474 (N_1474,In_412,In_626);
nor U1475 (N_1475,In_557,In_588);
nand U1476 (N_1476,In_260,In_150);
nor U1477 (N_1477,In_670,In_139);
nand U1478 (N_1478,In_648,In_342);
and U1479 (N_1479,In_457,In_115);
nor U1480 (N_1480,In_448,In_284);
nand U1481 (N_1481,In_536,In_267);
nand U1482 (N_1482,In_417,In_61);
and U1483 (N_1483,In_30,In_222);
or U1484 (N_1484,In_533,In_390);
nor U1485 (N_1485,In_562,In_113);
nand U1486 (N_1486,In_71,In_584);
nor U1487 (N_1487,In_219,In_514);
nand U1488 (N_1488,In_432,In_593);
nor U1489 (N_1489,In_535,In_276);
nand U1490 (N_1490,In_24,In_564);
nor U1491 (N_1491,In_149,In_269);
nand U1492 (N_1492,In_150,In_640);
nor U1493 (N_1493,In_559,In_440);
nor U1494 (N_1494,In_79,In_539);
nand U1495 (N_1495,In_32,In_551);
xor U1496 (N_1496,In_159,In_157);
nand U1497 (N_1497,In_121,In_570);
nor U1498 (N_1498,In_602,In_38);
and U1499 (N_1499,In_199,In_629);
nor U1500 (N_1500,In_709,In_394);
xor U1501 (N_1501,In_250,In_97);
nor U1502 (N_1502,In_594,In_96);
and U1503 (N_1503,In_147,In_410);
nand U1504 (N_1504,In_63,In_548);
and U1505 (N_1505,In_649,In_416);
and U1506 (N_1506,In_145,In_379);
and U1507 (N_1507,In_257,In_627);
nand U1508 (N_1508,In_662,In_153);
and U1509 (N_1509,In_392,In_718);
xnor U1510 (N_1510,In_351,In_618);
and U1511 (N_1511,In_542,In_191);
xor U1512 (N_1512,In_748,In_375);
nand U1513 (N_1513,In_223,In_299);
or U1514 (N_1514,In_531,In_6);
and U1515 (N_1515,In_712,In_201);
nand U1516 (N_1516,In_357,In_540);
nor U1517 (N_1517,In_735,In_473);
or U1518 (N_1518,In_448,In_319);
and U1519 (N_1519,In_682,In_673);
and U1520 (N_1520,In_357,In_290);
nor U1521 (N_1521,In_689,In_701);
nor U1522 (N_1522,In_615,In_112);
or U1523 (N_1523,In_631,In_27);
and U1524 (N_1524,In_263,In_179);
or U1525 (N_1525,In_545,In_596);
nor U1526 (N_1526,In_100,In_579);
and U1527 (N_1527,In_392,In_194);
and U1528 (N_1528,In_571,In_464);
and U1529 (N_1529,In_261,In_736);
nor U1530 (N_1530,In_506,In_238);
or U1531 (N_1531,In_317,In_621);
nor U1532 (N_1532,In_652,In_192);
nand U1533 (N_1533,In_40,In_542);
nor U1534 (N_1534,In_352,In_69);
or U1535 (N_1535,In_344,In_469);
nor U1536 (N_1536,In_714,In_120);
and U1537 (N_1537,In_230,In_494);
and U1538 (N_1538,In_67,In_107);
nor U1539 (N_1539,In_166,In_562);
or U1540 (N_1540,In_234,In_249);
or U1541 (N_1541,In_341,In_58);
or U1542 (N_1542,In_242,In_465);
or U1543 (N_1543,In_465,In_398);
and U1544 (N_1544,In_564,In_146);
nand U1545 (N_1545,In_479,In_743);
and U1546 (N_1546,In_245,In_500);
and U1547 (N_1547,In_199,In_706);
and U1548 (N_1548,In_701,In_56);
nand U1549 (N_1549,In_735,In_503);
and U1550 (N_1550,In_13,In_314);
nor U1551 (N_1551,In_94,In_669);
or U1552 (N_1552,In_181,In_416);
nor U1553 (N_1553,In_749,In_44);
nand U1554 (N_1554,In_733,In_545);
or U1555 (N_1555,In_741,In_498);
nor U1556 (N_1556,In_394,In_112);
or U1557 (N_1557,In_198,In_100);
xnor U1558 (N_1558,In_445,In_460);
nor U1559 (N_1559,In_374,In_358);
and U1560 (N_1560,In_215,In_191);
nand U1561 (N_1561,In_24,In_238);
or U1562 (N_1562,In_585,In_316);
nand U1563 (N_1563,In_487,In_89);
and U1564 (N_1564,In_23,In_335);
and U1565 (N_1565,In_191,In_529);
nand U1566 (N_1566,In_357,In_410);
nand U1567 (N_1567,In_387,In_13);
and U1568 (N_1568,In_381,In_280);
nand U1569 (N_1569,In_224,In_360);
nor U1570 (N_1570,In_523,In_72);
or U1571 (N_1571,In_131,In_310);
or U1572 (N_1572,In_66,In_105);
or U1573 (N_1573,In_722,In_498);
and U1574 (N_1574,In_378,In_203);
and U1575 (N_1575,In_686,In_353);
nor U1576 (N_1576,In_659,In_297);
or U1577 (N_1577,In_70,In_282);
and U1578 (N_1578,In_403,In_309);
nand U1579 (N_1579,In_368,In_243);
nand U1580 (N_1580,In_477,In_111);
or U1581 (N_1581,In_274,In_0);
or U1582 (N_1582,In_110,In_143);
nand U1583 (N_1583,In_195,In_632);
and U1584 (N_1584,In_133,In_334);
nor U1585 (N_1585,In_133,In_72);
nand U1586 (N_1586,In_381,In_70);
nor U1587 (N_1587,In_60,In_105);
and U1588 (N_1588,In_599,In_702);
and U1589 (N_1589,In_592,In_13);
nand U1590 (N_1590,In_309,In_604);
or U1591 (N_1591,In_416,In_615);
nor U1592 (N_1592,In_547,In_366);
nand U1593 (N_1593,In_738,In_627);
nand U1594 (N_1594,In_420,In_300);
and U1595 (N_1595,In_520,In_397);
nor U1596 (N_1596,In_717,In_2);
nor U1597 (N_1597,In_122,In_80);
nor U1598 (N_1598,In_365,In_381);
and U1599 (N_1599,In_702,In_202);
nand U1600 (N_1600,In_490,In_153);
and U1601 (N_1601,In_656,In_513);
nor U1602 (N_1602,In_304,In_234);
nor U1603 (N_1603,In_535,In_527);
or U1604 (N_1604,In_35,In_701);
nor U1605 (N_1605,In_604,In_121);
nor U1606 (N_1606,In_552,In_537);
nor U1607 (N_1607,In_366,In_513);
nand U1608 (N_1608,In_277,In_280);
or U1609 (N_1609,In_330,In_730);
nor U1610 (N_1610,In_263,In_441);
nor U1611 (N_1611,In_308,In_604);
or U1612 (N_1612,In_42,In_314);
nand U1613 (N_1613,In_258,In_539);
nor U1614 (N_1614,In_356,In_720);
nand U1615 (N_1615,In_252,In_447);
or U1616 (N_1616,In_83,In_701);
nand U1617 (N_1617,In_652,In_370);
and U1618 (N_1618,In_303,In_459);
or U1619 (N_1619,In_298,In_293);
and U1620 (N_1620,In_341,In_30);
nand U1621 (N_1621,In_640,In_582);
nand U1622 (N_1622,In_511,In_629);
and U1623 (N_1623,In_273,In_469);
and U1624 (N_1624,In_229,In_540);
and U1625 (N_1625,In_575,In_613);
and U1626 (N_1626,In_555,In_124);
nand U1627 (N_1627,In_668,In_621);
nand U1628 (N_1628,In_445,In_214);
nor U1629 (N_1629,In_637,In_591);
nor U1630 (N_1630,In_464,In_434);
or U1631 (N_1631,In_156,In_644);
nand U1632 (N_1632,In_536,In_67);
or U1633 (N_1633,In_497,In_304);
or U1634 (N_1634,In_548,In_615);
nand U1635 (N_1635,In_117,In_72);
nor U1636 (N_1636,In_407,In_597);
nand U1637 (N_1637,In_625,In_743);
and U1638 (N_1638,In_173,In_500);
nor U1639 (N_1639,In_294,In_713);
nor U1640 (N_1640,In_316,In_310);
and U1641 (N_1641,In_295,In_508);
nand U1642 (N_1642,In_357,In_226);
or U1643 (N_1643,In_1,In_748);
nand U1644 (N_1644,In_64,In_528);
nand U1645 (N_1645,In_453,In_285);
nor U1646 (N_1646,In_441,In_282);
nor U1647 (N_1647,In_599,In_541);
and U1648 (N_1648,In_36,In_212);
nor U1649 (N_1649,In_345,In_78);
or U1650 (N_1650,In_318,In_734);
xor U1651 (N_1651,In_233,In_589);
or U1652 (N_1652,In_417,In_657);
nand U1653 (N_1653,In_508,In_109);
nand U1654 (N_1654,In_713,In_611);
nand U1655 (N_1655,In_533,In_175);
nor U1656 (N_1656,In_252,In_227);
nor U1657 (N_1657,In_56,In_575);
nand U1658 (N_1658,In_226,In_114);
nor U1659 (N_1659,In_272,In_333);
and U1660 (N_1660,In_363,In_295);
nand U1661 (N_1661,In_679,In_544);
nand U1662 (N_1662,In_329,In_662);
and U1663 (N_1663,In_196,In_72);
xor U1664 (N_1664,In_498,In_321);
or U1665 (N_1665,In_573,In_376);
and U1666 (N_1666,In_312,In_65);
or U1667 (N_1667,In_400,In_252);
nor U1668 (N_1668,In_336,In_554);
and U1669 (N_1669,In_638,In_387);
or U1670 (N_1670,In_708,In_367);
nand U1671 (N_1671,In_78,In_559);
nor U1672 (N_1672,In_572,In_256);
or U1673 (N_1673,In_155,In_336);
nor U1674 (N_1674,In_457,In_556);
or U1675 (N_1675,In_534,In_724);
nor U1676 (N_1676,In_270,In_197);
nor U1677 (N_1677,In_589,In_395);
and U1678 (N_1678,In_191,In_282);
nand U1679 (N_1679,In_174,In_19);
or U1680 (N_1680,In_360,In_517);
nand U1681 (N_1681,In_134,In_40);
and U1682 (N_1682,In_732,In_496);
nand U1683 (N_1683,In_139,In_503);
nand U1684 (N_1684,In_461,In_79);
nor U1685 (N_1685,In_366,In_466);
and U1686 (N_1686,In_277,In_664);
nor U1687 (N_1687,In_235,In_243);
nor U1688 (N_1688,In_580,In_561);
nor U1689 (N_1689,In_527,In_83);
nand U1690 (N_1690,In_294,In_252);
and U1691 (N_1691,In_468,In_37);
and U1692 (N_1692,In_443,In_722);
and U1693 (N_1693,In_230,In_400);
or U1694 (N_1694,In_446,In_223);
or U1695 (N_1695,In_79,In_673);
nand U1696 (N_1696,In_8,In_123);
nor U1697 (N_1697,In_583,In_377);
nand U1698 (N_1698,In_470,In_302);
and U1699 (N_1699,In_425,In_45);
or U1700 (N_1700,In_564,In_683);
and U1701 (N_1701,In_680,In_382);
nor U1702 (N_1702,In_716,In_72);
xnor U1703 (N_1703,In_526,In_146);
and U1704 (N_1704,In_715,In_127);
and U1705 (N_1705,In_439,In_24);
nor U1706 (N_1706,In_205,In_417);
and U1707 (N_1707,In_706,In_574);
or U1708 (N_1708,In_364,In_443);
nand U1709 (N_1709,In_720,In_72);
or U1710 (N_1710,In_595,In_28);
nor U1711 (N_1711,In_149,In_609);
nand U1712 (N_1712,In_515,In_153);
or U1713 (N_1713,In_641,In_204);
or U1714 (N_1714,In_421,In_352);
nand U1715 (N_1715,In_732,In_596);
nor U1716 (N_1716,In_16,In_489);
and U1717 (N_1717,In_91,In_545);
and U1718 (N_1718,In_730,In_580);
nor U1719 (N_1719,In_143,In_202);
nand U1720 (N_1720,In_375,In_493);
or U1721 (N_1721,In_207,In_256);
nand U1722 (N_1722,In_436,In_379);
or U1723 (N_1723,In_202,In_645);
and U1724 (N_1724,In_214,In_619);
nand U1725 (N_1725,In_541,In_82);
nor U1726 (N_1726,In_374,In_586);
and U1727 (N_1727,In_638,In_462);
and U1728 (N_1728,In_56,In_689);
or U1729 (N_1729,In_736,In_9);
nor U1730 (N_1730,In_359,In_356);
or U1731 (N_1731,In_383,In_420);
and U1732 (N_1732,In_83,In_611);
nor U1733 (N_1733,In_162,In_235);
or U1734 (N_1734,In_87,In_275);
nand U1735 (N_1735,In_305,In_285);
or U1736 (N_1736,In_6,In_427);
and U1737 (N_1737,In_238,In_397);
nand U1738 (N_1738,In_540,In_84);
nor U1739 (N_1739,In_495,In_716);
nor U1740 (N_1740,In_72,In_621);
or U1741 (N_1741,In_330,In_181);
and U1742 (N_1742,In_89,In_387);
or U1743 (N_1743,In_128,In_659);
nand U1744 (N_1744,In_479,In_719);
or U1745 (N_1745,In_519,In_620);
and U1746 (N_1746,In_671,In_86);
nand U1747 (N_1747,In_206,In_714);
or U1748 (N_1748,In_343,In_212);
or U1749 (N_1749,In_290,In_689);
or U1750 (N_1750,In_53,In_503);
and U1751 (N_1751,In_566,In_6);
nand U1752 (N_1752,In_46,In_371);
and U1753 (N_1753,In_630,In_190);
or U1754 (N_1754,In_100,In_320);
or U1755 (N_1755,In_152,In_52);
nor U1756 (N_1756,In_124,In_322);
or U1757 (N_1757,In_153,In_67);
nor U1758 (N_1758,In_303,In_301);
or U1759 (N_1759,In_304,In_467);
or U1760 (N_1760,In_30,In_510);
and U1761 (N_1761,In_286,In_340);
nand U1762 (N_1762,In_40,In_261);
nor U1763 (N_1763,In_191,In_702);
nor U1764 (N_1764,In_499,In_458);
nand U1765 (N_1765,In_341,In_297);
or U1766 (N_1766,In_622,In_36);
or U1767 (N_1767,In_268,In_611);
nor U1768 (N_1768,In_92,In_124);
and U1769 (N_1769,In_17,In_609);
nor U1770 (N_1770,In_581,In_88);
nor U1771 (N_1771,In_671,In_513);
and U1772 (N_1772,In_733,In_227);
or U1773 (N_1773,In_654,In_540);
or U1774 (N_1774,In_653,In_283);
or U1775 (N_1775,In_309,In_328);
nor U1776 (N_1776,In_623,In_579);
or U1777 (N_1777,In_153,In_141);
and U1778 (N_1778,In_431,In_122);
and U1779 (N_1779,In_1,In_212);
and U1780 (N_1780,In_261,In_179);
nand U1781 (N_1781,In_124,In_471);
or U1782 (N_1782,In_452,In_607);
and U1783 (N_1783,In_452,In_355);
and U1784 (N_1784,In_301,In_374);
or U1785 (N_1785,In_323,In_114);
nor U1786 (N_1786,In_646,In_355);
nand U1787 (N_1787,In_388,In_40);
and U1788 (N_1788,In_418,In_468);
or U1789 (N_1789,In_21,In_657);
nor U1790 (N_1790,In_595,In_611);
nand U1791 (N_1791,In_19,In_93);
and U1792 (N_1792,In_542,In_104);
and U1793 (N_1793,In_724,In_715);
nand U1794 (N_1794,In_211,In_703);
nand U1795 (N_1795,In_504,In_107);
nand U1796 (N_1796,In_575,In_128);
or U1797 (N_1797,In_592,In_731);
and U1798 (N_1798,In_647,In_284);
nor U1799 (N_1799,In_76,In_365);
or U1800 (N_1800,In_679,In_270);
nor U1801 (N_1801,In_399,In_565);
nor U1802 (N_1802,In_611,In_637);
or U1803 (N_1803,In_474,In_181);
and U1804 (N_1804,In_116,In_84);
nor U1805 (N_1805,In_286,In_587);
nand U1806 (N_1806,In_27,In_38);
nor U1807 (N_1807,In_209,In_375);
or U1808 (N_1808,In_144,In_130);
nand U1809 (N_1809,In_522,In_591);
and U1810 (N_1810,In_663,In_506);
nand U1811 (N_1811,In_116,In_554);
or U1812 (N_1812,In_712,In_368);
nand U1813 (N_1813,In_35,In_594);
nor U1814 (N_1814,In_425,In_327);
and U1815 (N_1815,In_268,In_645);
or U1816 (N_1816,In_411,In_665);
nand U1817 (N_1817,In_163,In_386);
and U1818 (N_1818,In_659,In_70);
nand U1819 (N_1819,In_214,In_229);
nor U1820 (N_1820,In_135,In_610);
or U1821 (N_1821,In_451,In_684);
nor U1822 (N_1822,In_592,In_21);
or U1823 (N_1823,In_377,In_724);
nor U1824 (N_1824,In_224,In_56);
or U1825 (N_1825,In_419,In_324);
or U1826 (N_1826,In_494,In_550);
nor U1827 (N_1827,In_6,In_203);
nor U1828 (N_1828,In_153,In_532);
nor U1829 (N_1829,In_88,In_252);
nand U1830 (N_1830,In_314,In_345);
or U1831 (N_1831,In_469,In_543);
xnor U1832 (N_1832,In_528,In_241);
nand U1833 (N_1833,In_42,In_642);
nand U1834 (N_1834,In_640,In_355);
and U1835 (N_1835,In_531,In_411);
and U1836 (N_1836,In_234,In_127);
and U1837 (N_1837,In_678,In_64);
nor U1838 (N_1838,In_378,In_214);
nor U1839 (N_1839,In_549,In_623);
nor U1840 (N_1840,In_577,In_505);
and U1841 (N_1841,In_260,In_252);
or U1842 (N_1842,In_393,In_53);
and U1843 (N_1843,In_506,In_130);
nor U1844 (N_1844,In_446,In_238);
or U1845 (N_1845,In_28,In_353);
or U1846 (N_1846,In_65,In_332);
and U1847 (N_1847,In_735,In_626);
and U1848 (N_1848,In_36,In_458);
and U1849 (N_1849,In_362,In_339);
and U1850 (N_1850,In_16,In_354);
nand U1851 (N_1851,In_660,In_51);
or U1852 (N_1852,In_290,In_36);
or U1853 (N_1853,In_526,In_595);
or U1854 (N_1854,In_279,In_598);
and U1855 (N_1855,In_667,In_675);
and U1856 (N_1856,In_38,In_226);
and U1857 (N_1857,In_629,In_129);
nand U1858 (N_1858,In_372,In_712);
nor U1859 (N_1859,In_460,In_687);
nor U1860 (N_1860,In_66,In_186);
and U1861 (N_1861,In_261,In_32);
and U1862 (N_1862,In_384,In_464);
and U1863 (N_1863,In_439,In_313);
or U1864 (N_1864,In_466,In_469);
or U1865 (N_1865,In_686,In_528);
or U1866 (N_1866,In_252,In_470);
and U1867 (N_1867,In_359,In_16);
nor U1868 (N_1868,In_334,In_694);
nand U1869 (N_1869,In_371,In_377);
or U1870 (N_1870,In_618,In_537);
or U1871 (N_1871,In_114,In_46);
and U1872 (N_1872,In_643,In_433);
nor U1873 (N_1873,In_299,In_65);
nand U1874 (N_1874,In_508,In_181);
nand U1875 (N_1875,In_0,In_295);
or U1876 (N_1876,In_214,In_213);
nor U1877 (N_1877,In_719,In_476);
nor U1878 (N_1878,In_59,In_398);
nor U1879 (N_1879,In_738,In_406);
and U1880 (N_1880,In_568,In_33);
nor U1881 (N_1881,In_175,In_29);
or U1882 (N_1882,In_169,In_376);
nand U1883 (N_1883,In_255,In_110);
and U1884 (N_1884,In_137,In_314);
nand U1885 (N_1885,In_631,In_319);
nor U1886 (N_1886,In_684,In_725);
or U1887 (N_1887,In_644,In_481);
nand U1888 (N_1888,In_362,In_77);
and U1889 (N_1889,In_522,In_604);
and U1890 (N_1890,In_436,In_701);
or U1891 (N_1891,In_563,In_601);
or U1892 (N_1892,In_315,In_647);
and U1893 (N_1893,In_526,In_144);
or U1894 (N_1894,In_459,In_441);
nand U1895 (N_1895,In_341,In_569);
nor U1896 (N_1896,In_477,In_309);
and U1897 (N_1897,In_722,In_692);
nor U1898 (N_1898,In_566,In_162);
nor U1899 (N_1899,In_659,In_360);
and U1900 (N_1900,In_427,In_122);
or U1901 (N_1901,In_188,In_553);
nand U1902 (N_1902,In_300,In_144);
xnor U1903 (N_1903,In_323,In_327);
nor U1904 (N_1904,In_147,In_222);
or U1905 (N_1905,In_678,In_359);
nor U1906 (N_1906,In_391,In_480);
or U1907 (N_1907,In_277,In_128);
and U1908 (N_1908,In_127,In_540);
and U1909 (N_1909,In_74,In_474);
nor U1910 (N_1910,In_546,In_13);
and U1911 (N_1911,In_576,In_251);
and U1912 (N_1912,In_656,In_195);
nor U1913 (N_1913,In_295,In_49);
and U1914 (N_1914,In_554,In_427);
nand U1915 (N_1915,In_108,In_431);
or U1916 (N_1916,In_6,In_429);
nor U1917 (N_1917,In_610,In_343);
nand U1918 (N_1918,In_584,In_188);
nand U1919 (N_1919,In_559,In_519);
and U1920 (N_1920,In_616,In_515);
nor U1921 (N_1921,In_213,In_361);
or U1922 (N_1922,In_389,In_187);
and U1923 (N_1923,In_329,In_19);
or U1924 (N_1924,In_492,In_725);
nor U1925 (N_1925,In_78,In_396);
nor U1926 (N_1926,In_358,In_503);
or U1927 (N_1927,In_579,In_229);
nand U1928 (N_1928,In_380,In_196);
or U1929 (N_1929,In_316,In_599);
nor U1930 (N_1930,In_467,In_276);
nor U1931 (N_1931,In_294,In_727);
and U1932 (N_1932,In_568,In_20);
nand U1933 (N_1933,In_371,In_617);
or U1934 (N_1934,In_354,In_121);
and U1935 (N_1935,In_13,In_702);
or U1936 (N_1936,In_279,In_104);
nor U1937 (N_1937,In_449,In_749);
nand U1938 (N_1938,In_525,In_107);
nand U1939 (N_1939,In_599,In_418);
and U1940 (N_1940,In_573,In_286);
nor U1941 (N_1941,In_102,In_280);
nand U1942 (N_1942,In_312,In_302);
nor U1943 (N_1943,In_22,In_49);
and U1944 (N_1944,In_283,In_87);
or U1945 (N_1945,In_209,In_264);
nand U1946 (N_1946,In_329,In_433);
or U1947 (N_1947,In_41,In_693);
nand U1948 (N_1948,In_645,In_225);
nand U1949 (N_1949,In_347,In_275);
nor U1950 (N_1950,In_51,In_288);
nor U1951 (N_1951,In_258,In_559);
nand U1952 (N_1952,In_138,In_392);
and U1953 (N_1953,In_654,In_343);
nand U1954 (N_1954,In_55,In_565);
or U1955 (N_1955,In_74,In_316);
nor U1956 (N_1956,In_152,In_81);
and U1957 (N_1957,In_597,In_321);
nand U1958 (N_1958,In_273,In_81);
nor U1959 (N_1959,In_158,In_256);
and U1960 (N_1960,In_341,In_636);
nand U1961 (N_1961,In_479,In_380);
nor U1962 (N_1962,In_737,In_331);
nand U1963 (N_1963,In_144,In_569);
and U1964 (N_1964,In_174,In_196);
nand U1965 (N_1965,In_573,In_367);
nand U1966 (N_1966,In_89,In_308);
nand U1967 (N_1967,In_184,In_741);
nand U1968 (N_1968,In_685,In_376);
nor U1969 (N_1969,In_37,In_721);
and U1970 (N_1970,In_237,In_520);
nand U1971 (N_1971,In_519,In_230);
nor U1972 (N_1972,In_549,In_475);
nand U1973 (N_1973,In_407,In_677);
nor U1974 (N_1974,In_368,In_585);
or U1975 (N_1975,In_91,In_82);
and U1976 (N_1976,In_201,In_143);
nor U1977 (N_1977,In_734,In_552);
nor U1978 (N_1978,In_438,In_395);
and U1979 (N_1979,In_564,In_202);
nand U1980 (N_1980,In_232,In_403);
and U1981 (N_1981,In_489,In_268);
nand U1982 (N_1982,In_569,In_401);
or U1983 (N_1983,In_129,In_157);
or U1984 (N_1984,In_57,In_634);
nand U1985 (N_1985,In_453,In_190);
or U1986 (N_1986,In_299,In_546);
or U1987 (N_1987,In_80,In_133);
and U1988 (N_1988,In_254,In_198);
and U1989 (N_1989,In_635,In_318);
and U1990 (N_1990,In_330,In_120);
nor U1991 (N_1991,In_197,In_89);
and U1992 (N_1992,In_156,In_310);
nor U1993 (N_1993,In_305,In_512);
and U1994 (N_1994,In_339,In_297);
nor U1995 (N_1995,In_388,In_327);
or U1996 (N_1996,In_504,In_432);
nand U1997 (N_1997,In_145,In_722);
nand U1998 (N_1998,In_648,In_676);
and U1999 (N_1999,In_445,In_89);
nor U2000 (N_2000,In_644,In_527);
nor U2001 (N_2001,In_197,In_264);
nand U2002 (N_2002,In_94,In_399);
and U2003 (N_2003,In_653,In_677);
nand U2004 (N_2004,In_149,In_313);
nand U2005 (N_2005,In_738,In_402);
or U2006 (N_2006,In_479,In_339);
and U2007 (N_2007,In_101,In_432);
nor U2008 (N_2008,In_456,In_549);
nand U2009 (N_2009,In_69,In_522);
or U2010 (N_2010,In_272,In_370);
or U2011 (N_2011,In_51,In_661);
and U2012 (N_2012,In_28,In_290);
nor U2013 (N_2013,In_292,In_273);
and U2014 (N_2014,In_65,In_274);
and U2015 (N_2015,In_184,In_730);
nand U2016 (N_2016,In_142,In_522);
nand U2017 (N_2017,In_253,In_538);
nor U2018 (N_2018,In_170,In_584);
nand U2019 (N_2019,In_439,In_90);
nor U2020 (N_2020,In_156,In_205);
and U2021 (N_2021,In_441,In_534);
or U2022 (N_2022,In_496,In_551);
and U2023 (N_2023,In_521,In_444);
nand U2024 (N_2024,In_340,In_436);
nor U2025 (N_2025,In_341,In_310);
nor U2026 (N_2026,In_398,In_115);
nand U2027 (N_2027,In_197,In_117);
nand U2028 (N_2028,In_2,In_449);
nand U2029 (N_2029,In_84,In_78);
nand U2030 (N_2030,In_130,In_594);
nand U2031 (N_2031,In_132,In_676);
and U2032 (N_2032,In_710,In_553);
xnor U2033 (N_2033,In_339,In_447);
nand U2034 (N_2034,In_165,In_661);
nand U2035 (N_2035,In_291,In_92);
and U2036 (N_2036,In_544,In_608);
nor U2037 (N_2037,In_536,In_400);
nor U2038 (N_2038,In_121,In_543);
xnor U2039 (N_2039,In_395,In_57);
nand U2040 (N_2040,In_497,In_445);
or U2041 (N_2041,In_537,In_324);
nand U2042 (N_2042,In_404,In_267);
nand U2043 (N_2043,In_79,In_683);
and U2044 (N_2044,In_604,In_614);
nand U2045 (N_2045,In_319,In_725);
or U2046 (N_2046,In_493,In_708);
nor U2047 (N_2047,In_91,In_405);
or U2048 (N_2048,In_595,In_316);
and U2049 (N_2049,In_145,In_98);
and U2050 (N_2050,In_13,In_222);
nand U2051 (N_2051,In_725,In_307);
and U2052 (N_2052,In_287,In_716);
or U2053 (N_2053,In_375,In_165);
nor U2054 (N_2054,In_474,In_15);
nor U2055 (N_2055,In_573,In_543);
nor U2056 (N_2056,In_606,In_274);
nand U2057 (N_2057,In_92,In_643);
or U2058 (N_2058,In_411,In_564);
and U2059 (N_2059,In_488,In_388);
nand U2060 (N_2060,In_170,In_442);
nor U2061 (N_2061,In_36,In_468);
xor U2062 (N_2062,In_370,In_441);
or U2063 (N_2063,In_14,In_464);
nand U2064 (N_2064,In_340,In_693);
nand U2065 (N_2065,In_55,In_302);
nor U2066 (N_2066,In_28,In_240);
and U2067 (N_2067,In_123,In_643);
nand U2068 (N_2068,In_470,In_93);
nor U2069 (N_2069,In_174,In_623);
and U2070 (N_2070,In_470,In_493);
or U2071 (N_2071,In_396,In_269);
and U2072 (N_2072,In_667,In_254);
and U2073 (N_2073,In_53,In_422);
nand U2074 (N_2074,In_178,In_24);
or U2075 (N_2075,In_104,In_651);
nor U2076 (N_2076,In_584,In_548);
nor U2077 (N_2077,In_718,In_55);
nor U2078 (N_2078,In_455,In_346);
nand U2079 (N_2079,In_0,In_361);
or U2080 (N_2080,In_319,In_616);
or U2081 (N_2081,In_377,In_191);
nor U2082 (N_2082,In_570,In_471);
or U2083 (N_2083,In_427,In_168);
and U2084 (N_2084,In_485,In_488);
or U2085 (N_2085,In_78,In_272);
nand U2086 (N_2086,In_278,In_617);
or U2087 (N_2087,In_362,In_166);
and U2088 (N_2088,In_208,In_663);
nand U2089 (N_2089,In_632,In_212);
or U2090 (N_2090,In_4,In_317);
or U2091 (N_2091,In_73,In_108);
and U2092 (N_2092,In_51,In_336);
or U2093 (N_2093,In_267,In_258);
or U2094 (N_2094,In_295,In_526);
nor U2095 (N_2095,In_130,In_29);
nand U2096 (N_2096,In_585,In_602);
nand U2097 (N_2097,In_24,In_142);
nor U2098 (N_2098,In_190,In_289);
or U2099 (N_2099,In_263,In_236);
and U2100 (N_2100,In_104,In_526);
or U2101 (N_2101,In_182,In_99);
or U2102 (N_2102,In_216,In_575);
or U2103 (N_2103,In_334,In_118);
nand U2104 (N_2104,In_627,In_68);
or U2105 (N_2105,In_725,In_544);
and U2106 (N_2106,In_493,In_243);
nand U2107 (N_2107,In_133,In_108);
nor U2108 (N_2108,In_284,In_186);
nand U2109 (N_2109,In_205,In_617);
and U2110 (N_2110,In_111,In_314);
or U2111 (N_2111,In_365,In_718);
nor U2112 (N_2112,In_553,In_114);
nor U2113 (N_2113,In_517,In_251);
and U2114 (N_2114,In_616,In_746);
nor U2115 (N_2115,In_81,In_55);
or U2116 (N_2116,In_713,In_82);
and U2117 (N_2117,In_689,In_742);
or U2118 (N_2118,In_730,In_734);
or U2119 (N_2119,In_31,In_73);
nand U2120 (N_2120,In_97,In_222);
and U2121 (N_2121,In_699,In_475);
or U2122 (N_2122,In_50,In_705);
or U2123 (N_2123,In_653,In_474);
and U2124 (N_2124,In_407,In_126);
nor U2125 (N_2125,In_375,In_455);
nor U2126 (N_2126,In_86,In_206);
nand U2127 (N_2127,In_265,In_528);
and U2128 (N_2128,In_225,In_547);
or U2129 (N_2129,In_733,In_237);
and U2130 (N_2130,In_651,In_522);
nor U2131 (N_2131,In_748,In_123);
nand U2132 (N_2132,In_413,In_232);
nor U2133 (N_2133,In_451,In_124);
or U2134 (N_2134,In_735,In_16);
nand U2135 (N_2135,In_252,In_572);
nor U2136 (N_2136,In_573,In_529);
nand U2137 (N_2137,In_272,In_193);
nor U2138 (N_2138,In_512,In_258);
or U2139 (N_2139,In_301,In_207);
nor U2140 (N_2140,In_569,In_600);
nor U2141 (N_2141,In_635,In_81);
or U2142 (N_2142,In_677,In_116);
or U2143 (N_2143,In_42,In_536);
nor U2144 (N_2144,In_445,In_190);
and U2145 (N_2145,In_296,In_237);
or U2146 (N_2146,In_368,In_682);
nand U2147 (N_2147,In_116,In_206);
nand U2148 (N_2148,In_113,In_743);
or U2149 (N_2149,In_517,In_298);
nand U2150 (N_2150,In_429,In_56);
nand U2151 (N_2151,In_2,In_419);
and U2152 (N_2152,In_147,In_680);
and U2153 (N_2153,In_561,In_2);
and U2154 (N_2154,In_290,In_563);
or U2155 (N_2155,In_521,In_255);
or U2156 (N_2156,In_335,In_502);
and U2157 (N_2157,In_440,In_324);
nand U2158 (N_2158,In_324,In_424);
and U2159 (N_2159,In_16,In_22);
nand U2160 (N_2160,In_57,In_430);
nor U2161 (N_2161,In_422,In_84);
or U2162 (N_2162,In_471,In_683);
nor U2163 (N_2163,In_250,In_524);
or U2164 (N_2164,In_313,In_592);
nor U2165 (N_2165,In_282,In_130);
and U2166 (N_2166,In_238,In_159);
xor U2167 (N_2167,In_91,In_211);
or U2168 (N_2168,In_205,In_89);
nor U2169 (N_2169,In_24,In_283);
or U2170 (N_2170,In_259,In_597);
and U2171 (N_2171,In_111,In_169);
nand U2172 (N_2172,In_397,In_583);
nand U2173 (N_2173,In_667,In_370);
nand U2174 (N_2174,In_407,In_709);
nand U2175 (N_2175,In_83,In_19);
nor U2176 (N_2176,In_661,In_436);
nor U2177 (N_2177,In_289,In_605);
or U2178 (N_2178,In_296,In_1);
nor U2179 (N_2179,In_313,In_401);
or U2180 (N_2180,In_390,In_557);
or U2181 (N_2181,In_4,In_579);
nand U2182 (N_2182,In_278,In_154);
or U2183 (N_2183,In_207,In_118);
nand U2184 (N_2184,In_151,In_504);
nand U2185 (N_2185,In_228,In_234);
nor U2186 (N_2186,In_190,In_156);
or U2187 (N_2187,In_169,In_235);
or U2188 (N_2188,In_524,In_582);
nor U2189 (N_2189,In_669,In_363);
nand U2190 (N_2190,In_605,In_213);
and U2191 (N_2191,In_307,In_166);
nand U2192 (N_2192,In_447,In_261);
nand U2193 (N_2193,In_227,In_680);
or U2194 (N_2194,In_704,In_610);
or U2195 (N_2195,In_749,In_467);
or U2196 (N_2196,In_299,In_191);
or U2197 (N_2197,In_396,In_533);
and U2198 (N_2198,In_580,In_407);
xnor U2199 (N_2199,In_622,In_130);
and U2200 (N_2200,In_321,In_574);
nand U2201 (N_2201,In_4,In_375);
nor U2202 (N_2202,In_278,In_602);
nor U2203 (N_2203,In_338,In_361);
nand U2204 (N_2204,In_195,In_391);
nand U2205 (N_2205,In_491,In_378);
nand U2206 (N_2206,In_67,In_663);
nor U2207 (N_2207,In_166,In_36);
nand U2208 (N_2208,In_144,In_274);
and U2209 (N_2209,In_733,In_587);
nor U2210 (N_2210,In_555,In_686);
and U2211 (N_2211,In_473,In_144);
and U2212 (N_2212,In_447,In_23);
nand U2213 (N_2213,In_216,In_5);
nor U2214 (N_2214,In_520,In_622);
or U2215 (N_2215,In_34,In_492);
nor U2216 (N_2216,In_514,In_535);
nand U2217 (N_2217,In_530,In_585);
nor U2218 (N_2218,In_381,In_429);
and U2219 (N_2219,In_307,In_227);
nand U2220 (N_2220,In_726,In_315);
or U2221 (N_2221,In_741,In_133);
nand U2222 (N_2222,In_8,In_690);
and U2223 (N_2223,In_29,In_338);
nand U2224 (N_2224,In_351,In_402);
nand U2225 (N_2225,In_432,In_368);
and U2226 (N_2226,In_536,In_639);
and U2227 (N_2227,In_680,In_584);
nor U2228 (N_2228,In_491,In_722);
nand U2229 (N_2229,In_494,In_513);
nor U2230 (N_2230,In_9,In_118);
nor U2231 (N_2231,In_606,In_240);
nand U2232 (N_2232,In_327,In_501);
or U2233 (N_2233,In_316,In_76);
nand U2234 (N_2234,In_603,In_104);
nor U2235 (N_2235,In_51,In_89);
or U2236 (N_2236,In_28,In_549);
and U2237 (N_2237,In_547,In_126);
nor U2238 (N_2238,In_72,In_606);
and U2239 (N_2239,In_197,In_492);
or U2240 (N_2240,In_49,In_627);
or U2241 (N_2241,In_141,In_327);
and U2242 (N_2242,In_25,In_501);
or U2243 (N_2243,In_191,In_9);
nor U2244 (N_2244,In_413,In_553);
and U2245 (N_2245,In_454,In_542);
and U2246 (N_2246,In_664,In_423);
and U2247 (N_2247,In_610,In_358);
nor U2248 (N_2248,In_408,In_635);
nor U2249 (N_2249,In_545,In_14);
nand U2250 (N_2250,In_1,In_684);
nand U2251 (N_2251,In_141,In_45);
nor U2252 (N_2252,In_512,In_225);
nor U2253 (N_2253,In_623,In_269);
and U2254 (N_2254,In_248,In_82);
and U2255 (N_2255,In_558,In_687);
and U2256 (N_2256,In_145,In_472);
nor U2257 (N_2257,In_159,In_227);
nand U2258 (N_2258,In_676,In_459);
and U2259 (N_2259,In_260,In_67);
nor U2260 (N_2260,In_336,In_233);
or U2261 (N_2261,In_361,In_290);
nor U2262 (N_2262,In_713,In_433);
or U2263 (N_2263,In_526,In_215);
and U2264 (N_2264,In_355,In_690);
and U2265 (N_2265,In_547,In_730);
or U2266 (N_2266,In_308,In_616);
or U2267 (N_2267,In_524,In_738);
nor U2268 (N_2268,In_138,In_659);
nor U2269 (N_2269,In_255,In_9);
nor U2270 (N_2270,In_727,In_225);
nor U2271 (N_2271,In_671,In_202);
and U2272 (N_2272,In_373,In_6);
and U2273 (N_2273,In_688,In_35);
nand U2274 (N_2274,In_735,In_526);
and U2275 (N_2275,In_77,In_561);
or U2276 (N_2276,In_149,In_718);
or U2277 (N_2277,In_380,In_537);
nand U2278 (N_2278,In_687,In_746);
or U2279 (N_2279,In_131,In_644);
or U2280 (N_2280,In_20,In_143);
and U2281 (N_2281,In_415,In_222);
xor U2282 (N_2282,In_353,In_407);
or U2283 (N_2283,In_611,In_341);
and U2284 (N_2284,In_703,In_60);
and U2285 (N_2285,In_273,In_137);
or U2286 (N_2286,In_527,In_11);
nand U2287 (N_2287,In_714,In_669);
nor U2288 (N_2288,In_56,In_693);
nor U2289 (N_2289,In_127,In_196);
and U2290 (N_2290,In_716,In_282);
or U2291 (N_2291,In_676,In_391);
xor U2292 (N_2292,In_36,In_601);
and U2293 (N_2293,In_434,In_215);
or U2294 (N_2294,In_704,In_599);
xnor U2295 (N_2295,In_192,In_549);
nand U2296 (N_2296,In_500,In_98);
nor U2297 (N_2297,In_246,In_344);
nand U2298 (N_2298,In_480,In_282);
nor U2299 (N_2299,In_699,In_8);
or U2300 (N_2300,In_560,In_267);
and U2301 (N_2301,In_356,In_53);
nor U2302 (N_2302,In_153,In_432);
nand U2303 (N_2303,In_404,In_308);
and U2304 (N_2304,In_425,In_144);
nand U2305 (N_2305,In_395,In_309);
or U2306 (N_2306,In_608,In_184);
or U2307 (N_2307,In_564,In_664);
or U2308 (N_2308,In_330,In_361);
and U2309 (N_2309,In_29,In_522);
and U2310 (N_2310,In_513,In_135);
nand U2311 (N_2311,In_644,In_183);
nor U2312 (N_2312,In_562,In_229);
nor U2313 (N_2313,In_414,In_689);
and U2314 (N_2314,In_517,In_450);
or U2315 (N_2315,In_312,In_611);
nand U2316 (N_2316,In_143,In_247);
and U2317 (N_2317,In_366,In_550);
nor U2318 (N_2318,In_731,In_29);
nor U2319 (N_2319,In_193,In_266);
or U2320 (N_2320,In_485,In_156);
and U2321 (N_2321,In_220,In_152);
or U2322 (N_2322,In_169,In_394);
and U2323 (N_2323,In_155,In_237);
and U2324 (N_2324,In_578,In_295);
nor U2325 (N_2325,In_344,In_554);
or U2326 (N_2326,In_493,In_161);
nor U2327 (N_2327,In_661,In_710);
and U2328 (N_2328,In_383,In_492);
nand U2329 (N_2329,In_10,In_358);
or U2330 (N_2330,In_453,In_204);
nand U2331 (N_2331,In_532,In_688);
and U2332 (N_2332,In_14,In_745);
or U2333 (N_2333,In_254,In_360);
or U2334 (N_2334,In_694,In_271);
nand U2335 (N_2335,In_163,In_735);
nor U2336 (N_2336,In_235,In_41);
nor U2337 (N_2337,In_175,In_73);
and U2338 (N_2338,In_720,In_424);
nand U2339 (N_2339,In_476,In_362);
nand U2340 (N_2340,In_291,In_119);
or U2341 (N_2341,In_686,In_333);
nor U2342 (N_2342,In_568,In_195);
and U2343 (N_2343,In_202,In_118);
nor U2344 (N_2344,In_17,In_473);
nor U2345 (N_2345,In_520,In_594);
or U2346 (N_2346,In_375,In_174);
and U2347 (N_2347,In_650,In_220);
and U2348 (N_2348,In_239,In_218);
or U2349 (N_2349,In_180,In_545);
nor U2350 (N_2350,In_222,In_9);
and U2351 (N_2351,In_462,In_291);
and U2352 (N_2352,In_702,In_326);
and U2353 (N_2353,In_64,In_536);
nand U2354 (N_2354,In_536,In_280);
or U2355 (N_2355,In_311,In_104);
and U2356 (N_2356,In_218,In_161);
or U2357 (N_2357,In_621,In_457);
nor U2358 (N_2358,In_188,In_447);
and U2359 (N_2359,In_0,In_585);
or U2360 (N_2360,In_493,In_422);
or U2361 (N_2361,In_386,In_459);
and U2362 (N_2362,In_379,In_113);
nor U2363 (N_2363,In_288,In_619);
or U2364 (N_2364,In_39,In_696);
and U2365 (N_2365,In_308,In_274);
and U2366 (N_2366,In_449,In_689);
nor U2367 (N_2367,In_329,In_748);
and U2368 (N_2368,In_112,In_334);
nand U2369 (N_2369,In_350,In_395);
or U2370 (N_2370,In_132,In_574);
nor U2371 (N_2371,In_243,In_110);
or U2372 (N_2372,In_58,In_257);
and U2373 (N_2373,In_357,In_86);
nand U2374 (N_2374,In_60,In_174);
and U2375 (N_2375,In_678,In_541);
and U2376 (N_2376,In_160,In_335);
or U2377 (N_2377,In_22,In_521);
nand U2378 (N_2378,In_207,In_191);
or U2379 (N_2379,In_675,In_108);
nor U2380 (N_2380,In_489,In_656);
and U2381 (N_2381,In_618,In_645);
or U2382 (N_2382,In_129,In_366);
nor U2383 (N_2383,In_495,In_100);
and U2384 (N_2384,In_447,In_480);
nor U2385 (N_2385,In_461,In_398);
nor U2386 (N_2386,In_51,In_599);
or U2387 (N_2387,In_631,In_222);
or U2388 (N_2388,In_247,In_293);
and U2389 (N_2389,In_99,In_384);
nand U2390 (N_2390,In_85,In_726);
nor U2391 (N_2391,In_390,In_573);
nor U2392 (N_2392,In_732,In_302);
nand U2393 (N_2393,In_625,In_333);
nand U2394 (N_2394,In_502,In_536);
nand U2395 (N_2395,In_299,In_146);
nand U2396 (N_2396,In_595,In_178);
or U2397 (N_2397,In_669,In_318);
or U2398 (N_2398,In_561,In_734);
nand U2399 (N_2399,In_702,In_695);
and U2400 (N_2400,In_432,In_606);
nand U2401 (N_2401,In_251,In_145);
nand U2402 (N_2402,In_656,In_134);
nand U2403 (N_2403,In_339,In_291);
nor U2404 (N_2404,In_371,In_290);
xor U2405 (N_2405,In_642,In_173);
nand U2406 (N_2406,In_588,In_357);
nor U2407 (N_2407,In_636,In_48);
and U2408 (N_2408,In_459,In_575);
nand U2409 (N_2409,In_187,In_42);
or U2410 (N_2410,In_532,In_534);
nand U2411 (N_2411,In_381,In_370);
nor U2412 (N_2412,In_304,In_307);
nand U2413 (N_2413,In_131,In_460);
or U2414 (N_2414,In_330,In_533);
and U2415 (N_2415,In_79,In_709);
nand U2416 (N_2416,In_293,In_44);
or U2417 (N_2417,In_650,In_512);
nand U2418 (N_2418,In_154,In_311);
nand U2419 (N_2419,In_602,In_110);
nand U2420 (N_2420,In_225,In_308);
nor U2421 (N_2421,In_95,In_470);
nand U2422 (N_2422,In_166,In_135);
nand U2423 (N_2423,In_419,In_674);
nor U2424 (N_2424,In_652,In_61);
nor U2425 (N_2425,In_305,In_293);
and U2426 (N_2426,In_391,In_700);
nor U2427 (N_2427,In_423,In_517);
or U2428 (N_2428,In_208,In_693);
nor U2429 (N_2429,In_366,In_388);
or U2430 (N_2430,In_373,In_601);
nand U2431 (N_2431,In_668,In_55);
and U2432 (N_2432,In_616,In_299);
and U2433 (N_2433,In_437,In_710);
and U2434 (N_2434,In_546,In_128);
and U2435 (N_2435,In_43,In_564);
and U2436 (N_2436,In_446,In_275);
and U2437 (N_2437,In_652,In_129);
nand U2438 (N_2438,In_248,In_679);
nand U2439 (N_2439,In_212,In_287);
and U2440 (N_2440,In_597,In_484);
nor U2441 (N_2441,In_568,In_446);
and U2442 (N_2442,In_493,In_290);
nand U2443 (N_2443,In_360,In_196);
nand U2444 (N_2444,In_514,In_502);
and U2445 (N_2445,In_14,In_470);
and U2446 (N_2446,In_680,In_79);
and U2447 (N_2447,In_533,In_33);
and U2448 (N_2448,In_357,In_457);
nand U2449 (N_2449,In_433,In_188);
nor U2450 (N_2450,In_479,In_504);
nor U2451 (N_2451,In_538,In_648);
nand U2452 (N_2452,In_634,In_553);
nand U2453 (N_2453,In_695,In_598);
nand U2454 (N_2454,In_623,In_587);
nor U2455 (N_2455,In_357,In_232);
nor U2456 (N_2456,In_285,In_24);
and U2457 (N_2457,In_448,In_682);
or U2458 (N_2458,In_43,In_547);
nor U2459 (N_2459,In_321,In_27);
or U2460 (N_2460,In_272,In_478);
and U2461 (N_2461,In_208,In_268);
nor U2462 (N_2462,In_513,In_64);
or U2463 (N_2463,In_243,In_238);
and U2464 (N_2464,In_681,In_361);
nor U2465 (N_2465,In_414,In_200);
nor U2466 (N_2466,In_619,In_350);
nor U2467 (N_2467,In_185,In_514);
or U2468 (N_2468,In_465,In_463);
and U2469 (N_2469,In_410,In_529);
and U2470 (N_2470,In_630,In_205);
or U2471 (N_2471,In_412,In_560);
and U2472 (N_2472,In_133,In_228);
or U2473 (N_2473,In_490,In_369);
nand U2474 (N_2474,In_417,In_482);
and U2475 (N_2475,In_572,In_98);
nor U2476 (N_2476,In_530,In_655);
and U2477 (N_2477,In_526,In_231);
and U2478 (N_2478,In_741,In_490);
or U2479 (N_2479,In_616,In_294);
nor U2480 (N_2480,In_620,In_603);
xor U2481 (N_2481,In_388,In_38);
nor U2482 (N_2482,In_347,In_613);
or U2483 (N_2483,In_199,In_203);
or U2484 (N_2484,In_483,In_181);
and U2485 (N_2485,In_645,In_127);
nand U2486 (N_2486,In_610,In_236);
nand U2487 (N_2487,In_241,In_407);
and U2488 (N_2488,In_736,In_579);
nor U2489 (N_2489,In_219,In_613);
or U2490 (N_2490,In_12,In_77);
nor U2491 (N_2491,In_205,In_509);
or U2492 (N_2492,In_121,In_245);
and U2493 (N_2493,In_214,In_242);
and U2494 (N_2494,In_712,In_494);
nand U2495 (N_2495,In_412,In_186);
nand U2496 (N_2496,In_534,In_41);
nor U2497 (N_2497,In_230,In_695);
or U2498 (N_2498,In_224,In_516);
xnor U2499 (N_2499,In_374,In_450);
and U2500 (N_2500,N_317,N_2461);
and U2501 (N_2501,N_2261,N_2164);
or U2502 (N_2502,N_1032,N_2017);
nor U2503 (N_2503,N_2379,N_2268);
and U2504 (N_2504,N_1413,N_620);
nor U2505 (N_2505,N_1126,N_344);
or U2506 (N_2506,N_694,N_1960);
and U2507 (N_2507,N_2051,N_1366);
nor U2508 (N_2508,N_618,N_70);
or U2509 (N_2509,N_1967,N_763);
or U2510 (N_2510,N_179,N_37);
nand U2511 (N_2511,N_2236,N_80);
nor U2512 (N_2512,N_2493,N_1769);
nand U2513 (N_2513,N_504,N_2464);
and U2514 (N_2514,N_2234,N_32);
and U2515 (N_2515,N_1014,N_211);
nor U2516 (N_2516,N_1172,N_2120);
or U2517 (N_2517,N_2310,N_217);
nor U2518 (N_2518,N_2292,N_1381);
or U2519 (N_2519,N_1723,N_2007);
nor U2520 (N_2520,N_564,N_227);
nand U2521 (N_2521,N_2099,N_1911);
nand U2522 (N_2522,N_2297,N_2455);
nor U2523 (N_2523,N_1080,N_1718);
or U2524 (N_2524,N_2313,N_2135);
nor U2525 (N_2525,N_1238,N_1886);
or U2526 (N_2526,N_1510,N_468);
nor U2527 (N_2527,N_734,N_316);
nand U2528 (N_2528,N_1362,N_2121);
nand U2529 (N_2529,N_666,N_1842);
nand U2530 (N_2530,N_2494,N_1936);
nand U2531 (N_2531,N_1865,N_2491);
and U2532 (N_2532,N_1878,N_263);
and U2533 (N_2533,N_932,N_1214);
xnor U2534 (N_2534,N_509,N_831);
and U2535 (N_2535,N_1262,N_327);
nor U2536 (N_2536,N_2417,N_552);
xor U2537 (N_2537,N_2492,N_1115);
and U2538 (N_2538,N_2406,N_1927);
or U2539 (N_2539,N_140,N_880);
and U2540 (N_2540,N_341,N_150);
and U2541 (N_2541,N_1902,N_1309);
or U2542 (N_2542,N_1016,N_496);
nand U2543 (N_2543,N_982,N_794);
or U2544 (N_2544,N_1734,N_2317);
xnor U2545 (N_2545,N_968,N_303);
and U2546 (N_2546,N_358,N_299);
and U2547 (N_2547,N_2114,N_1209);
nor U2548 (N_2548,N_1537,N_2133);
nor U2549 (N_2549,N_2361,N_1290);
nand U2550 (N_2550,N_2032,N_1876);
or U2551 (N_2551,N_2411,N_124);
or U2552 (N_2552,N_44,N_1867);
or U2553 (N_2553,N_1010,N_1849);
or U2554 (N_2554,N_605,N_1604);
or U2555 (N_2555,N_2260,N_1012);
or U2556 (N_2556,N_2288,N_2278);
or U2557 (N_2557,N_759,N_951);
or U2558 (N_2558,N_1311,N_2239);
nand U2559 (N_2559,N_2356,N_43);
nand U2560 (N_2560,N_877,N_2423);
nand U2561 (N_2561,N_349,N_626);
and U2562 (N_2562,N_209,N_659);
or U2563 (N_2563,N_410,N_1836);
nand U2564 (N_2564,N_174,N_1190);
nand U2565 (N_2565,N_1647,N_1475);
nand U2566 (N_2566,N_1673,N_130);
nand U2567 (N_2567,N_1184,N_17);
nand U2568 (N_2568,N_1706,N_1577);
or U2569 (N_2569,N_205,N_478);
and U2570 (N_2570,N_1061,N_1280);
nor U2571 (N_2571,N_979,N_2081);
and U2572 (N_2572,N_1151,N_1027);
and U2573 (N_2573,N_15,N_2187);
and U2574 (N_2574,N_107,N_2372);
and U2575 (N_2575,N_1662,N_2308);
nand U2576 (N_2576,N_2086,N_1654);
nor U2577 (N_2577,N_1197,N_1194);
nor U2578 (N_2578,N_2340,N_490);
and U2579 (N_2579,N_2197,N_1843);
nor U2580 (N_2580,N_1198,N_99);
nand U2581 (N_2581,N_288,N_2496);
and U2582 (N_2582,N_1720,N_2090);
nand U2583 (N_2583,N_1065,N_1685);
nand U2584 (N_2584,N_1295,N_352);
nand U2585 (N_2585,N_1155,N_1778);
or U2586 (N_2586,N_1074,N_840);
nor U2587 (N_2587,N_2141,N_2025);
and U2588 (N_2588,N_1868,N_573);
nor U2589 (N_2589,N_1226,N_531);
and U2590 (N_2590,N_2254,N_1260);
nor U2591 (N_2591,N_2403,N_260);
nand U2592 (N_2592,N_297,N_1269);
nor U2593 (N_2593,N_1367,N_952);
nor U2594 (N_2594,N_2235,N_2365);
or U2595 (N_2595,N_821,N_1009);
nor U2596 (N_2596,N_1177,N_828);
nor U2597 (N_2597,N_23,N_399);
nor U2598 (N_2598,N_440,N_801);
nand U2599 (N_2599,N_2440,N_2243);
nor U2600 (N_2600,N_296,N_1751);
nand U2601 (N_2601,N_266,N_1330);
and U2602 (N_2602,N_1946,N_558);
and U2603 (N_2603,N_2183,N_1548);
or U2604 (N_2604,N_575,N_2251);
nand U2605 (N_2605,N_2298,N_646);
nor U2606 (N_2606,N_2155,N_1030);
and U2607 (N_2607,N_616,N_64);
nor U2608 (N_2608,N_1643,N_760);
nor U2609 (N_2609,N_2448,N_1468);
xor U2610 (N_2610,N_180,N_886);
nand U2611 (N_2611,N_1363,N_1301);
and U2612 (N_2612,N_1013,N_2005);
nand U2613 (N_2613,N_2466,N_1120);
nor U2614 (N_2614,N_1979,N_1526);
and U2615 (N_2615,N_948,N_1265);
or U2616 (N_2616,N_1651,N_781);
nand U2617 (N_2617,N_2302,N_1429);
nor U2618 (N_2618,N_1002,N_1561);
nand U2619 (N_2619,N_1212,N_515);
or U2620 (N_2620,N_1037,N_768);
or U2621 (N_2621,N_2161,N_1839);
or U2622 (N_2622,N_1375,N_795);
or U2623 (N_2623,N_2381,N_936);
or U2624 (N_2624,N_1442,N_2219);
or U2625 (N_2625,N_127,N_973);
or U2626 (N_2626,N_2035,N_2256);
nand U2627 (N_2627,N_556,N_1140);
nand U2628 (N_2628,N_2212,N_108);
and U2629 (N_2629,N_940,N_1050);
or U2630 (N_2630,N_4,N_45);
or U2631 (N_2631,N_587,N_1182);
and U2632 (N_2632,N_83,N_1848);
and U2633 (N_2633,N_2281,N_1292);
nor U2634 (N_2634,N_1554,N_397);
nand U2635 (N_2635,N_1056,N_2449);
and U2636 (N_2636,N_2163,N_2453);
nand U2637 (N_2637,N_577,N_2162);
nor U2638 (N_2638,N_79,N_2429);
nor U2639 (N_2639,N_163,N_1063);
nor U2640 (N_2640,N_2244,N_2101);
or U2641 (N_2641,N_2459,N_1488);
or U2642 (N_2642,N_1502,N_2412);
nor U2643 (N_2643,N_345,N_1499);
and U2644 (N_2644,N_1327,N_1138);
and U2645 (N_2645,N_2003,N_1255);
nand U2646 (N_2646,N_2369,N_1904);
nor U2647 (N_2647,N_849,N_1915);
nor U2648 (N_2648,N_870,N_2354);
nand U2649 (N_2649,N_1321,N_2432);
nor U2650 (N_2650,N_396,N_2143);
or U2651 (N_2651,N_1620,N_194);
nand U2652 (N_2652,N_1603,N_1071);
nor U2653 (N_2653,N_571,N_756);
or U2654 (N_2654,N_1830,N_1696);
nor U2655 (N_2655,N_773,N_1459);
and U2656 (N_2656,N_993,N_1952);
nor U2657 (N_2657,N_914,N_1305);
or U2658 (N_2658,N_340,N_2434);
and U2659 (N_2659,N_1476,N_162);
nor U2660 (N_2660,N_856,N_1175);
and U2661 (N_2661,N_1855,N_422);
nand U2662 (N_2662,N_2217,N_950);
or U2663 (N_2663,N_851,N_1500);
nand U2664 (N_2664,N_1087,N_301);
nand U2665 (N_2665,N_101,N_680);
or U2666 (N_2666,N_1397,N_133);
nor U2667 (N_2667,N_2039,N_780);
and U2668 (N_2668,N_1853,N_1004);
or U2669 (N_2669,N_505,N_1707);
or U2670 (N_2670,N_1046,N_2064);
nor U2671 (N_2671,N_783,N_61);
nor U2672 (N_2672,N_1111,N_1273);
or U2673 (N_2673,N_1792,N_2377);
or U2674 (N_2674,N_290,N_579);
or U2675 (N_2675,N_1891,N_2425);
and U2676 (N_2676,N_727,N_1586);
nand U2677 (N_2677,N_2480,N_1726);
or U2678 (N_2678,N_1371,N_1732);
and U2679 (N_2679,N_1672,N_24);
nand U2680 (N_2680,N_750,N_2332);
or U2681 (N_2681,N_181,N_1395);
xor U2682 (N_2682,N_192,N_1569);
or U2683 (N_2683,N_216,N_723);
nand U2684 (N_2684,N_224,N_364);
nand U2685 (N_2685,N_741,N_2222);
nand U2686 (N_2686,N_1020,N_852);
or U2687 (N_2687,N_772,N_1096);
or U2688 (N_2688,N_1545,N_1387);
nor U2689 (N_2689,N_976,N_1248);
nor U2690 (N_2690,N_602,N_649);
or U2691 (N_2691,N_755,N_1391);
and U2692 (N_2692,N_2198,N_566);
and U2693 (N_2693,N_2285,N_1044);
and U2694 (N_2694,N_782,N_252);
or U2695 (N_2695,N_1088,N_307);
nand U2696 (N_2696,N_165,N_890);
or U2697 (N_2697,N_1105,N_2240);
or U2698 (N_2698,N_2274,N_678);
nor U2699 (N_2699,N_1462,N_189);
and U2700 (N_2700,N_1243,N_2123);
or U2701 (N_2701,N_1498,N_1642);
or U2702 (N_2702,N_958,N_758);
or U2703 (N_2703,N_2037,N_803);
xnor U2704 (N_2704,N_1690,N_386);
nand U2705 (N_2705,N_1609,N_608);
or U2706 (N_2706,N_1340,N_1926);
nand U2707 (N_2707,N_2087,N_1179);
nand U2708 (N_2708,N_1602,N_551);
nor U2709 (N_2709,N_1329,N_2151);
and U2710 (N_2710,N_2264,N_2168);
or U2711 (N_2711,N_40,N_2207);
or U2712 (N_2712,N_1378,N_1316);
and U2713 (N_2713,N_1912,N_1221);
nand U2714 (N_2714,N_231,N_2074);
and U2715 (N_2715,N_1337,N_2205);
or U2716 (N_2716,N_1547,N_116);
nand U2717 (N_2717,N_1517,N_1064);
nand U2718 (N_2718,N_1683,N_534);
or U2719 (N_2719,N_1796,N_2034);
nand U2720 (N_2720,N_1596,N_722);
or U2721 (N_2721,N_2248,N_2220);
nor U2722 (N_2722,N_1688,N_146);
nor U2723 (N_2723,N_1567,N_420);
nand U2724 (N_2724,N_1298,N_2293);
nor U2725 (N_2725,N_1006,N_1324);
nand U2726 (N_2726,N_631,N_469);
or U2727 (N_2727,N_2136,N_2036);
nand U2728 (N_2728,N_2495,N_817);
nand U2729 (N_2729,N_1990,N_406);
and U2730 (N_2730,N_1947,N_2328);
nor U2731 (N_2731,N_569,N_1208);
nor U2732 (N_2732,N_1572,N_1542);
nand U2733 (N_2733,N_1522,N_2223);
and U2734 (N_2734,N_152,N_2213);
nand U2735 (N_2735,N_1342,N_766);
or U2736 (N_2736,N_844,N_1241);
and U2737 (N_2737,N_647,N_2079);
nor U2738 (N_2738,N_1347,N_2478);
and U2739 (N_2739,N_1060,N_1514);
or U2740 (N_2740,N_221,N_1850);
nand U2741 (N_2741,N_1800,N_2375);
nand U2742 (N_2742,N_400,N_1808);
or U2743 (N_2743,N_540,N_2069);
nand U2744 (N_2744,N_819,N_925);
or U2745 (N_2745,N_319,N_2066);
nand U2746 (N_2746,N_1388,N_2176);
and U2747 (N_2747,N_241,N_675);
nand U2748 (N_2748,N_875,N_687);
nand U2749 (N_2749,N_2134,N_2218);
nor U2750 (N_2750,N_545,N_466);
nand U2751 (N_2751,N_1598,N_242);
or U2752 (N_2752,N_1213,N_1047);
nand U2753 (N_2753,N_351,N_1288);
nand U2754 (N_2754,N_970,N_1229);
nand U2755 (N_2755,N_1963,N_832);
nand U2756 (N_2756,N_141,N_1538);
or U2757 (N_2757,N_10,N_1453);
nand U2758 (N_2758,N_554,N_1760);
and U2759 (N_2759,N_2124,N_786);
nand U2760 (N_2760,N_621,N_1756);
or U2761 (N_2761,N_2345,N_506);
nand U2762 (N_2762,N_1021,N_2013);
or U2763 (N_2763,N_1112,N_1113);
and U2764 (N_2764,N_2108,N_16);
and U2765 (N_2765,N_1318,N_543);
or U2766 (N_2766,N_1159,N_1656);
nor U2767 (N_2767,N_1658,N_2247);
and U2768 (N_2768,N_962,N_1251);
nor U2769 (N_2769,N_873,N_2324);
or U2770 (N_2770,N_1998,N_1158);
nand U2771 (N_2771,N_492,N_1872);
and U2772 (N_2772,N_1948,N_735);
nand U2773 (N_2773,N_1621,N_1296);
nand U2774 (N_2774,N_1671,N_567);
and U2775 (N_2775,N_1232,N_670);
and U2776 (N_2776,N_804,N_673);
xnor U2777 (N_2777,N_395,N_1059);
and U2778 (N_2778,N_657,N_311);
and U2779 (N_2779,N_1247,N_167);
and U2780 (N_2780,N_1953,N_1687);
and U2781 (N_2781,N_517,N_206);
nor U2782 (N_2782,N_906,N_428);
or U2783 (N_2783,N_633,N_1802);
and U2784 (N_2784,N_2452,N_300);
nand U2785 (N_2785,N_1995,N_432);
and U2786 (N_2786,N_1349,N_2422);
nor U2787 (N_2787,N_60,N_557);
or U2788 (N_2788,N_156,N_595);
or U2789 (N_2789,N_113,N_894);
nor U2790 (N_2790,N_1583,N_1078);
nand U2791 (N_2791,N_1424,N_1315);
nand U2792 (N_2792,N_1574,N_1485);
nor U2793 (N_2793,N_1312,N_25);
nand U2794 (N_2794,N_915,N_363);
nor U2795 (N_2795,N_1306,N_1471);
nor U2796 (N_2796,N_1794,N_1245);
and U2797 (N_2797,N_818,N_1432);
and U2798 (N_2798,N_2267,N_2202);
nand U2799 (N_2799,N_453,N_939);
and U2800 (N_2800,N_2337,N_207);
and U2801 (N_2801,N_709,N_2242);
or U2802 (N_2802,N_953,N_2311);
nor U2803 (N_2803,N_1763,N_1085);
or U2804 (N_2804,N_1692,N_524);
nand U2805 (N_2805,N_771,N_2132);
nand U2806 (N_2806,N_1267,N_1225);
or U2807 (N_2807,N_1599,N_479);
or U2808 (N_2808,N_8,N_1370);
or U2809 (N_2809,N_474,N_1043);
nand U2810 (N_2810,N_1668,N_1667);
xor U2811 (N_2811,N_1202,N_2263);
nand U2812 (N_2812,N_1834,N_414);
nand U2813 (N_2813,N_2330,N_1530);
nor U2814 (N_2814,N_685,N_1240);
and U2815 (N_2815,N_847,N_865);
and U2816 (N_2816,N_2094,N_1768);
and U2817 (N_2817,N_1965,N_1093);
nor U2818 (N_2818,N_1752,N_2072);
nor U2819 (N_2819,N_640,N_2049);
and U2820 (N_2820,N_2472,N_681);
or U2821 (N_2821,N_14,N_1108);
or U2822 (N_2822,N_1540,N_1480);
or U2823 (N_2823,N_95,N_0);
nand U2824 (N_2824,N_1484,N_320);
nand U2825 (N_2825,N_1497,N_777);
or U2826 (N_2826,N_1258,N_1483);
and U2827 (N_2827,N_1369,N_2169);
or U2828 (N_2828,N_2258,N_825);
nand U2829 (N_2829,N_134,N_262);
nand U2830 (N_2830,N_1632,N_1610);
nand U2831 (N_2831,N_1581,N_472);
or U2832 (N_2832,N_1943,N_2450);
and U2833 (N_2833,N_829,N_994);
nand U2834 (N_2834,N_1351,N_1536);
nand U2835 (N_2835,N_1930,N_1116);
and U2836 (N_2836,N_1274,N_606);
nand U2837 (N_2837,N_1425,N_1431);
and U2838 (N_2838,N_999,N_425);
nor U2839 (N_2839,N_1680,N_2360);
nand U2840 (N_2840,N_1132,N_270);
nor U2841 (N_2841,N_368,N_934);
or U2842 (N_2842,N_1666,N_2301);
and U2843 (N_2843,N_792,N_991);
nor U2844 (N_2844,N_738,N_1293);
nor U2845 (N_2845,N_177,N_234);
nand U2846 (N_2846,N_1496,N_960);
or U2847 (N_2847,N_1961,N_1339);
and U2848 (N_2848,N_375,N_1304);
or U2849 (N_2849,N_417,N_615);
and U2850 (N_2850,N_2109,N_2409);
nand U2851 (N_2851,N_816,N_2019);
nand U2852 (N_2852,N_328,N_1747);
nand U2853 (N_2853,N_1049,N_280);
nor U2854 (N_2854,N_1029,N_1154);
nor U2855 (N_2855,N_596,N_928);
and U2856 (N_2856,N_1383,N_389);
nand U2857 (N_2857,N_1674,N_1552);
nand U2858 (N_2858,N_1460,N_411);
and U2859 (N_2859,N_1435,N_809);
and U2860 (N_2860,N_1719,N_1863);
or U2861 (N_2861,N_1508,N_1959);
nand U2862 (N_2862,N_2282,N_1977);
and U2863 (N_2863,N_1294,N_69);
or U2864 (N_2864,N_715,N_1031);
nand U2865 (N_2865,N_542,N_2250);
nor U2866 (N_2866,N_471,N_784);
or U2867 (N_2867,N_2320,N_1094);
or U2868 (N_2868,N_995,N_66);
nor U2869 (N_2869,N_1789,N_129);
or U2870 (N_2870,N_576,N_1535);
and U2871 (N_2871,N_2026,N_2245);
nor U2872 (N_2872,N_2100,N_1386);
and U2873 (N_2873,N_2184,N_87);
or U2874 (N_2874,N_942,N_720);
nor U2875 (N_2875,N_1277,N_700);
nand U2876 (N_2876,N_806,N_1938);
or U2877 (N_2877,N_31,N_2041);
or U2878 (N_2878,N_1167,N_767);
nor U2879 (N_2879,N_861,N_905);
or U2880 (N_2880,N_2352,N_1954);
nor U2881 (N_2881,N_717,N_2392);
and U2882 (N_2882,N_75,N_429);
nand U2883 (N_2883,N_1018,N_2346);
or U2884 (N_2884,N_961,N_2071);
nor U2885 (N_2885,N_1940,N_1474);
nand U2886 (N_2886,N_30,N_1841);
and U2887 (N_2887,N_1829,N_793);
nand U2888 (N_2888,N_897,N_1);
nand U2889 (N_2889,N_2287,N_1698);
and U2890 (N_2890,N_2269,N_398);
and U2891 (N_2891,N_1670,N_1454);
and U2892 (N_2892,N_998,N_1437);
or U2893 (N_2893,N_1578,N_312);
nor U2894 (N_2894,N_2393,N_2359);
and U2895 (N_2895,N_1219,N_1200);
nor U2896 (N_2896,N_529,N_2209);
or U2897 (N_2897,N_2195,N_359);
nor U2898 (N_2898,N_353,N_1308);
nor U2899 (N_2899,N_1119,N_516);
or U2900 (N_2900,N_665,N_71);
or U2901 (N_2901,N_1793,N_987);
or U2902 (N_2902,N_1407,N_1600);
or U2903 (N_2903,N_1636,N_1605);
or U2904 (N_2904,N_2150,N_2052);
and U2905 (N_2905,N_2126,N_1450);
xnor U2906 (N_2906,N_1479,N_1851);
and U2907 (N_2907,N_690,N_1585);
nor U2908 (N_2908,N_1206,N_1253);
nor U2909 (N_2909,N_650,N_2181);
nand U2910 (N_2910,N_1944,N_2068);
xor U2911 (N_2911,N_1562,N_222);
and U2912 (N_2912,N_1045,N_29);
nand U2913 (N_2913,N_1406,N_1822);
and U2914 (N_2914,N_1895,N_1576);
or U2915 (N_2915,N_1644,N_1019);
or U2916 (N_2916,N_585,N_2487);
or U2917 (N_2917,N_1958,N_1528);
or U2918 (N_2918,N_318,N_704);
and U2919 (N_2919,N_1379,N_1169);
nor U2920 (N_2920,N_1787,N_1127);
or U2921 (N_2921,N_2210,N_1591);
nand U2922 (N_2922,N_302,N_597);
xor U2923 (N_2923,N_1623,N_1814);
or U2924 (N_2924,N_698,N_1594);
xor U2925 (N_2925,N_811,N_1153);
nor U2926 (N_2926,N_2433,N_2498);
nor U2927 (N_2927,N_947,N_1580);
or U2928 (N_2928,N_989,N_697);
nand U2929 (N_2929,N_2055,N_1884);
and U2930 (N_2930,N_2447,N_1612);
nand U2931 (N_2931,N_1571,N_1457);
or U2932 (N_2932,N_35,N_689);
nand U2933 (N_2933,N_2018,N_1550);
nor U2934 (N_2934,N_151,N_1055);
nand U2935 (N_2935,N_2058,N_1317);
or U2936 (N_2936,N_1481,N_1187);
nand U2937 (N_2937,N_1412,N_2385);
nor U2938 (N_2938,N_1837,N_1054);
nand U2939 (N_2939,N_106,N_981);
and U2940 (N_2940,N_808,N_1652);
or U2941 (N_2941,N_568,N_355);
nand U2942 (N_2942,N_1721,N_480);
nor U2943 (N_2943,N_1630,N_1356);
and U2944 (N_2944,N_1336,N_1070);
and U2945 (N_2945,N_1909,N_2331);
and U2946 (N_2946,N_513,N_419);
nand U2947 (N_2947,N_1495,N_1211);
and U2948 (N_2948,N_1440,N_1051);
and U2949 (N_2949,N_1973,N_2065);
nor U2950 (N_2950,N_228,N_283);
nor U2951 (N_2951,N_244,N_1236);
and U2952 (N_2952,N_1482,N_1428);
or U2953 (N_2953,N_350,N_785);
nand U2954 (N_2954,N_1490,N_836);
nand U2955 (N_2955,N_272,N_1434);
and U2956 (N_2956,N_1874,N_2273);
or U2957 (N_2957,N_1465,N_1478);
or U2958 (N_2958,N_1282,N_1518);
nand U2959 (N_2959,N_1102,N_1803);
or U2960 (N_2960,N_2057,N_256);
and U2961 (N_2961,N_196,N_1828);
or U2962 (N_2962,N_1716,N_2386);
nand U2963 (N_2963,N_1168,N_2341);
nor U2964 (N_2964,N_1053,N_1871);
and U2965 (N_2965,N_1928,N_157);
nand U2966 (N_2966,N_889,N_2060);
nor U2967 (N_2967,N_22,N_154);
or U2968 (N_2968,N_210,N_1446);
and U2969 (N_2969,N_1712,N_424);
nand U2970 (N_2970,N_1728,N_1161);
or U2971 (N_2971,N_1185,N_853);
nor U2972 (N_2972,N_645,N_1131);
nand U2973 (N_2973,N_1157,N_88);
xor U2974 (N_2974,N_1813,N_295);
nand U2975 (N_2975,N_142,N_1109);
or U2976 (N_2976,N_1801,N_1798);
nand U2977 (N_2977,N_1117,N_1042);
nor U2978 (N_2978,N_706,N_1584);
and U2979 (N_2979,N_949,N_390);
and U2980 (N_2980,N_1854,N_243);
or U2981 (N_2981,N_1207,N_1352);
nor U2982 (N_2982,N_126,N_2063);
and U2983 (N_2983,N_761,N_562);
and U2984 (N_2984,N_102,N_185);
and U2985 (N_2985,N_837,N_1757);
nand U2986 (N_2986,N_439,N_751);
or U2987 (N_2987,N_2314,N_686);
and U2988 (N_2988,N_269,N_2130);
and U2989 (N_2989,N_525,N_1427);
and U2990 (N_2990,N_444,N_2174);
or U2991 (N_2991,N_611,N_1557);
xor U2992 (N_2992,N_245,N_1470);
or U2993 (N_2993,N_470,N_1896);
nand U2994 (N_2994,N_884,N_2445);
nor U2995 (N_2995,N_1637,N_202);
and U2996 (N_2996,N_21,N_1777);
nor U2997 (N_2997,N_139,N_1847);
nor U2998 (N_2998,N_1524,N_2465);
or U2999 (N_2999,N_1512,N_438);
nor U3000 (N_3000,N_123,N_111);
or U3001 (N_3001,N_459,N_1669);
nand U3002 (N_3002,N_708,N_1971);
and U3003 (N_3003,N_560,N_521);
nor U3004 (N_3004,N_1786,N_497);
nand U3005 (N_3005,N_2230,N_1001);
or U3006 (N_3006,N_27,N_84);
or U3007 (N_3007,N_1815,N_1141);
or U3008 (N_3008,N_1844,N_1195);
nor U3009 (N_3009,N_862,N_743);
nor U3010 (N_3010,N_1350,N_2280);
or U3011 (N_3011,N_774,N_1887);
nand U3012 (N_3012,N_2462,N_332);
nor U3013 (N_3013,N_1357,N_931);
and U3014 (N_3014,N_292,N_522);
nor U3015 (N_3015,N_1970,N_572);
or U3016 (N_3016,N_2061,N_391);
xor U3017 (N_3017,N_1641,N_11);
nor U3018 (N_3018,N_2175,N_433);
or U3019 (N_3019,N_1389,N_456);
or U3020 (N_3020,N_1693,N_2200);
nand U3021 (N_3021,N_212,N_1744);
nor U3022 (N_3022,N_122,N_2371);
xnor U3023 (N_3023,N_465,N_1589);
nor U3024 (N_3024,N_2325,N_985);
or U3025 (N_3025,N_1400,N_1754);
nor U3026 (N_3026,N_1558,N_1869);
and U3027 (N_3027,N_499,N_2115);
and U3028 (N_3028,N_1319,N_1076);
and U3029 (N_3029,N_199,N_2272);
nand U3030 (N_3030,N_2499,N_2275);
or U3031 (N_3031,N_1039,N_1272);
or U3032 (N_3032,N_776,N_2042);
and U3033 (N_3033,N_943,N_1422);
or U3034 (N_3034,N_1655,N_247);
or U3035 (N_3035,N_1361,N_2300);
nand U3036 (N_3036,N_1799,N_2388);
nand U3037 (N_3037,N_96,N_143);
or U3038 (N_3038,N_2421,N_2118);
or U3039 (N_3039,N_1941,N_1264);
or U3040 (N_3040,N_799,N_1722);
or U3041 (N_3041,N_166,N_1903);
nor U3042 (N_3042,N_764,N_36);
nand U3043 (N_3043,N_520,N_2395);
nor U3044 (N_3044,N_966,N_436);
and U3045 (N_3045,N_1727,N_1417);
nor U3046 (N_3046,N_502,N_2246);
or U3047 (N_3047,N_2128,N_1544);
nand U3048 (N_3048,N_1919,N_1564);
and U3049 (N_3049,N_1974,N_1783);
or U3050 (N_3050,N_528,N_1890);
or U3051 (N_3051,N_731,N_537);
or U3052 (N_3052,N_376,N_1714);
and U3053 (N_3053,N_171,N_2249);
nand U3054 (N_3054,N_712,N_1993);
nand U3055 (N_3055,N_2075,N_1742);
nor U3056 (N_3056,N_604,N_864);
and U3057 (N_3057,N_1403,N_2188);
nor U3058 (N_3058,N_2299,N_339);
or U3059 (N_3059,N_1077,N_1216);
nor U3060 (N_3060,N_2228,N_854);
and U3061 (N_3061,N_314,N_491);
nand U3062 (N_3062,N_239,N_1880);
and U3063 (N_3063,N_2316,N_791);
nor U3064 (N_3064,N_1934,N_1942);
nand U3065 (N_3065,N_775,N_1899);
nand U3066 (N_3066,N_1331,N_184);
and U3067 (N_3067,N_2252,N_85);
nand U3068 (N_3068,N_251,N_613);
xor U3069 (N_3069,N_484,N_49);
or U3070 (N_3070,N_1289,N_1447);
or U3071 (N_3071,N_2399,N_752);
and U3072 (N_3072,N_488,N_1401);
or U3073 (N_3073,N_1753,N_1156);
or U3074 (N_3074,N_749,N_872);
nor U3075 (N_3075,N_1989,N_813);
and U3076 (N_3076,N_1160,N_2376);
and U3077 (N_3077,N_1575,N_1040);
nand U3078 (N_3078,N_1631,N_737);
or U3079 (N_3079,N_278,N_1246);
or U3080 (N_3080,N_1617,N_1992);
xor U3081 (N_3081,N_1023,N_2321);
nor U3082 (N_3082,N_1533,N_1394);
and U3083 (N_3083,N_2418,N_1507);
and U3084 (N_3084,N_1663,N_2334);
nor U3085 (N_3085,N_1067,N_121);
nand U3086 (N_3086,N_1504,N_2323);
nand U3087 (N_3087,N_2015,N_1531);
and U3088 (N_3088,N_1354,N_2454);
or U3089 (N_3089,N_322,N_1924);
nor U3090 (N_3090,N_1566,N_51);
and U3091 (N_3091,N_2333,N_2306);
or U3092 (N_3092,N_175,N_628);
nand U3093 (N_3093,N_1494,N_1750);
nor U3094 (N_3094,N_1519,N_2231);
and U3095 (N_3095,N_1925,N_805);
nor U3096 (N_3096,N_1618,N_1263);
nand U3097 (N_3097,N_2259,N_2097);
or U3098 (N_3098,N_1149,N_1917);
nor U3099 (N_3099,N_407,N_695);
nand U3100 (N_3100,N_2318,N_1083);
and U3101 (N_3101,N_1196,N_200);
nand U3102 (N_3102,N_426,N_2428);
and U3103 (N_3103,N_1313,N_892);
or U3104 (N_3104,N_1755,N_68);
or U3105 (N_3105,N_500,N_294);
nor U3106 (N_3106,N_2398,N_1439);
nand U3107 (N_3107,N_178,N_1606);
or U3108 (N_3108,N_2257,N_2167);
or U3109 (N_3109,N_699,N_519);
and U3110 (N_3110,N_1913,N_1748);
nor U3111 (N_3111,N_888,N_1908);
nor U3112 (N_3112,N_898,N_1436);
nand U3113 (N_3113,N_2366,N_323);
nand U3114 (N_3114,N_2490,N_2489);
and U3115 (N_3115,N_693,N_530);
nand U3116 (N_3116,N_1449,N_33);
or U3117 (N_3117,N_1443,N_1334);
or U3118 (N_3118,N_2374,N_779);
nor U3119 (N_3119,N_1870,N_638);
nand U3120 (N_3120,N_574,N_923);
and U3121 (N_3121,N_1877,N_1950);
nand U3122 (N_3122,N_172,N_921);
nand U3123 (N_3123,N_219,N_2067);
or U3124 (N_3124,N_2145,N_1066);
nand U3125 (N_3125,N_2295,N_1660);
nand U3126 (N_3126,N_830,N_431);
or U3127 (N_3127,N_1174,N_26);
and U3128 (N_3128,N_1615,N_2111);
nor U3129 (N_3129,N_2457,N_963);
nor U3130 (N_3130,N_2098,N_1461);
or U3131 (N_3131,N_1710,N_273);
and U3132 (N_3132,N_2347,N_553);
nor U3133 (N_3133,N_97,N_878);
nor U3134 (N_3134,N_2107,N_369);
or U3135 (N_3135,N_56,N_2102);
and U3136 (N_3136,N_827,N_213);
or U3137 (N_3137,N_1415,N_676);
nor U3138 (N_3138,N_1858,N_2214);
nand U3139 (N_3139,N_2192,N_1758);
nand U3140 (N_3140,N_1682,N_1242);
nand U3141 (N_3141,N_2336,N_423);
or U3142 (N_3142,N_413,N_2451);
nand U3143 (N_3143,N_895,N_1729);
and U3144 (N_3144,N_1003,N_977);
and U3145 (N_3145,N_1073,N_986);
or U3146 (N_3146,N_1181,N_826);
or U3147 (N_3147,N_1840,N_2216);
nor U3148 (N_3148,N_1980,N_2400);
and U3149 (N_3149,N_661,N_430);
or U3150 (N_3150,N_1419,N_238);
nor U3151 (N_3151,N_972,N_1996);
or U3152 (N_3152,N_434,N_2238);
nor U3153 (N_3153,N_1089,N_2482);
and U3154 (N_3154,N_144,N_1467);
nand U3155 (N_3155,N_2125,N_1343);
or U3156 (N_3156,N_546,N_1227);
and U3157 (N_3157,N_1964,N_683);
nor U3158 (N_3158,N_739,N_1588);
nand U3159 (N_3159,N_1675,N_1008);
nand U3160 (N_3160,N_281,N_1824);
nor U3161 (N_3161,N_822,N_944);
nor U3162 (N_3162,N_2054,N_2131);
nand U3163 (N_3163,N_1717,N_2009);
xnor U3164 (N_3164,N_2046,N_916);
and U3165 (N_3165,N_1303,N_688);
nor U3166 (N_3166,N_2363,N_361);
or U3167 (N_3167,N_1164,N_421);
and U3168 (N_3168,N_198,N_1888);
nor U3169 (N_3169,N_744,N_89);
nor U3170 (N_3170,N_2326,N_2229);
xnor U3171 (N_3171,N_1825,N_1393);
and U3172 (N_3172,N_1595,N_1806);
nor U3173 (N_3173,N_669,N_326);
nand U3174 (N_3174,N_2002,N_2170);
nor U3175 (N_3175,N_1657,N_2062);
nand U3176 (N_3176,N_2348,N_711);
and U3177 (N_3177,N_726,N_2225);
xnor U3178 (N_3178,N_1137,N_1404);
and U3179 (N_3179,N_374,N_362);
nor U3180 (N_3180,N_912,N_1041);
nand U3181 (N_3181,N_1859,N_220);
and U3182 (N_3182,N_2226,N_1746);
nand U3183 (N_3183,N_2177,N_753);
or U3184 (N_3184,N_2303,N_2266);
and U3185 (N_3185,N_1582,N_2179);
nand U3186 (N_3186,N_47,N_812);
and U3187 (N_3187,N_2182,N_2437);
nor U3188 (N_3188,N_839,N_2355);
or U3189 (N_3189,N_237,N_2148);
or U3190 (N_3190,N_2085,N_1593);
nor U3191 (N_3191,N_1410,N_1015);
and U3192 (N_3192,N_493,N_2439);
nand U3193 (N_3193,N_2485,N_2294);
or U3194 (N_3194,N_330,N_2001);
nand U3195 (N_3195,N_2160,N_347);
nand U3196 (N_3196,N_807,N_2405);
nor U3197 (N_3197,N_1521,N_2224);
nand U3198 (N_3198,N_1268,N_1935);
nand U3199 (N_3199,N_536,N_1420);
nand U3200 (N_3200,N_1776,N_487);
and U3201 (N_3201,N_135,N_2389);
nand U3202 (N_3202,N_2185,N_1322);
nand U3203 (N_3203,N_971,N_1646);
or U3204 (N_3204,N_2327,N_1703);
and U3205 (N_3205,N_846,N_589);
nor U3206 (N_3206,N_1901,N_403);
nand U3207 (N_3207,N_1501,N_1987);
and U3208 (N_3208,N_277,N_721);
nand U3209 (N_3209,N_1894,N_476);
nand U3210 (N_3210,N_1250,N_482);
nand U3211 (N_3211,N_909,N_757);
or U3212 (N_3212,N_1900,N_334);
or U3213 (N_3213,N_1384,N_2172);
nand U3214 (N_3214,N_86,N_860);
and U3215 (N_3215,N_1788,N_2383);
or U3216 (N_3216,N_1118,N_891);
nor U3217 (N_3217,N_1114,N_1364);
or U3218 (N_3218,N_1715,N_1739);
and U3219 (N_3219,N_2394,N_230);
or U3220 (N_3220,N_388,N_1058);
and U3221 (N_3221,N_2382,N_1816);
or U3222 (N_3222,N_920,N_356);
or U3223 (N_3223,N_1705,N_1281);
or U3224 (N_3224,N_1451,N_246);
or U3225 (N_3225,N_959,N_929);
nor U3226 (N_3226,N_1176,N_1770);
nor U3227 (N_3227,N_2180,N_1122);
nor U3228 (N_3228,N_1133,N_2186);
nand U3229 (N_3229,N_2416,N_104);
and U3230 (N_3230,N_2040,N_477);
nand U3231 (N_3231,N_578,N_1810);
and U3232 (N_3232,N_610,N_1697);
and U3233 (N_3233,N_1882,N_2191);
nand U3234 (N_3234,N_20,N_276);
and U3235 (N_3235,N_1270,N_2157);
nand U3236 (N_3236,N_232,N_1555);
or U3237 (N_3237,N_842,N_1130);
xnor U3238 (N_3238,N_810,N_383);
nor U3239 (N_3239,N_1325,N_625);
and U3240 (N_3240,N_918,N_1966);
nor U3241 (N_3241,N_696,N_1635);
and U3242 (N_3242,N_448,N_1456);
nand U3243 (N_3243,N_984,N_451);
and U3244 (N_3244,N_160,N_308);
nor U3245 (N_3245,N_634,N_1741);
and U3246 (N_3246,N_2029,N_473);
nor U3247 (N_3247,N_539,N_769);
nand U3248 (N_3248,N_1759,N_1579);
nand U3249 (N_3249,N_149,N_729);
and U3250 (N_3250,N_654,N_28);
or U3251 (N_3251,N_2446,N_1835);
nand U3252 (N_3252,N_1740,N_483);
or U3253 (N_3253,N_65,N_1139);
nor U3254 (N_3254,N_549,N_1234);
nand U3255 (N_3255,N_1228,N_1222);
or U3256 (N_3256,N_2270,N_820);
nand U3257 (N_3257,N_78,N_367);
nor U3258 (N_3258,N_1679,N_5);
nand U3259 (N_3259,N_858,N_899);
nor U3260 (N_3260,N_481,N_2022);
or U3261 (N_3261,N_583,N_110);
nor U3262 (N_3262,N_903,N_885);
nor U3263 (N_3263,N_1689,N_105);
nand U3264 (N_3264,N_937,N_1873);
nand U3265 (N_3265,N_191,N_1186);
or U3266 (N_3266,N_1982,N_630);
xor U3267 (N_3267,N_1441,N_705);
and U3268 (N_3268,N_823,N_1861);
nand U3269 (N_3269,N_1145,N_1135);
nor U3270 (N_3270,N_1897,N_1984);
nand U3271 (N_3271,N_1418,N_798);
nand U3272 (N_3272,N_1005,N_2391);
nor U3273 (N_3273,N_348,N_935);
and U3274 (N_3274,N_401,N_1864);
nor U3275 (N_3275,N_2030,N_1099);
nor U3276 (N_3276,N_1541,N_523);
or U3277 (N_3277,N_1784,N_145);
or U3278 (N_3278,N_800,N_2276);
nor U3279 (N_3279,N_1527,N_716);
nor U3280 (N_3280,N_674,N_732);
nand U3281 (N_3281,N_2368,N_684);
xor U3282 (N_3282,N_1279,N_2023);
or U3283 (N_3283,N_1625,N_2153);
or U3284 (N_3284,N_2483,N_850);
nand U3285 (N_3285,N_1081,N_463);
nor U3286 (N_3286,N_1807,N_561);
and U3287 (N_3287,N_1183,N_1626);
nor U3288 (N_3288,N_2396,N_692);
or U3289 (N_3289,N_1286,N_617);
nand U3290 (N_3290,N_1291,N_1192);
or U3291 (N_3291,N_1314,N_1563);
and U3292 (N_3292,N_1146,N_623);
or U3293 (N_3293,N_2122,N_745);
nand U3294 (N_3294,N_371,N_2038);
and U3295 (N_3295,N_164,N_291);
xnor U3296 (N_3296,N_1028,N_187);
nor U3297 (N_3297,N_412,N_1881);
nand U3298 (N_3298,N_402,N_1565);
or U3299 (N_3299,N_2080,N_1818);
or U3300 (N_3300,N_725,N_833);
or U3301 (N_3301,N_1601,N_1376);
nand U3302 (N_3302,N_974,N_1539);
or U3303 (N_3303,N_1650,N_1421);
and U3304 (N_3304,N_416,N_1189);
nor U3305 (N_3305,N_538,N_2144);
nand U3306 (N_3306,N_235,N_261);
nand U3307 (N_3307,N_1949,N_1489);
nor U3308 (N_3308,N_1405,N_624);
or U3309 (N_3309,N_1191,N_1695);
or U3310 (N_3310,N_445,N_1627);
or U3311 (N_3311,N_1086,N_1780);
nand U3312 (N_3312,N_1011,N_188);
and U3313 (N_3313,N_956,N_619);
or U3314 (N_3314,N_1414,N_2441);
nand U3315 (N_3315,N_1101,N_1616);
or U3316 (N_3316,N_236,N_360);
nand U3317 (N_3317,N_874,N_1811);
nor U3318 (N_3318,N_1981,N_1052);
or U3319 (N_3319,N_1832,N_336);
nand U3320 (N_3320,N_679,N_1922);
and U3321 (N_3321,N_298,N_607);
and U3322 (N_3322,N_306,N_1075);
nand U3323 (N_3323,N_329,N_957);
nor U3324 (N_3324,N_1205,N_2158);
and U3325 (N_3325,N_1945,N_2028);
nand U3326 (N_3326,N_1173,N_1180);
nor U3327 (N_3327,N_2473,N_1463);
and U3328 (N_3328,N_346,N_643);
or U3329 (N_3329,N_1889,N_748);
nor U3330 (N_3330,N_195,N_1898);
and U3331 (N_3331,N_778,N_713);
nand U3332 (N_3332,N_1452,N_2353);
and U3333 (N_3333,N_1491,N_2468);
or U3334 (N_3334,N_1091,N_841);
or U3335 (N_3335,N_1866,N_1493);
nand U3336 (N_3336,N_193,N_2232);
and U3337 (N_3337,N_1433,N_2073);
and U3338 (N_3338,N_1920,N_2410);
nor U3339 (N_3339,N_2000,N_1856);
nor U3340 (N_3340,N_1857,N_310);
nand U3341 (N_3341,N_254,N_983);
or U3342 (N_3342,N_315,N_2142);
and U3343 (N_3343,N_1411,N_1092);
nand U3344 (N_3344,N_462,N_1385);
nor U3345 (N_3345,N_2414,N_910);
or U3346 (N_3346,N_1553,N_526);
and U3347 (N_3347,N_394,N_12);
nor U3348 (N_3348,N_2138,N_2307);
nand U3349 (N_3349,N_1516,N_598);
and U3350 (N_3350,N_1691,N_967);
nor U3351 (N_3351,N_331,N_1738);
nand U3352 (N_3352,N_718,N_1398);
nor U3353 (N_3353,N_730,N_1372);
nand U3354 (N_3354,N_2093,N_1505);
nand U3355 (N_3355,N_667,N_1134);
nand U3356 (N_3356,N_1929,N_1556);
xnor U3357 (N_3357,N_2431,N_2289);
nand U3358 (N_3358,N_1188,N_3);
nor U3359 (N_3359,N_1374,N_1233);
or U3360 (N_3360,N_1906,N_2027);
nor U3361 (N_3361,N_467,N_1166);
and U3362 (N_3362,N_714,N_2117);
or U3363 (N_3363,N_2233,N_1676);
and U3364 (N_3364,N_215,N_1110);
nor U3365 (N_3365,N_1883,N_1817);
nor U3366 (N_3366,N_1923,N_1223);
and U3367 (N_3367,N_475,N_1344);
nor U3368 (N_3368,N_2277,N_2402);
and U3369 (N_3369,N_765,N_924);
nand U3370 (N_3370,N_1885,N_535);
and U3371 (N_3371,N_2349,N_1597);
nor U3372 (N_3372,N_2201,N_115);
nand U3373 (N_3373,N_226,N_788);
and U3374 (N_3374,N_1731,N_354);
nand U3375 (N_3375,N_724,N_258);
and U3376 (N_3376,N_1775,N_103);
or U3377 (N_3377,N_922,N_1022);
or U3378 (N_3378,N_1487,N_507);
or U3379 (N_3379,N_338,N_1916);
nor U3380 (N_3380,N_1568,N_385);
or U3381 (N_3381,N_2291,N_1951);
or U3382 (N_3382,N_2350,N_1244);
and U3383 (N_3383,N_1095,N_53);
and U3384 (N_3384,N_2140,N_2435);
or U3385 (N_3385,N_2284,N_599);
or U3386 (N_3386,N_100,N_627);
nand U3387 (N_3387,N_2370,N_1472);
nor U3388 (N_3388,N_1335,N_1237);
or U3389 (N_3389,N_662,N_1968);
and U3390 (N_3390,N_2059,N_590);
or U3391 (N_3391,N_392,N_879);
nor U3392 (N_3392,N_119,N_580);
and U3393 (N_3393,N_614,N_1664);
nor U3394 (N_3394,N_1745,N_2315);
or U3395 (N_3395,N_1283,N_2484);
or U3396 (N_3396,N_1782,N_457);
and U3397 (N_3397,N_1905,N_1638);
nand U3398 (N_3398,N_1057,N_2384);
or U3399 (N_3399,N_2474,N_1103);
nor U3400 (N_3400,N_1100,N_1838);
nor U3401 (N_3401,N_427,N_158);
nand U3402 (N_3402,N_1346,N_1034);
nand U3403 (N_3403,N_2283,N_644);
and U3404 (N_3404,N_1106,N_1152);
and U3405 (N_3405,N_2089,N_136);
or U3406 (N_3406,N_900,N_2165);
and U3407 (N_3407,N_927,N_887);
or U3408 (N_3408,N_2011,N_1231);
or U3409 (N_3409,N_591,N_1653);
or U3410 (N_3410,N_510,N_415);
nand U3411 (N_3411,N_1000,N_790);
or U3412 (N_3412,N_408,N_1147);
nand U3413 (N_3413,N_1678,N_271);
or U3414 (N_3414,N_2206,N_1026);
and U3415 (N_3415,N_997,N_1875);
and U3416 (N_3416,N_2470,N_117);
nor U3417 (N_3417,N_1932,N_1771);
nand U3418 (N_3418,N_447,N_1148);
nor U3419 (N_3419,N_988,N_1276);
nor U3420 (N_3420,N_1918,N_203);
or U3421 (N_3421,N_1062,N_1464);
nand U3422 (N_3422,N_286,N_1713);
and U3423 (N_3423,N_1975,N_267);
nand U3424 (N_3424,N_1017,N_639);
or U3425 (N_3425,N_92,N_2467);
nor U3426 (N_3426,N_1708,N_1445);
and U3427 (N_3427,N_293,N_1038);
nand U3428 (N_3428,N_1271,N_1284);
nand U3429 (N_3429,N_655,N_582);
nand U3430 (N_3430,N_2048,N_59);
nor U3431 (N_3431,N_1097,N_1123);
nand U3432 (N_3432,N_2045,N_902);
nor U3433 (N_3433,N_1629,N_18);
nor U3434 (N_3434,N_1007,N_1937);
or U3435 (N_3435,N_1699,N_2112);
nor U3436 (N_3436,N_2415,N_1737);
or U3437 (N_3437,N_176,N_703);
nand U3438 (N_3438,N_57,N_229);
nor U3439 (N_3439,N_1999,N_2103);
or U3440 (N_3440,N_2104,N_460);
nor U3441 (N_3441,N_2373,N_50);
nor U3442 (N_3442,N_642,N_186);
and U3443 (N_3443,N_603,N_54);
nand U3444 (N_3444,N_1805,N_274);
nand U3445 (N_3445,N_1458,N_1749);
nand U3446 (N_3446,N_137,N_2488);
and U3447 (N_3447,N_285,N_719);
nor U3448 (N_3448,N_109,N_265);
nand U3449 (N_3449,N_1220,N_1257);
or U3450 (N_3450,N_2367,N_1570);
or U3451 (N_3451,N_1931,N_501);
or U3452 (N_3452,N_2043,N_2408);
nand U3453 (N_3453,N_2199,N_2265);
nor U3454 (N_3454,N_1513,N_1239);
and U3455 (N_3455,N_1645,N_1543);
xor U3456 (N_3456,N_1622,N_641);
or U3457 (N_3457,N_1204,N_2012);
nand U3458 (N_3458,N_1163,N_789);
and U3459 (N_3459,N_1359,N_1767);
or U3460 (N_3460,N_2020,N_2237);
or U3461 (N_3461,N_379,N_325);
and U3462 (N_3462,N_1515,N_1772);
and U3463 (N_3463,N_2427,N_1390);
nand U3464 (N_3464,N_867,N_1628);
nor U3465 (N_3465,N_1302,N_2091);
and U3466 (N_3466,N_1733,N_668);
nand U3467 (N_3467,N_2016,N_512);
and U3468 (N_3468,N_1358,N_857);
and U3469 (N_3469,N_2173,N_1700);
or U3470 (N_3470,N_393,N_257);
nand U3471 (N_3471,N_1845,N_2286);
nor U3472 (N_3472,N_1549,N_287);
and U3473 (N_3473,N_2227,N_2262);
or U3474 (N_3474,N_2419,N_250);
nor U3475 (N_3475,N_2319,N_90);
nor U3476 (N_3476,N_2271,N_2477);
nand U3477 (N_3477,N_1827,N_2178);
nand U3478 (N_3478,N_486,N_1178);
and U3479 (N_3479,N_120,N_945);
and U3480 (N_3480,N_2082,N_147);
nor U3481 (N_3481,N_2241,N_2095);
nand U3482 (N_3482,N_2443,N_594);
nand U3483 (N_3483,N_1278,N_2127);
nor U3484 (N_3484,N_2078,N_946);
nand U3485 (N_3485,N_1473,N_1819);
nand U3486 (N_3486,N_370,N_1338);
and U3487 (N_3487,N_372,N_876);
nor U3488 (N_3488,N_450,N_682);
nor U3489 (N_3489,N_1323,N_1107);
or U3490 (N_3490,N_282,N_1129);
nand U3491 (N_3491,N_485,N_1254);
nand U3492 (N_3492,N_1252,N_183);
and U3493 (N_3493,N_1820,N_1661);
nor U3494 (N_3494,N_1520,N_592);
or U3495 (N_3495,N_305,N_1320);
and U3496 (N_3496,N_1307,N_652);
and U3497 (N_3497,N_321,N_565);
nor U3498 (N_3498,N_34,N_802);
nand U3499 (N_3499,N_1939,N_2137);
and U3500 (N_3500,N_1035,N_304);
or U3501 (N_3501,N_2193,N_664);
and U3502 (N_3502,N_548,N_559);
or U3503 (N_3503,N_555,N_593);
or U3504 (N_3504,N_2203,N_2296);
and U3505 (N_3505,N_223,N_275);
or U3506 (N_3506,N_2397,N_868);
nand U3507 (N_3507,N_1826,N_1907);
and U3508 (N_3508,N_67,N_446);
or U3509 (N_3509,N_1762,N_1624);
and U3510 (N_3510,N_1275,N_2008);
and U3511 (N_3511,N_2166,N_2070);
nor U3512 (N_3512,N_635,N_1297);
nor U3513 (N_3513,N_1546,N_218);
nand U3514 (N_3514,N_1300,N_387);
nand U3515 (N_3515,N_1761,N_980);
nand U3516 (N_3516,N_637,N_1128);
nor U3517 (N_3517,N_736,N_1079);
or U3518 (N_3518,N_2088,N_2006);
and U3519 (N_3519,N_1969,N_896);
nor U3520 (N_3520,N_2021,N_441);
and U3521 (N_3521,N_1193,N_1523);
nor U3522 (N_3522,N_955,N_919);
nor U3523 (N_3523,N_1781,N_2004);
or U3524 (N_3524,N_1036,N_343);
and U3525 (N_3525,N_1224,N_489);
nand U3526 (N_3526,N_55,N_550);
nor U3527 (N_3527,N_2424,N_1215);
nor U3528 (N_3528,N_495,N_859);
nand U3529 (N_3529,N_954,N_52);
and U3530 (N_3530,N_2364,N_1590);
and U3531 (N_3531,N_42,N_2084);
or U3532 (N_3532,N_1355,N_138);
nand U3533 (N_3533,N_1852,N_2116);
nand U3534 (N_3534,N_118,N_1466);
or U3535 (N_3535,N_1525,N_240);
nand U3536 (N_3536,N_1048,N_2105);
or U3537 (N_3537,N_1310,N_1285);
nor U3538 (N_3538,N_357,N_2014);
nand U3539 (N_3539,N_2335,N_1333);
nand U3540 (N_3540,N_2456,N_881);
and U3541 (N_3541,N_648,N_651);
nor U3542 (N_3542,N_740,N_869);
nor U3543 (N_3543,N_1534,N_1341);
and U3544 (N_3544,N_508,N_609);
nor U3545 (N_3545,N_2204,N_2196);
and U3546 (N_3546,N_1659,N_1833);
nand U3547 (N_3547,N_309,N_1509);
and U3548 (N_3548,N_1068,N_863);
or U3549 (N_3549,N_2343,N_2342);
nand U3550 (N_3550,N_1365,N_464);
nand U3551 (N_3551,N_452,N_824);
nand U3552 (N_3552,N_835,N_1978);
or U3553 (N_3553,N_964,N_2010);
and U3554 (N_3554,N_1831,N_1033);
nor U3555 (N_3555,N_1972,N_313);
and U3556 (N_3556,N_1677,N_259);
or U3557 (N_3557,N_2344,N_48);
and U3558 (N_3558,N_1613,N_1392);
and U3559 (N_3559,N_996,N_381);
nand U3560 (N_3560,N_612,N_170);
or U3561 (N_3561,N_855,N_733);
xnor U3562 (N_3562,N_1104,N_1409);
nand U3563 (N_3563,N_511,N_1611);
or U3564 (N_3564,N_1448,N_255);
or U3565 (N_3565,N_1684,N_380);
or U3566 (N_3566,N_2305,N_443);
nand U3567 (N_3567,N_38,N_843);
and U3568 (N_3568,N_2110,N_742);
nor U3569 (N_3569,N_1809,N_2279);
nor U3570 (N_3570,N_2047,N_125);
and U3571 (N_3571,N_746,N_93);
and U3572 (N_3572,N_707,N_677);
and U3573 (N_3573,N_1396,N_933);
nand U3574 (N_3574,N_1024,N_1587);
and U3575 (N_3575,N_581,N_454);
or U3576 (N_3576,N_1210,N_2076);
nand U3577 (N_3577,N_1299,N_6);
nor U3578 (N_3578,N_1988,N_1764);
nand U3579 (N_3579,N_201,N_1348);
or U3580 (N_3580,N_893,N_132);
nand U3581 (N_3581,N_2339,N_1701);
nand U3582 (N_3582,N_527,N_112);
and U3583 (N_3583,N_173,N_814);
nor U3584 (N_3584,N_159,N_671);
nand U3585 (N_3585,N_1773,N_1469);
nor U3586 (N_3586,N_588,N_1879);
and U3587 (N_3587,N_365,N_2358);
and U3588 (N_3588,N_1665,N_1529);
or U3589 (N_3589,N_131,N_656);
and U3590 (N_3590,N_1025,N_1259);
nor U3591 (N_3591,N_1506,N_1962);
or U3592 (N_3592,N_1143,N_1266);
nand U3593 (N_3593,N_1649,N_1933);
nor U3594 (N_3594,N_1235,N_930);
or U3595 (N_3595,N_563,N_63);
nor U3596 (N_3596,N_1991,N_161);
nand U3597 (N_3597,N_658,N_2312);
nor U3598 (N_3598,N_1402,N_418);
nand U3599 (N_3599,N_2407,N_1560);
and U3600 (N_3600,N_913,N_1735);
and U3601 (N_3601,N_1914,N_547);
nor U3602 (N_3602,N_73,N_2044);
or U3603 (N_3603,N_225,N_663);
nand U3604 (N_3604,N_584,N_1455);
or U3605 (N_3605,N_2221,N_2056);
and U3606 (N_3606,N_1170,N_2413);
nor U3607 (N_3607,N_289,N_1328);
or U3608 (N_3608,N_2438,N_378);
xnor U3609 (N_3609,N_2253,N_2149);
or U3610 (N_3610,N_2194,N_2460);
nand U3611 (N_3611,N_1503,N_2481);
and U3612 (N_3612,N_1812,N_7);
and U3613 (N_3613,N_1423,N_9);
nor U3614 (N_3614,N_2329,N_155);
nor U3615 (N_3615,N_1162,N_2119);
nand U3616 (N_3616,N_1765,N_2401);
or U3617 (N_3617,N_532,N_926);
and U3618 (N_3618,N_969,N_710);
nor U3619 (N_3619,N_2050,N_2208);
nand U3620 (N_3620,N_701,N_1332);
nor U3621 (N_3621,N_19,N_1957);
and U3622 (N_3622,N_2211,N_2430);
nor U3623 (N_3623,N_449,N_1702);
and U3624 (N_3624,N_1199,N_264);
nand U3625 (N_3625,N_834,N_1072);
or U3626 (N_3626,N_366,N_1639);
nand U3627 (N_3627,N_754,N_2442);
and U3628 (N_3628,N_883,N_46);
and U3629 (N_3629,N_1360,N_660);
nand U3630 (N_3630,N_1373,N_728);
nand U3631 (N_3631,N_384,N_405);
nor U3632 (N_3632,N_2129,N_622);
or U3633 (N_3633,N_2290,N_838);
nand U3634 (N_3634,N_2390,N_1892);
nand U3635 (N_3635,N_796,N_1956);
nand U3636 (N_3636,N_197,N_1551);
and U3637 (N_3637,N_342,N_1142);
nand U3638 (N_3638,N_503,N_1326);
and U3639 (N_3639,N_702,N_1426);
and U3640 (N_3640,N_1862,N_1082);
nand U3641 (N_3641,N_442,N_214);
nor U3642 (N_3642,N_1218,N_248);
and U3643 (N_3643,N_1256,N_1559);
nor U3644 (N_3644,N_1607,N_249);
nor U3645 (N_3645,N_901,N_190);
nor U3646 (N_3646,N_1430,N_2338);
nand U3647 (N_3647,N_1795,N_1694);
or U3648 (N_3648,N_1532,N_409);
nor U3649 (N_3649,N_1592,N_1492);
and U3650 (N_3650,N_1399,N_1124);
nand U3651 (N_3651,N_2096,N_337);
and U3652 (N_3652,N_1090,N_978);
or U3653 (N_3653,N_458,N_1704);
nor U3654 (N_3654,N_62,N_2380);
and U3655 (N_3655,N_153,N_1619);
and U3656 (N_3656,N_1681,N_882);
and U3657 (N_3657,N_871,N_1573);
and U3658 (N_3658,N_2476,N_1686);
and U3659 (N_3659,N_94,N_58);
nand U3660 (N_3660,N_2463,N_82);
or U3661 (N_3661,N_1382,N_1444);
or U3662 (N_3662,N_2190,N_787);
nor U3663 (N_3663,N_2426,N_941);
and U3664 (N_3664,N_333,N_461);
nand U3665 (N_3665,N_2479,N_76);
or U3666 (N_3666,N_1614,N_762);
and U3667 (N_3667,N_815,N_1797);
nand U3668 (N_3668,N_1955,N_148);
nand U3669 (N_3669,N_1790,N_284);
or U3670 (N_3670,N_2497,N_2362);
or U3671 (N_3671,N_2351,N_114);
nor U3672 (N_3672,N_514,N_1997);
nor U3673 (N_3673,N_2147,N_770);
and U3674 (N_3674,N_975,N_1921);
nand U3675 (N_3675,N_1477,N_1353);
nor U3676 (N_3676,N_1860,N_1791);
or U3677 (N_3677,N_797,N_437);
nand U3678 (N_3678,N_2255,N_636);
or U3679 (N_3679,N_72,N_1203);
or U3680 (N_3680,N_268,N_1249);
and U3681 (N_3681,N_204,N_1994);
or U3682 (N_3682,N_1711,N_233);
nor U3683 (N_3683,N_2106,N_1633);
nor U3684 (N_3684,N_1165,N_1136);
or U3685 (N_3685,N_1201,N_335);
nor U3686 (N_3686,N_848,N_904);
nand U3687 (N_3687,N_498,N_1634);
nand U3688 (N_3688,N_2,N_1893);
nor U3689 (N_3689,N_1098,N_2304);
nand U3690 (N_3690,N_1171,N_2092);
nand U3691 (N_3691,N_570,N_653);
xor U3692 (N_3692,N_908,N_1804);
or U3693 (N_3693,N_77,N_182);
nor U3694 (N_3694,N_601,N_1725);
and U3695 (N_3695,N_2469,N_2404);
nor U3696 (N_3696,N_128,N_2113);
or U3697 (N_3697,N_992,N_2420);
and U3698 (N_3698,N_2436,N_1976);
nor U3699 (N_3699,N_1069,N_169);
and U3700 (N_3700,N_691,N_2146);
nand U3701 (N_3701,N_917,N_2053);
and U3702 (N_3702,N_2458,N_541);
nand U3703 (N_3703,N_1730,N_98);
or U3704 (N_3704,N_208,N_1736);
and U3705 (N_3705,N_2189,N_866);
or U3706 (N_3706,N_629,N_518);
and U3707 (N_3707,N_13,N_1983);
or U3708 (N_3708,N_1608,N_747);
nand U3709 (N_3709,N_2471,N_1766);
nand U3710 (N_3710,N_845,N_74);
and U3711 (N_3711,N_2024,N_911);
nand U3712 (N_3712,N_324,N_2215);
or U3713 (N_3713,N_2387,N_2322);
or U3714 (N_3714,N_2171,N_672);
or U3715 (N_3715,N_1345,N_1121);
nand U3716 (N_3716,N_1416,N_494);
nand U3717 (N_3717,N_600,N_1380);
nand U3718 (N_3718,N_2077,N_2031);
nand U3719 (N_3719,N_1368,N_1486);
or U3720 (N_3720,N_435,N_2159);
nor U3721 (N_3721,N_455,N_533);
or U3722 (N_3722,N_1985,N_1774);
nand U3723 (N_3723,N_168,N_1823);
nor U3724 (N_3724,N_41,N_81);
and U3725 (N_3725,N_377,N_2152);
and U3726 (N_3726,N_2475,N_1230);
and U3727 (N_3727,N_544,N_1785);
nor U3728 (N_3728,N_990,N_1743);
nor U3729 (N_3729,N_1150,N_253);
and U3730 (N_3730,N_938,N_1125);
nor U3731 (N_3731,N_1986,N_2033);
or U3732 (N_3732,N_1640,N_2357);
or U3733 (N_3733,N_91,N_39);
nand U3734 (N_3734,N_1084,N_2486);
nor U3735 (N_3735,N_2378,N_1287);
xor U3736 (N_3736,N_1910,N_586);
or U3737 (N_3737,N_1144,N_1408);
nand U3738 (N_3738,N_1779,N_2139);
nand U3739 (N_3739,N_1261,N_1377);
and U3740 (N_3740,N_2156,N_2444);
nand U3741 (N_3741,N_1709,N_1846);
nor U3742 (N_3742,N_965,N_1511);
and U3743 (N_3743,N_2083,N_279);
nor U3744 (N_3744,N_382,N_1821);
or U3745 (N_3745,N_404,N_2309);
and U3746 (N_3746,N_632,N_1438);
nand U3747 (N_3747,N_1648,N_1724);
nor U3748 (N_3748,N_2154,N_907);
and U3749 (N_3749,N_1217,N_373);
or U3750 (N_3750,N_229,N_843);
and U3751 (N_3751,N_462,N_518);
or U3752 (N_3752,N_1420,N_759);
and U3753 (N_3753,N_1608,N_762);
nand U3754 (N_3754,N_1635,N_2449);
nor U3755 (N_3755,N_1776,N_680);
or U3756 (N_3756,N_1056,N_2311);
nor U3757 (N_3757,N_418,N_2448);
or U3758 (N_3758,N_989,N_2316);
nor U3759 (N_3759,N_1218,N_1237);
or U3760 (N_3760,N_1088,N_883);
and U3761 (N_3761,N_1922,N_1954);
and U3762 (N_3762,N_2440,N_351);
nor U3763 (N_3763,N_1452,N_411);
nand U3764 (N_3764,N_850,N_1232);
or U3765 (N_3765,N_779,N_615);
and U3766 (N_3766,N_901,N_401);
or U3767 (N_3767,N_1344,N_1413);
nor U3768 (N_3768,N_548,N_1491);
nor U3769 (N_3769,N_2432,N_588);
or U3770 (N_3770,N_1453,N_558);
nand U3771 (N_3771,N_1363,N_67);
nor U3772 (N_3772,N_1330,N_2188);
and U3773 (N_3773,N_2075,N_1283);
nor U3774 (N_3774,N_763,N_790);
and U3775 (N_3775,N_220,N_343);
or U3776 (N_3776,N_1873,N_548);
nor U3777 (N_3777,N_1029,N_989);
nor U3778 (N_3778,N_906,N_1086);
and U3779 (N_3779,N_2401,N_1511);
nand U3780 (N_3780,N_2326,N_1691);
nand U3781 (N_3781,N_1814,N_2410);
or U3782 (N_3782,N_132,N_2491);
nor U3783 (N_3783,N_889,N_1818);
nand U3784 (N_3784,N_1137,N_2471);
nand U3785 (N_3785,N_2435,N_1791);
or U3786 (N_3786,N_647,N_1349);
nor U3787 (N_3787,N_899,N_150);
and U3788 (N_3788,N_1890,N_2181);
and U3789 (N_3789,N_1077,N_1554);
nand U3790 (N_3790,N_1440,N_1337);
nor U3791 (N_3791,N_2051,N_2496);
nor U3792 (N_3792,N_197,N_1708);
nand U3793 (N_3793,N_2324,N_1366);
or U3794 (N_3794,N_2025,N_486);
or U3795 (N_3795,N_1282,N_1127);
nand U3796 (N_3796,N_208,N_855);
nand U3797 (N_3797,N_490,N_1272);
and U3798 (N_3798,N_1224,N_1069);
or U3799 (N_3799,N_970,N_1504);
and U3800 (N_3800,N_1060,N_1105);
and U3801 (N_3801,N_240,N_1193);
nor U3802 (N_3802,N_235,N_147);
xnor U3803 (N_3803,N_1522,N_1833);
and U3804 (N_3804,N_1871,N_293);
nor U3805 (N_3805,N_270,N_1759);
or U3806 (N_3806,N_1107,N_1540);
nand U3807 (N_3807,N_1871,N_489);
nand U3808 (N_3808,N_1181,N_2172);
or U3809 (N_3809,N_626,N_2450);
nand U3810 (N_3810,N_1914,N_1084);
or U3811 (N_3811,N_270,N_105);
nand U3812 (N_3812,N_1195,N_1136);
nor U3813 (N_3813,N_1934,N_432);
or U3814 (N_3814,N_1142,N_1630);
nor U3815 (N_3815,N_1173,N_425);
nand U3816 (N_3816,N_359,N_2076);
and U3817 (N_3817,N_117,N_651);
nand U3818 (N_3818,N_1839,N_2309);
or U3819 (N_3819,N_2419,N_70);
or U3820 (N_3820,N_245,N_1286);
nand U3821 (N_3821,N_824,N_1958);
nor U3822 (N_3822,N_624,N_665);
or U3823 (N_3823,N_1472,N_1225);
and U3824 (N_3824,N_2029,N_66);
or U3825 (N_3825,N_2114,N_1346);
or U3826 (N_3826,N_2490,N_2125);
and U3827 (N_3827,N_1387,N_1643);
nand U3828 (N_3828,N_646,N_421);
nand U3829 (N_3829,N_392,N_647);
nor U3830 (N_3830,N_1567,N_1513);
and U3831 (N_3831,N_1570,N_370);
nand U3832 (N_3832,N_1189,N_1621);
or U3833 (N_3833,N_417,N_1936);
nand U3834 (N_3834,N_890,N_436);
nor U3835 (N_3835,N_455,N_2209);
and U3836 (N_3836,N_0,N_895);
and U3837 (N_3837,N_186,N_2057);
nand U3838 (N_3838,N_2430,N_2484);
nand U3839 (N_3839,N_615,N_307);
or U3840 (N_3840,N_1930,N_2072);
or U3841 (N_3841,N_2048,N_950);
nand U3842 (N_3842,N_1709,N_206);
nor U3843 (N_3843,N_1574,N_1366);
or U3844 (N_3844,N_1921,N_2295);
or U3845 (N_3845,N_47,N_2285);
and U3846 (N_3846,N_2444,N_979);
nand U3847 (N_3847,N_803,N_1026);
nor U3848 (N_3848,N_504,N_2323);
nand U3849 (N_3849,N_566,N_968);
and U3850 (N_3850,N_112,N_1519);
nor U3851 (N_3851,N_1260,N_2364);
and U3852 (N_3852,N_2339,N_1536);
and U3853 (N_3853,N_1606,N_1277);
or U3854 (N_3854,N_1869,N_379);
and U3855 (N_3855,N_1335,N_653);
or U3856 (N_3856,N_1226,N_957);
nor U3857 (N_3857,N_464,N_712);
or U3858 (N_3858,N_1701,N_1995);
and U3859 (N_3859,N_1018,N_1834);
nand U3860 (N_3860,N_726,N_2262);
or U3861 (N_3861,N_2262,N_786);
nand U3862 (N_3862,N_856,N_1080);
nor U3863 (N_3863,N_2135,N_528);
or U3864 (N_3864,N_16,N_856);
and U3865 (N_3865,N_1647,N_87);
nand U3866 (N_3866,N_411,N_985);
or U3867 (N_3867,N_463,N_603);
and U3868 (N_3868,N_1164,N_403);
nor U3869 (N_3869,N_544,N_2367);
nor U3870 (N_3870,N_953,N_2163);
or U3871 (N_3871,N_1485,N_162);
nor U3872 (N_3872,N_1173,N_2061);
and U3873 (N_3873,N_577,N_2089);
nand U3874 (N_3874,N_929,N_1090);
and U3875 (N_3875,N_1370,N_1367);
nand U3876 (N_3876,N_2199,N_2468);
and U3877 (N_3877,N_2349,N_746);
and U3878 (N_3878,N_2445,N_1916);
and U3879 (N_3879,N_54,N_2336);
and U3880 (N_3880,N_1361,N_1024);
or U3881 (N_3881,N_2268,N_602);
nand U3882 (N_3882,N_199,N_989);
or U3883 (N_3883,N_1382,N_1680);
and U3884 (N_3884,N_711,N_342);
nand U3885 (N_3885,N_48,N_776);
nand U3886 (N_3886,N_1138,N_2290);
nor U3887 (N_3887,N_1014,N_1595);
nor U3888 (N_3888,N_682,N_2026);
nand U3889 (N_3889,N_652,N_421);
or U3890 (N_3890,N_591,N_1882);
nor U3891 (N_3891,N_148,N_1666);
nand U3892 (N_3892,N_846,N_2063);
nor U3893 (N_3893,N_2305,N_1047);
nand U3894 (N_3894,N_686,N_1576);
nand U3895 (N_3895,N_1378,N_1358);
or U3896 (N_3896,N_228,N_68);
and U3897 (N_3897,N_1465,N_220);
or U3898 (N_3898,N_785,N_346);
nor U3899 (N_3899,N_1104,N_2247);
nor U3900 (N_3900,N_561,N_1730);
or U3901 (N_3901,N_1770,N_1542);
and U3902 (N_3902,N_1541,N_493);
nand U3903 (N_3903,N_987,N_29);
or U3904 (N_3904,N_572,N_605);
nand U3905 (N_3905,N_399,N_27);
nor U3906 (N_3906,N_939,N_1530);
nand U3907 (N_3907,N_486,N_1003);
and U3908 (N_3908,N_441,N_703);
nor U3909 (N_3909,N_481,N_1697);
nand U3910 (N_3910,N_2333,N_1306);
nand U3911 (N_3911,N_34,N_1269);
or U3912 (N_3912,N_2023,N_1265);
nand U3913 (N_3913,N_2358,N_717);
or U3914 (N_3914,N_2358,N_2282);
nand U3915 (N_3915,N_1618,N_2029);
or U3916 (N_3916,N_2112,N_1084);
or U3917 (N_3917,N_2452,N_893);
or U3918 (N_3918,N_461,N_1218);
or U3919 (N_3919,N_1004,N_1219);
nand U3920 (N_3920,N_2256,N_353);
and U3921 (N_3921,N_21,N_424);
nor U3922 (N_3922,N_1340,N_1647);
or U3923 (N_3923,N_2282,N_1552);
nand U3924 (N_3924,N_1728,N_264);
nand U3925 (N_3925,N_148,N_758);
nand U3926 (N_3926,N_2048,N_1640);
or U3927 (N_3927,N_2225,N_1209);
or U3928 (N_3928,N_758,N_257);
or U3929 (N_3929,N_590,N_1460);
nand U3930 (N_3930,N_893,N_618);
or U3931 (N_3931,N_1843,N_60);
nor U3932 (N_3932,N_471,N_718);
nor U3933 (N_3933,N_1060,N_2264);
and U3934 (N_3934,N_2266,N_706);
and U3935 (N_3935,N_671,N_1634);
and U3936 (N_3936,N_112,N_1818);
and U3937 (N_3937,N_459,N_572);
and U3938 (N_3938,N_2122,N_1420);
nor U3939 (N_3939,N_1061,N_1320);
or U3940 (N_3940,N_1552,N_2065);
and U3941 (N_3941,N_2416,N_2109);
nor U3942 (N_3942,N_1627,N_2287);
and U3943 (N_3943,N_518,N_70);
or U3944 (N_3944,N_666,N_346);
or U3945 (N_3945,N_241,N_2094);
nor U3946 (N_3946,N_1787,N_367);
nor U3947 (N_3947,N_862,N_966);
or U3948 (N_3948,N_315,N_838);
nand U3949 (N_3949,N_1772,N_202);
nand U3950 (N_3950,N_18,N_1910);
nand U3951 (N_3951,N_1942,N_2237);
nand U3952 (N_3952,N_327,N_2461);
and U3953 (N_3953,N_2052,N_1947);
nor U3954 (N_3954,N_677,N_286);
or U3955 (N_3955,N_1082,N_1771);
or U3956 (N_3956,N_720,N_2038);
or U3957 (N_3957,N_1994,N_238);
or U3958 (N_3958,N_1900,N_2314);
and U3959 (N_3959,N_1866,N_2353);
and U3960 (N_3960,N_1930,N_38);
or U3961 (N_3961,N_2096,N_1585);
or U3962 (N_3962,N_2470,N_2103);
xor U3963 (N_3963,N_2310,N_1170);
nand U3964 (N_3964,N_429,N_923);
and U3965 (N_3965,N_1041,N_1957);
and U3966 (N_3966,N_2016,N_2038);
and U3967 (N_3967,N_2466,N_1917);
and U3968 (N_3968,N_69,N_142);
nor U3969 (N_3969,N_2287,N_526);
and U3970 (N_3970,N_401,N_151);
nor U3971 (N_3971,N_483,N_209);
or U3972 (N_3972,N_880,N_1444);
or U3973 (N_3973,N_227,N_370);
nand U3974 (N_3974,N_2076,N_1402);
nor U3975 (N_3975,N_1197,N_783);
or U3976 (N_3976,N_2388,N_267);
nor U3977 (N_3977,N_404,N_2220);
or U3978 (N_3978,N_1788,N_1237);
or U3979 (N_3979,N_2215,N_2138);
nand U3980 (N_3980,N_544,N_26);
or U3981 (N_3981,N_1844,N_2232);
and U3982 (N_3982,N_520,N_633);
nor U3983 (N_3983,N_704,N_1617);
nand U3984 (N_3984,N_736,N_1754);
nor U3985 (N_3985,N_407,N_1580);
nand U3986 (N_3986,N_924,N_1629);
or U3987 (N_3987,N_1826,N_2078);
nor U3988 (N_3988,N_18,N_1937);
nor U3989 (N_3989,N_1445,N_422);
nand U3990 (N_3990,N_591,N_1958);
or U3991 (N_3991,N_577,N_2304);
nand U3992 (N_3992,N_399,N_1626);
or U3993 (N_3993,N_295,N_419);
or U3994 (N_3994,N_55,N_1180);
and U3995 (N_3995,N_2229,N_1160);
or U3996 (N_3996,N_710,N_830);
xor U3997 (N_3997,N_2381,N_225);
nand U3998 (N_3998,N_2353,N_1492);
and U3999 (N_3999,N_943,N_1287);
and U4000 (N_4000,N_2449,N_1557);
nand U4001 (N_4001,N_2261,N_14);
and U4002 (N_4002,N_2019,N_2169);
nor U4003 (N_4003,N_2336,N_21);
nor U4004 (N_4004,N_1256,N_649);
and U4005 (N_4005,N_1053,N_564);
nand U4006 (N_4006,N_1596,N_339);
and U4007 (N_4007,N_2218,N_2335);
and U4008 (N_4008,N_520,N_1239);
nor U4009 (N_4009,N_845,N_246);
nand U4010 (N_4010,N_450,N_1556);
nand U4011 (N_4011,N_1537,N_1982);
and U4012 (N_4012,N_270,N_968);
or U4013 (N_4013,N_898,N_1258);
or U4014 (N_4014,N_2463,N_1490);
and U4015 (N_4015,N_657,N_394);
nand U4016 (N_4016,N_674,N_2375);
nand U4017 (N_4017,N_1232,N_1447);
nor U4018 (N_4018,N_2224,N_758);
nor U4019 (N_4019,N_1262,N_2173);
or U4020 (N_4020,N_242,N_1314);
nor U4021 (N_4021,N_537,N_1377);
or U4022 (N_4022,N_1460,N_1637);
nand U4023 (N_4023,N_375,N_1643);
nand U4024 (N_4024,N_1120,N_1466);
or U4025 (N_4025,N_1919,N_756);
or U4026 (N_4026,N_883,N_2431);
and U4027 (N_4027,N_1259,N_580);
nor U4028 (N_4028,N_889,N_620);
and U4029 (N_4029,N_571,N_2457);
nand U4030 (N_4030,N_1208,N_1111);
nor U4031 (N_4031,N_1219,N_183);
and U4032 (N_4032,N_1231,N_304);
nand U4033 (N_4033,N_919,N_1618);
nor U4034 (N_4034,N_407,N_1897);
or U4035 (N_4035,N_536,N_2096);
or U4036 (N_4036,N_1631,N_1770);
nor U4037 (N_4037,N_2341,N_1814);
nand U4038 (N_4038,N_2406,N_826);
nand U4039 (N_4039,N_374,N_781);
or U4040 (N_4040,N_1101,N_1898);
or U4041 (N_4041,N_2490,N_956);
nor U4042 (N_4042,N_1026,N_715);
or U4043 (N_4043,N_2160,N_1071);
nor U4044 (N_4044,N_2268,N_675);
nand U4045 (N_4045,N_451,N_2331);
nand U4046 (N_4046,N_919,N_742);
or U4047 (N_4047,N_2210,N_1302);
and U4048 (N_4048,N_849,N_1693);
nor U4049 (N_4049,N_864,N_2426);
nand U4050 (N_4050,N_1882,N_982);
or U4051 (N_4051,N_1891,N_1609);
nand U4052 (N_4052,N_646,N_643);
nor U4053 (N_4053,N_1135,N_1182);
or U4054 (N_4054,N_2349,N_980);
and U4055 (N_4055,N_1273,N_1986);
or U4056 (N_4056,N_1816,N_564);
or U4057 (N_4057,N_2453,N_842);
nor U4058 (N_4058,N_1298,N_2432);
and U4059 (N_4059,N_1744,N_2035);
or U4060 (N_4060,N_611,N_744);
and U4061 (N_4061,N_227,N_2256);
or U4062 (N_4062,N_1918,N_2380);
nand U4063 (N_4063,N_1232,N_1502);
nand U4064 (N_4064,N_752,N_1210);
nand U4065 (N_4065,N_1466,N_900);
nor U4066 (N_4066,N_1133,N_1870);
or U4067 (N_4067,N_148,N_1659);
nand U4068 (N_4068,N_1077,N_1568);
nor U4069 (N_4069,N_1467,N_891);
and U4070 (N_4070,N_2080,N_946);
or U4071 (N_4071,N_932,N_156);
nand U4072 (N_4072,N_2054,N_307);
and U4073 (N_4073,N_2413,N_83);
or U4074 (N_4074,N_1878,N_595);
and U4075 (N_4075,N_771,N_2351);
nor U4076 (N_4076,N_343,N_899);
and U4077 (N_4077,N_1075,N_1492);
nand U4078 (N_4078,N_929,N_1973);
or U4079 (N_4079,N_2444,N_1585);
nand U4080 (N_4080,N_2361,N_1442);
nor U4081 (N_4081,N_550,N_1808);
nor U4082 (N_4082,N_2460,N_2200);
or U4083 (N_4083,N_1874,N_1070);
or U4084 (N_4084,N_2099,N_617);
nand U4085 (N_4085,N_1963,N_2462);
nor U4086 (N_4086,N_1871,N_1995);
and U4087 (N_4087,N_699,N_163);
nor U4088 (N_4088,N_2418,N_273);
and U4089 (N_4089,N_1571,N_983);
or U4090 (N_4090,N_611,N_2437);
nand U4091 (N_4091,N_391,N_780);
and U4092 (N_4092,N_2197,N_1813);
or U4093 (N_4093,N_520,N_1523);
nand U4094 (N_4094,N_344,N_469);
and U4095 (N_4095,N_1921,N_159);
and U4096 (N_4096,N_1933,N_986);
nor U4097 (N_4097,N_994,N_2170);
nor U4098 (N_4098,N_1309,N_2435);
nor U4099 (N_4099,N_2351,N_1771);
nand U4100 (N_4100,N_2248,N_1267);
nand U4101 (N_4101,N_2226,N_1915);
nor U4102 (N_4102,N_726,N_392);
and U4103 (N_4103,N_967,N_467);
nand U4104 (N_4104,N_911,N_1727);
and U4105 (N_4105,N_622,N_1900);
nand U4106 (N_4106,N_1279,N_1465);
nand U4107 (N_4107,N_518,N_1795);
and U4108 (N_4108,N_1926,N_1136);
nor U4109 (N_4109,N_2490,N_360);
and U4110 (N_4110,N_1426,N_1013);
nor U4111 (N_4111,N_239,N_1595);
or U4112 (N_4112,N_1603,N_1691);
or U4113 (N_4113,N_229,N_630);
and U4114 (N_4114,N_125,N_105);
and U4115 (N_4115,N_1105,N_995);
or U4116 (N_4116,N_1479,N_837);
nand U4117 (N_4117,N_1973,N_1677);
and U4118 (N_4118,N_1253,N_1480);
nand U4119 (N_4119,N_844,N_221);
nand U4120 (N_4120,N_2373,N_1980);
or U4121 (N_4121,N_484,N_2248);
nand U4122 (N_4122,N_1478,N_902);
nor U4123 (N_4123,N_758,N_2399);
nand U4124 (N_4124,N_1345,N_1962);
nor U4125 (N_4125,N_1283,N_2496);
or U4126 (N_4126,N_2044,N_302);
nand U4127 (N_4127,N_1084,N_1101);
nand U4128 (N_4128,N_2463,N_1542);
nand U4129 (N_4129,N_987,N_1949);
nand U4130 (N_4130,N_567,N_2499);
nor U4131 (N_4131,N_1074,N_299);
nand U4132 (N_4132,N_724,N_1575);
or U4133 (N_4133,N_1257,N_1105);
or U4134 (N_4134,N_822,N_1321);
nor U4135 (N_4135,N_1640,N_70);
nand U4136 (N_4136,N_995,N_1507);
or U4137 (N_4137,N_248,N_402);
nand U4138 (N_4138,N_1785,N_2322);
or U4139 (N_4139,N_1060,N_1524);
nand U4140 (N_4140,N_2306,N_1256);
nand U4141 (N_4141,N_1107,N_2183);
or U4142 (N_4142,N_2486,N_1595);
and U4143 (N_4143,N_1704,N_1333);
nor U4144 (N_4144,N_222,N_811);
nand U4145 (N_4145,N_1951,N_1267);
xor U4146 (N_4146,N_647,N_2103);
nand U4147 (N_4147,N_1545,N_326);
and U4148 (N_4148,N_939,N_883);
or U4149 (N_4149,N_945,N_1108);
nor U4150 (N_4150,N_943,N_1772);
and U4151 (N_4151,N_1317,N_1627);
nor U4152 (N_4152,N_401,N_965);
nor U4153 (N_4153,N_754,N_1911);
or U4154 (N_4154,N_431,N_311);
nand U4155 (N_4155,N_1461,N_2248);
nand U4156 (N_4156,N_1915,N_1582);
nand U4157 (N_4157,N_1792,N_2165);
and U4158 (N_4158,N_710,N_2060);
or U4159 (N_4159,N_1481,N_2131);
or U4160 (N_4160,N_2385,N_349);
and U4161 (N_4161,N_2476,N_2076);
and U4162 (N_4162,N_499,N_1679);
and U4163 (N_4163,N_2306,N_997);
nor U4164 (N_4164,N_944,N_33);
nand U4165 (N_4165,N_106,N_2122);
or U4166 (N_4166,N_1997,N_82);
or U4167 (N_4167,N_833,N_2084);
nor U4168 (N_4168,N_1620,N_1384);
nor U4169 (N_4169,N_1458,N_1998);
or U4170 (N_4170,N_798,N_1040);
nor U4171 (N_4171,N_1622,N_1028);
and U4172 (N_4172,N_1093,N_1813);
nand U4173 (N_4173,N_1274,N_981);
and U4174 (N_4174,N_1520,N_199);
nand U4175 (N_4175,N_2127,N_1205);
nor U4176 (N_4176,N_253,N_991);
or U4177 (N_4177,N_1557,N_299);
nor U4178 (N_4178,N_558,N_2188);
xnor U4179 (N_4179,N_595,N_55);
nor U4180 (N_4180,N_1334,N_1353);
and U4181 (N_4181,N_10,N_388);
nand U4182 (N_4182,N_2239,N_1820);
or U4183 (N_4183,N_246,N_1384);
and U4184 (N_4184,N_113,N_2033);
or U4185 (N_4185,N_828,N_2444);
nor U4186 (N_4186,N_1713,N_613);
xor U4187 (N_4187,N_281,N_522);
and U4188 (N_4188,N_2198,N_863);
or U4189 (N_4189,N_1260,N_759);
or U4190 (N_4190,N_2287,N_2105);
and U4191 (N_4191,N_2248,N_1568);
and U4192 (N_4192,N_1845,N_1240);
nand U4193 (N_4193,N_1638,N_11);
or U4194 (N_4194,N_2034,N_1645);
and U4195 (N_4195,N_1698,N_2499);
and U4196 (N_4196,N_1040,N_298);
and U4197 (N_4197,N_844,N_1761);
and U4198 (N_4198,N_896,N_1898);
nand U4199 (N_4199,N_32,N_507);
and U4200 (N_4200,N_2456,N_857);
or U4201 (N_4201,N_1343,N_2121);
nor U4202 (N_4202,N_1871,N_150);
nand U4203 (N_4203,N_1858,N_97);
nand U4204 (N_4204,N_950,N_2204);
or U4205 (N_4205,N_1841,N_1399);
nor U4206 (N_4206,N_1196,N_291);
or U4207 (N_4207,N_2294,N_1490);
nor U4208 (N_4208,N_1843,N_1678);
or U4209 (N_4209,N_44,N_706);
nand U4210 (N_4210,N_1309,N_2181);
nand U4211 (N_4211,N_2263,N_341);
and U4212 (N_4212,N_937,N_1780);
nor U4213 (N_4213,N_793,N_1393);
and U4214 (N_4214,N_1800,N_357);
nand U4215 (N_4215,N_2023,N_595);
or U4216 (N_4216,N_124,N_1090);
and U4217 (N_4217,N_787,N_2173);
nor U4218 (N_4218,N_1389,N_1844);
nor U4219 (N_4219,N_2046,N_46);
nand U4220 (N_4220,N_1183,N_713);
xnor U4221 (N_4221,N_216,N_259);
nor U4222 (N_4222,N_51,N_999);
and U4223 (N_4223,N_1000,N_989);
or U4224 (N_4224,N_585,N_2331);
nand U4225 (N_4225,N_1260,N_1886);
nand U4226 (N_4226,N_918,N_1940);
or U4227 (N_4227,N_190,N_1592);
or U4228 (N_4228,N_2363,N_1288);
and U4229 (N_4229,N_2293,N_66);
nor U4230 (N_4230,N_86,N_325);
or U4231 (N_4231,N_203,N_745);
or U4232 (N_4232,N_638,N_2286);
and U4233 (N_4233,N_1102,N_2068);
and U4234 (N_4234,N_933,N_2179);
or U4235 (N_4235,N_981,N_348);
or U4236 (N_4236,N_293,N_197);
nand U4237 (N_4237,N_461,N_2091);
or U4238 (N_4238,N_1925,N_1013);
or U4239 (N_4239,N_1877,N_567);
nor U4240 (N_4240,N_1958,N_847);
nand U4241 (N_4241,N_1965,N_106);
and U4242 (N_4242,N_255,N_1115);
nand U4243 (N_4243,N_1223,N_1697);
nor U4244 (N_4244,N_2165,N_677);
or U4245 (N_4245,N_1825,N_2423);
nand U4246 (N_4246,N_2213,N_1764);
or U4247 (N_4247,N_2359,N_1264);
and U4248 (N_4248,N_1138,N_636);
nand U4249 (N_4249,N_1466,N_2409);
or U4250 (N_4250,N_1697,N_1342);
or U4251 (N_4251,N_466,N_610);
or U4252 (N_4252,N_1805,N_859);
or U4253 (N_4253,N_818,N_440);
or U4254 (N_4254,N_1942,N_566);
nor U4255 (N_4255,N_1432,N_742);
and U4256 (N_4256,N_833,N_2117);
or U4257 (N_4257,N_258,N_1757);
and U4258 (N_4258,N_416,N_260);
or U4259 (N_4259,N_285,N_1717);
nand U4260 (N_4260,N_2493,N_167);
or U4261 (N_4261,N_888,N_225);
or U4262 (N_4262,N_1499,N_208);
nor U4263 (N_4263,N_429,N_600);
or U4264 (N_4264,N_2305,N_1736);
or U4265 (N_4265,N_894,N_809);
nand U4266 (N_4266,N_2305,N_146);
and U4267 (N_4267,N_479,N_283);
nand U4268 (N_4268,N_1886,N_68);
nor U4269 (N_4269,N_112,N_80);
nor U4270 (N_4270,N_1042,N_2416);
and U4271 (N_4271,N_864,N_2481);
nor U4272 (N_4272,N_884,N_873);
and U4273 (N_4273,N_1828,N_2420);
or U4274 (N_4274,N_1761,N_1396);
or U4275 (N_4275,N_1355,N_2288);
or U4276 (N_4276,N_627,N_1892);
nand U4277 (N_4277,N_1843,N_292);
nor U4278 (N_4278,N_985,N_2318);
and U4279 (N_4279,N_683,N_1082);
nor U4280 (N_4280,N_1234,N_571);
nand U4281 (N_4281,N_1369,N_476);
nor U4282 (N_4282,N_2191,N_1987);
and U4283 (N_4283,N_1926,N_90);
nand U4284 (N_4284,N_1952,N_975);
nor U4285 (N_4285,N_2110,N_2218);
nor U4286 (N_4286,N_1184,N_6);
and U4287 (N_4287,N_1639,N_1879);
and U4288 (N_4288,N_2164,N_2054);
or U4289 (N_4289,N_2477,N_245);
nor U4290 (N_4290,N_1661,N_1310);
and U4291 (N_4291,N_2091,N_444);
or U4292 (N_4292,N_1904,N_1161);
and U4293 (N_4293,N_655,N_1437);
and U4294 (N_4294,N_613,N_1203);
nand U4295 (N_4295,N_396,N_888);
nor U4296 (N_4296,N_448,N_1735);
or U4297 (N_4297,N_2114,N_2250);
nor U4298 (N_4298,N_112,N_1607);
nor U4299 (N_4299,N_910,N_1432);
or U4300 (N_4300,N_1608,N_454);
nor U4301 (N_4301,N_1828,N_1270);
and U4302 (N_4302,N_1136,N_1382);
or U4303 (N_4303,N_1150,N_930);
nor U4304 (N_4304,N_1643,N_2400);
or U4305 (N_4305,N_1994,N_1138);
nand U4306 (N_4306,N_1083,N_1275);
or U4307 (N_4307,N_970,N_2224);
nand U4308 (N_4308,N_1963,N_2227);
or U4309 (N_4309,N_979,N_459);
nor U4310 (N_4310,N_717,N_1241);
or U4311 (N_4311,N_2474,N_1848);
and U4312 (N_4312,N_1049,N_423);
or U4313 (N_4313,N_944,N_1913);
nand U4314 (N_4314,N_909,N_721);
and U4315 (N_4315,N_1241,N_932);
nor U4316 (N_4316,N_2157,N_2197);
or U4317 (N_4317,N_643,N_31);
or U4318 (N_4318,N_2472,N_423);
nor U4319 (N_4319,N_2107,N_1627);
nand U4320 (N_4320,N_1779,N_1658);
nor U4321 (N_4321,N_384,N_2192);
or U4322 (N_4322,N_1412,N_987);
or U4323 (N_4323,N_4,N_936);
and U4324 (N_4324,N_1113,N_314);
nor U4325 (N_4325,N_588,N_2169);
nand U4326 (N_4326,N_854,N_1025);
or U4327 (N_4327,N_1161,N_2436);
nand U4328 (N_4328,N_832,N_3);
and U4329 (N_4329,N_564,N_379);
and U4330 (N_4330,N_1398,N_3);
nand U4331 (N_4331,N_913,N_1875);
or U4332 (N_4332,N_67,N_1025);
and U4333 (N_4333,N_790,N_2294);
or U4334 (N_4334,N_690,N_1153);
nor U4335 (N_4335,N_1489,N_1385);
and U4336 (N_4336,N_1426,N_1044);
or U4337 (N_4337,N_1008,N_125);
nand U4338 (N_4338,N_1,N_1386);
nor U4339 (N_4339,N_1821,N_881);
nor U4340 (N_4340,N_125,N_1319);
nand U4341 (N_4341,N_470,N_1483);
xnor U4342 (N_4342,N_2320,N_1248);
nand U4343 (N_4343,N_1924,N_1951);
and U4344 (N_4344,N_1583,N_978);
and U4345 (N_4345,N_601,N_2135);
nor U4346 (N_4346,N_88,N_1233);
nand U4347 (N_4347,N_1766,N_509);
nand U4348 (N_4348,N_1922,N_2318);
nor U4349 (N_4349,N_1453,N_1549);
nor U4350 (N_4350,N_1573,N_2003);
and U4351 (N_4351,N_824,N_1560);
nand U4352 (N_4352,N_2157,N_2151);
and U4353 (N_4353,N_658,N_1561);
or U4354 (N_4354,N_1638,N_467);
nor U4355 (N_4355,N_310,N_2124);
or U4356 (N_4356,N_2491,N_1454);
and U4357 (N_4357,N_271,N_996);
and U4358 (N_4358,N_1829,N_1908);
nor U4359 (N_4359,N_744,N_125);
and U4360 (N_4360,N_72,N_92);
nand U4361 (N_4361,N_293,N_478);
nor U4362 (N_4362,N_2068,N_252);
nand U4363 (N_4363,N_1756,N_663);
and U4364 (N_4364,N_1560,N_2058);
or U4365 (N_4365,N_2156,N_2230);
nand U4366 (N_4366,N_1159,N_1939);
or U4367 (N_4367,N_2009,N_509);
and U4368 (N_4368,N_363,N_910);
nor U4369 (N_4369,N_1283,N_2478);
nand U4370 (N_4370,N_198,N_1164);
and U4371 (N_4371,N_1418,N_1187);
nand U4372 (N_4372,N_1981,N_1003);
and U4373 (N_4373,N_1677,N_1862);
nor U4374 (N_4374,N_1953,N_719);
or U4375 (N_4375,N_132,N_340);
nand U4376 (N_4376,N_2162,N_2393);
and U4377 (N_4377,N_2178,N_521);
nor U4378 (N_4378,N_2399,N_760);
or U4379 (N_4379,N_1559,N_2455);
nand U4380 (N_4380,N_859,N_2049);
and U4381 (N_4381,N_2072,N_966);
or U4382 (N_4382,N_1203,N_2026);
nor U4383 (N_4383,N_2484,N_980);
and U4384 (N_4384,N_1714,N_56);
or U4385 (N_4385,N_1746,N_898);
nand U4386 (N_4386,N_175,N_1621);
and U4387 (N_4387,N_1131,N_781);
and U4388 (N_4388,N_848,N_2079);
nand U4389 (N_4389,N_2028,N_1824);
or U4390 (N_4390,N_2090,N_21);
nor U4391 (N_4391,N_2097,N_576);
or U4392 (N_4392,N_104,N_1962);
nand U4393 (N_4393,N_2465,N_1194);
nor U4394 (N_4394,N_700,N_396);
nor U4395 (N_4395,N_291,N_1731);
or U4396 (N_4396,N_1910,N_2015);
or U4397 (N_4397,N_1530,N_1811);
nand U4398 (N_4398,N_2190,N_262);
and U4399 (N_4399,N_1558,N_1519);
or U4400 (N_4400,N_1036,N_1877);
or U4401 (N_4401,N_1627,N_2466);
nand U4402 (N_4402,N_1954,N_2226);
nand U4403 (N_4403,N_248,N_1298);
nor U4404 (N_4404,N_1002,N_1010);
and U4405 (N_4405,N_479,N_698);
nor U4406 (N_4406,N_1737,N_942);
xnor U4407 (N_4407,N_1350,N_584);
and U4408 (N_4408,N_2065,N_1122);
and U4409 (N_4409,N_286,N_1923);
nor U4410 (N_4410,N_1775,N_1072);
nand U4411 (N_4411,N_2336,N_561);
nor U4412 (N_4412,N_2086,N_1187);
or U4413 (N_4413,N_609,N_26);
and U4414 (N_4414,N_9,N_446);
or U4415 (N_4415,N_1176,N_2345);
nor U4416 (N_4416,N_1199,N_1779);
or U4417 (N_4417,N_1140,N_854);
and U4418 (N_4418,N_2102,N_261);
or U4419 (N_4419,N_1028,N_861);
nand U4420 (N_4420,N_124,N_1508);
and U4421 (N_4421,N_774,N_1227);
or U4422 (N_4422,N_1564,N_501);
nor U4423 (N_4423,N_1473,N_429);
and U4424 (N_4424,N_337,N_316);
nor U4425 (N_4425,N_1955,N_472);
and U4426 (N_4426,N_217,N_670);
nand U4427 (N_4427,N_101,N_2442);
and U4428 (N_4428,N_1506,N_2093);
or U4429 (N_4429,N_591,N_1356);
nand U4430 (N_4430,N_1154,N_998);
nor U4431 (N_4431,N_1821,N_859);
nand U4432 (N_4432,N_1986,N_32);
nor U4433 (N_4433,N_1615,N_240);
or U4434 (N_4434,N_990,N_719);
nor U4435 (N_4435,N_972,N_1436);
and U4436 (N_4436,N_180,N_265);
and U4437 (N_4437,N_280,N_284);
nor U4438 (N_4438,N_732,N_244);
nor U4439 (N_4439,N_1354,N_630);
and U4440 (N_4440,N_1700,N_721);
nand U4441 (N_4441,N_1663,N_998);
nor U4442 (N_4442,N_626,N_1138);
or U4443 (N_4443,N_2415,N_124);
and U4444 (N_4444,N_1751,N_2364);
nand U4445 (N_4445,N_1987,N_1888);
or U4446 (N_4446,N_2368,N_2023);
or U4447 (N_4447,N_1832,N_2103);
nor U4448 (N_4448,N_846,N_2221);
nand U4449 (N_4449,N_2226,N_1600);
nand U4450 (N_4450,N_477,N_200);
and U4451 (N_4451,N_2202,N_1748);
nand U4452 (N_4452,N_980,N_1182);
nor U4453 (N_4453,N_1030,N_2058);
nand U4454 (N_4454,N_1111,N_1186);
or U4455 (N_4455,N_2471,N_2376);
nor U4456 (N_4456,N_557,N_1069);
nor U4457 (N_4457,N_1901,N_826);
nand U4458 (N_4458,N_1376,N_1589);
or U4459 (N_4459,N_2459,N_1771);
and U4460 (N_4460,N_2095,N_1784);
nand U4461 (N_4461,N_1864,N_2230);
or U4462 (N_4462,N_7,N_2045);
nor U4463 (N_4463,N_2182,N_1090);
and U4464 (N_4464,N_2331,N_1898);
nor U4465 (N_4465,N_182,N_387);
or U4466 (N_4466,N_621,N_577);
and U4467 (N_4467,N_2429,N_2066);
or U4468 (N_4468,N_1548,N_397);
or U4469 (N_4469,N_1489,N_21);
nor U4470 (N_4470,N_1370,N_2376);
nand U4471 (N_4471,N_590,N_1711);
and U4472 (N_4472,N_1504,N_1526);
nor U4473 (N_4473,N_2042,N_1946);
nand U4474 (N_4474,N_2043,N_305);
and U4475 (N_4475,N_839,N_2388);
nor U4476 (N_4476,N_1603,N_1893);
nor U4477 (N_4477,N_413,N_2429);
xnor U4478 (N_4478,N_1723,N_2084);
and U4479 (N_4479,N_246,N_1383);
or U4480 (N_4480,N_1438,N_1293);
xor U4481 (N_4481,N_629,N_327);
nand U4482 (N_4482,N_963,N_1220);
nor U4483 (N_4483,N_644,N_939);
nor U4484 (N_4484,N_2098,N_760);
nand U4485 (N_4485,N_288,N_791);
nand U4486 (N_4486,N_1824,N_592);
and U4487 (N_4487,N_2497,N_1451);
or U4488 (N_4488,N_1635,N_2360);
or U4489 (N_4489,N_546,N_232);
and U4490 (N_4490,N_1253,N_760);
nand U4491 (N_4491,N_2135,N_32);
nor U4492 (N_4492,N_2092,N_105);
or U4493 (N_4493,N_31,N_163);
nor U4494 (N_4494,N_1716,N_1525);
nor U4495 (N_4495,N_1399,N_292);
and U4496 (N_4496,N_98,N_1144);
nor U4497 (N_4497,N_1945,N_1136);
and U4498 (N_4498,N_2104,N_1232);
and U4499 (N_4499,N_1838,N_1987);
or U4500 (N_4500,N_1214,N_1253);
and U4501 (N_4501,N_13,N_2117);
or U4502 (N_4502,N_2068,N_2353);
and U4503 (N_4503,N_1115,N_1151);
nand U4504 (N_4504,N_2312,N_1122);
and U4505 (N_4505,N_1924,N_948);
and U4506 (N_4506,N_35,N_914);
or U4507 (N_4507,N_1590,N_787);
nand U4508 (N_4508,N_2341,N_1048);
or U4509 (N_4509,N_2382,N_978);
nor U4510 (N_4510,N_1683,N_376);
and U4511 (N_4511,N_1396,N_1991);
nand U4512 (N_4512,N_425,N_320);
nand U4513 (N_4513,N_1281,N_917);
nand U4514 (N_4514,N_78,N_958);
and U4515 (N_4515,N_1584,N_634);
nand U4516 (N_4516,N_913,N_2326);
or U4517 (N_4517,N_1560,N_301);
nand U4518 (N_4518,N_2331,N_843);
nand U4519 (N_4519,N_2116,N_1410);
nand U4520 (N_4520,N_2469,N_678);
and U4521 (N_4521,N_918,N_1929);
or U4522 (N_4522,N_1118,N_2340);
and U4523 (N_4523,N_1375,N_418);
or U4524 (N_4524,N_1198,N_1537);
or U4525 (N_4525,N_771,N_1210);
or U4526 (N_4526,N_2217,N_1982);
nor U4527 (N_4527,N_289,N_816);
and U4528 (N_4528,N_1734,N_1572);
or U4529 (N_4529,N_1366,N_640);
xnor U4530 (N_4530,N_1818,N_2292);
and U4531 (N_4531,N_1650,N_785);
nor U4532 (N_4532,N_2060,N_356);
and U4533 (N_4533,N_2336,N_997);
or U4534 (N_4534,N_53,N_2487);
or U4535 (N_4535,N_1323,N_2374);
or U4536 (N_4536,N_1241,N_651);
nand U4537 (N_4537,N_1143,N_2368);
and U4538 (N_4538,N_117,N_1586);
nand U4539 (N_4539,N_1732,N_468);
nand U4540 (N_4540,N_1609,N_644);
and U4541 (N_4541,N_646,N_491);
xnor U4542 (N_4542,N_684,N_1524);
nand U4543 (N_4543,N_1039,N_617);
or U4544 (N_4544,N_1023,N_438);
or U4545 (N_4545,N_497,N_1929);
nand U4546 (N_4546,N_1557,N_1537);
or U4547 (N_4547,N_1349,N_2352);
nand U4548 (N_4548,N_1621,N_1609);
and U4549 (N_4549,N_1721,N_63);
nor U4550 (N_4550,N_417,N_2041);
or U4551 (N_4551,N_2487,N_2292);
or U4552 (N_4552,N_1210,N_162);
nor U4553 (N_4553,N_1040,N_1795);
nor U4554 (N_4554,N_1528,N_1921);
and U4555 (N_4555,N_225,N_796);
or U4556 (N_4556,N_2051,N_2249);
nand U4557 (N_4557,N_696,N_2480);
nor U4558 (N_4558,N_1678,N_2477);
nor U4559 (N_4559,N_12,N_1258);
or U4560 (N_4560,N_1704,N_1899);
and U4561 (N_4561,N_1463,N_1352);
or U4562 (N_4562,N_12,N_156);
or U4563 (N_4563,N_1048,N_1418);
and U4564 (N_4564,N_1530,N_445);
and U4565 (N_4565,N_457,N_2155);
nor U4566 (N_4566,N_2349,N_1836);
or U4567 (N_4567,N_106,N_1151);
nand U4568 (N_4568,N_1963,N_274);
nor U4569 (N_4569,N_2324,N_785);
nand U4570 (N_4570,N_121,N_180);
nand U4571 (N_4571,N_1739,N_164);
or U4572 (N_4572,N_656,N_191);
or U4573 (N_4573,N_201,N_1925);
xnor U4574 (N_4574,N_502,N_2471);
nor U4575 (N_4575,N_1767,N_1009);
and U4576 (N_4576,N_2179,N_564);
or U4577 (N_4577,N_396,N_1026);
and U4578 (N_4578,N_459,N_2064);
nand U4579 (N_4579,N_634,N_453);
nand U4580 (N_4580,N_119,N_583);
nand U4581 (N_4581,N_885,N_1095);
or U4582 (N_4582,N_157,N_1380);
nand U4583 (N_4583,N_1284,N_2069);
nand U4584 (N_4584,N_1965,N_990);
and U4585 (N_4585,N_2072,N_946);
and U4586 (N_4586,N_371,N_594);
nand U4587 (N_4587,N_1649,N_39);
nand U4588 (N_4588,N_2284,N_2027);
or U4589 (N_4589,N_408,N_855);
and U4590 (N_4590,N_710,N_1529);
or U4591 (N_4591,N_1071,N_1880);
or U4592 (N_4592,N_331,N_1703);
nor U4593 (N_4593,N_1318,N_2064);
nand U4594 (N_4594,N_1238,N_1691);
or U4595 (N_4595,N_379,N_691);
nor U4596 (N_4596,N_420,N_1887);
or U4597 (N_4597,N_603,N_1536);
nor U4598 (N_4598,N_2051,N_705);
and U4599 (N_4599,N_1174,N_1126);
nor U4600 (N_4600,N_1385,N_1611);
or U4601 (N_4601,N_399,N_2204);
and U4602 (N_4602,N_311,N_149);
nor U4603 (N_4603,N_414,N_1736);
and U4604 (N_4604,N_1401,N_1149);
and U4605 (N_4605,N_904,N_1667);
nor U4606 (N_4606,N_737,N_286);
or U4607 (N_4607,N_151,N_2483);
or U4608 (N_4608,N_1927,N_2146);
nor U4609 (N_4609,N_1788,N_2466);
nand U4610 (N_4610,N_1469,N_629);
nand U4611 (N_4611,N_388,N_1339);
nor U4612 (N_4612,N_1242,N_2389);
nor U4613 (N_4613,N_2242,N_1857);
and U4614 (N_4614,N_2314,N_2009);
and U4615 (N_4615,N_638,N_2040);
nor U4616 (N_4616,N_1040,N_2297);
nand U4617 (N_4617,N_822,N_935);
nand U4618 (N_4618,N_1655,N_1920);
nand U4619 (N_4619,N_819,N_1353);
nor U4620 (N_4620,N_40,N_2164);
nor U4621 (N_4621,N_1927,N_1151);
and U4622 (N_4622,N_543,N_621);
nand U4623 (N_4623,N_2222,N_1528);
and U4624 (N_4624,N_2400,N_1327);
nand U4625 (N_4625,N_2428,N_12);
and U4626 (N_4626,N_1111,N_1001);
nor U4627 (N_4627,N_469,N_1407);
nor U4628 (N_4628,N_1030,N_0);
nand U4629 (N_4629,N_2206,N_335);
or U4630 (N_4630,N_447,N_2338);
and U4631 (N_4631,N_623,N_1075);
nand U4632 (N_4632,N_835,N_606);
nor U4633 (N_4633,N_2471,N_1705);
and U4634 (N_4634,N_684,N_1578);
nor U4635 (N_4635,N_673,N_52);
nor U4636 (N_4636,N_1822,N_2032);
nand U4637 (N_4637,N_876,N_1022);
or U4638 (N_4638,N_1348,N_586);
nand U4639 (N_4639,N_1809,N_363);
and U4640 (N_4640,N_1232,N_1476);
nand U4641 (N_4641,N_2077,N_965);
and U4642 (N_4642,N_1844,N_2273);
or U4643 (N_4643,N_1748,N_2377);
nand U4644 (N_4644,N_405,N_1681);
and U4645 (N_4645,N_355,N_1523);
or U4646 (N_4646,N_1706,N_1177);
nor U4647 (N_4647,N_1096,N_225);
nor U4648 (N_4648,N_565,N_1832);
nor U4649 (N_4649,N_1397,N_807);
nand U4650 (N_4650,N_322,N_2457);
nand U4651 (N_4651,N_2155,N_1160);
nand U4652 (N_4652,N_2097,N_1851);
or U4653 (N_4653,N_915,N_1984);
nand U4654 (N_4654,N_418,N_1690);
or U4655 (N_4655,N_398,N_2409);
or U4656 (N_4656,N_1160,N_1974);
nor U4657 (N_4657,N_565,N_2007);
or U4658 (N_4658,N_1409,N_713);
or U4659 (N_4659,N_1299,N_2176);
nor U4660 (N_4660,N_1698,N_1054);
and U4661 (N_4661,N_1932,N_1335);
nor U4662 (N_4662,N_2452,N_132);
or U4663 (N_4663,N_2187,N_1853);
or U4664 (N_4664,N_222,N_164);
or U4665 (N_4665,N_2287,N_1810);
or U4666 (N_4666,N_31,N_2372);
and U4667 (N_4667,N_2222,N_263);
nand U4668 (N_4668,N_257,N_748);
or U4669 (N_4669,N_2013,N_2050);
or U4670 (N_4670,N_833,N_959);
nand U4671 (N_4671,N_600,N_2038);
nand U4672 (N_4672,N_1003,N_945);
and U4673 (N_4673,N_1994,N_395);
and U4674 (N_4674,N_951,N_1753);
nand U4675 (N_4675,N_125,N_2303);
nand U4676 (N_4676,N_2219,N_819);
nor U4677 (N_4677,N_93,N_826);
nand U4678 (N_4678,N_307,N_1317);
nor U4679 (N_4679,N_1778,N_2217);
nand U4680 (N_4680,N_2084,N_1683);
nand U4681 (N_4681,N_1924,N_550);
nand U4682 (N_4682,N_1829,N_2296);
and U4683 (N_4683,N_2004,N_1270);
nand U4684 (N_4684,N_806,N_290);
nor U4685 (N_4685,N_2361,N_1305);
and U4686 (N_4686,N_931,N_848);
and U4687 (N_4687,N_1344,N_1229);
nor U4688 (N_4688,N_716,N_2331);
and U4689 (N_4689,N_870,N_960);
or U4690 (N_4690,N_1548,N_494);
nand U4691 (N_4691,N_1589,N_2260);
and U4692 (N_4692,N_1334,N_637);
and U4693 (N_4693,N_440,N_696);
nand U4694 (N_4694,N_59,N_490);
nor U4695 (N_4695,N_1710,N_100);
nand U4696 (N_4696,N_2186,N_140);
and U4697 (N_4697,N_1011,N_2421);
nor U4698 (N_4698,N_2384,N_1490);
and U4699 (N_4699,N_2400,N_1705);
and U4700 (N_4700,N_1856,N_612);
nor U4701 (N_4701,N_2178,N_216);
or U4702 (N_4702,N_1977,N_1566);
and U4703 (N_4703,N_2371,N_60);
nor U4704 (N_4704,N_322,N_531);
or U4705 (N_4705,N_1277,N_1886);
nand U4706 (N_4706,N_835,N_802);
nand U4707 (N_4707,N_1773,N_642);
nand U4708 (N_4708,N_900,N_798);
and U4709 (N_4709,N_1673,N_2110);
or U4710 (N_4710,N_195,N_225);
nor U4711 (N_4711,N_1010,N_2091);
nor U4712 (N_4712,N_1899,N_437);
nand U4713 (N_4713,N_1575,N_701);
nand U4714 (N_4714,N_1451,N_1038);
and U4715 (N_4715,N_2472,N_1086);
or U4716 (N_4716,N_1807,N_799);
nor U4717 (N_4717,N_1180,N_1290);
nand U4718 (N_4718,N_232,N_1781);
or U4719 (N_4719,N_765,N_99);
or U4720 (N_4720,N_788,N_1753);
and U4721 (N_4721,N_1162,N_1880);
nand U4722 (N_4722,N_406,N_1694);
and U4723 (N_4723,N_10,N_1391);
or U4724 (N_4724,N_751,N_793);
and U4725 (N_4725,N_1439,N_1617);
nand U4726 (N_4726,N_354,N_1764);
nor U4727 (N_4727,N_2462,N_1876);
or U4728 (N_4728,N_2190,N_2457);
nor U4729 (N_4729,N_2093,N_2032);
nand U4730 (N_4730,N_1521,N_1712);
or U4731 (N_4731,N_2499,N_363);
or U4732 (N_4732,N_1445,N_428);
or U4733 (N_4733,N_1052,N_2261);
and U4734 (N_4734,N_1822,N_887);
and U4735 (N_4735,N_1288,N_755);
or U4736 (N_4736,N_257,N_2074);
and U4737 (N_4737,N_2361,N_1855);
or U4738 (N_4738,N_2207,N_1639);
or U4739 (N_4739,N_2440,N_2042);
and U4740 (N_4740,N_842,N_214);
nand U4741 (N_4741,N_372,N_680);
nor U4742 (N_4742,N_467,N_35);
and U4743 (N_4743,N_194,N_2454);
and U4744 (N_4744,N_108,N_2012);
or U4745 (N_4745,N_2223,N_1077);
nor U4746 (N_4746,N_953,N_350);
nor U4747 (N_4747,N_670,N_2281);
nand U4748 (N_4748,N_47,N_2291);
or U4749 (N_4749,N_205,N_1291);
or U4750 (N_4750,N_863,N_1102);
nor U4751 (N_4751,N_1090,N_1653);
nor U4752 (N_4752,N_799,N_1053);
or U4753 (N_4753,N_1961,N_2016);
or U4754 (N_4754,N_560,N_1474);
or U4755 (N_4755,N_1127,N_261);
or U4756 (N_4756,N_1908,N_240);
nor U4757 (N_4757,N_1661,N_336);
nor U4758 (N_4758,N_1928,N_2086);
and U4759 (N_4759,N_1742,N_468);
nand U4760 (N_4760,N_230,N_294);
or U4761 (N_4761,N_1210,N_2302);
nand U4762 (N_4762,N_1056,N_1433);
and U4763 (N_4763,N_1607,N_1524);
and U4764 (N_4764,N_1394,N_1642);
and U4765 (N_4765,N_1320,N_60);
nor U4766 (N_4766,N_1568,N_265);
nor U4767 (N_4767,N_1983,N_2397);
nand U4768 (N_4768,N_697,N_875);
and U4769 (N_4769,N_1255,N_1829);
nor U4770 (N_4770,N_2182,N_557);
nor U4771 (N_4771,N_2276,N_9);
nand U4772 (N_4772,N_999,N_747);
nor U4773 (N_4773,N_286,N_1066);
and U4774 (N_4774,N_1096,N_2005);
or U4775 (N_4775,N_1429,N_2369);
and U4776 (N_4776,N_744,N_351);
or U4777 (N_4777,N_655,N_2211);
nand U4778 (N_4778,N_1840,N_256);
or U4779 (N_4779,N_1293,N_1250);
nand U4780 (N_4780,N_669,N_80);
nand U4781 (N_4781,N_1380,N_1868);
nand U4782 (N_4782,N_1116,N_459);
and U4783 (N_4783,N_1833,N_2113);
nor U4784 (N_4784,N_676,N_747);
and U4785 (N_4785,N_252,N_198);
nor U4786 (N_4786,N_2110,N_1346);
and U4787 (N_4787,N_1397,N_815);
or U4788 (N_4788,N_156,N_1709);
nor U4789 (N_4789,N_1092,N_99);
nand U4790 (N_4790,N_1938,N_768);
nor U4791 (N_4791,N_804,N_2173);
xor U4792 (N_4792,N_278,N_1994);
nor U4793 (N_4793,N_1355,N_883);
or U4794 (N_4794,N_277,N_1293);
nand U4795 (N_4795,N_391,N_2426);
nand U4796 (N_4796,N_893,N_2413);
nand U4797 (N_4797,N_495,N_1856);
and U4798 (N_4798,N_563,N_2427);
nand U4799 (N_4799,N_236,N_377);
nand U4800 (N_4800,N_924,N_1423);
and U4801 (N_4801,N_2042,N_2373);
nand U4802 (N_4802,N_269,N_48);
nand U4803 (N_4803,N_362,N_1165);
and U4804 (N_4804,N_1783,N_1874);
or U4805 (N_4805,N_2416,N_1722);
nand U4806 (N_4806,N_2311,N_1960);
and U4807 (N_4807,N_2348,N_1512);
and U4808 (N_4808,N_1365,N_962);
nor U4809 (N_4809,N_1569,N_753);
nor U4810 (N_4810,N_2126,N_2175);
or U4811 (N_4811,N_1191,N_1180);
nand U4812 (N_4812,N_1274,N_847);
or U4813 (N_4813,N_649,N_1940);
nor U4814 (N_4814,N_1752,N_899);
nand U4815 (N_4815,N_1148,N_51);
nor U4816 (N_4816,N_1899,N_111);
and U4817 (N_4817,N_154,N_1019);
or U4818 (N_4818,N_2151,N_857);
and U4819 (N_4819,N_656,N_401);
nand U4820 (N_4820,N_1760,N_232);
nor U4821 (N_4821,N_1324,N_1420);
nor U4822 (N_4822,N_2127,N_1020);
nor U4823 (N_4823,N_709,N_1981);
nor U4824 (N_4824,N_1293,N_990);
nor U4825 (N_4825,N_1179,N_1998);
or U4826 (N_4826,N_716,N_12);
or U4827 (N_4827,N_500,N_395);
and U4828 (N_4828,N_1050,N_1173);
nor U4829 (N_4829,N_173,N_2149);
and U4830 (N_4830,N_1216,N_729);
nor U4831 (N_4831,N_1228,N_163);
nor U4832 (N_4832,N_1006,N_409);
or U4833 (N_4833,N_2,N_578);
nand U4834 (N_4834,N_1912,N_1240);
nand U4835 (N_4835,N_733,N_866);
and U4836 (N_4836,N_137,N_309);
nand U4837 (N_4837,N_1291,N_335);
and U4838 (N_4838,N_2490,N_2377);
nor U4839 (N_4839,N_2424,N_759);
and U4840 (N_4840,N_153,N_289);
or U4841 (N_4841,N_556,N_376);
nor U4842 (N_4842,N_1623,N_1332);
and U4843 (N_4843,N_1857,N_1009);
or U4844 (N_4844,N_1396,N_1970);
nand U4845 (N_4845,N_2212,N_664);
nor U4846 (N_4846,N_1120,N_2037);
or U4847 (N_4847,N_1279,N_816);
or U4848 (N_4848,N_1341,N_371);
or U4849 (N_4849,N_1638,N_1149);
and U4850 (N_4850,N_752,N_625);
or U4851 (N_4851,N_2463,N_1193);
or U4852 (N_4852,N_1352,N_1551);
or U4853 (N_4853,N_483,N_1910);
nand U4854 (N_4854,N_528,N_1834);
nor U4855 (N_4855,N_644,N_2405);
or U4856 (N_4856,N_1928,N_2436);
and U4857 (N_4857,N_132,N_1062);
nand U4858 (N_4858,N_2426,N_748);
and U4859 (N_4859,N_27,N_390);
nand U4860 (N_4860,N_352,N_1412);
or U4861 (N_4861,N_1206,N_503);
xnor U4862 (N_4862,N_821,N_2479);
nor U4863 (N_4863,N_1405,N_905);
nor U4864 (N_4864,N_1428,N_2094);
or U4865 (N_4865,N_1440,N_2479);
nor U4866 (N_4866,N_2243,N_886);
nand U4867 (N_4867,N_804,N_1970);
and U4868 (N_4868,N_1608,N_1838);
nand U4869 (N_4869,N_65,N_2236);
nor U4870 (N_4870,N_2030,N_923);
or U4871 (N_4871,N_300,N_2089);
nand U4872 (N_4872,N_585,N_1160);
nand U4873 (N_4873,N_1318,N_1259);
nor U4874 (N_4874,N_227,N_1930);
or U4875 (N_4875,N_66,N_525);
or U4876 (N_4876,N_2042,N_1178);
nand U4877 (N_4877,N_51,N_1373);
or U4878 (N_4878,N_2445,N_247);
or U4879 (N_4879,N_1320,N_2039);
nor U4880 (N_4880,N_660,N_2399);
and U4881 (N_4881,N_1153,N_2446);
nand U4882 (N_4882,N_486,N_431);
and U4883 (N_4883,N_770,N_840);
nand U4884 (N_4884,N_188,N_1463);
and U4885 (N_4885,N_894,N_701);
or U4886 (N_4886,N_1657,N_1287);
and U4887 (N_4887,N_1112,N_1234);
or U4888 (N_4888,N_235,N_1151);
or U4889 (N_4889,N_234,N_2229);
nor U4890 (N_4890,N_2239,N_731);
nor U4891 (N_4891,N_2016,N_772);
nor U4892 (N_4892,N_1624,N_1868);
or U4893 (N_4893,N_1713,N_2142);
or U4894 (N_4894,N_610,N_2000);
nor U4895 (N_4895,N_1391,N_35);
or U4896 (N_4896,N_8,N_1786);
nor U4897 (N_4897,N_1702,N_1350);
and U4898 (N_4898,N_1592,N_1612);
nand U4899 (N_4899,N_1732,N_76);
nor U4900 (N_4900,N_793,N_1342);
and U4901 (N_4901,N_1461,N_1894);
and U4902 (N_4902,N_1448,N_2356);
and U4903 (N_4903,N_454,N_1178);
xor U4904 (N_4904,N_1650,N_283);
xnor U4905 (N_4905,N_73,N_893);
nand U4906 (N_4906,N_1300,N_562);
nor U4907 (N_4907,N_149,N_842);
or U4908 (N_4908,N_150,N_2370);
nand U4909 (N_4909,N_2103,N_1480);
or U4910 (N_4910,N_1634,N_2469);
and U4911 (N_4911,N_1577,N_503);
and U4912 (N_4912,N_2072,N_2185);
and U4913 (N_4913,N_435,N_1261);
nor U4914 (N_4914,N_1085,N_2193);
nand U4915 (N_4915,N_377,N_1557);
and U4916 (N_4916,N_508,N_1940);
nor U4917 (N_4917,N_2193,N_312);
or U4918 (N_4918,N_1278,N_875);
nor U4919 (N_4919,N_1154,N_1055);
nor U4920 (N_4920,N_539,N_2493);
nand U4921 (N_4921,N_2491,N_712);
or U4922 (N_4922,N_991,N_2234);
and U4923 (N_4923,N_1003,N_1528);
or U4924 (N_4924,N_966,N_2300);
nand U4925 (N_4925,N_822,N_2180);
and U4926 (N_4926,N_563,N_1156);
nor U4927 (N_4927,N_1088,N_1984);
and U4928 (N_4928,N_1197,N_1556);
and U4929 (N_4929,N_625,N_796);
nand U4930 (N_4930,N_1201,N_1659);
and U4931 (N_4931,N_1442,N_2444);
nand U4932 (N_4932,N_1498,N_300);
and U4933 (N_4933,N_2094,N_2169);
or U4934 (N_4934,N_2304,N_90);
nand U4935 (N_4935,N_1619,N_1738);
nor U4936 (N_4936,N_869,N_1118);
nand U4937 (N_4937,N_2092,N_800);
nor U4938 (N_4938,N_2444,N_202);
or U4939 (N_4939,N_1277,N_2360);
and U4940 (N_4940,N_57,N_2194);
or U4941 (N_4941,N_1683,N_465);
nand U4942 (N_4942,N_1345,N_1681);
and U4943 (N_4943,N_1284,N_2470);
nor U4944 (N_4944,N_1165,N_1621);
or U4945 (N_4945,N_856,N_1438);
or U4946 (N_4946,N_410,N_669);
nor U4947 (N_4947,N_1298,N_972);
nand U4948 (N_4948,N_739,N_2308);
nand U4949 (N_4949,N_349,N_314);
or U4950 (N_4950,N_1567,N_274);
and U4951 (N_4951,N_2106,N_1852);
nor U4952 (N_4952,N_1171,N_337);
nand U4953 (N_4953,N_1629,N_832);
nor U4954 (N_4954,N_1203,N_520);
or U4955 (N_4955,N_1451,N_724);
nor U4956 (N_4956,N_577,N_521);
nor U4957 (N_4957,N_2418,N_1522);
or U4958 (N_4958,N_2100,N_422);
nand U4959 (N_4959,N_792,N_1754);
nor U4960 (N_4960,N_73,N_1251);
or U4961 (N_4961,N_168,N_301);
and U4962 (N_4962,N_1232,N_1655);
and U4963 (N_4963,N_1226,N_815);
and U4964 (N_4964,N_1063,N_1255);
nand U4965 (N_4965,N_1143,N_1507);
and U4966 (N_4966,N_1694,N_2026);
nand U4967 (N_4967,N_2499,N_1892);
nor U4968 (N_4968,N_885,N_734);
nor U4969 (N_4969,N_2094,N_2036);
and U4970 (N_4970,N_950,N_1533);
nor U4971 (N_4971,N_1916,N_1348);
nor U4972 (N_4972,N_1460,N_2412);
or U4973 (N_4973,N_1399,N_1132);
nand U4974 (N_4974,N_147,N_143);
nand U4975 (N_4975,N_2031,N_1455);
nor U4976 (N_4976,N_2121,N_2153);
nand U4977 (N_4977,N_188,N_1310);
nand U4978 (N_4978,N_837,N_38);
nor U4979 (N_4979,N_1195,N_642);
nor U4980 (N_4980,N_1067,N_2362);
or U4981 (N_4981,N_2095,N_116);
nor U4982 (N_4982,N_1372,N_67);
or U4983 (N_4983,N_1792,N_807);
and U4984 (N_4984,N_2372,N_1272);
or U4985 (N_4985,N_1900,N_1512);
nand U4986 (N_4986,N_1038,N_2320);
or U4987 (N_4987,N_241,N_2299);
and U4988 (N_4988,N_634,N_955);
or U4989 (N_4989,N_2297,N_1519);
nand U4990 (N_4990,N_1999,N_537);
and U4991 (N_4991,N_939,N_663);
or U4992 (N_4992,N_2275,N_244);
or U4993 (N_4993,N_1111,N_605);
nand U4994 (N_4994,N_29,N_237);
and U4995 (N_4995,N_1412,N_2434);
and U4996 (N_4996,N_1760,N_2302);
nand U4997 (N_4997,N_321,N_2028);
nand U4998 (N_4998,N_64,N_1259);
and U4999 (N_4999,N_723,N_2232);
nand UO_0 (O_0,N_4080,N_3841);
nand UO_1 (O_1,N_2625,N_3710);
nor UO_2 (O_2,N_4269,N_4583);
nor UO_3 (O_3,N_2507,N_3644);
or UO_4 (O_4,N_3804,N_4564);
nor UO_5 (O_5,N_4664,N_4549);
or UO_6 (O_6,N_3747,N_4657);
nand UO_7 (O_7,N_4576,N_4753);
nand UO_8 (O_8,N_3491,N_4963);
or UO_9 (O_9,N_3611,N_4676);
and UO_10 (O_10,N_3879,N_3248);
nand UO_11 (O_11,N_3893,N_4422);
and UO_12 (O_12,N_4369,N_2954);
nand UO_13 (O_13,N_4988,N_3303);
nand UO_14 (O_14,N_4058,N_4671);
nand UO_15 (O_15,N_2675,N_2980);
nor UO_16 (O_16,N_3053,N_3913);
nand UO_17 (O_17,N_4218,N_3363);
and UO_18 (O_18,N_4955,N_2944);
nand UO_19 (O_19,N_2732,N_4613);
or UO_20 (O_20,N_4112,N_4870);
nand UO_21 (O_21,N_3267,N_4879);
nor UO_22 (O_22,N_4293,N_2901);
nand UO_23 (O_23,N_3471,N_2882);
nor UO_24 (O_24,N_3726,N_4352);
and UO_25 (O_25,N_3230,N_3135);
nor UO_26 (O_26,N_3353,N_4244);
or UO_27 (O_27,N_3950,N_3348);
nand UO_28 (O_28,N_4105,N_4783);
or UO_29 (O_29,N_4641,N_2928);
and UO_30 (O_30,N_4715,N_4891);
and UO_31 (O_31,N_3555,N_4979);
or UO_32 (O_32,N_4277,N_4554);
nand UO_33 (O_33,N_3826,N_4805);
and UO_34 (O_34,N_3497,N_3049);
and UO_35 (O_35,N_3408,N_3423);
nand UO_36 (O_36,N_3101,N_2547);
nor UO_37 (O_37,N_2829,N_4827);
and UO_38 (O_38,N_2966,N_3270);
nand UO_39 (O_39,N_4441,N_3444);
or UO_40 (O_40,N_4268,N_3823);
or UO_41 (O_41,N_2607,N_4832);
nor UO_42 (O_42,N_3144,N_4781);
xnor UO_43 (O_43,N_4969,N_3265);
nor UO_44 (O_44,N_3551,N_2649);
nor UO_45 (O_45,N_3006,N_4308);
nand UO_46 (O_46,N_2674,N_4651);
and UO_47 (O_47,N_2932,N_4221);
and UO_48 (O_48,N_2704,N_4959);
nand UO_49 (O_49,N_4289,N_2616);
and UO_50 (O_50,N_3852,N_2773);
and UO_51 (O_51,N_4329,N_3050);
nor UO_52 (O_52,N_2924,N_4019);
nor UO_53 (O_53,N_4724,N_3436);
and UO_54 (O_54,N_2981,N_2782);
nand UO_55 (O_55,N_4767,N_2650);
and UO_56 (O_56,N_4201,N_4663);
nand UO_57 (O_57,N_4039,N_3920);
nor UO_58 (O_58,N_3309,N_3389);
and UO_59 (O_59,N_3732,N_2852);
nor UO_60 (O_60,N_2589,N_4726);
nand UO_61 (O_61,N_3880,N_4187);
or UO_62 (O_62,N_3662,N_2819);
or UO_63 (O_63,N_4932,N_4883);
xor UO_64 (O_64,N_4947,N_3717);
nor UO_65 (O_65,N_3973,N_3794);
nor UO_66 (O_66,N_3818,N_3466);
nand UO_67 (O_67,N_2731,N_2703);
and UO_68 (O_68,N_4113,N_3928);
and UO_69 (O_69,N_4319,N_4785);
and UO_70 (O_70,N_4371,N_2525);
nor UO_71 (O_71,N_3882,N_2824);
nand UO_72 (O_72,N_2919,N_2835);
and UO_73 (O_73,N_3399,N_3148);
and UO_74 (O_74,N_2569,N_2548);
nand UO_75 (O_75,N_3979,N_3812);
and UO_76 (O_76,N_3917,N_3001);
nand UO_77 (O_77,N_4440,N_2777);
nor UO_78 (O_78,N_4594,N_4779);
nor UO_79 (O_79,N_3697,N_3220);
nand UO_80 (O_80,N_4706,N_3429);
and UO_81 (O_81,N_2620,N_3617);
nor UO_82 (O_82,N_3250,N_3520);
nor UO_83 (O_83,N_4833,N_4603);
nand UO_84 (O_84,N_3825,N_3218);
and UO_85 (O_85,N_4235,N_2791);
or UO_86 (O_86,N_3881,N_3819);
and UO_87 (O_87,N_3528,N_4001);
and UO_88 (O_88,N_2770,N_3264);
or UO_89 (O_89,N_2979,N_2694);
nor UO_90 (O_90,N_4752,N_3407);
or UO_91 (O_91,N_3039,N_4200);
nand UO_92 (O_92,N_2817,N_4614);
nor UO_93 (O_93,N_4630,N_2603);
or UO_94 (O_94,N_3482,N_3495);
or UO_95 (O_95,N_3022,N_3426);
or UO_96 (O_96,N_4669,N_4341);
nor UO_97 (O_97,N_4881,N_3015);
and UO_98 (O_98,N_3573,N_3569);
and UO_99 (O_99,N_4210,N_3134);
nor UO_100 (O_100,N_2858,N_2804);
nand UO_101 (O_101,N_3319,N_3074);
nand UO_102 (O_102,N_3425,N_4089);
nand UO_103 (O_103,N_3963,N_4294);
or UO_104 (O_104,N_2952,N_3875);
and UO_105 (O_105,N_3775,N_3061);
nand UO_106 (O_106,N_3970,N_3923);
and UO_107 (O_107,N_3978,N_4658);
or UO_108 (O_108,N_3318,N_4342);
or UO_109 (O_109,N_3051,N_4976);
or UO_110 (O_110,N_2526,N_4683);
nand UO_111 (O_111,N_4184,N_3308);
and UO_112 (O_112,N_2628,N_4751);
nor UO_113 (O_113,N_3713,N_2577);
and UO_114 (O_114,N_4364,N_3412);
nor UO_115 (O_115,N_3900,N_4954);
or UO_116 (O_116,N_3846,N_2629);
and UO_117 (O_117,N_3515,N_3162);
nand UO_118 (O_118,N_4729,N_4607);
nand UO_119 (O_119,N_3871,N_3510);
nor UO_120 (O_120,N_3339,N_2502);
nor UO_121 (O_121,N_3208,N_4018);
and UO_122 (O_122,N_4190,N_4445);
nand UO_123 (O_123,N_3373,N_4575);
or UO_124 (O_124,N_2527,N_2830);
or UO_125 (O_125,N_2641,N_4497);
nor UO_126 (O_126,N_4232,N_2522);
nor UO_127 (O_127,N_2592,N_4578);
nand UO_128 (O_128,N_4132,N_2812);
nand UO_129 (O_129,N_3452,N_4983);
nand UO_130 (O_130,N_3185,N_3140);
nand UO_131 (O_131,N_3811,N_4646);
nand UO_132 (O_132,N_3563,N_3219);
or UO_133 (O_133,N_3236,N_4798);
nand UO_134 (O_134,N_4066,N_3902);
and UO_135 (O_135,N_3851,N_2900);
nor UO_136 (O_136,N_4337,N_3519);
nand UO_137 (O_137,N_3561,N_3623);
or UO_138 (O_138,N_3651,N_3990);
or UO_139 (O_139,N_4709,N_2786);
and UO_140 (O_140,N_3387,N_4175);
or UO_141 (O_141,N_3406,N_4192);
nor UO_142 (O_142,N_3695,N_2754);
nor UO_143 (O_143,N_2842,N_3885);
and UO_144 (O_144,N_4609,N_4937);
nor UO_145 (O_145,N_3079,N_4622);
and UO_146 (O_146,N_4860,N_3763);
nand UO_147 (O_147,N_3457,N_3667);
or UO_148 (O_148,N_4303,N_3098);
or UO_149 (O_149,N_4920,N_4307);
and UO_150 (O_150,N_4114,N_3987);
or UO_151 (O_151,N_4276,N_3118);
nor UO_152 (O_152,N_4209,N_3405);
or UO_153 (O_153,N_3146,N_2977);
or UO_154 (O_154,N_2575,N_3580);
or UO_155 (O_155,N_2585,N_3108);
or UO_156 (O_156,N_2506,N_4822);
nand UO_157 (O_157,N_3817,N_4814);
nand UO_158 (O_158,N_4507,N_2716);
or UO_159 (O_159,N_3957,N_3099);
nor UO_160 (O_160,N_3947,N_4797);
nor UO_161 (O_161,N_3206,N_4903);
or UO_162 (O_162,N_3532,N_4081);
and UO_163 (O_163,N_2908,N_4629);
or UO_164 (O_164,N_3512,N_2586);
and UO_165 (O_165,N_3592,N_4413);
nand UO_166 (O_166,N_4156,N_3513);
nand UO_167 (O_167,N_3223,N_3715);
or UO_168 (O_168,N_3566,N_4710);
nor UO_169 (O_169,N_4766,N_2560);
or UO_170 (O_170,N_3562,N_3071);
nor UO_171 (O_171,N_4618,N_3474);
nor UO_172 (O_172,N_3411,N_3523);
nor UO_173 (O_173,N_4368,N_2596);
nand UO_174 (O_174,N_3261,N_4402);
nand UO_175 (O_175,N_2771,N_4202);
nor UO_176 (O_176,N_4452,N_4301);
nand UO_177 (O_177,N_4215,N_3455);
nand UO_178 (O_178,N_2869,N_3390);
nor UO_179 (O_179,N_3785,N_3699);
or UO_180 (O_180,N_4263,N_4640);
nand UO_181 (O_181,N_3921,N_4907);
nand UO_182 (O_182,N_2965,N_2783);
and UO_183 (O_183,N_4272,N_2836);
nand UO_184 (O_184,N_2728,N_2530);
and UO_185 (O_185,N_3136,N_3683);
or UO_186 (O_186,N_4558,N_3493);
nand UO_187 (O_187,N_4249,N_2573);
nand UO_188 (O_188,N_4064,N_2802);
and UO_189 (O_189,N_4626,N_3126);
and UO_190 (O_190,N_4942,N_4031);
nand UO_191 (O_191,N_3091,N_4078);
nand UO_192 (O_192,N_4333,N_4160);
nor UO_193 (O_193,N_4107,N_3470);
and UO_194 (O_194,N_4043,N_3692);
nand UO_195 (O_195,N_4668,N_2893);
or UO_196 (O_196,N_3367,N_3756);
nand UO_197 (O_197,N_4734,N_2511);
nand UO_198 (O_198,N_4138,N_4258);
nand UO_199 (O_199,N_4864,N_4556);
or UO_200 (O_200,N_2659,N_3906);
nand UO_201 (O_201,N_3680,N_4525);
nand UO_202 (O_202,N_3127,N_3149);
nor UO_203 (O_203,N_3023,N_4322);
or UO_204 (O_204,N_3294,N_2753);
nor UO_205 (O_205,N_4890,N_4389);
and UO_206 (O_206,N_3832,N_4938);
nand UO_207 (O_207,N_3321,N_4665);
nor UO_208 (O_208,N_3518,N_4690);
nand UO_209 (O_209,N_4635,N_3451);
nand UO_210 (O_210,N_3431,N_3332);
or UO_211 (O_211,N_4648,N_3840);
nand UO_212 (O_212,N_3650,N_4170);
and UO_213 (O_213,N_4973,N_4625);
or UO_214 (O_214,N_2899,N_3031);
nor UO_215 (O_215,N_4291,N_4586);
nor UO_216 (O_216,N_2599,N_4611);
nor UO_217 (O_217,N_3361,N_3191);
and UO_218 (O_218,N_3069,N_3287);
or UO_219 (O_219,N_2672,N_4387);
nand UO_220 (O_220,N_4863,N_2706);
and UO_221 (O_221,N_4824,N_2680);
or UO_222 (O_222,N_3235,N_3085);
and UO_223 (O_223,N_4419,N_4844);
nand UO_224 (O_224,N_3612,N_3285);
nor UO_225 (O_225,N_4104,N_4197);
nand UO_226 (O_226,N_4155,N_4813);
and UO_227 (O_227,N_4165,N_4529);
or UO_228 (O_228,N_3268,N_4252);
nand UO_229 (O_229,N_4163,N_3066);
nor UO_230 (O_230,N_4807,N_2745);
nand UO_231 (O_231,N_3861,N_2790);
or UO_232 (O_232,N_4906,N_4216);
and UO_233 (O_233,N_4040,N_4977);
and UO_234 (O_234,N_4998,N_4801);
nor UO_235 (O_235,N_2904,N_3059);
nor UO_236 (O_236,N_3995,N_4590);
xor UO_237 (O_237,N_3454,N_3831);
nand UO_238 (O_238,N_4003,N_4966);
nor UO_239 (O_239,N_4070,N_4188);
nand UO_240 (O_240,N_4696,N_4129);
and UO_241 (O_241,N_2514,N_3105);
and UO_242 (O_242,N_4479,N_2545);
nor UO_243 (O_243,N_2637,N_3952);
nor UO_244 (O_244,N_4345,N_4711);
and UO_245 (O_245,N_3167,N_3117);
xor UO_246 (O_246,N_4012,N_3196);
or UO_247 (O_247,N_4968,N_4051);
nand UO_248 (O_248,N_2841,N_3577);
nor UO_249 (O_249,N_3057,N_2591);
nand UO_250 (O_250,N_3111,N_4817);
nor UO_251 (O_251,N_4426,N_3251);
nor UO_252 (O_252,N_4340,N_4872);
or UO_253 (O_253,N_4171,N_4544);
and UO_254 (O_254,N_2837,N_3988);
nand UO_255 (O_255,N_4220,N_4453);
or UO_256 (O_256,N_4999,N_4045);
and UO_257 (O_257,N_4458,N_3002);
nand UO_258 (O_258,N_4808,N_2763);
nor UO_259 (O_259,N_4972,N_2963);
nand UO_260 (O_260,N_3645,N_3366);
nor UO_261 (O_261,N_3298,N_4555);
or UO_262 (O_262,N_2666,N_2871);
or UO_263 (O_263,N_3745,N_3021);
nor UO_264 (O_264,N_3033,N_2877);
nand UO_265 (O_265,N_4261,N_2799);
nand UO_266 (O_266,N_3273,N_2998);
nand UO_267 (O_267,N_4526,N_4073);
nor UO_268 (O_268,N_4634,N_4795);
nand UO_269 (O_269,N_3578,N_3310);
and UO_270 (O_270,N_3511,N_3976);
and UO_271 (O_271,N_2950,N_4508);
or UO_272 (O_272,N_4559,N_4666);
or UO_273 (O_273,N_4986,N_3173);
and UO_274 (O_274,N_4898,N_4985);
nor UO_275 (O_275,N_4207,N_3008);
or UO_276 (O_276,N_4299,N_4224);
or UO_277 (O_277,N_4425,N_3720);
or UO_278 (O_278,N_4122,N_3796);
xnor UO_279 (O_279,N_4598,N_3686);
nor UO_280 (O_280,N_2554,N_3170);
nand UO_281 (O_281,N_4738,N_4563);
and UO_282 (O_282,N_4357,N_4480);
nand UO_283 (O_283,N_4628,N_4915);
nand UO_284 (O_284,N_3249,N_2984);
and UO_285 (O_285,N_2606,N_2559);
nor UO_286 (O_286,N_3247,N_3172);
nor UO_287 (O_287,N_4284,N_3567);
nor UO_288 (O_288,N_3601,N_3489);
or UO_289 (O_289,N_2682,N_2911);
nor UO_290 (O_290,N_2513,N_3914);
nor UO_291 (O_291,N_4455,N_3216);
nor UO_292 (O_292,N_4536,N_3279);
and UO_293 (O_293,N_3682,N_4530);
and UO_294 (O_294,N_3202,N_2537);
or UO_295 (O_295,N_4941,N_2809);
nor UO_296 (O_296,N_3739,N_4523);
nand UO_297 (O_297,N_3393,N_2797);
nand UO_298 (O_298,N_3487,N_2821);
nand UO_299 (O_299,N_3940,N_4137);
nand UO_300 (O_300,N_2721,N_3838);
xor UO_301 (O_301,N_3222,N_4444);
nand UO_302 (O_302,N_3536,N_4853);
nand UO_303 (O_303,N_3859,N_2558);
nand UO_304 (O_304,N_3169,N_3590);
and UO_305 (O_305,N_4067,N_3388);
nand UO_306 (O_306,N_2712,N_4957);
and UO_307 (O_307,N_4296,N_4323);
or UO_308 (O_308,N_4353,N_2807);
nand UO_309 (O_309,N_4348,N_2915);
nor UO_310 (O_310,N_2598,N_3582);
nand UO_311 (O_311,N_2536,N_2538);
xor UO_312 (O_312,N_4873,N_3538);
nor UO_313 (O_313,N_3807,N_4580);
or UO_314 (O_314,N_3965,N_3176);
or UO_315 (O_315,N_4737,N_3701);
and UO_316 (O_316,N_2631,N_4505);
nor UO_317 (O_317,N_4700,N_3727);
nand UO_318 (O_318,N_4180,N_2818);
nor UO_319 (O_319,N_3938,N_3576);
or UO_320 (O_320,N_2781,N_3320);
or UO_321 (O_321,N_4325,N_4673);
nand UO_322 (O_322,N_3596,N_2964);
nor UO_323 (O_323,N_3032,N_2889);
and UO_324 (O_324,N_4749,N_3437);
and UO_325 (O_325,N_4270,N_4532);
or UO_326 (O_326,N_4926,N_3659);
xor UO_327 (O_327,N_3174,N_4406);
nor UO_328 (O_328,N_2879,N_3936);
and UO_329 (O_329,N_4153,N_4971);
nor UO_330 (O_330,N_2746,N_3164);
and UO_331 (O_331,N_2774,N_3631);
and UO_332 (O_332,N_4764,N_2738);
and UO_333 (O_333,N_2635,N_3992);
nand UO_334 (O_334,N_3438,N_3029);
nor UO_335 (O_335,N_4214,N_3931);
nand UO_336 (O_336,N_4395,N_4405);
nand UO_337 (O_337,N_4408,N_3089);
and UO_338 (O_338,N_2542,N_3045);
and UO_339 (O_339,N_2761,N_2697);
and UO_340 (O_340,N_4740,N_3381);
nor UO_341 (O_341,N_4211,N_4878);
or UO_342 (O_342,N_3907,N_2846);
nand UO_343 (O_343,N_4819,N_2923);
nand UO_344 (O_344,N_3205,N_3314);
nor UO_345 (O_345,N_3056,N_3755);
nor UO_346 (O_346,N_2811,N_3442);
nand UO_347 (O_347,N_3060,N_3449);
nor UO_348 (O_348,N_4837,N_3100);
nor UO_349 (O_349,N_4421,N_3820);
nand UO_350 (O_350,N_4639,N_4135);
nand UO_351 (O_351,N_4437,N_4065);
nor UO_352 (O_352,N_4615,N_2700);
and UO_353 (O_353,N_3669,N_2634);
nor UO_354 (O_354,N_4116,N_4140);
nand UO_355 (O_355,N_3737,N_2941);
nand UO_356 (O_356,N_3554,N_4351);
or UO_357 (O_357,N_4855,N_3629);
nor UO_358 (O_358,N_3055,N_4484);
or UO_359 (O_359,N_3028,N_4489);
nor UO_360 (O_360,N_4531,N_3565);
nor UO_361 (O_361,N_3277,N_3621);
and UO_362 (O_362,N_4806,N_3549);
or UO_363 (O_363,N_4546,N_3943);
and UO_364 (O_364,N_3194,N_4791);
and UO_365 (O_365,N_3553,N_3731);
and UO_366 (O_366,N_2764,N_2698);
nor UO_367 (O_367,N_3613,N_4894);
nor UO_368 (O_368,N_3684,N_3080);
nor UO_369 (O_369,N_3283,N_4693);
nand UO_370 (O_370,N_2667,N_3537);
and UO_371 (O_371,N_4191,N_3062);
nor UO_372 (O_372,N_4794,N_3327);
or UO_373 (O_373,N_3276,N_3730);
or UO_374 (O_374,N_4145,N_4183);
and UO_375 (O_375,N_3847,N_2887);
or UO_376 (O_376,N_3469,N_4354);
and UO_377 (O_377,N_2524,N_4811);
or UO_378 (O_378,N_4584,N_3719);
nand UO_379 (O_379,N_4702,N_4223);
nor UO_380 (O_380,N_4945,N_3614);
nand UO_381 (O_381,N_4483,N_3989);
and UO_382 (O_382,N_3560,N_3912);
nor UO_383 (O_383,N_3122,N_3648);
and UO_384 (O_384,N_3378,N_2902);
nor UO_385 (O_385,N_3234,N_4158);
nor UO_386 (O_386,N_3688,N_4880);
nor UO_387 (O_387,N_4747,N_3307);
nand UO_388 (O_388,N_4757,N_4705);
nand UO_389 (O_389,N_2884,N_2665);
and UO_390 (O_390,N_4804,N_3878);
and UO_391 (O_391,N_3910,N_3357);
and UO_392 (O_392,N_4786,N_2897);
nand UO_393 (O_393,N_3646,N_3890);
and UO_394 (O_394,N_3675,N_2689);
nor UO_395 (O_395,N_3043,N_3114);
and UO_396 (O_396,N_4335,N_4098);
or UO_397 (O_397,N_4835,N_2710);
nand UO_398 (O_398,N_2517,N_4472);
nand UO_399 (O_399,N_3761,N_3119);
nand UO_400 (O_400,N_2910,N_3991);
and UO_401 (O_401,N_3783,N_3759);
nand UO_402 (O_402,N_2692,N_4150);
xor UO_403 (O_403,N_2520,N_2734);
or UO_404 (O_404,N_4871,N_4476);
and UO_405 (O_405,N_4346,N_2744);
or UO_406 (O_406,N_3770,N_3131);
nor UO_407 (O_407,N_4416,N_3805);
or UO_408 (O_408,N_3128,N_3213);
nand UO_409 (O_409,N_4305,N_3721);
nor UO_410 (O_410,N_4130,N_4256);
or UO_411 (O_411,N_4278,N_4290);
and UO_412 (O_412,N_3142,N_3556);
or UO_413 (O_413,N_3150,N_3974);
and UO_414 (O_414,N_2556,N_4091);
xor UO_415 (O_415,N_3003,N_3225);
nor UO_416 (O_416,N_4362,N_3679);
nand UO_417 (O_417,N_2916,N_3981);
or UO_418 (O_418,N_3415,N_4044);
nor UO_419 (O_419,N_3464,N_2742);
nor UO_420 (O_420,N_2539,N_2593);
nand UO_421 (O_421,N_2623,N_3020);
or UO_422 (O_422,N_3384,N_4516);
nand UO_423 (O_423,N_3937,N_3171);
nor UO_424 (O_424,N_3640,N_3997);
nand UO_425 (O_425,N_2519,N_3499);
nand UO_426 (O_426,N_3058,N_4317);
nand UO_427 (O_427,N_2588,N_4688);
nand UO_428 (O_428,N_2733,N_4493);
or UO_429 (O_429,N_3143,N_2864);
and UO_430 (O_430,N_3839,N_3445);
nand UO_431 (O_431,N_2737,N_4877);
nand UO_432 (O_432,N_4830,N_4931);
or UO_433 (O_433,N_4025,N_3665);
or UO_434 (O_434,N_3559,N_4796);
or UO_435 (O_435,N_4084,N_3120);
or UO_436 (O_436,N_2800,N_2845);
nor UO_437 (O_437,N_3795,N_4131);
nand UO_438 (O_438,N_3822,N_4203);
nand UO_439 (O_439,N_4285,N_4498);
and UO_440 (O_440,N_3490,N_4522);
nor UO_441 (O_441,N_2740,N_4016);
nand UO_442 (O_442,N_4103,N_4339);
or UO_443 (O_443,N_4265,N_4962);
and UO_444 (O_444,N_3157,N_4446);
and UO_445 (O_445,N_3281,N_3776);
nand UO_446 (O_446,N_4432,N_2801);
or UO_447 (O_447,N_3960,N_4773);
or UO_448 (O_448,N_3282,N_2578);
and UO_449 (O_449,N_2974,N_4225);
nor UO_450 (O_450,N_3121,N_2855);
or UO_451 (O_451,N_3753,N_3063);
and UO_452 (O_452,N_4002,N_3401);
nor UO_453 (O_453,N_4143,N_3246);
nor UO_454 (O_454,N_4958,N_2670);
nand UO_455 (O_455,N_2550,N_4101);
nand UO_456 (O_456,N_3954,N_3942);
nor UO_457 (O_457,N_4481,N_2794);
nor UO_458 (O_458,N_4519,N_4179);
nand UO_459 (O_459,N_3124,N_3221);
nor UO_460 (O_460,N_2883,N_2945);
and UO_461 (O_461,N_3813,N_4541);
and UO_462 (O_462,N_4714,N_2833);
nand UO_463 (O_463,N_3165,N_4311);
or UO_464 (O_464,N_4185,N_2688);
nand UO_465 (O_465,N_2867,N_2814);
nand UO_466 (O_466,N_3703,N_2508);
and UO_467 (O_467,N_3472,N_2961);
and UO_468 (O_468,N_3369,N_3244);
and UO_469 (O_469,N_2565,N_3193);
or UO_470 (O_470,N_3004,N_3227);
nor UO_471 (O_471,N_4733,N_3242);
nor UO_472 (O_472,N_2626,N_4241);
nand UO_473 (O_473,N_2678,N_4009);
nor UO_474 (O_474,N_3382,N_2662);
nand UO_475 (O_475,N_2892,N_2832);
or UO_476 (O_476,N_4398,N_4910);
or UO_477 (O_477,N_2958,N_4631);
and UO_478 (O_478,N_2638,N_4074);
nand UO_479 (O_479,N_3799,N_3712);
nor UO_480 (O_480,N_3866,N_4816);
nor UO_481 (O_481,N_4071,N_3856);
and UO_482 (O_482,N_3535,N_4857);
nand UO_483 (O_483,N_2999,N_3919);
nand UO_484 (O_484,N_4698,N_4028);
and UO_485 (O_485,N_3414,N_4491);
or UO_486 (O_486,N_4637,N_4858);
or UO_487 (O_487,N_4072,N_4647);
nand UO_488 (O_488,N_3312,N_3342);
nor UO_489 (O_489,N_4049,N_2762);
nand UO_490 (O_490,N_2562,N_3198);
nand UO_491 (O_491,N_4701,N_2553);
or UO_492 (O_492,N_4088,N_3935);
or UO_493 (O_493,N_3463,N_3531);
and UO_494 (O_494,N_2948,N_4984);
or UO_495 (O_495,N_3133,N_4314);
nand UO_496 (O_496,N_2654,N_3286);
and UO_497 (O_497,N_3955,N_4704);
or UO_498 (O_498,N_2555,N_3752);
and UO_499 (O_499,N_4238,N_4246);
and UO_500 (O_500,N_4090,N_2549);
and UO_501 (O_501,N_3266,N_4273);
nand UO_502 (O_502,N_2660,N_4077);
or UO_503 (O_503,N_3527,N_2857);
nor UO_504 (O_504,N_4513,N_4744);
nand UO_505 (O_505,N_3263,N_2834);
or UO_506 (O_506,N_4597,N_3096);
or UO_507 (O_507,N_4230,N_2656);
nor UO_508 (O_508,N_3850,N_4083);
nor UO_509 (O_509,N_4026,N_4868);
nand UO_510 (O_510,N_2827,N_4633);
and UO_511 (O_511,N_3529,N_3864);
nor UO_512 (O_512,N_4562,N_3417);
nor UO_513 (O_513,N_2690,N_4274);
nand UO_514 (O_514,N_3356,N_3272);
nand UO_515 (O_515,N_4247,N_4475);
nor UO_516 (O_516,N_4788,N_2760);
nor UO_517 (O_517,N_3226,N_4151);
and UO_518 (O_518,N_3395,N_4259);
nor UO_519 (O_519,N_2695,N_3698);
or UO_520 (O_520,N_4699,N_2655);
and UO_521 (O_521,N_4126,N_2701);
nand UO_522 (O_522,N_3801,N_4087);
nor UO_523 (O_523,N_4852,N_4375);
and UO_524 (O_524,N_3241,N_3725);
nand UO_525 (O_525,N_4599,N_4940);
or UO_526 (O_526,N_2714,N_3504);
and UO_527 (O_527,N_2810,N_4075);
or UO_528 (O_528,N_3778,N_4917);
nor UO_529 (O_529,N_4347,N_4503);
nor UO_530 (O_530,N_4385,N_4320);
nand UO_531 (O_531,N_4330,N_3998);
and UO_532 (O_532,N_3605,N_4948);
or UO_533 (O_533,N_3478,N_4499);
nand UO_534 (O_534,N_4770,N_4839);
or UO_535 (O_535,N_4279,N_4349);
nor UO_536 (O_536,N_4888,N_2587);
or UO_537 (O_537,N_4502,N_2613);
nor UO_538 (O_538,N_3481,N_3754);
nand UO_539 (O_539,N_3867,N_3828);
nand UO_540 (O_540,N_3588,N_3652);
or UO_541 (O_541,N_4079,N_2936);
nor UO_542 (O_542,N_4228,N_2859);
nand UO_543 (O_543,N_2563,N_3476);
and UO_544 (O_544,N_4685,N_4537);
or UO_545 (O_545,N_2939,N_4856);
and UO_546 (O_546,N_4254,N_3780);
and UO_547 (O_547,N_2906,N_4845);
nor UO_548 (O_548,N_3690,N_4474);
nor UO_549 (O_549,N_3600,N_2574);
and UO_550 (O_550,N_4774,N_4233);
or UO_551 (O_551,N_4050,N_3873);
and UO_552 (O_552,N_2970,N_3154);
and UO_553 (O_553,N_4978,N_4547);
nand UO_554 (O_554,N_2888,N_3137);
nand UO_555 (O_555,N_3837,N_4778);
or UO_556 (O_556,N_3083,N_4099);
nand UO_557 (O_557,N_2645,N_2572);
nor UO_558 (O_558,N_3422,N_3550);
nand UO_559 (O_559,N_2815,N_4588);
or UO_560 (O_560,N_3232,N_4161);
nor UO_561 (O_561,N_4534,N_3594);
or UO_562 (O_562,N_2567,N_3238);
and UO_563 (O_563,N_4694,N_3428);
nor UO_564 (O_564,N_4282,N_2788);
nor UO_565 (O_565,N_3017,N_3728);
or UO_566 (O_566,N_2813,N_4849);
and UO_567 (O_567,N_4149,N_4443);
and UO_568 (O_568,N_3371,N_3636);
nor UO_569 (O_569,N_4391,N_4922);
or UO_570 (O_570,N_3257,N_4538);
and UO_571 (O_571,N_4939,N_2926);
nand UO_572 (O_572,N_4846,N_4415);
and UO_573 (O_573,N_3534,N_4380);
or UO_574 (O_574,N_2624,N_3655);
nand UO_575 (O_575,N_4501,N_3358);
nor UO_576 (O_576,N_3953,N_4409);
and UO_577 (O_577,N_3868,N_4956);
nand UO_578 (O_578,N_4927,N_2789);
nor UO_579 (O_579,N_4198,N_2776);
nor UO_580 (O_580,N_4048,N_4524);
nand UO_581 (O_581,N_3635,N_4036);
and UO_582 (O_582,N_4407,N_3163);
and UO_583 (O_583,N_3815,N_3380);
or UO_584 (O_584,N_4396,N_3933);
or UO_585 (O_585,N_4141,N_2956);
or UO_586 (O_586,N_3231,N_2972);
nor UO_587 (O_587,N_3610,N_4271);
nand UO_588 (O_588,N_3427,N_3315);
and UO_589 (O_589,N_4728,N_3188);
or UO_590 (O_590,N_3259,N_4068);
and UO_591 (O_591,N_4394,N_2868);
nand UO_592 (O_592,N_2600,N_4430);
or UO_593 (O_593,N_2685,N_3894);
or UO_594 (O_594,N_4392,N_2983);
and UO_595 (O_595,N_3830,N_2653);
nand UO_596 (O_596,N_4251,N_3525);
nor UO_597 (O_597,N_2651,N_3052);
nand UO_598 (O_598,N_3994,N_4361);
nor UO_599 (O_599,N_4373,N_3674);
nand UO_600 (O_600,N_3608,N_3641);
or UO_601 (O_601,N_2995,N_2529);
nor UO_602 (O_602,N_2957,N_2920);
or UO_603 (O_603,N_3199,N_3985);
and UO_604 (O_604,N_3762,N_3435);
nor UO_605 (O_605,N_3040,N_2766);
nand UO_606 (O_606,N_2921,N_3139);
nand UO_607 (O_607,N_3901,N_2848);
nor UO_608 (O_608,N_3322,N_2561);
and UO_609 (O_609,N_2707,N_4176);
nor UO_610 (O_610,N_3258,N_2579);
nand UO_611 (O_611,N_3983,N_4466);
and UO_612 (O_612,N_2551,N_3506);
nor UO_613 (O_613,N_3552,N_4359);
nand UO_614 (O_614,N_3706,N_3649);
nor UO_615 (O_615,N_4239,N_3168);
or UO_616 (O_616,N_4435,N_3691);
nand UO_617 (O_617,N_4055,N_2978);
nand UO_618 (O_618,N_2501,N_3333);
nand UO_619 (O_619,N_3240,N_3833);
or UO_620 (O_620,N_4784,N_4100);
nor UO_621 (O_621,N_3011,N_4936);
and UO_622 (O_622,N_2727,N_3824);
and UO_623 (O_623,N_4275,N_3076);
or UO_624 (O_624,N_4605,N_3178);
or UO_625 (O_625,N_4029,N_4226);
and UO_626 (O_626,N_3597,N_3486);
and UO_627 (O_627,N_3044,N_3758);
nand UO_628 (O_628,N_3197,N_4540);
nand UO_629 (O_629,N_3779,N_4754);
and UO_630 (O_630,N_3364,N_3152);
nor UO_631 (O_631,N_4836,N_2711);
or UO_632 (O_632,N_3845,N_3498);
nor UO_633 (O_633,N_3911,N_4449);
xor UO_634 (O_634,N_3934,N_4181);
and UO_635 (O_635,N_4309,N_2953);
nor UO_636 (O_636,N_2748,N_3295);
nand UO_637 (O_637,N_3654,N_3477);
nand UO_638 (O_638,N_4434,N_4731);
nand UO_639 (O_639,N_2933,N_2994);
nor UO_640 (O_640,N_3354,N_3742);
or UO_641 (O_641,N_2891,N_4790);
or UO_642 (O_642,N_4617,N_2912);
or UO_643 (O_643,N_3966,N_2975);
nor UO_644 (O_644,N_2860,N_3360);
nand UO_645 (O_645,N_2838,N_2726);
or UO_646 (O_646,N_3980,N_3372);
and UO_647 (O_647,N_4004,N_4159);
nor UO_648 (O_648,N_2566,N_3302);
nand UO_649 (O_649,N_2808,N_4060);
or UO_650 (O_650,N_3237,N_3630);
nand UO_651 (O_651,N_4379,N_2935);
nand UO_652 (O_652,N_3228,N_3325);
nand UO_653 (O_653,N_2500,N_4900);
nand UO_654 (O_654,N_3424,N_3109);
and UO_655 (O_655,N_3696,N_4454);
nor UO_656 (O_656,N_3639,N_3115);
or UO_657 (O_657,N_4924,N_2854);
or UO_658 (O_658,N_4334,N_3892);
nor UO_659 (O_659,N_2552,N_4655);
nand UO_660 (O_660,N_3810,N_3624);
nand UO_661 (O_661,N_2741,N_2540);
and UO_662 (O_662,N_3962,N_2785);
nor UO_663 (O_663,N_4866,N_4264);
nand UO_664 (O_664,N_4952,N_4763);
nor UO_665 (O_665,N_2987,N_4602);
nand UO_666 (O_666,N_3808,N_3704);
nor UO_667 (O_667,N_3255,N_4492);
nand UO_668 (O_668,N_4459,N_3189);
nand UO_669 (O_669,N_3094,N_4436);
nor UO_670 (O_670,N_3179,N_4326);
nor UO_671 (O_671,N_4417,N_4495);
nand UO_672 (O_672,N_3024,N_4777);
nand UO_673 (O_673,N_3620,N_4841);
and UO_674 (O_674,N_2851,N_3723);
nand UO_675 (O_675,N_2960,N_3037);
nand UO_676 (O_676,N_2609,N_3192);
nor UO_677 (O_677,N_3009,N_2823);
xnor UO_678 (O_678,N_4382,N_4967);
or UO_679 (O_679,N_4295,N_3500);
nand UO_680 (O_680,N_3503,N_3897);
nor UO_681 (O_681,N_2880,N_3433);
xnor UO_682 (O_682,N_4234,N_2803);
nand UO_683 (O_683,N_4020,N_2875);
or UO_684 (O_684,N_2535,N_4062);
nor UO_685 (O_685,N_4916,N_4730);
or UO_686 (O_686,N_2597,N_3386);
nor UO_687 (O_687,N_3760,N_4933);
nor UO_688 (O_688,N_4697,N_4612);
and UO_689 (O_689,N_3093,N_4177);
or UO_690 (O_690,N_4390,N_2595);
nor UO_691 (O_691,N_4035,N_4017);
or UO_692 (O_692,N_4950,N_3284);
and UO_693 (O_693,N_4042,N_3702);
nand UO_694 (O_694,N_3862,N_3262);
nand UO_695 (O_695,N_4266,N_3175);
nor UO_696 (O_696,N_3082,N_3155);
or UO_697 (O_697,N_3465,N_3769);
or UO_698 (O_698,N_4769,N_2601);
nor UO_699 (O_699,N_3711,N_4616);
nand UO_700 (O_700,N_3161,N_3673);
or UO_701 (O_701,N_4799,N_4344);
nor UO_702 (O_702,N_4450,N_3328);
nor UO_703 (O_703,N_4338,N_2792);
and UO_704 (O_704,N_4011,N_4010);
nor UO_705 (O_705,N_4818,N_4995);
and UO_706 (O_706,N_3949,N_4343);
nor UO_707 (O_707,N_3663,N_3744);
or UO_708 (O_708,N_4527,N_4494);
nand UO_709 (O_709,N_3038,N_4196);
or UO_710 (O_710,N_2940,N_2604);
and UO_711 (O_711,N_3541,N_4069);
and UO_712 (O_712,N_4606,N_2664);
or UO_713 (O_713,N_3829,N_3925);
nor UO_714 (O_714,N_3458,N_2768);
or UO_715 (O_715,N_4742,N_3473);
nand UO_716 (O_716,N_4756,N_4205);
nand UO_717 (O_717,N_4515,N_3786);
and UO_718 (O_718,N_2705,N_4381);
and UO_719 (O_719,N_3685,N_4248);
nand UO_720 (O_720,N_4585,N_3095);
and UO_721 (O_721,N_2683,N_3996);
nand UO_722 (O_722,N_4401,N_2927);
or UO_723 (O_723,N_4925,N_4128);
nand UO_724 (O_724,N_3587,N_4782);
and UO_725 (O_725,N_4092,N_2739);
or UO_726 (O_726,N_3413,N_4713);
nand UO_727 (O_727,N_2582,N_3557);
nor UO_728 (O_728,N_4759,N_2796);
or UO_729 (O_729,N_4720,N_2826);
or UO_730 (O_730,N_4281,N_4378);
and UO_731 (O_731,N_3615,N_3622);
and UO_732 (O_732,N_4884,N_3306);
nor UO_733 (O_733,N_4260,N_3750);
and UO_734 (O_734,N_4034,N_4620);
or UO_735 (O_735,N_4332,N_3666);
nand UO_736 (O_736,N_3903,N_3889);
nor UO_737 (O_737,N_3888,N_2715);
nand UO_738 (O_738,N_3922,N_4775);
nor UO_739 (O_739,N_2820,N_3245);
nand UO_740 (O_740,N_2967,N_4262);
nand UO_741 (O_741,N_4550,N_3292);
nand UO_742 (O_742,N_4981,N_3589);
nor UO_743 (O_743,N_3125,N_3872);
nor UO_744 (O_744,N_3334,N_4243);
or UO_745 (O_745,N_4134,N_3151);
nor UO_746 (O_746,N_4964,N_4388);
nand UO_747 (O_747,N_4568,N_4118);
nand UO_748 (O_748,N_4195,N_4287);
or UO_749 (O_749,N_4052,N_2946);
nand UO_750 (O_750,N_3809,N_4240);
nor UO_751 (O_751,N_4461,N_4420);
nor UO_752 (O_752,N_4776,N_4997);
nand UO_753 (O_753,N_3505,N_4736);
nor UO_754 (O_754,N_3869,N_4154);
and UO_755 (O_755,N_4674,N_4566);
nand UO_756 (O_756,N_4692,N_4245);
nand UO_757 (O_757,N_3558,N_3398);
and UO_758 (O_758,N_2713,N_2856);
and UO_759 (O_759,N_2985,N_4661);
nor UO_760 (O_760,N_3564,N_2885);
or UO_761 (O_761,N_4046,N_3626);
or UO_762 (O_762,N_4928,N_4911);
nand UO_763 (O_763,N_4253,N_3288);
nand UO_764 (O_764,N_2509,N_3460);
nor UO_765 (O_765,N_4032,N_3676);
or UO_766 (O_766,N_2862,N_4231);
or UO_767 (O_767,N_3792,N_4076);
nand UO_768 (O_768,N_4596,N_3468);
nor UO_769 (O_769,N_2917,N_3441);
and UO_770 (O_770,N_4557,N_3274);
nand UO_771 (O_771,N_4120,N_3377);
or UO_772 (O_772,N_3088,N_4306);
nor UO_773 (O_773,N_4360,N_3331);
nor UO_774 (O_774,N_3440,N_4283);
or UO_775 (O_775,N_3214,N_4242);
nand UO_776 (O_776,N_4063,N_3772);
nor UO_777 (O_777,N_4869,N_4096);
or UO_778 (O_778,N_3000,N_4053);
nor UO_779 (O_779,N_2639,N_3843);
nor UO_780 (O_780,N_3068,N_3479);
and UO_781 (O_781,N_2925,N_4644);
xnor UO_782 (O_782,N_3280,N_3533);
nor UO_783 (O_783,N_3064,N_3329);
or UO_784 (O_784,N_2735,N_2993);
nor UO_785 (O_785,N_3656,N_3586);
or UO_786 (O_786,N_3526,N_2863);
and UO_787 (O_787,N_4237,N_3416);
or UO_788 (O_788,N_3293,N_3400);
or UO_789 (O_789,N_3443,N_3432);
nor UO_790 (O_790,N_4930,N_3607);
nor UO_791 (O_791,N_3112,N_4212);
nor UO_792 (O_792,N_3705,N_3501);
and UO_793 (O_793,N_4982,N_4834);
nand UO_794 (O_794,N_4935,N_2505);
nand UO_795 (O_795,N_3271,N_3956);
and UO_796 (O_796,N_4148,N_2775);
or UO_797 (O_797,N_4451,N_3797);
and UO_798 (O_798,N_2504,N_2648);
nor UO_799 (O_799,N_4681,N_2630);
nand UO_800 (O_800,N_4567,N_3791);
xor UO_801 (O_801,N_2636,N_4946);
or UO_802 (O_802,N_2991,N_2533);
xor UO_803 (O_803,N_4164,N_3858);
or UO_804 (O_804,N_3439,N_3383);
or UO_805 (O_805,N_2612,N_4178);
and UO_806 (O_806,N_4005,N_2778);
nand UO_807 (O_807,N_4462,N_2898);
or UO_808 (O_808,N_3187,N_3821);
and UO_809 (O_809,N_4094,N_3718);
and UO_810 (O_810,N_4227,N_3599);
nor UO_811 (O_811,N_3545,N_4886);
and UO_812 (O_812,N_4642,N_3113);
or UO_813 (O_813,N_4204,N_4762);
nor UO_814 (O_814,N_4893,N_4182);
nor UO_815 (O_815,N_2699,N_3102);
and UO_816 (O_816,N_4919,N_4991);
nand UO_817 (O_817,N_4117,N_4124);
nor UO_818 (O_818,N_2633,N_3546);
or UO_819 (O_819,N_2521,N_4429);
or UO_820 (O_820,N_3583,N_3835);
nand UO_821 (O_821,N_3410,N_3800);
nor UO_822 (O_822,N_4194,N_3252);
or UO_823 (O_823,N_4173,N_4980);
nand UO_824 (O_824,N_3450,N_3190);
nand UO_825 (O_825,N_3853,N_3041);
and UO_826 (O_826,N_2843,N_2730);
or UO_827 (O_827,N_4500,N_3317);
nor UO_828 (O_828,N_3816,N_4686);
and UO_829 (O_829,N_4431,N_2686);
nand UO_830 (O_830,N_3430,N_2729);
nor UO_831 (O_831,N_3670,N_4718);
nor UO_832 (O_832,N_2755,N_4944);
nor UO_833 (O_833,N_4393,N_3421);
nor UO_834 (O_834,N_3047,N_2532);
and UO_835 (O_835,N_4624,N_4623);
nor UO_836 (O_836,N_4302,N_4403);
and UO_837 (O_837,N_4372,N_3048);
nor UO_838 (O_838,N_3982,N_4427);
nor UO_839 (O_839,N_3183,N_3547);
nor UO_840 (O_840,N_4545,N_3977);
nor UO_841 (O_841,N_4848,N_2673);
nor UO_842 (O_842,N_3036,N_4636);
nand UO_843 (O_843,N_4383,N_4842);
nand UO_844 (O_844,N_4438,N_2853);
nor UO_845 (O_845,N_3324,N_2614);
nand UO_846 (O_846,N_3299,N_4572);
and UO_847 (O_847,N_4298,N_3201);
and UO_848 (O_848,N_3514,N_3330);
or UO_849 (O_849,N_3507,N_2615);
nand UO_850 (O_850,N_3301,N_2990);
or UO_851 (O_851,N_2719,N_4280);
or UO_852 (O_852,N_3700,N_4660);
and UO_853 (O_853,N_4367,N_4521);
xnor UO_854 (O_854,N_3757,N_3999);
or UO_855 (O_855,N_2969,N_3362);
and UO_856 (O_856,N_3658,N_3834);
and UO_857 (O_857,N_4024,N_2594);
or UO_858 (O_858,N_3110,N_4115);
or UO_859 (O_859,N_3418,N_3899);
nor UO_860 (O_860,N_4000,N_3773);
nor UO_861 (O_861,N_3077,N_3876);
nand UO_862 (O_862,N_4960,N_4414);
or UO_863 (O_863,N_4478,N_4815);
nand UO_864 (O_864,N_4167,N_4111);
and UO_865 (O_865,N_4574,N_3072);
nand UO_866 (O_866,N_4577,N_4831);
or UO_867 (O_867,N_4327,N_4533);
nor UO_868 (O_868,N_2822,N_3735);
nor UO_869 (O_869,N_3595,N_4712);
nand UO_870 (O_870,N_4682,N_2751);
and UO_871 (O_871,N_4504,N_4632);
nand UO_872 (O_872,N_3269,N_4030);
nand UO_873 (O_873,N_3521,N_4721);
or UO_874 (O_874,N_4918,N_4297);
and UO_875 (O_875,N_3738,N_4654);
nor UO_876 (O_876,N_4675,N_2931);
xor UO_877 (O_877,N_4059,N_4162);
nand UO_878 (O_878,N_4022,N_4468);
and UO_879 (O_879,N_4768,N_4913);
and UO_880 (O_880,N_4889,N_3857);
and UO_881 (O_881,N_3016,N_2627);
nand UO_882 (O_882,N_4560,N_4412);
nor UO_883 (O_883,N_3627,N_4146);
nand UO_884 (O_884,N_3932,N_3103);
nor UO_885 (O_885,N_3177,N_3494);
nor UO_886 (O_886,N_3767,N_4037);
nor UO_887 (O_887,N_4653,N_4199);
or UO_888 (O_888,N_4970,N_3260);
and UO_889 (O_889,N_3905,N_3186);
or UO_890 (O_890,N_3827,N_3335);
nand UO_891 (O_891,N_4312,N_4974);
nor UO_892 (O_892,N_4851,N_2878);
or UO_893 (O_893,N_4464,N_4582);
nor UO_894 (O_894,N_4953,N_3969);
or UO_895 (O_895,N_2722,N_2693);
or UO_896 (O_896,N_4901,N_4595);
or UO_897 (O_897,N_2872,N_4512);
or UO_898 (O_898,N_3475,N_3180);
or UO_899 (O_899,N_4677,N_4876);
and UO_900 (O_900,N_3968,N_4561);
or UO_901 (O_901,N_4097,N_3181);
nor UO_902 (O_902,N_4789,N_4467);
or UO_903 (O_903,N_3524,N_4318);
and UO_904 (O_904,N_4509,N_3379);
or UO_905 (O_905,N_2531,N_2992);
and UO_906 (O_906,N_2584,N_3316);
or UO_907 (O_907,N_3341,N_3806);
or UO_908 (O_908,N_2602,N_4717);
nor UO_909 (O_909,N_4899,N_3661);
nand UO_910 (O_910,N_3870,N_4085);
and UO_911 (O_911,N_4914,N_4439);
nor UO_912 (O_912,N_2605,N_3539);
nor UO_913 (O_913,N_4356,N_4679);
nor UO_914 (O_914,N_4656,N_4961);
and UO_915 (O_915,N_3971,N_3337);
nand UO_916 (O_916,N_4168,N_4033);
and UO_917 (O_917,N_4418,N_4650);
or UO_918 (O_918,N_3485,N_2825);
and UO_919 (O_919,N_3311,N_2687);
or UO_920 (O_920,N_3446,N_3209);
nor UO_921 (O_921,N_3860,N_4904);
nand UO_922 (O_922,N_4645,N_4331);
nor UO_923 (O_923,N_2971,N_3215);
and UO_924 (O_924,N_3278,N_2866);
and UO_925 (O_925,N_2590,N_4592);
nand UO_926 (O_926,N_3740,N_3347);
and UO_927 (O_927,N_4217,N_2640);
nand UO_928 (O_928,N_4485,N_2955);
nor UO_929 (O_929,N_3736,N_2805);
nand UO_930 (O_930,N_2643,N_4292);
and UO_931 (O_931,N_3027,N_3898);
and UO_932 (O_932,N_2876,N_4771);
or UO_933 (O_933,N_3355,N_3239);
nand UO_934 (O_934,N_4838,N_4895);
nor UO_935 (O_935,N_4949,N_3887);
nand UO_936 (O_936,N_2581,N_2752);
nor UO_937 (O_937,N_4310,N_3138);
nand UO_938 (O_938,N_2913,N_2724);
nand UO_939 (O_939,N_3018,N_3370);
nor UO_940 (O_940,N_4047,N_3606);
nor UO_941 (O_941,N_3909,N_4934);
nand UO_942 (O_942,N_2756,N_3014);
nand UO_943 (O_943,N_3087,N_3634);
or UO_944 (O_944,N_4826,N_4056);
nand UO_945 (O_945,N_4847,N_3067);
or UO_946 (O_946,N_3734,N_2968);
nor UO_947 (O_947,N_4765,N_4707);
or UO_948 (O_948,N_4772,N_4703);
nor UO_949 (O_949,N_4638,N_2784);
or UO_950 (O_950,N_3375,N_3729);
nor UO_951 (O_951,N_3884,N_4610);
and UO_952 (O_952,N_3010,N_2541);
or UO_953 (O_953,N_4678,N_3958);
nand UO_954 (O_954,N_4397,N_2621);
or UO_955 (O_955,N_3182,N_2896);
nor UO_956 (O_956,N_3160,N_4222);
and UO_957 (O_957,N_3233,N_4133);
nand UO_958 (O_958,N_3993,N_4670);
or UO_959 (O_959,N_3842,N_2515);
and UO_960 (O_960,N_4746,N_3748);
or UO_961 (O_961,N_4127,N_3653);
nor UO_962 (O_962,N_4014,N_4627);
and UO_963 (O_963,N_3603,N_3678);
and UO_964 (O_964,N_4433,N_3116);
and UO_965 (O_965,N_3253,N_3212);
or UO_966 (O_966,N_2743,N_4897);
or UO_967 (O_967,N_2929,N_2795);
or UO_968 (O_968,N_3863,N_3855);
nor UO_969 (O_969,N_4007,N_3709);
nor UO_970 (O_970,N_2949,N_4821);
nand UO_971 (O_971,N_3030,N_4328);
and UO_972 (O_972,N_2723,N_4810);
nor UO_973 (O_973,N_4106,N_4643);
nor UO_974 (O_974,N_3598,N_2988);
and UO_975 (O_975,N_4400,N_3448);
nor UO_976 (O_976,N_3159,N_3166);
or UO_977 (O_977,N_4581,N_3781);
and UO_978 (O_978,N_3275,N_3689);
and UO_979 (O_979,N_3848,N_3865);
nor UO_980 (O_980,N_2681,N_3789);
or UO_981 (O_981,N_4365,N_4865);
xor UO_982 (O_982,N_3203,N_3542);
or UO_983 (O_983,N_3790,N_4570);
nor UO_984 (O_984,N_4374,N_2759);
nand UO_985 (O_985,N_3313,N_3746);
nand UO_986 (O_986,N_4553,N_2608);
nand UO_987 (O_987,N_4750,N_4350);
or UO_988 (O_988,N_3918,N_3340);
and UO_989 (O_989,N_3618,N_3374);
nor UO_990 (O_990,N_2720,N_2780);
nand UO_991 (O_991,N_3509,N_4708);
nand UO_992 (O_992,N_4460,N_4208);
nor UO_993 (O_993,N_3814,N_3522);
and UO_994 (O_994,N_4267,N_2570);
nand UO_995 (O_995,N_4206,N_3078);
nor UO_996 (O_996,N_4528,N_2828);
nor UO_997 (O_997,N_2951,N_2564);
and UO_998 (O_998,N_3625,N_4739);
nor UO_999 (O_999,N_3891,N_4812);
endmodule