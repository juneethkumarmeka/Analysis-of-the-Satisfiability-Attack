module basic_1500_15000_2000_50_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_768,In_1067);
and U1 (N_1,In_1255,In_684);
xor U2 (N_2,In_1234,In_1425);
and U3 (N_3,In_245,In_129);
xnor U4 (N_4,In_695,In_1185);
nor U5 (N_5,In_1250,In_102);
and U6 (N_6,In_1410,In_602);
and U7 (N_7,In_1267,In_276);
xor U8 (N_8,In_1082,In_985);
and U9 (N_9,In_422,In_429);
or U10 (N_10,In_1162,In_1358);
and U11 (N_11,In_740,In_809);
or U12 (N_12,In_1188,In_577);
or U13 (N_13,In_352,In_901);
nand U14 (N_14,In_1291,In_241);
nand U15 (N_15,In_887,In_1137);
xnor U16 (N_16,In_708,In_337);
or U17 (N_17,In_304,In_555);
nand U18 (N_18,In_675,In_1089);
nand U19 (N_19,In_1120,In_842);
nand U20 (N_20,In_1406,In_867);
or U21 (N_21,In_1353,In_355);
xnor U22 (N_22,In_882,In_915);
nand U23 (N_23,In_1369,In_759);
or U24 (N_24,In_939,In_1157);
nand U25 (N_25,In_356,In_1233);
nor U26 (N_26,In_2,In_153);
or U27 (N_27,In_1390,In_1294);
xor U28 (N_28,In_1438,In_820);
nand U29 (N_29,In_1262,In_667);
nand U30 (N_30,In_539,In_335);
nor U31 (N_31,In_664,In_475);
nor U32 (N_32,In_916,In_285);
nand U33 (N_33,In_24,In_1346);
or U34 (N_34,In_793,In_636);
xor U35 (N_35,In_1257,In_609);
and U36 (N_36,In_169,In_767);
nand U37 (N_37,In_907,In_1416);
nand U38 (N_38,In_604,In_1434);
xnor U39 (N_39,In_1393,In_653);
nand U40 (N_40,In_479,In_472);
or U41 (N_41,In_1072,In_1027);
or U42 (N_42,In_1460,In_775);
and U43 (N_43,In_681,In_607);
nand U44 (N_44,In_891,In_384);
xnor U45 (N_45,In_453,In_417);
nor U46 (N_46,In_535,In_207);
or U47 (N_47,In_909,In_175);
and U48 (N_48,In_154,In_1236);
and U49 (N_49,In_856,In_430);
nor U50 (N_50,In_1321,In_381);
xor U51 (N_51,In_630,In_934);
and U52 (N_52,In_1190,In_506);
nand U53 (N_53,In_427,In_493);
and U54 (N_54,In_1465,In_1286);
nor U55 (N_55,In_1242,In_1090);
or U56 (N_56,In_197,In_263);
or U57 (N_57,In_124,In_1145);
nand U58 (N_58,In_251,In_502);
or U59 (N_59,In_77,In_394);
and U60 (N_60,In_596,In_1117);
or U61 (N_61,In_103,In_1037);
and U62 (N_62,In_1453,In_974);
nor U63 (N_63,In_1379,In_1340);
nor U64 (N_64,In_1451,In_970);
nand U65 (N_65,In_1287,In_371);
xor U66 (N_66,In_801,In_1450);
xnor U67 (N_67,In_266,In_733);
xor U68 (N_68,In_1354,In_1490);
nand U69 (N_69,In_404,In_271);
or U70 (N_70,In_1179,In_520);
or U71 (N_71,In_1079,In_550);
xor U72 (N_72,In_813,In_803);
nand U73 (N_73,In_126,In_998);
nand U74 (N_74,In_327,In_328);
or U75 (N_75,In_996,In_713);
nor U76 (N_76,In_306,In_652);
nand U77 (N_77,In_869,In_81);
or U78 (N_78,In_42,In_886);
or U79 (N_79,In_43,In_61);
nand U80 (N_80,In_936,In_1182);
nor U81 (N_81,In_331,In_325);
nand U82 (N_82,In_38,In_569);
xor U83 (N_83,In_938,In_552);
nand U84 (N_84,In_829,In_487);
and U85 (N_85,In_1183,In_1070);
or U86 (N_86,In_255,In_572);
xnor U87 (N_87,In_534,In_150);
nand U88 (N_88,In_185,In_1311);
xnor U89 (N_89,In_471,In_1337);
xor U90 (N_90,In_946,In_835);
or U91 (N_91,In_1269,In_1094);
xnor U92 (N_92,In_12,In_774);
and U93 (N_93,In_74,In_1423);
nor U94 (N_94,In_1122,In_359);
or U95 (N_95,In_498,In_1331);
and U96 (N_96,In_1196,In_1116);
and U97 (N_97,In_615,In_1228);
and U98 (N_98,In_1436,In_106);
xnor U99 (N_99,In_1235,In_629);
and U100 (N_100,In_318,In_1356);
nand U101 (N_101,In_1433,In_966);
nand U102 (N_102,In_1386,In_388);
and U103 (N_103,In_620,In_123);
nor U104 (N_104,In_613,In_884);
xnor U105 (N_105,In_156,In_1109);
nand U106 (N_106,In_1350,In_990);
or U107 (N_107,In_346,In_1456);
or U108 (N_108,In_899,In_1132);
and U109 (N_109,In_568,In_727);
nand U110 (N_110,In_277,In_987);
and U111 (N_111,In_895,In_4);
nor U112 (N_112,In_1298,In_195);
or U113 (N_113,In_456,In_1034);
or U114 (N_114,In_1470,In_1177);
and U115 (N_115,In_576,In_1243);
nand U116 (N_116,In_942,In_315);
and U117 (N_117,In_832,In_405);
or U118 (N_118,In_1485,In_904);
or U119 (N_119,In_779,In_1086);
and U120 (N_120,In_1428,In_75);
xor U121 (N_121,In_616,In_1483);
nor U122 (N_122,In_953,In_619);
and U123 (N_123,In_228,In_997);
and U124 (N_124,In_1268,In_413);
and U125 (N_125,In_965,In_208);
nand U126 (N_126,In_962,In_1279);
nor U127 (N_127,In_1031,In_1056);
nand U128 (N_128,In_1186,In_1080);
and U129 (N_129,In_284,In_724);
xor U130 (N_130,In_741,In_1351);
nor U131 (N_131,In_736,In_608);
xnor U132 (N_132,In_324,In_849);
xor U133 (N_133,In_1096,In_551);
and U134 (N_134,In_448,In_326);
xnor U135 (N_135,In_1408,In_1395);
or U136 (N_136,In_811,In_357);
and U137 (N_137,In_612,In_191);
and U138 (N_138,In_682,In_1105);
or U139 (N_139,In_709,In_1322);
xnor U140 (N_140,In_1493,In_1481);
or U141 (N_141,In_17,In_898);
or U142 (N_142,In_287,In_848);
or U143 (N_143,In_580,In_1161);
and U144 (N_144,In_386,In_605);
nor U145 (N_145,In_362,In_1240);
nand U146 (N_146,In_1285,In_193);
xor U147 (N_147,In_194,In_749);
or U148 (N_148,In_1441,In_766);
xnor U149 (N_149,In_138,In_1019);
and U150 (N_150,In_3,In_223);
nand U151 (N_151,In_575,In_288);
xnor U152 (N_152,In_136,In_678);
nand U153 (N_153,In_1176,In_1316);
nand U154 (N_154,In_82,In_703);
nor U155 (N_155,In_585,In_1159);
nand U156 (N_156,In_745,In_1057);
nand U157 (N_157,In_747,In_1223);
nand U158 (N_158,In_227,In_541);
and U159 (N_159,In_579,In_390);
and U160 (N_160,In_725,In_1076);
nor U161 (N_161,In_802,In_94);
and U162 (N_162,In_19,In_701);
xnor U163 (N_163,In_31,In_746);
xnor U164 (N_164,In_217,In_1131);
nor U165 (N_165,In_1388,In_624);
or U166 (N_166,In_1175,In_240);
or U167 (N_167,In_1209,In_952);
nand U168 (N_168,In_864,In_521);
nand U169 (N_169,In_37,In_1025);
and U170 (N_170,In_96,In_560);
xnor U171 (N_171,In_299,In_190);
nor U172 (N_172,In_317,In_256);
xor U173 (N_173,In_603,In_235);
and U174 (N_174,In_483,In_1457);
and U175 (N_175,In_507,In_1478);
nand U176 (N_176,In_463,In_488);
xnor U177 (N_177,In_651,In_1221);
or U178 (N_178,In_1083,In_178);
and U179 (N_179,In_338,In_1227);
xnor U180 (N_180,In_280,In_1426);
nand U181 (N_181,In_204,In_748);
xor U182 (N_182,In_268,In_329);
or U183 (N_183,In_819,In_111);
xor U184 (N_184,In_189,In_125);
xor U185 (N_185,In_1211,In_844);
nor U186 (N_186,In_1018,In_214);
and U187 (N_187,In_1274,In_1181);
nor U188 (N_188,In_501,In_1259);
and U189 (N_189,In_409,In_314);
or U190 (N_190,In_719,In_1210);
nor U191 (N_191,In_1320,In_1381);
and U192 (N_192,In_1173,In_344);
nand U193 (N_193,In_1380,In_1058);
xnor U194 (N_194,In_689,In_489);
xor U195 (N_195,In_598,In_1224);
nor U196 (N_196,In_1016,In_559);
nor U197 (N_197,In_234,In_1184);
or U198 (N_198,In_236,In_374);
and U199 (N_199,In_1146,In_248);
or U200 (N_200,In_392,In_657);
nand U201 (N_201,In_457,In_406);
nand U202 (N_202,In_101,In_145);
nor U203 (N_203,In_918,In_1030);
nand U204 (N_204,In_797,In_441);
or U205 (N_205,In_592,In_574);
and U206 (N_206,In_1197,In_1392);
or U207 (N_207,In_361,In_229);
nor U208 (N_208,In_1226,In_1147);
or U209 (N_209,In_1213,In_1344);
or U210 (N_210,In_673,In_1212);
nand U211 (N_211,In_52,In_130);
nand U212 (N_212,In_98,In_503);
xor U213 (N_213,In_807,In_1254);
xnor U214 (N_214,In_122,In_812);
and U215 (N_215,In_643,In_1239);
and U216 (N_216,In_732,In_211);
and U217 (N_217,In_290,In_66);
nand U218 (N_218,In_64,In_715);
nor U219 (N_219,In_1497,In_843);
nor U220 (N_220,In_999,In_1253);
and U221 (N_221,In_387,In_54);
or U222 (N_222,In_1052,In_1202);
nand U223 (N_223,In_1222,In_894);
xor U224 (N_224,In_542,In_1472);
or U225 (N_225,In_308,In_90);
nor U226 (N_226,In_866,In_1012);
and U227 (N_227,In_511,In_72);
or U228 (N_228,In_1092,In_1302);
nand U229 (N_229,In_705,In_92);
xor U230 (N_230,In_1313,In_310);
xor U231 (N_231,In_470,In_1238);
or U232 (N_232,In_637,In_726);
nor U233 (N_233,In_1093,In_1376);
nor U234 (N_234,In_182,In_1138);
nand U235 (N_235,In_638,In_890);
xnor U236 (N_236,In_912,In_1219);
or U237 (N_237,In_1015,In_671);
nor U238 (N_238,In_845,In_1060);
or U239 (N_239,In_1366,In_691);
nor U240 (N_240,In_1263,In_963);
or U241 (N_241,In_582,In_139);
or U242 (N_242,In_345,In_646);
nor U243 (N_243,In_599,In_1251);
xnor U244 (N_244,In_1178,In_1325);
or U245 (N_245,In_1373,In_1050);
and U246 (N_246,In_1283,In_1091);
nor U247 (N_247,In_1062,In_631);
or U248 (N_248,In_723,In_220);
and U249 (N_249,In_635,In_436);
nor U250 (N_250,In_1494,In_1192);
and U251 (N_251,In_972,In_547);
nor U252 (N_252,In_698,In_333);
and U253 (N_253,In_781,In_558);
and U254 (N_254,In_951,In_313);
and U255 (N_255,In_1409,In_931);
or U256 (N_256,In_1498,In_261);
nor U257 (N_257,In_640,In_1260);
and U258 (N_258,In_519,In_595);
nand U259 (N_259,In_971,In_380);
nor U260 (N_260,In_654,In_578);
xor U261 (N_261,In_137,In_1135);
nor U262 (N_262,In_859,In_1010);
nor U263 (N_263,In_399,In_922);
nor U264 (N_264,In_570,In_791);
xor U265 (N_265,In_908,In_1167);
and U266 (N_266,In_920,In_1486);
nor U267 (N_267,In_1479,In_1098);
xnor U268 (N_268,In_788,In_258);
xnor U269 (N_269,In_481,In_1336);
or U270 (N_270,In_1001,In_330);
xor U271 (N_271,In_954,In_57);
and U272 (N_272,In_656,In_35);
xnor U273 (N_273,In_597,In_933);
or U274 (N_274,In_243,In_210);
and U275 (N_275,In_460,In_286);
xnor U276 (N_276,In_545,In_593);
xor U277 (N_277,In_897,In_414);
or U278 (N_278,In_989,In_142);
or U279 (N_279,In_633,In_1435);
nor U280 (N_280,In_1134,In_1489);
or U281 (N_281,In_22,In_425);
and U282 (N_282,In_179,In_53);
nand U283 (N_283,In_716,In_1318);
nand U284 (N_284,In_1398,In_1458);
xnor U285 (N_285,In_1277,In_969);
xor U286 (N_286,In_165,In_1415);
and U287 (N_287,In_676,In_1252);
nand U288 (N_288,In_27,In_1371);
and U289 (N_289,In_275,In_739);
nand U290 (N_290,In_1207,In_979);
xor U291 (N_291,In_1011,In_369);
nor U292 (N_292,In_202,In_647);
nor U293 (N_293,In_209,In_515);
and U294 (N_294,In_737,In_1403);
xor U295 (N_295,In_68,In_108);
xor U296 (N_296,In_29,In_244);
nor U297 (N_297,In_1278,In_1115);
nand U298 (N_298,In_1174,In_232);
nand U299 (N_299,In_1201,In_1169);
nand U300 (N_300,N_88,N_284);
nand U301 (N_301,In_700,In_1156);
xnor U302 (N_302,In_239,N_195);
and U303 (N_303,In_563,In_400);
or U304 (N_304,In_571,In_1036);
or U305 (N_305,In_567,In_188);
and U306 (N_306,N_32,N_7);
and U307 (N_307,In_1021,N_200);
nor U308 (N_308,In_63,In_459);
and U309 (N_309,In_995,In_282);
or U310 (N_310,In_1163,In_836);
xor U311 (N_311,In_370,In_588);
xor U312 (N_312,N_140,In_762);
xor U313 (N_313,In_350,In_91);
nand U314 (N_314,N_90,N_136);
xnor U315 (N_315,N_43,In_1281);
nand U316 (N_316,In_1246,In_623);
or U317 (N_317,In_9,In_365);
or U318 (N_318,N_93,N_56);
and U319 (N_319,N_76,N_13);
nand U320 (N_320,In_1151,In_878);
nand U321 (N_321,In_442,In_1264);
xnor U322 (N_322,In_823,In_1312);
nand U323 (N_323,In_690,In_561);
nor U324 (N_324,In_752,In_1114);
or U325 (N_325,In_1496,N_27);
and U326 (N_326,N_154,In_1101);
nor U327 (N_327,In_1155,In_921);
nand U328 (N_328,In_517,In_249);
nand U329 (N_329,In_135,In_761);
and U330 (N_330,In_611,In_546);
nand U331 (N_331,In_549,In_1124);
or U332 (N_332,N_165,N_221);
and U333 (N_333,In_300,In_1108);
xnor U334 (N_334,In_484,In_1204);
and U335 (N_335,In_439,N_170);
nor U336 (N_336,N_191,N_10);
xor U337 (N_337,In_1049,In_469);
or U338 (N_338,In_816,In_548);
nor U339 (N_339,N_156,In_412);
or U340 (N_340,N_261,In_1007);
nand U341 (N_341,In_385,N_83);
or U342 (N_342,N_141,In_617);
or U343 (N_343,In_465,In_1112);
nand U344 (N_344,In_444,In_391);
and U345 (N_345,N_163,In_1225);
or U346 (N_346,N_73,N_180);
nor U347 (N_347,In_783,N_67);
xor U348 (N_348,In_289,N_58);
nor U349 (N_349,In_80,In_26);
xnor U350 (N_350,In_1334,In_1389);
or U351 (N_351,In_1153,In_1073);
or U352 (N_352,N_131,In_846);
nand U353 (N_353,In_1314,In_1061);
nand U354 (N_354,In_874,In_993);
xnor U355 (N_355,N_197,In_218);
nor U356 (N_356,In_397,In_410);
nor U357 (N_357,In_134,In_1013);
nor U358 (N_358,N_212,In_1249);
or U359 (N_359,In_447,In_1208);
nand U360 (N_360,In_784,In_685);
nand U361 (N_361,N_133,In_451);
nor U362 (N_362,In_1349,In_1247);
and U363 (N_363,N_142,In_537);
nor U364 (N_364,In_644,In_18);
and U365 (N_365,N_292,In_452);
or U366 (N_366,In_937,In_1300);
nand U367 (N_367,N_169,In_763);
nand U368 (N_368,In_786,In_113);
nand U369 (N_369,N_230,In_1273);
nor U370 (N_370,In_85,In_364);
xnor U371 (N_371,In_888,In_1029);
xor U372 (N_372,N_41,In_1044);
or U373 (N_373,N_295,In_530);
nand U374 (N_374,In_246,In_693);
nor U375 (N_375,In_1140,In_1048);
and U376 (N_376,In_929,In_1437);
nand U377 (N_377,In_1372,In_1459);
nand U378 (N_378,In_104,In_564);
xnor U379 (N_379,In_1121,In_932);
nor U380 (N_380,In_1377,In_1172);
xor U381 (N_381,In_1327,In_935);
and U382 (N_382,In_688,In_69);
xor U383 (N_383,In_283,N_188);
and U384 (N_384,N_35,In_1348);
nand U385 (N_385,In_707,N_79);
nor U386 (N_386,N_196,In_1271);
or U387 (N_387,In_911,In_1480);
xnor U388 (N_388,In_166,In_320);
xor U389 (N_389,N_171,In_642);
xnor U390 (N_390,N_273,N_247);
xnor U391 (N_391,N_246,In_1203);
and U392 (N_392,In_877,N_66);
nand U393 (N_393,In_1104,In_1288);
and U394 (N_394,In_292,In_769);
and U395 (N_395,In_1378,N_143);
or U396 (N_396,N_104,In_1464);
nor U397 (N_397,In_403,In_1168);
xnor U398 (N_398,N_152,In_927);
or U399 (N_399,In_712,In_312);
xnor U400 (N_400,In_1187,N_270);
and U401 (N_401,N_289,In_440);
nand U402 (N_402,In_1040,In_155);
or U403 (N_403,In_296,In_159);
nand U404 (N_404,In_957,In_349);
nand U405 (N_405,In_839,In_434);
or U406 (N_406,In_100,In_1200);
nand U407 (N_407,In_1374,In_148);
nand U408 (N_408,In_1148,N_106);
nor U409 (N_409,In_423,In_119);
xnor U410 (N_410,In_254,N_118);
or U411 (N_411,In_1136,In_260);
and U412 (N_412,In_529,In_34);
and U413 (N_413,In_1244,In_847);
xor U414 (N_414,In_662,In_267);
nor U415 (N_415,In_944,N_126);
and U416 (N_416,N_42,In_33);
nor U417 (N_417,In_1333,In_372);
nor U418 (N_418,In_177,N_29);
or U419 (N_419,In_508,In_1303);
or U420 (N_420,In_321,In_379);
or U421 (N_421,In_1017,In_272);
and U422 (N_422,In_59,In_494);
xnor U423 (N_423,N_14,N_81);
or U424 (N_424,N_241,N_294);
xor U425 (N_425,In_799,In_509);
or U426 (N_426,In_474,In_573);
nor U427 (N_427,N_45,In_1422);
or U428 (N_428,In_1342,N_281);
or U429 (N_429,In_853,N_291);
xnor U430 (N_430,N_12,N_272);
xnor U431 (N_431,In_114,In_1319);
and U432 (N_432,In_183,In_1129);
xor U433 (N_433,In_525,N_147);
nor U434 (N_434,In_309,In_1326);
nor U435 (N_435,N_250,In_87);
xnor U436 (N_436,In_1332,In_40);
xor U437 (N_437,In_196,In_557);
and U438 (N_438,In_860,N_185);
nand U439 (N_439,In_994,In_1078);
nand U440 (N_440,In_224,In_1362);
nand U441 (N_441,In_1054,N_211);
nor U442 (N_442,In_461,In_132);
nor U443 (N_443,In_259,In_913);
and U444 (N_444,N_122,In_1495);
xor U445 (N_445,In_950,In_632);
or U446 (N_446,N_245,In_1119);
nand U447 (N_447,In_1431,N_276);
and U448 (N_448,N_264,N_251);
and U449 (N_449,N_127,N_189);
xor U450 (N_450,In_1357,N_112);
xor U451 (N_451,In_661,N_124);
xor U452 (N_452,In_672,In_107);
nor U453 (N_453,In_1206,N_249);
nor U454 (N_454,In_1248,N_19);
or U455 (N_455,In_645,In_622);
nor U456 (N_456,In_433,In_626);
or U457 (N_457,In_168,N_204);
nand U458 (N_458,In_1055,N_297);
nand U459 (N_459,In_482,In_212);
nand U460 (N_460,N_62,In_174);
nor U461 (N_461,In_714,In_162);
xor U462 (N_462,In_201,In_25);
or U463 (N_463,In_1305,In_1069);
nor U464 (N_464,In_1469,N_4);
xor U465 (N_465,In_322,In_1166);
or U466 (N_466,In_868,N_225);
xor U467 (N_467,In_294,In_659);
nand U468 (N_468,In_875,In_62);
nor U469 (N_469,In_706,N_207);
nor U470 (N_470,In_295,N_107);
or U471 (N_471,N_116,In_751);
and U472 (N_472,In_586,In_1484);
xnor U473 (N_473,In_892,In_591);
xnor U474 (N_474,In_1488,In_1215);
and U475 (N_475,In_432,In_1359);
or U476 (N_476,In_893,In_928);
xnor U477 (N_477,In_238,In_758);
nand U478 (N_478,In_1158,In_301);
or U479 (N_479,In_1180,In_841);
and U480 (N_480,In_279,In_792);
nand U481 (N_481,In_213,In_1022);
or U482 (N_482,In_41,N_176);
xor U483 (N_483,In_1282,In_872);
or U484 (N_484,In_917,In_854);
and U485 (N_485,N_259,In_734);
and U486 (N_486,N_17,In_144);
and U487 (N_487,N_227,N_172);
and U488 (N_488,In_677,In_354);
nand U489 (N_489,N_82,N_193);
nor U490 (N_490,In_499,In_21);
xnor U491 (N_491,In_163,In_486);
xnor U492 (N_492,N_206,In_735);
and U493 (N_493,In_641,In_1152);
or U494 (N_494,In_1003,In_851);
nand U495 (N_495,N_216,In_787);
nor U496 (N_496,In_1063,In_226);
nand U497 (N_497,In_445,In_1084);
or U498 (N_498,In_589,In_1364);
nor U499 (N_499,In_800,N_239);
nor U500 (N_500,N_153,In_71);
or U501 (N_501,In_1476,N_265);
xor U502 (N_502,In_721,In_858);
and U503 (N_503,In_305,In_110);
or U504 (N_504,In_808,In_1445);
and U505 (N_505,In_1391,In_473);
xor U506 (N_506,N_20,N_24);
xor U507 (N_507,In_1330,In_1487);
nand U508 (N_508,In_900,In_1448);
and U509 (N_509,N_215,In_581);
or U510 (N_510,In_167,In_533);
or U511 (N_511,In_1006,In_342);
and U512 (N_512,In_961,In_1143);
nor U513 (N_513,In_902,In_1068);
nand U514 (N_514,N_25,In_44);
nand U515 (N_515,In_772,In_311);
or U516 (N_516,In_421,In_1165);
and U517 (N_517,In_905,N_285);
or U518 (N_518,In_1468,In_1429);
nand U519 (N_519,In_668,N_44);
and U520 (N_520,In_11,In_97);
xor U521 (N_521,In_958,In_366);
nor U522 (N_522,In_683,N_123);
and U523 (N_523,In_544,In_1154);
xnor U524 (N_524,In_527,In_1407);
or U525 (N_525,In_118,In_378);
xor U526 (N_526,In_206,In_1455);
xor U527 (N_527,N_128,In_840);
or U528 (N_528,N_162,In_269);
xnor U529 (N_529,N_108,In_340);
or U530 (N_530,In_358,In_30);
nor U531 (N_531,N_296,In_32);
and U532 (N_532,In_225,In_1009);
or U533 (N_533,N_248,In_1245);
nor U534 (N_534,In_584,In_192);
xor U535 (N_535,In_704,In_1074);
nor U536 (N_536,N_59,In_1130);
xor U537 (N_537,N_235,In_1047);
xor U538 (N_538,N_0,In_1420);
xnor U539 (N_539,In_496,In_341);
xor U540 (N_540,In_826,In_416);
and U541 (N_541,In_1042,N_18);
nor U542 (N_542,In_1375,In_634);
xor U543 (N_543,In_606,N_268);
nand U544 (N_544,In_1195,In_1046);
xnor U545 (N_545,In_437,In_583);
nor U546 (N_546,In_1237,In_323);
and U547 (N_547,N_37,In_1232);
nor U548 (N_548,N_11,In_1482);
or U549 (N_549,N_155,N_262);
nand U550 (N_550,N_63,N_208);
or U551 (N_551,In_1113,In_924);
xnor U552 (N_552,In_1355,N_22);
nor U553 (N_553,In_1404,In_828);
xor U554 (N_554,N_223,In_180);
and U555 (N_555,In_804,In_1418);
and U556 (N_556,N_49,In_1149);
nor U557 (N_557,In_222,N_217);
and U558 (N_558,In_200,In_837);
or U559 (N_559,In_1065,In_536);
nor U560 (N_560,In_1144,In_1307);
and U561 (N_561,In_665,N_6);
xnor U562 (N_562,In_984,In_814);
nand U563 (N_563,In_553,N_137);
or U564 (N_564,In_556,N_202);
nand U565 (N_565,In_722,In_13);
nand U566 (N_566,N_77,In_601);
nand U567 (N_567,In_231,In_426);
or U568 (N_568,N_115,In_70);
xor U569 (N_569,In_1241,N_51);
and U570 (N_570,N_219,N_102);
and U571 (N_571,N_47,In_1309);
xnor U572 (N_572,N_120,In_639);
xnor U573 (N_573,In_1290,N_95);
or U574 (N_574,In_83,N_298);
and U575 (N_575,In_562,In_711);
or U576 (N_576,In_16,N_64);
nor U577 (N_577,In_1284,In_274);
and U578 (N_578,In_1110,N_65);
nand U579 (N_579,N_275,In_120);
nand U580 (N_580,In_348,In_367);
xor U581 (N_581,In_14,N_125);
or U582 (N_582,In_1261,In_1111);
nand U583 (N_583,N_28,N_151);
nand U584 (N_584,N_30,In_298);
or U585 (N_585,In_1365,In_492);
nor U586 (N_586,In_184,In_147);
xor U587 (N_587,In_418,In_1014);
nand U588 (N_588,In_755,In_490);
xor U589 (N_589,N_114,In_247);
xor U590 (N_590,N_38,In_1411);
and U591 (N_591,In_164,In_88);
nor U592 (N_592,In_862,N_69);
nand U593 (N_593,In_99,In_115);
or U594 (N_594,In_1081,In_464);
and U595 (N_595,In_680,N_236);
or U596 (N_596,In_1000,In_960);
and U597 (N_597,N_199,In_1440);
and U598 (N_598,In_109,In_293);
xor U599 (N_599,In_879,In_1217);
and U600 (N_600,In_1396,N_383);
or U601 (N_601,In_830,In_1039);
and U602 (N_602,In_1280,In_334);
or U603 (N_603,N_220,N_557);
xnor U604 (N_604,In_1306,In_273);
or U605 (N_605,In_941,N_362);
and U606 (N_606,N_594,N_1);
and U607 (N_607,N_414,N_307);
and U608 (N_608,N_585,N_425);
or U609 (N_609,N_559,In_760);
or U610 (N_610,N_316,In_687);
nand U611 (N_611,In_393,N_483);
xnor U612 (N_612,N_543,N_564);
or U613 (N_613,N_74,N_121);
nand U614 (N_614,N_537,In_982);
or U615 (N_615,In_176,N_554);
and U616 (N_616,In_187,N_228);
nor U617 (N_617,In_1352,In_270);
nor U618 (N_618,N_87,In_1128);
and U619 (N_619,In_628,N_139);
and U620 (N_620,N_214,In_618);
xor U621 (N_621,N_203,In_1100);
nor U622 (N_622,N_263,In_1194);
and U623 (N_623,N_492,In_1041);
nor U624 (N_624,In_827,N_462);
nand U625 (N_625,N_591,In_1439);
and U626 (N_626,N_509,In_822);
or U627 (N_627,N_504,In_750);
or U628 (N_628,In_649,In_1258);
nor U629 (N_629,N_570,N_198);
nor U630 (N_630,In_281,In_1);
nand U631 (N_631,In_360,N_55);
or U632 (N_632,N_513,N_86);
xor U633 (N_633,N_105,N_448);
nand U634 (N_634,In_697,In_510);
nand U635 (N_635,In_988,N_562);
xnor U636 (N_636,In_411,In_297);
and U637 (N_637,N_407,In_1276);
nor U638 (N_638,In_855,In_945);
nor U639 (N_639,N_532,In_663);
or U640 (N_640,In_1419,N_103);
xnor U641 (N_641,N_571,In_1275);
xnor U642 (N_642,N_326,N_333);
nor U643 (N_643,In_264,In_590);
and U644 (N_644,N_387,In_1370);
nor U645 (N_645,In_1462,N_338);
and U646 (N_646,In_86,N_381);
nand U647 (N_647,In_850,N_368);
nor U648 (N_648,In_742,N_369);
nand U649 (N_649,In_203,In_1417);
or U650 (N_650,N_302,In_1266);
nand U651 (N_651,N_237,In_1107);
nor U652 (N_652,In_1103,In_896);
or U653 (N_653,N_377,N_517);
nor U654 (N_654,N_472,In_964);
and U655 (N_655,In_720,In_1033);
and U656 (N_656,N_502,In_532);
xnor U657 (N_657,N_413,N_382);
xnor U658 (N_658,N_468,N_441);
or U659 (N_659,In_815,In_1367);
nor U660 (N_660,N_466,N_342);
nor U661 (N_661,In_610,N_205);
nand U662 (N_662,In_738,In_764);
and U663 (N_663,N_288,N_53);
and U664 (N_664,In_117,In_408);
or U665 (N_665,N_488,In_824);
nor U666 (N_666,N_346,In_1399);
xnor U667 (N_667,In_127,In_458);
nand U668 (N_668,In_133,In_1189);
and U669 (N_669,In_1199,N_356);
nand U670 (N_670,N_315,N_555);
nand U671 (N_671,N_395,N_563);
xor U672 (N_672,In_513,N_380);
nor U673 (N_673,N_339,N_224);
or U674 (N_674,N_160,N_506);
or U675 (N_675,In_821,N_523);
and U676 (N_676,N_218,N_75);
xnor U677 (N_677,In_428,In_1421);
nor U678 (N_678,In_1265,In_870);
xor U679 (N_679,N_351,N_486);
nor U680 (N_680,N_187,In_810);
xnor U681 (N_681,In_1087,In_1430);
nand U682 (N_682,In_1347,N_447);
and U683 (N_683,N_491,N_129);
and U684 (N_684,N_580,In_955);
nand U685 (N_685,N_98,In_291);
nor U686 (N_686,In_468,In_377);
and U687 (N_687,In_140,In_873);
nor U688 (N_688,N_310,N_416);
nand U689 (N_689,N_23,N_91);
or U690 (N_690,In_543,In_351);
nand U691 (N_691,In_852,In_407);
or U692 (N_692,N_283,In_480);
or U693 (N_693,N_375,N_231);
or U694 (N_694,N_402,N_135);
and U695 (N_695,N_560,In_594);
and U696 (N_696,In_478,N_391);
nor U697 (N_697,In_600,In_1171);
nor U698 (N_698,N_438,N_490);
nand U699 (N_699,In_903,N_460);
xor U700 (N_700,N_400,In_1383);
nand U701 (N_701,N_399,In_777);
nor U702 (N_702,N_54,In_798);
or U703 (N_703,N_430,N_595);
or U704 (N_704,In_565,N_344);
xnor U705 (N_705,In_1412,N_109);
and U706 (N_706,In_524,In_23);
and U707 (N_707,In_1452,In_28);
xnor U708 (N_708,In_58,N_432);
nand U709 (N_709,N_279,In_1339);
nor U710 (N_710,In_1384,N_252);
or U711 (N_711,In_790,In_1475);
and U712 (N_712,N_92,N_545);
and U713 (N_713,N_327,In_655);
xnor U714 (N_714,In_956,N_159);
and U715 (N_715,In_398,In_1123);
nand U716 (N_716,N_280,In_36);
and U717 (N_717,N_94,In_1051);
xnor U718 (N_718,N_145,In_1304);
and U719 (N_719,In_1231,N_436);
xor U720 (N_720,N_319,N_524);
or U721 (N_721,N_324,In_173);
and U722 (N_722,In_538,In_316);
xor U723 (N_723,N_100,In_1397);
or U724 (N_724,In_1170,N_5);
nor U725 (N_725,In_731,N_520);
nor U726 (N_726,In_6,N_321);
nand U727 (N_727,N_577,N_183);
or U728 (N_728,In_415,In_625);
or U729 (N_729,N_579,In_717);
xnor U730 (N_730,N_458,N_325);
and U731 (N_731,N_452,In_5);
or U732 (N_732,N_359,In_157);
nor U733 (N_733,N_385,In_658);
or U734 (N_734,N_164,In_60);
and U735 (N_735,In_817,N_406);
xor U736 (N_736,N_372,In_670);
or U737 (N_737,N_299,In_20);
nand U738 (N_738,N_464,N_16);
and U739 (N_739,N_522,In_1473);
and U740 (N_740,N_179,N_161);
or U741 (N_741,N_113,In_1368);
xor U742 (N_742,In_795,N_192);
xor U743 (N_743,N_158,In_476);
xor U744 (N_744,In_1085,In_1095);
nand U745 (N_745,In_1032,In_1028);
xor U746 (N_746,N_593,N_511);
nor U747 (N_747,N_348,N_444);
nand U748 (N_748,N_434,In_215);
nor U749 (N_749,N_455,N_499);
and U750 (N_750,N_61,In_959);
nand U751 (N_751,N_15,N_393);
nand U752 (N_752,In_729,N_478);
nand U753 (N_753,N_361,N_345);
nand U754 (N_754,In_368,In_1125);
or U755 (N_755,In_1299,N_363);
nand U756 (N_756,In_865,N_213);
or U757 (N_757,In_773,N_255);
xnor U758 (N_758,N_487,N_417);
nand U759 (N_759,In_614,In_116);
nor U760 (N_760,In_949,In_554);
nand U761 (N_761,In_660,In_455);
nor U762 (N_762,N_515,In_514);
nand U763 (N_763,N_415,In_796);
nand U764 (N_764,N_548,In_666);
and U765 (N_765,N_508,In_79);
and U766 (N_766,In_1295,N_445);
xnor U767 (N_767,In_376,N_148);
and U768 (N_768,N_8,In_230);
nor U769 (N_769,N_232,N_467);
or U770 (N_770,In_375,In_980);
xor U771 (N_771,N_349,In_1466);
or U772 (N_772,In_1064,In_1077);
nand U773 (N_773,N_489,In_1401);
nor U774 (N_774,N_598,N_493);
nor U775 (N_775,In_128,In_818);
or U776 (N_776,N_238,In_914);
and U777 (N_777,N_586,In_1446);
or U778 (N_778,In_756,In_771);
nor U779 (N_779,In_172,In_55);
or U780 (N_780,N_328,In_1053);
or U781 (N_781,In_1141,In_252);
or U782 (N_782,N_335,In_1447);
or U783 (N_783,N_446,In_1345);
or U784 (N_784,In_923,N_456);
or U785 (N_785,In_93,In_171);
xor U786 (N_786,In_910,N_552);
nand U787 (N_787,N_599,N_269);
nor U788 (N_788,In_1193,N_34);
or U789 (N_789,N_388,In_992);
and U790 (N_790,N_427,N_461);
nor U791 (N_791,N_510,In_149);
nand U792 (N_792,In_861,In_84);
nand U793 (N_793,In_1024,In_1323);
xnor U794 (N_794,In_744,In_1297);
and U795 (N_795,In_233,N_130);
nand U796 (N_796,N_497,In_497);
nor U797 (N_797,In_871,N_366);
nand U798 (N_798,In_1198,In_382);
xor U799 (N_799,In_1382,In_76);
xnor U800 (N_800,N_309,In_765);
and U801 (N_801,N_479,In_466);
nor U802 (N_802,In_237,In_531);
and U803 (N_803,In_491,N_556);
or U804 (N_804,In_307,N_551);
xnor U805 (N_805,N_186,In_1338);
nor U806 (N_806,N_566,N_21);
nand U807 (N_807,N_3,N_306);
and U808 (N_808,In_47,N_561);
nand U809 (N_809,In_540,In_1317);
or U810 (N_810,In_1471,In_395);
nand U811 (N_811,In_1139,In_880);
nand U812 (N_812,N_166,N_553);
and U813 (N_813,N_409,In_757);
xnor U814 (N_814,N_132,In_431);
nand U815 (N_815,N_494,N_168);
xor U816 (N_816,N_226,In_780);
and U817 (N_817,N_449,N_512);
and U818 (N_818,N_150,N_260);
or U819 (N_819,In_485,N_39);
nor U820 (N_820,N_244,N_442);
nor U821 (N_821,In_696,In_794);
xnor U822 (N_822,N_450,N_533);
and U823 (N_823,In_838,N_111);
xor U824 (N_824,N_394,In_679);
xor U825 (N_825,N_470,In_1491);
nand U826 (N_826,N_290,In_976);
nor U827 (N_827,In_968,In_242);
and U828 (N_828,N_209,N_174);
nor U829 (N_829,N_429,N_48);
and U830 (N_830,In_1361,In_1454);
nor U831 (N_831,In_89,In_221);
nor U832 (N_832,N_419,N_519);
nor U833 (N_833,In_754,In_753);
xor U834 (N_834,In_1008,In_477);
and U835 (N_835,In_0,N_78);
xor U836 (N_836,In_710,N_330);
nor U837 (N_837,In_435,N_347);
and U838 (N_838,N_482,In_181);
and U839 (N_839,N_389,In_919);
and U840 (N_840,In_1142,N_542);
or U841 (N_841,N_329,N_80);
nor U842 (N_842,In_967,N_587);
and U843 (N_843,N_474,In_1106);
xnor U844 (N_844,N_36,In_857);
or U845 (N_845,In_1230,N_317);
xnor U846 (N_846,N_451,In_699);
nand U847 (N_847,In_505,In_926);
nor U848 (N_848,In_262,In_977);
xor U849 (N_849,N_424,N_40);
nand U850 (N_850,In_983,N_463);
nor U851 (N_851,N_352,In_105);
xor U852 (N_852,In_219,In_343);
nor U853 (N_853,N_398,N_536);
xnor U854 (N_854,N_96,In_302);
and U855 (N_855,N_313,N_340);
or U856 (N_856,N_374,N_146);
nand U857 (N_857,N_596,In_383);
nand U858 (N_858,N_287,In_1394);
xor U859 (N_859,In_1402,In_363);
nor U860 (N_860,N_157,N_473);
nor U861 (N_861,In_199,In_462);
xor U862 (N_862,N_392,N_574);
or U863 (N_863,In_522,In_303);
and U864 (N_864,N_350,N_360);
nand U865 (N_865,N_404,In_50);
or U866 (N_866,N_234,In_121);
nor U867 (N_867,N_89,In_730);
nand U868 (N_868,In_48,In_141);
nor U869 (N_869,In_806,N_282);
xor U870 (N_870,In_73,N_84);
nor U871 (N_871,N_355,N_274);
nand U872 (N_872,N_527,N_516);
and U873 (N_873,In_1133,N_567);
and U874 (N_874,N_278,N_526);
xnor U875 (N_875,In_250,N_343);
and U876 (N_876,N_97,N_439);
nor U877 (N_877,In_1424,In_1385);
and U878 (N_878,In_46,N_433);
and U879 (N_879,In_1150,N_459);
xnor U880 (N_880,N_412,N_33);
and U881 (N_881,N_314,N_341);
or U882 (N_882,N_465,In_1035);
nor U883 (N_883,In_1449,In_718);
nand U884 (N_884,N_332,N_367);
xor U885 (N_885,N_194,In_419);
nor U886 (N_886,In_925,In_1301);
and U887 (N_887,In_692,In_863);
xor U888 (N_888,In_1292,N_254);
or U889 (N_889,In_973,N_371);
nand U890 (N_890,In_831,N_364);
and U891 (N_891,N_311,N_379);
nor U892 (N_892,In_834,N_201);
or U893 (N_893,In_770,In_78);
nand U894 (N_894,In_885,N_437);
xor U895 (N_895,In_1043,In_991);
nand U896 (N_896,In_15,In_95);
nor U897 (N_897,N_322,N_401);
nand U898 (N_898,In_1020,In_67);
nor U899 (N_899,In_1442,N_453);
nor U900 (N_900,N_578,N_318);
xnor U901 (N_901,N_806,In_1477);
nand U902 (N_902,N_184,In_805);
nand U903 (N_903,N_761,N_897);
xor U904 (N_904,N_810,N_711);
nand U905 (N_905,N_657,N_378);
nor U906 (N_906,In_319,In_1427);
and U907 (N_907,N_681,N_805);
xor U908 (N_908,In_278,N_633);
nor U909 (N_909,N_708,N_850);
and U910 (N_910,N_669,N_614);
nor U911 (N_911,N_426,N_786);
nand U912 (N_912,N_167,N_610);
xor U913 (N_913,N_778,N_420);
nand U914 (N_914,In_1220,N_480);
xor U915 (N_915,N_619,In_446);
and U916 (N_916,N_210,N_688);
and U917 (N_917,N_550,N_797);
or U918 (N_918,N_606,In_1005);
xor U919 (N_919,N_767,N_788);
nor U920 (N_920,In_1443,In_1467);
or U921 (N_921,In_940,In_1256);
nor U922 (N_922,In_49,N_624);
and U923 (N_923,N_660,N_791);
xnor U924 (N_924,In_1444,N_878);
or U925 (N_925,N_46,In_131);
and U926 (N_926,In_778,N_883);
nand U927 (N_927,N_719,N_655);
and U928 (N_928,N_645,N_881);
or U929 (N_929,N_770,N_809);
and U930 (N_930,N_588,N_754);
and U931 (N_931,In_1004,N_626);
or U932 (N_932,In_694,N_469);
xor U933 (N_933,N_884,N_741);
xnor U934 (N_934,In_1270,N_410);
xor U935 (N_935,N_757,In_1329);
and U936 (N_936,N_531,In_1400);
and U937 (N_937,N_825,N_484);
xnor U938 (N_938,N_304,In_930);
nand U939 (N_939,In_516,In_151);
xor U940 (N_940,N_780,N_738);
nand U941 (N_941,N_609,N_530);
or U942 (N_942,N_589,N_846);
and U943 (N_943,In_1205,In_216);
nor U944 (N_944,N_683,In_674);
and U945 (N_945,N_686,N_707);
nor U946 (N_946,N_827,N_838);
nand U947 (N_947,N_431,In_347);
xnor U948 (N_948,N_665,In_336);
or U949 (N_949,N_411,N_743);
and U950 (N_950,In_1328,In_825);
nand U951 (N_951,N_898,N_869);
nor U952 (N_952,N_501,N_783);
nand U953 (N_953,N_173,N_829);
nor U954 (N_954,N_454,N_749);
or U955 (N_955,In_1102,N_177);
xnor U956 (N_956,N_569,N_572);
and U957 (N_957,N_664,N_811);
nor U958 (N_958,N_408,N_576);
xnor U959 (N_959,N_744,N_751);
and U960 (N_960,N_632,In_1296);
nand U961 (N_961,N_676,N_784);
nor U962 (N_962,N_857,N_608);
and U963 (N_963,N_613,N_766);
nor U964 (N_964,N_842,In_1272);
and U965 (N_965,In_1343,N_390);
and U966 (N_966,In_889,N_618);
xor U967 (N_967,N_540,N_758);
nor U968 (N_968,N_734,N_286);
xnor U969 (N_969,In_45,In_1229);
nand U970 (N_970,In_1414,N_724);
or U971 (N_971,N_423,N_649);
nor U972 (N_972,N_695,N_860);
nor U973 (N_973,N_485,In_56);
or U974 (N_974,N_752,N_776);
nand U975 (N_975,In_112,N_405);
nand U976 (N_976,N_885,N_746);
xor U977 (N_977,N_726,N_182);
xor U978 (N_978,N_768,N_354);
and U979 (N_979,N_175,N_888);
xor U980 (N_980,N_243,N_815);
or U981 (N_981,N_833,N_320);
and U982 (N_982,N_590,N_795);
nor U983 (N_983,N_856,N_762);
xnor U984 (N_984,In_512,N_617);
nand U985 (N_985,In_353,In_1463);
nand U986 (N_986,N_643,In_152);
nor U987 (N_987,In_1308,N_803);
nand U988 (N_988,N_841,N_721);
or U989 (N_989,In_205,N_661);
nor U990 (N_990,In_947,N_547);
or U991 (N_991,N_772,N_773);
nand U992 (N_992,N_634,N_134);
nand U993 (N_993,N_861,N_774);
and U994 (N_994,N_854,In_402);
and U995 (N_995,N_222,N_877);
nor U996 (N_996,N_706,N_687);
nand U997 (N_997,N_794,N_812);
and U998 (N_998,N_895,In_1341);
and U999 (N_999,N_740,N_759);
or U1000 (N_1000,N_421,In_785);
nor U1001 (N_1001,N_828,N_853);
nand U1002 (N_1002,N_514,N_300);
nand U1003 (N_1003,N_498,N_575);
or U1004 (N_1004,In_1099,N_60);
nand U1005 (N_1005,N_495,N_832);
nor U1006 (N_1006,N_745,N_779);
nand U1007 (N_1007,N_808,N_673);
nand U1008 (N_1008,In_702,In_1216);
or U1009 (N_1009,In_146,In_253);
and U1010 (N_1010,N_851,In_1324);
xor U1011 (N_1011,N_521,N_879);
and U1012 (N_1012,In_265,N_790);
nor U1013 (N_1013,N_813,N_696);
xnor U1014 (N_1014,N_600,N_544);
or U1015 (N_1015,In_449,N_682);
nand U1016 (N_1016,N_739,N_691);
nand U1017 (N_1017,In_495,N_871);
and U1018 (N_1018,N_685,N_893);
xnor U1019 (N_1019,N_804,In_401);
nor U1020 (N_1020,In_1360,N_777);
nor U1021 (N_1021,N_365,In_450);
nand U1022 (N_1022,N_736,N_693);
xnor U1023 (N_1023,N_271,N_144);
or U1024 (N_1024,N_709,N_820);
or U1025 (N_1025,In_373,N_680);
nand U1026 (N_1026,N_558,In_621);
and U1027 (N_1027,N_612,N_865);
nor U1028 (N_1028,N_679,In_1126);
or U1029 (N_1029,In_424,N_240);
nand U1030 (N_1030,N_830,N_831);
and U1031 (N_1031,N_892,N_714);
nand U1032 (N_1032,N_336,N_859);
nand U1033 (N_1033,In_170,N_638);
and U1034 (N_1034,N_755,In_833);
and U1035 (N_1035,In_789,In_1289);
nand U1036 (N_1036,N_789,N_764);
nand U1037 (N_1037,N_821,N_800);
or U1038 (N_1038,N_763,N_722);
nor U1039 (N_1039,N_622,In_523);
nor U1040 (N_1040,N_640,N_525);
nor U1041 (N_1041,N_658,In_906);
nand U1042 (N_1042,In_669,N_443);
nand U1043 (N_1043,N_9,N_698);
and U1044 (N_1044,In_1164,N_2);
nand U1045 (N_1045,N_847,N_796);
nand U1046 (N_1046,N_697,N_376);
nor U1047 (N_1047,N_475,N_704);
and U1048 (N_1048,N_644,N_656);
nand U1049 (N_1049,In_650,N_592);
xor U1050 (N_1050,N_720,N_358);
or U1051 (N_1051,N_500,N_886);
and U1052 (N_1052,In_1474,N_597);
nor U1053 (N_1053,N_541,N_546);
or U1054 (N_1054,In_1038,In_1218);
nand U1055 (N_1055,In_1499,N_816);
nand U1056 (N_1056,N_735,N_650);
and U1057 (N_1057,N_257,N_627);
and U1058 (N_1058,N_99,In_648);
xnor U1059 (N_1059,N_712,N_647);
nor U1060 (N_1060,N_242,N_801);
nand U1061 (N_1061,N_119,In_396);
nand U1062 (N_1062,N_57,N_642);
nor U1063 (N_1063,N_689,In_1461);
or U1064 (N_1064,In_1335,N_277);
or U1065 (N_1065,N_864,N_601);
nor U1066 (N_1066,N_611,N_384);
xnor U1067 (N_1067,N_666,N_403);
nor U1068 (N_1068,N_616,N_872);
nand U1069 (N_1069,N_68,N_357);
or U1070 (N_1070,N_716,N_457);
and U1071 (N_1071,N_615,In_504);
or U1072 (N_1072,N_675,N_435);
nand U1073 (N_1073,N_573,N_715);
or U1074 (N_1074,N_737,N_72);
nor U1075 (N_1075,In_528,N_837);
nand U1076 (N_1076,In_975,N_769);
and U1077 (N_1077,N_418,N_713);
and U1078 (N_1078,In_158,N_807);
xnor U1079 (N_1079,N_750,N_890);
nor U1080 (N_1080,N_692,N_646);
and U1081 (N_1081,N_725,In_948);
nand U1082 (N_1082,N_625,N_814);
nand U1083 (N_1083,N_760,N_641);
xnor U1084 (N_1084,N_699,N_568);
and U1085 (N_1085,N_781,N_256);
and U1086 (N_1086,N_710,In_160);
or U1087 (N_1087,N_732,In_1387);
nand U1088 (N_1088,N_659,In_467);
xnor U1089 (N_1089,N_874,N_862);
nand U1090 (N_1090,N_817,In_443);
or U1091 (N_1091,In_1059,N_396);
and U1092 (N_1092,N_181,In_943);
xnor U1093 (N_1093,N_428,N_582);
and U1094 (N_1094,N_742,N_663);
nor U1095 (N_1095,N_765,N_840);
nand U1096 (N_1096,N_476,N_631);
and U1097 (N_1097,N_787,N_305);
nor U1098 (N_1098,N_397,In_627);
nand U1099 (N_1099,N_896,N_621);
and U1100 (N_1100,N_353,N_639);
xor U1101 (N_1101,N_891,In_332);
xor U1102 (N_1102,N_440,N_834);
nand U1103 (N_1103,N_802,N_867);
and U1104 (N_1104,In_1002,In_389);
nand U1105 (N_1105,N_334,N_845);
nor U1106 (N_1106,N_538,In_743);
xnor U1107 (N_1107,N_799,N_528);
nor U1108 (N_1108,N_529,N_694);
xor U1109 (N_1109,N_836,N_700);
or U1110 (N_1110,N_718,N_782);
and U1111 (N_1111,N_826,N_843);
nor U1112 (N_1112,N_775,N_662);
and U1113 (N_1113,N_539,N_668);
nor U1114 (N_1114,N_518,N_233);
nor U1115 (N_1115,N_863,N_727);
nor U1116 (N_1116,N_581,N_635);
nor U1117 (N_1117,In_1315,N_651);
nand U1118 (N_1118,N_337,N_729);
xor U1119 (N_1119,N_31,In_198);
or U1120 (N_1120,N_702,N_672);
and U1121 (N_1121,N_178,In_10);
and U1122 (N_1122,N_705,N_138);
xor U1123 (N_1123,In_1066,N_835);
nor U1124 (N_1124,N_671,N_653);
and U1125 (N_1125,N_747,In_782);
nor U1126 (N_1126,N_50,N_534);
and U1127 (N_1127,N_858,N_267);
nor U1128 (N_1128,N_604,N_756);
or U1129 (N_1129,N_496,N_819);
nand U1130 (N_1130,N_882,N_844);
nand U1131 (N_1131,N_785,In_526);
or U1132 (N_1132,N_701,N_868);
nand U1133 (N_1133,In_1310,N_549);
and U1134 (N_1134,N_583,N_894);
xnor U1135 (N_1135,N_703,N_70);
or U1136 (N_1136,N_602,In_876);
nor U1137 (N_1137,In_1045,N_690);
or U1138 (N_1138,N_748,N_258);
or U1139 (N_1139,N_880,N_229);
and U1140 (N_1140,In_1097,N_110);
xor U1141 (N_1141,N_373,N_730);
xor U1142 (N_1142,N_605,In_566);
and U1143 (N_1143,In_986,N_565);
nor U1144 (N_1144,In_1023,N_422);
or U1145 (N_1145,In_500,N_717);
xor U1146 (N_1146,N_848,N_818);
nand U1147 (N_1147,N_386,In_39);
or U1148 (N_1148,N_677,In_161);
and U1149 (N_1149,N_652,In_978);
xnor U1150 (N_1150,N_678,N_875);
nor U1151 (N_1151,In_1363,N_824);
xnor U1152 (N_1152,In_686,In_143);
nor U1153 (N_1153,N_481,In_65);
or U1154 (N_1154,In_186,In_587);
and U1155 (N_1155,N_607,N_26);
or U1156 (N_1156,N_684,N_648);
nor U1157 (N_1157,In_438,In_1160);
nor U1158 (N_1158,In_51,In_1071);
nand U1159 (N_1159,N_293,In_1432);
xnor U1160 (N_1160,In_981,N_630);
nor U1161 (N_1161,In_1492,In_881);
xor U1162 (N_1162,N_637,In_1413);
and U1163 (N_1163,N_149,N_301);
nor U1164 (N_1164,N_266,N_303);
nor U1165 (N_1165,N_629,In_728);
or U1166 (N_1166,N_866,N_101);
and U1167 (N_1167,N_873,N_793);
nor U1168 (N_1168,In_1293,In_420);
and U1169 (N_1169,N_889,N_117);
and U1170 (N_1170,N_636,N_535);
nor U1171 (N_1171,N_620,N_308);
xnor U1172 (N_1172,In_1026,In_1118);
xnor U1173 (N_1173,N_855,N_507);
and U1174 (N_1174,N_674,N_190);
and U1175 (N_1175,In_257,N_731);
and U1176 (N_1176,N_52,In_1191);
or U1177 (N_1177,N_471,N_723);
xnor U1178 (N_1178,N_505,In_1405);
nor U1179 (N_1179,In_518,N_623);
nand U1180 (N_1180,N_899,N_370);
xor U1181 (N_1181,N_85,N_839);
and U1182 (N_1182,In_454,N_253);
nand U1183 (N_1183,In_7,N_477);
xnor U1184 (N_1184,In_1214,N_71);
and U1185 (N_1185,N_323,N_728);
or U1186 (N_1186,N_792,In_1075);
nor U1187 (N_1187,In_339,In_1127);
and U1188 (N_1188,N_312,N_503);
and U1189 (N_1189,N_603,In_1088);
or U1190 (N_1190,In_883,N_584);
xor U1191 (N_1191,In_776,N_852);
and U1192 (N_1192,N_870,N_771);
and U1193 (N_1193,N_654,N_733);
xor U1194 (N_1194,In_8,N_887);
and U1195 (N_1195,N_628,N_798);
and U1196 (N_1196,N_667,N_822);
nand U1197 (N_1197,N_876,N_331);
nor U1198 (N_1198,N_753,N_670);
or U1199 (N_1199,N_849,N_823);
xnor U1200 (N_1200,N_994,N_1078);
or U1201 (N_1201,N_1133,N_945);
nor U1202 (N_1202,N_912,N_1135);
nand U1203 (N_1203,N_1000,N_900);
nor U1204 (N_1204,N_1087,N_1083);
and U1205 (N_1205,N_1187,N_933);
xor U1206 (N_1206,N_990,N_1104);
and U1207 (N_1207,N_902,N_975);
nand U1208 (N_1208,N_1139,N_1075);
xnor U1209 (N_1209,N_1151,N_949);
xor U1210 (N_1210,N_937,N_928);
and U1211 (N_1211,N_1026,N_1108);
and U1212 (N_1212,N_986,N_977);
xnor U1213 (N_1213,N_1048,N_991);
and U1214 (N_1214,N_954,N_1006);
xor U1215 (N_1215,N_1084,N_913);
nor U1216 (N_1216,N_1118,N_988);
nand U1217 (N_1217,N_1145,N_1093);
xor U1218 (N_1218,N_1132,N_976);
nand U1219 (N_1219,N_970,N_1022);
nor U1220 (N_1220,N_1057,N_1003);
nor U1221 (N_1221,N_916,N_1122);
nand U1222 (N_1222,N_1036,N_1111);
xor U1223 (N_1223,N_1046,N_1090);
nand U1224 (N_1224,N_1156,N_917);
xor U1225 (N_1225,N_1007,N_944);
or U1226 (N_1226,N_1146,N_974);
and U1227 (N_1227,N_972,N_1134);
and U1228 (N_1228,N_1159,N_968);
or U1229 (N_1229,N_1021,N_1189);
nor U1230 (N_1230,N_1106,N_1171);
xnor U1231 (N_1231,N_1193,N_1163);
or U1232 (N_1232,N_1054,N_1028);
and U1233 (N_1233,N_1141,N_1005);
and U1234 (N_1234,N_1095,N_1085);
xnor U1235 (N_1235,N_1168,N_1025);
xnor U1236 (N_1236,N_1130,N_1154);
or U1237 (N_1237,N_983,N_1155);
or U1238 (N_1238,N_1060,N_907);
or U1239 (N_1239,N_966,N_1181);
xnor U1240 (N_1240,N_936,N_1113);
nand U1241 (N_1241,N_1004,N_1055);
xnor U1242 (N_1242,N_980,N_1016);
nor U1243 (N_1243,N_919,N_1024);
and U1244 (N_1244,N_958,N_1065);
nand U1245 (N_1245,N_1010,N_962);
nor U1246 (N_1246,N_973,N_940);
nor U1247 (N_1247,N_1053,N_1008);
nand U1248 (N_1248,N_1039,N_1009);
or U1249 (N_1249,N_1119,N_1032);
xor U1250 (N_1250,N_1176,N_1161);
xnor U1251 (N_1251,N_1081,N_1012);
or U1252 (N_1252,N_1038,N_1027);
nor U1253 (N_1253,N_901,N_1037);
nand U1254 (N_1254,N_947,N_952);
nand U1255 (N_1255,N_946,N_943);
xor U1256 (N_1256,N_1011,N_1063);
xnor U1257 (N_1257,N_1002,N_1014);
nor U1258 (N_1258,N_984,N_1018);
nand U1259 (N_1259,N_1077,N_982);
and U1260 (N_1260,N_1061,N_938);
nor U1261 (N_1261,N_1047,N_992);
or U1262 (N_1262,N_1058,N_1126);
nand U1263 (N_1263,N_1033,N_1042);
xor U1264 (N_1264,N_1149,N_1082);
or U1265 (N_1265,N_1115,N_960);
and U1266 (N_1266,N_1172,N_1192);
xnor U1267 (N_1267,N_1147,N_911);
xnor U1268 (N_1268,N_926,N_905);
or U1269 (N_1269,N_1191,N_1158);
nor U1270 (N_1270,N_1092,N_1101);
or U1271 (N_1271,N_998,N_1109);
nand U1272 (N_1272,N_932,N_1001);
xnor U1273 (N_1273,N_922,N_1040);
nor U1274 (N_1274,N_1100,N_1180);
or U1275 (N_1275,N_1067,N_921);
or U1276 (N_1276,N_1050,N_1013);
or U1277 (N_1277,N_1088,N_1170);
nor U1278 (N_1278,N_1105,N_964);
nor U1279 (N_1279,N_1031,N_1079);
nor U1280 (N_1280,N_1175,N_1023);
and U1281 (N_1281,N_1103,N_1052);
nand U1282 (N_1282,N_959,N_1188);
and U1283 (N_1283,N_1064,N_1177);
and U1284 (N_1284,N_1072,N_1157);
and U1285 (N_1285,N_923,N_903);
or U1286 (N_1286,N_1080,N_1173);
nand U1287 (N_1287,N_929,N_1029);
and U1288 (N_1288,N_953,N_978);
xor U1289 (N_1289,N_935,N_1062);
xor U1290 (N_1290,N_1128,N_1096);
nand U1291 (N_1291,N_908,N_930);
nor U1292 (N_1292,N_1099,N_1110);
nand U1293 (N_1293,N_934,N_941);
nor U1294 (N_1294,N_1107,N_1034);
nor U1295 (N_1295,N_1117,N_927);
nand U1296 (N_1296,N_1166,N_1068);
nor U1297 (N_1297,N_1169,N_963);
and U1298 (N_1298,N_920,N_1094);
xnor U1299 (N_1299,N_1121,N_931);
and U1300 (N_1300,N_1059,N_1199);
and U1301 (N_1301,N_1086,N_997);
nor U1302 (N_1302,N_1020,N_1041);
nand U1303 (N_1303,N_925,N_914);
nand U1304 (N_1304,N_1196,N_939);
nor U1305 (N_1305,N_1116,N_1138);
xnor U1306 (N_1306,N_1198,N_1136);
and U1307 (N_1307,N_996,N_942);
nor U1308 (N_1308,N_1150,N_1164);
or U1309 (N_1309,N_1194,N_1183);
or U1310 (N_1310,N_987,N_1162);
xnor U1311 (N_1311,N_1112,N_961);
xnor U1312 (N_1312,N_1035,N_1049);
xnor U1313 (N_1313,N_1127,N_999);
or U1314 (N_1314,N_967,N_1070);
and U1315 (N_1315,N_915,N_1017);
and U1316 (N_1316,N_1153,N_1066);
xnor U1317 (N_1317,N_1144,N_1179);
or U1318 (N_1318,N_1167,N_1131);
and U1319 (N_1319,N_1069,N_1097);
or U1320 (N_1320,N_981,N_1184);
nand U1321 (N_1321,N_1185,N_1152);
or U1322 (N_1322,N_1030,N_969);
and U1323 (N_1323,N_1073,N_957);
nand U1324 (N_1324,N_1015,N_985);
or U1325 (N_1325,N_909,N_956);
xor U1326 (N_1326,N_1120,N_1186);
xor U1327 (N_1327,N_1165,N_951);
xnor U1328 (N_1328,N_1195,N_1190);
or U1329 (N_1329,N_1044,N_1124);
or U1330 (N_1330,N_918,N_995);
nor U1331 (N_1331,N_1051,N_1074);
and U1332 (N_1332,N_1043,N_1178);
and U1333 (N_1333,N_906,N_1148);
nor U1334 (N_1334,N_1129,N_1140);
nor U1335 (N_1335,N_1102,N_1019);
and U1336 (N_1336,N_1182,N_910);
nand U1337 (N_1337,N_950,N_1091);
and U1338 (N_1338,N_971,N_948);
xor U1339 (N_1339,N_955,N_989);
nor U1340 (N_1340,N_1076,N_1056);
xor U1341 (N_1341,N_924,N_1137);
and U1342 (N_1342,N_1089,N_1045);
and U1343 (N_1343,N_1142,N_1143);
xor U1344 (N_1344,N_1123,N_1098);
nor U1345 (N_1345,N_965,N_1125);
nand U1346 (N_1346,N_1197,N_979);
and U1347 (N_1347,N_993,N_1114);
nor U1348 (N_1348,N_1160,N_1071);
xnor U1349 (N_1349,N_904,N_1174);
and U1350 (N_1350,N_1118,N_1078);
and U1351 (N_1351,N_919,N_1143);
and U1352 (N_1352,N_1072,N_1143);
and U1353 (N_1353,N_1006,N_1174);
nor U1354 (N_1354,N_1124,N_1018);
or U1355 (N_1355,N_1196,N_1171);
and U1356 (N_1356,N_1144,N_1098);
xor U1357 (N_1357,N_1179,N_1006);
xnor U1358 (N_1358,N_932,N_904);
xnor U1359 (N_1359,N_1084,N_901);
nand U1360 (N_1360,N_995,N_1135);
xor U1361 (N_1361,N_1044,N_1012);
xor U1362 (N_1362,N_1043,N_1144);
and U1363 (N_1363,N_947,N_924);
or U1364 (N_1364,N_1103,N_1005);
and U1365 (N_1365,N_1113,N_1040);
xnor U1366 (N_1366,N_1175,N_992);
nand U1367 (N_1367,N_1155,N_1010);
and U1368 (N_1368,N_1066,N_1046);
nor U1369 (N_1369,N_1163,N_1140);
xnor U1370 (N_1370,N_913,N_1082);
or U1371 (N_1371,N_927,N_1005);
and U1372 (N_1372,N_1137,N_1054);
nand U1373 (N_1373,N_1010,N_924);
nor U1374 (N_1374,N_984,N_1179);
nor U1375 (N_1375,N_1199,N_1060);
nand U1376 (N_1376,N_1127,N_983);
nand U1377 (N_1377,N_986,N_968);
and U1378 (N_1378,N_1180,N_902);
nor U1379 (N_1379,N_957,N_971);
and U1380 (N_1380,N_944,N_1038);
or U1381 (N_1381,N_983,N_1088);
nor U1382 (N_1382,N_911,N_902);
nand U1383 (N_1383,N_1039,N_914);
or U1384 (N_1384,N_910,N_1083);
nor U1385 (N_1385,N_1024,N_1066);
or U1386 (N_1386,N_976,N_1037);
nand U1387 (N_1387,N_1098,N_1091);
and U1388 (N_1388,N_1039,N_1049);
and U1389 (N_1389,N_1192,N_1057);
nor U1390 (N_1390,N_950,N_912);
nor U1391 (N_1391,N_1047,N_1139);
and U1392 (N_1392,N_974,N_1113);
nand U1393 (N_1393,N_1158,N_1184);
nand U1394 (N_1394,N_1043,N_1097);
nand U1395 (N_1395,N_1162,N_1170);
nor U1396 (N_1396,N_1073,N_1020);
nor U1397 (N_1397,N_927,N_922);
nand U1398 (N_1398,N_981,N_1019);
and U1399 (N_1399,N_903,N_1095);
and U1400 (N_1400,N_916,N_1007);
or U1401 (N_1401,N_1067,N_975);
nor U1402 (N_1402,N_927,N_949);
or U1403 (N_1403,N_1027,N_1199);
and U1404 (N_1404,N_1093,N_1142);
xor U1405 (N_1405,N_1160,N_907);
or U1406 (N_1406,N_1092,N_1033);
and U1407 (N_1407,N_954,N_970);
or U1408 (N_1408,N_987,N_1141);
xnor U1409 (N_1409,N_1031,N_1006);
xor U1410 (N_1410,N_1054,N_1039);
or U1411 (N_1411,N_958,N_1147);
xnor U1412 (N_1412,N_1191,N_1096);
nor U1413 (N_1413,N_1050,N_972);
nand U1414 (N_1414,N_1027,N_1085);
nand U1415 (N_1415,N_1119,N_1115);
xnor U1416 (N_1416,N_928,N_1048);
xnor U1417 (N_1417,N_943,N_1199);
xor U1418 (N_1418,N_961,N_1139);
nor U1419 (N_1419,N_1162,N_1153);
xor U1420 (N_1420,N_1078,N_970);
nand U1421 (N_1421,N_1176,N_934);
and U1422 (N_1422,N_1192,N_1014);
and U1423 (N_1423,N_1005,N_1173);
or U1424 (N_1424,N_1177,N_1153);
or U1425 (N_1425,N_909,N_1012);
nand U1426 (N_1426,N_911,N_1167);
or U1427 (N_1427,N_1096,N_1087);
nand U1428 (N_1428,N_1053,N_1046);
or U1429 (N_1429,N_922,N_949);
xnor U1430 (N_1430,N_1106,N_994);
xnor U1431 (N_1431,N_1013,N_935);
nor U1432 (N_1432,N_1092,N_1079);
nor U1433 (N_1433,N_1118,N_1063);
and U1434 (N_1434,N_1182,N_989);
and U1435 (N_1435,N_1069,N_916);
xor U1436 (N_1436,N_1182,N_1185);
nor U1437 (N_1437,N_932,N_1023);
xor U1438 (N_1438,N_1132,N_960);
or U1439 (N_1439,N_1087,N_983);
nand U1440 (N_1440,N_1044,N_1079);
and U1441 (N_1441,N_1077,N_1016);
nand U1442 (N_1442,N_959,N_1131);
nor U1443 (N_1443,N_1021,N_1079);
and U1444 (N_1444,N_961,N_1169);
or U1445 (N_1445,N_1000,N_980);
nor U1446 (N_1446,N_965,N_1032);
or U1447 (N_1447,N_1119,N_1012);
xnor U1448 (N_1448,N_1047,N_1049);
xor U1449 (N_1449,N_1018,N_1121);
nand U1450 (N_1450,N_1093,N_933);
xnor U1451 (N_1451,N_1151,N_929);
xnor U1452 (N_1452,N_1096,N_972);
and U1453 (N_1453,N_1139,N_1101);
xor U1454 (N_1454,N_1150,N_1156);
and U1455 (N_1455,N_1033,N_1044);
xnor U1456 (N_1456,N_1165,N_1038);
or U1457 (N_1457,N_1087,N_1011);
nand U1458 (N_1458,N_935,N_1098);
xor U1459 (N_1459,N_1161,N_935);
or U1460 (N_1460,N_1006,N_914);
and U1461 (N_1461,N_1020,N_1087);
nand U1462 (N_1462,N_1106,N_943);
or U1463 (N_1463,N_1182,N_1021);
xor U1464 (N_1464,N_912,N_993);
and U1465 (N_1465,N_1015,N_1137);
nand U1466 (N_1466,N_925,N_1156);
nand U1467 (N_1467,N_1043,N_1090);
xnor U1468 (N_1468,N_1078,N_1068);
nand U1469 (N_1469,N_1051,N_1014);
and U1470 (N_1470,N_1039,N_962);
xnor U1471 (N_1471,N_1197,N_935);
xor U1472 (N_1472,N_929,N_1039);
and U1473 (N_1473,N_975,N_1041);
xnor U1474 (N_1474,N_1122,N_1048);
and U1475 (N_1475,N_1027,N_1164);
nand U1476 (N_1476,N_1181,N_928);
or U1477 (N_1477,N_1116,N_900);
and U1478 (N_1478,N_914,N_1049);
or U1479 (N_1479,N_1086,N_1170);
nand U1480 (N_1480,N_1097,N_963);
nand U1481 (N_1481,N_965,N_1195);
or U1482 (N_1482,N_1063,N_1065);
or U1483 (N_1483,N_1026,N_1037);
nor U1484 (N_1484,N_1150,N_1152);
nor U1485 (N_1485,N_934,N_1197);
nor U1486 (N_1486,N_926,N_1153);
xor U1487 (N_1487,N_945,N_1050);
xor U1488 (N_1488,N_1110,N_1109);
nand U1489 (N_1489,N_1112,N_1153);
or U1490 (N_1490,N_1056,N_1093);
or U1491 (N_1491,N_1081,N_958);
nand U1492 (N_1492,N_1080,N_1087);
nor U1493 (N_1493,N_940,N_1020);
xor U1494 (N_1494,N_1127,N_1028);
and U1495 (N_1495,N_1193,N_1097);
and U1496 (N_1496,N_1023,N_1188);
and U1497 (N_1497,N_927,N_1049);
xnor U1498 (N_1498,N_994,N_957);
nor U1499 (N_1499,N_1091,N_1008);
nor U1500 (N_1500,N_1473,N_1336);
xnor U1501 (N_1501,N_1449,N_1474);
and U1502 (N_1502,N_1226,N_1382);
nor U1503 (N_1503,N_1267,N_1229);
xor U1504 (N_1504,N_1466,N_1215);
and U1505 (N_1505,N_1470,N_1419);
nor U1506 (N_1506,N_1270,N_1365);
nand U1507 (N_1507,N_1445,N_1414);
nor U1508 (N_1508,N_1420,N_1494);
xnor U1509 (N_1509,N_1206,N_1236);
xor U1510 (N_1510,N_1303,N_1252);
nor U1511 (N_1511,N_1332,N_1313);
nor U1512 (N_1512,N_1289,N_1264);
nor U1513 (N_1513,N_1245,N_1388);
and U1514 (N_1514,N_1385,N_1295);
xor U1515 (N_1515,N_1492,N_1342);
and U1516 (N_1516,N_1395,N_1352);
xnor U1517 (N_1517,N_1323,N_1450);
and U1518 (N_1518,N_1446,N_1468);
nor U1519 (N_1519,N_1374,N_1490);
nor U1520 (N_1520,N_1242,N_1339);
nor U1521 (N_1521,N_1308,N_1348);
xnor U1522 (N_1522,N_1321,N_1418);
or U1523 (N_1523,N_1408,N_1256);
xnor U1524 (N_1524,N_1328,N_1320);
nor U1525 (N_1525,N_1377,N_1478);
nand U1526 (N_1526,N_1220,N_1265);
or U1527 (N_1527,N_1269,N_1307);
or U1528 (N_1528,N_1412,N_1326);
nor U1529 (N_1529,N_1370,N_1378);
xor U1530 (N_1530,N_1399,N_1330);
and U1531 (N_1531,N_1393,N_1467);
nor U1532 (N_1532,N_1260,N_1356);
nand U1533 (N_1533,N_1325,N_1223);
or U1534 (N_1534,N_1361,N_1274);
or U1535 (N_1535,N_1431,N_1235);
nor U1536 (N_1536,N_1425,N_1331);
nor U1537 (N_1537,N_1358,N_1479);
xor U1538 (N_1538,N_1278,N_1271);
and U1539 (N_1539,N_1394,N_1211);
xnor U1540 (N_1540,N_1246,N_1448);
nand U1541 (N_1541,N_1230,N_1324);
nand U1542 (N_1542,N_1241,N_1337);
xnor U1543 (N_1543,N_1417,N_1345);
nand U1544 (N_1544,N_1469,N_1403);
and U1545 (N_1545,N_1222,N_1231);
nor U1546 (N_1546,N_1369,N_1463);
xor U1547 (N_1547,N_1224,N_1259);
and U1548 (N_1548,N_1362,N_1288);
and U1549 (N_1549,N_1329,N_1316);
nor U1550 (N_1550,N_1272,N_1327);
nor U1551 (N_1551,N_1407,N_1373);
xnor U1552 (N_1552,N_1305,N_1263);
nor U1553 (N_1553,N_1472,N_1453);
nor U1554 (N_1554,N_1451,N_1411);
xor U1555 (N_1555,N_1281,N_1301);
nor U1556 (N_1556,N_1415,N_1386);
or U1557 (N_1557,N_1335,N_1484);
xor U1558 (N_1558,N_1338,N_1317);
and U1559 (N_1559,N_1239,N_1475);
xor U1560 (N_1560,N_1404,N_1402);
and U1561 (N_1561,N_1423,N_1319);
or U1562 (N_1562,N_1253,N_1396);
xnor U1563 (N_1563,N_1461,N_1353);
nor U1564 (N_1564,N_1243,N_1410);
nand U1565 (N_1565,N_1218,N_1481);
and U1566 (N_1566,N_1294,N_1392);
or U1567 (N_1567,N_1304,N_1432);
and U1568 (N_1568,N_1233,N_1428);
nor U1569 (N_1569,N_1217,N_1255);
xnor U1570 (N_1570,N_1207,N_1401);
and U1571 (N_1571,N_1314,N_1208);
nor U1572 (N_1572,N_1292,N_1375);
nand U1573 (N_1573,N_1216,N_1363);
and U1574 (N_1574,N_1455,N_1427);
xnor U1575 (N_1575,N_1257,N_1486);
nand U1576 (N_1576,N_1234,N_1202);
or U1577 (N_1577,N_1340,N_1387);
and U1578 (N_1578,N_1477,N_1483);
xnor U1579 (N_1579,N_1232,N_1351);
and U1580 (N_1580,N_1435,N_1444);
xor U1581 (N_1581,N_1489,N_1371);
nand U1582 (N_1582,N_1341,N_1498);
xnor U1583 (N_1583,N_1383,N_1300);
nand U1584 (N_1584,N_1280,N_1282);
nor U1585 (N_1585,N_1344,N_1276);
or U1586 (N_1586,N_1397,N_1460);
nand U1587 (N_1587,N_1452,N_1426);
xor U1588 (N_1588,N_1203,N_1249);
nor U1589 (N_1589,N_1476,N_1464);
nor U1590 (N_1590,N_1380,N_1268);
nand U1591 (N_1591,N_1422,N_1279);
nor U1592 (N_1592,N_1251,N_1299);
or U1593 (N_1593,N_1424,N_1346);
and U1594 (N_1594,N_1438,N_1277);
and U1595 (N_1595,N_1248,N_1379);
nor U1596 (N_1596,N_1360,N_1409);
nand U1597 (N_1597,N_1493,N_1482);
xnor U1598 (N_1598,N_1350,N_1290);
or U1599 (N_1599,N_1298,N_1497);
or U1600 (N_1600,N_1244,N_1405);
nor U1601 (N_1601,N_1254,N_1293);
nand U1602 (N_1602,N_1368,N_1367);
xnor U1603 (N_1603,N_1436,N_1390);
or U1604 (N_1604,N_1496,N_1357);
nor U1605 (N_1605,N_1439,N_1389);
nor U1606 (N_1606,N_1366,N_1430);
or U1607 (N_1607,N_1355,N_1413);
or U1608 (N_1608,N_1487,N_1406);
and U1609 (N_1609,N_1376,N_1364);
or U1610 (N_1610,N_1441,N_1462);
nor U1611 (N_1611,N_1354,N_1247);
xor U1612 (N_1612,N_1238,N_1212);
and U1613 (N_1613,N_1447,N_1310);
or U1614 (N_1614,N_1359,N_1287);
or U1615 (N_1615,N_1297,N_1458);
nand U1616 (N_1616,N_1491,N_1398);
nor U1617 (N_1617,N_1454,N_1286);
nor U1618 (N_1618,N_1209,N_1210);
nor U1619 (N_1619,N_1201,N_1349);
or U1620 (N_1620,N_1381,N_1457);
or U1621 (N_1621,N_1456,N_1266);
or U1622 (N_1622,N_1291,N_1429);
and U1623 (N_1623,N_1302,N_1400);
nor U1624 (N_1624,N_1273,N_1347);
nor U1625 (N_1625,N_1205,N_1221);
and U1626 (N_1626,N_1284,N_1285);
xor U1627 (N_1627,N_1333,N_1275);
or U1628 (N_1628,N_1204,N_1309);
nor U1629 (N_1629,N_1237,N_1322);
nand U1630 (N_1630,N_1262,N_1214);
or U1631 (N_1631,N_1480,N_1437);
and U1632 (N_1632,N_1440,N_1485);
and U1633 (N_1633,N_1343,N_1306);
xnor U1634 (N_1634,N_1495,N_1213);
and U1635 (N_1635,N_1372,N_1283);
nand U1636 (N_1636,N_1488,N_1384);
nor U1637 (N_1637,N_1296,N_1228);
xor U1638 (N_1638,N_1318,N_1311);
nand U1639 (N_1639,N_1240,N_1219);
xor U1640 (N_1640,N_1433,N_1465);
and U1641 (N_1641,N_1200,N_1391);
nor U1642 (N_1642,N_1442,N_1434);
or U1643 (N_1643,N_1225,N_1315);
nand U1644 (N_1644,N_1261,N_1421);
nor U1645 (N_1645,N_1459,N_1334);
xnor U1646 (N_1646,N_1258,N_1471);
and U1647 (N_1647,N_1227,N_1443);
nand U1648 (N_1648,N_1250,N_1416);
nor U1649 (N_1649,N_1312,N_1499);
xnor U1650 (N_1650,N_1368,N_1493);
xor U1651 (N_1651,N_1349,N_1351);
xor U1652 (N_1652,N_1212,N_1352);
nor U1653 (N_1653,N_1369,N_1238);
and U1654 (N_1654,N_1383,N_1207);
or U1655 (N_1655,N_1215,N_1287);
nor U1656 (N_1656,N_1207,N_1310);
or U1657 (N_1657,N_1412,N_1380);
nor U1658 (N_1658,N_1330,N_1335);
and U1659 (N_1659,N_1398,N_1479);
nand U1660 (N_1660,N_1443,N_1268);
nand U1661 (N_1661,N_1472,N_1351);
and U1662 (N_1662,N_1417,N_1421);
nor U1663 (N_1663,N_1276,N_1264);
and U1664 (N_1664,N_1346,N_1473);
nor U1665 (N_1665,N_1229,N_1257);
xor U1666 (N_1666,N_1495,N_1276);
or U1667 (N_1667,N_1410,N_1452);
nor U1668 (N_1668,N_1479,N_1415);
or U1669 (N_1669,N_1395,N_1326);
nand U1670 (N_1670,N_1261,N_1312);
nor U1671 (N_1671,N_1416,N_1265);
nor U1672 (N_1672,N_1398,N_1274);
nor U1673 (N_1673,N_1232,N_1250);
nand U1674 (N_1674,N_1461,N_1239);
or U1675 (N_1675,N_1294,N_1376);
nor U1676 (N_1676,N_1217,N_1448);
and U1677 (N_1677,N_1209,N_1331);
nand U1678 (N_1678,N_1308,N_1406);
xnor U1679 (N_1679,N_1391,N_1271);
nor U1680 (N_1680,N_1376,N_1241);
or U1681 (N_1681,N_1389,N_1374);
xor U1682 (N_1682,N_1294,N_1363);
nor U1683 (N_1683,N_1348,N_1396);
nand U1684 (N_1684,N_1458,N_1457);
xnor U1685 (N_1685,N_1352,N_1260);
and U1686 (N_1686,N_1262,N_1373);
and U1687 (N_1687,N_1373,N_1221);
nand U1688 (N_1688,N_1344,N_1363);
or U1689 (N_1689,N_1352,N_1232);
xnor U1690 (N_1690,N_1461,N_1352);
nor U1691 (N_1691,N_1352,N_1226);
nor U1692 (N_1692,N_1292,N_1406);
and U1693 (N_1693,N_1200,N_1341);
nand U1694 (N_1694,N_1342,N_1298);
and U1695 (N_1695,N_1455,N_1379);
or U1696 (N_1696,N_1317,N_1347);
and U1697 (N_1697,N_1347,N_1460);
nand U1698 (N_1698,N_1337,N_1249);
nand U1699 (N_1699,N_1231,N_1207);
xor U1700 (N_1700,N_1224,N_1234);
and U1701 (N_1701,N_1333,N_1395);
xor U1702 (N_1702,N_1447,N_1313);
nand U1703 (N_1703,N_1385,N_1204);
nand U1704 (N_1704,N_1450,N_1241);
nand U1705 (N_1705,N_1494,N_1470);
or U1706 (N_1706,N_1362,N_1348);
xnor U1707 (N_1707,N_1371,N_1406);
and U1708 (N_1708,N_1410,N_1311);
or U1709 (N_1709,N_1392,N_1255);
nor U1710 (N_1710,N_1370,N_1433);
nor U1711 (N_1711,N_1226,N_1246);
and U1712 (N_1712,N_1398,N_1350);
nor U1713 (N_1713,N_1480,N_1376);
or U1714 (N_1714,N_1353,N_1326);
nand U1715 (N_1715,N_1450,N_1398);
or U1716 (N_1716,N_1380,N_1240);
or U1717 (N_1717,N_1212,N_1426);
or U1718 (N_1718,N_1426,N_1381);
or U1719 (N_1719,N_1286,N_1491);
xor U1720 (N_1720,N_1438,N_1468);
xnor U1721 (N_1721,N_1491,N_1281);
xnor U1722 (N_1722,N_1392,N_1243);
or U1723 (N_1723,N_1296,N_1310);
and U1724 (N_1724,N_1386,N_1227);
nor U1725 (N_1725,N_1452,N_1337);
nand U1726 (N_1726,N_1361,N_1317);
or U1727 (N_1727,N_1277,N_1221);
and U1728 (N_1728,N_1425,N_1236);
nor U1729 (N_1729,N_1319,N_1239);
nand U1730 (N_1730,N_1316,N_1330);
xor U1731 (N_1731,N_1261,N_1386);
nand U1732 (N_1732,N_1363,N_1210);
or U1733 (N_1733,N_1277,N_1385);
nand U1734 (N_1734,N_1390,N_1293);
or U1735 (N_1735,N_1211,N_1262);
or U1736 (N_1736,N_1485,N_1397);
or U1737 (N_1737,N_1429,N_1233);
nand U1738 (N_1738,N_1488,N_1226);
nand U1739 (N_1739,N_1279,N_1357);
or U1740 (N_1740,N_1351,N_1306);
xor U1741 (N_1741,N_1468,N_1302);
xor U1742 (N_1742,N_1249,N_1453);
and U1743 (N_1743,N_1463,N_1394);
and U1744 (N_1744,N_1380,N_1403);
and U1745 (N_1745,N_1393,N_1332);
or U1746 (N_1746,N_1347,N_1386);
nand U1747 (N_1747,N_1499,N_1482);
and U1748 (N_1748,N_1490,N_1289);
or U1749 (N_1749,N_1365,N_1460);
xnor U1750 (N_1750,N_1363,N_1237);
nor U1751 (N_1751,N_1212,N_1378);
nor U1752 (N_1752,N_1372,N_1441);
nand U1753 (N_1753,N_1324,N_1413);
nor U1754 (N_1754,N_1222,N_1370);
and U1755 (N_1755,N_1456,N_1358);
nor U1756 (N_1756,N_1474,N_1470);
nand U1757 (N_1757,N_1361,N_1212);
nand U1758 (N_1758,N_1428,N_1200);
and U1759 (N_1759,N_1380,N_1451);
nor U1760 (N_1760,N_1340,N_1353);
xor U1761 (N_1761,N_1323,N_1365);
and U1762 (N_1762,N_1285,N_1313);
nand U1763 (N_1763,N_1417,N_1423);
and U1764 (N_1764,N_1433,N_1476);
xnor U1765 (N_1765,N_1315,N_1419);
and U1766 (N_1766,N_1390,N_1292);
nand U1767 (N_1767,N_1424,N_1471);
nand U1768 (N_1768,N_1473,N_1451);
xnor U1769 (N_1769,N_1499,N_1259);
or U1770 (N_1770,N_1323,N_1215);
and U1771 (N_1771,N_1275,N_1473);
xor U1772 (N_1772,N_1216,N_1449);
or U1773 (N_1773,N_1356,N_1298);
or U1774 (N_1774,N_1436,N_1273);
nand U1775 (N_1775,N_1320,N_1307);
nand U1776 (N_1776,N_1471,N_1425);
or U1777 (N_1777,N_1356,N_1237);
xor U1778 (N_1778,N_1230,N_1313);
nor U1779 (N_1779,N_1328,N_1445);
nor U1780 (N_1780,N_1335,N_1200);
nor U1781 (N_1781,N_1433,N_1337);
or U1782 (N_1782,N_1370,N_1495);
or U1783 (N_1783,N_1251,N_1244);
nor U1784 (N_1784,N_1200,N_1310);
nand U1785 (N_1785,N_1345,N_1207);
or U1786 (N_1786,N_1244,N_1230);
nand U1787 (N_1787,N_1228,N_1363);
nor U1788 (N_1788,N_1437,N_1300);
or U1789 (N_1789,N_1303,N_1328);
xor U1790 (N_1790,N_1458,N_1322);
or U1791 (N_1791,N_1471,N_1357);
nand U1792 (N_1792,N_1357,N_1266);
or U1793 (N_1793,N_1330,N_1291);
xor U1794 (N_1794,N_1387,N_1480);
nand U1795 (N_1795,N_1271,N_1485);
and U1796 (N_1796,N_1413,N_1314);
nor U1797 (N_1797,N_1273,N_1462);
nor U1798 (N_1798,N_1461,N_1483);
and U1799 (N_1799,N_1277,N_1283);
nor U1800 (N_1800,N_1513,N_1653);
and U1801 (N_1801,N_1688,N_1736);
and U1802 (N_1802,N_1745,N_1743);
and U1803 (N_1803,N_1531,N_1590);
xor U1804 (N_1804,N_1710,N_1526);
xor U1805 (N_1805,N_1703,N_1640);
nand U1806 (N_1806,N_1606,N_1671);
nand U1807 (N_1807,N_1681,N_1524);
xor U1808 (N_1808,N_1641,N_1540);
and U1809 (N_1809,N_1503,N_1594);
and U1810 (N_1810,N_1670,N_1793);
xnor U1811 (N_1811,N_1648,N_1636);
nand U1812 (N_1812,N_1677,N_1795);
or U1813 (N_1813,N_1601,N_1785);
or U1814 (N_1814,N_1551,N_1610);
or U1815 (N_1815,N_1635,N_1578);
or U1816 (N_1816,N_1798,N_1669);
xor U1817 (N_1817,N_1779,N_1598);
xor U1818 (N_1818,N_1783,N_1738);
or U1819 (N_1819,N_1548,N_1697);
xnor U1820 (N_1820,N_1559,N_1542);
xor U1821 (N_1821,N_1532,N_1799);
or U1822 (N_1822,N_1607,N_1692);
and U1823 (N_1823,N_1569,N_1570);
and U1824 (N_1824,N_1682,N_1660);
xor U1825 (N_1825,N_1603,N_1505);
nor U1826 (N_1826,N_1634,N_1719);
xor U1827 (N_1827,N_1666,N_1612);
and U1828 (N_1828,N_1756,N_1538);
nor U1829 (N_1829,N_1528,N_1623);
and U1830 (N_1830,N_1575,N_1584);
nand U1831 (N_1831,N_1545,N_1797);
nand U1832 (N_1832,N_1512,N_1775);
and U1833 (N_1833,N_1737,N_1760);
nand U1834 (N_1834,N_1502,N_1546);
and U1835 (N_1835,N_1701,N_1791);
xor U1836 (N_1836,N_1672,N_1732);
nand U1837 (N_1837,N_1630,N_1698);
xor U1838 (N_1838,N_1611,N_1708);
or U1839 (N_1839,N_1553,N_1766);
nor U1840 (N_1840,N_1683,N_1566);
and U1841 (N_1841,N_1789,N_1758);
nor U1842 (N_1842,N_1508,N_1574);
or U1843 (N_1843,N_1723,N_1582);
nor U1844 (N_1844,N_1744,N_1721);
nand U1845 (N_1845,N_1638,N_1767);
xnor U1846 (N_1846,N_1739,N_1534);
nor U1847 (N_1847,N_1725,N_1765);
and U1848 (N_1848,N_1763,N_1517);
nand U1849 (N_1849,N_1749,N_1773);
nand U1850 (N_1850,N_1622,N_1509);
nand U1851 (N_1851,N_1750,N_1595);
or U1852 (N_1852,N_1714,N_1709);
nand U1853 (N_1853,N_1627,N_1693);
and U1854 (N_1854,N_1695,N_1533);
nor U1855 (N_1855,N_1746,N_1652);
nand U1856 (N_1856,N_1718,N_1620);
nand U1857 (N_1857,N_1777,N_1615);
xnor U1858 (N_1858,N_1572,N_1511);
nand U1859 (N_1859,N_1587,N_1522);
and U1860 (N_1860,N_1729,N_1792);
nor U1861 (N_1861,N_1631,N_1514);
or U1862 (N_1862,N_1519,N_1597);
and U1863 (N_1863,N_1618,N_1573);
or U1864 (N_1864,N_1702,N_1550);
nand U1865 (N_1865,N_1751,N_1501);
or U1866 (N_1866,N_1796,N_1716);
xnor U1867 (N_1867,N_1543,N_1518);
nor U1868 (N_1868,N_1699,N_1794);
and U1869 (N_1869,N_1654,N_1642);
and U1870 (N_1870,N_1711,N_1764);
nor U1871 (N_1871,N_1571,N_1656);
and U1872 (N_1872,N_1537,N_1753);
nand U1873 (N_1873,N_1724,N_1759);
or U1874 (N_1874,N_1678,N_1625);
or U1875 (N_1875,N_1771,N_1772);
and U1876 (N_1876,N_1757,N_1655);
or U1877 (N_1877,N_1673,N_1589);
and U1878 (N_1878,N_1609,N_1722);
or U1879 (N_1879,N_1782,N_1593);
and U1880 (N_1880,N_1646,N_1628);
and U1881 (N_1881,N_1617,N_1561);
xor U1882 (N_1882,N_1696,N_1774);
or U1883 (N_1883,N_1727,N_1668);
nand U1884 (N_1884,N_1536,N_1544);
xor U1885 (N_1885,N_1715,N_1780);
xnor U1886 (N_1886,N_1563,N_1592);
nor U1887 (N_1887,N_1784,N_1755);
nor U1888 (N_1888,N_1776,N_1700);
nor U1889 (N_1889,N_1781,N_1658);
nor U1890 (N_1890,N_1735,N_1730);
xnor U1891 (N_1891,N_1649,N_1748);
nor U1892 (N_1892,N_1579,N_1787);
nand U1893 (N_1893,N_1619,N_1676);
xnor U1894 (N_1894,N_1786,N_1500);
xor U1895 (N_1895,N_1637,N_1687);
xnor U1896 (N_1896,N_1567,N_1564);
and U1897 (N_1897,N_1675,N_1560);
nand U1898 (N_1898,N_1521,N_1539);
nand U1899 (N_1899,N_1565,N_1728);
nand U1900 (N_1900,N_1506,N_1614);
xnor U1901 (N_1901,N_1643,N_1516);
xnor U1902 (N_1902,N_1568,N_1588);
nand U1903 (N_1903,N_1510,N_1562);
or U1904 (N_1904,N_1555,N_1591);
xor U1905 (N_1905,N_1769,N_1768);
and U1906 (N_1906,N_1788,N_1604);
or U1907 (N_1907,N_1661,N_1742);
xnor U1908 (N_1908,N_1527,N_1600);
xor U1909 (N_1909,N_1713,N_1694);
xor U1910 (N_1910,N_1645,N_1651);
or U1911 (N_1911,N_1552,N_1583);
or U1912 (N_1912,N_1667,N_1541);
nand U1913 (N_1913,N_1690,N_1712);
nand U1914 (N_1914,N_1525,N_1685);
nand U1915 (N_1915,N_1686,N_1680);
nand U1916 (N_1916,N_1613,N_1717);
nor U1917 (N_1917,N_1762,N_1639);
nor U1918 (N_1918,N_1657,N_1577);
and U1919 (N_1919,N_1644,N_1535);
nand U1920 (N_1920,N_1608,N_1504);
nor U1921 (N_1921,N_1752,N_1741);
nor U1922 (N_1922,N_1720,N_1679);
and U1923 (N_1923,N_1529,N_1520);
xnor U1924 (N_1924,N_1556,N_1778);
nor U1925 (N_1925,N_1705,N_1733);
nor U1926 (N_1926,N_1707,N_1629);
nor U1927 (N_1927,N_1547,N_1665);
or U1928 (N_1928,N_1616,N_1747);
nand U1929 (N_1929,N_1621,N_1599);
nor U1930 (N_1930,N_1576,N_1706);
xnor U1931 (N_1931,N_1558,N_1659);
nand U1932 (N_1932,N_1596,N_1585);
nor U1933 (N_1933,N_1726,N_1740);
nand U1934 (N_1934,N_1626,N_1754);
nor U1935 (N_1935,N_1530,N_1790);
nand U1936 (N_1936,N_1580,N_1586);
nor U1937 (N_1937,N_1704,N_1650);
and U1938 (N_1938,N_1523,N_1770);
nor U1939 (N_1939,N_1761,N_1674);
xor U1940 (N_1940,N_1647,N_1557);
or U1941 (N_1941,N_1734,N_1684);
xor U1942 (N_1942,N_1691,N_1602);
and U1943 (N_1943,N_1689,N_1664);
or U1944 (N_1944,N_1515,N_1605);
xnor U1945 (N_1945,N_1633,N_1731);
nand U1946 (N_1946,N_1662,N_1507);
and U1947 (N_1947,N_1549,N_1624);
or U1948 (N_1948,N_1554,N_1663);
and U1949 (N_1949,N_1632,N_1581);
nor U1950 (N_1950,N_1587,N_1710);
nand U1951 (N_1951,N_1763,N_1783);
xnor U1952 (N_1952,N_1545,N_1502);
nor U1953 (N_1953,N_1633,N_1715);
and U1954 (N_1954,N_1567,N_1792);
nand U1955 (N_1955,N_1793,N_1679);
nor U1956 (N_1956,N_1778,N_1564);
nand U1957 (N_1957,N_1774,N_1540);
nand U1958 (N_1958,N_1569,N_1723);
nand U1959 (N_1959,N_1554,N_1791);
nor U1960 (N_1960,N_1778,N_1557);
and U1961 (N_1961,N_1532,N_1692);
or U1962 (N_1962,N_1798,N_1548);
nand U1963 (N_1963,N_1591,N_1523);
nand U1964 (N_1964,N_1641,N_1675);
and U1965 (N_1965,N_1756,N_1752);
and U1966 (N_1966,N_1592,N_1775);
and U1967 (N_1967,N_1554,N_1542);
xor U1968 (N_1968,N_1747,N_1690);
and U1969 (N_1969,N_1621,N_1576);
xnor U1970 (N_1970,N_1516,N_1782);
and U1971 (N_1971,N_1629,N_1621);
xor U1972 (N_1972,N_1528,N_1507);
xnor U1973 (N_1973,N_1554,N_1683);
nor U1974 (N_1974,N_1553,N_1515);
or U1975 (N_1975,N_1510,N_1500);
or U1976 (N_1976,N_1627,N_1598);
or U1977 (N_1977,N_1684,N_1526);
nand U1978 (N_1978,N_1786,N_1673);
and U1979 (N_1979,N_1726,N_1758);
or U1980 (N_1980,N_1724,N_1656);
nor U1981 (N_1981,N_1531,N_1634);
and U1982 (N_1982,N_1782,N_1798);
and U1983 (N_1983,N_1762,N_1631);
nor U1984 (N_1984,N_1552,N_1762);
and U1985 (N_1985,N_1794,N_1646);
and U1986 (N_1986,N_1717,N_1523);
or U1987 (N_1987,N_1655,N_1542);
and U1988 (N_1988,N_1640,N_1789);
nand U1989 (N_1989,N_1545,N_1619);
nand U1990 (N_1990,N_1787,N_1567);
or U1991 (N_1991,N_1603,N_1584);
or U1992 (N_1992,N_1523,N_1798);
nand U1993 (N_1993,N_1797,N_1740);
xor U1994 (N_1994,N_1699,N_1670);
nand U1995 (N_1995,N_1627,N_1674);
or U1996 (N_1996,N_1556,N_1666);
nor U1997 (N_1997,N_1608,N_1587);
xor U1998 (N_1998,N_1523,N_1748);
or U1999 (N_1999,N_1678,N_1669);
or U2000 (N_2000,N_1784,N_1523);
nor U2001 (N_2001,N_1541,N_1655);
nand U2002 (N_2002,N_1560,N_1527);
nand U2003 (N_2003,N_1719,N_1534);
or U2004 (N_2004,N_1762,N_1541);
xor U2005 (N_2005,N_1622,N_1753);
or U2006 (N_2006,N_1661,N_1572);
nor U2007 (N_2007,N_1770,N_1533);
or U2008 (N_2008,N_1749,N_1695);
and U2009 (N_2009,N_1524,N_1633);
xnor U2010 (N_2010,N_1651,N_1715);
nor U2011 (N_2011,N_1595,N_1540);
nor U2012 (N_2012,N_1525,N_1535);
nor U2013 (N_2013,N_1754,N_1531);
and U2014 (N_2014,N_1577,N_1512);
xnor U2015 (N_2015,N_1689,N_1526);
xor U2016 (N_2016,N_1523,N_1719);
xnor U2017 (N_2017,N_1668,N_1542);
nor U2018 (N_2018,N_1708,N_1573);
xor U2019 (N_2019,N_1667,N_1649);
nor U2020 (N_2020,N_1761,N_1597);
nand U2021 (N_2021,N_1530,N_1622);
or U2022 (N_2022,N_1592,N_1707);
and U2023 (N_2023,N_1775,N_1694);
or U2024 (N_2024,N_1591,N_1649);
nand U2025 (N_2025,N_1708,N_1736);
nor U2026 (N_2026,N_1512,N_1607);
xor U2027 (N_2027,N_1585,N_1615);
nand U2028 (N_2028,N_1606,N_1611);
nor U2029 (N_2029,N_1791,N_1526);
xor U2030 (N_2030,N_1629,N_1675);
nor U2031 (N_2031,N_1577,N_1658);
and U2032 (N_2032,N_1523,N_1560);
nand U2033 (N_2033,N_1569,N_1653);
nor U2034 (N_2034,N_1721,N_1660);
xnor U2035 (N_2035,N_1721,N_1756);
or U2036 (N_2036,N_1536,N_1669);
nand U2037 (N_2037,N_1586,N_1653);
nand U2038 (N_2038,N_1631,N_1605);
and U2039 (N_2039,N_1707,N_1500);
and U2040 (N_2040,N_1642,N_1502);
or U2041 (N_2041,N_1569,N_1688);
nor U2042 (N_2042,N_1659,N_1717);
or U2043 (N_2043,N_1526,N_1721);
nor U2044 (N_2044,N_1511,N_1641);
xor U2045 (N_2045,N_1550,N_1649);
xor U2046 (N_2046,N_1776,N_1777);
or U2047 (N_2047,N_1729,N_1590);
or U2048 (N_2048,N_1570,N_1651);
nor U2049 (N_2049,N_1510,N_1787);
xnor U2050 (N_2050,N_1515,N_1556);
and U2051 (N_2051,N_1721,N_1705);
and U2052 (N_2052,N_1600,N_1759);
xnor U2053 (N_2053,N_1522,N_1508);
xnor U2054 (N_2054,N_1776,N_1510);
xor U2055 (N_2055,N_1562,N_1670);
and U2056 (N_2056,N_1725,N_1744);
nand U2057 (N_2057,N_1653,N_1576);
nor U2058 (N_2058,N_1745,N_1629);
nand U2059 (N_2059,N_1559,N_1692);
nor U2060 (N_2060,N_1512,N_1699);
and U2061 (N_2061,N_1795,N_1552);
nor U2062 (N_2062,N_1585,N_1645);
and U2063 (N_2063,N_1592,N_1792);
xnor U2064 (N_2064,N_1794,N_1772);
nand U2065 (N_2065,N_1623,N_1765);
xnor U2066 (N_2066,N_1582,N_1526);
nor U2067 (N_2067,N_1539,N_1598);
xnor U2068 (N_2068,N_1512,N_1588);
and U2069 (N_2069,N_1647,N_1511);
xnor U2070 (N_2070,N_1546,N_1683);
and U2071 (N_2071,N_1721,N_1538);
nand U2072 (N_2072,N_1620,N_1534);
nor U2073 (N_2073,N_1653,N_1705);
or U2074 (N_2074,N_1602,N_1616);
nand U2075 (N_2075,N_1527,N_1733);
or U2076 (N_2076,N_1565,N_1572);
nand U2077 (N_2077,N_1783,N_1718);
or U2078 (N_2078,N_1629,N_1588);
or U2079 (N_2079,N_1520,N_1799);
nand U2080 (N_2080,N_1614,N_1749);
xor U2081 (N_2081,N_1659,N_1667);
nor U2082 (N_2082,N_1601,N_1659);
nor U2083 (N_2083,N_1766,N_1598);
nor U2084 (N_2084,N_1731,N_1517);
or U2085 (N_2085,N_1764,N_1695);
xor U2086 (N_2086,N_1745,N_1702);
and U2087 (N_2087,N_1637,N_1612);
xor U2088 (N_2088,N_1591,N_1556);
nor U2089 (N_2089,N_1711,N_1562);
and U2090 (N_2090,N_1572,N_1615);
or U2091 (N_2091,N_1744,N_1637);
nor U2092 (N_2092,N_1574,N_1534);
nand U2093 (N_2093,N_1575,N_1512);
or U2094 (N_2094,N_1653,N_1736);
or U2095 (N_2095,N_1597,N_1567);
nor U2096 (N_2096,N_1684,N_1794);
nor U2097 (N_2097,N_1698,N_1581);
nand U2098 (N_2098,N_1662,N_1575);
and U2099 (N_2099,N_1671,N_1516);
nand U2100 (N_2100,N_2001,N_1844);
or U2101 (N_2101,N_2007,N_2081);
nand U2102 (N_2102,N_1857,N_2017);
nor U2103 (N_2103,N_1838,N_1864);
xor U2104 (N_2104,N_2028,N_2025);
nand U2105 (N_2105,N_1831,N_1980);
and U2106 (N_2106,N_1904,N_2098);
or U2107 (N_2107,N_1893,N_2011);
nand U2108 (N_2108,N_1919,N_1861);
nand U2109 (N_2109,N_1916,N_2002);
nor U2110 (N_2110,N_1821,N_1848);
and U2111 (N_2111,N_2064,N_1906);
nor U2112 (N_2112,N_1932,N_1955);
and U2113 (N_2113,N_1994,N_1886);
xnor U2114 (N_2114,N_2022,N_2016);
and U2115 (N_2115,N_2049,N_1997);
and U2116 (N_2116,N_2031,N_1850);
nor U2117 (N_2117,N_1926,N_2026);
nor U2118 (N_2118,N_1967,N_1824);
and U2119 (N_2119,N_1996,N_2055);
and U2120 (N_2120,N_2008,N_1858);
nand U2121 (N_2121,N_2003,N_1877);
or U2122 (N_2122,N_1975,N_1934);
and U2123 (N_2123,N_1827,N_2018);
nand U2124 (N_2124,N_1900,N_1897);
nand U2125 (N_2125,N_2070,N_1878);
nand U2126 (N_2126,N_1914,N_1887);
xnor U2127 (N_2127,N_2073,N_1960);
xor U2128 (N_2128,N_1944,N_1936);
nand U2129 (N_2129,N_1981,N_2060);
or U2130 (N_2130,N_2024,N_1851);
nand U2131 (N_2131,N_1933,N_1840);
nand U2132 (N_2132,N_1847,N_1825);
or U2133 (N_2133,N_2078,N_1938);
nor U2134 (N_2134,N_1884,N_2051);
nor U2135 (N_2135,N_1963,N_2086);
xnor U2136 (N_2136,N_1855,N_2095);
or U2137 (N_2137,N_2054,N_1950);
nor U2138 (N_2138,N_2039,N_1905);
nor U2139 (N_2139,N_2043,N_1957);
and U2140 (N_2140,N_2034,N_1874);
nor U2141 (N_2141,N_1930,N_2061);
and U2142 (N_2142,N_1985,N_1839);
nand U2143 (N_2143,N_1983,N_2096);
and U2144 (N_2144,N_1803,N_1818);
or U2145 (N_2145,N_2085,N_1856);
xnor U2146 (N_2146,N_1849,N_1920);
nand U2147 (N_2147,N_1860,N_2058);
nor U2148 (N_2148,N_1999,N_1812);
or U2149 (N_2149,N_1846,N_1987);
nor U2150 (N_2150,N_1881,N_1941);
nor U2151 (N_2151,N_1937,N_1829);
nor U2152 (N_2152,N_2077,N_1830);
xnor U2153 (N_2153,N_2084,N_2092);
xnor U2154 (N_2154,N_2027,N_2030);
nand U2155 (N_2155,N_1809,N_2075);
or U2156 (N_2156,N_2072,N_1989);
nor U2157 (N_2157,N_2059,N_1947);
nand U2158 (N_2158,N_1880,N_1842);
and U2159 (N_2159,N_2014,N_2029);
and U2160 (N_2160,N_2065,N_1823);
nand U2161 (N_2161,N_2089,N_1899);
nor U2162 (N_2162,N_1929,N_1984);
and U2163 (N_2163,N_2038,N_1833);
and U2164 (N_2164,N_1925,N_2010);
nor U2165 (N_2165,N_1896,N_1986);
nor U2166 (N_2166,N_2071,N_1807);
xnor U2167 (N_2167,N_1806,N_2040);
or U2168 (N_2168,N_1974,N_1907);
nor U2169 (N_2169,N_2094,N_2053);
xnor U2170 (N_2170,N_2020,N_1924);
xnor U2171 (N_2171,N_1992,N_1837);
nor U2172 (N_2172,N_1802,N_2093);
nand U2173 (N_2173,N_1968,N_2090);
and U2174 (N_2174,N_2056,N_2033);
nand U2175 (N_2175,N_1854,N_2009);
or U2176 (N_2176,N_1993,N_2006);
nor U2177 (N_2177,N_1921,N_2015);
or U2178 (N_2178,N_1971,N_1804);
and U2179 (N_2179,N_1909,N_1853);
or U2180 (N_2180,N_1903,N_1942);
nand U2181 (N_2181,N_1964,N_1954);
nor U2182 (N_2182,N_1814,N_1943);
nor U2183 (N_2183,N_2050,N_2052);
and U2184 (N_2184,N_2091,N_1908);
nand U2185 (N_2185,N_2041,N_1889);
and U2186 (N_2186,N_2099,N_1841);
and U2187 (N_2187,N_2057,N_2083);
nand U2188 (N_2188,N_1946,N_2019);
and U2189 (N_2189,N_1902,N_1965);
or U2190 (N_2190,N_1977,N_2035);
or U2191 (N_2191,N_2068,N_1952);
and U2192 (N_2192,N_1868,N_1927);
nor U2193 (N_2193,N_2021,N_1923);
or U2194 (N_2194,N_1962,N_1826);
xor U2195 (N_2195,N_2004,N_1958);
nand U2196 (N_2196,N_2069,N_1917);
and U2197 (N_2197,N_1998,N_1948);
and U2198 (N_2198,N_1911,N_1969);
and U2199 (N_2199,N_1872,N_2032);
or U2200 (N_2200,N_1871,N_1888);
nand U2201 (N_2201,N_1990,N_2087);
xnor U2202 (N_2202,N_1913,N_1813);
nor U2203 (N_2203,N_1939,N_1800);
nand U2204 (N_2204,N_1862,N_1879);
nor U2205 (N_2205,N_1845,N_1956);
or U2206 (N_2206,N_1895,N_1953);
nor U2207 (N_2207,N_1865,N_1912);
or U2208 (N_2208,N_1940,N_2013);
nor U2209 (N_2209,N_2042,N_1931);
nand U2210 (N_2210,N_2023,N_2000);
nor U2211 (N_2211,N_1918,N_2045);
nor U2212 (N_2212,N_1910,N_1915);
xnor U2213 (N_2213,N_1805,N_2082);
or U2214 (N_2214,N_1959,N_1834);
and U2215 (N_2215,N_1973,N_1843);
and U2216 (N_2216,N_1898,N_1882);
and U2217 (N_2217,N_1970,N_1972);
xor U2218 (N_2218,N_1863,N_1810);
xnor U2219 (N_2219,N_1949,N_1966);
xnor U2220 (N_2220,N_1869,N_1891);
and U2221 (N_2221,N_1935,N_2067);
nor U2222 (N_2222,N_2036,N_2048);
nand U2223 (N_2223,N_1811,N_2066);
and U2224 (N_2224,N_2046,N_1988);
nand U2225 (N_2225,N_1820,N_2047);
nor U2226 (N_2226,N_2097,N_1928);
xor U2227 (N_2227,N_1819,N_1892);
or U2228 (N_2228,N_1817,N_1816);
or U2229 (N_2229,N_2005,N_2079);
or U2230 (N_2230,N_1870,N_1922);
or U2231 (N_2231,N_1875,N_1867);
or U2232 (N_2232,N_1995,N_1815);
and U2233 (N_2233,N_1808,N_2076);
nor U2234 (N_2234,N_1894,N_1876);
or U2235 (N_2235,N_1859,N_1945);
xor U2236 (N_2236,N_1852,N_1991);
xor U2237 (N_2237,N_2063,N_1951);
nand U2238 (N_2238,N_1978,N_2012);
or U2239 (N_2239,N_1982,N_2037);
xnor U2240 (N_2240,N_1979,N_1801);
xor U2241 (N_2241,N_1822,N_1890);
and U2242 (N_2242,N_2062,N_1883);
or U2243 (N_2243,N_1885,N_1961);
nor U2244 (N_2244,N_1828,N_1866);
xnor U2245 (N_2245,N_2044,N_2088);
and U2246 (N_2246,N_2074,N_1832);
xnor U2247 (N_2247,N_1835,N_1901);
nor U2248 (N_2248,N_1836,N_1873);
nor U2249 (N_2249,N_2080,N_1976);
nand U2250 (N_2250,N_1859,N_1957);
and U2251 (N_2251,N_1834,N_1884);
nor U2252 (N_2252,N_2074,N_2061);
nand U2253 (N_2253,N_2032,N_1898);
or U2254 (N_2254,N_2067,N_1924);
nand U2255 (N_2255,N_2088,N_1842);
nor U2256 (N_2256,N_1866,N_1867);
nor U2257 (N_2257,N_2035,N_1979);
nand U2258 (N_2258,N_2063,N_2077);
or U2259 (N_2259,N_1954,N_1931);
or U2260 (N_2260,N_2029,N_1893);
xnor U2261 (N_2261,N_1998,N_1886);
xor U2262 (N_2262,N_1885,N_2020);
nor U2263 (N_2263,N_1815,N_1903);
nor U2264 (N_2264,N_1878,N_1889);
nor U2265 (N_2265,N_2099,N_1819);
nor U2266 (N_2266,N_2001,N_1818);
nor U2267 (N_2267,N_1934,N_1863);
nor U2268 (N_2268,N_1996,N_2023);
xor U2269 (N_2269,N_2035,N_2055);
nand U2270 (N_2270,N_1822,N_2094);
nand U2271 (N_2271,N_2046,N_1937);
and U2272 (N_2272,N_2064,N_1981);
xor U2273 (N_2273,N_2030,N_1942);
xnor U2274 (N_2274,N_1968,N_1812);
xor U2275 (N_2275,N_1868,N_1984);
nor U2276 (N_2276,N_2076,N_1944);
nand U2277 (N_2277,N_1824,N_1936);
xnor U2278 (N_2278,N_2035,N_1976);
xor U2279 (N_2279,N_1982,N_1844);
or U2280 (N_2280,N_1834,N_1913);
nor U2281 (N_2281,N_1977,N_1857);
or U2282 (N_2282,N_1819,N_2029);
nand U2283 (N_2283,N_1855,N_1866);
nor U2284 (N_2284,N_1984,N_2031);
and U2285 (N_2285,N_1988,N_2089);
xnor U2286 (N_2286,N_1973,N_1841);
nand U2287 (N_2287,N_2028,N_1927);
xnor U2288 (N_2288,N_1937,N_2000);
nand U2289 (N_2289,N_2008,N_1864);
or U2290 (N_2290,N_2097,N_1982);
and U2291 (N_2291,N_1848,N_1826);
nor U2292 (N_2292,N_1896,N_1931);
nand U2293 (N_2293,N_1915,N_1928);
or U2294 (N_2294,N_1893,N_1974);
nor U2295 (N_2295,N_2016,N_1829);
or U2296 (N_2296,N_1831,N_2037);
or U2297 (N_2297,N_1853,N_1845);
nor U2298 (N_2298,N_2071,N_1874);
nor U2299 (N_2299,N_2087,N_2061);
or U2300 (N_2300,N_2093,N_1933);
nand U2301 (N_2301,N_1817,N_1836);
xor U2302 (N_2302,N_1919,N_2022);
xnor U2303 (N_2303,N_2058,N_1936);
and U2304 (N_2304,N_1886,N_2006);
and U2305 (N_2305,N_2070,N_1974);
xor U2306 (N_2306,N_2034,N_1945);
and U2307 (N_2307,N_1954,N_1941);
nand U2308 (N_2308,N_1809,N_1807);
and U2309 (N_2309,N_1897,N_1978);
nand U2310 (N_2310,N_1996,N_2057);
and U2311 (N_2311,N_1881,N_1986);
nand U2312 (N_2312,N_1949,N_1926);
or U2313 (N_2313,N_2020,N_2008);
and U2314 (N_2314,N_1848,N_1926);
nand U2315 (N_2315,N_1954,N_2008);
nor U2316 (N_2316,N_1806,N_1945);
or U2317 (N_2317,N_1971,N_1836);
xnor U2318 (N_2318,N_2092,N_2017);
or U2319 (N_2319,N_1824,N_1820);
nor U2320 (N_2320,N_1840,N_1846);
nor U2321 (N_2321,N_1913,N_2068);
nor U2322 (N_2322,N_1951,N_1962);
and U2323 (N_2323,N_2036,N_1846);
xor U2324 (N_2324,N_1850,N_1913);
xor U2325 (N_2325,N_1882,N_1945);
nand U2326 (N_2326,N_2072,N_1866);
and U2327 (N_2327,N_1933,N_1891);
and U2328 (N_2328,N_2098,N_1823);
nor U2329 (N_2329,N_2042,N_1917);
xor U2330 (N_2330,N_2096,N_2051);
and U2331 (N_2331,N_1848,N_1999);
and U2332 (N_2332,N_1989,N_1812);
xor U2333 (N_2333,N_1872,N_1815);
nor U2334 (N_2334,N_1953,N_2093);
and U2335 (N_2335,N_2021,N_1984);
or U2336 (N_2336,N_1871,N_1959);
and U2337 (N_2337,N_1900,N_1844);
or U2338 (N_2338,N_1941,N_1879);
or U2339 (N_2339,N_1902,N_2032);
and U2340 (N_2340,N_1911,N_1879);
or U2341 (N_2341,N_1964,N_2066);
xor U2342 (N_2342,N_1972,N_2013);
and U2343 (N_2343,N_1867,N_1964);
nand U2344 (N_2344,N_1835,N_1825);
nand U2345 (N_2345,N_2055,N_2046);
xnor U2346 (N_2346,N_1814,N_1935);
or U2347 (N_2347,N_2099,N_1971);
and U2348 (N_2348,N_1951,N_2027);
xnor U2349 (N_2349,N_2069,N_1939);
or U2350 (N_2350,N_1848,N_1897);
and U2351 (N_2351,N_2000,N_1809);
nand U2352 (N_2352,N_1866,N_1976);
and U2353 (N_2353,N_1994,N_1967);
or U2354 (N_2354,N_1844,N_1823);
xor U2355 (N_2355,N_1841,N_1855);
or U2356 (N_2356,N_1997,N_1970);
or U2357 (N_2357,N_1956,N_1831);
and U2358 (N_2358,N_1922,N_1985);
or U2359 (N_2359,N_1900,N_1870);
or U2360 (N_2360,N_1885,N_1912);
nand U2361 (N_2361,N_2013,N_1865);
xor U2362 (N_2362,N_1950,N_1930);
xnor U2363 (N_2363,N_1975,N_2032);
nor U2364 (N_2364,N_1814,N_2045);
nor U2365 (N_2365,N_2087,N_1988);
xnor U2366 (N_2366,N_2042,N_1916);
and U2367 (N_2367,N_2070,N_1982);
or U2368 (N_2368,N_1823,N_1833);
or U2369 (N_2369,N_1884,N_1964);
or U2370 (N_2370,N_2000,N_1964);
nand U2371 (N_2371,N_1897,N_2045);
nor U2372 (N_2372,N_1899,N_1809);
or U2373 (N_2373,N_1896,N_1980);
and U2374 (N_2374,N_1839,N_2081);
and U2375 (N_2375,N_1957,N_1904);
nand U2376 (N_2376,N_1909,N_1840);
xnor U2377 (N_2377,N_1962,N_2053);
nand U2378 (N_2378,N_1872,N_1817);
or U2379 (N_2379,N_2080,N_1981);
xor U2380 (N_2380,N_2042,N_1804);
and U2381 (N_2381,N_1902,N_2073);
nand U2382 (N_2382,N_1855,N_2048);
nor U2383 (N_2383,N_1844,N_1906);
or U2384 (N_2384,N_1992,N_1812);
or U2385 (N_2385,N_2012,N_1903);
nand U2386 (N_2386,N_2031,N_1997);
and U2387 (N_2387,N_1997,N_1853);
nor U2388 (N_2388,N_2095,N_1844);
and U2389 (N_2389,N_1917,N_1912);
and U2390 (N_2390,N_2056,N_1867);
nand U2391 (N_2391,N_1916,N_1958);
nor U2392 (N_2392,N_1843,N_2042);
nor U2393 (N_2393,N_2059,N_1917);
or U2394 (N_2394,N_1838,N_1825);
nand U2395 (N_2395,N_1827,N_2068);
and U2396 (N_2396,N_2088,N_1912);
xnor U2397 (N_2397,N_1849,N_1834);
and U2398 (N_2398,N_2001,N_1858);
xor U2399 (N_2399,N_2028,N_1861);
nor U2400 (N_2400,N_2336,N_2189);
xor U2401 (N_2401,N_2131,N_2371);
nor U2402 (N_2402,N_2350,N_2232);
or U2403 (N_2403,N_2139,N_2345);
nor U2404 (N_2404,N_2134,N_2164);
nand U2405 (N_2405,N_2317,N_2275);
nor U2406 (N_2406,N_2160,N_2279);
xnor U2407 (N_2407,N_2215,N_2354);
and U2408 (N_2408,N_2274,N_2294);
nor U2409 (N_2409,N_2281,N_2322);
nand U2410 (N_2410,N_2302,N_2168);
nor U2411 (N_2411,N_2321,N_2363);
nor U2412 (N_2412,N_2397,N_2228);
or U2413 (N_2413,N_2209,N_2153);
xor U2414 (N_2414,N_2102,N_2187);
or U2415 (N_2415,N_2188,N_2283);
and U2416 (N_2416,N_2148,N_2115);
nand U2417 (N_2417,N_2375,N_2185);
nand U2418 (N_2418,N_2266,N_2123);
xnor U2419 (N_2419,N_2229,N_2258);
nand U2420 (N_2420,N_2328,N_2181);
nand U2421 (N_2421,N_2137,N_2373);
nand U2422 (N_2422,N_2374,N_2313);
xnor U2423 (N_2423,N_2344,N_2101);
nor U2424 (N_2424,N_2211,N_2332);
or U2425 (N_2425,N_2305,N_2262);
or U2426 (N_2426,N_2169,N_2117);
xor U2427 (N_2427,N_2120,N_2203);
nor U2428 (N_2428,N_2114,N_2323);
xnor U2429 (N_2429,N_2360,N_2179);
nor U2430 (N_2430,N_2394,N_2196);
nand U2431 (N_2431,N_2106,N_2361);
or U2432 (N_2432,N_2233,N_2204);
xnor U2433 (N_2433,N_2158,N_2105);
xnor U2434 (N_2434,N_2273,N_2263);
or U2435 (N_2435,N_2355,N_2248);
xnor U2436 (N_2436,N_2372,N_2167);
nor U2437 (N_2437,N_2175,N_2316);
xor U2438 (N_2438,N_2369,N_2132);
xor U2439 (N_2439,N_2172,N_2260);
and U2440 (N_2440,N_2318,N_2380);
nor U2441 (N_2441,N_2225,N_2383);
xnor U2442 (N_2442,N_2385,N_2240);
xor U2443 (N_2443,N_2100,N_2338);
and U2444 (N_2444,N_2220,N_2312);
nand U2445 (N_2445,N_2370,N_2269);
or U2446 (N_2446,N_2112,N_2346);
nand U2447 (N_2447,N_2116,N_2184);
xor U2448 (N_2448,N_2324,N_2251);
nor U2449 (N_2449,N_2339,N_2253);
nor U2450 (N_2450,N_2108,N_2288);
nor U2451 (N_2451,N_2280,N_2300);
nand U2452 (N_2452,N_2238,N_2265);
or U2453 (N_2453,N_2191,N_2311);
nor U2454 (N_2454,N_2314,N_2118);
xnor U2455 (N_2455,N_2208,N_2237);
and U2456 (N_2456,N_2119,N_2310);
nand U2457 (N_2457,N_2366,N_2340);
nand U2458 (N_2458,N_2190,N_2195);
or U2459 (N_2459,N_2287,N_2277);
or U2460 (N_2460,N_2399,N_2392);
xor U2461 (N_2461,N_2296,N_2149);
nor U2462 (N_2462,N_2103,N_2154);
nor U2463 (N_2463,N_2387,N_2356);
xor U2464 (N_2464,N_2290,N_2192);
nor U2465 (N_2465,N_2161,N_2171);
xnor U2466 (N_2466,N_2284,N_2271);
and U2467 (N_2467,N_2197,N_2291);
xor U2468 (N_2468,N_2259,N_2176);
and U2469 (N_2469,N_2157,N_2151);
nor U2470 (N_2470,N_2330,N_2140);
or U2471 (N_2471,N_2236,N_2341);
nand U2472 (N_2472,N_2303,N_2193);
xnor U2473 (N_2473,N_2173,N_2264);
and U2474 (N_2474,N_2217,N_2395);
nor U2475 (N_2475,N_2145,N_2147);
nor U2476 (N_2476,N_2272,N_2194);
nand U2477 (N_2477,N_2143,N_2234);
nor U2478 (N_2478,N_2342,N_2122);
and U2479 (N_2479,N_2301,N_2216);
nand U2480 (N_2480,N_2349,N_2390);
and U2481 (N_2481,N_2141,N_2227);
nand U2482 (N_2482,N_2268,N_2249);
xor U2483 (N_2483,N_2327,N_2389);
and U2484 (N_2484,N_2252,N_2396);
or U2485 (N_2485,N_2309,N_2335);
or U2486 (N_2486,N_2221,N_2368);
xor U2487 (N_2487,N_2223,N_2359);
nand U2488 (N_2488,N_2174,N_2198);
and U2489 (N_2489,N_2384,N_2130);
nand U2490 (N_2490,N_2230,N_2376);
and U2491 (N_2491,N_2150,N_2207);
xnor U2492 (N_2492,N_2166,N_2186);
and U2493 (N_2493,N_2124,N_2126);
and U2494 (N_2494,N_2241,N_2121);
xor U2495 (N_2495,N_2333,N_2261);
nor U2496 (N_2496,N_2243,N_2177);
and U2497 (N_2497,N_2381,N_2199);
nand U2498 (N_2498,N_2136,N_2180);
nor U2499 (N_2499,N_2170,N_2247);
nand U2500 (N_2500,N_2152,N_2325);
nand U2501 (N_2501,N_2178,N_2348);
nand U2502 (N_2502,N_2182,N_2214);
xnor U2503 (N_2503,N_2365,N_2398);
and U2504 (N_2504,N_2219,N_2289);
xnor U2505 (N_2505,N_2377,N_2210);
or U2506 (N_2506,N_2133,N_2319);
or U2507 (N_2507,N_2218,N_2297);
or U2508 (N_2508,N_2292,N_2304);
and U2509 (N_2509,N_2326,N_2200);
nor U2510 (N_2510,N_2162,N_2267);
xnor U2511 (N_2511,N_2226,N_2125);
and U2512 (N_2512,N_2293,N_2159);
and U2513 (N_2513,N_2331,N_2308);
xor U2514 (N_2514,N_2347,N_2183);
xor U2515 (N_2515,N_2382,N_2111);
nand U2516 (N_2516,N_2250,N_2224);
nand U2517 (N_2517,N_2128,N_2282);
and U2518 (N_2518,N_2129,N_2343);
or U2519 (N_2519,N_2286,N_2276);
xnor U2520 (N_2520,N_2127,N_2353);
nand U2521 (N_2521,N_2242,N_2142);
nor U2522 (N_2522,N_2155,N_2379);
xor U2523 (N_2523,N_2107,N_2367);
and U2524 (N_2524,N_2222,N_2144);
and U2525 (N_2525,N_2388,N_2205);
nand U2526 (N_2526,N_2138,N_2362);
and U2527 (N_2527,N_2270,N_2206);
nor U2528 (N_2528,N_2163,N_2306);
nor U2529 (N_2529,N_2358,N_2231);
and U2530 (N_2530,N_2254,N_2298);
nand U2531 (N_2531,N_2256,N_2299);
and U2532 (N_2532,N_2351,N_2255);
xor U2533 (N_2533,N_2235,N_2165);
xnor U2534 (N_2534,N_2391,N_2334);
xnor U2535 (N_2535,N_2386,N_2320);
xor U2536 (N_2536,N_2295,N_2245);
or U2537 (N_2537,N_2357,N_2239);
and U2538 (N_2538,N_2109,N_2156);
nand U2539 (N_2539,N_2244,N_2246);
nand U2540 (N_2540,N_2337,N_2278);
or U2541 (N_2541,N_2202,N_2104);
or U2542 (N_2542,N_2329,N_2201);
nor U2543 (N_2543,N_2285,N_2110);
or U2544 (N_2544,N_2257,N_2352);
xor U2545 (N_2545,N_2315,N_2307);
nor U2546 (N_2546,N_2393,N_2378);
nor U2547 (N_2547,N_2213,N_2135);
xnor U2548 (N_2548,N_2146,N_2212);
nor U2549 (N_2549,N_2113,N_2364);
xnor U2550 (N_2550,N_2184,N_2173);
nor U2551 (N_2551,N_2115,N_2396);
and U2552 (N_2552,N_2295,N_2277);
nand U2553 (N_2553,N_2124,N_2291);
nor U2554 (N_2554,N_2243,N_2175);
xnor U2555 (N_2555,N_2314,N_2188);
or U2556 (N_2556,N_2223,N_2229);
nor U2557 (N_2557,N_2301,N_2214);
xnor U2558 (N_2558,N_2272,N_2228);
and U2559 (N_2559,N_2218,N_2129);
xor U2560 (N_2560,N_2308,N_2102);
nand U2561 (N_2561,N_2114,N_2160);
or U2562 (N_2562,N_2256,N_2186);
nor U2563 (N_2563,N_2386,N_2330);
and U2564 (N_2564,N_2300,N_2177);
xor U2565 (N_2565,N_2111,N_2118);
nor U2566 (N_2566,N_2314,N_2142);
or U2567 (N_2567,N_2329,N_2225);
nor U2568 (N_2568,N_2229,N_2349);
nand U2569 (N_2569,N_2142,N_2274);
or U2570 (N_2570,N_2319,N_2240);
nor U2571 (N_2571,N_2360,N_2267);
nand U2572 (N_2572,N_2346,N_2254);
nand U2573 (N_2573,N_2101,N_2105);
and U2574 (N_2574,N_2214,N_2355);
nor U2575 (N_2575,N_2148,N_2271);
and U2576 (N_2576,N_2248,N_2113);
and U2577 (N_2577,N_2236,N_2343);
xnor U2578 (N_2578,N_2349,N_2395);
nand U2579 (N_2579,N_2231,N_2274);
xor U2580 (N_2580,N_2397,N_2261);
or U2581 (N_2581,N_2350,N_2269);
nand U2582 (N_2582,N_2177,N_2200);
and U2583 (N_2583,N_2249,N_2378);
nor U2584 (N_2584,N_2326,N_2248);
nand U2585 (N_2585,N_2287,N_2148);
nand U2586 (N_2586,N_2256,N_2383);
nand U2587 (N_2587,N_2239,N_2211);
or U2588 (N_2588,N_2334,N_2257);
nand U2589 (N_2589,N_2154,N_2167);
nor U2590 (N_2590,N_2224,N_2327);
nand U2591 (N_2591,N_2238,N_2335);
nand U2592 (N_2592,N_2224,N_2309);
and U2593 (N_2593,N_2395,N_2207);
or U2594 (N_2594,N_2128,N_2288);
and U2595 (N_2595,N_2298,N_2338);
nor U2596 (N_2596,N_2320,N_2282);
nand U2597 (N_2597,N_2142,N_2148);
or U2598 (N_2598,N_2240,N_2244);
and U2599 (N_2599,N_2100,N_2262);
and U2600 (N_2600,N_2111,N_2174);
and U2601 (N_2601,N_2262,N_2110);
and U2602 (N_2602,N_2345,N_2104);
nand U2603 (N_2603,N_2243,N_2165);
xor U2604 (N_2604,N_2305,N_2235);
nand U2605 (N_2605,N_2254,N_2338);
nand U2606 (N_2606,N_2137,N_2202);
or U2607 (N_2607,N_2188,N_2194);
xor U2608 (N_2608,N_2248,N_2331);
xor U2609 (N_2609,N_2141,N_2226);
and U2610 (N_2610,N_2144,N_2125);
or U2611 (N_2611,N_2227,N_2310);
nor U2612 (N_2612,N_2171,N_2365);
xnor U2613 (N_2613,N_2169,N_2229);
xor U2614 (N_2614,N_2137,N_2267);
nor U2615 (N_2615,N_2195,N_2388);
nand U2616 (N_2616,N_2218,N_2347);
nor U2617 (N_2617,N_2138,N_2370);
and U2618 (N_2618,N_2242,N_2310);
xnor U2619 (N_2619,N_2176,N_2388);
xnor U2620 (N_2620,N_2273,N_2134);
xnor U2621 (N_2621,N_2348,N_2188);
or U2622 (N_2622,N_2174,N_2183);
nand U2623 (N_2623,N_2150,N_2358);
xor U2624 (N_2624,N_2251,N_2107);
nor U2625 (N_2625,N_2269,N_2318);
and U2626 (N_2626,N_2203,N_2195);
xor U2627 (N_2627,N_2104,N_2349);
xor U2628 (N_2628,N_2363,N_2209);
nand U2629 (N_2629,N_2374,N_2280);
or U2630 (N_2630,N_2279,N_2341);
xor U2631 (N_2631,N_2332,N_2217);
or U2632 (N_2632,N_2188,N_2167);
nand U2633 (N_2633,N_2148,N_2321);
or U2634 (N_2634,N_2232,N_2386);
and U2635 (N_2635,N_2196,N_2118);
xnor U2636 (N_2636,N_2293,N_2267);
xnor U2637 (N_2637,N_2191,N_2147);
xnor U2638 (N_2638,N_2307,N_2179);
nor U2639 (N_2639,N_2192,N_2179);
or U2640 (N_2640,N_2112,N_2198);
or U2641 (N_2641,N_2182,N_2255);
nor U2642 (N_2642,N_2173,N_2335);
nand U2643 (N_2643,N_2316,N_2322);
nor U2644 (N_2644,N_2190,N_2242);
xnor U2645 (N_2645,N_2241,N_2300);
nor U2646 (N_2646,N_2398,N_2346);
and U2647 (N_2647,N_2173,N_2276);
and U2648 (N_2648,N_2309,N_2393);
xor U2649 (N_2649,N_2376,N_2351);
and U2650 (N_2650,N_2332,N_2356);
xnor U2651 (N_2651,N_2308,N_2167);
and U2652 (N_2652,N_2364,N_2138);
or U2653 (N_2653,N_2333,N_2212);
or U2654 (N_2654,N_2396,N_2254);
xor U2655 (N_2655,N_2399,N_2149);
nor U2656 (N_2656,N_2195,N_2184);
nor U2657 (N_2657,N_2181,N_2156);
and U2658 (N_2658,N_2197,N_2372);
or U2659 (N_2659,N_2357,N_2179);
nor U2660 (N_2660,N_2234,N_2368);
xor U2661 (N_2661,N_2216,N_2317);
xor U2662 (N_2662,N_2138,N_2118);
xnor U2663 (N_2663,N_2199,N_2164);
or U2664 (N_2664,N_2102,N_2323);
xnor U2665 (N_2665,N_2162,N_2274);
or U2666 (N_2666,N_2347,N_2253);
or U2667 (N_2667,N_2391,N_2344);
and U2668 (N_2668,N_2282,N_2161);
or U2669 (N_2669,N_2283,N_2248);
or U2670 (N_2670,N_2279,N_2312);
xor U2671 (N_2671,N_2325,N_2334);
and U2672 (N_2672,N_2126,N_2134);
nor U2673 (N_2673,N_2149,N_2233);
nand U2674 (N_2674,N_2318,N_2133);
xnor U2675 (N_2675,N_2273,N_2112);
or U2676 (N_2676,N_2355,N_2270);
xor U2677 (N_2677,N_2343,N_2271);
nor U2678 (N_2678,N_2109,N_2312);
nor U2679 (N_2679,N_2195,N_2261);
nor U2680 (N_2680,N_2128,N_2138);
xor U2681 (N_2681,N_2379,N_2262);
or U2682 (N_2682,N_2354,N_2204);
nor U2683 (N_2683,N_2391,N_2191);
nor U2684 (N_2684,N_2245,N_2379);
nand U2685 (N_2685,N_2275,N_2234);
nand U2686 (N_2686,N_2161,N_2268);
nor U2687 (N_2687,N_2127,N_2321);
and U2688 (N_2688,N_2153,N_2259);
nor U2689 (N_2689,N_2313,N_2252);
nor U2690 (N_2690,N_2132,N_2376);
xnor U2691 (N_2691,N_2250,N_2340);
or U2692 (N_2692,N_2310,N_2236);
nor U2693 (N_2693,N_2129,N_2195);
nor U2694 (N_2694,N_2262,N_2323);
nand U2695 (N_2695,N_2251,N_2311);
or U2696 (N_2696,N_2361,N_2353);
xnor U2697 (N_2697,N_2397,N_2174);
or U2698 (N_2698,N_2253,N_2274);
xnor U2699 (N_2699,N_2175,N_2287);
xnor U2700 (N_2700,N_2533,N_2687);
and U2701 (N_2701,N_2625,N_2597);
xor U2702 (N_2702,N_2556,N_2476);
or U2703 (N_2703,N_2524,N_2509);
nand U2704 (N_2704,N_2599,N_2691);
xor U2705 (N_2705,N_2628,N_2418);
nor U2706 (N_2706,N_2560,N_2645);
nor U2707 (N_2707,N_2589,N_2424);
nand U2708 (N_2708,N_2467,N_2483);
nand U2709 (N_2709,N_2477,N_2499);
nor U2710 (N_2710,N_2671,N_2505);
and U2711 (N_2711,N_2596,N_2503);
xor U2712 (N_2712,N_2595,N_2683);
nor U2713 (N_2713,N_2571,N_2496);
xnor U2714 (N_2714,N_2416,N_2414);
nor U2715 (N_2715,N_2634,N_2449);
and U2716 (N_2716,N_2610,N_2504);
xnor U2717 (N_2717,N_2549,N_2622);
nand U2718 (N_2718,N_2619,N_2434);
nand U2719 (N_2719,N_2605,N_2540);
nand U2720 (N_2720,N_2576,N_2603);
xor U2721 (N_2721,N_2523,N_2400);
xor U2722 (N_2722,N_2647,N_2402);
and U2723 (N_2723,N_2561,N_2443);
or U2724 (N_2724,N_2427,N_2641);
nand U2725 (N_2725,N_2696,N_2470);
nor U2726 (N_2726,N_2694,N_2654);
nor U2727 (N_2727,N_2425,N_2543);
nand U2728 (N_2728,N_2542,N_2611);
nor U2729 (N_2729,N_2629,N_2659);
xnor U2730 (N_2730,N_2612,N_2668);
xor U2731 (N_2731,N_2472,N_2649);
nand U2732 (N_2732,N_2521,N_2495);
nand U2733 (N_2733,N_2604,N_2493);
xnor U2734 (N_2734,N_2453,N_2591);
and U2735 (N_2735,N_2441,N_2490);
and U2736 (N_2736,N_2422,N_2586);
nor U2737 (N_2737,N_2455,N_2460);
xor U2738 (N_2738,N_2680,N_2658);
nor U2739 (N_2739,N_2466,N_2436);
nor U2740 (N_2740,N_2590,N_2579);
nand U2741 (N_2741,N_2473,N_2551);
nand U2742 (N_2742,N_2512,N_2581);
and U2743 (N_2743,N_2567,N_2428);
or U2744 (N_2744,N_2663,N_2463);
nor U2745 (N_2745,N_2617,N_2577);
xnor U2746 (N_2746,N_2609,N_2423);
xor U2747 (N_2747,N_2410,N_2624);
nand U2748 (N_2748,N_2502,N_2620);
xor U2749 (N_2749,N_2479,N_2448);
xor U2750 (N_2750,N_2475,N_2646);
and U2751 (N_2751,N_2638,N_2644);
and U2752 (N_2752,N_2553,N_2614);
nor U2753 (N_2753,N_2451,N_2534);
nand U2754 (N_2754,N_2661,N_2537);
xor U2755 (N_2755,N_2676,N_2606);
nor U2756 (N_2756,N_2440,N_2584);
nor U2757 (N_2757,N_2552,N_2690);
or U2758 (N_2758,N_2627,N_2678);
xnor U2759 (N_2759,N_2615,N_2442);
and U2760 (N_2760,N_2421,N_2562);
nor U2761 (N_2761,N_2471,N_2665);
or U2762 (N_2762,N_2573,N_2588);
xnor U2763 (N_2763,N_2404,N_2631);
or U2764 (N_2764,N_2454,N_2517);
nand U2765 (N_2765,N_2693,N_2653);
and U2766 (N_2766,N_2594,N_2420);
nand U2767 (N_2767,N_2557,N_2510);
nand U2768 (N_2768,N_2593,N_2569);
nor U2769 (N_2769,N_2616,N_2530);
nor U2770 (N_2770,N_2488,N_2478);
xnor U2771 (N_2771,N_2667,N_2408);
xnor U2772 (N_2772,N_2640,N_2623);
or U2773 (N_2773,N_2585,N_2600);
nor U2774 (N_2774,N_2660,N_2575);
nand U2775 (N_2775,N_2608,N_2698);
or U2776 (N_2776,N_2635,N_2452);
or U2777 (N_2777,N_2474,N_2480);
nand U2778 (N_2778,N_2511,N_2558);
xor U2779 (N_2779,N_2679,N_2652);
xnor U2780 (N_2780,N_2431,N_2547);
or U2781 (N_2781,N_2633,N_2695);
nand U2782 (N_2782,N_2529,N_2626);
xnor U2783 (N_2783,N_2648,N_2458);
nand U2784 (N_2784,N_2437,N_2439);
nand U2785 (N_2785,N_2486,N_2692);
nand U2786 (N_2786,N_2566,N_2525);
and U2787 (N_2787,N_2592,N_2446);
xnor U2788 (N_2788,N_2494,N_2528);
and U2789 (N_2789,N_2681,N_2580);
xnor U2790 (N_2790,N_2492,N_2587);
and U2791 (N_2791,N_2657,N_2674);
nor U2792 (N_2792,N_2430,N_2539);
or U2793 (N_2793,N_2656,N_2447);
nor U2794 (N_2794,N_2618,N_2482);
xnor U2795 (N_2795,N_2429,N_2677);
xnor U2796 (N_2796,N_2670,N_2438);
or U2797 (N_2797,N_2484,N_2538);
nand U2798 (N_2798,N_2456,N_2563);
nand U2799 (N_2799,N_2415,N_2621);
and U2800 (N_2800,N_2426,N_2630);
xor U2801 (N_2801,N_2675,N_2544);
xor U2802 (N_2802,N_2672,N_2464);
xor U2803 (N_2803,N_2686,N_2527);
and U2804 (N_2804,N_2688,N_2462);
or U2805 (N_2805,N_2444,N_2574);
xnor U2806 (N_2806,N_2699,N_2637);
nand U2807 (N_2807,N_2459,N_2532);
and U2808 (N_2808,N_2689,N_2445);
nand U2809 (N_2809,N_2412,N_2497);
and U2810 (N_2810,N_2664,N_2519);
nand U2811 (N_2811,N_2601,N_2669);
or U2812 (N_2812,N_2536,N_2406);
nor U2813 (N_2813,N_2651,N_2632);
nor U2814 (N_2814,N_2465,N_2643);
and U2815 (N_2815,N_2541,N_2583);
nand U2816 (N_2816,N_2468,N_2531);
and U2817 (N_2817,N_2535,N_2582);
xnor U2818 (N_2818,N_2507,N_2401);
nor U2819 (N_2819,N_2554,N_2602);
nor U2820 (N_2820,N_2433,N_2548);
nand U2821 (N_2821,N_2489,N_2682);
or U2822 (N_2822,N_2650,N_2491);
nor U2823 (N_2823,N_2550,N_2508);
xnor U2824 (N_2824,N_2545,N_2405);
xnor U2825 (N_2825,N_2655,N_2501);
or U2826 (N_2826,N_2555,N_2515);
or U2827 (N_2827,N_2513,N_2565);
or U2828 (N_2828,N_2435,N_2498);
and U2829 (N_2829,N_2673,N_2526);
xnor U2830 (N_2830,N_2636,N_2432);
or U2831 (N_2831,N_2559,N_2411);
nor U2832 (N_2832,N_2546,N_2607);
and U2833 (N_2833,N_2578,N_2516);
nand U2834 (N_2834,N_2572,N_2485);
nor U2835 (N_2835,N_2518,N_2666);
nand U2836 (N_2836,N_2662,N_2685);
xor U2837 (N_2837,N_2413,N_2570);
xor U2838 (N_2838,N_2642,N_2568);
or U2839 (N_2839,N_2417,N_2461);
and U2840 (N_2840,N_2520,N_2409);
xor U2841 (N_2841,N_2500,N_2481);
xnor U2842 (N_2842,N_2506,N_2450);
nand U2843 (N_2843,N_2457,N_2564);
and U2844 (N_2844,N_2487,N_2522);
nor U2845 (N_2845,N_2613,N_2598);
nor U2846 (N_2846,N_2514,N_2639);
and U2847 (N_2847,N_2407,N_2684);
nand U2848 (N_2848,N_2419,N_2403);
and U2849 (N_2849,N_2697,N_2469);
nand U2850 (N_2850,N_2575,N_2686);
xnor U2851 (N_2851,N_2403,N_2550);
nand U2852 (N_2852,N_2453,N_2568);
xor U2853 (N_2853,N_2629,N_2524);
nand U2854 (N_2854,N_2587,N_2653);
xnor U2855 (N_2855,N_2684,N_2678);
and U2856 (N_2856,N_2468,N_2491);
nor U2857 (N_2857,N_2565,N_2603);
nand U2858 (N_2858,N_2417,N_2498);
nor U2859 (N_2859,N_2476,N_2628);
nand U2860 (N_2860,N_2545,N_2640);
nor U2861 (N_2861,N_2643,N_2457);
or U2862 (N_2862,N_2531,N_2588);
nand U2863 (N_2863,N_2588,N_2574);
xnor U2864 (N_2864,N_2621,N_2574);
and U2865 (N_2865,N_2516,N_2660);
and U2866 (N_2866,N_2584,N_2402);
nand U2867 (N_2867,N_2427,N_2457);
nor U2868 (N_2868,N_2558,N_2522);
and U2869 (N_2869,N_2545,N_2425);
xnor U2870 (N_2870,N_2698,N_2431);
nor U2871 (N_2871,N_2667,N_2616);
nor U2872 (N_2872,N_2511,N_2516);
nor U2873 (N_2873,N_2511,N_2648);
xnor U2874 (N_2874,N_2525,N_2491);
xnor U2875 (N_2875,N_2612,N_2622);
nand U2876 (N_2876,N_2531,N_2426);
and U2877 (N_2877,N_2503,N_2423);
and U2878 (N_2878,N_2514,N_2511);
nor U2879 (N_2879,N_2629,N_2621);
and U2880 (N_2880,N_2557,N_2561);
nand U2881 (N_2881,N_2556,N_2518);
xnor U2882 (N_2882,N_2548,N_2602);
nand U2883 (N_2883,N_2695,N_2573);
nor U2884 (N_2884,N_2458,N_2578);
xnor U2885 (N_2885,N_2468,N_2408);
and U2886 (N_2886,N_2657,N_2552);
xnor U2887 (N_2887,N_2489,N_2494);
xor U2888 (N_2888,N_2534,N_2602);
nand U2889 (N_2889,N_2648,N_2560);
and U2890 (N_2890,N_2590,N_2528);
nor U2891 (N_2891,N_2657,N_2589);
nor U2892 (N_2892,N_2418,N_2530);
and U2893 (N_2893,N_2666,N_2555);
nor U2894 (N_2894,N_2499,N_2419);
nor U2895 (N_2895,N_2440,N_2631);
nor U2896 (N_2896,N_2571,N_2629);
xor U2897 (N_2897,N_2672,N_2687);
nor U2898 (N_2898,N_2473,N_2666);
xor U2899 (N_2899,N_2467,N_2566);
nand U2900 (N_2900,N_2623,N_2588);
or U2901 (N_2901,N_2454,N_2430);
or U2902 (N_2902,N_2569,N_2480);
nor U2903 (N_2903,N_2478,N_2652);
and U2904 (N_2904,N_2574,N_2667);
or U2905 (N_2905,N_2574,N_2440);
nand U2906 (N_2906,N_2668,N_2557);
or U2907 (N_2907,N_2659,N_2461);
nand U2908 (N_2908,N_2593,N_2588);
xor U2909 (N_2909,N_2649,N_2430);
or U2910 (N_2910,N_2580,N_2517);
and U2911 (N_2911,N_2672,N_2463);
or U2912 (N_2912,N_2490,N_2574);
xor U2913 (N_2913,N_2695,N_2694);
or U2914 (N_2914,N_2655,N_2550);
xor U2915 (N_2915,N_2508,N_2493);
or U2916 (N_2916,N_2410,N_2570);
or U2917 (N_2917,N_2637,N_2657);
and U2918 (N_2918,N_2552,N_2462);
nor U2919 (N_2919,N_2515,N_2523);
nand U2920 (N_2920,N_2480,N_2497);
and U2921 (N_2921,N_2692,N_2551);
or U2922 (N_2922,N_2644,N_2523);
xor U2923 (N_2923,N_2599,N_2479);
or U2924 (N_2924,N_2400,N_2538);
nor U2925 (N_2925,N_2514,N_2513);
and U2926 (N_2926,N_2619,N_2691);
or U2927 (N_2927,N_2429,N_2587);
nor U2928 (N_2928,N_2535,N_2616);
xor U2929 (N_2929,N_2448,N_2552);
and U2930 (N_2930,N_2578,N_2674);
and U2931 (N_2931,N_2475,N_2556);
nor U2932 (N_2932,N_2440,N_2503);
xnor U2933 (N_2933,N_2669,N_2622);
nor U2934 (N_2934,N_2541,N_2507);
xnor U2935 (N_2935,N_2489,N_2517);
and U2936 (N_2936,N_2691,N_2429);
or U2937 (N_2937,N_2612,N_2527);
nand U2938 (N_2938,N_2674,N_2661);
nor U2939 (N_2939,N_2554,N_2539);
and U2940 (N_2940,N_2452,N_2506);
nand U2941 (N_2941,N_2494,N_2565);
nand U2942 (N_2942,N_2643,N_2560);
nor U2943 (N_2943,N_2427,N_2414);
xor U2944 (N_2944,N_2467,N_2536);
nand U2945 (N_2945,N_2488,N_2443);
xnor U2946 (N_2946,N_2674,N_2478);
nor U2947 (N_2947,N_2564,N_2433);
or U2948 (N_2948,N_2453,N_2486);
nand U2949 (N_2949,N_2612,N_2606);
and U2950 (N_2950,N_2664,N_2697);
nor U2951 (N_2951,N_2495,N_2502);
or U2952 (N_2952,N_2545,N_2662);
and U2953 (N_2953,N_2439,N_2570);
nand U2954 (N_2954,N_2446,N_2431);
or U2955 (N_2955,N_2631,N_2570);
xor U2956 (N_2956,N_2572,N_2476);
nor U2957 (N_2957,N_2578,N_2625);
nand U2958 (N_2958,N_2692,N_2549);
or U2959 (N_2959,N_2663,N_2599);
and U2960 (N_2960,N_2468,N_2585);
nand U2961 (N_2961,N_2453,N_2630);
nand U2962 (N_2962,N_2444,N_2403);
and U2963 (N_2963,N_2691,N_2576);
nor U2964 (N_2964,N_2575,N_2519);
nor U2965 (N_2965,N_2527,N_2521);
or U2966 (N_2966,N_2521,N_2616);
and U2967 (N_2967,N_2667,N_2617);
xnor U2968 (N_2968,N_2565,N_2509);
or U2969 (N_2969,N_2432,N_2411);
and U2970 (N_2970,N_2459,N_2486);
or U2971 (N_2971,N_2581,N_2485);
nor U2972 (N_2972,N_2490,N_2518);
xnor U2973 (N_2973,N_2674,N_2439);
xor U2974 (N_2974,N_2594,N_2663);
xnor U2975 (N_2975,N_2440,N_2477);
and U2976 (N_2976,N_2617,N_2599);
xor U2977 (N_2977,N_2481,N_2570);
xnor U2978 (N_2978,N_2581,N_2464);
nor U2979 (N_2979,N_2415,N_2549);
nand U2980 (N_2980,N_2472,N_2439);
xor U2981 (N_2981,N_2508,N_2557);
nor U2982 (N_2982,N_2451,N_2516);
or U2983 (N_2983,N_2617,N_2630);
xnor U2984 (N_2984,N_2590,N_2486);
and U2985 (N_2985,N_2693,N_2663);
nand U2986 (N_2986,N_2445,N_2428);
or U2987 (N_2987,N_2526,N_2543);
and U2988 (N_2988,N_2574,N_2527);
xnor U2989 (N_2989,N_2614,N_2679);
nand U2990 (N_2990,N_2518,N_2661);
xnor U2991 (N_2991,N_2576,N_2639);
or U2992 (N_2992,N_2632,N_2477);
nand U2993 (N_2993,N_2547,N_2596);
xor U2994 (N_2994,N_2563,N_2416);
and U2995 (N_2995,N_2601,N_2656);
nand U2996 (N_2996,N_2535,N_2498);
nand U2997 (N_2997,N_2505,N_2557);
nand U2998 (N_2998,N_2438,N_2671);
and U2999 (N_2999,N_2521,N_2617);
nand U3000 (N_3000,N_2847,N_2807);
nor U3001 (N_3001,N_2950,N_2990);
or U3002 (N_3002,N_2968,N_2984);
nor U3003 (N_3003,N_2930,N_2805);
xor U3004 (N_3004,N_2779,N_2709);
and U3005 (N_3005,N_2786,N_2795);
nor U3006 (N_3006,N_2980,N_2820);
xnor U3007 (N_3007,N_2725,N_2946);
xor U3008 (N_3008,N_2918,N_2977);
xnor U3009 (N_3009,N_2824,N_2745);
xor U3010 (N_3010,N_2874,N_2838);
and U3011 (N_3011,N_2762,N_2986);
and U3012 (N_3012,N_2922,N_2799);
nor U3013 (N_3013,N_2826,N_2700);
and U3014 (N_3014,N_2976,N_2815);
and U3015 (N_3015,N_2858,N_2731);
xnor U3016 (N_3016,N_2963,N_2706);
and U3017 (N_3017,N_2929,N_2956);
or U3018 (N_3018,N_2909,N_2836);
xnor U3019 (N_3019,N_2937,N_2942);
or U3020 (N_3020,N_2865,N_2734);
xnor U3021 (N_3021,N_2948,N_2943);
nor U3022 (N_3022,N_2926,N_2790);
and U3023 (N_3023,N_2778,N_2845);
or U3024 (N_3024,N_2832,N_2800);
or U3025 (N_3025,N_2787,N_2712);
nand U3026 (N_3026,N_2961,N_2710);
xnor U3027 (N_3027,N_2884,N_2707);
nor U3028 (N_3028,N_2705,N_2822);
or U3029 (N_3029,N_2857,N_2966);
nand U3030 (N_3030,N_2839,N_2877);
xnor U3031 (N_3031,N_2780,N_2866);
nand U3032 (N_3032,N_2987,N_2947);
xnor U3033 (N_3033,N_2830,N_2978);
or U3034 (N_3034,N_2856,N_2837);
nor U3035 (N_3035,N_2999,N_2843);
nand U3036 (N_3036,N_2788,N_2809);
and U3037 (N_3037,N_2776,N_2841);
or U3038 (N_3038,N_2952,N_2803);
xnor U3039 (N_3039,N_2798,N_2913);
nor U3040 (N_3040,N_2938,N_2738);
and U3041 (N_3041,N_2719,N_2796);
and U3042 (N_3042,N_2936,N_2821);
nor U3043 (N_3043,N_2997,N_2829);
or U3044 (N_3044,N_2993,N_2825);
nor U3045 (N_3045,N_2872,N_2804);
or U3046 (N_3046,N_2729,N_2876);
nor U3047 (N_3047,N_2982,N_2998);
and U3048 (N_3048,N_2765,N_2751);
xor U3049 (N_3049,N_2823,N_2891);
xor U3050 (N_3050,N_2873,N_2991);
or U3051 (N_3051,N_2958,N_2750);
or U3052 (N_3052,N_2960,N_2771);
or U3053 (N_3053,N_2813,N_2728);
nand U3054 (N_3054,N_2878,N_2708);
and U3055 (N_3055,N_2811,N_2890);
xor U3056 (N_3056,N_2717,N_2908);
xnor U3057 (N_3057,N_2896,N_2816);
xor U3058 (N_3058,N_2867,N_2868);
nand U3059 (N_3059,N_2899,N_2768);
nor U3060 (N_3060,N_2933,N_2785);
or U3061 (N_3061,N_2715,N_2921);
or U3062 (N_3062,N_2949,N_2885);
nand U3063 (N_3063,N_2880,N_2802);
nand U3064 (N_3064,N_2740,N_2840);
xnor U3065 (N_3065,N_2848,N_2774);
and U3066 (N_3066,N_2742,N_2975);
or U3067 (N_3067,N_2903,N_2923);
nand U3068 (N_3068,N_2741,N_2760);
and U3069 (N_3069,N_2905,N_2919);
nor U3070 (N_3070,N_2912,N_2863);
nor U3071 (N_3071,N_2844,N_2965);
xnor U3072 (N_3072,N_2941,N_2994);
or U3073 (N_3073,N_2931,N_2851);
and U3074 (N_3074,N_2988,N_2764);
and U3075 (N_3075,N_2748,N_2962);
or U3076 (N_3076,N_2894,N_2730);
xor U3077 (N_3077,N_2945,N_2792);
nand U3078 (N_3078,N_2833,N_2846);
xor U3079 (N_3079,N_2722,N_2985);
xor U3080 (N_3080,N_2781,N_2739);
xor U3081 (N_3081,N_2861,N_2871);
xor U3082 (N_3082,N_2951,N_2910);
and U3083 (N_3083,N_2889,N_2911);
xor U3084 (N_3084,N_2784,N_2892);
nand U3085 (N_3085,N_2972,N_2959);
or U3086 (N_3086,N_2814,N_2969);
nor U3087 (N_3087,N_2749,N_2902);
and U3088 (N_3088,N_2732,N_2860);
nor U3089 (N_3089,N_2720,N_2743);
nand U3090 (N_3090,N_2967,N_2835);
xor U3091 (N_3091,N_2763,N_2714);
and U3092 (N_3092,N_2723,N_2828);
or U3093 (N_3093,N_2995,N_2754);
or U3094 (N_3094,N_2907,N_2974);
or U3095 (N_3095,N_2897,N_2983);
and U3096 (N_3096,N_2701,N_2920);
nand U3097 (N_3097,N_2746,N_2756);
and U3098 (N_3098,N_2859,N_2870);
xnor U3099 (N_3099,N_2914,N_2834);
or U3100 (N_3100,N_2855,N_2989);
or U3101 (N_3101,N_2753,N_2953);
nor U3102 (N_3102,N_2758,N_2992);
nor U3103 (N_3103,N_2819,N_2721);
and U3104 (N_3104,N_2996,N_2932);
nor U3105 (N_3105,N_2726,N_2713);
or U3106 (N_3106,N_2883,N_2864);
or U3107 (N_3107,N_2971,N_2727);
xor U3108 (N_3108,N_2744,N_2973);
or U3109 (N_3109,N_2703,N_2917);
nor U3110 (N_3110,N_2702,N_2812);
nor U3111 (N_3111,N_2789,N_2827);
nand U3112 (N_3112,N_2769,N_2853);
nand U3113 (N_3113,N_2934,N_2793);
or U3114 (N_3114,N_2818,N_2900);
nor U3115 (N_3115,N_2737,N_2794);
nand U3116 (N_3116,N_2783,N_2752);
and U3117 (N_3117,N_2981,N_2964);
nor U3118 (N_3118,N_2782,N_2718);
nor U3119 (N_3119,N_2970,N_2736);
xnor U3120 (N_3120,N_2759,N_2879);
nand U3121 (N_3121,N_2770,N_2957);
xor U3122 (N_3122,N_2801,N_2940);
xnor U3123 (N_3123,N_2755,N_2772);
and U3124 (N_3124,N_2898,N_2927);
or U3125 (N_3125,N_2895,N_2906);
nand U3126 (N_3126,N_2817,N_2882);
and U3127 (N_3127,N_2854,N_2916);
nand U3128 (N_3128,N_2767,N_2761);
and U3129 (N_3129,N_2928,N_2797);
xnor U3130 (N_3130,N_2711,N_2831);
or U3131 (N_3131,N_2808,N_2886);
and U3132 (N_3132,N_2852,N_2904);
nand U3133 (N_3133,N_2810,N_2766);
and U3134 (N_3134,N_2775,N_2747);
and U3135 (N_3135,N_2925,N_2724);
nand U3136 (N_3136,N_2733,N_2849);
nor U3137 (N_3137,N_2979,N_2954);
nand U3138 (N_3138,N_2901,N_2704);
nand U3139 (N_3139,N_2915,N_2735);
or U3140 (N_3140,N_2888,N_2875);
or U3141 (N_3141,N_2777,N_2806);
nor U3142 (N_3142,N_2955,N_2773);
and U3143 (N_3143,N_2716,N_2757);
nor U3144 (N_3144,N_2939,N_2881);
and U3145 (N_3145,N_2869,N_2791);
or U3146 (N_3146,N_2924,N_2887);
and U3147 (N_3147,N_2850,N_2893);
nor U3148 (N_3148,N_2944,N_2935);
and U3149 (N_3149,N_2842,N_2862);
nor U3150 (N_3150,N_2701,N_2706);
nor U3151 (N_3151,N_2909,N_2954);
and U3152 (N_3152,N_2875,N_2871);
nand U3153 (N_3153,N_2807,N_2743);
nor U3154 (N_3154,N_2974,N_2915);
or U3155 (N_3155,N_2925,N_2748);
xnor U3156 (N_3156,N_2708,N_2890);
xor U3157 (N_3157,N_2846,N_2964);
or U3158 (N_3158,N_2855,N_2754);
nor U3159 (N_3159,N_2920,N_2962);
xnor U3160 (N_3160,N_2960,N_2903);
nor U3161 (N_3161,N_2864,N_2923);
nand U3162 (N_3162,N_2934,N_2859);
xor U3163 (N_3163,N_2752,N_2981);
nand U3164 (N_3164,N_2969,N_2986);
xor U3165 (N_3165,N_2773,N_2927);
or U3166 (N_3166,N_2955,N_2767);
xnor U3167 (N_3167,N_2847,N_2701);
xor U3168 (N_3168,N_2776,N_2983);
and U3169 (N_3169,N_2987,N_2874);
nand U3170 (N_3170,N_2875,N_2774);
xor U3171 (N_3171,N_2770,N_2990);
nand U3172 (N_3172,N_2977,N_2959);
and U3173 (N_3173,N_2974,N_2890);
or U3174 (N_3174,N_2790,N_2722);
or U3175 (N_3175,N_2859,N_2724);
nor U3176 (N_3176,N_2983,N_2885);
nor U3177 (N_3177,N_2791,N_2744);
or U3178 (N_3178,N_2835,N_2901);
and U3179 (N_3179,N_2894,N_2833);
nor U3180 (N_3180,N_2734,N_2832);
xor U3181 (N_3181,N_2863,N_2792);
xnor U3182 (N_3182,N_2748,N_2976);
nand U3183 (N_3183,N_2977,N_2759);
or U3184 (N_3184,N_2962,N_2958);
nor U3185 (N_3185,N_2710,N_2770);
nand U3186 (N_3186,N_2957,N_2954);
and U3187 (N_3187,N_2780,N_2755);
or U3188 (N_3188,N_2973,N_2923);
nor U3189 (N_3189,N_2950,N_2896);
xnor U3190 (N_3190,N_2792,N_2942);
xnor U3191 (N_3191,N_2850,N_2906);
and U3192 (N_3192,N_2831,N_2731);
xor U3193 (N_3193,N_2729,N_2836);
nand U3194 (N_3194,N_2744,N_2813);
xor U3195 (N_3195,N_2982,N_2942);
and U3196 (N_3196,N_2749,N_2949);
xnor U3197 (N_3197,N_2885,N_2904);
or U3198 (N_3198,N_2993,N_2988);
nor U3199 (N_3199,N_2753,N_2877);
and U3200 (N_3200,N_2707,N_2906);
nand U3201 (N_3201,N_2924,N_2951);
and U3202 (N_3202,N_2861,N_2832);
or U3203 (N_3203,N_2897,N_2819);
or U3204 (N_3204,N_2857,N_2886);
nor U3205 (N_3205,N_2708,N_2896);
xnor U3206 (N_3206,N_2949,N_2802);
and U3207 (N_3207,N_2860,N_2838);
nand U3208 (N_3208,N_2776,N_2911);
nor U3209 (N_3209,N_2795,N_2963);
xnor U3210 (N_3210,N_2939,N_2908);
nor U3211 (N_3211,N_2752,N_2768);
nand U3212 (N_3212,N_2965,N_2718);
nor U3213 (N_3213,N_2998,N_2799);
or U3214 (N_3214,N_2860,N_2881);
or U3215 (N_3215,N_2861,N_2727);
nand U3216 (N_3216,N_2810,N_2841);
xor U3217 (N_3217,N_2792,N_2790);
xor U3218 (N_3218,N_2863,N_2837);
nor U3219 (N_3219,N_2881,N_2795);
nand U3220 (N_3220,N_2716,N_2808);
nand U3221 (N_3221,N_2957,N_2729);
and U3222 (N_3222,N_2898,N_2779);
xor U3223 (N_3223,N_2979,N_2973);
or U3224 (N_3224,N_2889,N_2865);
xor U3225 (N_3225,N_2817,N_2993);
nand U3226 (N_3226,N_2706,N_2780);
nand U3227 (N_3227,N_2955,N_2740);
xor U3228 (N_3228,N_2734,N_2805);
or U3229 (N_3229,N_2794,N_2714);
or U3230 (N_3230,N_2870,N_2723);
and U3231 (N_3231,N_2789,N_2888);
or U3232 (N_3232,N_2764,N_2952);
xor U3233 (N_3233,N_2943,N_2751);
and U3234 (N_3234,N_2960,N_2833);
and U3235 (N_3235,N_2801,N_2751);
or U3236 (N_3236,N_2825,N_2763);
nor U3237 (N_3237,N_2910,N_2938);
nand U3238 (N_3238,N_2992,N_2740);
and U3239 (N_3239,N_2943,N_2863);
or U3240 (N_3240,N_2723,N_2913);
nand U3241 (N_3241,N_2821,N_2721);
nand U3242 (N_3242,N_2755,N_2852);
nand U3243 (N_3243,N_2961,N_2991);
and U3244 (N_3244,N_2808,N_2733);
and U3245 (N_3245,N_2819,N_2746);
nand U3246 (N_3246,N_2764,N_2702);
and U3247 (N_3247,N_2901,N_2967);
and U3248 (N_3248,N_2754,N_2874);
xnor U3249 (N_3249,N_2889,N_2713);
nand U3250 (N_3250,N_2939,N_2996);
xor U3251 (N_3251,N_2717,N_2875);
or U3252 (N_3252,N_2884,N_2986);
and U3253 (N_3253,N_2892,N_2823);
nor U3254 (N_3254,N_2867,N_2801);
and U3255 (N_3255,N_2971,N_2769);
or U3256 (N_3256,N_2707,N_2782);
or U3257 (N_3257,N_2772,N_2935);
and U3258 (N_3258,N_2965,N_2870);
or U3259 (N_3259,N_2989,N_2712);
or U3260 (N_3260,N_2850,N_2948);
and U3261 (N_3261,N_2828,N_2825);
or U3262 (N_3262,N_2809,N_2987);
nor U3263 (N_3263,N_2722,N_2769);
nor U3264 (N_3264,N_2909,N_2975);
nand U3265 (N_3265,N_2760,N_2730);
xnor U3266 (N_3266,N_2885,N_2850);
nand U3267 (N_3267,N_2761,N_2864);
or U3268 (N_3268,N_2956,N_2822);
nor U3269 (N_3269,N_2760,N_2824);
and U3270 (N_3270,N_2927,N_2984);
xor U3271 (N_3271,N_2864,N_2951);
xor U3272 (N_3272,N_2747,N_2945);
xnor U3273 (N_3273,N_2729,N_2981);
nand U3274 (N_3274,N_2811,N_2753);
nand U3275 (N_3275,N_2905,N_2917);
xnor U3276 (N_3276,N_2991,N_2715);
xnor U3277 (N_3277,N_2957,N_2838);
or U3278 (N_3278,N_2832,N_2799);
nand U3279 (N_3279,N_2855,N_2950);
nor U3280 (N_3280,N_2999,N_2951);
nor U3281 (N_3281,N_2919,N_2776);
and U3282 (N_3282,N_2954,N_2746);
and U3283 (N_3283,N_2859,N_2881);
nand U3284 (N_3284,N_2937,N_2747);
nand U3285 (N_3285,N_2840,N_2803);
nand U3286 (N_3286,N_2969,N_2935);
nand U3287 (N_3287,N_2794,N_2996);
nand U3288 (N_3288,N_2721,N_2966);
xnor U3289 (N_3289,N_2759,N_2929);
or U3290 (N_3290,N_2742,N_2974);
xnor U3291 (N_3291,N_2802,N_2983);
or U3292 (N_3292,N_2799,N_2794);
xnor U3293 (N_3293,N_2709,N_2784);
and U3294 (N_3294,N_2704,N_2874);
nand U3295 (N_3295,N_2823,N_2709);
nor U3296 (N_3296,N_2807,N_2923);
and U3297 (N_3297,N_2780,N_2967);
nand U3298 (N_3298,N_2802,N_2971);
or U3299 (N_3299,N_2814,N_2952);
xor U3300 (N_3300,N_3009,N_3024);
or U3301 (N_3301,N_3000,N_3166);
nand U3302 (N_3302,N_3163,N_3016);
nand U3303 (N_3303,N_3251,N_3122);
and U3304 (N_3304,N_3219,N_3136);
nand U3305 (N_3305,N_3228,N_3220);
and U3306 (N_3306,N_3098,N_3084);
xnor U3307 (N_3307,N_3225,N_3152);
xor U3308 (N_3308,N_3222,N_3049);
xor U3309 (N_3309,N_3202,N_3139);
and U3310 (N_3310,N_3297,N_3253);
xor U3311 (N_3311,N_3211,N_3204);
or U3312 (N_3312,N_3028,N_3217);
or U3313 (N_3313,N_3143,N_3153);
nor U3314 (N_3314,N_3106,N_3147);
xor U3315 (N_3315,N_3275,N_3276);
nor U3316 (N_3316,N_3118,N_3117);
or U3317 (N_3317,N_3190,N_3013);
nand U3318 (N_3318,N_3002,N_3103);
xor U3319 (N_3319,N_3281,N_3142);
or U3320 (N_3320,N_3296,N_3230);
nor U3321 (N_3321,N_3160,N_3114);
xor U3322 (N_3322,N_3283,N_3124);
and U3323 (N_3323,N_3191,N_3111);
or U3324 (N_3324,N_3027,N_3260);
nor U3325 (N_3325,N_3259,N_3074);
xnor U3326 (N_3326,N_3039,N_3145);
nand U3327 (N_3327,N_3177,N_3042);
nor U3328 (N_3328,N_3001,N_3258);
nor U3329 (N_3329,N_3216,N_3268);
xor U3330 (N_3330,N_3080,N_3026);
xnor U3331 (N_3331,N_3183,N_3223);
nor U3332 (N_3332,N_3244,N_3203);
and U3333 (N_3333,N_3113,N_3077);
nor U3334 (N_3334,N_3252,N_3261);
nand U3335 (N_3335,N_3286,N_3107);
nor U3336 (N_3336,N_3291,N_3178);
nand U3337 (N_3337,N_3115,N_3184);
xnor U3338 (N_3338,N_3198,N_3110);
xnor U3339 (N_3339,N_3087,N_3004);
and U3340 (N_3340,N_3227,N_3194);
nand U3341 (N_3341,N_3037,N_3130);
and U3342 (N_3342,N_3003,N_3018);
and U3343 (N_3343,N_3020,N_3277);
and U3344 (N_3344,N_3092,N_3287);
nand U3345 (N_3345,N_3012,N_3280);
and U3346 (N_3346,N_3066,N_3174);
or U3347 (N_3347,N_3047,N_3025);
and U3348 (N_3348,N_3085,N_3173);
nor U3349 (N_3349,N_3298,N_3165);
and U3350 (N_3350,N_3148,N_3046);
or U3351 (N_3351,N_3053,N_3059);
nor U3352 (N_3352,N_3062,N_3133);
and U3353 (N_3353,N_3040,N_3019);
nor U3354 (N_3354,N_3294,N_3180);
nor U3355 (N_3355,N_3068,N_3195);
nand U3356 (N_3356,N_3181,N_3104);
xnor U3357 (N_3357,N_3140,N_3093);
or U3358 (N_3358,N_3058,N_3167);
xor U3359 (N_3359,N_3127,N_3196);
or U3360 (N_3360,N_3015,N_3236);
nor U3361 (N_3361,N_3029,N_3238);
or U3362 (N_3362,N_3185,N_3200);
xnor U3363 (N_3363,N_3069,N_3237);
or U3364 (N_3364,N_3101,N_3060);
or U3365 (N_3365,N_3242,N_3155);
nor U3366 (N_3366,N_3299,N_3067);
xor U3367 (N_3367,N_3179,N_3096);
or U3368 (N_3368,N_3005,N_3064);
nor U3369 (N_3369,N_3097,N_3006);
xnor U3370 (N_3370,N_3109,N_3161);
nand U3371 (N_3371,N_3149,N_3288);
nand U3372 (N_3372,N_3150,N_3126);
or U3373 (N_3373,N_3156,N_3017);
and U3374 (N_3374,N_3116,N_3205);
nor U3375 (N_3375,N_3008,N_3246);
nand U3376 (N_3376,N_3076,N_3041);
or U3377 (N_3377,N_3055,N_3144);
xor U3378 (N_3378,N_3257,N_3090);
nand U3379 (N_3379,N_3129,N_3050);
nand U3380 (N_3380,N_3256,N_3121);
nand U3381 (N_3381,N_3197,N_3081);
or U3382 (N_3382,N_3250,N_3188);
nand U3383 (N_3383,N_3135,N_3295);
and U3384 (N_3384,N_3199,N_3154);
nor U3385 (N_3385,N_3033,N_3247);
or U3386 (N_3386,N_3293,N_3245);
nand U3387 (N_3387,N_3141,N_3065);
nor U3388 (N_3388,N_3078,N_3213);
and U3389 (N_3389,N_3207,N_3169);
and U3390 (N_3390,N_3137,N_3057);
nand U3391 (N_3391,N_3038,N_3285);
nand U3392 (N_3392,N_3239,N_3229);
xnor U3393 (N_3393,N_3171,N_3138);
nor U3394 (N_3394,N_3048,N_3157);
nor U3395 (N_3395,N_3262,N_3045);
or U3396 (N_3396,N_3070,N_3108);
or U3397 (N_3397,N_3176,N_3168);
or U3398 (N_3398,N_3254,N_3290);
nand U3399 (N_3399,N_3270,N_3051);
and U3400 (N_3400,N_3146,N_3233);
nor U3401 (N_3401,N_3273,N_3201);
and U3402 (N_3402,N_3241,N_3063);
or U3403 (N_3403,N_3075,N_3035);
or U3404 (N_3404,N_3030,N_3100);
nor U3405 (N_3405,N_3264,N_3132);
and U3406 (N_3406,N_3079,N_3011);
nor U3407 (N_3407,N_3243,N_3231);
nand U3408 (N_3408,N_3267,N_3218);
and U3409 (N_3409,N_3189,N_3105);
nand U3410 (N_3410,N_3182,N_3224);
or U3411 (N_3411,N_3172,N_3021);
and U3412 (N_3412,N_3091,N_3120);
or U3413 (N_3413,N_3263,N_3255);
or U3414 (N_3414,N_3014,N_3234);
xor U3415 (N_3415,N_3215,N_3272);
nand U3416 (N_3416,N_3099,N_3187);
or U3417 (N_3417,N_3134,N_3044);
nor U3418 (N_3418,N_3284,N_3056);
nand U3419 (N_3419,N_3054,N_3086);
or U3420 (N_3420,N_3061,N_3036);
or U3421 (N_3421,N_3289,N_3095);
nor U3422 (N_3422,N_3131,N_3279);
nor U3423 (N_3423,N_3265,N_3089);
and U3424 (N_3424,N_3072,N_3226);
xor U3425 (N_3425,N_3125,N_3162);
xnor U3426 (N_3426,N_3032,N_3266);
nor U3427 (N_3427,N_3240,N_3102);
xnor U3428 (N_3428,N_3034,N_3206);
nor U3429 (N_3429,N_3292,N_3007);
xnor U3430 (N_3430,N_3249,N_3128);
or U3431 (N_3431,N_3159,N_3186);
nor U3432 (N_3432,N_3209,N_3282);
and U3433 (N_3433,N_3192,N_3221);
xor U3434 (N_3434,N_3071,N_3271);
xnor U3435 (N_3435,N_3031,N_3119);
nand U3436 (N_3436,N_3170,N_3164);
or U3437 (N_3437,N_3083,N_3082);
or U3438 (N_3438,N_3088,N_3248);
xor U3439 (N_3439,N_3235,N_3043);
or U3440 (N_3440,N_3210,N_3214);
or U3441 (N_3441,N_3123,N_3151);
nor U3442 (N_3442,N_3010,N_3269);
nor U3443 (N_3443,N_3232,N_3094);
and U3444 (N_3444,N_3175,N_3212);
nand U3445 (N_3445,N_3193,N_3208);
or U3446 (N_3446,N_3158,N_3022);
nor U3447 (N_3447,N_3023,N_3052);
nor U3448 (N_3448,N_3278,N_3112);
xor U3449 (N_3449,N_3073,N_3274);
nor U3450 (N_3450,N_3148,N_3031);
and U3451 (N_3451,N_3096,N_3262);
nor U3452 (N_3452,N_3011,N_3199);
nand U3453 (N_3453,N_3215,N_3225);
and U3454 (N_3454,N_3289,N_3287);
nor U3455 (N_3455,N_3178,N_3262);
and U3456 (N_3456,N_3017,N_3006);
or U3457 (N_3457,N_3100,N_3000);
nor U3458 (N_3458,N_3263,N_3138);
or U3459 (N_3459,N_3131,N_3297);
and U3460 (N_3460,N_3161,N_3069);
xor U3461 (N_3461,N_3121,N_3266);
or U3462 (N_3462,N_3253,N_3262);
xnor U3463 (N_3463,N_3035,N_3033);
or U3464 (N_3464,N_3211,N_3252);
nand U3465 (N_3465,N_3087,N_3041);
nand U3466 (N_3466,N_3195,N_3039);
xor U3467 (N_3467,N_3125,N_3161);
xnor U3468 (N_3468,N_3133,N_3197);
nor U3469 (N_3469,N_3064,N_3083);
and U3470 (N_3470,N_3247,N_3067);
xnor U3471 (N_3471,N_3247,N_3244);
or U3472 (N_3472,N_3048,N_3149);
xor U3473 (N_3473,N_3120,N_3247);
nand U3474 (N_3474,N_3227,N_3273);
xnor U3475 (N_3475,N_3240,N_3283);
and U3476 (N_3476,N_3087,N_3188);
nor U3477 (N_3477,N_3086,N_3022);
xnor U3478 (N_3478,N_3137,N_3065);
or U3479 (N_3479,N_3208,N_3221);
nor U3480 (N_3480,N_3177,N_3194);
nand U3481 (N_3481,N_3020,N_3085);
nor U3482 (N_3482,N_3006,N_3050);
xor U3483 (N_3483,N_3260,N_3271);
or U3484 (N_3484,N_3039,N_3009);
xor U3485 (N_3485,N_3142,N_3173);
nor U3486 (N_3486,N_3251,N_3169);
nand U3487 (N_3487,N_3028,N_3155);
nor U3488 (N_3488,N_3023,N_3093);
and U3489 (N_3489,N_3083,N_3216);
xnor U3490 (N_3490,N_3003,N_3025);
and U3491 (N_3491,N_3264,N_3247);
nand U3492 (N_3492,N_3086,N_3170);
xor U3493 (N_3493,N_3203,N_3164);
nand U3494 (N_3494,N_3125,N_3071);
xnor U3495 (N_3495,N_3118,N_3160);
or U3496 (N_3496,N_3143,N_3122);
nor U3497 (N_3497,N_3127,N_3118);
nor U3498 (N_3498,N_3071,N_3035);
nand U3499 (N_3499,N_3017,N_3290);
and U3500 (N_3500,N_3008,N_3275);
nand U3501 (N_3501,N_3241,N_3054);
nor U3502 (N_3502,N_3291,N_3094);
and U3503 (N_3503,N_3028,N_3128);
and U3504 (N_3504,N_3144,N_3275);
and U3505 (N_3505,N_3238,N_3237);
xor U3506 (N_3506,N_3069,N_3156);
xor U3507 (N_3507,N_3174,N_3005);
nand U3508 (N_3508,N_3145,N_3215);
or U3509 (N_3509,N_3064,N_3197);
and U3510 (N_3510,N_3177,N_3195);
xor U3511 (N_3511,N_3108,N_3102);
nor U3512 (N_3512,N_3250,N_3040);
nand U3513 (N_3513,N_3169,N_3278);
and U3514 (N_3514,N_3054,N_3106);
xor U3515 (N_3515,N_3098,N_3220);
nor U3516 (N_3516,N_3166,N_3083);
nor U3517 (N_3517,N_3233,N_3059);
xnor U3518 (N_3518,N_3271,N_3228);
or U3519 (N_3519,N_3216,N_3154);
or U3520 (N_3520,N_3271,N_3092);
or U3521 (N_3521,N_3181,N_3168);
and U3522 (N_3522,N_3175,N_3150);
xor U3523 (N_3523,N_3253,N_3213);
xor U3524 (N_3524,N_3176,N_3227);
and U3525 (N_3525,N_3179,N_3204);
nor U3526 (N_3526,N_3263,N_3258);
nor U3527 (N_3527,N_3079,N_3001);
nand U3528 (N_3528,N_3293,N_3112);
nand U3529 (N_3529,N_3116,N_3102);
and U3530 (N_3530,N_3123,N_3110);
nor U3531 (N_3531,N_3118,N_3196);
or U3532 (N_3532,N_3066,N_3275);
or U3533 (N_3533,N_3071,N_3127);
xnor U3534 (N_3534,N_3285,N_3063);
and U3535 (N_3535,N_3105,N_3288);
nand U3536 (N_3536,N_3215,N_3104);
or U3537 (N_3537,N_3173,N_3281);
and U3538 (N_3538,N_3278,N_3060);
nand U3539 (N_3539,N_3215,N_3078);
or U3540 (N_3540,N_3016,N_3084);
nor U3541 (N_3541,N_3265,N_3136);
nand U3542 (N_3542,N_3074,N_3223);
and U3543 (N_3543,N_3227,N_3192);
or U3544 (N_3544,N_3105,N_3252);
and U3545 (N_3545,N_3004,N_3141);
xor U3546 (N_3546,N_3077,N_3008);
nand U3547 (N_3547,N_3284,N_3045);
and U3548 (N_3548,N_3084,N_3086);
nand U3549 (N_3549,N_3128,N_3237);
xnor U3550 (N_3550,N_3054,N_3071);
nor U3551 (N_3551,N_3199,N_3139);
or U3552 (N_3552,N_3018,N_3101);
and U3553 (N_3553,N_3106,N_3055);
and U3554 (N_3554,N_3172,N_3188);
nor U3555 (N_3555,N_3066,N_3259);
nor U3556 (N_3556,N_3152,N_3272);
nand U3557 (N_3557,N_3272,N_3146);
nand U3558 (N_3558,N_3074,N_3098);
xnor U3559 (N_3559,N_3031,N_3229);
or U3560 (N_3560,N_3293,N_3105);
nand U3561 (N_3561,N_3295,N_3080);
xor U3562 (N_3562,N_3053,N_3261);
xor U3563 (N_3563,N_3267,N_3216);
or U3564 (N_3564,N_3280,N_3192);
nand U3565 (N_3565,N_3158,N_3224);
nor U3566 (N_3566,N_3245,N_3023);
and U3567 (N_3567,N_3136,N_3152);
and U3568 (N_3568,N_3149,N_3045);
nand U3569 (N_3569,N_3041,N_3105);
nor U3570 (N_3570,N_3088,N_3030);
and U3571 (N_3571,N_3185,N_3230);
nand U3572 (N_3572,N_3101,N_3195);
and U3573 (N_3573,N_3202,N_3124);
and U3574 (N_3574,N_3021,N_3049);
xnor U3575 (N_3575,N_3067,N_3145);
or U3576 (N_3576,N_3081,N_3006);
or U3577 (N_3577,N_3257,N_3284);
xnor U3578 (N_3578,N_3196,N_3044);
nand U3579 (N_3579,N_3173,N_3157);
xor U3580 (N_3580,N_3026,N_3285);
or U3581 (N_3581,N_3244,N_3267);
and U3582 (N_3582,N_3101,N_3153);
or U3583 (N_3583,N_3184,N_3272);
nand U3584 (N_3584,N_3213,N_3095);
or U3585 (N_3585,N_3075,N_3173);
or U3586 (N_3586,N_3171,N_3169);
nor U3587 (N_3587,N_3191,N_3158);
or U3588 (N_3588,N_3076,N_3133);
xor U3589 (N_3589,N_3142,N_3245);
xor U3590 (N_3590,N_3011,N_3044);
or U3591 (N_3591,N_3126,N_3240);
or U3592 (N_3592,N_3155,N_3096);
and U3593 (N_3593,N_3000,N_3011);
xor U3594 (N_3594,N_3120,N_3011);
or U3595 (N_3595,N_3216,N_3208);
and U3596 (N_3596,N_3091,N_3280);
xnor U3597 (N_3597,N_3256,N_3199);
xnor U3598 (N_3598,N_3199,N_3075);
nor U3599 (N_3599,N_3114,N_3136);
nand U3600 (N_3600,N_3494,N_3520);
and U3601 (N_3601,N_3422,N_3343);
and U3602 (N_3602,N_3579,N_3478);
xor U3603 (N_3603,N_3593,N_3338);
and U3604 (N_3604,N_3370,N_3389);
nand U3605 (N_3605,N_3335,N_3590);
and U3606 (N_3606,N_3372,N_3591);
xnor U3607 (N_3607,N_3477,N_3391);
or U3608 (N_3608,N_3547,N_3313);
nand U3609 (N_3609,N_3421,N_3566);
and U3610 (N_3610,N_3560,N_3513);
or U3611 (N_3611,N_3401,N_3581);
or U3612 (N_3612,N_3525,N_3431);
or U3613 (N_3613,N_3497,N_3385);
or U3614 (N_3614,N_3527,N_3564);
or U3615 (N_3615,N_3426,N_3555);
or U3616 (N_3616,N_3532,N_3443);
and U3617 (N_3617,N_3577,N_3589);
xnor U3618 (N_3618,N_3363,N_3423);
or U3619 (N_3619,N_3432,N_3466);
nor U3620 (N_3620,N_3379,N_3378);
nor U3621 (N_3621,N_3514,N_3573);
xor U3622 (N_3622,N_3377,N_3530);
nand U3623 (N_3623,N_3320,N_3515);
and U3624 (N_3624,N_3462,N_3390);
xnor U3625 (N_3625,N_3471,N_3369);
nand U3626 (N_3626,N_3472,N_3481);
nor U3627 (N_3627,N_3449,N_3425);
xor U3628 (N_3628,N_3561,N_3460);
xnor U3629 (N_3629,N_3455,N_3428);
nand U3630 (N_3630,N_3578,N_3387);
or U3631 (N_3631,N_3339,N_3307);
nand U3632 (N_3632,N_3444,N_3588);
and U3633 (N_3633,N_3308,N_3550);
xor U3634 (N_3634,N_3465,N_3381);
and U3635 (N_3635,N_3475,N_3410);
nor U3636 (N_3636,N_3576,N_3479);
nor U3637 (N_3637,N_3340,N_3533);
xnor U3638 (N_3638,N_3345,N_3583);
or U3639 (N_3639,N_3540,N_3434);
nand U3640 (N_3640,N_3382,N_3341);
and U3641 (N_3641,N_3453,N_3556);
or U3642 (N_3642,N_3427,N_3498);
and U3643 (N_3643,N_3534,N_3388);
nor U3644 (N_3644,N_3473,N_3330);
nand U3645 (N_3645,N_3344,N_3480);
and U3646 (N_3646,N_3597,N_3580);
nor U3647 (N_3647,N_3539,N_3327);
nor U3648 (N_3648,N_3446,N_3463);
and U3649 (N_3649,N_3399,N_3417);
and U3650 (N_3650,N_3304,N_3439);
nand U3651 (N_3651,N_3476,N_3366);
xor U3652 (N_3652,N_3502,N_3456);
or U3653 (N_3653,N_3505,N_3524);
xor U3654 (N_3654,N_3300,N_3474);
nor U3655 (N_3655,N_3383,N_3450);
or U3656 (N_3656,N_3408,N_3324);
xor U3657 (N_3657,N_3375,N_3484);
nor U3658 (N_3658,N_3482,N_3565);
nand U3659 (N_3659,N_3436,N_3485);
nand U3660 (N_3660,N_3352,N_3569);
nand U3661 (N_3661,N_3404,N_3403);
and U3662 (N_3662,N_3325,N_3311);
or U3663 (N_3663,N_3356,N_3572);
nand U3664 (N_3664,N_3328,N_3337);
nand U3665 (N_3665,N_3364,N_3342);
nand U3666 (N_3666,N_3518,N_3458);
and U3667 (N_3667,N_3509,N_3402);
and U3668 (N_3668,N_3586,N_3575);
or U3669 (N_3669,N_3570,N_3568);
nand U3670 (N_3670,N_3412,N_3558);
nand U3671 (N_3671,N_3396,N_3430);
or U3672 (N_3672,N_3549,N_3470);
nand U3673 (N_3673,N_3414,N_3585);
nand U3674 (N_3674,N_3347,N_3506);
or U3675 (N_3675,N_3537,N_3467);
nand U3676 (N_3676,N_3316,N_3405);
nor U3677 (N_3677,N_3424,N_3321);
xnor U3678 (N_3678,N_3397,N_3409);
xnor U3679 (N_3679,N_3411,N_3329);
xor U3680 (N_3680,N_3309,N_3503);
xnor U3681 (N_3681,N_3571,N_3528);
nor U3682 (N_3682,N_3461,N_3454);
xor U3683 (N_3683,N_3457,N_3416);
and U3684 (N_3684,N_3319,N_3314);
or U3685 (N_3685,N_3542,N_3452);
nand U3686 (N_3686,N_3336,N_3357);
xnor U3687 (N_3687,N_3594,N_3406);
or U3688 (N_3688,N_3507,N_3362);
nand U3689 (N_3689,N_3333,N_3531);
xor U3690 (N_3690,N_3459,N_3490);
or U3691 (N_3691,N_3374,N_3551);
xnor U3692 (N_3692,N_3538,N_3371);
nor U3693 (N_3693,N_3504,N_3488);
nand U3694 (N_3694,N_3322,N_3492);
nand U3695 (N_3695,N_3511,N_3418);
or U3696 (N_3696,N_3315,N_3348);
and U3697 (N_3697,N_3440,N_3493);
and U3698 (N_3698,N_3361,N_3510);
nand U3699 (N_3699,N_3413,N_3301);
and U3700 (N_3700,N_3529,N_3451);
or U3701 (N_3701,N_3496,N_3419);
nand U3702 (N_3702,N_3415,N_3522);
xor U3703 (N_3703,N_3435,N_3574);
xor U3704 (N_3704,N_3365,N_3429);
nand U3705 (N_3705,N_3442,N_3305);
xnor U3706 (N_3706,N_3317,N_3351);
or U3707 (N_3707,N_3407,N_3582);
or U3708 (N_3708,N_3508,N_3554);
or U3709 (N_3709,N_3441,N_3541);
and U3710 (N_3710,N_3400,N_3310);
nand U3711 (N_3711,N_3584,N_3331);
and U3712 (N_3712,N_3326,N_3376);
nand U3713 (N_3713,N_3302,N_3398);
and U3714 (N_3714,N_3516,N_3536);
and U3715 (N_3715,N_3445,N_3367);
nor U3716 (N_3716,N_3448,N_3501);
nor U3717 (N_3717,N_3512,N_3354);
or U3718 (N_3718,N_3360,N_3433);
xor U3719 (N_3719,N_3567,N_3437);
nand U3720 (N_3720,N_3306,N_3386);
and U3721 (N_3721,N_3323,N_3350);
nand U3722 (N_3722,N_3546,N_3499);
nand U3723 (N_3723,N_3563,N_3447);
nor U3724 (N_3724,N_3517,N_3334);
or U3725 (N_3725,N_3303,N_3521);
or U3726 (N_3726,N_3373,N_3438);
nor U3727 (N_3727,N_3545,N_3349);
nor U3728 (N_3728,N_3393,N_3526);
xnor U3729 (N_3729,N_3519,N_3359);
nand U3730 (N_3730,N_3392,N_3487);
nor U3731 (N_3731,N_3312,N_3557);
and U3732 (N_3732,N_3535,N_3562);
xor U3733 (N_3733,N_3495,N_3353);
nor U3734 (N_3734,N_3500,N_3559);
nor U3735 (N_3735,N_3358,N_3368);
xnor U3736 (N_3736,N_3592,N_3332);
or U3737 (N_3737,N_3491,N_3394);
and U3738 (N_3738,N_3596,N_3552);
xor U3739 (N_3739,N_3483,N_3489);
or U3740 (N_3740,N_3464,N_3523);
nand U3741 (N_3741,N_3384,N_3355);
nand U3742 (N_3742,N_3469,N_3395);
xor U3743 (N_3743,N_3468,N_3486);
nor U3744 (N_3744,N_3598,N_3346);
xor U3745 (N_3745,N_3553,N_3420);
nor U3746 (N_3746,N_3599,N_3380);
nand U3747 (N_3747,N_3548,N_3318);
nor U3748 (N_3748,N_3543,N_3544);
nand U3749 (N_3749,N_3595,N_3587);
nor U3750 (N_3750,N_3440,N_3444);
nand U3751 (N_3751,N_3592,N_3459);
and U3752 (N_3752,N_3445,N_3300);
nand U3753 (N_3753,N_3545,N_3372);
and U3754 (N_3754,N_3396,N_3581);
xor U3755 (N_3755,N_3406,N_3553);
nand U3756 (N_3756,N_3480,N_3582);
nor U3757 (N_3757,N_3445,N_3541);
nor U3758 (N_3758,N_3309,N_3527);
or U3759 (N_3759,N_3582,N_3440);
or U3760 (N_3760,N_3537,N_3503);
xnor U3761 (N_3761,N_3498,N_3478);
and U3762 (N_3762,N_3555,N_3498);
xnor U3763 (N_3763,N_3445,N_3303);
and U3764 (N_3764,N_3329,N_3354);
or U3765 (N_3765,N_3512,N_3532);
nor U3766 (N_3766,N_3474,N_3412);
or U3767 (N_3767,N_3586,N_3500);
or U3768 (N_3768,N_3397,N_3510);
xnor U3769 (N_3769,N_3440,N_3320);
xor U3770 (N_3770,N_3401,N_3344);
and U3771 (N_3771,N_3444,N_3313);
nor U3772 (N_3772,N_3547,N_3311);
nor U3773 (N_3773,N_3595,N_3308);
and U3774 (N_3774,N_3491,N_3318);
and U3775 (N_3775,N_3312,N_3439);
and U3776 (N_3776,N_3485,N_3315);
or U3777 (N_3777,N_3329,N_3422);
and U3778 (N_3778,N_3490,N_3307);
nor U3779 (N_3779,N_3411,N_3403);
and U3780 (N_3780,N_3551,N_3588);
nand U3781 (N_3781,N_3422,N_3390);
or U3782 (N_3782,N_3538,N_3321);
nand U3783 (N_3783,N_3306,N_3354);
or U3784 (N_3784,N_3510,N_3381);
nand U3785 (N_3785,N_3377,N_3413);
or U3786 (N_3786,N_3464,N_3454);
or U3787 (N_3787,N_3416,N_3314);
and U3788 (N_3788,N_3576,N_3350);
or U3789 (N_3789,N_3414,N_3566);
nor U3790 (N_3790,N_3436,N_3357);
nand U3791 (N_3791,N_3548,N_3541);
nand U3792 (N_3792,N_3583,N_3511);
xnor U3793 (N_3793,N_3543,N_3337);
nand U3794 (N_3794,N_3317,N_3371);
or U3795 (N_3795,N_3509,N_3464);
and U3796 (N_3796,N_3463,N_3400);
or U3797 (N_3797,N_3322,N_3487);
nor U3798 (N_3798,N_3536,N_3337);
and U3799 (N_3799,N_3337,N_3390);
nor U3800 (N_3800,N_3556,N_3515);
xnor U3801 (N_3801,N_3460,N_3328);
xnor U3802 (N_3802,N_3517,N_3321);
xor U3803 (N_3803,N_3490,N_3338);
nor U3804 (N_3804,N_3576,N_3585);
or U3805 (N_3805,N_3400,N_3458);
xor U3806 (N_3806,N_3579,N_3477);
or U3807 (N_3807,N_3338,N_3462);
and U3808 (N_3808,N_3440,N_3306);
or U3809 (N_3809,N_3340,N_3514);
xnor U3810 (N_3810,N_3524,N_3336);
or U3811 (N_3811,N_3563,N_3586);
nand U3812 (N_3812,N_3539,N_3385);
and U3813 (N_3813,N_3577,N_3393);
nor U3814 (N_3814,N_3460,N_3597);
nand U3815 (N_3815,N_3524,N_3334);
xor U3816 (N_3816,N_3585,N_3549);
nand U3817 (N_3817,N_3428,N_3460);
xor U3818 (N_3818,N_3531,N_3563);
nand U3819 (N_3819,N_3553,N_3529);
or U3820 (N_3820,N_3434,N_3303);
or U3821 (N_3821,N_3444,N_3327);
nand U3822 (N_3822,N_3402,N_3574);
nor U3823 (N_3823,N_3408,N_3436);
xnor U3824 (N_3824,N_3505,N_3545);
nor U3825 (N_3825,N_3496,N_3591);
xor U3826 (N_3826,N_3323,N_3401);
or U3827 (N_3827,N_3435,N_3475);
and U3828 (N_3828,N_3302,N_3416);
nor U3829 (N_3829,N_3313,N_3591);
or U3830 (N_3830,N_3368,N_3300);
xnor U3831 (N_3831,N_3489,N_3372);
or U3832 (N_3832,N_3450,N_3486);
nand U3833 (N_3833,N_3469,N_3586);
and U3834 (N_3834,N_3491,N_3362);
nor U3835 (N_3835,N_3408,N_3396);
and U3836 (N_3836,N_3489,N_3362);
xnor U3837 (N_3837,N_3595,N_3437);
and U3838 (N_3838,N_3324,N_3423);
nand U3839 (N_3839,N_3372,N_3470);
nor U3840 (N_3840,N_3572,N_3543);
nor U3841 (N_3841,N_3536,N_3392);
xnor U3842 (N_3842,N_3361,N_3437);
xor U3843 (N_3843,N_3316,N_3330);
nand U3844 (N_3844,N_3333,N_3522);
or U3845 (N_3845,N_3433,N_3311);
and U3846 (N_3846,N_3326,N_3559);
or U3847 (N_3847,N_3594,N_3547);
nor U3848 (N_3848,N_3432,N_3594);
xor U3849 (N_3849,N_3549,N_3392);
and U3850 (N_3850,N_3343,N_3541);
nor U3851 (N_3851,N_3407,N_3529);
or U3852 (N_3852,N_3474,N_3347);
or U3853 (N_3853,N_3304,N_3380);
nand U3854 (N_3854,N_3571,N_3584);
and U3855 (N_3855,N_3591,N_3479);
xor U3856 (N_3856,N_3303,N_3372);
nand U3857 (N_3857,N_3583,N_3405);
or U3858 (N_3858,N_3457,N_3528);
xnor U3859 (N_3859,N_3512,N_3421);
nor U3860 (N_3860,N_3576,N_3332);
xor U3861 (N_3861,N_3433,N_3407);
nor U3862 (N_3862,N_3369,N_3373);
nand U3863 (N_3863,N_3397,N_3573);
or U3864 (N_3864,N_3519,N_3477);
nand U3865 (N_3865,N_3309,N_3512);
nor U3866 (N_3866,N_3411,N_3425);
nand U3867 (N_3867,N_3446,N_3453);
nor U3868 (N_3868,N_3399,N_3342);
nor U3869 (N_3869,N_3455,N_3452);
xnor U3870 (N_3870,N_3393,N_3402);
and U3871 (N_3871,N_3417,N_3554);
or U3872 (N_3872,N_3340,N_3456);
or U3873 (N_3873,N_3551,N_3379);
nand U3874 (N_3874,N_3311,N_3358);
or U3875 (N_3875,N_3417,N_3513);
nand U3876 (N_3876,N_3501,N_3401);
nand U3877 (N_3877,N_3325,N_3508);
xor U3878 (N_3878,N_3411,N_3432);
nor U3879 (N_3879,N_3419,N_3500);
xor U3880 (N_3880,N_3383,N_3392);
nor U3881 (N_3881,N_3421,N_3484);
or U3882 (N_3882,N_3375,N_3518);
and U3883 (N_3883,N_3418,N_3525);
xor U3884 (N_3884,N_3466,N_3496);
or U3885 (N_3885,N_3334,N_3390);
xnor U3886 (N_3886,N_3370,N_3549);
or U3887 (N_3887,N_3402,N_3533);
xor U3888 (N_3888,N_3402,N_3598);
nand U3889 (N_3889,N_3330,N_3368);
nor U3890 (N_3890,N_3387,N_3358);
and U3891 (N_3891,N_3567,N_3590);
and U3892 (N_3892,N_3321,N_3479);
or U3893 (N_3893,N_3379,N_3525);
and U3894 (N_3894,N_3459,N_3457);
xor U3895 (N_3895,N_3341,N_3481);
xor U3896 (N_3896,N_3336,N_3469);
or U3897 (N_3897,N_3582,N_3439);
nand U3898 (N_3898,N_3356,N_3477);
or U3899 (N_3899,N_3579,N_3448);
nand U3900 (N_3900,N_3813,N_3661);
nor U3901 (N_3901,N_3642,N_3764);
or U3902 (N_3902,N_3768,N_3864);
nand U3903 (N_3903,N_3629,N_3613);
nor U3904 (N_3904,N_3710,N_3848);
xnor U3905 (N_3905,N_3638,N_3670);
and U3906 (N_3906,N_3627,N_3677);
and U3907 (N_3907,N_3798,N_3622);
nor U3908 (N_3908,N_3636,N_3749);
xnor U3909 (N_3909,N_3787,N_3603);
nor U3910 (N_3910,N_3635,N_3759);
or U3911 (N_3911,N_3832,N_3879);
xnor U3912 (N_3912,N_3608,N_3857);
nand U3913 (N_3913,N_3872,N_3658);
or U3914 (N_3914,N_3789,N_3646);
and U3915 (N_3915,N_3688,N_3895);
or U3916 (N_3916,N_3678,N_3890);
nand U3917 (N_3917,N_3632,N_3831);
nor U3918 (N_3918,N_3656,N_3793);
nand U3919 (N_3919,N_3682,N_3711);
and U3920 (N_3920,N_3626,N_3833);
and U3921 (N_3921,N_3610,N_3891);
and U3922 (N_3922,N_3862,N_3617);
and U3923 (N_3923,N_3756,N_3845);
or U3924 (N_3924,N_3628,N_3820);
nand U3925 (N_3925,N_3790,N_3795);
xnor U3926 (N_3926,N_3648,N_3738);
nand U3927 (N_3927,N_3676,N_3691);
nand U3928 (N_3928,N_3666,N_3619);
xor U3929 (N_3929,N_3722,N_3814);
nand U3930 (N_3930,N_3762,N_3777);
nor U3931 (N_3931,N_3750,N_3887);
nor U3932 (N_3932,N_3866,N_3884);
nor U3933 (N_3933,N_3611,N_3624);
or U3934 (N_3934,N_3746,N_3708);
or U3935 (N_3935,N_3853,N_3838);
nor U3936 (N_3936,N_3870,N_3659);
nor U3937 (N_3937,N_3671,N_3729);
and U3938 (N_3938,N_3614,N_3788);
and U3939 (N_3939,N_3769,N_3669);
xnor U3940 (N_3940,N_3747,N_3655);
or U3941 (N_3941,N_3782,N_3732);
xor U3942 (N_3942,N_3804,N_3826);
nor U3943 (N_3943,N_3728,N_3612);
nor U3944 (N_3944,N_3821,N_3690);
nand U3945 (N_3945,N_3753,N_3720);
xnor U3946 (N_3946,N_3886,N_3835);
and U3947 (N_3947,N_3637,N_3745);
xor U3948 (N_3948,N_3640,N_3686);
and U3949 (N_3949,N_3776,N_3773);
xnor U3950 (N_3950,N_3606,N_3707);
nand U3951 (N_3951,N_3727,N_3885);
or U3952 (N_3952,N_3644,N_3693);
nor U3953 (N_3953,N_3701,N_3819);
nor U3954 (N_3954,N_3761,N_3868);
nor U3955 (N_3955,N_3726,N_3616);
nor U3956 (N_3956,N_3844,N_3781);
and U3957 (N_3957,N_3816,N_3704);
or U3958 (N_3958,N_3755,N_3631);
and U3959 (N_3959,N_3660,N_3639);
xnor U3960 (N_3960,N_3700,N_3687);
nor U3961 (N_3961,N_3775,N_3695);
xor U3962 (N_3962,N_3874,N_3730);
nor U3963 (N_3963,N_3852,N_3675);
and U3964 (N_3964,N_3892,N_3800);
nand U3965 (N_3965,N_3736,N_3683);
nor U3966 (N_3966,N_3758,N_3633);
nand U3967 (N_3967,N_3829,N_3618);
nor U3968 (N_3968,N_3815,N_3713);
or U3969 (N_3969,N_3880,N_3641);
xor U3970 (N_3970,N_3662,N_3876);
xnor U3971 (N_3971,N_3873,N_3602);
and U3972 (N_3972,N_3698,N_3609);
nand U3973 (N_3973,N_3794,N_3651);
or U3974 (N_3974,N_3785,N_3825);
and U3975 (N_3975,N_3812,N_3881);
and U3976 (N_3976,N_3858,N_3767);
or U3977 (N_3977,N_3652,N_3634);
or U3978 (N_3978,N_3799,N_3672);
or U3979 (N_3979,N_3893,N_3664);
xor U3980 (N_3980,N_3889,N_3780);
xor U3981 (N_3981,N_3654,N_3860);
or U3982 (N_3982,N_3807,N_3801);
and U3983 (N_3983,N_3869,N_3696);
nor U3984 (N_3984,N_3620,N_3742);
xor U3985 (N_3985,N_3605,N_3630);
xnor U3986 (N_3986,N_3843,N_3607);
or U3987 (N_3987,N_3875,N_3706);
nand U3988 (N_3988,N_3859,N_3604);
nand U3989 (N_3989,N_3667,N_3718);
xnor U3990 (N_3990,N_3725,N_3601);
nor U3991 (N_3991,N_3770,N_3863);
and U3992 (N_3992,N_3754,N_3673);
and U3993 (N_3993,N_3846,N_3830);
nand U3994 (N_3994,N_3663,N_3822);
nor U3995 (N_3995,N_3806,N_3811);
or U3996 (N_3996,N_3809,N_3600);
nor U3997 (N_3997,N_3842,N_3802);
and U3998 (N_3998,N_3680,N_3810);
or U3999 (N_3999,N_3847,N_3737);
nand U4000 (N_4000,N_3694,N_3739);
or U4001 (N_4001,N_3836,N_3766);
nand U4002 (N_4002,N_3703,N_3724);
xnor U4003 (N_4003,N_3784,N_3837);
nand U4004 (N_4004,N_3740,N_3861);
nor U4005 (N_4005,N_3897,N_3883);
xnor U4006 (N_4006,N_3625,N_3796);
nand U4007 (N_4007,N_3685,N_3772);
or U4008 (N_4008,N_3763,N_3689);
or U4009 (N_4009,N_3733,N_3615);
or U4010 (N_4010,N_3854,N_3679);
xnor U4011 (N_4011,N_3834,N_3856);
nor U4012 (N_4012,N_3741,N_3898);
or U4013 (N_4013,N_3878,N_3851);
and U4014 (N_4014,N_3734,N_3839);
and U4015 (N_4015,N_3896,N_3643);
nor U4016 (N_4016,N_3850,N_3668);
or U4017 (N_4017,N_3681,N_3716);
and U4018 (N_4018,N_3645,N_3827);
nand U4019 (N_4019,N_3748,N_3849);
nor U4020 (N_4020,N_3649,N_3817);
xnor U4021 (N_4021,N_3867,N_3744);
or U4022 (N_4022,N_3712,N_3808);
nand U4023 (N_4023,N_3692,N_3714);
and U4024 (N_4024,N_3778,N_3882);
nand U4025 (N_4025,N_3805,N_3697);
and U4026 (N_4026,N_3786,N_3877);
or U4027 (N_4027,N_3865,N_3871);
nor U4028 (N_4028,N_3894,N_3824);
nor U4029 (N_4029,N_3751,N_3647);
xnor U4030 (N_4030,N_3840,N_3650);
and U4031 (N_4031,N_3828,N_3705);
and U4032 (N_4032,N_3702,N_3899);
nand U4033 (N_4033,N_3757,N_3783);
nand U4034 (N_4034,N_3719,N_3653);
nand U4035 (N_4035,N_3735,N_3888);
nor U4036 (N_4036,N_3855,N_3743);
or U4037 (N_4037,N_3723,N_3774);
or U4038 (N_4038,N_3792,N_3731);
or U4039 (N_4039,N_3841,N_3623);
nand U4040 (N_4040,N_3699,N_3721);
xnor U4041 (N_4041,N_3803,N_3823);
nor U4042 (N_4042,N_3818,N_3797);
xnor U4043 (N_4043,N_3791,N_3779);
xnor U4044 (N_4044,N_3765,N_3621);
or U4045 (N_4045,N_3771,N_3684);
or U4046 (N_4046,N_3709,N_3715);
or U4047 (N_4047,N_3752,N_3657);
or U4048 (N_4048,N_3674,N_3717);
xnor U4049 (N_4049,N_3760,N_3665);
and U4050 (N_4050,N_3695,N_3799);
xor U4051 (N_4051,N_3812,N_3884);
nor U4052 (N_4052,N_3844,N_3829);
nand U4053 (N_4053,N_3835,N_3840);
nor U4054 (N_4054,N_3838,N_3820);
or U4055 (N_4055,N_3634,N_3854);
nor U4056 (N_4056,N_3697,N_3655);
or U4057 (N_4057,N_3819,N_3863);
or U4058 (N_4058,N_3845,N_3748);
nor U4059 (N_4059,N_3775,N_3663);
or U4060 (N_4060,N_3703,N_3816);
xor U4061 (N_4061,N_3872,N_3826);
xor U4062 (N_4062,N_3750,N_3650);
xnor U4063 (N_4063,N_3626,N_3868);
and U4064 (N_4064,N_3724,N_3758);
nand U4065 (N_4065,N_3797,N_3753);
xnor U4066 (N_4066,N_3806,N_3787);
and U4067 (N_4067,N_3866,N_3602);
nor U4068 (N_4068,N_3668,N_3809);
xnor U4069 (N_4069,N_3785,N_3783);
nor U4070 (N_4070,N_3603,N_3841);
or U4071 (N_4071,N_3871,N_3647);
nand U4072 (N_4072,N_3776,N_3834);
or U4073 (N_4073,N_3695,N_3814);
nand U4074 (N_4074,N_3740,N_3634);
or U4075 (N_4075,N_3858,N_3692);
nand U4076 (N_4076,N_3715,N_3714);
or U4077 (N_4077,N_3855,N_3878);
nand U4078 (N_4078,N_3781,N_3811);
nand U4079 (N_4079,N_3812,N_3723);
nor U4080 (N_4080,N_3681,N_3658);
or U4081 (N_4081,N_3703,N_3698);
xor U4082 (N_4082,N_3717,N_3692);
nor U4083 (N_4083,N_3853,N_3806);
xnor U4084 (N_4084,N_3721,N_3656);
and U4085 (N_4085,N_3842,N_3654);
nand U4086 (N_4086,N_3600,N_3761);
and U4087 (N_4087,N_3787,N_3656);
and U4088 (N_4088,N_3716,N_3621);
or U4089 (N_4089,N_3823,N_3816);
or U4090 (N_4090,N_3782,N_3873);
nor U4091 (N_4091,N_3857,N_3708);
or U4092 (N_4092,N_3718,N_3626);
nor U4093 (N_4093,N_3693,N_3625);
nand U4094 (N_4094,N_3785,N_3738);
nor U4095 (N_4095,N_3679,N_3771);
xor U4096 (N_4096,N_3851,N_3611);
xor U4097 (N_4097,N_3889,N_3724);
xnor U4098 (N_4098,N_3782,N_3843);
or U4099 (N_4099,N_3782,N_3854);
or U4100 (N_4100,N_3694,N_3836);
nand U4101 (N_4101,N_3601,N_3721);
nor U4102 (N_4102,N_3672,N_3811);
and U4103 (N_4103,N_3737,N_3835);
or U4104 (N_4104,N_3758,N_3778);
nand U4105 (N_4105,N_3710,N_3613);
nand U4106 (N_4106,N_3633,N_3624);
and U4107 (N_4107,N_3835,N_3848);
nand U4108 (N_4108,N_3791,N_3897);
and U4109 (N_4109,N_3795,N_3639);
nor U4110 (N_4110,N_3893,N_3853);
nand U4111 (N_4111,N_3828,N_3868);
nor U4112 (N_4112,N_3663,N_3675);
nand U4113 (N_4113,N_3747,N_3741);
nand U4114 (N_4114,N_3677,N_3705);
nand U4115 (N_4115,N_3777,N_3821);
nand U4116 (N_4116,N_3669,N_3820);
xor U4117 (N_4117,N_3875,N_3634);
or U4118 (N_4118,N_3795,N_3673);
or U4119 (N_4119,N_3657,N_3728);
or U4120 (N_4120,N_3601,N_3664);
and U4121 (N_4121,N_3736,N_3647);
nand U4122 (N_4122,N_3872,N_3862);
nor U4123 (N_4123,N_3797,N_3871);
xor U4124 (N_4124,N_3653,N_3635);
nor U4125 (N_4125,N_3744,N_3747);
and U4126 (N_4126,N_3631,N_3884);
xnor U4127 (N_4127,N_3856,N_3641);
nor U4128 (N_4128,N_3743,N_3812);
xor U4129 (N_4129,N_3610,N_3770);
nand U4130 (N_4130,N_3856,N_3774);
or U4131 (N_4131,N_3704,N_3794);
and U4132 (N_4132,N_3766,N_3762);
nor U4133 (N_4133,N_3765,N_3856);
nand U4134 (N_4134,N_3635,N_3697);
or U4135 (N_4135,N_3871,N_3600);
or U4136 (N_4136,N_3757,N_3691);
nor U4137 (N_4137,N_3897,N_3739);
xnor U4138 (N_4138,N_3800,N_3815);
xnor U4139 (N_4139,N_3630,N_3794);
xor U4140 (N_4140,N_3696,N_3629);
nor U4141 (N_4141,N_3860,N_3870);
and U4142 (N_4142,N_3734,N_3745);
nand U4143 (N_4143,N_3796,N_3604);
xor U4144 (N_4144,N_3749,N_3656);
nand U4145 (N_4145,N_3669,N_3632);
and U4146 (N_4146,N_3605,N_3704);
and U4147 (N_4147,N_3693,N_3852);
xor U4148 (N_4148,N_3693,N_3626);
nand U4149 (N_4149,N_3700,N_3750);
and U4150 (N_4150,N_3746,N_3626);
nand U4151 (N_4151,N_3744,N_3808);
nand U4152 (N_4152,N_3603,N_3602);
nand U4153 (N_4153,N_3827,N_3796);
or U4154 (N_4154,N_3796,N_3757);
and U4155 (N_4155,N_3660,N_3839);
and U4156 (N_4156,N_3895,N_3741);
and U4157 (N_4157,N_3875,N_3835);
xor U4158 (N_4158,N_3680,N_3754);
or U4159 (N_4159,N_3650,N_3734);
nor U4160 (N_4160,N_3742,N_3628);
nand U4161 (N_4161,N_3750,N_3623);
and U4162 (N_4162,N_3808,N_3896);
xor U4163 (N_4163,N_3636,N_3858);
xnor U4164 (N_4164,N_3864,N_3744);
and U4165 (N_4165,N_3730,N_3794);
and U4166 (N_4166,N_3857,N_3770);
xor U4167 (N_4167,N_3803,N_3689);
nor U4168 (N_4168,N_3874,N_3799);
and U4169 (N_4169,N_3619,N_3650);
nor U4170 (N_4170,N_3747,N_3688);
nor U4171 (N_4171,N_3777,N_3801);
nand U4172 (N_4172,N_3713,N_3790);
and U4173 (N_4173,N_3797,N_3621);
nor U4174 (N_4174,N_3658,N_3831);
or U4175 (N_4175,N_3645,N_3734);
nand U4176 (N_4176,N_3782,N_3866);
or U4177 (N_4177,N_3794,N_3762);
nor U4178 (N_4178,N_3821,N_3710);
xor U4179 (N_4179,N_3760,N_3601);
nor U4180 (N_4180,N_3694,N_3644);
and U4181 (N_4181,N_3601,N_3864);
nor U4182 (N_4182,N_3801,N_3853);
nand U4183 (N_4183,N_3732,N_3707);
or U4184 (N_4184,N_3761,N_3627);
xnor U4185 (N_4185,N_3628,N_3666);
xnor U4186 (N_4186,N_3806,N_3763);
or U4187 (N_4187,N_3882,N_3898);
and U4188 (N_4188,N_3828,N_3752);
nor U4189 (N_4189,N_3628,N_3836);
xor U4190 (N_4190,N_3835,N_3820);
xnor U4191 (N_4191,N_3647,N_3791);
xnor U4192 (N_4192,N_3835,N_3885);
and U4193 (N_4193,N_3775,N_3621);
or U4194 (N_4194,N_3689,N_3753);
nand U4195 (N_4195,N_3890,N_3746);
xnor U4196 (N_4196,N_3835,N_3892);
or U4197 (N_4197,N_3623,N_3866);
nand U4198 (N_4198,N_3783,N_3812);
and U4199 (N_4199,N_3732,N_3777);
or U4200 (N_4200,N_3967,N_4096);
nor U4201 (N_4201,N_3921,N_4023);
xnor U4202 (N_4202,N_4127,N_3934);
xnor U4203 (N_4203,N_4042,N_4006);
nand U4204 (N_4204,N_4155,N_3994);
nor U4205 (N_4205,N_4116,N_4074);
nor U4206 (N_4206,N_3902,N_4114);
nand U4207 (N_4207,N_4095,N_4022);
xnor U4208 (N_4208,N_4109,N_3963);
and U4209 (N_4209,N_4036,N_4170);
or U4210 (N_4210,N_4012,N_4041);
and U4211 (N_4211,N_4164,N_4083);
xnor U4212 (N_4212,N_4001,N_4134);
or U4213 (N_4213,N_3952,N_4058);
xor U4214 (N_4214,N_3936,N_4043);
nand U4215 (N_4215,N_4004,N_4141);
xor U4216 (N_4216,N_3907,N_3944);
or U4217 (N_4217,N_3983,N_4091);
nand U4218 (N_4218,N_4077,N_4026);
and U4219 (N_4219,N_3964,N_4173);
or U4220 (N_4220,N_4171,N_3953);
and U4221 (N_4221,N_4158,N_3935);
and U4222 (N_4222,N_4092,N_4069);
xnor U4223 (N_4223,N_3969,N_3979);
nand U4224 (N_4224,N_3943,N_3937);
nor U4225 (N_4225,N_3916,N_4197);
nand U4226 (N_4226,N_3957,N_4190);
nand U4227 (N_4227,N_4169,N_4038);
nor U4228 (N_4228,N_4107,N_4048);
and U4229 (N_4229,N_3974,N_4059);
or U4230 (N_4230,N_4143,N_4099);
xnor U4231 (N_4231,N_4049,N_4102);
nand U4232 (N_4232,N_4000,N_4184);
and U4233 (N_4233,N_4100,N_4024);
nor U4234 (N_4234,N_4124,N_3993);
nor U4235 (N_4235,N_4054,N_4185);
nor U4236 (N_4236,N_4090,N_3932);
or U4237 (N_4237,N_4167,N_4113);
xor U4238 (N_4238,N_3999,N_4084);
nand U4239 (N_4239,N_4050,N_4097);
or U4240 (N_4240,N_4039,N_4125);
xor U4241 (N_4241,N_3947,N_3978);
xnor U4242 (N_4242,N_4017,N_4192);
xor U4243 (N_4243,N_3903,N_3991);
nor U4244 (N_4244,N_4014,N_4176);
nor U4245 (N_4245,N_3939,N_4052);
nor U4246 (N_4246,N_4101,N_4019);
and U4247 (N_4247,N_3985,N_3931);
nand U4248 (N_4248,N_4007,N_4168);
nand U4249 (N_4249,N_4159,N_4104);
and U4250 (N_4250,N_3954,N_4189);
nor U4251 (N_4251,N_4162,N_4132);
and U4252 (N_4252,N_3990,N_3960);
nand U4253 (N_4253,N_4029,N_4073);
xor U4254 (N_4254,N_3904,N_4191);
and U4255 (N_4255,N_4016,N_3927);
or U4256 (N_4256,N_4053,N_4064);
and U4257 (N_4257,N_3901,N_3971);
or U4258 (N_4258,N_3988,N_3913);
xor U4259 (N_4259,N_4030,N_3946);
nand U4260 (N_4260,N_4149,N_4133);
xor U4261 (N_4261,N_3919,N_4117);
and U4262 (N_4262,N_4089,N_4070);
nand U4263 (N_4263,N_3980,N_3926);
nand U4264 (N_4264,N_3912,N_4122);
nand U4265 (N_4265,N_4151,N_4130);
and U4266 (N_4266,N_3970,N_4055);
nor U4267 (N_4267,N_4172,N_4156);
nor U4268 (N_4268,N_4182,N_4121);
or U4269 (N_4269,N_3924,N_4140);
or U4270 (N_4270,N_3949,N_4137);
xnor U4271 (N_4271,N_4015,N_3911);
nand U4272 (N_4272,N_3996,N_4161);
and U4273 (N_4273,N_3925,N_3928);
and U4274 (N_4274,N_3975,N_4174);
nand U4275 (N_4275,N_3917,N_4098);
nor U4276 (N_4276,N_4166,N_4136);
nor U4277 (N_4277,N_3909,N_4163);
or U4278 (N_4278,N_4106,N_4087);
nand U4279 (N_4279,N_4119,N_3973);
nor U4280 (N_4280,N_4123,N_3920);
nor U4281 (N_4281,N_4034,N_4131);
or U4282 (N_4282,N_4021,N_3976);
or U4283 (N_4283,N_4111,N_4148);
nor U4284 (N_4284,N_4088,N_3956);
or U4285 (N_4285,N_4018,N_4080);
nand U4286 (N_4286,N_3987,N_3992);
nand U4287 (N_4287,N_3945,N_4085);
nand U4288 (N_4288,N_3961,N_4196);
nor U4289 (N_4289,N_4175,N_4093);
and U4290 (N_4290,N_4033,N_4027);
xor U4291 (N_4291,N_4005,N_3972);
nand U4292 (N_4292,N_3959,N_4110);
xnor U4293 (N_4293,N_4179,N_4198);
xnor U4294 (N_4294,N_3968,N_4195);
and U4295 (N_4295,N_4081,N_4150);
and U4296 (N_4296,N_4051,N_4188);
and U4297 (N_4297,N_4037,N_4068);
nand U4298 (N_4298,N_4177,N_4115);
nor U4299 (N_4299,N_4160,N_4146);
or U4300 (N_4300,N_3915,N_3929);
nand U4301 (N_4301,N_4186,N_4011);
or U4302 (N_4302,N_4046,N_3905);
nor U4303 (N_4303,N_4028,N_4010);
and U4304 (N_4304,N_4067,N_4056);
or U4305 (N_4305,N_4082,N_4076);
and U4306 (N_4306,N_3998,N_3906);
and U4307 (N_4307,N_3938,N_4057);
and U4308 (N_4308,N_4199,N_4181);
xnor U4309 (N_4309,N_4144,N_4013);
nand U4310 (N_4310,N_4032,N_4060);
and U4311 (N_4311,N_4129,N_4066);
and U4312 (N_4312,N_3914,N_3923);
xnor U4313 (N_4313,N_4079,N_3951);
or U4314 (N_4314,N_4065,N_4062);
xor U4315 (N_4315,N_4126,N_3962);
xor U4316 (N_4316,N_4105,N_4047);
nand U4317 (N_4317,N_4139,N_4120);
or U4318 (N_4318,N_3955,N_3986);
xor U4319 (N_4319,N_4135,N_4154);
and U4320 (N_4320,N_3940,N_4086);
or U4321 (N_4321,N_3984,N_4193);
and U4322 (N_4322,N_4075,N_3965);
and U4323 (N_4323,N_4187,N_4180);
xnor U4324 (N_4324,N_4044,N_3948);
or U4325 (N_4325,N_3958,N_4145);
xor U4326 (N_4326,N_4071,N_3950);
or U4327 (N_4327,N_4009,N_4142);
nand U4328 (N_4328,N_4094,N_3910);
xor U4329 (N_4329,N_3966,N_4072);
and U4330 (N_4330,N_4153,N_3941);
and U4331 (N_4331,N_3942,N_4035);
or U4332 (N_4332,N_4002,N_3922);
xor U4333 (N_4333,N_4157,N_4147);
or U4334 (N_4334,N_3930,N_3977);
or U4335 (N_4335,N_4040,N_4118);
or U4336 (N_4336,N_4103,N_3908);
and U4337 (N_4337,N_4025,N_4020);
nor U4338 (N_4338,N_4003,N_4128);
nand U4339 (N_4339,N_3933,N_4045);
nand U4340 (N_4340,N_4031,N_4138);
nor U4341 (N_4341,N_3918,N_3997);
nor U4342 (N_4342,N_4061,N_4165);
xnor U4343 (N_4343,N_4078,N_4063);
xor U4344 (N_4344,N_3981,N_4008);
nor U4345 (N_4345,N_3900,N_4183);
xor U4346 (N_4346,N_4178,N_4108);
and U4347 (N_4347,N_4112,N_3989);
xor U4348 (N_4348,N_4194,N_3982);
and U4349 (N_4349,N_4152,N_3995);
nand U4350 (N_4350,N_4012,N_4017);
or U4351 (N_4351,N_4010,N_3910);
or U4352 (N_4352,N_4029,N_4036);
and U4353 (N_4353,N_4198,N_4114);
nor U4354 (N_4354,N_3932,N_3963);
nand U4355 (N_4355,N_4101,N_3914);
nand U4356 (N_4356,N_3961,N_3988);
xnor U4357 (N_4357,N_3927,N_4070);
and U4358 (N_4358,N_4132,N_4042);
or U4359 (N_4359,N_4128,N_4130);
or U4360 (N_4360,N_4124,N_3954);
nand U4361 (N_4361,N_3960,N_4121);
nor U4362 (N_4362,N_4086,N_4025);
nor U4363 (N_4363,N_3911,N_3913);
or U4364 (N_4364,N_3955,N_3950);
nand U4365 (N_4365,N_3998,N_4007);
nor U4366 (N_4366,N_4004,N_4172);
or U4367 (N_4367,N_4000,N_3989);
or U4368 (N_4368,N_3930,N_4060);
or U4369 (N_4369,N_3984,N_3965);
nand U4370 (N_4370,N_4078,N_4124);
or U4371 (N_4371,N_3944,N_4098);
and U4372 (N_4372,N_3963,N_3966);
nand U4373 (N_4373,N_4112,N_4064);
and U4374 (N_4374,N_4105,N_3905);
nand U4375 (N_4375,N_4188,N_3906);
nand U4376 (N_4376,N_4057,N_3925);
nand U4377 (N_4377,N_4177,N_4061);
or U4378 (N_4378,N_3975,N_3927);
or U4379 (N_4379,N_4033,N_4188);
xor U4380 (N_4380,N_4056,N_4057);
nand U4381 (N_4381,N_4125,N_4106);
nor U4382 (N_4382,N_4038,N_4098);
nand U4383 (N_4383,N_3940,N_4119);
nand U4384 (N_4384,N_4169,N_4172);
nor U4385 (N_4385,N_3939,N_3915);
nor U4386 (N_4386,N_4131,N_3924);
nor U4387 (N_4387,N_3989,N_4070);
nor U4388 (N_4388,N_4003,N_4123);
and U4389 (N_4389,N_4022,N_4155);
xnor U4390 (N_4390,N_3931,N_3957);
and U4391 (N_4391,N_4183,N_4120);
or U4392 (N_4392,N_4046,N_4080);
xor U4393 (N_4393,N_4021,N_3934);
or U4394 (N_4394,N_3956,N_4006);
and U4395 (N_4395,N_4111,N_3960);
xor U4396 (N_4396,N_4038,N_3909);
xor U4397 (N_4397,N_4101,N_4187);
nor U4398 (N_4398,N_3959,N_4165);
and U4399 (N_4399,N_4114,N_4016);
nor U4400 (N_4400,N_3967,N_3958);
and U4401 (N_4401,N_3931,N_4174);
nand U4402 (N_4402,N_3914,N_4021);
nand U4403 (N_4403,N_4162,N_4185);
and U4404 (N_4404,N_4169,N_4167);
nand U4405 (N_4405,N_4016,N_4001);
or U4406 (N_4406,N_3922,N_3923);
xnor U4407 (N_4407,N_3915,N_3903);
or U4408 (N_4408,N_4006,N_3925);
xor U4409 (N_4409,N_4103,N_4135);
nand U4410 (N_4410,N_4065,N_4172);
or U4411 (N_4411,N_3951,N_4040);
and U4412 (N_4412,N_3923,N_3945);
nor U4413 (N_4413,N_3953,N_3934);
and U4414 (N_4414,N_4071,N_3921);
nor U4415 (N_4415,N_4096,N_4009);
nor U4416 (N_4416,N_4150,N_3951);
nor U4417 (N_4417,N_4124,N_4051);
and U4418 (N_4418,N_4067,N_4131);
nor U4419 (N_4419,N_3906,N_3920);
nor U4420 (N_4420,N_4171,N_3954);
xor U4421 (N_4421,N_4097,N_4087);
nand U4422 (N_4422,N_4035,N_4008);
or U4423 (N_4423,N_4193,N_3999);
nand U4424 (N_4424,N_4196,N_4097);
nand U4425 (N_4425,N_3974,N_3935);
or U4426 (N_4426,N_4017,N_4188);
nand U4427 (N_4427,N_4104,N_4197);
xnor U4428 (N_4428,N_4171,N_4085);
and U4429 (N_4429,N_4021,N_4137);
xor U4430 (N_4430,N_3992,N_3909);
nor U4431 (N_4431,N_4013,N_4004);
xor U4432 (N_4432,N_3994,N_3971);
xnor U4433 (N_4433,N_4157,N_4050);
nand U4434 (N_4434,N_4029,N_3901);
nand U4435 (N_4435,N_4072,N_4086);
xnor U4436 (N_4436,N_4024,N_3911);
and U4437 (N_4437,N_3921,N_3996);
and U4438 (N_4438,N_4092,N_4174);
nor U4439 (N_4439,N_3938,N_3939);
nor U4440 (N_4440,N_4083,N_4059);
and U4441 (N_4441,N_4085,N_4087);
xnor U4442 (N_4442,N_3963,N_3905);
nor U4443 (N_4443,N_4019,N_4108);
or U4444 (N_4444,N_4120,N_3943);
nand U4445 (N_4445,N_4074,N_4018);
nand U4446 (N_4446,N_4145,N_3953);
nor U4447 (N_4447,N_3934,N_4118);
nand U4448 (N_4448,N_3969,N_4148);
or U4449 (N_4449,N_3936,N_4175);
nand U4450 (N_4450,N_3941,N_3948);
and U4451 (N_4451,N_4192,N_3973);
nand U4452 (N_4452,N_4000,N_4084);
nor U4453 (N_4453,N_4015,N_3971);
xnor U4454 (N_4454,N_4192,N_4123);
and U4455 (N_4455,N_3964,N_3989);
nor U4456 (N_4456,N_4087,N_4111);
xnor U4457 (N_4457,N_4105,N_4154);
nand U4458 (N_4458,N_4172,N_3911);
and U4459 (N_4459,N_4150,N_4172);
nor U4460 (N_4460,N_4140,N_4125);
and U4461 (N_4461,N_4087,N_4046);
nor U4462 (N_4462,N_3952,N_4054);
nor U4463 (N_4463,N_4052,N_3969);
and U4464 (N_4464,N_3901,N_4057);
nand U4465 (N_4465,N_4051,N_3948);
or U4466 (N_4466,N_4198,N_4135);
xor U4467 (N_4467,N_3902,N_4008);
nor U4468 (N_4468,N_4190,N_4095);
nor U4469 (N_4469,N_4167,N_4175);
or U4470 (N_4470,N_4195,N_3914);
nor U4471 (N_4471,N_3981,N_4090);
and U4472 (N_4472,N_4093,N_4185);
nor U4473 (N_4473,N_4111,N_4091);
and U4474 (N_4474,N_4012,N_4010);
and U4475 (N_4475,N_4041,N_4161);
xnor U4476 (N_4476,N_3902,N_4141);
and U4477 (N_4477,N_4133,N_4138);
xnor U4478 (N_4478,N_4086,N_3979);
nor U4479 (N_4479,N_4162,N_4106);
or U4480 (N_4480,N_4195,N_4012);
or U4481 (N_4481,N_4045,N_3903);
and U4482 (N_4482,N_3955,N_3975);
xnor U4483 (N_4483,N_3911,N_4083);
and U4484 (N_4484,N_4049,N_4192);
and U4485 (N_4485,N_3974,N_4128);
nor U4486 (N_4486,N_4018,N_4136);
nor U4487 (N_4487,N_3956,N_4014);
and U4488 (N_4488,N_4104,N_4002);
nor U4489 (N_4489,N_4180,N_4039);
nor U4490 (N_4490,N_4031,N_4027);
xnor U4491 (N_4491,N_4092,N_4196);
nor U4492 (N_4492,N_3956,N_4145);
or U4493 (N_4493,N_4050,N_4098);
or U4494 (N_4494,N_3990,N_4166);
and U4495 (N_4495,N_3953,N_4104);
nor U4496 (N_4496,N_4195,N_4123);
xnor U4497 (N_4497,N_4055,N_4190);
or U4498 (N_4498,N_4051,N_4163);
or U4499 (N_4499,N_4084,N_4190);
xnor U4500 (N_4500,N_4410,N_4346);
xnor U4501 (N_4501,N_4318,N_4235);
nand U4502 (N_4502,N_4280,N_4276);
xnor U4503 (N_4503,N_4489,N_4224);
nor U4504 (N_4504,N_4422,N_4454);
nor U4505 (N_4505,N_4494,N_4286);
nor U4506 (N_4506,N_4369,N_4474);
or U4507 (N_4507,N_4433,N_4309);
or U4508 (N_4508,N_4336,N_4365);
and U4509 (N_4509,N_4353,N_4428);
and U4510 (N_4510,N_4371,N_4442);
nand U4511 (N_4511,N_4348,N_4443);
and U4512 (N_4512,N_4388,N_4403);
and U4513 (N_4513,N_4421,N_4273);
nor U4514 (N_4514,N_4229,N_4269);
or U4515 (N_4515,N_4383,N_4225);
or U4516 (N_4516,N_4393,N_4206);
nor U4517 (N_4517,N_4375,N_4387);
and U4518 (N_4518,N_4304,N_4331);
xnor U4519 (N_4519,N_4244,N_4475);
nand U4520 (N_4520,N_4426,N_4352);
or U4521 (N_4521,N_4354,N_4482);
nor U4522 (N_4522,N_4469,N_4347);
nor U4523 (N_4523,N_4342,N_4262);
nor U4524 (N_4524,N_4481,N_4314);
nor U4525 (N_4525,N_4201,N_4243);
and U4526 (N_4526,N_4408,N_4351);
xnor U4527 (N_4527,N_4302,N_4332);
or U4528 (N_4528,N_4333,N_4356);
xor U4529 (N_4529,N_4226,N_4278);
nand U4530 (N_4530,N_4233,N_4487);
xnor U4531 (N_4531,N_4258,N_4259);
and U4532 (N_4532,N_4435,N_4452);
nand U4533 (N_4533,N_4294,N_4247);
or U4534 (N_4534,N_4207,N_4495);
xnor U4535 (N_4535,N_4219,N_4218);
nand U4536 (N_4536,N_4239,N_4432);
or U4537 (N_4537,N_4330,N_4293);
nor U4538 (N_4538,N_4400,N_4252);
nand U4539 (N_4539,N_4215,N_4251);
and U4540 (N_4540,N_4287,N_4405);
nor U4541 (N_4541,N_4412,N_4493);
or U4542 (N_4542,N_4463,N_4484);
xnor U4543 (N_4543,N_4476,N_4312);
and U4544 (N_4544,N_4277,N_4498);
or U4545 (N_4545,N_4456,N_4288);
and U4546 (N_4546,N_4217,N_4291);
or U4547 (N_4547,N_4292,N_4289);
or U4548 (N_4548,N_4439,N_4389);
xor U4549 (N_4549,N_4234,N_4246);
nor U4550 (N_4550,N_4430,N_4395);
xor U4551 (N_4551,N_4397,N_4458);
xor U4552 (N_4552,N_4460,N_4431);
and U4553 (N_4553,N_4253,N_4488);
nor U4554 (N_4554,N_4416,N_4324);
or U4555 (N_4555,N_4473,N_4265);
and U4556 (N_4556,N_4222,N_4268);
and U4557 (N_4557,N_4241,N_4228);
xor U4558 (N_4558,N_4419,N_4462);
or U4559 (N_4559,N_4376,N_4470);
or U4560 (N_4560,N_4447,N_4394);
nand U4561 (N_4561,N_4212,N_4308);
or U4562 (N_4562,N_4305,N_4295);
nor U4563 (N_4563,N_4425,N_4396);
and U4564 (N_4564,N_4231,N_4338);
nor U4565 (N_4565,N_4402,N_4471);
xnor U4566 (N_4566,N_4209,N_4372);
nor U4567 (N_4567,N_4380,N_4451);
nand U4568 (N_4568,N_4260,N_4378);
xnor U4569 (N_4569,N_4464,N_4491);
and U4570 (N_4570,N_4370,N_4381);
nand U4571 (N_4571,N_4423,N_4264);
xor U4572 (N_4572,N_4414,N_4275);
nand U4573 (N_4573,N_4361,N_4202);
xor U4574 (N_4574,N_4216,N_4325);
xnor U4575 (N_4575,N_4240,N_4407);
and U4576 (N_4576,N_4497,N_4359);
nand U4577 (N_4577,N_4398,N_4210);
nor U4578 (N_4578,N_4329,N_4320);
nor U4579 (N_4579,N_4284,N_4364);
or U4580 (N_4580,N_4281,N_4413);
or U4581 (N_4581,N_4390,N_4467);
or U4582 (N_4582,N_4249,N_4335);
xor U4583 (N_4583,N_4257,N_4386);
or U4584 (N_4584,N_4344,N_4440);
nand U4585 (N_4585,N_4434,N_4411);
nand U4586 (N_4586,N_4349,N_4261);
nand U4587 (N_4587,N_4340,N_4418);
nor U4588 (N_4588,N_4271,N_4437);
or U4589 (N_4589,N_4366,N_4367);
xor U4590 (N_4590,N_4382,N_4254);
nor U4591 (N_4591,N_4230,N_4444);
and U4592 (N_4592,N_4242,N_4450);
xor U4593 (N_4593,N_4420,N_4360);
and U4594 (N_4594,N_4377,N_4399);
and U4595 (N_4595,N_4424,N_4345);
and U4596 (N_4596,N_4499,N_4221);
or U4597 (N_4597,N_4483,N_4427);
nor U4598 (N_4598,N_4448,N_4256);
and U4599 (N_4599,N_4379,N_4313);
xnor U4600 (N_4600,N_4266,N_4350);
or U4601 (N_4601,N_4391,N_4203);
xor U4602 (N_4602,N_4323,N_4373);
nor U4603 (N_4603,N_4208,N_4339);
nand U4604 (N_4604,N_4417,N_4446);
xor U4605 (N_4605,N_4457,N_4328);
and U4606 (N_4606,N_4401,N_4415);
or U4607 (N_4607,N_4274,N_4449);
xnor U4608 (N_4608,N_4200,N_4409);
xnor U4609 (N_4609,N_4213,N_4404);
or U4610 (N_4610,N_4283,N_4272);
nor U4611 (N_4611,N_4429,N_4285);
xor U4612 (N_4612,N_4468,N_4465);
xor U4613 (N_4613,N_4214,N_4459);
nand U4614 (N_4614,N_4461,N_4327);
nor U4615 (N_4615,N_4374,N_4343);
nand U4616 (N_4616,N_4301,N_4445);
nand U4617 (N_4617,N_4438,N_4472);
nor U4618 (N_4618,N_4300,N_4279);
and U4619 (N_4619,N_4392,N_4306);
nand U4620 (N_4620,N_4322,N_4267);
or U4621 (N_4621,N_4238,N_4490);
xor U4622 (N_4622,N_4492,N_4236);
or U4623 (N_4623,N_4321,N_4357);
xor U4624 (N_4624,N_4303,N_4436);
xor U4625 (N_4625,N_4310,N_4385);
and U4626 (N_4626,N_4319,N_4455);
xor U4627 (N_4627,N_4248,N_4316);
xnor U4628 (N_4628,N_4307,N_4311);
nand U4629 (N_4629,N_4223,N_4315);
and U4630 (N_4630,N_4466,N_4479);
xor U4631 (N_4631,N_4290,N_4296);
nor U4632 (N_4632,N_4297,N_4270);
nand U4633 (N_4633,N_4245,N_4480);
or U4634 (N_4634,N_4477,N_4237);
and U4635 (N_4635,N_4232,N_4317);
and U4636 (N_4636,N_4362,N_4255);
and U4637 (N_4637,N_4298,N_4441);
or U4638 (N_4638,N_4358,N_4496);
nor U4639 (N_4639,N_4406,N_4250);
xnor U4640 (N_4640,N_4453,N_4485);
nor U4641 (N_4641,N_4326,N_4334);
or U4642 (N_4642,N_4299,N_4355);
xnor U4643 (N_4643,N_4337,N_4478);
nor U4644 (N_4644,N_4205,N_4211);
and U4645 (N_4645,N_4363,N_4227);
xnor U4646 (N_4646,N_4384,N_4282);
nor U4647 (N_4647,N_4368,N_4204);
xnor U4648 (N_4648,N_4341,N_4263);
nand U4649 (N_4649,N_4220,N_4486);
nor U4650 (N_4650,N_4417,N_4200);
xnor U4651 (N_4651,N_4279,N_4231);
or U4652 (N_4652,N_4416,N_4299);
xor U4653 (N_4653,N_4315,N_4476);
nand U4654 (N_4654,N_4429,N_4497);
nand U4655 (N_4655,N_4450,N_4436);
and U4656 (N_4656,N_4388,N_4365);
nand U4657 (N_4657,N_4318,N_4360);
nand U4658 (N_4658,N_4379,N_4310);
and U4659 (N_4659,N_4201,N_4372);
xor U4660 (N_4660,N_4490,N_4365);
xnor U4661 (N_4661,N_4422,N_4232);
nor U4662 (N_4662,N_4333,N_4271);
and U4663 (N_4663,N_4435,N_4333);
xor U4664 (N_4664,N_4396,N_4449);
or U4665 (N_4665,N_4470,N_4472);
xor U4666 (N_4666,N_4293,N_4458);
nor U4667 (N_4667,N_4397,N_4381);
nand U4668 (N_4668,N_4274,N_4289);
xnor U4669 (N_4669,N_4480,N_4232);
nand U4670 (N_4670,N_4294,N_4365);
or U4671 (N_4671,N_4473,N_4231);
and U4672 (N_4672,N_4461,N_4206);
nand U4673 (N_4673,N_4346,N_4389);
and U4674 (N_4674,N_4264,N_4252);
or U4675 (N_4675,N_4369,N_4344);
nor U4676 (N_4676,N_4233,N_4410);
xor U4677 (N_4677,N_4479,N_4477);
and U4678 (N_4678,N_4390,N_4466);
xnor U4679 (N_4679,N_4388,N_4474);
nand U4680 (N_4680,N_4458,N_4302);
nand U4681 (N_4681,N_4265,N_4315);
and U4682 (N_4682,N_4356,N_4431);
or U4683 (N_4683,N_4204,N_4348);
nor U4684 (N_4684,N_4400,N_4211);
nand U4685 (N_4685,N_4307,N_4434);
and U4686 (N_4686,N_4217,N_4303);
xor U4687 (N_4687,N_4329,N_4283);
nand U4688 (N_4688,N_4299,N_4407);
nor U4689 (N_4689,N_4375,N_4481);
and U4690 (N_4690,N_4497,N_4344);
nor U4691 (N_4691,N_4457,N_4347);
nor U4692 (N_4692,N_4368,N_4441);
nand U4693 (N_4693,N_4342,N_4315);
or U4694 (N_4694,N_4481,N_4308);
nand U4695 (N_4695,N_4300,N_4354);
xor U4696 (N_4696,N_4435,N_4466);
nand U4697 (N_4697,N_4472,N_4294);
xnor U4698 (N_4698,N_4296,N_4246);
xor U4699 (N_4699,N_4342,N_4326);
xnor U4700 (N_4700,N_4476,N_4459);
xor U4701 (N_4701,N_4383,N_4449);
and U4702 (N_4702,N_4449,N_4259);
and U4703 (N_4703,N_4397,N_4216);
and U4704 (N_4704,N_4459,N_4470);
nand U4705 (N_4705,N_4221,N_4484);
or U4706 (N_4706,N_4296,N_4219);
or U4707 (N_4707,N_4217,N_4486);
and U4708 (N_4708,N_4339,N_4460);
and U4709 (N_4709,N_4285,N_4356);
and U4710 (N_4710,N_4230,N_4250);
and U4711 (N_4711,N_4245,N_4290);
nor U4712 (N_4712,N_4230,N_4345);
xor U4713 (N_4713,N_4324,N_4221);
and U4714 (N_4714,N_4383,N_4386);
xor U4715 (N_4715,N_4308,N_4404);
and U4716 (N_4716,N_4278,N_4358);
nor U4717 (N_4717,N_4313,N_4341);
xor U4718 (N_4718,N_4486,N_4211);
nor U4719 (N_4719,N_4424,N_4217);
nor U4720 (N_4720,N_4368,N_4210);
nand U4721 (N_4721,N_4376,N_4408);
nand U4722 (N_4722,N_4386,N_4336);
xnor U4723 (N_4723,N_4200,N_4379);
or U4724 (N_4724,N_4235,N_4417);
nand U4725 (N_4725,N_4417,N_4398);
xnor U4726 (N_4726,N_4413,N_4483);
nor U4727 (N_4727,N_4428,N_4351);
nor U4728 (N_4728,N_4233,N_4286);
and U4729 (N_4729,N_4262,N_4479);
and U4730 (N_4730,N_4319,N_4422);
xor U4731 (N_4731,N_4338,N_4445);
xor U4732 (N_4732,N_4288,N_4242);
and U4733 (N_4733,N_4218,N_4463);
or U4734 (N_4734,N_4348,N_4219);
nor U4735 (N_4735,N_4459,N_4488);
xnor U4736 (N_4736,N_4363,N_4404);
and U4737 (N_4737,N_4265,N_4241);
or U4738 (N_4738,N_4422,N_4381);
or U4739 (N_4739,N_4350,N_4285);
nor U4740 (N_4740,N_4346,N_4495);
nor U4741 (N_4741,N_4248,N_4331);
nand U4742 (N_4742,N_4388,N_4438);
nand U4743 (N_4743,N_4480,N_4425);
xor U4744 (N_4744,N_4397,N_4432);
nor U4745 (N_4745,N_4242,N_4477);
xor U4746 (N_4746,N_4421,N_4321);
or U4747 (N_4747,N_4303,N_4237);
nor U4748 (N_4748,N_4231,N_4491);
nand U4749 (N_4749,N_4387,N_4271);
nand U4750 (N_4750,N_4323,N_4355);
and U4751 (N_4751,N_4424,N_4383);
and U4752 (N_4752,N_4269,N_4285);
and U4753 (N_4753,N_4383,N_4415);
nor U4754 (N_4754,N_4413,N_4472);
nor U4755 (N_4755,N_4491,N_4333);
and U4756 (N_4756,N_4478,N_4395);
nand U4757 (N_4757,N_4375,N_4293);
and U4758 (N_4758,N_4379,N_4284);
nand U4759 (N_4759,N_4438,N_4313);
or U4760 (N_4760,N_4224,N_4380);
xnor U4761 (N_4761,N_4465,N_4214);
xor U4762 (N_4762,N_4478,N_4287);
and U4763 (N_4763,N_4466,N_4384);
or U4764 (N_4764,N_4204,N_4352);
and U4765 (N_4765,N_4263,N_4277);
nand U4766 (N_4766,N_4443,N_4450);
xor U4767 (N_4767,N_4437,N_4293);
xor U4768 (N_4768,N_4454,N_4234);
nor U4769 (N_4769,N_4344,N_4351);
xor U4770 (N_4770,N_4260,N_4356);
or U4771 (N_4771,N_4291,N_4485);
and U4772 (N_4772,N_4416,N_4372);
or U4773 (N_4773,N_4211,N_4312);
xnor U4774 (N_4774,N_4480,N_4319);
xnor U4775 (N_4775,N_4276,N_4227);
nand U4776 (N_4776,N_4458,N_4367);
or U4777 (N_4777,N_4272,N_4401);
nand U4778 (N_4778,N_4265,N_4482);
or U4779 (N_4779,N_4364,N_4331);
xor U4780 (N_4780,N_4270,N_4312);
or U4781 (N_4781,N_4365,N_4376);
nor U4782 (N_4782,N_4495,N_4230);
nand U4783 (N_4783,N_4418,N_4406);
nor U4784 (N_4784,N_4229,N_4287);
and U4785 (N_4785,N_4441,N_4445);
and U4786 (N_4786,N_4260,N_4282);
nor U4787 (N_4787,N_4392,N_4356);
and U4788 (N_4788,N_4297,N_4238);
nor U4789 (N_4789,N_4342,N_4430);
and U4790 (N_4790,N_4309,N_4224);
xor U4791 (N_4791,N_4411,N_4202);
nor U4792 (N_4792,N_4251,N_4489);
nand U4793 (N_4793,N_4359,N_4453);
nand U4794 (N_4794,N_4363,N_4268);
xnor U4795 (N_4795,N_4483,N_4366);
nor U4796 (N_4796,N_4435,N_4202);
nand U4797 (N_4797,N_4385,N_4258);
nor U4798 (N_4798,N_4297,N_4293);
and U4799 (N_4799,N_4319,N_4331);
and U4800 (N_4800,N_4660,N_4600);
xor U4801 (N_4801,N_4552,N_4673);
nand U4802 (N_4802,N_4645,N_4696);
xnor U4803 (N_4803,N_4727,N_4774);
or U4804 (N_4804,N_4702,N_4598);
and U4805 (N_4805,N_4732,N_4761);
or U4806 (N_4806,N_4567,N_4762);
nor U4807 (N_4807,N_4728,N_4664);
nor U4808 (N_4808,N_4522,N_4618);
or U4809 (N_4809,N_4576,N_4633);
nand U4810 (N_4810,N_4563,N_4776);
xor U4811 (N_4811,N_4646,N_4791);
nand U4812 (N_4812,N_4580,N_4715);
and U4813 (N_4813,N_4675,N_4655);
nor U4814 (N_4814,N_4706,N_4595);
xnor U4815 (N_4815,N_4579,N_4513);
xnor U4816 (N_4816,N_4694,N_4765);
or U4817 (N_4817,N_4764,N_4500);
or U4818 (N_4818,N_4773,N_4707);
and U4819 (N_4819,N_4797,N_4687);
xor U4820 (N_4820,N_4748,N_4670);
and U4821 (N_4821,N_4672,N_4653);
or U4822 (N_4822,N_4789,N_4690);
nor U4823 (N_4823,N_4516,N_4740);
xnor U4824 (N_4824,N_4657,N_4613);
nand U4825 (N_4825,N_4527,N_4794);
nor U4826 (N_4826,N_4544,N_4724);
xnor U4827 (N_4827,N_4753,N_4575);
and U4828 (N_4828,N_4640,N_4685);
or U4829 (N_4829,N_4713,N_4754);
nor U4830 (N_4830,N_4506,N_4784);
and U4831 (N_4831,N_4622,N_4757);
nand U4832 (N_4832,N_4572,N_4532);
nor U4833 (N_4833,N_4537,N_4631);
or U4834 (N_4834,N_4708,N_4635);
xor U4835 (N_4835,N_4534,N_4693);
xnor U4836 (N_4836,N_4745,N_4529);
or U4837 (N_4837,N_4746,N_4712);
or U4838 (N_4838,N_4570,N_4790);
xor U4839 (N_4839,N_4744,N_4663);
nor U4840 (N_4840,N_4583,N_4639);
or U4841 (N_4841,N_4584,N_4768);
nand U4842 (N_4842,N_4667,N_4709);
and U4843 (N_4843,N_4629,N_4799);
and U4844 (N_4844,N_4602,N_4559);
nor U4845 (N_4845,N_4671,N_4772);
and U4846 (N_4846,N_4738,N_4551);
nor U4847 (N_4847,N_4780,N_4502);
nand U4848 (N_4848,N_4592,N_4758);
xnor U4849 (N_4849,N_4662,N_4766);
xor U4850 (N_4850,N_4620,N_4603);
nor U4851 (N_4851,N_4718,N_4778);
nand U4852 (N_4852,N_4755,N_4628);
and U4853 (N_4853,N_4651,N_4779);
or U4854 (N_4854,N_4553,N_4697);
and U4855 (N_4855,N_4535,N_4734);
or U4856 (N_4856,N_4782,N_4607);
xor U4857 (N_4857,N_4679,N_4538);
and U4858 (N_4858,N_4616,N_4688);
nand U4859 (N_4859,N_4573,N_4684);
or U4860 (N_4860,N_4503,N_4523);
and U4861 (N_4861,N_4601,N_4669);
nand U4862 (N_4862,N_4710,N_4723);
and U4863 (N_4863,N_4548,N_4650);
and U4864 (N_4864,N_4652,N_4729);
nor U4865 (N_4865,N_4659,N_4704);
and U4866 (N_4866,N_4725,N_4751);
nor U4867 (N_4867,N_4788,N_4641);
xor U4868 (N_4868,N_4610,N_4519);
nor U4869 (N_4869,N_4599,N_4731);
nand U4870 (N_4870,N_4756,N_4624);
and U4871 (N_4871,N_4666,N_4578);
and U4872 (N_4872,N_4643,N_4648);
xor U4873 (N_4873,N_4569,N_4665);
and U4874 (N_4874,N_4531,N_4759);
or U4875 (N_4875,N_4589,N_4509);
and U4876 (N_4876,N_4545,N_4526);
xnor U4877 (N_4877,N_4504,N_4783);
and U4878 (N_4878,N_4582,N_4689);
nand U4879 (N_4879,N_4612,N_4614);
or U4880 (N_4880,N_4590,N_4507);
and U4881 (N_4881,N_4515,N_4717);
or U4882 (N_4882,N_4777,N_4763);
and U4883 (N_4883,N_4542,N_4514);
or U4884 (N_4884,N_4691,N_4550);
nor U4885 (N_4885,N_4739,N_4543);
xnor U4886 (N_4886,N_4656,N_4677);
nor U4887 (N_4887,N_4686,N_4742);
xor U4888 (N_4888,N_4521,N_4591);
nand U4889 (N_4889,N_4554,N_4637);
xnor U4890 (N_4890,N_4597,N_4647);
or U4891 (N_4891,N_4747,N_4668);
nand U4892 (N_4892,N_4501,N_4781);
xor U4893 (N_4893,N_4630,N_4661);
nand U4894 (N_4894,N_4626,N_4604);
nor U4895 (N_4895,N_4741,N_4611);
xnor U4896 (N_4896,N_4769,N_4508);
nand U4897 (N_4897,N_4593,N_4528);
and U4898 (N_4898,N_4596,N_4556);
nand U4899 (N_4899,N_4692,N_4705);
or U4900 (N_4900,N_4505,N_4581);
or U4901 (N_4901,N_4649,N_4566);
nor U4902 (N_4902,N_4703,N_4736);
or U4903 (N_4903,N_4577,N_4638);
nand U4904 (N_4904,N_4644,N_4619);
xnor U4905 (N_4905,N_4726,N_4564);
and U4906 (N_4906,N_4711,N_4609);
xor U4907 (N_4907,N_4750,N_4621);
nand U4908 (N_4908,N_4558,N_4512);
and U4909 (N_4909,N_4634,N_4733);
xnor U4910 (N_4910,N_4721,N_4615);
nand U4911 (N_4911,N_4796,N_4605);
nor U4912 (N_4912,N_4795,N_4625);
and U4913 (N_4913,N_4700,N_4520);
xor U4914 (N_4914,N_4525,N_4722);
or U4915 (N_4915,N_4682,N_4561);
xnor U4916 (N_4916,N_4536,N_4557);
nor U4917 (N_4917,N_4793,N_4524);
and U4918 (N_4918,N_4530,N_4540);
nor U4919 (N_4919,N_4585,N_4658);
xnor U4920 (N_4920,N_4719,N_4760);
and U4921 (N_4921,N_4623,N_4771);
xnor U4922 (N_4922,N_4517,N_4632);
nand U4923 (N_4923,N_4586,N_4786);
or U4924 (N_4924,N_4730,N_4720);
or U4925 (N_4925,N_4716,N_4627);
or U4926 (N_4926,N_4701,N_4565);
or U4927 (N_4927,N_4606,N_4608);
nor U4928 (N_4928,N_4792,N_4574);
nand U4929 (N_4929,N_4533,N_4511);
nor U4930 (N_4930,N_4555,N_4699);
or U4931 (N_4931,N_4737,N_4695);
xor U4932 (N_4932,N_4588,N_4642);
and U4933 (N_4933,N_4743,N_4510);
xor U4934 (N_4934,N_4676,N_4680);
nand U4935 (N_4935,N_4678,N_4518);
nand U4936 (N_4936,N_4541,N_4549);
or U4937 (N_4937,N_4767,N_4539);
or U4938 (N_4938,N_4798,N_4546);
nor U4939 (N_4939,N_4587,N_4571);
xnor U4940 (N_4940,N_4547,N_4594);
nor U4941 (N_4941,N_4714,N_4787);
nor U4942 (N_4942,N_4749,N_4674);
and U4943 (N_4943,N_4698,N_4681);
and U4944 (N_4944,N_4683,N_4562);
nand U4945 (N_4945,N_4636,N_4654);
xnor U4946 (N_4946,N_4735,N_4785);
xor U4947 (N_4947,N_4617,N_4775);
and U4948 (N_4948,N_4560,N_4770);
nor U4949 (N_4949,N_4752,N_4568);
and U4950 (N_4950,N_4621,N_4507);
nand U4951 (N_4951,N_4564,N_4518);
or U4952 (N_4952,N_4768,N_4534);
nand U4953 (N_4953,N_4751,N_4612);
nand U4954 (N_4954,N_4593,N_4588);
or U4955 (N_4955,N_4726,N_4729);
nand U4956 (N_4956,N_4607,N_4670);
xor U4957 (N_4957,N_4695,N_4634);
nand U4958 (N_4958,N_4511,N_4779);
or U4959 (N_4959,N_4761,N_4700);
xnor U4960 (N_4960,N_4561,N_4605);
nand U4961 (N_4961,N_4708,N_4641);
or U4962 (N_4962,N_4797,N_4656);
or U4963 (N_4963,N_4652,N_4586);
xor U4964 (N_4964,N_4745,N_4640);
and U4965 (N_4965,N_4616,N_4710);
or U4966 (N_4966,N_4751,N_4519);
nand U4967 (N_4967,N_4741,N_4503);
nand U4968 (N_4968,N_4786,N_4594);
nor U4969 (N_4969,N_4632,N_4585);
nor U4970 (N_4970,N_4533,N_4779);
nand U4971 (N_4971,N_4588,N_4549);
xnor U4972 (N_4972,N_4523,N_4664);
or U4973 (N_4973,N_4732,N_4796);
or U4974 (N_4974,N_4774,N_4687);
and U4975 (N_4975,N_4599,N_4586);
and U4976 (N_4976,N_4529,N_4793);
or U4977 (N_4977,N_4592,N_4793);
or U4978 (N_4978,N_4659,N_4547);
and U4979 (N_4979,N_4794,N_4776);
nor U4980 (N_4980,N_4676,N_4799);
nor U4981 (N_4981,N_4726,N_4577);
and U4982 (N_4982,N_4720,N_4744);
xnor U4983 (N_4983,N_4611,N_4773);
nor U4984 (N_4984,N_4645,N_4785);
nand U4985 (N_4985,N_4779,N_4529);
nor U4986 (N_4986,N_4552,N_4609);
nand U4987 (N_4987,N_4738,N_4565);
nor U4988 (N_4988,N_4615,N_4589);
xor U4989 (N_4989,N_4642,N_4550);
or U4990 (N_4990,N_4787,N_4771);
xor U4991 (N_4991,N_4517,N_4672);
nand U4992 (N_4992,N_4766,N_4682);
nor U4993 (N_4993,N_4689,N_4778);
xnor U4994 (N_4994,N_4586,N_4527);
xor U4995 (N_4995,N_4794,N_4540);
nand U4996 (N_4996,N_4752,N_4785);
and U4997 (N_4997,N_4568,N_4700);
nor U4998 (N_4998,N_4513,N_4582);
nand U4999 (N_4999,N_4585,N_4789);
and U5000 (N_5000,N_4607,N_4701);
xor U5001 (N_5001,N_4548,N_4777);
and U5002 (N_5002,N_4700,N_4547);
nor U5003 (N_5003,N_4788,N_4724);
and U5004 (N_5004,N_4608,N_4503);
xnor U5005 (N_5005,N_4693,N_4600);
or U5006 (N_5006,N_4612,N_4691);
xnor U5007 (N_5007,N_4755,N_4697);
nor U5008 (N_5008,N_4724,N_4746);
or U5009 (N_5009,N_4570,N_4794);
xnor U5010 (N_5010,N_4762,N_4770);
xor U5011 (N_5011,N_4629,N_4534);
xnor U5012 (N_5012,N_4738,N_4639);
nand U5013 (N_5013,N_4525,N_4772);
nand U5014 (N_5014,N_4523,N_4569);
and U5015 (N_5015,N_4534,N_4597);
or U5016 (N_5016,N_4545,N_4507);
or U5017 (N_5017,N_4578,N_4558);
or U5018 (N_5018,N_4522,N_4577);
nand U5019 (N_5019,N_4583,N_4552);
nor U5020 (N_5020,N_4745,N_4521);
and U5021 (N_5021,N_4760,N_4727);
xnor U5022 (N_5022,N_4790,N_4512);
nor U5023 (N_5023,N_4670,N_4636);
or U5024 (N_5024,N_4703,N_4578);
nor U5025 (N_5025,N_4794,N_4761);
xnor U5026 (N_5026,N_4678,N_4782);
nand U5027 (N_5027,N_4632,N_4625);
nand U5028 (N_5028,N_4705,N_4568);
nor U5029 (N_5029,N_4548,N_4780);
nand U5030 (N_5030,N_4502,N_4766);
xor U5031 (N_5031,N_4643,N_4577);
and U5032 (N_5032,N_4709,N_4723);
xor U5033 (N_5033,N_4709,N_4610);
and U5034 (N_5034,N_4620,N_4661);
nor U5035 (N_5035,N_4642,N_4685);
xnor U5036 (N_5036,N_4701,N_4557);
or U5037 (N_5037,N_4538,N_4699);
and U5038 (N_5038,N_4748,N_4702);
or U5039 (N_5039,N_4753,N_4549);
nor U5040 (N_5040,N_4576,N_4594);
nor U5041 (N_5041,N_4723,N_4769);
xnor U5042 (N_5042,N_4697,N_4585);
nor U5043 (N_5043,N_4549,N_4689);
and U5044 (N_5044,N_4798,N_4638);
xor U5045 (N_5045,N_4782,N_4618);
and U5046 (N_5046,N_4683,N_4536);
nand U5047 (N_5047,N_4744,N_4555);
nor U5048 (N_5048,N_4796,N_4542);
xnor U5049 (N_5049,N_4616,N_4746);
and U5050 (N_5050,N_4786,N_4731);
nand U5051 (N_5051,N_4739,N_4790);
or U5052 (N_5052,N_4676,N_4697);
or U5053 (N_5053,N_4508,N_4507);
xor U5054 (N_5054,N_4656,N_4643);
and U5055 (N_5055,N_4506,N_4543);
or U5056 (N_5056,N_4503,N_4621);
nand U5057 (N_5057,N_4753,N_4764);
nand U5058 (N_5058,N_4638,N_4657);
or U5059 (N_5059,N_4679,N_4527);
and U5060 (N_5060,N_4770,N_4576);
nor U5061 (N_5061,N_4568,N_4633);
or U5062 (N_5062,N_4757,N_4794);
nand U5063 (N_5063,N_4551,N_4678);
xnor U5064 (N_5064,N_4661,N_4704);
and U5065 (N_5065,N_4611,N_4657);
nor U5066 (N_5066,N_4789,N_4703);
nand U5067 (N_5067,N_4582,N_4503);
xor U5068 (N_5068,N_4689,N_4572);
xor U5069 (N_5069,N_4648,N_4770);
or U5070 (N_5070,N_4665,N_4655);
or U5071 (N_5071,N_4698,N_4787);
and U5072 (N_5072,N_4700,N_4639);
and U5073 (N_5073,N_4667,N_4763);
and U5074 (N_5074,N_4555,N_4749);
nor U5075 (N_5075,N_4730,N_4533);
or U5076 (N_5076,N_4603,N_4796);
or U5077 (N_5077,N_4609,N_4624);
nand U5078 (N_5078,N_4688,N_4604);
nand U5079 (N_5079,N_4765,N_4727);
or U5080 (N_5080,N_4636,N_4647);
or U5081 (N_5081,N_4799,N_4518);
xor U5082 (N_5082,N_4771,N_4683);
nor U5083 (N_5083,N_4553,N_4544);
or U5084 (N_5084,N_4673,N_4648);
nor U5085 (N_5085,N_4646,N_4518);
nand U5086 (N_5086,N_4595,N_4575);
nor U5087 (N_5087,N_4644,N_4695);
xor U5088 (N_5088,N_4603,N_4554);
and U5089 (N_5089,N_4524,N_4586);
and U5090 (N_5090,N_4709,N_4632);
nor U5091 (N_5091,N_4639,N_4510);
and U5092 (N_5092,N_4749,N_4731);
and U5093 (N_5093,N_4672,N_4754);
nor U5094 (N_5094,N_4673,N_4694);
nor U5095 (N_5095,N_4706,N_4546);
nor U5096 (N_5096,N_4543,N_4666);
and U5097 (N_5097,N_4513,N_4710);
and U5098 (N_5098,N_4519,N_4609);
xnor U5099 (N_5099,N_4620,N_4537);
or U5100 (N_5100,N_5007,N_5091);
and U5101 (N_5101,N_5002,N_4813);
and U5102 (N_5102,N_5063,N_4970);
nor U5103 (N_5103,N_5065,N_4869);
or U5104 (N_5104,N_4887,N_5028);
xor U5105 (N_5105,N_4845,N_4913);
xor U5106 (N_5106,N_4877,N_5039);
nand U5107 (N_5107,N_5046,N_5030);
or U5108 (N_5108,N_5029,N_4925);
or U5109 (N_5109,N_4908,N_4894);
or U5110 (N_5110,N_4800,N_4885);
or U5111 (N_5111,N_5000,N_4884);
or U5112 (N_5112,N_4814,N_4860);
or U5113 (N_5113,N_4927,N_5097);
and U5114 (N_5114,N_4902,N_5021);
or U5115 (N_5115,N_4909,N_4937);
or U5116 (N_5116,N_4967,N_5053);
xnor U5117 (N_5117,N_4897,N_4947);
nand U5118 (N_5118,N_5026,N_4898);
xor U5119 (N_5119,N_5008,N_4963);
nand U5120 (N_5120,N_4899,N_5031);
nand U5121 (N_5121,N_4969,N_5050);
xnor U5122 (N_5122,N_4951,N_4900);
xnor U5123 (N_5123,N_5015,N_5069);
nand U5124 (N_5124,N_4914,N_4838);
nor U5125 (N_5125,N_4819,N_5057);
and U5126 (N_5126,N_4916,N_5013);
nor U5127 (N_5127,N_4843,N_4961);
xnor U5128 (N_5128,N_4934,N_4857);
nand U5129 (N_5129,N_5019,N_5098);
nand U5130 (N_5130,N_4805,N_4818);
nor U5131 (N_5131,N_4865,N_5062);
and U5132 (N_5132,N_4972,N_4985);
nand U5133 (N_5133,N_4876,N_5092);
xor U5134 (N_5134,N_4991,N_4935);
xor U5135 (N_5135,N_4923,N_5090);
or U5136 (N_5136,N_4983,N_4821);
nor U5137 (N_5137,N_4945,N_5049);
nor U5138 (N_5138,N_5014,N_4835);
and U5139 (N_5139,N_4825,N_4806);
nor U5140 (N_5140,N_4979,N_5075);
or U5141 (N_5141,N_4901,N_4872);
nor U5142 (N_5142,N_4842,N_4816);
and U5143 (N_5143,N_5051,N_4809);
nor U5144 (N_5144,N_4994,N_5085);
nor U5145 (N_5145,N_4988,N_4866);
nor U5146 (N_5146,N_4933,N_5009);
nor U5147 (N_5147,N_4943,N_4826);
nand U5148 (N_5148,N_4807,N_5079);
nor U5149 (N_5149,N_4941,N_4839);
nand U5150 (N_5150,N_4893,N_4989);
and U5151 (N_5151,N_4949,N_4803);
and U5152 (N_5152,N_4980,N_4844);
and U5153 (N_5153,N_4811,N_5033);
nor U5154 (N_5154,N_4827,N_5006);
or U5155 (N_5155,N_4862,N_5083);
xor U5156 (N_5156,N_5077,N_4948);
or U5157 (N_5157,N_4837,N_5059);
nor U5158 (N_5158,N_4846,N_5074);
or U5159 (N_5159,N_4931,N_4956);
xnor U5160 (N_5160,N_5099,N_4996);
nor U5161 (N_5161,N_4804,N_4997);
or U5162 (N_5162,N_4836,N_5052);
nand U5163 (N_5163,N_4929,N_5066);
nor U5164 (N_5164,N_4995,N_5071);
nand U5165 (N_5165,N_5094,N_4822);
nand U5166 (N_5166,N_4964,N_4832);
or U5167 (N_5167,N_4848,N_5016);
nand U5168 (N_5168,N_4841,N_5034);
or U5169 (N_5169,N_5023,N_4858);
or U5170 (N_5170,N_5073,N_4810);
or U5171 (N_5171,N_4875,N_5048);
xor U5172 (N_5172,N_4856,N_4871);
nand U5173 (N_5173,N_4957,N_4987);
and U5174 (N_5174,N_4863,N_4958);
and U5175 (N_5175,N_4984,N_4840);
nor U5176 (N_5176,N_5084,N_4878);
nand U5177 (N_5177,N_4801,N_5078);
and U5178 (N_5178,N_4944,N_4938);
xnor U5179 (N_5179,N_4855,N_4920);
nor U5180 (N_5180,N_4939,N_5025);
and U5181 (N_5181,N_4880,N_5080);
nand U5182 (N_5182,N_4918,N_4881);
or U5183 (N_5183,N_5041,N_5087);
nand U5184 (N_5184,N_4829,N_4982);
nor U5185 (N_5185,N_4946,N_5045);
nand U5186 (N_5186,N_4867,N_4890);
or U5187 (N_5187,N_4849,N_4990);
and U5188 (N_5188,N_4930,N_4873);
and U5189 (N_5189,N_5093,N_4993);
or U5190 (N_5190,N_4895,N_5040);
or U5191 (N_5191,N_4952,N_4815);
and U5192 (N_5192,N_4975,N_5038);
or U5193 (N_5193,N_4905,N_4828);
nand U5194 (N_5194,N_5043,N_5003);
or U5195 (N_5195,N_5012,N_4955);
or U5196 (N_5196,N_4824,N_4977);
nor U5197 (N_5197,N_4959,N_4820);
and U5198 (N_5198,N_5064,N_5067);
nor U5199 (N_5199,N_5035,N_5095);
and U5200 (N_5200,N_4896,N_4864);
or U5201 (N_5201,N_5068,N_5061);
nand U5202 (N_5202,N_4892,N_4850);
xnor U5203 (N_5203,N_5024,N_4907);
nand U5204 (N_5204,N_5047,N_4962);
and U5205 (N_5205,N_4879,N_4942);
xor U5206 (N_5206,N_4834,N_5044);
nand U5207 (N_5207,N_5017,N_4999);
xnor U5208 (N_5208,N_4974,N_5005);
nor U5209 (N_5209,N_4953,N_4868);
nand U5210 (N_5210,N_5060,N_4919);
xor U5211 (N_5211,N_4992,N_4926);
xnor U5212 (N_5212,N_4861,N_5001);
or U5213 (N_5213,N_4903,N_5055);
and U5214 (N_5214,N_4928,N_5010);
nand U5215 (N_5215,N_4888,N_4817);
nor U5216 (N_5216,N_5096,N_5042);
nand U5217 (N_5217,N_4954,N_4833);
and U5218 (N_5218,N_4976,N_5058);
or U5219 (N_5219,N_4906,N_4950);
and U5220 (N_5220,N_4981,N_5032);
nor U5221 (N_5221,N_4965,N_4853);
nor U5222 (N_5222,N_5037,N_5082);
nor U5223 (N_5223,N_5036,N_5086);
and U5224 (N_5224,N_4940,N_5004);
xor U5225 (N_5225,N_4859,N_4851);
and U5226 (N_5226,N_4973,N_4823);
nor U5227 (N_5227,N_4917,N_4922);
nand U5228 (N_5228,N_4911,N_4870);
or U5229 (N_5229,N_4912,N_4936);
and U5230 (N_5230,N_4854,N_5076);
xnor U5231 (N_5231,N_4889,N_5056);
or U5232 (N_5232,N_5022,N_4904);
and U5233 (N_5233,N_5011,N_4966);
and U5234 (N_5234,N_4847,N_4831);
and U5235 (N_5235,N_4915,N_4971);
nor U5236 (N_5236,N_5088,N_5072);
xnor U5237 (N_5237,N_4812,N_4891);
or U5238 (N_5238,N_4998,N_4830);
nand U5239 (N_5239,N_4968,N_5070);
or U5240 (N_5240,N_4921,N_5081);
nor U5241 (N_5241,N_4986,N_4808);
xor U5242 (N_5242,N_4882,N_4802);
nand U5243 (N_5243,N_4910,N_5018);
and U5244 (N_5244,N_5027,N_4883);
nor U5245 (N_5245,N_5020,N_4874);
nor U5246 (N_5246,N_5089,N_4924);
or U5247 (N_5247,N_4978,N_4932);
nor U5248 (N_5248,N_4960,N_4852);
and U5249 (N_5249,N_4886,N_5054);
nand U5250 (N_5250,N_4871,N_4829);
nand U5251 (N_5251,N_4974,N_5041);
or U5252 (N_5252,N_5020,N_4993);
xor U5253 (N_5253,N_4954,N_4865);
xnor U5254 (N_5254,N_4833,N_5022);
and U5255 (N_5255,N_4899,N_4952);
or U5256 (N_5256,N_4994,N_5017);
nor U5257 (N_5257,N_4966,N_4971);
or U5258 (N_5258,N_5059,N_4907);
and U5259 (N_5259,N_5092,N_4891);
nor U5260 (N_5260,N_4840,N_5073);
or U5261 (N_5261,N_4816,N_4808);
nor U5262 (N_5262,N_4968,N_4949);
nand U5263 (N_5263,N_4915,N_5053);
nor U5264 (N_5264,N_4887,N_5024);
nand U5265 (N_5265,N_4915,N_4964);
xor U5266 (N_5266,N_4961,N_5050);
and U5267 (N_5267,N_4852,N_5071);
nor U5268 (N_5268,N_4978,N_4973);
or U5269 (N_5269,N_4951,N_4845);
nand U5270 (N_5270,N_5028,N_4858);
or U5271 (N_5271,N_4976,N_4855);
xnor U5272 (N_5272,N_4996,N_4997);
nand U5273 (N_5273,N_5081,N_5057);
or U5274 (N_5274,N_4938,N_5062);
and U5275 (N_5275,N_5059,N_4856);
and U5276 (N_5276,N_4831,N_4941);
xor U5277 (N_5277,N_4859,N_4937);
xor U5278 (N_5278,N_4942,N_4869);
xor U5279 (N_5279,N_4943,N_4919);
xnor U5280 (N_5280,N_4948,N_5036);
nor U5281 (N_5281,N_4827,N_4895);
and U5282 (N_5282,N_5003,N_5041);
or U5283 (N_5283,N_5035,N_5069);
nor U5284 (N_5284,N_5090,N_4981);
xnor U5285 (N_5285,N_4885,N_4964);
or U5286 (N_5286,N_4844,N_4929);
nand U5287 (N_5287,N_4960,N_4927);
nand U5288 (N_5288,N_4847,N_4865);
xor U5289 (N_5289,N_4896,N_4819);
xor U5290 (N_5290,N_4999,N_4930);
or U5291 (N_5291,N_4939,N_4966);
nor U5292 (N_5292,N_4923,N_4983);
or U5293 (N_5293,N_5012,N_5087);
nand U5294 (N_5294,N_4846,N_4983);
xor U5295 (N_5295,N_4812,N_4966);
nor U5296 (N_5296,N_4836,N_4904);
nand U5297 (N_5297,N_4911,N_4827);
nor U5298 (N_5298,N_4800,N_4809);
or U5299 (N_5299,N_5059,N_5093);
or U5300 (N_5300,N_4837,N_4843);
nand U5301 (N_5301,N_4997,N_5086);
nand U5302 (N_5302,N_5050,N_5034);
and U5303 (N_5303,N_5059,N_4803);
nand U5304 (N_5304,N_4963,N_5095);
xnor U5305 (N_5305,N_4878,N_5055);
nor U5306 (N_5306,N_5072,N_4958);
or U5307 (N_5307,N_4909,N_4933);
or U5308 (N_5308,N_4942,N_4963);
xor U5309 (N_5309,N_4889,N_5026);
nor U5310 (N_5310,N_4984,N_4997);
nor U5311 (N_5311,N_5003,N_4901);
and U5312 (N_5312,N_4934,N_4923);
and U5313 (N_5313,N_4948,N_4875);
and U5314 (N_5314,N_4956,N_5010);
xnor U5315 (N_5315,N_4844,N_4840);
nor U5316 (N_5316,N_4832,N_4958);
and U5317 (N_5317,N_4813,N_5062);
and U5318 (N_5318,N_4961,N_4853);
nor U5319 (N_5319,N_4970,N_4820);
and U5320 (N_5320,N_5086,N_4927);
or U5321 (N_5321,N_4836,N_5084);
nand U5322 (N_5322,N_4871,N_4875);
nor U5323 (N_5323,N_4901,N_4937);
or U5324 (N_5324,N_4854,N_4943);
nor U5325 (N_5325,N_4892,N_4927);
and U5326 (N_5326,N_5023,N_4902);
nand U5327 (N_5327,N_4911,N_5081);
nor U5328 (N_5328,N_5096,N_4916);
xor U5329 (N_5329,N_5028,N_5007);
or U5330 (N_5330,N_5065,N_5063);
nand U5331 (N_5331,N_4891,N_4984);
nor U5332 (N_5332,N_4906,N_4876);
xnor U5333 (N_5333,N_5005,N_4959);
or U5334 (N_5334,N_4930,N_4915);
or U5335 (N_5335,N_5004,N_4905);
and U5336 (N_5336,N_5022,N_4891);
and U5337 (N_5337,N_4824,N_4995);
and U5338 (N_5338,N_4940,N_4835);
nand U5339 (N_5339,N_4926,N_4815);
or U5340 (N_5340,N_4958,N_4984);
or U5341 (N_5341,N_4920,N_4876);
nor U5342 (N_5342,N_4974,N_4818);
nor U5343 (N_5343,N_4869,N_5053);
and U5344 (N_5344,N_4864,N_4911);
nand U5345 (N_5345,N_4924,N_5002);
xor U5346 (N_5346,N_5006,N_4881);
and U5347 (N_5347,N_5040,N_4993);
and U5348 (N_5348,N_4819,N_4827);
xor U5349 (N_5349,N_5086,N_4889);
nand U5350 (N_5350,N_5023,N_4995);
or U5351 (N_5351,N_4865,N_4980);
nand U5352 (N_5352,N_4970,N_4804);
nand U5353 (N_5353,N_5075,N_4854);
and U5354 (N_5354,N_5083,N_5003);
and U5355 (N_5355,N_4850,N_4945);
and U5356 (N_5356,N_5028,N_4812);
and U5357 (N_5357,N_4858,N_4990);
and U5358 (N_5358,N_5058,N_4857);
nand U5359 (N_5359,N_4914,N_4886);
nand U5360 (N_5360,N_5044,N_5096);
or U5361 (N_5361,N_4877,N_5067);
nand U5362 (N_5362,N_5032,N_5008);
or U5363 (N_5363,N_4872,N_4834);
xnor U5364 (N_5364,N_4987,N_5053);
nor U5365 (N_5365,N_5031,N_5016);
nor U5366 (N_5366,N_4825,N_4970);
or U5367 (N_5367,N_4931,N_4872);
xor U5368 (N_5368,N_4849,N_5045);
nand U5369 (N_5369,N_5079,N_4987);
or U5370 (N_5370,N_5014,N_4978);
xnor U5371 (N_5371,N_4934,N_5032);
nor U5372 (N_5372,N_5062,N_5066);
and U5373 (N_5373,N_4892,N_5044);
or U5374 (N_5374,N_4824,N_4876);
or U5375 (N_5375,N_4943,N_4918);
nand U5376 (N_5376,N_5003,N_4859);
and U5377 (N_5377,N_5076,N_5045);
xnor U5378 (N_5378,N_4857,N_4963);
xnor U5379 (N_5379,N_4935,N_5036);
xor U5380 (N_5380,N_4822,N_4817);
xnor U5381 (N_5381,N_4826,N_4913);
nor U5382 (N_5382,N_5089,N_4929);
nor U5383 (N_5383,N_4847,N_5026);
or U5384 (N_5384,N_5027,N_4896);
and U5385 (N_5385,N_5070,N_4867);
nor U5386 (N_5386,N_4827,N_5037);
nand U5387 (N_5387,N_4939,N_5006);
and U5388 (N_5388,N_5017,N_4909);
and U5389 (N_5389,N_4954,N_5051);
nor U5390 (N_5390,N_4913,N_4956);
nand U5391 (N_5391,N_4949,N_4893);
or U5392 (N_5392,N_4992,N_4894);
and U5393 (N_5393,N_4912,N_4944);
or U5394 (N_5394,N_4994,N_5063);
xor U5395 (N_5395,N_4889,N_4853);
and U5396 (N_5396,N_4989,N_5011);
and U5397 (N_5397,N_5098,N_4822);
nand U5398 (N_5398,N_4969,N_5007);
xor U5399 (N_5399,N_4956,N_4827);
and U5400 (N_5400,N_5354,N_5293);
or U5401 (N_5401,N_5390,N_5223);
and U5402 (N_5402,N_5149,N_5148);
or U5403 (N_5403,N_5271,N_5369);
nand U5404 (N_5404,N_5257,N_5196);
or U5405 (N_5405,N_5353,N_5222);
nand U5406 (N_5406,N_5343,N_5101);
or U5407 (N_5407,N_5323,N_5305);
xor U5408 (N_5408,N_5307,N_5247);
and U5409 (N_5409,N_5238,N_5392);
nand U5410 (N_5410,N_5302,N_5251);
nor U5411 (N_5411,N_5322,N_5108);
xnor U5412 (N_5412,N_5180,N_5132);
or U5413 (N_5413,N_5349,N_5113);
nand U5414 (N_5414,N_5172,N_5378);
and U5415 (N_5415,N_5304,N_5135);
nand U5416 (N_5416,N_5208,N_5275);
nor U5417 (N_5417,N_5311,N_5170);
nor U5418 (N_5418,N_5255,N_5258);
nor U5419 (N_5419,N_5127,N_5168);
xor U5420 (N_5420,N_5204,N_5233);
and U5421 (N_5421,N_5285,N_5174);
and U5422 (N_5422,N_5143,N_5176);
and U5423 (N_5423,N_5294,N_5391);
and U5424 (N_5424,N_5296,N_5229);
or U5425 (N_5425,N_5125,N_5318);
and U5426 (N_5426,N_5279,N_5320);
nand U5427 (N_5427,N_5341,N_5260);
nor U5428 (N_5428,N_5201,N_5188);
and U5429 (N_5429,N_5380,N_5191);
xor U5430 (N_5430,N_5252,N_5206);
or U5431 (N_5431,N_5399,N_5144);
xor U5432 (N_5432,N_5227,N_5331);
or U5433 (N_5433,N_5129,N_5230);
nor U5434 (N_5434,N_5335,N_5287);
nand U5435 (N_5435,N_5240,N_5209);
nor U5436 (N_5436,N_5126,N_5321);
xor U5437 (N_5437,N_5315,N_5217);
xnor U5438 (N_5438,N_5379,N_5398);
xor U5439 (N_5439,N_5329,N_5396);
nor U5440 (N_5440,N_5363,N_5151);
and U5441 (N_5441,N_5376,N_5266);
or U5442 (N_5442,N_5212,N_5122);
nand U5443 (N_5443,N_5102,N_5199);
xor U5444 (N_5444,N_5225,N_5189);
xor U5445 (N_5445,N_5393,N_5310);
nand U5446 (N_5446,N_5181,N_5193);
or U5447 (N_5447,N_5299,N_5339);
xor U5448 (N_5448,N_5364,N_5138);
nor U5449 (N_5449,N_5219,N_5270);
nand U5450 (N_5450,N_5207,N_5185);
or U5451 (N_5451,N_5348,N_5337);
xor U5452 (N_5452,N_5194,N_5111);
or U5453 (N_5453,N_5355,N_5152);
xor U5454 (N_5454,N_5274,N_5309);
nor U5455 (N_5455,N_5298,N_5159);
nor U5456 (N_5456,N_5277,N_5308);
xnor U5457 (N_5457,N_5192,N_5130);
or U5458 (N_5458,N_5216,N_5248);
xnor U5459 (N_5459,N_5316,N_5384);
nor U5460 (N_5460,N_5328,N_5134);
nor U5461 (N_5461,N_5179,N_5205);
and U5462 (N_5462,N_5203,N_5358);
nand U5463 (N_5463,N_5182,N_5351);
nand U5464 (N_5464,N_5186,N_5190);
or U5465 (N_5465,N_5202,N_5360);
xor U5466 (N_5466,N_5116,N_5264);
nand U5467 (N_5467,N_5104,N_5361);
nor U5468 (N_5468,N_5115,N_5338);
or U5469 (N_5469,N_5110,N_5128);
and U5470 (N_5470,N_5246,N_5156);
and U5471 (N_5471,N_5383,N_5187);
xnor U5472 (N_5472,N_5166,N_5288);
nor U5473 (N_5473,N_5243,N_5342);
nand U5474 (N_5474,N_5231,N_5261);
or U5475 (N_5475,N_5220,N_5362);
and U5476 (N_5476,N_5386,N_5313);
nor U5477 (N_5477,N_5344,N_5367);
xor U5478 (N_5478,N_5214,N_5112);
nor U5479 (N_5479,N_5356,N_5385);
or U5480 (N_5480,N_5119,N_5280);
and U5481 (N_5481,N_5211,N_5276);
nand U5482 (N_5482,N_5306,N_5325);
and U5483 (N_5483,N_5177,N_5210);
nor U5484 (N_5484,N_5103,N_5366);
xor U5485 (N_5485,N_5373,N_5272);
nor U5486 (N_5486,N_5388,N_5265);
and U5487 (N_5487,N_5105,N_5273);
nand U5488 (N_5488,N_5224,N_5160);
or U5489 (N_5489,N_5142,N_5200);
or U5490 (N_5490,N_5334,N_5154);
nand U5491 (N_5491,N_5368,N_5282);
or U5492 (N_5492,N_5336,N_5359);
or U5493 (N_5493,N_5153,N_5352);
nor U5494 (N_5494,N_5133,N_5340);
nand U5495 (N_5495,N_5256,N_5242);
nand U5496 (N_5496,N_5232,N_5345);
nand U5497 (N_5497,N_5381,N_5145);
xor U5498 (N_5498,N_5281,N_5213);
nor U5499 (N_5499,N_5297,N_5195);
nand U5500 (N_5500,N_5218,N_5162);
nor U5501 (N_5501,N_5124,N_5249);
and U5502 (N_5502,N_5371,N_5150);
or U5503 (N_5503,N_5158,N_5239);
or U5504 (N_5504,N_5165,N_5184);
nor U5505 (N_5505,N_5314,N_5241);
or U5506 (N_5506,N_5161,N_5109);
or U5507 (N_5507,N_5291,N_5327);
nor U5508 (N_5508,N_5155,N_5215);
xor U5509 (N_5509,N_5300,N_5183);
nor U5510 (N_5510,N_5139,N_5235);
nor U5511 (N_5511,N_5147,N_5395);
xor U5512 (N_5512,N_5263,N_5295);
xor U5513 (N_5513,N_5394,N_5167);
nand U5514 (N_5514,N_5346,N_5303);
xor U5515 (N_5515,N_5146,N_5120);
nor U5516 (N_5516,N_5136,N_5245);
or U5517 (N_5517,N_5269,N_5283);
nor U5518 (N_5518,N_5253,N_5157);
or U5519 (N_5519,N_5326,N_5237);
nor U5520 (N_5520,N_5317,N_5301);
or U5521 (N_5521,N_5123,N_5140);
nand U5522 (N_5522,N_5169,N_5357);
or U5523 (N_5523,N_5333,N_5289);
and U5524 (N_5524,N_5100,N_5374);
nor U5525 (N_5525,N_5290,N_5228);
and U5526 (N_5526,N_5106,N_5312);
nor U5527 (N_5527,N_5197,N_5121);
xor U5528 (N_5528,N_5330,N_5382);
or U5529 (N_5529,N_5278,N_5267);
nor U5530 (N_5530,N_5319,N_5365);
xor U5531 (N_5531,N_5163,N_5131);
nor U5532 (N_5532,N_5286,N_5198);
nand U5533 (N_5533,N_5332,N_5221);
and U5534 (N_5534,N_5372,N_5244);
or U5535 (N_5535,N_5175,N_5377);
nor U5536 (N_5536,N_5114,N_5226);
and U5537 (N_5537,N_5178,N_5236);
xor U5538 (N_5538,N_5171,N_5137);
or U5539 (N_5539,N_5324,N_5117);
xnor U5540 (N_5540,N_5234,N_5292);
or U5541 (N_5541,N_5268,N_5347);
and U5542 (N_5542,N_5387,N_5389);
nor U5543 (N_5543,N_5375,N_5254);
nand U5544 (N_5544,N_5397,N_5284);
or U5545 (N_5545,N_5173,N_5107);
or U5546 (N_5546,N_5370,N_5118);
xnor U5547 (N_5547,N_5259,N_5164);
xor U5548 (N_5548,N_5250,N_5262);
nand U5549 (N_5549,N_5141,N_5350);
nor U5550 (N_5550,N_5216,N_5157);
nor U5551 (N_5551,N_5239,N_5361);
or U5552 (N_5552,N_5157,N_5349);
or U5553 (N_5553,N_5134,N_5369);
nand U5554 (N_5554,N_5176,N_5391);
nor U5555 (N_5555,N_5225,N_5245);
nor U5556 (N_5556,N_5227,N_5105);
xor U5557 (N_5557,N_5208,N_5385);
and U5558 (N_5558,N_5276,N_5281);
xnor U5559 (N_5559,N_5101,N_5332);
nor U5560 (N_5560,N_5328,N_5154);
xor U5561 (N_5561,N_5352,N_5225);
xnor U5562 (N_5562,N_5163,N_5371);
nand U5563 (N_5563,N_5270,N_5203);
and U5564 (N_5564,N_5391,N_5210);
and U5565 (N_5565,N_5158,N_5217);
nand U5566 (N_5566,N_5148,N_5361);
and U5567 (N_5567,N_5260,N_5196);
nor U5568 (N_5568,N_5153,N_5264);
nor U5569 (N_5569,N_5181,N_5264);
and U5570 (N_5570,N_5171,N_5233);
xnor U5571 (N_5571,N_5214,N_5388);
nor U5572 (N_5572,N_5133,N_5111);
nand U5573 (N_5573,N_5274,N_5308);
nand U5574 (N_5574,N_5365,N_5348);
xor U5575 (N_5575,N_5214,N_5320);
and U5576 (N_5576,N_5275,N_5242);
and U5577 (N_5577,N_5197,N_5257);
nand U5578 (N_5578,N_5184,N_5139);
or U5579 (N_5579,N_5103,N_5314);
xor U5580 (N_5580,N_5108,N_5215);
or U5581 (N_5581,N_5193,N_5224);
or U5582 (N_5582,N_5258,N_5326);
and U5583 (N_5583,N_5347,N_5159);
nand U5584 (N_5584,N_5175,N_5104);
or U5585 (N_5585,N_5120,N_5251);
or U5586 (N_5586,N_5241,N_5370);
xor U5587 (N_5587,N_5166,N_5338);
and U5588 (N_5588,N_5211,N_5208);
or U5589 (N_5589,N_5218,N_5320);
and U5590 (N_5590,N_5366,N_5304);
xnor U5591 (N_5591,N_5178,N_5122);
or U5592 (N_5592,N_5280,N_5305);
xnor U5593 (N_5593,N_5231,N_5275);
nand U5594 (N_5594,N_5200,N_5139);
nor U5595 (N_5595,N_5234,N_5299);
and U5596 (N_5596,N_5352,N_5365);
or U5597 (N_5597,N_5277,N_5132);
xnor U5598 (N_5598,N_5242,N_5155);
xor U5599 (N_5599,N_5112,N_5341);
and U5600 (N_5600,N_5303,N_5208);
and U5601 (N_5601,N_5384,N_5269);
nand U5602 (N_5602,N_5213,N_5347);
and U5603 (N_5603,N_5133,N_5121);
or U5604 (N_5604,N_5273,N_5252);
or U5605 (N_5605,N_5337,N_5365);
nand U5606 (N_5606,N_5100,N_5322);
nor U5607 (N_5607,N_5314,N_5164);
and U5608 (N_5608,N_5165,N_5233);
nor U5609 (N_5609,N_5286,N_5158);
xnor U5610 (N_5610,N_5268,N_5105);
or U5611 (N_5611,N_5353,N_5133);
and U5612 (N_5612,N_5316,N_5272);
nand U5613 (N_5613,N_5249,N_5349);
xnor U5614 (N_5614,N_5296,N_5265);
nor U5615 (N_5615,N_5238,N_5317);
and U5616 (N_5616,N_5134,N_5309);
and U5617 (N_5617,N_5398,N_5216);
nand U5618 (N_5618,N_5180,N_5128);
or U5619 (N_5619,N_5344,N_5126);
or U5620 (N_5620,N_5102,N_5286);
nor U5621 (N_5621,N_5200,N_5140);
and U5622 (N_5622,N_5386,N_5244);
xor U5623 (N_5623,N_5348,N_5382);
nand U5624 (N_5624,N_5117,N_5300);
or U5625 (N_5625,N_5310,N_5307);
nor U5626 (N_5626,N_5104,N_5282);
and U5627 (N_5627,N_5373,N_5139);
or U5628 (N_5628,N_5157,N_5315);
xor U5629 (N_5629,N_5140,N_5366);
nor U5630 (N_5630,N_5347,N_5158);
xor U5631 (N_5631,N_5368,N_5297);
or U5632 (N_5632,N_5133,N_5209);
nor U5633 (N_5633,N_5312,N_5288);
nand U5634 (N_5634,N_5204,N_5399);
nand U5635 (N_5635,N_5382,N_5214);
nand U5636 (N_5636,N_5150,N_5200);
and U5637 (N_5637,N_5103,N_5273);
nand U5638 (N_5638,N_5318,N_5258);
or U5639 (N_5639,N_5238,N_5116);
and U5640 (N_5640,N_5337,N_5356);
nor U5641 (N_5641,N_5268,N_5108);
xnor U5642 (N_5642,N_5176,N_5225);
nand U5643 (N_5643,N_5309,N_5373);
xnor U5644 (N_5644,N_5118,N_5141);
nand U5645 (N_5645,N_5199,N_5208);
and U5646 (N_5646,N_5204,N_5167);
or U5647 (N_5647,N_5133,N_5371);
xnor U5648 (N_5648,N_5185,N_5378);
or U5649 (N_5649,N_5251,N_5344);
xnor U5650 (N_5650,N_5266,N_5129);
nor U5651 (N_5651,N_5195,N_5102);
and U5652 (N_5652,N_5153,N_5156);
nor U5653 (N_5653,N_5123,N_5242);
nand U5654 (N_5654,N_5108,N_5300);
xnor U5655 (N_5655,N_5146,N_5328);
nand U5656 (N_5656,N_5389,N_5216);
and U5657 (N_5657,N_5374,N_5262);
or U5658 (N_5658,N_5128,N_5317);
nand U5659 (N_5659,N_5289,N_5171);
nor U5660 (N_5660,N_5298,N_5361);
or U5661 (N_5661,N_5305,N_5364);
or U5662 (N_5662,N_5340,N_5287);
or U5663 (N_5663,N_5223,N_5262);
xor U5664 (N_5664,N_5143,N_5108);
nand U5665 (N_5665,N_5331,N_5211);
nor U5666 (N_5666,N_5275,N_5382);
nand U5667 (N_5667,N_5115,N_5295);
nand U5668 (N_5668,N_5195,N_5294);
or U5669 (N_5669,N_5345,N_5294);
xor U5670 (N_5670,N_5272,N_5127);
or U5671 (N_5671,N_5370,N_5105);
xor U5672 (N_5672,N_5173,N_5146);
or U5673 (N_5673,N_5288,N_5339);
and U5674 (N_5674,N_5101,N_5303);
nand U5675 (N_5675,N_5283,N_5394);
xor U5676 (N_5676,N_5171,N_5161);
and U5677 (N_5677,N_5199,N_5166);
and U5678 (N_5678,N_5208,N_5283);
and U5679 (N_5679,N_5302,N_5319);
nand U5680 (N_5680,N_5260,N_5163);
or U5681 (N_5681,N_5214,N_5173);
and U5682 (N_5682,N_5150,N_5157);
xor U5683 (N_5683,N_5352,N_5321);
nor U5684 (N_5684,N_5305,N_5114);
and U5685 (N_5685,N_5331,N_5215);
nor U5686 (N_5686,N_5277,N_5360);
xor U5687 (N_5687,N_5379,N_5353);
xnor U5688 (N_5688,N_5274,N_5346);
or U5689 (N_5689,N_5363,N_5327);
xor U5690 (N_5690,N_5291,N_5392);
nand U5691 (N_5691,N_5313,N_5295);
or U5692 (N_5692,N_5151,N_5191);
or U5693 (N_5693,N_5131,N_5382);
or U5694 (N_5694,N_5204,N_5128);
nand U5695 (N_5695,N_5150,N_5151);
and U5696 (N_5696,N_5160,N_5329);
or U5697 (N_5697,N_5270,N_5383);
nor U5698 (N_5698,N_5335,N_5298);
nor U5699 (N_5699,N_5195,N_5242);
or U5700 (N_5700,N_5639,N_5580);
nor U5701 (N_5701,N_5505,N_5583);
and U5702 (N_5702,N_5608,N_5551);
and U5703 (N_5703,N_5656,N_5582);
nand U5704 (N_5704,N_5662,N_5695);
and U5705 (N_5705,N_5464,N_5684);
nand U5706 (N_5706,N_5462,N_5453);
nand U5707 (N_5707,N_5439,N_5431);
or U5708 (N_5708,N_5641,N_5459);
nand U5709 (N_5709,N_5502,N_5491);
or U5710 (N_5710,N_5616,N_5541);
nor U5711 (N_5711,N_5496,N_5680);
nand U5712 (N_5712,N_5411,N_5460);
or U5713 (N_5713,N_5660,N_5487);
nand U5714 (N_5714,N_5628,N_5403);
or U5715 (N_5715,N_5685,N_5657);
and U5716 (N_5716,N_5558,N_5696);
and U5717 (N_5717,N_5532,N_5517);
nor U5718 (N_5718,N_5671,N_5678);
nor U5719 (N_5719,N_5446,N_5570);
nor U5720 (N_5720,N_5448,N_5699);
nor U5721 (N_5721,N_5621,N_5620);
nor U5722 (N_5722,N_5400,N_5412);
nor U5723 (N_5723,N_5474,N_5596);
nor U5724 (N_5724,N_5676,N_5625);
xor U5725 (N_5725,N_5447,N_5607);
nand U5726 (N_5726,N_5504,N_5690);
or U5727 (N_5727,N_5511,N_5594);
nor U5728 (N_5728,N_5408,N_5528);
or U5729 (N_5729,N_5575,N_5568);
xor U5730 (N_5730,N_5563,N_5689);
nand U5731 (N_5731,N_5544,N_5605);
nor U5732 (N_5732,N_5632,N_5651);
nor U5733 (N_5733,N_5434,N_5470);
nor U5734 (N_5734,N_5590,N_5424);
and U5735 (N_5735,N_5556,N_5486);
and U5736 (N_5736,N_5609,N_5546);
and U5737 (N_5737,N_5661,N_5539);
nand U5738 (N_5738,N_5573,N_5553);
nor U5739 (N_5739,N_5407,N_5577);
nor U5740 (N_5740,N_5510,N_5694);
and U5741 (N_5741,N_5449,N_5427);
and U5742 (N_5742,N_5451,N_5497);
and U5743 (N_5743,N_5418,N_5643);
nand U5744 (N_5744,N_5578,N_5697);
and U5745 (N_5745,N_5547,N_5428);
xor U5746 (N_5746,N_5457,N_5499);
or U5747 (N_5747,N_5549,N_5597);
or U5748 (N_5748,N_5581,N_5513);
and U5749 (N_5749,N_5498,N_5554);
nand U5750 (N_5750,N_5534,N_5598);
and U5751 (N_5751,N_5444,N_5617);
or U5752 (N_5752,N_5477,N_5409);
or U5753 (N_5753,N_5426,N_5530);
xnor U5754 (N_5754,N_5630,N_5698);
xor U5755 (N_5755,N_5545,N_5614);
and U5756 (N_5756,N_5509,N_5693);
and U5757 (N_5757,N_5592,N_5465);
nand U5758 (N_5758,N_5645,N_5619);
xnor U5759 (N_5759,N_5519,N_5673);
or U5760 (N_5760,N_5419,N_5672);
xor U5761 (N_5761,N_5623,N_5668);
or U5762 (N_5762,N_5537,N_5422);
or U5763 (N_5763,N_5461,N_5664);
and U5764 (N_5764,N_5515,N_5522);
or U5765 (N_5765,N_5479,N_5473);
nand U5766 (N_5766,N_5654,N_5529);
nor U5767 (N_5767,N_5591,N_5518);
xnor U5768 (N_5768,N_5501,N_5445);
and U5769 (N_5769,N_5599,N_5561);
nor U5770 (N_5770,N_5480,N_5482);
or U5771 (N_5771,N_5631,N_5681);
nor U5772 (N_5772,N_5593,N_5489);
xnor U5773 (N_5773,N_5441,N_5600);
nand U5774 (N_5774,N_5514,N_5548);
nand U5775 (N_5775,N_5533,N_5523);
nand U5776 (N_5776,N_5633,N_5521);
xnor U5777 (N_5777,N_5543,N_5435);
nand U5778 (N_5778,N_5567,N_5624);
and U5779 (N_5779,N_5443,N_5535);
nor U5780 (N_5780,N_5559,N_5669);
or U5781 (N_5781,N_5458,N_5610);
nor U5782 (N_5782,N_5503,N_5647);
nand U5783 (N_5783,N_5524,N_5478);
or U5784 (N_5784,N_5564,N_5469);
or U5785 (N_5785,N_5490,N_5508);
and U5786 (N_5786,N_5438,N_5601);
and U5787 (N_5787,N_5576,N_5674);
nand U5788 (N_5788,N_5436,N_5667);
and U5789 (N_5789,N_5562,N_5637);
xor U5790 (N_5790,N_5557,N_5655);
nand U5791 (N_5791,N_5440,N_5485);
nor U5792 (N_5792,N_5584,N_5542);
and U5793 (N_5793,N_5683,N_5626);
and U5794 (N_5794,N_5682,N_5467);
nand U5795 (N_5795,N_5423,N_5494);
xor U5796 (N_5796,N_5415,N_5405);
nand U5797 (N_5797,N_5500,N_5471);
and U5798 (N_5798,N_5615,N_5429);
nand U5799 (N_5799,N_5455,N_5606);
nor U5800 (N_5800,N_5538,N_5506);
nor U5801 (N_5801,N_5520,N_5579);
nor U5802 (N_5802,N_5468,N_5665);
and U5803 (N_5803,N_5613,N_5686);
or U5804 (N_5804,N_5492,N_5481);
xor U5805 (N_5805,N_5569,N_5466);
xnor U5806 (N_5806,N_5622,N_5574);
or U5807 (N_5807,N_5463,N_5475);
nand U5808 (N_5808,N_5536,N_5603);
or U5809 (N_5809,N_5653,N_5659);
or U5810 (N_5810,N_5618,N_5437);
xor U5811 (N_5811,N_5410,N_5646);
nor U5812 (N_5812,N_5452,N_5433);
or U5813 (N_5813,N_5611,N_5636);
and U5814 (N_5814,N_5414,N_5677);
xor U5815 (N_5815,N_5404,N_5692);
or U5816 (N_5816,N_5488,N_5663);
nand U5817 (N_5817,N_5572,N_5450);
nor U5818 (N_5818,N_5472,N_5687);
xor U5819 (N_5819,N_5602,N_5420);
nor U5820 (N_5820,N_5640,N_5526);
nor U5821 (N_5821,N_5666,N_5627);
nand U5822 (N_5822,N_5629,N_5442);
nor U5823 (N_5823,N_5516,N_5421);
nand U5824 (N_5824,N_5688,N_5652);
and U5825 (N_5825,N_5402,N_5507);
nand U5826 (N_5826,N_5454,N_5648);
xnor U5827 (N_5827,N_5691,N_5540);
nor U5828 (N_5828,N_5493,N_5644);
and U5829 (N_5829,N_5555,N_5585);
and U5830 (N_5830,N_5413,N_5586);
xor U5831 (N_5831,N_5416,N_5675);
or U5832 (N_5832,N_5531,N_5483);
nor U5833 (N_5833,N_5650,N_5525);
nor U5834 (N_5834,N_5456,N_5512);
xnor U5835 (N_5835,N_5560,N_5595);
xor U5836 (N_5836,N_5587,N_5670);
xor U5837 (N_5837,N_5432,N_5634);
and U5838 (N_5838,N_5638,N_5476);
and U5839 (N_5839,N_5527,N_5401);
nand U5840 (N_5840,N_5658,N_5571);
nand U5841 (N_5841,N_5649,N_5425);
and U5842 (N_5842,N_5588,N_5550);
or U5843 (N_5843,N_5484,N_5430);
xor U5844 (N_5844,N_5604,N_5589);
xnor U5845 (N_5845,N_5612,N_5417);
nor U5846 (N_5846,N_5406,N_5495);
nor U5847 (N_5847,N_5566,N_5552);
xor U5848 (N_5848,N_5635,N_5565);
or U5849 (N_5849,N_5642,N_5679);
and U5850 (N_5850,N_5504,N_5558);
nor U5851 (N_5851,N_5606,N_5490);
xor U5852 (N_5852,N_5541,N_5530);
or U5853 (N_5853,N_5583,N_5436);
nor U5854 (N_5854,N_5539,N_5571);
xnor U5855 (N_5855,N_5636,N_5447);
or U5856 (N_5856,N_5665,N_5660);
nand U5857 (N_5857,N_5676,N_5462);
nand U5858 (N_5858,N_5649,N_5572);
nor U5859 (N_5859,N_5674,N_5514);
xnor U5860 (N_5860,N_5683,N_5652);
and U5861 (N_5861,N_5646,N_5499);
xor U5862 (N_5862,N_5562,N_5418);
nor U5863 (N_5863,N_5634,N_5503);
nor U5864 (N_5864,N_5552,N_5417);
nor U5865 (N_5865,N_5480,N_5511);
xor U5866 (N_5866,N_5418,N_5547);
nand U5867 (N_5867,N_5538,N_5609);
nand U5868 (N_5868,N_5465,N_5454);
xnor U5869 (N_5869,N_5492,N_5408);
xnor U5870 (N_5870,N_5670,N_5400);
nand U5871 (N_5871,N_5519,N_5415);
nor U5872 (N_5872,N_5587,N_5539);
nand U5873 (N_5873,N_5636,N_5565);
or U5874 (N_5874,N_5659,N_5476);
or U5875 (N_5875,N_5464,N_5640);
nand U5876 (N_5876,N_5570,N_5615);
or U5877 (N_5877,N_5448,N_5487);
nand U5878 (N_5878,N_5627,N_5696);
or U5879 (N_5879,N_5485,N_5646);
and U5880 (N_5880,N_5483,N_5500);
and U5881 (N_5881,N_5404,N_5430);
nor U5882 (N_5882,N_5456,N_5652);
nor U5883 (N_5883,N_5646,N_5487);
and U5884 (N_5884,N_5537,N_5421);
xor U5885 (N_5885,N_5520,N_5686);
nand U5886 (N_5886,N_5493,N_5568);
and U5887 (N_5887,N_5557,N_5443);
nor U5888 (N_5888,N_5460,N_5688);
xnor U5889 (N_5889,N_5572,N_5563);
xor U5890 (N_5890,N_5567,N_5551);
or U5891 (N_5891,N_5438,N_5532);
nor U5892 (N_5892,N_5498,N_5530);
and U5893 (N_5893,N_5418,N_5697);
or U5894 (N_5894,N_5453,N_5666);
nor U5895 (N_5895,N_5530,N_5522);
nor U5896 (N_5896,N_5568,N_5512);
xor U5897 (N_5897,N_5601,N_5523);
nand U5898 (N_5898,N_5521,N_5457);
and U5899 (N_5899,N_5616,N_5536);
or U5900 (N_5900,N_5687,N_5498);
or U5901 (N_5901,N_5626,N_5484);
xor U5902 (N_5902,N_5590,N_5578);
and U5903 (N_5903,N_5574,N_5508);
nand U5904 (N_5904,N_5507,N_5610);
nor U5905 (N_5905,N_5525,N_5598);
nor U5906 (N_5906,N_5672,N_5538);
nor U5907 (N_5907,N_5696,N_5479);
nand U5908 (N_5908,N_5442,N_5473);
xnor U5909 (N_5909,N_5435,N_5496);
xor U5910 (N_5910,N_5689,N_5529);
nor U5911 (N_5911,N_5416,N_5669);
and U5912 (N_5912,N_5476,N_5446);
and U5913 (N_5913,N_5546,N_5588);
and U5914 (N_5914,N_5606,N_5569);
or U5915 (N_5915,N_5580,N_5679);
and U5916 (N_5916,N_5442,N_5512);
nand U5917 (N_5917,N_5521,N_5537);
and U5918 (N_5918,N_5419,N_5484);
and U5919 (N_5919,N_5461,N_5656);
and U5920 (N_5920,N_5685,N_5686);
or U5921 (N_5921,N_5562,N_5676);
and U5922 (N_5922,N_5686,N_5561);
and U5923 (N_5923,N_5636,N_5533);
or U5924 (N_5924,N_5411,N_5632);
or U5925 (N_5925,N_5467,N_5410);
nor U5926 (N_5926,N_5484,N_5513);
and U5927 (N_5927,N_5591,N_5443);
xnor U5928 (N_5928,N_5479,N_5512);
or U5929 (N_5929,N_5460,N_5556);
xnor U5930 (N_5930,N_5410,N_5641);
or U5931 (N_5931,N_5512,N_5551);
or U5932 (N_5932,N_5553,N_5546);
and U5933 (N_5933,N_5642,N_5488);
and U5934 (N_5934,N_5559,N_5484);
and U5935 (N_5935,N_5604,N_5431);
nand U5936 (N_5936,N_5496,N_5623);
or U5937 (N_5937,N_5618,N_5597);
nand U5938 (N_5938,N_5481,N_5462);
nand U5939 (N_5939,N_5454,N_5443);
xnor U5940 (N_5940,N_5674,N_5688);
nor U5941 (N_5941,N_5591,N_5673);
nor U5942 (N_5942,N_5577,N_5605);
nor U5943 (N_5943,N_5590,N_5645);
nor U5944 (N_5944,N_5592,N_5482);
or U5945 (N_5945,N_5495,N_5582);
nand U5946 (N_5946,N_5475,N_5438);
nor U5947 (N_5947,N_5546,N_5593);
nor U5948 (N_5948,N_5538,N_5414);
nand U5949 (N_5949,N_5608,N_5584);
nand U5950 (N_5950,N_5481,N_5512);
nor U5951 (N_5951,N_5607,N_5676);
or U5952 (N_5952,N_5503,N_5461);
nand U5953 (N_5953,N_5518,N_5418);
xnor U5954 (N_5954,N_5681,N_5523);
nor U5955 (N_5955,N_5512,N_5491);
and U5956 (N_5956,N_5601,N_5441);
xnor U5957 (N_5957,N_5615,N_5618);
or U5958 (N_5958,N_5621,N_5593);
and U5959 (N_5959,N_5649,N_5691);
and U5960 (N_5960,N_5416,N_5630);
nand U5961 (N_5961,N_5404,N_5558);
and U5962 (N_5962,N_5698,N_5444);
or U5963 (N_5963,N_5513,N_5551);
xor U5964 (N_5964,N_5491,N_5646);
nand U5965 (N_5965,N_5616,N_5429);
xnor U5966 (N_5966,N_5433,N_5629);
nor U5967 (N_5967,N_5544,N_5476);
or U5968 (N_5968,N_5614,N_5593);
xnor U5969 (N_5969,N_5608,N_5508);
nand U5970 (N_5970,N_5677,N_5549);
nand U5971 (N_5971,N_5634,N_5487);
nor U5972 (N_5972,N_5668,N_5457);
nor U5973 (N_5973,N_5602,N_5444);
and U5974 (N_5974,N_5629,N_5455);
and U5975 (N_5975,N_5610,N_5493);
nand U5976 (N_5976,N_5519,N_5459);
xor U5977 (N_5977,N_5571,N_5538);
and U5978 (N_5978,N_5632,N_5471);
xnor U5979 (N_5979,N_5600,N_5606);
nand U5980 (N_5980,N_5556,N_5547);
nor U5981 (N_5981,N_5691,N_5631);
nand U5982 (N_5982,N_5688,N_5482);
nor U5983 (N_5983,N_5608,N_5428);
nand U5984 (N_5984,N_5516,N_5509);
and U5985 (N_5985,N_5409,N_5472);
and U5986 (N_5986,N_5572,N_5533);
or U5987 (N_5987,N_5525,N_5594);
xnor U5988 (N_5988,N_5616,N_5475);
nor U5989 (N_5989,N_5614,N_5669);
nor U5990 (N_5990,N_5660,N_5470);
and U5991 (N_5991,N_5477,N_5475);
or U5992 (N_5992,N_5446,N_5450);
nor U5993 (N_5993,N_5470,N_5452);
nor U5994 (N_5994,N_5600,N_5446);
nor U5995 (N_5995,N_5644,N_5538);
xnor U5996 (N_5996,N_5428,N_5486);
xnor U5997 (N_5997,N_5516,N_5497);
xor U5998 (N_5998,N_5565,N_5527);
nand U5999 (N_5999,N_5424,N_5476);
or U6000 (N_6000,N_5945,N_5810);
or U6001 (N_6001,N_5720,N_5886);
and U6002 (N_6002,N_5837,N_5982);
or U6003 (N_6003,N_5955,N_5890);
xnor U6004 (N_6004,N_5996,N_5828);
and U6005 (N_6005,N_5781,N_5752);
nor U6006 (N_6006,N_5899,N_5873);
or U6007 (N_6007,N_5824,N_5746);
or U6008 (N_6008,N_5999,N_5813);
and U6009 (N_6009,N_5965,N_5950);
nand U6010 (N_6010,N_5845,N_5758);
xor U6011 (N_6011,N_5876,N_5714);
nand U6012 (N_6012,N_5862,N_5869);
xnor U6013 (N_6013,N_5737,N_5958);
xnor U6014 (N_6014,N_5860,N_5791);
xnor U6015 (N_6015,N_5794,N_5902);
nand U6016 (N_6016,N_5855,N_5966);
nor U6017 (N_6017,N_5983,N_5708);
and U6018 (N_6018,N_5974,N_5948);
nor U6019 (N_6019,N_5935,N_5921);
nor U6020 (N_6020,N_5814,N_5911);
xor U6021 (N_6021,N_5721,N_5884);
nand U6022 (N_6022,N_5887,N_5874);
and U6023 (N_6023,N_5780,N_5970);
nor U6024 (N_6024,N_5733,N_5768);
xor U6025 (N_6025,N_5798,N_5909);
and U6026 (N_6026,N_5701,N_5782);
nor U6027 (N_6027,N_5880,N_5809);
nor U6028 (N_6028,N_5981,N_5994);
nand U6029 (N_6029,N_5846,N_5932);
nand U6030 (N_6030,N_5826,N_5971);
nor U6031 (N_6031,N_5803,N_5934);
or U6032 (N_6032,N_5872,N_5764);
nand U6033 (N_6033,N_5787,N_5953);
nor U6034 (N_6034,N_5849,N_5906);
or U6035 (N_6035,N_5933,N_5741);
xnor U6036 (N_6036,N_5841,N_5865);
xnor U6037 (N_6037,N_5829,N_5986);
xnor U6038 (N_6038,N_5804,N_5875);
nand U6039 (N_6039,N_5770,N_5785);
or U6040 (N_6040,N_5928,N_5738);
nor U6041 (N_6041,N_5918,N_5942);
nor U6042 (N_6042,N_5844,N_5892);
nand U6043 (N_6043,N_5894,N_5867);
xnor U6044 (N_6044,N_5774,N_5743);
or U6045 (N_6045,N_5730,N_5938);
nand U6046 (N_6046,N_5960,N_5987);
nor U6047 (N_6047,N_5985,N_5812);
xor U6048 (N_6048,N_5757,N_5700);
and U6049 (N_6049,N_5946,N_5908);
and U6050 (N_6050,N_5724,N_5717);
nor U6051 (N_6051,N_5795,N_5786);
or U6052 (N_6052,N_5761,N_5889);
or U6053 (N_6053,N_5788,N_5878);
nor U6054 (N_6054,N_5951,N_5759);
or U6055 (N_6055,N_5995,N_5883);
and U6056 (N_6056,N_5926,N_5962);
or U6057 (N_6057,N_5895,N_5710);
and U6058 (N_6058,N_5992,N_5838);
xor U6059 (N_6059,N_5858,N_5704);
nand U6060 (N_6060,N_5832,N_5818);
or U6061 (N_6061,N_5972,N_5968);
and U6062 (N_6062,N_5997,N_5731);
and U6063 (N_6063,N_5879,N_5913);
nand U6064 (N_6064,N_5796,N_5989);
nor U6065 (N_6065,N_5919,N_5922);
or U6066 (N_6066,N_5726,N_5808);
or U6067 (N_6067,N_5760,N_5949);
nand U6068 (N_6068,N_5920,N_5973);
and U6069 (N_6069,N_5707,N_5712);
nand U6070 (N_6070,N_5929,N_5825);
or U6071 (N_6071,N_5854,N_5917);
or U6072 (N_6072,N_5963,N_5939);
or U6073 (N_6073,N_5871,N_5961);
nand U6074 (N_6074,N_5771,N_5891);
nand U6075 (N_6075,N_5836,N_5923);
or U6076 (N_6076,N_5705,N_5772);
and U6077 (N_6077,N_5975,N_5900);
xnor U6078 (N_6078,N_5840,N_5993);
nor U6079 (N_6079,N_5978,N_5801);
xnor U6080 (N_6080,N_5776,N_5967);
or U6081 (N_6081,N_5979,N_5756);
xor U6082 (N_6082,N_5936,N_5976);
xnor U6083 (N_6083,N_5819,N_5893);
nor U6084 (N_6084,N_5784,N_5722);
or U6085 (N_6085,N_5751,N_5745);
or U6086 (N_6086,N_5903,N_5842);
xnor U6087 (N_6087,N_5897,N_5943);
or U6088 (N_6088,N_5988,N_5910);
nand U6089 (N_6089,N_5767,N_5739);
nor U6090 (N_6090,N_5898,N_5940);
nand U6091 (N_6091,N_5885,N_5853);
and U6092 (N_6092,N_5980,N_5789);
xnor U6093 (N_6093,N_5927,N_5916);
or U6094 (N_6094,N_5896,N_5792);
nor U6095 (N_6095,N_5777,N_5850);
or U6096 (N_6096,N_5969,N_5740);
and U6097 (N_6097,N_5835,N_5715);
and U6098 (N_6098,N_5706,N_5870);
or U6099 (N_6099,N_5763,N_5834);
or U6100 (N_6100,N_5852,N_5881);
nor U6101 (N_6101,N_5831,N_5959);
xor U6102 (N_6102,N_5930,N_5747);
nor U6103 (N_6103,N_5817,N_5843);
nand U6104 (N_6104,N_5947,N_5823);
xnor U6105 (N_6105,N_5857,N_5742);
nor U6106 (N_6106,N_5944,N_5713);
nand U6107 (N_6107,N_5822,N_5991);
or U6108 (N_6108,N_5790,N_5877);
and U6109 (N_6109,N_5778,N_5709);
nor U6110 (N_6110,N_5851,N_5866);
xnor U6111 (N_6111,N_5732,N_5748);
and U6112 (N_6112,N_5863,N_5816);
xnor U6113 (N_6113,N_5802,N_5749);
and U6114 (N_6114,N_5806,N_5769);
or U6115 (N_6115,N_5901,N_5703);
nor U6116 (N_6116,N_5762,N_5848);
and U6117 (N_6117,N_5727,N_5723);
nand U6118 (N_6118,N_5716,N_5905);
xor U6119 (N_6119,N_5779,N_5775);
or U6120 (N_6120,N_5977,N_5800);
nand U6121 (N_6121,N_5839,N_5937);
or U6122 (N_6122,N_5998,N_5755);
and U6123 (N_6123,N_5957,N_5734);
xnor U6124 (N_6124,N_5736,N_5754);
nand U6125 (N_6125,N_5805,N_5833);
nand U6126 (N_6126,N_5793,N_5956);
and U6127 (N_6127,N_5904,N_5859);
nor U6128 (N_6128,N_5868,N_5912);
xnor U6129 (N_6129,N_5766,N_5924);
xnor U6130 (N_6130,N_5750,N_5882);
nand U6131 (N_6131,N_5711,N_5807);
and U6132 (N_6132,N_5931,N_5914);
nor U6133 (N_6133,N_5864,N_5861);
xor U6134 (N_6134,N_5915,N_5735);
xor U6135 (N_6135,N_5952,N_5719);
and U6136 (N_6136,N_5827,N_5925);
nand U6137 (N_6137,N_5820,N_5765);
or U6138 (N_6138,N_5954,N_5811);
nor U6139 (N_6139,N_5847,N_5964);
or U6140 (N_6140,N_5729,N_5744);
nor U6141 (N_6141,N_5888,N_5830);
or U6142 (N_6142,N_5941,N_5984);
xnor U6143 (N_6143,N_5753,N_5725);
xor U6144 (N_6144,N_5728,N_5773);
or U6145 (N_6145,N_5990,N_5907);
nor U6146 (N_6146,N_5815,N_5821);
xnor U6147 (N_6147,N_5783,N_5797);
or U6148 (N_6148,N_5718,N_5702);
nor U6149 (N_6149,N_5856,N_5799);
or U6150 (N_6150,N_5727,N_5869);
nand U6151 (N_6151,N_5982,N_5782);
or U6152 (N_6152,N_5963,N_5826);
or U6153 (N_6153,N_5735,N_5999);
and U6154 (N_6154,N_5933,N_5951);
or U6155 (N_6155,N_5876,N_5829);
xor U6156 (N_6156,N_5810,N_5977);
or U6157 (N_6157,N_5769,N_5966);
xor U6158 (N_6158,N_5766,N_5746);
nand U6159 (N_6159,N_5971,N_5732);
and U6160 (N_6160,N_5881,N_5860);
nand U6161 (N_6161,N_5804,N_5876);
xor U6162 (N_6162,N_5925,N_5829);
xnor U6163 (N_6163,N_5818,N_5824);
nor U6164 (N_6164,N_5947,N_5970);
nor U6165 (N_6165,N_5911,N_5915);
xnor U6166 (N_6166,N_5993,N_5988);
and U6167 (N_6167,N_5871,N_5793);
nor U6168 (N_6168,N_5877,N_5788);
nor U6169 (N_6169,N_5981,N_5855);
and U6170 (N_6170,N_5858,N_5866);
and U6171 (N_6171,N_5795,N_5790);
and U6172 (N_6172,N_5984,N_5872);
xor U6173 (N_6173,N_5974,N_5767);
nor U6174 (N_6174,N_5842,N_5844);
nor U6175 (N_6175,N_5831,N_5768);
xor U6176 (N_6176,N_5743,N_5746);
xor U6177 (N_6177,N_5735,N_5953);
nor U6178 (N_6178,N_5823,N_5921);
or U6179 (N_6179,N_5863,N_5763);
nand U6180 (N_6180,N_5914,N_5959);
xor U6181 (N_6181,N_5891,N_5883);
and U6182 (N_6182,N_5924,N_5919);
and U6183 (N_6183,N_5932,N_5763);
nand U6184 (N_6184,N_5847,N_5967);
or U6185 (N_6185,N_5831,N_5811);
and U6186 (N_6186,N_5700,N_5791);
nand U6187 (N_6187,N_5831,N_5838);
and U6188 (N_6188,N_5733,N_5717);
xnor U6189 (N_6189,N_5958,N_5700);
nor U6190 (N_6190,N_5902,N_5946);
nor U6191 (N_6191,N_5910,N_5798);
and U6192 (N_6192,N_5934,N_5835);
or U6193 (N_6193,N_5769,N_5997);
xnor U6194 (N_6194,N_5877,N_5757);
nor U6195 (N_6195,N_5791,N_5893);
nor U6196 (N_6196,N_5954,N_5837);
or U6197 (N_6197,N_5785,N_5886);
xnor U6198 (N_6198,N_5703,N_5834);
and U6199 (N_6199,N_5998,N_5912);
nand U6200 (N_6200,N_5806,N_5996);
and U6201 (N_6201,N_5926,N_5964);
or U6202 (N_6202,N_5754,N_5750);
nand U6203 (N_6203,N_5801,N_5845);
nor U6204 (N_6204,N_5937,N_5916);
nand U6205 (N_6205,N_5892,N_5912);
nor U6206 (N_6206,N_5959,N_5759);
and U6207 (N_6207,N_5758,N_5937);
xor U6208 (N_6208,N_5753,N_5813);
nor U6209 (N_6209,N_5747,N_5720);
and U6210 (N_6210,N_5980,N_5949);
nor U6211 (N_6211,N_5707,N_5842);
nor U6212 (N_6212,N_5967,N_5851);
and U6213 (N_6213,N_5879,N_5911);
or U6214 (N_6214,N_5838,N_5840);
nor U6215 (N_6215,N_5739,N_5983);
nand U6216 (N_6216,N_5916,N_5788);
and U6217 (N_6217,N_5865,N_5947);
or U6218 (N_6218,N_5908,N_5897);
nand U6219 (N_6219,N_5715,N_5933);
and U6220 (N_6220,N_5831,N_5975);
nor U6221 (N_6221,N_5775,N_5865);
nand U6222 (N_6222,N_5756,N_5899);
nor U6223 (N_6223,N_5817,N_5765);
and U6224 (N_6224,N_5737,N_5972);
and U6225 (N_6225,N_5838,N_5850);
nor U6226 (N_6226,N_5929,N_5839);
nor U6227 (N_6227,N_5905,N_5973);
xnor U6228 (N_6228,N_5875,N_5860);
nor U6229 (N_6229,N_5752,N_5760);
and U6230 (N_6230,N_5861,N_5927);
and U6231 (N_6231,N_5702,N_5996);
nor U6232 (N_6232,N_5898,N_5778);
and U6233 (N_6233,N_5772,N_5958);
nand U6234 (N_6234,N_5911,N_5909);
nor U6235 (N_6235,N_5896,N_5987);
nor U6236 (N_6236,N_5744,N_5852);
xor U6237 (N_6237,N_5962,N_5915);
or U6238 (N_6238,N_5768,N_5726);
xnor U6239 (N_6239,N_5822,N_5941);
nand U6240 (N_6240,N_5747,N_5934);
xnor U6241 (N_6241,N_5703,N_5877);
or U6242 (N_6242,N_5815,N_5932);
nor U6243 (N_6243,N_5802,N_5773);
and U6244 (N_6244,N_5989,N_5801);
and U6245 (N_6245,N_5867,N_5759);
and U6246 (N_6246,N_5738,N_5885);
xnor U6247 (N_6247,N_5826,N_5970);
and U6248 (N_6248,N_5990,N_5861);
xor U6249 (N_6249,N_5727,N_5855);
or U6250 (N_6250,N_5729,N_5941);
nor U6251 (N_6251,N_5998,N_5928);
or U6252 (N_6252,N_5889,N_5903);
xnor U6253 (N_6253,N_5766,N_5826);
xor U6254 (N_6254,N_5993,N_5745);
xnor U6255 (N_6255,N_5778,N_5807);
or U6256 (N_6256,N_5813,N_5815);
nor U6257 (N_6257,N_5995,N_5807);
nand U6258 (N_6258,N_5893,N_5792);
or U6259 (N_6259,N_5971,N_5799);
nor U6260 (N_6260,N_5927,N_5952);
and U6261 (N_6261,N_5724,N_5855);
xor U6262 (N_6262,N_5806,N_5894);
nand U6263 (N_6263,N_5855,N_5712);
nand U6264 (N_6264,N_5779,N_5979);
or U6265 (N_6265,N_5983,N_5926);
xor U6266 (N_6266,N_5885,N_5777);
nor U6267 (N_6267,N_5972,N_5731);
and U6268 (N_6268,N_5822,N_5881);
or U6269 (N_6269,N_5861,N_5903);
xor U6270 (N_6270,N_5708,N_5947);
xor U6271 (N_6271,N_5959,N_5920);
nor U6272 (N_6272,N_5890,N_5907);
and U6273 (N_6273,N_5800,N_5949);
nand U6274 (N_6274,N_5731,N_5713);
nand U6275 (N_6275,N_5714,N_5742);
and U6276 (N_6276,N_5717,N_5837);
nor U6277 (N_6277,N_5807,N_5727);
nand U6278 (N_6278,N_5836,N_5718);
and U6279 (N_6279,N_5739,N_5751);
nor U6280 (N_6280,N_5765,N_5752);
nor U6281 (N_6281,N_5951,N_5750);
and U6282 (N_6282,N_5994,N_5709);
xnor U6283 (N_6283,N_5917,N_5726);
or U6284 (N_6284,N_5779,N_5763);
nor U6285 (N_6285,N_5974,N_5787);
and U6286 (N_6286,N_5972,N_5738);
or U6287 (N_6287,N_5798,N_5720);
nand U6288 (N_6288,N_5997,N_5987);
xnor U6289 (N_6289,N_5992,N_5873);
nor U6290 (N_6290,N_5987,N_5797);
and U6291 (N_6291,N_5705,N_5879);
nor U6292 (N_6292,N_5912,N_5878);
or U6293 (N_6293,N_5887,N_5762);
and U6294 (N_6294,N_5712,N_5737);
and U6295 (N_6295,N_5864,N_5781);
and U6296 (N_6296,N_5911,N_5872);
nand U6297 (N_6297,N_5918,N_5790);
and U6298 (N_6298,N_5754,N_5972);
and U6299 (N_6299,N_5804,N_5838);
nand U6300 (N_6300,N_6048,N_6165);
or U6301 (N_6301,N_6085,N_6279);
nand U6302 (N_6302,N_6275,N_6025);
nand U6303 (N_6303,N_6122,N_6169);
nor U6304 (N_6304,N_6128,N_6217);
nand U6305 (N_6305,N_6102,N_6298);
or U6306 (N_6306,N_6182,N_6192);
or U6307 (N_6307,N_6181,N_6117);
xnor U6308 (N_6308,N_6155,N_6129);
nor U6309 (N_6309,N_6009,N_6259);
and U6310 (N_6310,N_6133,N_6072);
or U6311 (N_6311,N_6067,N_6290);
and U6312 (N_6312,N_6171,N_6112);
nor U6313 (N_6313,N_6212,N_6091);
xor U6314 (N_6314,N_6017,N_6191);
xor U6315 (N_6315,N_6105,N_6253);
and U6316 (N_6316,N_6127,N_6119);
nand U6317 (N_6317,N_6106,N_6077);
and U6318 (N_6318,N_6222,N_6226);
or U6319 (N_6319,N_6244,N_6052);
or U6320 (N_6320,N_6154,N_6096);
nor U6321 (N_6321,N_6076,N_6138);
or U6322 (N_6322,N_6124,N_6135);
and U6323 (N_6323,N_6250,N_6002);
nor U6324 (N_6324,N_6203,N_6208);
xnor U6325 (N_6325,N_6199,N_6287);
or U6326 (N_6326,N_6243,N_6115);
nor U6327 (N_6327,N_6121,N_6209);
nor U6328 (N_6328,N_6031,N_6104);
nand U6329 (N_6329,N_6254,N_6190);
and U6330 (N_6330,N_6123,N_6299);
and U6331 (N_6331,N_6198,N_6225);
or U6332 (N_6332,N_6200,N_6255);
xnor U6333 (N_6333,N_6189,N_6173);
nor U6334 (N_6334,N_6187,N_6204);
and U6335 (N_6335,N_6042,N_6266);
or U6336 (N_6336,N_6248,N_6185);
xor U6337 (N_6337,N_6053,N_6224);
xor U6338 (N_6338,N_6110,N_6281);
nor U6339 (N_6339,N_6016,N_6295);
or U6340 (N_6340,N_6120,N_6000);
and U6341 (N_6341,N_6062,N_6152);
and U6342 (N_6342,N_6214,N_6088);
and U6343 (N_6343,N_6178,N_6147);
or U6344 (N_6344,N_6058,N_6194);
nor U6345 (N_6345,N_6164,N_6113);
nand U6346 (N_6346,N_6028,N_6068);
nor U6347 (N_6347,N_6261,N_6294);
nor U6348 (N_6348,N_6007,N_6297);
xor U6349 (N_6349,N_6083,N_6219);
and U6350 (N_6350,N_6196,N_6246);
xnor U6351 (N_6351,N_6131,N_6267);
or U6352 (N_6352,N_6015,N_6293);
xor U6353 (N_6353,N_6235,N_6086);
or U6354 (N_6354,N_6288,N_6159);
nor U6355 (N_6355,N_6276,N_6089);
and U6356 (N_6356,N_6056,N_6220);
nor U6357 (N_6357,N_6065,N_6045);
nand U6358 (N_6358,N_6073,N_6040);
or U6359 (N_6359,N_6139,N_6251);
xor U6360 (N_6360,N_6280,N_6075);
nand U6361 (N_6361,N_6237,N_6061);
nand U6362 (N_6362,N_6082,N_6114);
and U6363 (N_6363,N_6006,N_6084);
or U6364 (N_6364,N_6232,N_6118);
nand U6365 (N_6365,N_6050,N_6183);
and U6366 (N_6366,N_6223,N_6146);
or U6367 (N_6367,N_6066,N_6210);
nor U6368 (N_6368,N_6109,N_6140);
or U6369 (N_6369,N_6010,N_6013);
nand U6370 (N_6370,N_6111,N_6206);
or U6371 (N_6371,N_6236,N_6218);
nor U6372 (N_6372,N_6263,N_6060);
or U6373 (N_6373,N_6260,N_6024);
and U6374 (N_6374,N_6292,N_6238);
or U6375 (N_6375,N_6230,N_6043);
nor U6376 (N_6376,N_6240,N_6074);
nor U6377 (N_6377,N_6285,N_6020);
nand U6378 (N_6378,N_6273,N_6151);
nor U6379 (N_6379,N_6262,N_6229);
xor U6380 (N_6380,N_6160,N_6247);
xnor U6381 (N_6381,N_6213,N_6033);
and U6382 (N_6382,N_6107,N_6195);
and U6383 (N_6383,N_6272,N_6277);
nor U6384 (N_6384,N_6079,N_6184);
nand U6385 (N_6385,N_6274,N_6282);
nor U6386 (N_6386,N_6047,N_6141);
xor U6387 (N_6387,N_6063,N_6202);
or U6388 (N_6388,N_6049,N_6039);
nand U6389 (N_6389,N_6090,N_6116);
nand U6390 (N_6390,N_6098,N_6142);
nand U6391 (N_6391,N_6021,N_6207);
nor U6392 (N_6392,N_6044,N_6046);
and U6393 (N_6393,N_6051,N_6150);
nor U6394 (N_6394,N_6080,N_6228);
and U6395 (N_6395,N_6180,N_6161);
nand U6396 (N_6396,N_6215,N_6071);
and U6397 (N_6397,N_6144,N_6162);
or U6398 (N_6398,N_6001,N_6099);
xor U6399 (N_6399,N_6069,N_6163);
nor U6400 (N_6400,N_6172,N_6003);
and U6401 (N_6401,N_6221,N_6241);
and U6402 (N_6402,N_6291,N_6100);
and U6403 (N_6403,N_6023,N_6059);
or U6404 (N_6404,N_6004,N_6137);
and U6405 (N_6405,N_6136,N_6087);
nand U6406 (N_6406,N_6174,N_6036);
xnor U6407 (N_6407,N_6242,N_6038);
xnor U6408 (N_6408,N_6097,N_6108);
or U6409 (N_6409,N_6078,N_6132);
and U6410 (N_6410,N_6256,N_6216);
xor U6411 (N_6411,N_6064,N_6027);
xor U6412 (N_6412,N_6081,N_6030);
and U6413 (N_6413,N_6249,N_6041);
nand U6414 (N_6414,N_6070,N_6026);
nor U6415 (N_6415,N_6166,N_6130);
nor U6416 (N_6416,N_6018,N_6193);
nor U6417 (N_6417,N_6035,N_6179);
and U6418 (N_6418,N_6265,N_6205);
or U6419 (N_6419,N_6158,N_6157);
nand U6420 (N_6420,N_6264,N_6126);
nand U6421 (N_6421,N_6055,N_6156);
nand U6422 (N_6422,N_6008,N_6168);
and U6423 (N_6423,N_6257,N_6170);
or U6424 (N_6424,N_6012,N_6188);
and U6425 (N_6425,N_6103,N_6145);
nor U6426 (N_6426,N_6092,N_6153);
nor U6427 (N_6427,N_6177,N_6283);
xnor U6428 (N_6428,N_6289,N_6148);
and U6429 (N_6429,N_6034,N_6197);
xor U6430 (N_6430,N_6278,N_6271);
nor U6431 (N_6431,N_6233,N_6286);
or U6432 (N_6432,N_6057,N_6054);
and U6433 (N_6433,N_6134,N_6037);
or U6434 (N_6434,N_6234,N_6245);
and U6435 (N_6435,N_6296,N_6252);
xnor U6436 (N_6436,N_6143,N_6149);
nand U6437 (N_6437,N_6101,N_6011);
or U6438 (N_6438,N_6125,N_6176);
xnor U6439 (N_6439,N_6032,N_6268);
and U6440 (N_6440,N_6258,N_6231);
nor U6441 (N_6441,N_6094,N_6019);
and U6442 (N_6442,N_6227,N_6211);
nand U6443 (N_6443,N_6201,N_6186);
xor U6444 (N_6444,N_6269,N_6014);
xnor U6445 (N_6445,N_6095,N_6005);
nand U6446 (N_6446,N_6093,N_6022);
xnor U6447 (N_6447,N_6175,N_6284);
nor U6448 (N_6448,N_6239,N_6167);
nand U6449 (N_6449,N_6270,N_6029);
or U6450 (N_6450,N_6279,N_6088);
xor U6451 (N_6451,N_6184,N_6205);
nand U6452 (N_6452,N_6020,N_6145);
xnor U6453 (N_6453,N_6158,N_6239);
and U6454 (N_6454,N_6224,N_6061);
nand U6455 (N_6455,N_6202,N_6168);
and U6456 (N_6456,N_6127,N_6017);
nand U6457 (N_6457,N_6277,N_6083);
or U6458 (N_6458,N_6272,N_6182);
nand U6459 (N_6459,N_6000,N_6256);
or U6460 (N_6460,N_6199,N_6119);
or U6461 (N_6461,N_6006,N_6111);
and U6462 (N_6462,N_6061,N_6274);
and U6463 (N_6463,N_6183,N_6005);
nand U6464 (N_6464,N_6137,N_6224);
or U6465 (N_6465,N_6271,N_6050);
xor U6466 (N_6466,N_6165,N_6247);
and U6467 (N_6467,N_6016,N_6061);
nand U6468 (N_6468,N_6258,N_6284);
xor U6469 (N_6469,N_6236,N_6041);
or U6470 (N_6470,N_6126,N_6232);
and U6471 (N_6471,N_6240,N_6149);
or U6472 (N_6472,N_6100,N_6069);
xor U6473 (N_6473,N_6233,N_6069);
and U6474 (N_6474,N_6250,N_6121);
xnor U6475 (N_6475,N_6016,N_6067);
xnor U6476 (N_6476,N_6211,N_6095);
nand U6477 (N_6477,N_6260,N_6273);
xor U6478 (N_6478,N_6099,N_6290);
or U6479 (N_6479,N_6095,N_6099);
and U6480 (N_6480,N_6202,N_6169);
and U6481 (N_6481,N_6252,N_6227);
and U6482 (N_6482,N_6046,N_6113);
or U6483 (N_6483,N_6260,N_6278);
or U6484 (N_6484,N_6211,N_6166);
or U6485 (N_6485,N_6195,N_6139);
nor U6486 (N_6486,N_6032,N_6274);
and U6487 (N_6487,N_6214,N_6157);
xor U6488 (N_6488,N_6156,N_6136);
nand U6489 (N_6489,N_6054,N_6138);
xor U6490 (N_6490,N_6130,N_6242);
and U6491 (N_6491,N_6113,N_6292);
or U6492 (N_6492,N_6281,N_6041);
nand U6493 (N_6493,N_6003,N_6162);
nand U6494 (N_6494,N_6245,N_6179);
nand U6495 (N_6495,N_6259,N_6275);
nand U6496 (N_6496,N_6229,N_6293);
xnor U6497 (N_6497,N_6066,N_6203);
nand U6498 (N_6498,N_6225,N_6084);
or U6499 (N_6499,N_6115,N_6059);
xnor U6500 (N_6500,N_6091,N_6026);
nand U6501 (N_6501,N_6102,N_6271);
or U6502 (N_6502,N_6157,N_6013);
and U6503 (N_6503,N_6226,N_6200);
and U6504 (N_6504,N_6117,N_6269);
nor U6505 (N_6505,N_6038,N_6019);
nor U6506 (N_6506,N_6135,N_6264);
and U6507 (N_6507,N_6156,N_6286);
nand U6508 (N_6508,N_6117,N_6141);
xor U6509 (N_6509,N_6151,N_6271);
nand U6510 (N_6510,N_6264,N_6143);
and U6511 (N_6511,N_6047,N_6082);
and U6512 (N_6512,N_6119,N_6072);
or U6513 (N_6513,N_6082,N_6074);
and U6514 (N_6514,N_6178,N_6243);
xnor U6515 (N_6515,N_6062,N_6143);
nand U6516 (N_6516,N_6066,N_6124);
and U6517 (N_6517,N_6292,N_6284);
nor U6518 (N_6518,N_6070,N_6240);
nor U6519 (N_6519,N_6291,N_6063);
nor U6520 (N_6520,N_6166,N_6160);
or U6521 (N_6521,N_6202,N_6224);
nor U6522 (N_6522,N_6252,N_6186);
nor U6523 (N_6523,N_6094,N_6249);
or U6524 (N_6524,N_6212,N_6207);
and U6525 (N_6525,N_6270,N_6239);
or U6526 (N_6526,N_6217,N_6132);
nand U6527 (N_6527,N_6216,N_6188);
xor U6528 (N_6528,N_6158,N_6052);
nor U6529 (N_6529,N_6293,N_6074);
and U6530 (N_6530,N_6238,N_6149);
and U6531 (N_6531,N_6275,N_6138);
nand U6532 (N_6532,N_6257,N_6011);
nand U6533 (N_6533,N_6255,N_6296);
nand U6534 (N_6534,N_6052,N_6018);
or U6535 (N_6535,N_6284,N_6179);
nor U6536 (N_6536,N_6038,N_6072);
nand U6537 (N_6537,N_6014,N_6265);
or U6538 (N_6538,N_6089,N_6247);
xnor U6539 (N_6539,N_6006,N_6177);
and U6540 (N_6540,N_6181,N_6173);
nand U6541 (N_6541,N_6118,N_6234);
nand U6542 (N_6542,N_6010,N_6026);
nand U6543 (N_6543,N_6258,N_6150);
and U6544 (N_6544,N_6192,N_6231);
nand U6545 (N_6545,N_6036,N_6027);
nor U6546 (N_6546,N_6120,N_6128);
and U6547 (N_6547,N_6065,N_6129);
xnor U6548 (N_6548,N_6155,N_6259);
and U6549 (N_6549,N_6165,N_6028);
nor U6550 (N_6550,N_6171,N_6034);
or U6551 (N_6551,N_6023,N_6036);
xor U6552 (N_6552,N_6178,N_6217);
or U6553 (N_6553,N_6227,N_6262);
nand U6554 (N_6554,N_6001,N_6202);
xor U6555 (N_6555,N_6158,N_6107);
xor U6556 (N_6556,N_6212,N_6266);
nand U6557 (N_6557,N_6061,N_6065);
nand U6558 (N_6558,N_6012,N_6293);
xor U6559 (N_6559,N_6091,N_6004);
xor U6560 (N_6560,N_6100,N_6171);
nor U6561 (N_6561,N_6126,N_6054);
or U6562 (N_6562,N_6282,N_6076);
nand U6563 (N_6563,N_6163,N_6033);
xor U6564 (N_6564,N_6191,N_6239);
nor U6565 (N_6565,N_6152,N_6058);
nand U6566 (N_6566,N_6067,N_6217);
nor U6567 (N_6567,N_6008,N_6033);
xor U6568 (N_6568,N_6058,N_6155);
or U6569 (N_6569,N_6164,N_6268);
or U6570 (N_6570,N_6180,N_6281);
nand U6571 (N_6571,N_6263,N_6039);
nor U6572 (N_6572,N_6284,N_6074);
or U6573 (N_6573,N_6288,N_6198);
or U6574 (N_6574,N_6023,N_6152);
and U6575 (N_6575,N_6266,N_6089);
or U6576 (N_6576,N_6132,N_6234);
nor U6577 (N_6577,N_6149,N_6106);
nor U6578 (N_6578,N_6150,N_6172);
nor U6579 (N_6579,N_6223,N_6217);
and U6580 (N_6580,N_6100,N_6063);
or U6581 (N_6581,N_6270,N_6035);
nand U6582 (N_6582,N_6072,N_6002);
nor U6583 (N_6583,N_6187,N_6234);
xor U6584 (N_6584,N_6012,N_6151);
or U6585 (N_6585,N_6007,N_6262);
and U6586 (N_6586,N_6225,N_6044);
and U6587 (N_6587,N_6082,N_6055);
nor U6588 (N_6588,N_6166,N_6101);
nor U6589 (N_6589,N_6296,N_6292);
or U6590 (N_6590,N_6259,N_6196);
and U6591 (N_6591,N_6236,N_6061);
nand U6592 (N_6592,N_6127,N_6234);
nand U6593 (N_6593,N_6021,N_6141);
xor U6594 (N_6594,N_6174,N_6100);
and U6595 (N_6595,N_6260,N_6047);
nand U6596 (N_6596,N_6035,N_6280);
or U6597 (N_6597,N_6187,N_6183);
and U6598 (N_6598,N_6103,N_6268);
nor U6599 (N_6599,N_6242,N_6150);
nor U6600 (N_6600,N_6413,N_6441);
xnor U6601 (N_6601,N_6443,N_6505);
nand U6602 (N_6602,N_6401,N_6481);
xor U6603 (N_6603,N_6367,N_6337);
or U6604 (N_6604,N_6327,N_6578);
xnor U6605 (N_6605,N_6406,N_6370);
nand U6606 (N_6606,N_6485,N_6597);
nand U6607 (N_6607,N_6586,N_6440);
or U6608 (N_6608,N_6416,N_6520);
xor U6609 (N_6609,N_6561,N_6487);
and U6610 (N_6610,N_6388,N_6421);
xnor U6611 (N_6611,N_6577,N_6400);
nand U6612 (N_6612,N_6403,N_6419);
xnor U6613 (N_6613,N_6471,N_6506);
nor U6614 (N_6614,N_6553,N_6596);
or U6615 (N_6615,N_6433,N_6306);
xor U6616 (N_6616,N_6531,N_6365);
and U6617 (N_6617,N_6303,N_6439);
nor U6618 (N_6618,N_6540,N_6530);
or U6619 (N_6619,N_6345,N_6323);
nand U6620 (N_6620,N_6305,N_6523);
nand U6621 (N_6621,N_6310,N_6491);
or U6622 (N_6622,N_6395,N_6591);
or U6623 (N_6623,N_6449,N_6516);
and U6624 (N_6624,N_6579,N_6386);
xor U6625 (N_6625,N_6428,N_6458);
nand U6626 (N_6626,N_6479,N_6363);
nor U6627 (N_6627,N_6353,N_6560);
xnor U6628 (N_6628,N_6372,N_6486);
or U6629 (N_6629,N_6338,N_6459);
nand U6630 (N_6630,N_6510,N_6430);
or U6631 (N_6631,N_6318,N_6456);
nor U6632 (N_6632,N_6326,N_6336);
nand U6633 (N_6633,N_6502,N_6394);
nor U6634 (N_6634,N_6349,N_6352);
nor U6635 (N_6635,N_6355,N_6442);
xor U6636 (N_6636,N_6474,N_6522);
xnor U6637 (N_6637,N_6521,N_6450);
and U6638 (N_6638,N_6311,N_6423);
and U6639 (N_6639,N_6564,N_6329);
and U6640 (N_6640,N_6472,N_6495);
nor U6641 (N_6641,N_6515,N_6374);
or U6642 (N_6642,N_6593,N_6420);
or U6643 (N_6643,N_6478,N_6599);
or U6644 (N_6644,N_6315,N_6504);
nand U6645 (N_6645,N_6470,N_6402);
and U6646 (N_6646,N_6542,N_6369);
nand U6647 (N_6647,N_6585,N_6565);
nor U6648 (N_6648,N_6525,N_6567);
xnor U6649 (N_6649,N_6431,N_6467);
and U6650 (N_6650,N_6508,N_6398);
nand U6651 (N_6651,N_6437,N_6387);
xnor U6652 (N_6652,N_6424,N_6497);
xor U6653 (N_6653,N_6528,N_6381);
nand U6654 (N_6654,N_6378,N_6408);
nand U6655 (N_6655,N_6538,N_6371);
and U6656 (N_6656,N_6598,N_6346);
nand U6657 (N_6657,N_6307,N_6526);
or U6658 (N_6658,N_6475,N_6463);
nor U6659 (N_6659,N_6314,N_6563);
nand U6660 (N_6660,N_6301,N_6536);
xnor U6661 (N_6661,N_6422,N_6569);
nand U6662 (N_6662,N_6350,N_6499);
nand U6663 (N_6663,N_6454,N_6583);
and U6664 (N_6664,N_6503,N_6366);
nor U6665 (N_6665,N_6317,N_6581);
xor U6666 (N_6666,N_6584,N_6405);
nand U6667 (N_6667,N_6488,N_6446);
nand U6668 (N_6668,N_6572,N_6376);
and U6669 (N_6669,N_6544,N_6348);
and U6670 (N_6670,N_6362,N_6529);
or U6671 (N_6671,N_6555,N_6432);
nand U6672 (N_6672,N_6385,N_6514);
or U6673 (N_6673,N_6466,N_6410);
nand U6674 (N_6674,N_6435,N_6556);
and U6675 (N_6675,N_6359,N_6332);
and U6676 (N_6676,N_6590,N_6429);
xor U6677 (N_6677,N_6546,N_6557);
nor U6678 (N_6678,N_6592,N_6302);
and U6679 (N_6679,N_6399,N_6507);
nand U6680 (N_6680,N_6483,N_6576);
xnor U6681 (N_6681,N_6460,N_6477);
xor U6682 (N_6682,N_6496,N_6316);
nand U6683 (N_6683,N_6451,N_6340);
nor U6684 (N_6684,N_6341,N_6574);
and U6685 (N_6685,N_6354,N_6453);
xnor U6686 (N_6686,N_6457,N_6547);
or U6687 (N_6687,N_6404,N_6489);
xor U6688 (N_6688,N_6589,N_6313);
nand U6689 (N_6689,N_6343,N_6462);
nand U6690 (N_6690,N_6415,N_6511);
nor U6691 (N_6691,N_6537,N_6490);
and U6692 (N_6692,N_6325,N_6300);
and U6693 (N_6693,N_6335,N_6309);
nor U6694 (N_6694,N_6364,N_6412);
and U6695 (N_6695,N_6445,N_6308);
nand U6696 (N_6696,N_6573,N_6319);
nor U6697 (N_6697,N_6494,N_6543);
nand U6698 (N_6698,N_6558,N_6562);
nor U6699 (N_6699,N_6551,N_6397);
nand U6700 (N_6700,N_6461,N_6541);
and U6701 (N_6701,N_6448,N_6358);
nor U6702 (N_6702,N_6407,N_6549);
and U6703 (N_6703,N_6357,N_6339);
and U6704 (N_6704,N_6333,N_6331);
and U6705 (N_6705,N_6492,N_6534);
nor U6706 (N_6706,N_6436,N_6351);
nand U6707 (N_6707,N_6361,N_6568);
nand U6708 (N_6708,N_6379,N_6392);
nor U6709 (N_6709,N_6512,N_6383);
nand U6710 (N_6710,N_6582,N_6390);
nand U6711 (N_6711,N_6334,N_6594);
xnor U6712 (N_6712,N_6513,N_6444);
nand U6713 (N_6713,N_6321,N_6587);
and U6714 (N_6714,N_6493,N_6535);
xnor U6715 (N_6715,N_6468,N_6476);
nand U6716 (N_6716,N_6465,N_6455);
nand U6717 (N_6717,N_6411,N_6548);
nor U6718 (N_6718,N_6391,N_6320);
or U6719 (N_6719,N_6377,N_6360);
nand U6720 (N_6720,N_6380,N_6588);
nor U6721 (N_6721,N_6595,N_6580);
xnor U6722 (N_6722,N_6356,N_6447);
and U6723 (N_6723,N_6519,N_6575);
nand U6724 (N_6724,N_6312,N_6552);
xor U6725 (N_6725,N_6389,N_6509);
nand U6726 (N_6726,N_6517,N_6524);
xnor U6727 (N_6727,N_6473,N_6469);
nor U6728 (N_6728,N_6342,N_6527);
nand U6729 (N_6729,N_6539,N_6368);
xnor U6730 (N_6730,N_6425,N_6427);
nand U6731 (N_6731,N_6452,N_6382);
and U6732 (N_6732,N_6393,N_6554);
nand U6733 (N_6733,N_6498,N_6396);
xnor U6734 (N_6734,N_6434,N_6417);
and U6735 (N_6735,N_6571,N_6500);
or U6736 (N_6736,N_6566,N_6373);
or U6737 (N_6737,N_6518,N_6559);
nand U6738 (N_6738,N_6418,N_6414);
xnor U6739 (N_6739,N_6482,N_6532);
or U6740 (N_6740,N_6545,N_6533);
xor U6741 (N_6741,N_6409,N_6501);
or U6742 (N_6742,N_6480,N_6328);
or U6743 (N_6743,N_6330,N_6550);
or U6744 (N_6744,N_6322,N_6375);
and U6745 (N_6745,N_6344,N_6484);
nand U6746 (N_6746,N_6324,N_6304);
nand U6747 (N_6747,N_6426,N_6384);
nor U6748 (N_6748,N_6570,N_6347);
nand U6749 (N_6749,N_6438,N_6464);
nor U6750 (N_6750,N_6482,N_6577);
nand U6751 (N_6751,N_6534,N_6538);
nand U6752 (N_6752,N_6335,N_6424);
or U6753 (N_6753,N_6468,N_6554);
xnor U6754 (N_6754,N_6586,N_6301);
nor U6755 (N_6755,N_6419,N_6439);
and U6756 (N_6756,N_6581,N_6334);
nand U6757 (N_6757,N_6476,N_6339);
or U6758 (N_6758,N_6505,N_6392);
xor U6759 (N_6759,N_6300,N_6399);
xor U6760 (N_6760,N_6331,N_6484);
nor U6761 (N_6761,N_6324,N_6339);
or U6762 (N_6762,N_6416,N_6577);
nor U6763 (N_6763,N_6329,N_6569);
nor U6764 (N_6764,N_6539,N_6352);
or U6765 (N_6765,N_6539,N_6487);
xnor U6766 (N_6766,N_6522,N_6545);
or U6767 (N_6767,N_6408,N_6572);
nand U6768 (N_6768,N_6347,N_6454);
and U6769 (N_6769,N_6553,N_6418);
nor U6770 (N_6770,N_6587,N_6444);
nor U6771 (N_6771,N_6367,N_6546);
or U6772 (N_6772,N_6426,N_6343);
nor U6773 (N_6773,N_6325,N_6317);
nand U6774 (N_6774,N_6341,N_6519);
and U6775 (N_6775,N_6597,N_6569);
and U6776 (N_6776,N_6550,N_6341);
or U6777 (N_6777,N_6524,N_6395);
nor U6778 (N_6778,N_6387,N_6445);
or U6779 (N_6779,N_6570,N_6505);
nand U6780 (N_6780,N_6431,N_6446);
xor U6781 (N_6781,N_6520,N_6516);
xor U6782 (N_6782,N_6390,N_6419);
nor U6783 (N_6783,N_6549,N_6452);
or U6784 (N_6784,N_6526,N_6486);
nand U6785 (N_6785,N_6346,N_6357);
or U6786 (N_6786,N_6329,N_6379);
xor U6787 (N_6787,N_6507,N_6369);
nor U6788 (N_6788,N_6474,N_6533);
nor U6789 (N_6789,N_6411,N_6540);
and U6790 (N_6790,N_6563,N_6474);
nor U6791 (N_6791,N_6558,N_6597);
and U6792 (N_6792,N_6484,N_6462);
and U6793 (N_6793,N_6366,N_6453);
or U6794 (N_6794,N_6573,N_6460);
and U6795 (N_6795,N_6421,N_6471);
or U6796 (N_6796,N_6364,N_6473);
xor U6797 (N_6797,N_6363,N_6588);
nand U6798 (N_6798,N_6555,N_6365);
nand U6799 (N_6799,N_6470,N_6537);
nand U6800 (N_6800,N_6573,N_6433);
xor U6801 (N_6801,N_6361,N_6370);
xnor U6802 (N_6802,N_6486,N_6301);
xor U6803 (N_6803,N_6359,N_6599);
xnor U6804 (N_6804,N_6472,N_6377);
nor U6805 (N_6805,N_6363,N_6496);
nand U6806 (N_6806,N_6347,N_6534);
or U6807 (N_6807,N_6518,N_6448);
and U6808 (N_6808,N_6505,N_6464);
xnor U6809 (N_6809,N_6553,N_6407);
or U6810 (N_6810,N_6465,N_6337);
or U6811 (N_6811,N_6310,N_6551);
nand U6812 (N_6812,N_6582,N_6371);
or U6813 (N_6813,N_6373,N_6583);
and U6814 (N_6814,N_6321,N_6470);
xor U6815 (N_6815,N_6353,N_6478);
nor U6816 (N_6816,N_6316,N_6336);
nor U6817 (N_6817,N_6446,N_6544);
and U6818 (N_6818,N_6495,N_6576);
xor U6819 (N_6819,N_6338,N_6396);
and U6820 (N_6820,N_6380,N_6566);
and U6821 (N_6821,N_6351,N_6379);
or U6822 (N_6822,N_6481,N_6550);
xor U6823 (N_6823,N_6408,N_6492);
and U6824 (N_6824,N_6436,N_6535);
xnor U6825 (N_6825,N_6508,N_6568);
nor U6826 (N_6826,N_6561,N_6456);
and U6827 (N_6827,N_6488,N_6375);
nor U6828 (N_6828,N_6307,N_6306);
or U6829 (N_6829,N_6487,N_6393);
nor U6830 (N_6830,N_6411,N_6415);
and U6831 (N_6831,N_6377,N_6537);
nor U6832 (N_6832,N_6337,N_6597);
or U6833 (N_6833,N_6429,N_6341);
or U6834 (N_6834,N_6448,N_6303);
and U6835 (N_6835,N_6344,N_6361);
xnor U6836 (N_6836,N_6534,N_6521);
nand U6837 (N_6837,N_6452,N_6319);
xnor U6838 (N_6838,N_6571,N_6341);
xor U6839 (N_6839,N_6355,N_6398);
xor U6840 (N_6840,N_6477,N_6360);
or U6841 (N_6841,N_6483,N_6402);
xor U6842 (N_6842,N_6316,N_6360);
and U6843 (N_6843,N_6584,N_6471);
nor U6844 (N_6844,N_6541,N_6438);
nor U6845 (N_6845,N_6499,N_6300);
or U6846 (N_6846,N_6521,N_6465);
xnor U6847 (N_6847,N_6453,N_6411);
nor U6848 (N_6848,N_6430,N_6572);
or U6849 (N_6849,N_6409,N_6450);
and U6850 (N_6850,N_6505,N_6499);
and U6851 (N_6851,N_6374,N_6314);
nor U6852 (N_6852,N_6444,N_6523);
nor U6853 (N_6853,N_6580,N_6562);
and U6854 (N_6854,N_6473,N_6423);
nor U6855 (N_6855,N_6572,N_6448);
nand U6856 (N_6856,N_6382,N_6537);
or U6857 (N_6857,N_6430,N_6483);
nand U6858 (N_6858,N_6381,N_6552);
or U6859 (N_6859,N_6421,N_6543);
and U6860 (N_6860,N_6572,N_6526);
and U6861 (N_6861,N_6488,N_6586);
and U6862 (N_6862,N_6554,N_6494);
xnor U6863 (N_6863,N_6330,N_6377);
xnor U6864 (N_6864,N_6565,N_6440);
nand U6865 (N_6865,N_6536,N_6363);
xnor U6866 (N_6866,N_6581,N_6432);
nand U6867 (N_6867,N_6371,N_6565);
nand U6868 (N_6868,N_6546,N_6405);
or U6869 (N_6869,N_6461,N_6416);
xor U6870 (N_6870,N_6314,N_6526);
nor U6871 (N_6871,N_6495,N_6551);
and U6872 (N_6872,N_6387,N_6335);
xnor U6873 (N_6873,N_6527,N_6515);
or U6874 (N_6874,N_6363,N_6452);
xnor U6875 (N_6875,N_6558,N_6301);
and U6876 (N_6876,N_6581,N_6375);
nand U6877 (N_6877,N_6459,N_6536);
xnor U6878 (N_6878,N_6594,N_6470);
or U6879 (N_6879,N_6395,N_6310);
or U6880 (N_6880,N_6460,N_6519);
xor U6881 (N_6881,N_6304,N_6386);
nand U6882 (N_6882,N_6454,N_6324);
xor U6883 (N_6883,N_6592,N_6575);
nor U6884 (N_6884,N_6395,N_6417);
and U6885 (N_6885,N_6585,N_6352);
and U6886 (N_6886,N_6572,N_6524);
and U6887 (N_6887,N_6381,N_6371);
nor U6888 (N_6888,N_6581,N_6356);
and U6889 (N_6889,N_6474,N_6531);
xor U6890 (N_6890,N_6519,N_6478);
nor U6891 (N_6891,N_6568,N_6523);
and U6892 (N_6892,N_6587,N_6409);
and U6893 (N_6893,N_6558,N_6376);
and U6894 (N_6894,N_6596,N_6410);
nor U6895 (N_6895,N_6467,N_6433);
nor U6896 (N_6896,N_6326,N_6352);
and U6897 (N_6897,N_6337,N_6529);
nand U6898 (N_6898,N_6384,N_6405);
or U6899 (N_6899,N_6564,N_6317);
nor U6900 (N_6900,N_6619,N_6804);
and U6901 (N_6901,N_6721,N_6730);
nor U6902 (N_6902,N_6883,N_6744);
and U6903 (N_6903,N_6766,N_6788);
xnor U6904 (N_6904,N_6647,N_6836);
xnor U6905 (N_6905,N_6839,N_6714);
nand U6906 (N_6906,N_6743,N_6603);
nand U6907 (N_6907,N_6728,N_6809);
nor U6908 (N_6908,N_6867,N_6848);
xor U6909 (N_6909,N_6843,N_6820);
and U6910 (N_6910,N_6754,N_6745);
or U6911 (N_6911,N_6801,N_6880);
nor U6912 (N_6912,N_6680,N_6733);
nand U6913 (N_6913,N_6897,N_6851);
and U6914 (N_6914,N_6856,N_6884);
nor U6915 (N_6915,N_6861,N_6854);
nand U6916 (N_6916,N_6660,N_6882);
or U6917 (N_6917,N_6677,N_6799);
or U6918 (N_6918,N_6739,N_6611);
xor U6919 (N_6919,N_6767,N_6890);
or U6920 (N_6920,N_6825,N_6702);
nand U6921 (N_6921,N_6841,N_6664);
or U6922 (N_6922,N_6698,N_6786);
or U6923 (N_6923,N_6625,N_6771);
nor U6924 (N_6924,N_6666,N_6668);
or U6925 (N_6925,N_6672,N_6830);
and U6926 (N_6926,N_6746,N_6876);
nand U6927 (N_6927,N_6859,N_6615);
nor U6928 (N_6928,N_6888,N_6895);
or U6929 (N_6929,N_6708,N_6777);
nor U6930 (N_6930,N_6738,N_6622);
nand U6931 (N_6931,N_6755,N_6640);
nand U6932 (N_6932,N_6759,N_6840);
nand U6933 (N_6933,N_6659,N_6782);
or U6934 (N_6934,N_6635,N_6600);
nor U6935 (N_6935,N_6661,N_6729);
or U6936 (N_6936,N_6627,N_6793);
nand U6937 (N_6937,N_6657,N_6797);
or U6938 (N_6938,N_6727,N_6826);
or U6939 (N_6939,N_6690,N_6697);
xnor U6940 (N_6940,N_6725,N_6893);
nor U6941 (N_6941,N_6869,N_6868);
or U6942 (N_6942,N_6631,N_6688);
nand U6943 (N_6943,N_6720,N_6683);
nand U6944 (N_6944,N_6696,N_6623);
and U6945 (N_6945,N_6773,N_6879);
xor U6946 (N_6946,N_6616,N_6673);
xor U6947 (N_6947,N_6858,N_6823);
nor U6948 (N_6948,N_6864,N_6860);
and U6949 (N_6949,N_6852,N_6734);
nand U6950 (N_6950,N_6781,N_6816);
or U6951 (N_6951,N_6682,N_6731);
and U6952 (N_6952,N_6662,N_6878);
nor U6953 (N_6953,N_6757,N_6792);
nor U6954 (N_6954,N_6607,N_6636);
nand U6955 (N_6955,N_6828,N_6686);
xor U6956 (N_6956,N_6772,N_6628);
and U6957 (N_6957,N_6778,N_6753);
or U6958 (N_6958,N_6703,N_6892);
xnor U6959 (N_6959,N_6694,N_6747);
nand U6960 (N_6960,N_6621,N_6751);
xnor U6961 (N_6961,N_6722,N_6775);
and U6962 (N_6962,N_6705,N_6761);
nor U6963 (N_6963,N_6613,N_6610);
and U6964 (N_6964,N_6704,N_6875);
nor U6965 (N_6965,N_6887,N_6667);
nand U6966 (N_6966,N_6764,N_6676);
nand U6967 (N_6967,N_6814,N_6762);
nor U6968 (N_6968,N_6630,N_6737);
nor U6969 (N_6969,N_6654,N_6700);
xor U6970 (N_6970,N_6871,N_6780);
nand U6971 (N_6971,N_6643,N_6711);
or U6972 (N_6972,N_6835,N_6629);
or U6973 (N_6973,N_6701,N_6857);
nor U6974 (N_6974,N_6715,N_6855);
and U6975 (N_6975,N_6606,N_6827);
or U6976 (N_6976,N_6609,N_6850);
and U6977 (N_6977,N_6834,N_6881);
or U6978 (N_6978,N_6644,N_6805);
and U6979 (N_6979,N_6832,N_6872);
and U6980 (N_6980,N_6874,N_6853);
xnor U6981 (N_6981,N_6679,N_6614);
nand U6982 (N_6982,N_6865,N_6655);
xor U6983 (N_6983,N_6763,N_6789);
nor U6984 (N_6984,N_6706,N_6646);
xnor U6985 (N_6985,N_6601,N_6674);
nor U6986 (N_6986,N_6724,N_6821);
and U6987 (N_6987,N_6695,N_6813);
and U6988 (N_6988,N_6692,N_6642);
xor U6989 (N_6989,N_6822,N_6651);
nand U6990 (N_6990,N_6794,N_6774);
or U6991 (N_6991,N_6784,N_6899);
nor U6992 (N_6992,N_6634,N_6829);
or U6993 (N_6993,N_6894,N_6663);
or U6994 (N_6994,N_6866,N_6817);
xnor U6995 (N_6995,N_6648,N_6624);
or U6996 (N_6996,N_6709,N_6633);
xor U6997 (N_6997,N_6833,N_6765);
xor U6998 (N_6998,N_6847,N_6741);
nand U6999 (N_6999,N_6842,N_6681);
nor U7000 (N_7000,N_6670,N_6810);
and U7001 (N_7001,N_6645,N_6618);
xor U7002 (N_7002,N_6653,N_6740);
nand U7003 (N_7003,N_6671,N_6849);
xor U7004 (N_7004,N_6718,N_6811);
or U7005 (N_7005,N_6838,N_6800);
and U7006 (N_7006,N_6803,N_6846);
and U7007 (N_7007,N_6873,N_6806);
xor U7008 (N_7008,N_6758,N_6769);
or U7009 (N_7009,N_6837,N_6815);
nand U7010 (N_7010,N_6626,N_6675);
nand U7011 (N_7011,N_6650,N_6768);
nand U7012 (N_7012,N_6604,N_6612);
nand U7013 (N_7013,N_6808,N_6641);
nand U7014 (N_7014,N_6691,N_6863);
and U7015 (N_7015,N_6844,N_6732);
or U7016 (N_7016,N_6742,N_6770);
nand U7017 (N_7017,N_6687,N_6713);
xnor U7018 (N_7018,N_6605,N_6812);
and U7019 (N_7019,N_6807,N_6752);
nand U7020 (N_7020,N_6710,N_6891);
xnor U7021 (N_7021,N_6886,N_6898);
xnor U7022 (N_7022,N_6776,N_6712);
and U7023 (N_7023,N_6723,N_6795);
nand U7024 (N_7024,N_6684,N_6783);
nor U7025 (N_7025,N_6870,N_6885);
nor U7026 (N_7026,N_6798,N_6699);
or U7027 (N_7027,N_6608,N_6750);
or U7028 (N_7028,N_6877,N_6735);
or U7029 (N_7029,N_6656,N_6748);
xnor U7030 (N_7030,N_6617,N_6749);
nor U7031 (N_7031,N_6796,N_6637);
and U7032 (N_7032,N_6818,N_6785);
nand U7033 (N_7033,N_6678,N_6620);
or U7034 (N_7034,N_6707,N_6889);
or U7035 (N_7035,N_6726,N_6756);
nor U7036 (N_7036,N_6652,N_6717);
nand U7037 (N_7037,N_6693,N_6791);
or U7038 (N_7038,N_6639,N_6649);
nand U7039 (N_7039,N_6669,N_6638);
nand U7040 (N_7040,N_6779,N_6719);
nor U7041 (N_7041,N_6716,N_6736);
nor U7042 (N_7042,N_6831,N_6685);
xnor U7043 (N_7043,N_6689,N_6602);
nand U7044 (N_7044,N_6862,N_6658);
xnor U7045 (N_7045,N_6824,N_6819);
xor U7046 (N_7046,N_6632,N_6896);
and U7047 (N_7047,N_6787,N_6802);
and U7048 (N_7048,N_6760,N_6790);
nor U7049 (N_7049,N_6665,N_6845);
and U7050 (N_7050,N_6884,N_6853);
xor U7051 (N_7051,N_6843,N_6609);
and U7052 (N_7052,N_6890,N_6781);
or U7053 (N_7053,N_6631,N_6866);
xnor U7054 (N_7054,N_6665,N_6869);
nand U7055 (N_7055,N_6725,N_6889);
and U7056 (N_7056,N_6769,N_6798);
or U7057 (N_7057,N_6631,N_6771);
nor U7058 (N_7058,N_6725,N_6758);
and U7059 (N_7059,N_6889,N_6667);
and U7060 (N_7060,N_6786,N_6799);
and U7061 (N_7061,N_6627,N_6722);
and U7062 (N_7062,N_6815,N_6777);
or U7063 (N_7063,N_6696,N_6809);
and U7064 (N_7064,N_6749,N_6695);
nand U7065 (N_7065,N_6774,N_6860);
or U7066 (N_7066,N_6605,N_6777);
nor U7067 (N_7067,N_6605,N_6708);
nand U7068 (N_7068,N_6626,N_6780);
xnor U7069 (N_7069,N_6704,N_6691);
nand U7070 (N_7070,N_6773,N_6887);
nand U7071 (N_7071,N_6829,N_6651);
or U7072 (N_7072,N_6715,N_6603);
and U7073 (N_7073,N_6668,N_6689);
nand U7074 (N_7074,N_6708,N_6624);
and U7075 (N_7075,N_6752,N_6675);
or U7076 (N_7076,N_6718,N_6705);
xor U7077 (N_7077,N_6866,N_6653);
xnor U7078 (N_7078,N_6851,N_6773);
nand U7079 (N_7079,N_6663,N_6858);
nor U7080 (N_7080,N_6770,N_6820);
xnor U7081 (N_7081,N_6703,N_6738);
nand U7082 (N_7082,N_6647,N_6656);
or U7083 (N_7083,N_6784,N_6839);
and U7084 (N_7084,N_6643,N_6878);
nor U7085 (N_7085,N_6661,N_6825);
or U7086 (N_7086,N_6741,N_6687);
and U7087 (N_7087,N_6808,N_6785);
nor U7088 (N_7088,N_6671,N_6889);
nor U7089 (N_7089,N_6704,N_6874);
nand U7090 (N_7090,N_6723,N_6792);
or U7091 (N_7091,N_6688,N_6642);
xnor U7092 (N_7092,N_6880,N_6657);
xor U7093 (N_7093,N_6796,N_6668);
or U7094 (N_7094,N_6608,N_6665);
nand U7095 (N_7095,N_6627,N_6678);
nor U7096 (N_7096,N_6627,N_6867);
and U7097 (N_7097,N_6882,N_6664);
and U7098 (N_7098,N_6787,N_6640);
nand U7099 (N_7099,N_6788,N_6792);
nand U7100 (N_7100,N_6690,N_6816);
xnor U7101 (N_7101,N_6626,N_6622);
or U7102 (N_7102,N_6716,N_6794);
nor U7103 (N_7103,N_6873,N_6613);
or U7104 (N_7104,N_6791,N_6722);
and U7105 (N_7105,N_6654,N_6616);
xnor U7106 (N_7106,N_6680,N_6725);
and U7107 (N_7107,N_6802,N_6724);
nor U7108 (N_7108,N_6672,N_6753);
or U7109 (N_7109,N_6881,N_6739);
nand U7110 (N_7110,N_6869,N_6745);
xnor U7111 (N_7111,N_6705,N_6782);
nand U7112 (N_7112,N_6746,N_6630);
nand U7113 (N_7113,N_6880,N_6797);
xor U7114 (N_7114,N_6709,N_6841);
or U7115 (N_7115,N_6643,N_6778);
xnor U7116 (N_7116,N_6646,N_6853);
nand U7117 (N_7117,N_6823,N_6678);
or U7118 (N_7118,N_6601,N_6715);
and U7119 (N_7119,N_6815,N_6751);
nand U7120 (N_7120,N_6705,N_6672);
nand U7121 (N_7121,N_6864,N_6710);
nand U7122 (N_7122,N_6891,N_6688);
xnor U7123 (N_7123,N_6661,N_6890);
and U7124 (N_7124,N_6647,N_6780);
xnor U7125 (N_7125,N_6601,N_6718);
nand U7126 (N_7126,N_6876,N_6741);
xor U7127 (N_7127,N_6629,N_6749);
or U7128 (N_7128,N_6680,N_6820);
and U7129 (N_7129,N_6776,N_6779);
nor U7130 (N_7130,N_6719,N_6646);
nand U7131 (N_7131,N_6605,N_6857);
or U7132 (N_7132,N_6785,N_6631);
xnor U7133 (N_7133,N_6725,N_6749);
xnor U7134 (N_7134,N_6709,N_6607);
nand U7135 (N_7135,N_6676,N_6888);
or U7136 (N_7136,N_6845,N_6848);
and U7137 (N_7137,N_6791,N_6665);
or U7138 (N_7138,N_6685,N_6602);
nand U7139 (N_7139,N_6760,N_6709);
or U7140 (N_7140,N_6763,N_6723);
and U7141 (N_7141,N_6722,N_6750);
nand U7142 (N_7142,N_6875,N_6766);
nor U7143 (N_7143,N_6867,N_6857);
nor U7144 (N_7144,N_6809,N_6725);
nor U7145 (N_7145,N_6828,N_6632);
or U7146 (N_7146,N_6777,N_6892);
nand U7147 (N_7147,N_6679,N_6746);
nand U7148 (N_7148,N_6878,N_6613);
nor U7149 (N_7149,N_6868,N_6670);
or U7150 (N_7150,N_6755,N_6622);
xnor U7151 (N_7151,N_6858,N_6632);
xor U7152 (N_7152,N_6881,N_6717);
or U7153 (N_7153,N_6724,N_6690);
or U7154 (N_7154,N_6848,N_6849);
nand U7155 (N_7155,N_6872,N_6715);
xor U7156 (N_7156,N_6859,N_6680);
nor U7157 (N_7157,N_6829,N_6773);
nor U7158 (N_7158,N_6836,N_6680);
and U7159 (N_7159,N_6810,N_6607);
nand U7160 (N_7160,N_6696,N_6674);
xor U7161 (N_7161,N_6686,N_6658);
and U7162 (N_7162,N_6799,N_6866);
and U7163 (N_7163,N_6869,N_6716);
nor U7164 (N_7164,N_6849,N_6687);
xnor U7165 (N_7165,N_6881,N_6829);
nor U7166 (N_7166,N_6897,N_6673);
nand U7167 (N_7167,N_6894,N_6604);
nand U7168 (N_7168,N_6871,N_6647);
or U7169 (N_7169,N_6786,N_6859);
xnor U7170 (N_7170,N_6685,N_6731);
nor U7171 (N_7171,N_6604,N_6606);
nand U7172 (N_7172,N_6823,N_6824);
or U7173 (N_7173,N_6622,N_6707);
or U7174 (N_7174,N_6696,N_6739);
or U7175 (N_7175,N_6815,N_6603);
or U7176 (N_7176,N_6877,N_6631);
and U7177 (N_7177,N_6675,N_6871);
nand U7178 (N_7178,N_6640,N_6811);
or U7179 (N_7179,N_6885,N_6809);
xor U7180 (N_7180,N_6704,N_6662);
and U7181 (N_7181,N_6777,N_6833);
nor U7182 (N_7182,N_6753,N_6777);
nor U7183 (N_7183,N_6856,N_6794);
xnor U7184 (N_7184,N_6875,N_6773);
xnor U7185 (N_7185,N_6725,N_6772);
nor U7186 (N_7186,N_6765,N_6614);
and U7187 (N_7187,N_6818,N_6843);
and U7188 (N_7188,N_6694,N_6868);
or U7189 (N_7189,N_6760,N_6762);
nor U7190 (N_7190,N_6898,N_6630);
xor U7191 (N_7191,N_6830,N_6613);
nor U7192 (N_7192,N_6749,N_6858);
xor U7193 (N_7193,N_6811,N_6741);
nor U7194 (N_7194,N_6782,N_6844);
nand U7195 (N_7195,N_6710,N_6740);
and U7196 (N_7196,N_6868,N_6831);
nor U7197 (N_7197,N_6855,N_6789);
or U7198 (N_7198,N_6605,N_6889);
or U7199 (N_7199,N_6679,N_6646);
nor U7200 (N_7200,N_7091,N_7123);
xnor U7201 (N_7201,N_7158,N_7116);
xnor U7202 (N_7202,N_7186,N_7055);
nor U7203 (N_7203,N_7028,N_7031);
nand U7204 (N_7204,N_7080,N_7019);
xnor U7205 (N_7205,N_6901,N_7046);
xor U7206 (N_7206,N_7069,N_6921);
and U7207 (N_7207,N_6920,N_7047);
xor U7208 (N_7208,N_6924,N_7197);
and U7209 (N_7209,N_7085,N_7119);
or U7210 (N_7210,N_7001,N_6900);
nand U7211 (N_7211,N_6982,N_7073);
nand U7212 (N_7212,N_7168,N_7065);
nor U7213 (N_7213,N_7102,N_7183);
nand U7214 (N_7214,N_7026,N_7188);
or U7215 (N_7215,N_7162,N_7193);
or U7216 (N_7216,N_7018,N_7045);
nand U7217 (N_7217,N_7023,N_7187);
or U7218 (N_7218,N_6918,N_7087);
nand U7219 (N_7219,N_7007,N_7052);
xor U7220 (N_7220,N_7191,N_6940);
or U7221 (N_7221,N_7160,N_7143);
and U7222 (N_7222,N_6917,N_7147);
xor U7223 (N_7223,N_7000,N_7051);
xor U7224 (N_7224,N_7092,N_6983);
and U7225 (N_7225,N_7159,N_6978);
nor U7226 (N_7226,N_7040,N_7189);
nand U7227 (N_7227,N_6987,N_7008);
nand U7228 (N_7228,N_6996,N_6999);
xnor U7229 (N_7229,N_7077,N_6991);
or U7230 (N_7230,N_7194,N_7120);
nand U7231 (N_7231,N_6923,N_6966);
and U7232 (N_7232,N_7009,N_7105);
xor U7233 (N_7233,N_7115,N_6937);
nand U7234 (N_7234,N_6947,N_6957);
xnor U7235 (N_7235,N_6922,N_7169);
nor U7236 (N_7236,N_7027,N_7070);
nor U7237 (N_7237,N_6960,N_7054);
or U7238 (N_7238,N_6968,N_6935);
nand U7239 (N_7239,N_7195,N_7131);
or U7240 (N_7240,N_6945,N_7185);
nor U7241 (N_7241,N_7100,N_6967);
xnor U7242 (N_7242,N_7012,N_7170);
or U7243 (N_7243,N_7049,N_7146);
nand U7244 (N_7244,N_7153,N_7083);
nor U7245 (N_7245,N_7056,N_7057);
nand U7246 (N_7246,N_6981,N_6906);
nand U7247 (N_7247,N_6969,N_7003);
nor U7248 (N_7248,N_6952,N_7048);
and U7249 (N_7249,N_7112,N_6926);
and U7250 (N_7250,N_6962,N_7122);
nand U7251 (N_7251,N_7064,N_7035);
nor U7252 (N_7252,N_7106,N_7068);
nor U7253 (N_7253,N_7075,N_6943);
nor U7254 (N_7254,N_7101,N_7103);
and U7255 (N_7255,N_6953,N_7182);
or U7256 (N_7256,N_6977,N_6914);
or U7257 (N_7257,N_6972,N_6958);
xnor U7258 (N_7258,N_7124,N_7174);
nor U7259 (N_7259,N_6976,N_7071);
and U7260 (N_7260,N_7020,N_7111);
nand U7261 (N_7261,N_7104,N_7139);
or U7262 (N_7262,N_7034,N_7044);
xor U7263 (N_7263,N_7021,N_7088);
nand U7264 (N_7264,N_7107,N_7173);
and U7265 (N_7265,N_7094,N_6990);
xor U7266 (N_7266,N_7011,N_7015);
nor U7267 (N_7267,N_7125,N_6995);
xnor U7268 (N_7268,N_7155,N_7133);
and U7269 (N_7269,N_6908,N_7099);
nand U7270 (N_7270,N_7144,N_6915);
nor U7271 (N_7271,N_6980,N_7072);
and U7272 (N_7272,N_7014,N_6949);
nand U7273 (N_7273,N_6964,N_7149);
and U7274 (N_7274,N_7117,N_7096);
nor U7275 (N_7275,N_6941,N_7150);
or U7276 (N_7276,N_7042,N_6904);
or U7277 (N_7277,N_6910,N_7050);
nor U7278 (N_7278,N_7062,N_7140);
or U7279 (N_7279,N_7178,N_7002);
or U7280 (N_7280,N_6913,N_6927);
nand U7281 (N_7281,N_6911,N_7137);
xor U7282 (N_7282,N_7037,N_7016);
or U7283 (N_7283,N_7126,N_7132);
or U7284 (N_7284,N_7164,N_7024);
xnor U7285 (N_7285,N_6942,N_7059);
nand U7286 (N_7286,N_7121,N_6989);
and U7287 (N_7287,N_7156,N_6932);
and U7288 (N_7288,N_6997,N_7175);
xor U7289 (N_7289,N_7081,N_7060);
nand U7290 (N_7290,N_7154,N_7098);
xnor U7291 (N_7291,N_6955,N_6903);
xor U7292 (N_7292,N_7029,N_6970);
nand U7293 (N_7293,N_6951,N_6938);
and U7294 (N_7294,N_7095,N_7030);
xor U7295 (N_7295,N_7127,N_7135);
and U7296 (N_7296,N_6973,N_6971);
nor U7297 (N_7297,N_6919,N_6946);
xnor U7298 (N_7298,N_6948,N_7198);
xor U7299 (N_7299,N_7084,N_7114);
and U7300 (N_7300,N_6905,N_7058);
or U7301 (N_7301,N_6930,N_6925);
xnor U7302 (N_7302,N_6907,N_6993);
xor U7303 (N_7303,N_7010,N_6975);
xnor U7304 (N_7304,N_7063,N_6954);
nand U7305 (N_7305,N_6988,N_7079);
or U7306 (N_7306,N_7134,N_7033);
xnor U7307 (N_7307,N_6950,N_7180);
xor U7308 (N_7308,N_7199,N_6928);
nor U7309 (N_7309,N_7192,N_7061);
nand U7310 (N_7310,N_7032,N_6992);
and U7311 (N_7311,N_7151,N_6933);
nand U7312 (N_7312,N_7097,N_7148);
and U7313 (N_7313,N_6998,N_6961);
nor U7314 (N_7314,N_7086,N_7141);
and U7315 (N_7315,N_6985,N_7053);
xor U7316 (N_7316,N_7025,N_7136);
nand U7317 (N_7317,N_7004,N_7179);
xnor U7318 (N_7318,N_7165,N_7129);
nand U7319 (N_7319,N_7036,N_7138);
or U7320 (N_7320,N_6944,N_7108);
xor U7321 (N_7321,N_7041,N_7017);
or U7322 (N_7322,N_7078,N_7172);
and U7323 (N_7323,N_7090,N_7118);
or U7324 (N_7324,N_7145,N_7157);
nor U7325 (N_7325,N_6916,N_7184);
nor U7326 (N_7326,N_7039,N_6934);
nor U7327 (N_7327,N_7166,N_6939);
xor U7328 (N_7328,N_7089,N_7043);
or U7329 (N_7329,N_7113,N_6974);
xnor U7330 (N_7330,N_7022,N_7093);
nor U7331 (N_7331,N_7130,N_6902);
or U7332 (N_7332,N_7177,N_7190);
and U7333 (N_7333,N_6984,N_6956);
xnor U7334 (N_7334,N_7152,N_7109);
and U7335 (N_7335,N_7013,N_7196);
or U7336 (N_7336,N_6994,N_7163);
xor U7337 (N_7337,N_6986,N_7176);
and U7338 (N_7338,N_6979,N_7074);
and U7339 (N_7339,N_7142,N_7167);
nor U7340 (N_7340,N_6931,N_7082);
or U7341 (N_7341,N_7128,N_6912);
and U7342 (N_7342,N_7181,N_7171);
and U7343 (N_7343,N_6929,N_6936);
or U7344 (N_7344,N_7005,N_6963);
nand U7345 (N_7345,N_7110,N_6959);
or U7346 (N_7346,N_7067,N_7066);
xor U7347 (N_7347,N_6909,N_7038);
or U7348 (N_7348,N_7076,N_6965);
nor U7349 (N_7349,N_7006,N_7161);
nor U7350 (N_7350,N_7177,N_7179);
xor U7351 (N_7351,N_7015,N_7142);
xnor U7352 (N_7352,N_6934,N_6901);
nor U7353 (N_7353,N_7138,N_6995);
xor U7354 (N_7354,N_6975,N_6911);
xnor U7355 (N_7355,N_6914,N_7106);
nor U7356 (N_7356,N_6999,N_6907);
nand U7357 (N_7357,N_7184,N_7006);
nand U7358 (N_7358,N_7115,N_7121);
or U7359 (N_7359,N_7107,N_6993);
or U7360 (N_7360,N_7029,N_7024);
nor U7361 (N_7361,N_7063,N_6911);
xor U7362 (N_7362,N_6953,N_6916);
and U7363 (N_7363,N_6937,N_6910);
or U7364 (N_7364,N_6986,N_7166);
and U7365 (N_7365,N_6958,N_7176);
nor U7366 (N_7366,N_7100,N_7162);
or U7367 (N_7367,N_7007,N_7092);
or U7368 (N_7368,N_6942,N_6965);
nand U7369 (N_7369,N_6912,N_7101);
or U7370 (N_7370,N_7075,N_6997);
or U7371 (N_7371,N_7071,N_7096);
and U7372 (N_7372,N_6952,N_7180);
nand U7373 (N_7373,N_7107,N_6915);
xnor U7374 (N_7374,N_7195,N_7055);
xor U7375 (N_7375,N_7070,N_7177);
nand U7376 (N_7376,N_7195,N_6924);
xnor U7377 (N_7377,N_7199,N_7065);
or U7378 (N_7378,N_6964,N_6942);
and U7379 (N_7379,N_7130,N_7045);
nor U7380 (N_7380,N_6944,N_7121);
nor U7381 (N_7381,N_7189,N_6912);
or U7382 (N_7382,N_7073,N_7004);
nand U7383 (N_7383,N_6965,N_7080);
nor U7384 (N_7384,N_7033,N_7077);
or U7385 (N_7385,N_7174,N_7181);
and U7386 (N_7386,N_6989,N_6937);
or U7387 (N_7387,N_6941,N_7003);
nand U7388 (N_7388,N_7152,N_6910);
nand U7389 (N_7389,N_7133,N_7071);
nor U7390 (N_7390,N_7080,N_7135);
or U7391 (N_7391,N_6949,N_6907);
xor U7392 (N_7392,N_7116,N_7182);
or U7393 (N_7393,N_6967,N_7058);
nand U7394 (N_7394,N_6905,N_7032);
or U7395 (N_7395,N_7135,N_6936);
nor U7396 (N_7396,N_7013,N_7112);
nor U7397 (N_7397,N_7100,N_6935);
xnor U7398 (N_7398,N_7146,N_6943);
nor U7399 (N_7399,N_6960,N_6970);
and U7400 (N_7400,N_7107,N_6914);
nor U7401 (N_7401,N_6925,N_7023);
and U7402 (N_7402,N_7070,N_7009);
nand U7403 (N_7403,N_7157,N_7013);
xnor U7404 (N_7404,N_7014,N_7020);
nor U7405 (N_7405,N_7106,N_7041);
nor U7406 (N_7406,N_7066,N_7178);
xor U7407 (N_7407,N_7132,N_7125);
and U7408 (N_7408,N_7149,N_7193);
xor U7409 (N_7409,N_7115,N_7004);
xor U7410 (N_7410,N_6935,N_6960);
or U7411 (N_7411,N_7080,N_6982);
nand U7412 (N_7412,N_6933,N_7086);
xnor U7413 (N_7413,N_7117,N_7019);
nand U7414 (N_7414,N_7190,N_7020);
and U7415 (N_7415,N_7101,N_6917);
or U7416 (N_7416,N_7066,N_6939);
nor U7417 (N_7417,N_7049,N_7097);
nor U7418 (N_7418,N_7081,N_7198);
and U7419 (N_7419,N_7133,N_6969);
or U7420 (N_7420,N_7085,N_7121);
nand U7421 (N_7421,N_6907,N_7173);
nor U7422 (N_7422,N_7021,N_7002);
or U7423 (N_7423,N_7099,N_6955);
nand U7424 (N_7424,N_6962,N_6949);
or U7425 (N_7425,N_7073,N_7161);
and U7426 (N_7426,N_7144,N_7111);
and U7427 (N_7427,N_7197,N_7025);
or U7428 (N_7428,N_7139,N_6932);
or U7429 (N_7429,N_6934,N_7153);
xor U7430 (N_7430,N_7051,N_7121);
nand U7431 (N_7431,N_7167,N_7160);
or U7432 (N_7432,N_7133,N_7134);
nor U7433 (N_7433,N_7133,N_7100);
xor U7434 (N_7434,N_7096,N_7034);
and U7435 (N_7435,N_7035,N_7042);
nor U7436 (N_7436,N_7151,N_6949);
nand U7437 (N_7437,N_7058,N_6920);
nand U7438 (N_7438,N_6984,N_7086);
or U7439 (N_7439,N_7159,N_6952);
or U7440 (N_7440,N_6945,N_7151);
nand U7441 (N_7441,N_7118,N_7091);
and U7442 (N_7442,N_7108,N_6941);
nand U7443 (N_7443,N_6963,N_6950);
or U7444 (N_7444,N_7043,N_7126);
and U7445 (N_7445,N_7194,N_7143);
or U7446 (N_7446,N_6915,N_7017);
xnor U7447 (N_7447,N_7104,N_6916);
xnor U7448 (N_7448,N_7192,N_6991);
and U7449 (N_7449,N_7148,N_7184);
xor U7450 (N_7450,N_7043,N_6937);
nand U7451 (N_7451,N_7015,N_6930);
and U7452 (N_7452,N_7032,N_7004);
xnor U7453 (N_7453,N_7137,N_7040);
nand U7454 (N_7454,N_7183,N_7016);
xor U7455 (N_7455,N_7018,N_6995);
and U7456 (N_7456,N_6931,N_6968);
nor U7457 (N_7457,N_7104,N_6998);
xor U7458 (N_7458,N_6923,N_6956);
nand U7459 (N_7459,N_6958,N_6998);
nand U7460 (N_7460,N_7036,N_7144);
or U7461 (N_7461,N_7142,N_6935);
or U7462 (N_7462,N_7165,N_7094);
or U7463 (N_7463,N_7155,N_7162);
and U7464 (N_7464,N_7077,N_7157);
nand U7465 (N_7465,N_7105,N_7149);
xor U7466 (N_7466,N_7042,N_7101);
nand U7467 (N_7467,N_7113,N_6965);
nand U7468 (N_7468,N_7180,N_7136);
and U7469 (N_7469,N_7167,N_6995);
and U7470 (N_7470,N_7154,N_7100);
or U7471 (N_7471,N_6996,N_7150);
nor U7472 (N_7472,N_7161,N_7139);
nor U7473 (N_7473,N_7092,N_6931);
nand U7474 (N_7474,N_6932,N_7072);
nand U7475 (N_7475,N_7005,N_7091);
or U7476 (N_7476,N_7089,N_7146);
or U7477 (N_7477,N_7187,N_6984);
nand U7478 (N_7478,N_7191,N_7081);
nand U7479 (N_7479,N_6982,N_7181);
xnor U7480 (N_7480,N_6963,N_6969);
xnor U7481 (N_7481,N_7021,N_6912);
and U7482 (N_7482,N_6935,N_7190);
and U7483 (N_7483,N_7107,N_6954);
or U7484 (N_7484,N_6941,N_6940);
and U7485 (N_7485,N_7106,N_7016);
or U7486 (N_7486,N_6925,N_7045);
and U7487 (N_7487,N_6945,N_6946);
nand U7488 (N_7488,N_7100,N_6919);
nand U7489 (N_7489,N_7071,N_7019);
xor U7490 (N_7490,N_6952,N_7158);
nor U7491 (N_7491,N_6959,N_7105);
nor U7492 (N_7492,N_7116,N_7110);
xor U7493 (N_7493,N_7092,N_7004);
nand U7494 (N_7494,N_6907,N_6996);
or U7495 (N_7495,N_6911,N_7040);
xor U7496 (N_7496,N_7181,N_6975);
xnor U7497 (N_7497,N_7043,N_7186);
or U7498 (N_7498,N_7149,N_6924);
or U7499 (N_7499,N_7113,N_6962);
or U7500 (N_7500,N_7379,N_7220);
xnor U7501 (N_7501,N_7229,N_7283);
or U7502 (N_7502,N_7307,N_7218);
nor U7503 (N_7503,N_7222,N_7387);
xnor U7504 (N_7504,N_7324,N_7395);
nand U7505 (N_7505,N_7391,N_7480);
or U7506 (N_7506,N_7421,N_7359);
nand U7507 (N_7507,N_7333,N_7228);
and U7508 (N_7508,N_7219,N_7373);
nand U7509 (N_7509,N_7315,N_7299);
or U7510 (N_7510,N_7204,N_7280);
and U7511 (N_7511,N_7331,N_7400);
or U7512 (N_7512,N_7304,N_7416);
xnor U7513 (N_7513,N_7383,N_7332);
and U7514 (N_7514,N_7362,N_7369);
nor U7515 (N_7515,N_7370,N_7368);
or U7516 (N_7516,N_7301,N_7216);
nor U7517 (N_7517,N_7436,N_7460);
xnor U7518 (N_7518,N_7429,N_7485);
and U7519 (N_7519,N_7310,N_7392);
or U7520 (N_7520,N_7442,N_7293);
and U7521 (N_7521,N_7457,N_7271);
or U7522 (N_7522,N_7206,N_7372);
and U7523 (N_7523,N_7358,N_7473);
xor U7524 (N_7524,N_7428,N_7462);
or U7525 (N_7525,N_7438,N_7406);
nand U7526 (N_7526,N_7207,N_7308);
and U7527 (N_7527,N_7361,N_7401);
and U7528 (N_7528,N_7217,N_7208);
and U7529 (N_7529,N_7330,N_7215);
and U7530 (N_7530,N_7491,N_7279);
xor U7531 (N_7531,N_7223,N_7212);
xnor U7532 (N_7532,N_7431,N_7479);
and U7533 (N_7533,N_7458,N_7487);
nand U7534 (N_7534,N_7482,N_7260);
and U7535 (N_7535,N_7341,N_7318);
or U7536 (N_7536,N_7264,N_7201);
nor U7537 (N_7537,N_7353,N_7478);
nor U7538 (N_7538,N_7337,N_7418);
xnor U7539 (N_7539,N_7495,N_7292);
or U7540 (N_7540,N_7481,N_7364);
and U7541 (N_7541,N_7242,N_7366);
xnor U7542 (N_7542,N_7407,N_7239);
nand U7543 (N_7543,N_7314,N_7261);
and U7544 (N_7544,N_7453,N_7465);
nand U7545 (N_7545,N_7302,N_7469);
nand U7546 (N_7546,N_7303,N_7329);
nand U7547 (N_7547,N_7237,N_7463);
nor U7548 (N_7548,N_7488,N_7384);
xnor U7549 (N_7549,N_7380,N_7371);
and U7550 (N_7550,N_7454,N_7266);
xor U7551 (N_7551,N_7238,N_7338);
and U7552 (N_7552,N_7270,N_7396);
nand U7553 (N_7553,N_7455,N_7496);
xor U7554 (N_7554,N_7464,N_7378);
nor U7555 (N_7555,N_7444,N_7357);
and U7556 (N_7556,N_7402,N_7425);
nor U7557 (N_7557,N_7413,N_7461);
xnor U7558 (N_7558,N_7347,N_7493);
nand U7559 (N_7559,N_7323,N_7398);
nor U7560 (N_7560,N_7348,N_7205);
and U7561 (N_7561,N_7472,N_7471);
xnor U7562 (N_7562,N_7352,N_7417);
and U7563 (N_7563,N_7450,N_7376);
or U7564 (N_7564,N_7268,N_7486);
xor U7565 (N_7565,N_7258,N_7351);
xor U7566 (N_7566,N_7349,N_7240);
nand U7567 (N_7567,N_7445,N_7403);
nor U7568 (N_7568,N_7397,N_7326);
and U7569 (N_7569,N_7499,N_7290);
or U7570 (N_7570,N_7382,N_7255);
and U7571 (N_7571,N_7325,N_7335);
xnor U7572 (N_7572,N_7286,N_7321);
and U7573 (N_7573,N_7483,N_7313);
nand U7574 (N_7574,N_7354,N_7251);
and U7575 (N_7575,N_7311,N_7297);
nor U7576 (N_7576,N_7451,N_7423);
or U7577 (N_7577,N_7257,N_7245);
xnor U7578 (N_7578,N_7278,N_7408);
xnor U7579 (N_7579,N_7411,N_7210);
or U7580 (N_7580,N_7225,N_7322);
and U7581 (N_7581,N_7389,N_7399);
and U7582 (N_7582,N_7433,N_7287);
or U7583 (N_7583,N_7443,N_7288);
nand U7584 (N_7584,N_7262,N_7284);
nor U7585 (N_7585,N_7494,N_7256);
or U7586 (N_7586,N_7340,N_7243);
or U7587 (N_7587,N_7441,N_7489);
nor U7588 (N_7588,N_7363,N_7319);
xnor U7589 (N_7589,N_7252,N_7226);
nand U7590 (N_7590,N_7422,N_7306);
xnor U7591 (N_7591,N_7381,N_7236);
or U7592 (N_7592,N_7447,N_7211);
and U7593 (N_7593,N_7439,N_7296);
xor U7594 (N_7594,N_7231,N_7275);
nand U7595 (N_7595,N_7435,N_7221);
or U7596 (N_7596,N_7437,N_7227);
or U7597 (N_7597,N_7232,N_7492);
or U7598 (N_7598,N_7336,N_7440);
or U7599 (N_7599,N_7388,N_7291);
xnor U7600 (N_7600,N_7356,N_7484);
xor U7601 (N_7601,N_7466,N_7498);
and U7602 (N_7602,N_7316,N_7214);
nor U7603 (N_7603,N_7320,N_7456);
or U7604 (N_7604,N_7432,N_7247);
nor U7605 (N_7605,N_7328,N_7298);
nand U7606 (N_7606,N_7360,N_7377);
or U7607 (N_7607,N_7374,N_7233);
and U7608 (N_7608,N_7241,N_7253);
nand U7609 (N_7609,N_7277,N_7434);
xor U7610 (N_7610,N_7295,N_7312);
xnor U7611 (N_7611,N_7339,N_7375);
xnor U7612 (N_7612,N_7209,N_7468);
nor U7613 (N_7613,N_7272,N_7459);
xor U7614 (N_7614,N_7249,N_7203);
xor U7615 (N_7615,N_7276,N_7365);
nand U7616 (N_7616,N_7274,N_7476);
and U7617 (N_7617,N_7367,N_7390);
and U7618 (N_7618,N_7317,N_7430);
and U7619 (N_7619,N_7265,N_7230);
nand U7620 (N_7620,N_7345,N_7234);
nand U7621 (N_7621,N_7254,N_7269);
nand U7622 (N_7622,N_7385,N_7474);
or U7623 (N_7623,N_7334,N_7224);
nand U7624 (N_7624,N_7410,N_7412);
nand U7625 (N_7625,N_7414,N_7281);
and U7626 (N_7626,N_7200,N_7490);
nand U7627 (N_7627,N_7246,N_7342);
or U7628 (N_7628,N_7446,N_7327);
nand U7629 (N_7629,N_7405,N_7250);
nor U7630 (N_7630,N_7244,N_7294);
nand U7631 (N_7631,N_7267,N_7420);
and U7632 (N_7632,N_7346,N_7475);
nand U7633 (N_7633,N_7394,N_7415);
nor U7634 (N_7634,N_7427,N_7477);
nor U7635 (N_7635,N_7470,N_7449);
nor U7636 (N_7636,N_7409,N_7213);
or U7637 (N_7637,N_7448,N_7386);
nor U7638 (N_7638,N_7273,N_7305);
nor U7639 (N_7639,N_7355,N_7202);
nor U7640 (N_7640,N_7263,N_7452);
nand U7641 (N_7641,N_7350,N_7497);
and U7642 (N_7642,N_7344,N_7285);
or U7643 (N_7643,N_7248,N_7235);
or U7644 (N_7644,N_7343,N_7259);
nand U7645 (N_7645,N_7426,N_7419);
xnor U7646 (N_7646,N_7467,N_7424);
and U7647 (N_7647,N_7309,N_7300);
or U7648 (N_7648,N_7289,N_7282);
xor U7649 (N_7649,N_7393,N_7404);
and U7650 (N_7650,N_7445,N_7254);
and U7651 (N_7651,N_7464,N_7451);
nor U7652 (N_7652,N_7205,N_7463);
xnor U7653 (N_7653,N_7234,N_7231);
xor U7654 (N_7654,N_7372,N_7238);
or U7655 (N_7655,N_7431,N_7202);
nand U7656 (N_7656,N_7396,N_7352);
and U7657 (N_7657,N_7238,N_7224);
xor U7658 (N_7658,N_7341,N_7389);
and U7659 (N_7659,N_7209,N_7226);
and U7660 (N_7660,N_7319,N_7314);
and U7661 (N_7661,N_7281,N_7280);
and U7662 (N_7662,N_7477,N_7266);
nand U7663 (N_7663,N_7356,N_7487);
nand U7664 (N_7664,N_7365,N_7454);
and U7665 (N_7665,N_7388,N_7419);
nand U7666 (N_7666,N_7304,N_7245);
nor U7667 (N_7667,N_7244,N_7360);
and U7668 (N_7668,N_7391,N_7251);
xor U7669 (N_7669,N_7221,N_7398);
or U7670 (N_7670,N_7237,N_7247);
and U7671 (N_7671,N_7313,N_7492);
nand U7672 (N_7672,N_7225,N_7313);
and U7673 (N_7673,N_7441,N_7492);
and U7674 (N_7674,N_7299,N_7417);
nor U7675 (N_7675,N_7369,N_7204);
xor U7676 (N_7676,N_7258,N_7246);
nor U7677 (N_7677,N_7364,N_7337);
nor U7678 (N_7678,N_7443,N_7266);
nor U7679 (N_7679,N_7378,N_7441);
and U7680 (N_7680,N_7282,N_7405);
and U7681 (N_7681,N_7406,N_7321);
or U7682 (N_7682,N_7377,N_7383);
nor U7683 (N_7683,N_7462,N_7226);
or U7684 (N_7684,N_7418,N_7217);
or U7685 (N_7685,N_7476,N_7246);
or U7686 (N_7686,N_7389,N_7285);
or U7687 (N_7687,N_7346,N_7228);
xnor U7688 (N_7688,N_7425,N_7343);
or U7689 (N_7689,N_7207,N_7401);
and U7690 (N_7690,N_7374,N_7225);
xor U7691 (N_7691,N_7265,N_7341);
and U7692 (N_7692,N_7455,N_7243);
xnor U7693 (N_7693,N_7267,N_7408);
xor U7694 (N_7694,N_7380,N_7278);
nand U7695 (N_7695,N_7425,N_7474);
and U7696 (N_7696,N_7248,N_7381);
nand U7697 (N_7697,N_7278,N_7443);
or U7698 (N_7698,N_7351,N_7284);
nand U7699 (N_7699,N_7318,N_7311);
or U7700 (N_7700,N_7338,N_7426);
and U7701 (N_7701,N_7384,N_7420);
and U7702 (N_7702,N_7335,N_7303);
and U7703 (N_7703,N_7382,N_7439);
and U7704 (N_7704,N_7266,N_7368);
and U7705 (N_7705,N_7337,N_7471);
nand U7706 (N_7706,N_7445,N_7304);
nand U7707 (N_7707,N_7257,N_7389);
nor U7708 (N_7708,N_7375,N_7482);
xnor U7709 (N_7709,N_7344,N_7392);
and U7710 (N_7710,N_7361,N_7278);
and U7711 (N_7711,N_7287,N_7302);
nor U7712 (N_7712,N_7410,N_7462);
nor U7713 (N_7713,N_7228,N_7390);
or U7714 (N_7714,N_7446,N_7328);
nor U7715 (N_7715,N_7324,N_7202);
nand U7716 (N_7716,N_7449,N_7307);
nand U7717 (N_7717,N_7470,N_7231);
or U7718 (N_7718,N_7471,N_7338);
xor U7719 (N_7719,N_7463,N_7448);
and U7720 (N_7720,N_7409,N_7446);
nor U7721 (N_7721,N_7202,N_7326);
xnor U7722 (N_7722,N_7430,N_7319);
and U7723 (N_7723,N_7426,N_7399);
nor U7724 (N_7724,N_7485,N_7227);
nor U7725 (N_7725,N_7297,N_7489);
or U7726 (N_7726,N_7293,N_7377);
nor U7727 (N_7727,N_7360,N_7415);
and U7728 (N_7728,N_7296,N_7416);
nor U7729 (N_7729,N_7479,N_7385);
nand U7730 (N_7730,N_7350,N_7336);
and U7731 (N_7731,N_7340,N_7222);
nand U7732 (N_7732,N_7444,N_7289);
nor U7733 (N_7733,N_7447,N_7247);
xor U7734 (N_7734,N_7477,N_7245);
xnor U7735 (N_7735,N_7313,N_7448);
or U7736 (N_7736,N_7222,N_7260);
xor U7737 (N_7737,N_7265,N_7379);
xnor U7738 (N_7738,N_7367,N_7478);
or U7739 (N_7739,N_7376,N_7216);
or U7740 (N_7740,N_7355,N_7366);
nand U7741 (N_7741,N_7449,N_7372);
and U7742 (N_7742,N_7341,N_7233);
or U7743 (N_7743,N_7415,N_7289);
or U7744 (N_7744,N_7415,N_7210);
nand U7745 (N_7745,N_7269,N_7289);
nor U7746 (N_7746,N_7455,N_7325);
nor U7747 (N_7747,N_7245,N_7223);
xor U7748 (N_7748,N_7489,N_7495);
or U7749 (N_7749,N_7498,N_7431);
or U7750 (N_7750,N_7270,N_7257);
xor U7751 (N_7751,N_7315,N_7293);
or U7752 (N_7752,N_7400,N_7433);
xor U7753 (N_7753,N_7342,N_7419);
xor U7754 (N_7754,N_7363,N_7453);
and U7755 (N_7755,N_7288,N_7352);
xor U7756 (N_7756,N_7475,N_7377);
nor U7757 (N_7757,N_7412,N_7320);
xor U7758 (N_7758,N_7393,N_7267);
nand U7759 (N_7759,N_7446,N_7232);
or U7760 (N_7760,N_7308,N_7282);
xor U7761 (N_7761,N_7220,N_7465);
or U7762 (N_7762,N_7312,N_7446);
nor U7763 (N_7763,N_7266,N_7330);
and U7764 (N_7764,N_7387,N_7224);
or U7765 (N_7765,N_7472,N_7268);
xor U7766 (N_7766,N_7217,N_7340);
and U7767 (N_7767,N_7277,N_7491);
xor U7768 (N_7768,N_7420,N_7321);
nand U7769 (N_7769,N_7244,N_7497);
nor U7770 (N_7770,N_7214,N_7226);
nor U7771 (N_7771,N_7404,N_7472);
and U7772 (N_7772,N_7479,N_7249);
and U7773 (N_7773,N_7305,N_7488);
nand U7774 (N_7774,N_7436,N_7331);
or U7775 (N_7775,N_7281,N_7264);
nor U7776 (N_7776,N_7293,N_7209);
and U7777 (N_7777,N_7431,N_7265);
nor U7778 (N_7778,N_7479,N_7330);
nor U7779 (N_7779,N_7456,N_7471);
or U7780 (N_7780,N_7305,N_7284);
or U7781 (N_7781,N_7310,N_7468);
xor U7782 (N_7782,N_7397,N_7462);
or U7783 (N_7783,N_7357,N_7323);
nand U7784 (N_7784,N_7347,N_7274);
or U7785 (N_7785,N_7413,N_7439);
and U7786 (N_7786,N_7350,N_7244);
and U7787 (N_7787,N_7289,N_7374);
and U7788 (N_7788,N_7392,N_7400);
or U7789 (N_7789,N_7255,N_7243);
and U7790 (N_7790,N_7316,N_7228);
nand U7791 (N_7791,N_7203,N_7450);
nand U7792 (N_7792,N_7327,N_7368);
nand U7793 (N_7793,N_7219,N_7374);
nand U7794 (N_7794,N_7396,N_7285);
and U7795 (N_7795,N_7339,N_7245);
and U7796 (N_7796,N_7493,N_7319);
xor U7797 (N_7797,N_7374,N_7243);
and U7798 (N_7798,N_7391,N_7255);
nor U7799 (N_7799,N_7377,N_7490);
xor U7800 (N_7800,N_7731,N_7780);
or U7801 (N_7801,N_7532,N_7736);
or U7802 (N_7802,N_7624,N_7641);
or U7803 (N_7803,N_7521,N_7786);
nor U7804 (N_7804,N_7748,N_7796);
or U7805 (N_7805,N_7631,N_7683);
nand U7806 (N_7806,N_7795,N_7746);
nor U7807 (N_7807,N_7600,N_7642);
nand U7808 (N_7808,N_7656,N_7615);
or U7809 (N_7809,N_7680,N_7516);
nand U7810 (N_7810,N_7534,N_7784);
xnor U7811 (N_7811,N_7639,N_7525);
and U7812 (N_7812,N_7640,N_7674);
or U7813 (N_7813,N_7609,N_7645);
or U7814 (N_7814,N_7566,N_7703);
nand U7815 (N_7815,N_7568,N_7774);
and U7816 (N_7816,N_7529,N_7794);
nand U7817 (N_7817,N_7638,N_7761);
xnor U7818 (N_7818,N_7760,N_7782);
nor U7819 (N_7819,N_7660,N_7507);
xor U7820 (N_7820,N_7653,N_7766);
nor U7821 (N_7821,N_7790,N_7730);
and U7822 (N_7822,N_7752,N_7553);
nand U7823 (N_7823,N_7739,N_7623);
nand U7824 (N_7824,N_7576,N_7517);
xor U7825 (N_7825,N_7626,N_7702);
xor U7826 (N_7826,N_7673,N_7539);
nand U7827 (N_7827,N_7548,N_7612);
nand U7828 (N_7828,N_7740,N_7617);
xor U7829 (N_7829,N_7754,N_7589);
xnor U7830 (N_7830,N_7599,N_7764);
xnor U7831 (N_7831,N_7561,N_7577);
nand U7832 (N_7832,N_7603,N_7585);
and U7833 (N_7833,N_7792,N_7592);
or U7834 (N_7834,N_7636,N_7565);
nand U7835 (N_7835,N_7671,N_7635);
and U7836 (N_7836,N_7533,N_7714);
or U7837 (N_7837,N_7750,N_7509);
and U7838 (N_7838,N_7727,N_7676);
xnor U7839 (N_7839,N_7717,N_7697);
nor U7840 (N_7840,N_7720,N_7707);
and U7841 (N_7841,N_7601,N_7513);
nand U7842 (N_7842,N_7772,N_7523);
nand U7843 (N_7843,N_7604,N_7527);
nor U7844 (N_7844,N_7745,N_7567);
or U7845 (N_7845,N_7569,N_7614);
or U7846 (N_7846,N_7651,N_7560);
nand U7847 (N_7847,N_7747,N_7751);
nand U7848 (N_7848,N_7749,N_7753);
nand U7849 (N_7849,N_7783,N_7520);
and U7850 (N_7850,N_7512,N_7771);
or U7851 (N_7851,N_7713,N_7552);
xnor U7852 (N_7852,N_7701,N_7789);
nor U7853 (N_7853,N_7555,N_7508);
and U7854 (N_7854,N_7578,N_7596);
nand U7855 (N_7855,N_7728,N_7598);
and U7856 (N_7856,N_7724,N_7506);
and U7857 (N_7857,N_7500,N_7594);
and U7858 (N_7858,N_7742,N_7545);
nor U7859 (N_7859,N_7510,N_7734);
xor U7860 (N_7860,N_7743,N_7778);
nand U7861 (N_7861,N_7770,N_7647);
or U7862 (N_7862,N_7538,N_7563);
xnor U7863 (N_7863,N_7712,N_7698);
and U7864 (N_7864,N_7665,N_7787);
or U7865 (N_7865,N_7652,N_7543);
nor U7866 (N_7866,N_7710,N_7721);
nor U7867 (N_7867,N_7515,N_7668);
nand U7868 (N_7868,N_7611,N_7556);
xor U7869 (N_7869,N_7708,N_7579);
and U7870 (N_7870,N_7776,N_7779);
xnor U7871 (N_7871,N_7646,N_7644);
xor U7872 (N_7872,N_7618,N_7629);
xor U7873 (N_7873,N_7670,N_7685);
or U7874 (N_7874,N_7602,N_7756);
and U7875 (N_7875,N_7726,N_7559);
xnor U7876 (N_7876,N_7706,N_7634);
nor U7877 (N_7877,N_7605,N_7524);
and U7878 (N_7878,N_7502,N_7661);
nand U7879 (N_7879,N_7658,N_7744);
nor U7880 (N_7880,N_7765,N_7622);
nor U7881 (N_7881,N_7590,N_7501);
and U7882 (N_7882,N_7530,N_7705);
xor U7883 (N_7883,N_7627,N_7704);
and U7884 (N_7884,N_7583,N_7700);
xor U7885 (N_7885,N_7672,N_7549);
nand U7886 (N_7886,N_7655,N_7630);
nor U7887 (N_7887,N_7554,N_7528);
nand U7888 (N_7888,N_7547,N_7608);
nor U7889 (N_7889,N_7562,N_7613);
nor U7890 (N_7890,N_7669,N_7620);
xor U7891 (N_7891,N_7628,N_7763);
or U7892 (N_7892,N_7711,N_7591);
and U7893 (N_7893,N_7649,N_7610);
and U7894 (N_7894,N_7518,N_7657);
nor U7895 (N_7895,N_7580,N_7632);
nor U7896 (N_7896,N_7755,N_7519);
and U7897 (N_7897,N_7675,N_7505);
or U7898 (N_7898,N_7769,N_7582);
xor U7899 (N_7899,N_7597,N_7682);
or U7900 (N_7900,N_7692,N_7575);
or U7901 (N_7901,N_7791,N_7619);
nor U7902 (N_7902,N_7664,N_7522);
nand U7903 (N_7903,N_7741,N_7551);
nand U7904 (N_7904,N_7695,N_7621);
xor U7905 (N_7905,N_7503,N_7722);
and U7906 (N_7906,N_7666,N_7526);
or U7907 (N_7907,N_7718,N_7775);
nand U7908 (N_7908,N_7633,N_7690);
nand U7909 (N_7909,N_7616,N_7587);
or U7910 (N_7910,N_7540,N_7537);
or U7911 (N_7911,N_7797,N_7696);
xor U7912 (N_7912,N_7662,N_7719);
xnor U7913 (N_7913,N_7684,N_7777);
and U7914 (N_7914,N_7699,N_7584);
nor U7915 (N_7915,N_7650,N_7678);
nor U7916 (N_7916,N_7758,N_7514);
and U7917 (N_7917,N_7781,N_7733);
xnor U7918 (N_7918,N_7738,N_7667);
and U7919 (N_7919,N_7564,N_7793);
nor U7920 (N_7920,N_7799,N_7536);
and U7921 (N_7921,N_7716,N_7574);
nor U7922 (N_7922,N_7725,N_7693);
nand U7923 (N_7923,N_7759,N_7773);
xor U7924 (N_7924,N_7542,N_7788);
or U7925 (N_7925,N_7798,N_7558);
nor U7926 (N_7926,N_7729,N_7606);
nand U7927 (N_7927,N_7643,N_7557);
or U7928 (N_7928,N_7694,N_7785);
xnor U7929 (N_7929,N_7637,N_7762);
nand U7930 (N_7930,N_7648,N_7723);
nand U7931 (N_7931,N_7570,N_7688);
or U7932 (N_7932,N_7546,N_7571);
or U7933 (N_7933,N_7541,N_7607);
nand U7934 (N_7934,N_7572,N_7691);
or U7935 (N_7935,N_7544,N_7625);
nor U7936 (N_7936,N_7595,N_7737);
nand U7937 (N_7937,N_7768,N_7686);
or U7938 (N_7938,N_7531,N_7593);
or U7939 (N_7939,N_7511,N_7687);
or U7940 (N_7940,N_7586,N_7504);
xnor U7941 (N_7941,N_7681,N_7654);
or U7942 (N_7942,N_7535,N_7679);
nor U7943 (N_7943,N_7715,N_7689);
and U7944 (N_7944,N_7735,N_7709);
nor U7945 (N_7945,N_7767,N_7581);
xor U7946 (N_7946,N_7663,N_7550);
nor U7947 (N_7947,N_7588,N_7677);
or U7948 (N_7948,N_7732,N_7757);
and U7949 (N_7949,N_7573,N_7659);
xor U7950 (N_7950,N_7508,N_7743);
nand U7951 (N_7951,N_7746,N_7715);
and U7952 (N_7952,N_7566,N_7609);
xor U7953 (N_7953,N_7675,N_7514);
xnor U7954 (N_7954,N_7587,N_7663);
or U7955 (N_7955,N_7725,N_7569);
xnor U7956 (N_7956,N_7523,N_7542);
nand U7957 (N_7957,N_7795,N_7557);
xor U7958 (N_7958,N_7575,N_7625);
nand U7959 (N_7959,N_7733,N_7667);
nor U7960 (N_7960,N_7690,N_7560);
and U7961 (N_7961,N_7794,N_7651);
nor U7962 (N_7962,N_7715,N_7560);
xor U7963 (N_7963,N_7579,N_7796);
xnor U7964 (N_7964,N_7549,N_7561);
and U7965 (N_7965,N_7752,N_7758);
xor U7966 (N_7966,N_7693,N_7504);
and U7967 (N_7967,N_7718,N_7621);
xor U7968 (N_7968,N_7660,N_7681);
xnor U7969 (N_7969,N_7686,N_7744);
nor U7970 (N_7970,N_7715,N_7513);
nor U7971 (N_7971,N_7780,N_7708);
and U7972 (N_7972,N_7630,N_7684);
nor U7973 (N_7973,N_7738,N_7637);
and U7974 (N_7974,N_7600,N_7503);
nand U7975 (N_7975,N_7565,N_7616);
or U7976 (N_7976,N_7551,N_7723);
xor U7977 (N_7977,N_7757,N_7711);
nor U7978 (N_7978,N_7583,N_7605);
nand U7979 (N_7979,N_7773,N_7686);
and U7980 (N_7980,N_7751,N_7701);
or U7981 (N_7981,N_7596,N_7609);
nand U7982 (N_7982,N_7593,N_7668);
nor U7983 (N_7983,N_7599,N_7534);
nor U7984 (N_7984,N_7550,N_7667);
xnor U7985 (N_7985,N_7641,N_7709);
nor U7986 (N_7986,N_7663,N_7626);
or U7987 (N_7987,N_7571,N_7530);
and U7988 (N_7988,N_7634,N_7713);
and U7989 (N_7989,N_7791,N_7580);
and U7990 (N_7990,N_7686,N_7543);
xnor U7991 (N_7991,N_7594,N_7702);
xnor U7992 (N_7992,N_7539,N_7544);
nand U7993 (N_7993,N_7777,N_7575);
and U7994 (N_7994,N_7633,N_7661);
nand U7995 (N_7995,N_7527,N_7519);
and U7996 (N_7996,N_7538,N_7638);
nand U7997 (N_7997,N_7722,N_7513);
nand U7998 (N_7998,N_7679,N_7556);
and U7999 (N_7999,N_7667,N_7637);
nand U8000 (N_8000,N_7794,N_7546);
nor U8001 (N_8001,N_7792,N_7634);
or U8002 (N_8002,N_7674,N_7799);
xor U8003 (N_8003,N_7763,N_7760);
and U8004 (N_8004,N_7550,N_7556);
or U8005 (N_8005,N_7776,N_7517);
and U8006 (N_8006,N_7573,N_7768);
nand U8007 (N_8007,N_7591,N_7564);
nor U8008 (N_8008,N_7789,N_7614);
nand U8009 (N_8009,N_7550,N_7623);
nor U8010 (N_8010,N_7633,N_7716);
nor U8011 (N_8011,N_7778,N_7716);
or U8012 (N_8012,N_7752,N_7780);
nor U8013 (N_8013,N_7663,N_7521);
nand U8014 (N_8014,N_7693,N_7751);
xnor U8015 (N_8015,N_7704,N_7589);
xnor U8016 (N_8016,N_7710,N_7660);
nand U8017 (N_8017,N_7662,N_7703);
and U8018 (N_8018,N_7780,N_7513);
nand U8019 (N_8019,N_7690,N_7650);
nand U8020 (N_8020,N_7687,N_7787);
nand U8021 (N_8021,N_7636,N_7631);
xnor U8022 (N_8022,N_7794,N_7704);
nor U8023 (N_8023,N_7673,N_7565);
nand U8024 (N_8024,N_7510,N_7659);
nor U8025 (N_8025,N_7765,N_7591);
or U8026 (N_8026,N_7777,N_7578);
or U8027 (N_8027,N_7683,N_7656);
and U8028 (N_8028,N_7769,N_7581);
xor U8029 (N_8029,N_7676,N_7677);
nand U8030 (N_8030,N_7580,N_7621);
nor U8031 (N_8031,N_7583,N_7746);
nand U8032 (N_8032,N_7576,N_7680);
or U8033 (N_8033,N_7614,N_7680);
nor U8034 (N_8034,N_7703,N_7785);
xor U8035 (N_8035,N_7589,N_7759);
nor U8036 (N_8036,N_7738,N_7662);
nor U8037 (N_8037,N_7580,N_7562);
nand U8038 (N_8038,N_7618,N_7738);
or U8039 (N_8039,N_7636,N_7564);
and U8040 (N_8040,N_7576,N_7627);
and U8041 (N_8041,N_7543,N_7704);
nor U8042 (N_8042,N_7572,N_7607);
or U8043 (N_8043,N_7687,N_7526);
xnor U8044 (N_8044,N_7770,N_7613);
and U8045 (N_8045,N_7530,N_7590);
nor U8046 (N_8046,N_7523,N_7649);
nand U8047 (N_8047,N_7540,N_7638);
nor U8048 (N_8048,N_7627,N_7602);
nor U8049 (N_8049,N_7765,N_7619);
nor U8050 (N_8050,N_7537,N_7789);
or U8051 (N_8051,N_7778,N_7714);
or U8052 (N_8052,N_7693,N_7625);
xnor U8053 (N_8053,N_7609,N_7501);
or U8054 (N_8054,N_7719,N_7773);
and U8055 (N_8055,N_7677,N_7567);
xnor U8056 (N_8056,N_7629,N_7510);
xor U8057 (N_8057,N_7799,N_7667);
xnor U8058 (N_8058,N_7524,N_7521);
nor U8059 (N_8059,N_7739,N_7597);
and U8060 (N_8060,N_7508,N_7553);
and U8061 (N_8061,N_7577,N_7670);
nand U8062 (N_8062,N_7582,N_7775);
nor U8063 (N_8063,N_7539,N_7533);
xor U8064 (N_8064,N_7737,N_7553);
and U8065 (N_8065,N_7614,N_7572);
nand U8066 (N_8066,N_7721,N_7716);
and U8067 (N_8067,N_7758,N_7600);
xor U8068 (N_8068,N_7797,N_7743);
or U8069 (N_8069,N_7542,N_7606);
nand U8070 (N_8070,N_7673,N_7786);
nand U8071 (N_8071,N_7755,N_7545);
nor U8072 (N_8072,N_7575,N_7717);
nand U8073 (N_8073,N_7671,N_7684);
or U8074 (N_8074,N_7572,N_7646);
or U8075 (N_8075,N_7531,N_7659);
nor U8076 (N_8076,N_7512,N_7558);
xnor U8077 (N_8077,N_7780,N_7798);
nor U8078 (N_8078,N_7659,N_7738);
nor U8079 (N_8079,N_7784,N_7724);
or U8080 (N_8080,N_7718,N_7594);
and U8081 (N_8081,N_7783,N_7669);
and U8082 (N_8082,N_7792,N_7503);
and U8083 (N_8083,N_7645,N_7757);
and U8084 (N_8084,N_7723,N_7707);
and U8085 (N_8085,N_7633,N_7590);
and U8086 (N_8086,N_7524,N_7660);
or U8087 (N_8087,N_7734,N_7747);
xor U8088 (N_8088,N_7624,N_7602);
nand U8089 (N_8089,N_7777,N_7620);
nand U8090 (N_8090,N_7618,N_7742);
and U8091 (N_8091,N_7656,N_7761);
nand U8092 (N_8092,N_7592,N_7649);
xor U8093 (N_8093,N_7767,N_7786);
and U8094 (N_8094,N_7768,N_7661);
and U8095 (N_8095,N_7587,N_7522);
and U8096 (N_8096,N_7784,N_7703);
and U8097 (N_8097,N_7702,N_7604);
nand U8098 (N_8098,N_7678,N_7511);
xnor U8099 (N_8099,N_7539,N_7604);
nand U8100 (N_8100,N_7953,N_8050);
nor U8101 (N_8101,N_7996,N_7803);
nand U8102 (N_8102,N_8041,N_7930);
nor U8103 (N_8103,N_7830,N_8048);
xor U8104 (N_8104,N_7977,N_7968);
nand U8105 (N_8105,N_7987,N_7989);
xor U8106 (N_8106,N_8082,N_7981);
xor U8107 (N_8107,N_7939,N_7837);
nand U8108 (N_8108,N_7894,N_8002);
nor U8109 (N_8109,N_8072,N_8015);
xnor U8110 (N_8110,N_8003,N_7958);
nor U8111 (N_8111,N_8047,N_8052);
nand U8112 (N_8112,N_7893,N_8009);
xor U8113 (N_8113,N_7844,N_7947);
and U8114 (N_8114,N_7880,N_7994);
xnor U8115 (N_8115,N_8049,N_8058);
nand U8116 (N_8116,N_8001,N_7806);
xnor U8117 (N_8117,N_7853,N_8054);
nand U8118 (N_8118,N_7805,N_7845);
nor U8119 (N_8119,N_7838,N_8020);
nor U8120 (N_8120,N_7962,N_7851);
nor U8121 (N_8121,N_7924,N_7869);
or U8122 (N_8122,N_7920,N_7857);
nand U8123 (N_8123,N_8027,N_7937);
xnor U8124 (N_8124,N_8066,N_7849);
nor U8125 (N_8125,N_7896,N_8080);
nor U8126 (N_8126,N_7943,N_7817);
and U8127 (N_8127,N_7909,N_7906);
or U8128 (N_8128,N_7951,N_7900);
xor U8129 (N_8129,N_7932,N_7864);
nor U8130 (N_8130,N_7917,N_7925);
nand U8131 (N_8131,N_8098,N_7928);
nor U8132 (N_8132,N_8095,N_7821);
nor U8133 (N_8133,N_7888,N_8033);
xor U8134 (N_8134,N_7948,N_8039);
and U8135 (N_8135,N_7867,N_7908);
and U8136 (N_8136,N_7833,N_8035);
nor U8137 (N_8137,N_7916,N_8069);
nor U8138 (N_8138,N_8060,N_8088);
nand U8139 (N_8139,N_7808,N_8030);
xnor U8140 (N_8140,N_7965,N_8016);
xnor U8141 (N_8141,N_8008,N_7855);
and U8142 (N_8142,N_7814,N_7938);
and U8143 (N_8143,N_8029,N_8018);
or U8144 (N_8144,N_8065,N_8005);
nor U8145 (N_8145,N_7865,N_7955);
nor U8146 (N_8146,N_8026,N_7990);
nand U8147 (N_8147,N_7941,N_7934);
nand U8148 (N_8148,N_7999,N_7966);
nand U8149 (N_8149,N_8099,N_8046);
nand U8150 (N_8150,N_8061,N_8021);
nand U8151 (N_8151,N_8006,N_7826);
or U8152 (N_8152,N_7991,N_7979);
and U8153 (N_8153,N_7829,N_7933);
nand U8154 (N_8154,N_7861,N_7970);
or U8155 (N_8155,N_7915,N_7828);
or U8156 (N_8156,N_7997,N_7822);
xor U8157 (N_8157,N_7863,N_7936);
nand U8158 (N_8158,N_8087,N_7842);
or U8159 (N_8159,N_7862,N_7903);
xor U8160 (N_8160,N_7910,N_7978);
or U8161 (N_8161,N_8056,N_7919);
xnor U8162 (N_8162,N_7887,N_8042);
nor U8163 (N_8163,N_8071,N_8079);
nand U8164 (N_8164,N_7813,N_7879);
xor U8165 (N_8165,N_7945,N_8004);
nand U8166 (N_8166,N_7975,N_8074);
and U8167 (N_8167,N_7804,N_7832);
nor U8168 (N_8168,N_8093,N_7971);
nand U8169 (N_8169,N_7839,N_8090);
nand U8170 (N_8170,N_7956,N_7843);
xor U8171 (N_8171,N_8025,N_7993);
nor U8172 (N_8172,N_7898,N_7995);
or U8173 (N_8173,N_8091,N_8059);
nand U8174 (N_8174,N_7847,N_7922);
or U8175 (N_8175,N_7964,N_7850);
nand U8176 (N_8176,N_7876,N_7834);
or U8177 (N_8177,N_8022,N_7960);
or U8178 (N_8178,N_8043,N_7949);
and U8179 (N_8179,N_7802,N_8064);
or U8180 (N_8180,N_7980,N_7877);
or U8181 (N_8181,N_7935,N_7882);
nand U8182 (N_8182,N_8014,N_7998);
nor U8183 (N_8183,N_8007,N_8032);
nand U8184 (N_8184,N_7889,N_7872);
xor U8185 (N_8185,N_8057,N_7890);
nand U8186 (N_8186,N_7874,N_8045);
or U8187 (N_8187,N_7897,N_7950);
nand U8188 (N_8188,N_8097,N_7818);
nand U8189 (N_8189,N_7883,N_7878);
nor U8190 (N_8190,N_8037,N_8051);
nor U8191 (N_8191,N_7940,N_7873);
xor U8192 (N_8192,N_8000,N_8034);
nor U8193 (N_8193,N_7901,N_7927);
and U8194 (N_8194,N_7866,N_7895);
xnor U8195 (N_8195,N_8086,N_7840);
nor U8196 (N_8196,N_7816,N_7807);
xnor U8197 (N_8197,N_7954,N_7820);
nor U8198 (N_8198,N_7836,N_7904);
nand U8199 (N_8199,N_7860,N_8068);
xor U8200 (N_8200,N_7913,N_7868);
nand U8201 (N_8201,N_7825,N_8094);
or U8202 (N_8202,N_7976,N_7858);
or U8203 (N_8203,N_8067,N_8044);
and U8204 (N_8204,N_7988,N_7815);
nand U8205 (N_8205,N_7944,N_7884);
or U8206 (N_8206,N_7923,N_7819);
nor U8207 (N_8207,N_7823,N_7946);
xnor U8208 (N_8208,N_7812,N_8092);
or U8209 (N_8209,N_7891,N_8055);
xnor U8210 (N_8210,N_7959,N_8031);
nand U8211 (N_8211,N_7871,N_7875);
or U8212 (N_8212,N_8019,N_7992);
nand U8213 (N_8213,N_7921,N_7899);
nand U8214 (N_8214,N_8023,N_8078);
nor U8215 (N_8215,N_8073,N_8028);
or U8216 (N_8216,N_7854,N_7926);
and U8217 (N_8217,N_8011,N_7810);
xnor U8218 (N_8218,N_7986,N_8038);
xnor U8219 (N_8219,N_8036,N_7800);
nor U8220 (N_8220,N_7982,N_8012);
xnor U8221 (N_8221,N_8053,N_7942);
xnor U8222 (N_8222,N_7952,N_7902);
or U8223 (N_8223,N_7912,N_7907);
xnor U8224 (N_8224,N_8085,N_8017);
or U8225 (N_8225,N_7881,N_8081);
nor U8226 (N_8226,N_7984,N_8083);
and U8227 (N_8227,N_7983,N_7831);
or U8228 (N_8228,N_7963,N_7973);
or U8229 (N_8229,N_7848,N_7985);
xor U8230 (N_8230,N_7852,N_7886);
xnor U8231 (N_8231,N_8013,N_7827);
nor U8232 (N_8232,N_7914,N_8075);
and U8233 (N_8233,N_7972,N_8010);
nor U8234 (N_8234,N_7856,N_8096);
nand U8235 (N_8235,N_7905,N_8070);
nor U8236 (N_8236,N_7957,N_8076);
nand U8237 (N_8237,N_7892,N_7974);
xnor U8238 (N_8238,N_7809,N_8062);
xor U8239 (N_8239,N_7911,N_7811);
and U8240 (N_8240,N_7846,N_8089);
nor U8241 (N_8241,N_8024,N_7929);
and U8242 (N_8242,N_7859,N_7969);
nor U8243 (N_8243,N_7824,N_8084);
xnor U8244 (N_8244,N_7870,N_8077);
xor U8245 (N_8245,N_8063,N_7801);
and U8246 (N_8246,N_8040,N_7931);
or U8247 (N_8247,N_7885,N_7841);
xnor U8248 (N_8248,N_7961,N_7835);
or U8249 (N_8249,N_7918,N_7967);
nand U8250 (N_8250,N_7885,N_7817);
nor U8251 (N_8251,N_8094,N_7896);
nand U8252 (N_8252,N_7802,N_7963);
or U8253 (N_8253,N_7996,N_7827);
or U8254 (N_8254,N_8052,N_7917);
nand U8255 (N_8255,N_8011,N_8072);
and U8256 (N_8256,N_7851,N_8076);
and U8257 (N_8257,N_8075,N_7834);
xor U8258 (N_8258,N_7904,N_7910);
and U8259 (N_8259,N_7813,N_7823);
nand U8260 (N_8260,N_7942,N_8009);
xnor U8261 (N_8261,N_7962,N_8038);
nor U8262 (N_8262,N_7825,N_7902);
nand U8263 (N_8263,N_8070,N_8078);
xnor U8264 (N_8264,N_8050,N_7969);
nor U8265 (N_8265,N_7953,N_8029);
nand U8266 (N_8266,N_7866,N_8005);
nand U8267 (N_8267,N_7963,N_8081);
nor U8268 (N_8268,N_7970,N_7807);
xnor U8269 (N_8269,N_7979,N_7916);
nand U8270 (N_8270,N_7810,N_7844);
nand U8271 (N_8271,N_8082,N_7944);
nor U8272 (N_8272,N_7947,N_7873);
nor U8273 (N_8273,N_8059,N_7882);
or U8274 (N_8274,N_7907,N_7877);
or U8275 (N_8275,N_8056,N_7971);
and U8276 (N_8276,N_7816,N_7919);
or U8277 (N_8277,N_7862,N_8064);
nand U8278 (N_8278,N_8023,N_7871);
and U8279 (N_8279,N_7946,N_8091);
nand U8280 (N_8280,N_7993,N_7833);
xor U8281 (N_8281,N_7871,N_7823);
xnor U8282 (N_8282,N_7970,N_7864);
nor U8283 (N_8283,N_8014,N_7940);
or U8284 (N_8284,N_8024,N_7858);
nand U8285 (N_8285,N_7827,N_7923);
nand U8286 (N_8286,N_7909,N_8048);
xnor U8287 (N_8287,N_7966,N_8022);
nor U8288 (N_8288,N_8056,N_8032);
nand U8289 (N_8289,N_8044,N_7910);
xor U8290 (N_8290,N_7865,N_7824);
or U8291 (N_8291,N_8079,N_7977);
nor U8292 (N_8292,N_8076,N_7893);
nand U8293 (N_8293,N_8080,N_7898);
nor U8294 (N_8294,N_7837,N_7817);
xnor U8295 (N_8295,N_8050,N_7826);
xnor U8296 (N_8296,N_7800,N_7806);
and U8297 (N_8297,N_7899,N_8029);
nor U8298 (N_8298,N_7819,N_7887);
or U8299 (N_8299,N_7907,N_8060);
nand U8300 (N_8300,N_7875,N_7967);
nor U8301 (N_8301,N_7926,N_7902);
xor U8302 (N_8302,N_7907,N_8053);
and U8303 (N_8303,N_8052,N_8071);
nand U8304 (N_8304,N_7950,N_7995);
xnor U8305 (N_8305,N_7880,N_7979);
xnor U8306 (N_8306,N_7988,N_7863);
nor U8307 (N_8307,N_8013,N_7815);
xnor U8308 (N_8308,N_7879,N_7867);
and U8309 (N_8309,N_8058,N_7978);
and U8310 (N_8310,N_7977,N_8089);
and U8311 (N_8311,N_8084,N_7877);
nor U8312 (N_8312,N_7897,N_7853);
nand U8313 (N_8313,N_8090,N_7880);
xor U8314 (N_8314,N_8064,N_7801);
and U8315 (N_8315,N_7835,N_7813);
xnor U8316 (N_8316,N_7840,N_7914);
and U8317 (N_8317,N_7889,N_8017);
nor U8318 (N_8318,N_7924,N_8011);
nor U8319 (N_8319,N_7948,N_7876);
nand U8320 (N_8320,N_7940,N_7911);
or U8321 (N_8321,N_7920,N_7800);
nand U8322 (N_8322,N_8003,N_7996);
xor U8323 (N_8323,N_7809,N_7909);
or U8324 (N_8324,N_8019,N_7842);
nand U8325 (N_8325,N_8019,N_7818);
or U8326 (N_8326,N_7978,N_8093);
or U8327 (N_8327,N_7834,N_8010);
and U8328 (N_8328,N_7920,N_7957);
and U8329 (N_8329,N_8029,N_7810);
or U8330 (N_8330,N_8081,N_8039);
and U8331 (N_8331,N_8061,N_7841);
and U8332 (N_8332,N_7847,N_8072);
or U8333 (N_8333,N_7837,N_7918);
nand U8334 (N_8334,N_8001,N_8071);
nand U8335 (N_8335,N_7901,N_7917);
xor U8336 (N_8336,N_7854,N_7865);
and U8337 (N_8337,N_8001,N_7825);
nand U8338 (N_8338,N_7866,N_8078);
nand U8339 (N_8339,N_8006,N_8009);
nand U8340 (N_8340,N_7984,N_7832);
nor U8341 (N_8341,N_7838,N_7852);
xor U8342 (N_8342,N_7821,N_7864);
nor U8343 (N_8343,N_8020,N_7893);
and U8344 (N_8344,N_7997,N_8055);
or U8345 (N_8345,N_8048,N_7907);
and U8346 (N_8346,N_8030,N_8003);
nor U8347 (N_8347,N_7824,N_8007);
or U8348 (N_8348,N_8090,N_8093);
xnor U8349 (N_8349,N_8027,N_7855);
xor U8350 (N_8350,N_7926,N_8096);
nand U8351 (N_8351,N_7947,N_7841);
or U8352 (N_8352,N_7990,N_8008);
nand U8353 (N_8353,N_8099,N_8028);
nand U8354 (N_8354,N_7969,N_8061);
and U8355 (N_8355,N_7992,N_7843);
and U8356 (N_8356,N_7993,N_7818);
or U8357 (N_8357,N_7846,N_7932);
and U8358 (N_8358,N_8045,N_7988);
xor U8359 (N_8359,N_7987,N_7812);
nand U8360 (N_8360,N_7987,N_7906);
or U8361 (N_8361,N_7868,N_7954);
or U8362 (N_8362,N_8041,N_8007);
or U8363 (N_8363,N_7825,N_8026);
xor U8364 (N_8364,N_7997,N_7949);
xnor U8365 (N_8365,N_8094,N_8018);
and U8366 (N_8366,N_8078,N_7901);
xnor U8367 (N_8367,N_8021,N_7803);
or U8368 (N_8368,N_7852,N_8017);
xor U8369 (N_8369,N_7929,N_7876);
and U8370 (N_8370,N_8069,N_7938);
xnor U8371 (N_8371,N_7891,N_7908);
nand U8372 (N_8372,N_7829,N_8063);
or U8373 (N_8373,N_8054,N_7865);
and U8374 (N_8374,N_7953,N_8013);
or U8375 (N_8375,N_7888,N_7825);
nand U8376 (N_8376,N_7849,N_7960);
nor U8377 (N_8377,N_8055,N_8030);
or U8378 (N_8378,N_8046,N_7809);
nand U8379 (N_8379,N_7839,N_7983);
xor U8380 (N_8380,N_8031,N_8046);
nand U8381 (N_8381,N_7809,N_8076);
and U8382 (N_8382,N_7917,N_7800);
xor U8383 (N_8383,N_7957,N_7807);
xor U8384 (N_8384,N_7935,N_7839);
and U8385 (N_8385,N_8022,N_7876);
xnor U8386 (N_8386,N_7964,N_7914);
nand U8387 (N_8387,N_7805,N_7909);
xor U8388 (N_8388,N_7806,N_7865);
nand U8389 (N_8389,N_8024,N_7863);
or U8390 (N_8390,N_7870,N_7940);
or U8391 (N_8391,N_7898,N_7845);
or U8392 (N_8392,N_8003,N_7908);
nor U8393 (N_8393,N_7946,N_8062);
nor U8394 (N_8394,N_8093,N_7949);
xor U8395 (N_8395,N_8022,N_7918);
and U8396 (N_8396,N_7864,N_7814);
xnor U8397 (N_8397,N_7977,N_7871);
nand U8398 (N_8398,N_7801,N_7849);
and U8399 (N_8399,N_7840,N_7920);
and U8400 (N_8400,N_8182,N_8240);
nand U8401 (N_8401,N_8104,N_8139);
xnor U8402 (N_8402,N_8229,N_8201);
and U8403 (N_8403,N_8347,N_8399);
nor U8404 (N_8404,N_8175,N_8381);
nand U8405 (N_8405,N_8141,N_8166);
nor U8406 (N_8406,N_8198,N_8327);
xor U8407 (N_8407,N_8164,N_8151);
nor U8408 (N_8408,N_8373,N_8336);
xor U8409 (N_8409,N_8316,N_8158);
and U8410 (N_8410,N_8185,N_8398);
nand U8411 (N_8411,N_8222,N_8226);
nor U8412 (N_8412,N_8156,N_8122);
nand U8413 (N_8413,N_8313,N_8136);
xnor U8414 (N_8414,N_8100,N_8211);
or U8415 (N_8415,N_8176,N_8333);
nand U8416 (N_8416,N_8110,N_8396);
xnor U8417 (N_8417,N_8249,N_8103);
and U8418 (N_8418,N_8271,N_8278);
nand U8419 (N_8419,N_8134,N_8173);
and U8420 (N_8420,N_8276,N_8304);
xor U8421 (N_8421,N_8135,N_8354);
nor U8422 (N_8422,N_8218,N_8317);
nor U8423 (N_8423,N_8338,N_8283);
and U8424 (N_8424,N_8309,N_8324);
xnor U8425 (N_8425,N_8294,N_8257);
nor U8426 (N_8426,N_8334,N_8183);
xor U8427 (N_8427,N_8128,N_8389);
nand U8428 (N_8428,N_8320,N_8132);
nand U8429 (N_8429,N_8267,N_8287);
nor U8430 (N_8430,N_8174,N_8146);
and U8431 (N_8431,N_8116,N_8125);
nand U8432 (N_8432,N_8179,N_8275);
xnor U8433 (N_8433,N_8351,N_8251);
nand U8434 (N_8434,N_8165,N_8379);
and U8435 (N_8435,N_8342,N_8353);
and U8436 (N_8436,N_8306,N_8344);
nand U8437 (N_8437,N_8207,N_8206);
or U8438 (N_8438,N_8299,N_8203);
and U8439 (N_8439,N_8140,N_8113);
nand U8440 (N_8440,N_8322,N_8177);
xnor U8441 (N_8441,N_8259,N_8239);
and U8442 (N_8442,N_8114,N_8314);
and U8443 (N_8443,N_8237,N_8231);
or U8444 (N_8444,N_8191,N_8170);
nand U8445 (N_8445,N_8199,N_8269);
nand U8446 (N_8446,N_8209,N_8377);
nand U8447 (N_8447,N_8321,N_8375);
nor U8448 (N_8448,N_8368,N_8210);
or U8449 (N_8449,N_8361,N_8169);
or U8450 (N_8450,N_8266,N_8325);
and U8451 (N_8451,N_8213,N_8350);
and U8452 (N_8452,N_8236,N_8129);
nand U8453 (N_8453,N_8323,N_8264);
and U8454 (N_8454,N_8247,N_8106);
or U8455 (N_8455,N_8118,N_8149);
nor U8456 (N_8456,N_8189,N_8292);
nor U8457 (N_8457,N_8367,N_8274);
xor U8458 (N_8458,N_8194,N_8296);
and U8459 (N_8459,N_8117,N_8348);
nor U8460 (N_8460,N_8248,N_8298);
xnor U8461 (N_8461,N_8310,N_8162);
or U8462 (N_8462,N_8131,N_8331);
nor U8463 (N_8463,N_8235,N_8355);
xor U8464 (N_8464,N_8150,N_8293);
or U8465 (N_8465,N_8246,N_8369);
nor U8466 (N_8466,N_8232,N_8153);
or U8467 (N_8467,N_8329,N_8378);
nor U8468 (N_8468,N_8187,N_8328);
xnor U8469 (N_8469,N_8288,N_8341);
xor U8470 (N_8470,N_8388,N_8291);
and U8471 (N_8471,N_8390,N_8301);
xor U8472 (N_8472,N_8282,N_8395);
nand U8473 (N_8473,N_8371,N_8343);
and U8474 (N_8474,N_8233,N_8385);
and U8475 (N_8475,N_8205,N_8124);
nand U8476 (N_8476,N_8238,N_8340);
nor U8477 (N_8477,N_8167,N_8252);
nand U8478 (N_8478,N_8305,N_8152);
and U8479 (N_8479,N_8302,N_8279);
xor U8480 (N_8480,N_8330,N_8258);
nand U8481 (N_8481,N_8145,N_8262);
xnor U8482 (N_8482,N_8184,N_8109);
nor U8483 (N_8483,N_8178,N_8391);
xnor U8484 (N_8484,N_8364,N_8360);
or U8485 (N_8485,N_8311,N_8332);
xor U8486 (N_8486,N_8380,N_8241);
or U8487 (N_8487,N_8171,N_8105);
nor U8488 (N_8488,N_8295,N_8228);
xnor U8489 (N_8489,N_8393,N_8190);
and U8490 (N_8490,N_8280,N_8133);
xnor U8491 (N_8491,N_8217,N_8244);
xnor U8492 (N_8492,N_8387,N_8215);
nand U8493 (N_8493,N_8358,N_8277);
xor U8494 (N_8494,N_8195,N_8337);
nand U8495 (N_8495,N_8245,N_8130);
nor U8496 (N_8496,N_8253,N_8144);
xnor U8497 (N_8497,N_8121,N_8386);
xnor U8498 (N_8498,N_8242,N_8202);
or U8499 (N_8499,N_8365,N_8359);
or U8500 (N_8500,N_8270,N_8273);
nor U8501 (N_8501,N_8374,N_8397);
nand U8502 (N_8502,N_8303,N_8286);
nand U8503 (N_8503,N_8260,N_8108);
or U8504 (N_8504,N_8221,N_8181);
nand U8505 (N_8505,N_8147,N_8155);
nor U8506 (N_8506,N_8256,N_8161);
or U8507 (N_8507,N_8339,N_8180);
and U8508 (N_8508,N_8297,N_8188);
or U8509 (N_8509,N_8312,N_8307);
and U8510 (N_8510,N_8230,N_8159);
or U8511 (N_8511,N_8261,N_8284);
or U8512 (N_8512,N_8308,N_8349);
nor U8513 (N_8513,N_8281,N_8326);
and U8514 (N_8514,N_8225,N_8392);
or U8515 (N_8515,N_8335,N_8372);
and U8516 (N_8516,N_8220,N_8120);
and U8517 (N_8517,N_8111,N_8160);
nand U8518 (N_8518,N_8148,N_8119);
nand U8519 (N_8519,N_8123,N_8234);
and U8520 (N_8520,N_8352,N_8383);
or U8521 (N_8521,N_8319,N_8289);
and U8522 (N_8522,N_8216,N_8197);
nand U8523 (N_8523,N_8127,N_8363);
or U8524 (N_8524,N_8346,N_8204);
nand U8525 (N_8525,N_8126,N_8186);
nor U8526 (N_8526,N_8272,N_8263);
nand U8527 (N_8527,N_8163,N_8243);
nor U8528 (N_8528,N_8172,N_8224);
or U8529 (N_8529,N_8102,N_8265);
and U8530 (N_8530,N_8315,N_8254);
nand U8531 (N_8531,N_8200,N_8219);
nand U8532 (N_8532,N_8223,N_8250);
nor U8533 (N_8533,N_8143,N_8138);
nand U8534 (N_8534,N_8366,N_8212);
xnor U8535 (N_8535,N_8300,N_8356);
nor U8536 (N_8536,N_8142,N_8196);
nor U8537 (N_8537,N_8384,N_8101);
nand U8538 (N_8538,N_8376,N_8137);
and U8539 (N_8539,N_8268,N_8362);
nor U8540 (N_8540,N_8227,N_8394);
nor U8541 (N_8541,N_8382,N_8192);
xor U8542 (N_8542,N_8193,N_8370);
nand U8543 (N_8543,N_8214,N_8357);
or U8544 (N_8544,N_8168,N_8112);
xor U8545 (N_8545,N_8318,N_8345);
nor U8546 (N_8546,N_8290,N_8285);
or U8547 (N_8547,N_8157,N_8107);
and U8548 (N_8548,N_8115,N_8255);
xnor U8549 (N_8549,N_8208,N_8154);
nand U8550 (N_8550,N_8196,N_8195);
nand U8551 (N_8551,N_8171,N_8330);
nor U8552 (N_8552,N_8237,N_8333);
xnor U8553 (N_8553,N_8322,N_8181);
nand U8554 (N_8554,N_8214,N_8355);
xnor U8555 (N_8555,N_8233,N_8210);
nand U8556 (N_8556,N_8396,N_8229);
nor U8557 (N_8557,N_8279,N_8249);
nor U8558 (N_8558,N_8196,N_8253);
nor U8559 (N_8559,N_8322,N_8151);
nor U8560 (N_8560,N_8251,N_8124);
nor U8561 (N_8561,N_8291,N_8354);
and U8562 (N_8562,N_8276,N_8328);
nand U8563 (N_8563,N_8102,N_8132);
nor U8564 (N_8564,N_8154,N_8204);
and U8565 (N_8565,N_8357,N_8379);
or U8566 (N_8566,N_8307,N_8126);
or U8567 (N_8567,N_8180,N_8323);
nand U8568 (N_8568,N_8112,N_8371);
or U8569 (N_8569,N_8202,N_8273);
nand U8570 (N_8570,N_8137,N_8112);
nor U8571 (N_8571,N_8170,N_8267);
nand U8572 (N_8572,N_8379,N_8323);
and U8573 (N_8573,N_8160,N_8276);
nand U8574 (N_8574,N_8214,N_8227);
nor U8575 (N_8575,N_8103,N_8148);
xnor U8576 (N_8576,N_8320,N_8250);
or U8577 (N_8577,N_8323,N_8355);
nand U8578 (N_8578,N_8209,N_8264);
xnor U8579 (N_8579,N_8104,N_8205);
xnor U8580 (N_8580,N_8111,N_8191);
or U8581 (N_8581,N_8342,N_8398);
nor U8582 (N_8582,N_8189,N_8117);
and U8583 (N_8583,N_8154,N_8306);
nand U8584 (N_8584,N_8293,N_8158);
nand U8585 (N_8585,N_8179,N_8305);
nand U8586 (N_8586,N_8317,N_8139);
xnor U8587 (N_8587,N_8372,N_8179);
nor U8588 (N_8588,N_8113,N_8365);
or U8589 (N_8589,N_8273,N_8224);
nor U8590 (N_8590,N_8312,N_8210);
nor U8591 (N_8591,N_8230,N_8375);
nor U8592 (N_8592,N_8285,N_8263);
nand U8593 (N_8593,N_8214,N_8157);
and U8594 (N_8594,N_8343,N_8129);
nor U8595 (N_8595,N_8211,N_8352);
nor U8596 (N_8596,N_8313,N_8269);
nand U8597 (N_8597,N_8144,N_8369);
or U8598 (N_8598,N_8189,N_8136);
nand U8599 (N_8599,N_8308,N_8264);
and U8600 (N_8600,N_8276,N_8124);
nand U8601 (N_8601,N_8321,N_8145);
or U8602 (N_8602,N_8128,N_8336);
or U8603 (N_8603,N_8138,N_8180);
and U8604 (N_8604,N_8120,N_8173);
nand U8605 (N_8605,N_8201,N_8282);
xnor U8606 (N_8606,N_8129,N_8356);
xnor U8607 (N_8607,N_8145,N_8125);
and U8608 (N_8608,N_8259,N_8185);
and U8609 (N_8609,N_8259,N_8157);
xnor U8610 (N_8610,N_8373,N_8249);
xnor U8611 (N_8611,N_8178,N_8145);
nor U8612 (N_8612,N_8380,N_8139);
and U8613 (N_8613,N_8273,N_8143);
nor U8614 (N_8614,N_8289,N_8306);
xnor U8615 (N_8615,N_8383,N_8348);
or U8616 (N_8616,N_8366,N_8355);
nand U8617 (N_8617,N_8208,N_8103);
xor U8618 (N_8618,N_8349,N_8385);
nor U8619 (N_8619,N_8101,N_8307);
nand U8620 (N_8620,N_8102,N_8313);
nor U8621 (N_8621,N_8385,N_8148);
xnor U8622 (N_8622,N_8226,N_8232);
xnor U8623 (N_8623,N_8388,N_8366);
nor U8624 (N_8624,N_8206,N_8176);
or U8625 (N_8625,N_8116,N_8342);
or U8626 (N_8626,N_8199,N_8289);
xnor U8627 (N_8627,N_8252,N_8107);
xor U8628 (N_8628,N_8300,N_8216);
xnor U8629 (N_8629,N_8270,N_8217);
and U8630 (N_8630,N_8258,N_8239);
nand U8631 (N_8631,N_8341,N_8376);
xnor U8632 (N_8632,N_8344,N_8192);
nand U8633 (N_8633,N_8153,N_8300);
xor U8634 (N_8634,N_8151,N_8326);
nand U8635 (N_8635,N_8293,N_8103);
xnor U8636 (N_8636,N_8308,N_8393);
nor U8637 (N_8637,N_8177,N_8338);
nor U8638 (N_8638,N_8229,N_8269);
xor U8639 (N_8639,N_8126,N_8393);
nand U8640 (N_8640,N_8375,N_8351);
and U8641 (N_8641,N_8317,N_8112);
nand U8642 (N_8642,N_8397,N_8217);
nand U8643 (N_8643,N_8256,N_8199);
and U8644 (N_8644,N_8306,N_8165);
and U8645 (N_8645,N_8385,N_8109);
nor U8646 (N_8646,N_8111,N_8177);
nand U8647 (N_8647,N_8356,N_8199);
xnor U8648 (N_8648,N_8190,N_8264);
or U8649 (N_8649,N_8298,N_8229);
xor U8650 (N_8650,N_8398,N_8204);
nor U8651 (N_8651,N_8333,N_8308);
nand U8652 (N_8652,N_8134,N_8379);
and U8653 (N_8653,N_8262,N_8396);
xor U8654 (N_8654,N_8127,N_8293);
and U8655 (N_8655,N_8177,N_8262);
nor U8656 (N_8656,N_8185,N_8116);
nor U8657 (N_8657,N_8117,N_8100);
xor U8658 (N_8658,N_8306,N_8221);
or U8659 (N_8659,N_8298,N_8155);
nand U8660 (N_8660,N_8150,N_8204);
nand U8661 (N_8661,N_8149,N_8209);
nor U8662 (N_8662,N_8315,N_8364);
and U8663 (N_8663,N_8170,N_8216);
nand U8664 (N_8664,N_8190,N_8363);
nand U8665 (N_8665,N_8372,N_8141);
nand U8666 (N_8666,N_8365,N_8166);
or U8667 (N_8667,N_8239,N_8218);
and U8668 (N_8668,N_8264,N_8351);
or U8669 (N_8669,N_8227,N_8186);
nand U8670 (N_8670,N_8369,N_8313);
xnor U8671 (N_8671,N_8262,N_8368);
and U8672 (N_8672,N_8364,N_8251);
or U8673 (N_8673,N_8255,N_8351);
nand U8674 (N_8674,N_8299,N_8160);
xor U8675 (N_8675,N_8180,N_8260);
nand U8676 (N_8676,N_8298,N_8381);
and U8677 (N_8677,N_8107,N_8267);
and U8678 (N_8678,N_8188,N_8364);
nand U8679 (N_8679,N_8180,N_8183);
xor U8680 (N_8680,N_8354,N_8257);
or U8681 (N_8681,N_8218,N_8265);
or U8682 (N_8682,N_8397,N_8285);
and U8683 (N_8683,N_8140,N_8149);
xnor U8684 (N_8684,N_8366,N_8210);
xor U8685 (N_8685,N_8124,N_8344);
or U8686 (N_8686,N_8257,N_8364);
or U8687 (N_8687,N_8200,N_8120);
nor U8688 (N_8688,N_8311,N_8165);
or U8689 (N_8689,N_8296,N_8243);
xnor U8690 (N_8690,N_8284,N_8263);
or U8691 (N_8691,N_8141,N_8158);
or U8692 (N_8692,N_8140,N_8371);
nor U8693 (N_8693,N_8201,N_8268);
nand U8694 (N_8694,N_8207,N_8174);
and U8695 (N_8695,N_8341,N_8269);
nand U8696 (N_8696,N_8203,N_8388);
and U8697 (N_8697,N_8331,N_8140);
or U8698 (N_8698,N_8265,N_8242);
xnor U8699 (N_8699,N_8335,N_8286);
nor U8700 (N_8700,N_8578,N_8444);
or U8701 (N_8701,N_8586,N_8605);
or U8702 (N_8702,N_8588,N_8447);
nand U8703 (N_8703,N_8419,N_8553);
and U8704 (N_8704,N_8493,N_8612);
and U8705 (N_8705,N_8417,N_8659);
or U8706 (N_8706,N_8457,N_8429);
and U8707 (N_8707,N_8585,N_8446);
nand U8708 (N_8708,N_8404,N_8531);
or U8709 (N_8709,N_8554,N_8480);
nand U8710 (N_8710,N_8563,N_8443);
or U8711 (N_8711,N_8547,N_8458);
nand U8712 (N_8712,N_8663,N_8473);
xnor U8713 (N_8713,N_8650,N_8652);
or U8714 (N_8714,N_8667,N_8522);
and U8715 (N_8715,N_8589,N_8475);
and U8716 (N_8716,N_8672,N_8519);
xnor U8717 (N_8717,N_8662,N_8539);
xnor U8718 (N_8718,N_8653,N_8540);
nand U8719 (N_8719,N_8565,N_8501);
nor U8720 (N_8720,N_8490,N_8476);
nor U8721 (N_8721,N_8409,N_8494);
nand U8722 (N_8722,N_8595,N_8421);
xnor U8723 (N_8723,N_8453,N_8546);
nand U8724 (N_8724,N_8425,N_8657);
nor U8725 (N_8725,N_8465,N_8602);
nand U8726 (N_8726,N_8575,N_8673);
xor U8727 (N_8727,N_8439,N_8509);
or U8728 (N_8728,N_8573,N_8402);
and U8729 (N_8729,N_8675,N_8526);
nor U8730 (N_8730,N_8536,N_8668);
and U8731 (N_8731,N_8503,N_8505);
nor U8732 (N_8732,N_8528,N_8572);
nand U8733 (N_8733,N_8568,N_8415);
nand U8734 (N_8734,N_8413,N_8628);
nor U8735 (N_8735,N_8431,N_8499);
nor U8736 (N_8736,N_8504,N_8643);
xnor U8737 (N_8737,N_8438,N_8464);
and U8738 (N_8738,N_8641,N_8613);
xor U8739 (N_8739,N_8689,N_8687);
xor U8740 (N_8740,N_8500,N_8508);
xnor U8741 (N_8741,N_8576,N_8681);
nand U8742 (N_8742,N_8460,N_8407);
nor U8743 (N_8743,N_8498,N_8455);
nor U8744 (N_8744,N_8511,N_8428);
nand U8745 (N_8745,N_8623,N_8635);
nand U8746 (N_8746,N_8424,N_8527);
nand U8747 (N_8747,N_8590,N_8558);
xor U8748 (N_8748,N_8485,N_8646);
nand U8749 (N_8749,N_8695,N_8597);
nor U8750 (N_8750,N_8412,N_8506);
or U8751 (N_8751,N_8640,N_8683);
xnor U8752 (N_8752,N_8607,N_8648);
or U8753 (N_8753,N_8682,N_8483);
and U8754 (N_8754,N_8693,N_8510);
nand U8755 (N_8755,N_8617,N_8456);
nor U8756 (N_8756,N_8618,N_8619);
and U8757 (N_8757,N_8434,N_8666);
or U8758 (N_8758,N_8684,N_8594);
xnor U8759 (N_8759,N_8474,N_8642);
nand U8760 (N_8760,N_8631,N_8552);
or U8761 (N_8761,N_8436,N_8468);
and U8762 (N_8762,N_8632,N_8598);
xor U8763 (N_8763,N_8604,N_8596);
and U8764 (N_8764,N_8537,N_8426);
nand U8765 (N_8765,N_8449,N_8654);
xor U8766 (N_8766,N_8678,N_8423);
xor U8767 (N_8767,N_8535,N_8410);
and U8768 (N_8768,N_8664,N_8452);
nand U8769 (N_8769,N_8420,N_8599);
nor U8770 (N_8770,N_8601,N_8451);
nand U8771 (N_8771,N_8430,N_8538);
nor U8772 (N_8772,N_8532,N_8471);
xor U8773 (N_8773,N_8524,N_8520);
nand U8774 (N_8774,N_8478,N_8679);
xor U8775 (N_8775,N_8685,N_8427);
nand U8776 (N_8776,N_8608,N_8658);
and U8777 (N_8777,N_8541,N_8516);
or U8778 (N_8778,N_8432,N_8656);
or U8779 (N_8779,N_8486,N_8669);
or U8780 (N_8780,N_8625,N_8561);
nand U8781 (N_8781,N_8611,N_8502);
and U8782 (N_8782,N_8651,N_8433);
or U8783 (N_8783,N_8661,N_8551);
xor U8784 (N_8784,N_8655,N_8512);
or U8785 (N_8785,N_8591,N_8448);
or U8786 (N_8786,N_8680,N_8636);
and U8787 (N_8787,N_8606,N_8569);
and U8788 (N_8788,N_8533,N_8530);
and U8789 (N_8789,N_8406,N_8521);
nor U8790 (N_8790,N_8699,N_8616);
nand U8791 (N_8791,N_8470,N_8484);
nand U8792 (N_8792,N_8624,N_8463);
nand U8793 (N_8793,N_8630,N_8697);
nand U8794 (N_8794,N_8534,N_8670);
nand U8795 (N_8795,N_8645,N_8497);
nand U8796 (N_8796,N_8644,N_8518);
xor U8797 (N_8797,N_8544,N_8462);
nand U8798 (N_8798,N_8639,N_8496);
xor U8799 (N_8799,N_8525,N_8593);
nor U8800 (N_8800,N_8564,N_8555);
and U8801 (N_8801,N_8517,N_8418);
nor U8802 (N_8802,N_8549,N_8400);
or U8803 (N_8803,N_8620,N_8514);
xnor U8804 (N_8804,N_8403,N_8691);
nor U8805 (N_8805,N_8548,N_8489);
nor U8806 (N_8806,N_8692,N_8582);
nand U8807 (N_8807,N_8515,N_8690);
nor U8808 (N_8808,N_8479,N_8556);
xnor U8809 (N_8809,N_8487,N_8686);
or U8810 (N_8810,N_8688,N_8583);
xnor U8811 (N_8811,N_8401,N_8492);
nor U8812 (N_8812,N_8621,N_8615);
nand U8813 (N_8813,N_8676,N_8580);
nor U8814 (N_8814,N_8482,N_8441);
and U8815 (N_8815,N_8408,N_8542);
and U8816 (N_8816,N_8507,N_8488);
and U8817 (N_8817,N_8629,N_8545);
xnor U8818 (N_8818,N_8466,N_8513);
and U8819 (N_8819,N_8647,N_8477);
and U8820 (N_8820,N_8469,N_8649);
and U8821 (N_8821,N_8622,N_8571);
xor U8822 (N_8822,N_8411,N_8435);
xor U8823 (N_8823,N_8461,N_8560);
xor U8824 (N_8824,N_8543,N_8638);
nand U8825 (N_8825,N_8592,N_8550);
and U8826 (N_8826,N_8416,N_8633);
nand U8827 (N_8827,N_8454,N_8696);
nor U8828 (N_8828,N_8467,N_8626);
and U8829 (N_8829,N_8529,N_8567);
nor U8830 (N_8830,N_8660,N_8495);
nor U8831 (N_8831,N_8442,N_8609);
or U8832 (N_8832,N_8637,N_8437);
and U8833 (N_8833,N_8694,N_8559);
nor U8834 (N_8834,N_8459,N_8677);
nand U8835 (N_8835,N_8566,N_8674);
xnor U8836 (N_8836,N_8445,N_8634);
and U8837 (N_8837,N_8665,N_8614);
nor U8838 (N_8838,N_8414,N_8577);
nand U8839 (N_8839,N_8491,N_8481);
xnor U8840 (N_8840,N_8627,N_8570);
xor U8841 (N_8841,N_8581,N_8584);
xor U8842 (N_8842,N_8698,N_8422);
and U8843 (N_8843,N_8671,N_8600);
nand U8844 (N_8844,N_8405,N_8587);
or U8845 (N_8845,N_8603,N_8579);
xor U8846 (N_8846,N_8610,N_8557);
xor U8847 (N_8847,N_8574,N_8523);
xor U8848 (N_8848,N_8472,N_8450);
and U8849 (N_8849,N_8440,N_8562);
nor U8850 (N_8850,N_8624,N_8608);
and U8851 (N_8851,N_8423,N_8651);
nand U8852 (N_8852,N_8520,N_8527);
xnor U8853 (N_8853,N_8445,N_8675);
or U8854 (N_8854,N_8646,N_8691);
xor U8855 (N_8855,N_8610,N_8571);
nor U8856 (N_8856,N_8601,N_8604);
xnor U8857 (N_8857,N_8556,N_8647);
nand U8858 (N_8858,N_8698,N_8666);
xor U8859 (N_8859,N_8518,N_8669);
xor U8860 (N_8860,N_8606,N_8432);
nor U8861 (N_8861,N_8607,N_8538);
nand U8862 (N_8862,N_8595,N_8523);
and U8863 (N_8863,N_8658,N_8458);
or U8864 (N_8864,N_8435,N_8582);
nor U8865 (N_8865,N_8448,N_8518);
nand U8866 (N_8866,N_8429,N_8453);
xor U8867 (N_8867,N_8680,N_8525);
and U8868 (N_8868,N_8611,N_8544);
xnor U8869 (N_8869,N_8465,N_8512);
and U8870 (N_8870,N_8536,N_8413);
nor U8871 (N_8871,N_8499,N_8547);
nand U8872 (N_8872,N_8621,N_8502);
and U8873 (N_8873,N_8681,N_8640);
and U8874 (N_8874,N_8527,N_8494);
or U8875 (N_8875,N_8458,N_8626);
nand U8876 (N_8876,N_8471,N_8450);
nor U8877 (N_8877,N_8681,N_8518);
and U8878 (N_8878,N_8555,N_8652);
xnor U8879 (N_8879,N_8480,N_8676);
nor U8880 (N_8880,N_8480,N_8429);
nor U8881 (N_8881,N_8498,N_8582);
nand U8882 (N_8882,N_8402,N_8430);
nor U8883 (N_8883,N_8522,N_8680);
nand U8884 (N_8884,N_8574,N_8404);
nand U8885 (N_8885,N_8549,N_8553);
and U8886 (N_8886,N_8402,N_8415);
and U8887 (N_8887,N_8483,N_8683);
and U8888 (N_8888,N_8486,N_8459);
xnor U8889 (N_8889,N_8651,N_8650);
nor U8890 (N_8890,N_8513,N_8417);
or U8891 (N_8891,N_8575,N_8478);
nor U8892 (N_8892,N_8553,N_8688);
xor U8893 (N_8893,N_8597,N_8415);
or U8894 (N_8894,N_8598,N_8684);
nand U8895 (N_8895,N_8490,N_8515);
and U8896 (N_8896,N_8680,N_8609);
and U8897 (N_8897,N_8409,N_8489);
nor U8898 (N_8898,N_8415,N_8652);
nand U8899 (N_8899,N_8647,N_8684);
xnor U8900 (N_8900,N_8663,N_8588);
nor U8901 (N_8901,N_8473,N_8566);
or U8902 (N_8902,N_8534,N_8466);
nand U8903 (N_8903,N_8673,N_8586);
nor U8904 (N_8904,N_8641,N_8605);
or U8905 (N_8905,N_8675,N_8513);
xnor U8906 (N_8906,N_8439,N_8628);
nand U8907 (N_8907,N_8617,N_8509);
and U8908 (N_8908,N_8550,N_8522);
nor U8909 (N_8909,N_8460,N_8572);
nor U8910 (N_8910,N_8584,N_8597);
or U8911 (N_8911,N_8693,N_8547);
nor U8912 (N_8912,N_8432,N_8697);
nor U8913 (N_8913,N_8451,N_8565);
xnor U8914 (N_8914,N_8689,N_8519);
xor U8915 (N_8915,N_8647,N_8683);
xnor U8916 (N_8916,N_8672,N_8667);
and U8917 (N_8917,N_8652,N_8470);
or U8918 (N_8918,N_8576,N_8491);
or U8919 (N_8919,N_8442,N_8682);
nor U8920 (N_8920,N_8491,N_8622);
xor U8921 (N_8921,N_8531,N_8485);
and U8922 (N_8922,N_8442,N_8562);
or U8923 (N_8923,N_8526,N_8694);
or U8924 (N_8924,N_8575,N_8696);
xor U8925 (N_8925,N_8593,N_8664);
and U8926 (N_8926,N_8603,N_8507);
xor U8927 (N_8927,N_8619,N_8610);
nand U8928 (N_8928,N_8629,N_8551);
and U8929 (N_8929,N_8602,N_8476);
xor U8930 (N_8930,N_8463,N_8565);
nor U8931 (N_8931,N_8586,N_8686);
nor U8932 (N_8932,N_8483,N_8402);
nor U8933 (N_8933,N_8513,N_8482);
and U8934 (N_8934,N_8666,N_8555);
and U8935 (N_8935,N_8629,N_8645);
nand U8936 (N_8936,N_8416,N_8442);
xor U8937 (N_8937,N_8442,N_8512);
nand U8938 (N_8938,N_8597,N_8605);
or U8939 (N_8939,N_8471,N_8625);
nand U8940 (N_8940,N_8424,N_8552);
or U8941 (N_8941,N_8457,N_8565);
and U8942 (N_8942,N_8467,N_8510);
and U8943 (N_8943,N_8525,N_8591);
and U8944 (N_8944,N_8644,N_8409);
xor U8945 (N_8945,N_8475,N_8480);
and U8946 (N_8946,N_8517,N_8446);
nand U8947 (N_8947,N_8454,N_8512);
or U8948 (N_8948,N_8584,N_8419);
xnor U8949 (N_8949,N_8561,N_8636);
nand U8950 (N_8950,N_8430,N_8582);
and U8951 (N_8951,N_8487,N_8479);
xor U8952 (N_8952,N_8656,N_8515);
or U8953 (N_8953,N_8611,N_8558);
and U8954 (N_8954,N_8428,N_8652);
xor U8955 (N_8955,N_8628,N_8554);
or U8956 (N_8956,N_8581,N_8537);
or U8957 (N_8957,N_8530,N_8619);
and U8958 (N_8958,N_8498,N_8444);
nor U8959 (N_8959,N_8614,N_8590);
and U8960 (N_8960,N_8500,N_8680);
or U8961 (N_8961,N_8495,N_8582);
or U8962 (N_8962,N_8479,N_8496);
or U8963 (N_8963,N_8496,N_8679);
and U8964 (N_8964,N_8688,N_8437);
xnor U8965 (N_8965,N_8572,N_8400);
xor U8966 (N_8966,N_8668,N_8530);
or U8967 (N_8967,N_8614,N_8493);
nor U8968 (N_8968,N_8506,N_8539);
xor U8969 (N_8969,N_8695,N_8490);
xor U8970 (N_8970,N_8416,N_8664);
nand U8971 (N_8971,N_8467,N_8578);
xor U8972 (N_8972,N_8680,N_8423);
xnor U8973 (N_8973,N_8573,N_8408);
xnor U8974 (N_8974,N_8679,N_8581);
and U8975 (N_8975,N_8532,N_8595);
and U8976 (N_8976,N_8535,N_8491);
or U8977 (N_8977,N_8553,N_8474);
xor U8978 (N_8978,N_8589,N_8506);
xor U8979 (N_8979,N_8487,N_8464);
and U8980 (N_8980,N_8557,N_8638);
and U8981 (N_8981,N_8496,N_8414);
nor U8982 (N_8982,N_8679,N_8563);
nand U8983 (N_8983,N_8440,N_8460);
xnor U8984 (N_8984,N_8693,N_8410);
and U8985 (N_8985,N_8607,N_8636);
xor U8986 (N_8986,N_8415,N_8620);
or U8987 (N_8987,N_8546,N_8640);
xnor U8988 (N_8988,N_8494,N_8515);
or U8989 (N_8989,N_8544,N_8675);
xor U8990 (N_8990,N_8617,N_8627);
and U8991 (N_8991,N_8527,N_8440);
or U8992 (N_8992,N_8565,N_8599);
xor U8993 (N_8993,N_8455,N_8474);
nor U8994 (N_8994,N_8582,N_8440);
or U8995 (N_8995,N_8480,N_8471);
or U8996 (N_8996,N_8405,N_8548);
or U8997 (N_8997,N_8655,N_8546);
nand U8998 (N_8998,N_8465,N_8483);
xnor U8999 (N_8999,N_8586,N_8652);
and U9000 (N_9000,N_8984,N_8710);
xnor U9001 (N_9001,N_8708,N_8960);
and U9002 (N_9002,N_8878,N_8797);
xnor U9003 (N_9003,N_8798,N_8873);
nand U9004 (N_9004,N_8906,N_8854);
nor U9005 (N_9005,N_8804,N_8808);
and U9006 (N_9006,N_8769,N_8875);
nor U9007 (N_9007,N_8755,N_8977);
xnor U9008 (N_9008,N_8774,N_8700);
xor U9009 (N_9009,N_8716,N_8794);
nand U9010 (N_9010,N_8968,N_8860);
and U9011 (N_9011,N_8999,N_8775);
xnor U9012 (N_9012,N_8861,N_8896);
xor U9013 (N_9013,N_8834,N_8949);
and U9014 (N_9014,N_8855,N_8891);
xnor U9015 (N_9015,N_8752,N_8868);
or U9016 (N_9016,N_8895,N_8777);
or U9017 (N_9017,N_8722,N_8840);
or U9018 (N_9018,N_8859,N_8835);
nor U9019 (N_9019,N_8836,N_8887);
nor U9020 (N_9020,N_8900,N_8731);
nand U9021 (N_9021,N_8729,N_8963);
nand U9022 (N_9022,N_8757,N_8701);
xnor U9023 (N_9023,N_8799,N_8718);
nand U9024 (N_9024,N_8947,N_8759);
xnor U9025 (N_9025,N_8918,N_8762);
and U9026 (N_9026,N_8974,N_8760);
xnor U9027 (N_9027,N_8998,N_8811);
nor U9028 (N_9028,N_8983,N_8733);
nand U9029 (N_9029,N_8886,N_8975);
nand U9030 (N_9030,N_8793,N_8819);
and U9031 (N_9031,N_8863,N_8969);
xnor U9032 (N_9032,N_8913,N_8862);
nor U9033 (N_9033,N_8806,N_8964);
and U9034 (N_9034,N_8931,N_8936);
or U9035 (N_9035,N_8736,N_8844);
nor U9036 (N_9036,N_8828,N_8935);
or U9037 (N_9037,N_8748,N_8781);
and U9038 (N_9038,N_8904,N_8989);
nor U9039 (N_9039,N_8986,N_8715);
nor U9040 (N_9040,N_8909,N_8917);
xor U9041 (N_9041,N_8948,N_8740);
xnor U9042 (N_9042,N_8761,N_8867);
nor U9043 (N_9043,N_8816,N_8962);
or U9044 (N_9044,N_8897,N_8877);
nand U9045 (N_9045,N_8884,N_8845);
nand U9046 (N_9046,N_8912,N_8823);
and U9047 (N_9047,N_8914,N_8952);
xor U9048 (N_9048,N_8915,N_8842);
or U9049 (N_9049,N_8837,N_8779);
nand U9050 (N_9050,N_8979,N_8832);
and U9051 (N_9051,N_8772,N_8782);
xnor U9052 (N_9052,N_8749,N_8869);
nor U9053 (N_9053,N_8871,N_8893);
nor U9054 (N_9054,N_8945,N_8780);
and U9055 (N_9055,N_8750,N_8714);
nand U9056 (N_9056,N_8805,N_8971);
or U9057 (N_9057,N_8751,N_8981);
xor U9058 (N_9058,N_8719,N_8851);
or U9059 (N_9059,N_8919,N_8928);
and U9060 (N_9060,N_8880,N_8728);
nor U9061 (N_9061,N_8902,N_8812);
or U9062 (N_9062,N_8784,N_8813);
nor U9063 (N_9063,N_8739,N_8747);
nor U9064 (N_9064,N_8857,N_8881);
or U9065 (N_9065,N_8786,N_8703);
nand U9066 (N_9066,N_8957,N_8792);
xnor U9067 (N_9067,N_8830,N_8734);
nand U9068 (N_9068,N_8717,N_8879);
xnor U9069 (N_9069,N_8820,N_8988);
or U9070 (N_9070,N_8892,N_8922);
nand U9071 (N_9071,N_8758,N_8985);
nor U9072 (N_9072,N_8724,N_8987);
and U9073 (N_9073,N_8911,N_8831);
xnor U9074 (N_9074,N_8940,N_8889);
and U9075 (N_9075,N_8991,N_8742);
xor U9076 (N_9076,N_8870,N_8932);
nor U9077 (N_9077,N_8982,N_8866);
nand U9078 (N_9078,N_8732,N_8796);
nand U9079 (N_9079,N_8905,N_8821);
xor U9080 (N_9080,N_8829,N_8921);
or U9081 (N_9081,N_8826,N_8966);
and U9082 (N_9082,N_8994,N_8803);
xor U9083 (N_9083,N_8920,N_8795);
or U9084 (N_9084,N_8705,N_8753);
nand U9085 (N_9085,N_8950,N_8980);
nor U9086 (N_9086,N_8815,N_8973);
or U9087 (N_9087,N_8771,N_8711);
and U9088 (N_9088,N_8888,N_8727);
nor U9089 (N_9089,N_8946,N_8843);
or U9090 (N_9090,N_8817,N_8925);
nand U9091 (N_9091,N_8965,N_8933);
xnor U9092 (N_9092,N_8953,N_8709);
xor U9093 (N_9093,N_8767,N_8783);
nor U9094 (N_9094,N_8814,N_8726);
xnor U9095 (N_9095,N_8995,N_8741);
and U9096 (N_9096,N_8926,N_8872);
and U9097 (N_9097,N_8941,N_8885);
and U9098 (N_9098,N_8942,N_8901);
xor U9099 (N_9099,N_8809,N_8944);
nand U9100 (N_9100,N_8930,N_8730);
or U9101 (N_9101,N_8756,N_8882);
or U9102 (N_9102,N_8744,N_8959);
or U9103 (N_9103,N_8849,N_8903);
xor U9104 (N_9104,N_8927,N_8838);
and U9105 (N_9105,N_8939,N_8800);
nand U9106 (N_9106,N_8787,N_8818);
nor U9107 (N_9107,N_8938,N_8990);
and U9108 (N_9108,N_8737,N_8883);
nand U9109 (N_9109,N_8707,N_8807);
or U9110 (N_9110,N_8763,N_8937);
nor U9111 (N_9111,N_8864,N_8721);
nand U9112 (N_9112,N_8955,N_8824);
nor U9113 (N_9113,N_8908,N_8746);
and U9114 (N_9114,N_8972,N_8778);
nand U9115 (N_9115,N_8773,N_8961);
nand U9116 (N_9116,N_8978,N_8704);
nand U9117 (N_9117,N_8791,N_8934);
or U9118 (N_9118,N_8993,N_8846);
and U9119 (N_9119,N_8833,N_8706);
nand U9120 (N_9120,N_8970,N_8720);
and U9121 (N_9121,N_8764,N_8850);
nor U9122 (N_9122,N_8874,N_8789);
xor U9123 (N_9123,N_8712,N_8743);
or U9124 (N_9124,N_8858,N_8992);
nand U9125 (N_9125,N_8827,N_8810);
nand U9126 (N_9126,N_8924,N_8856);
xnor U9127 (N_9127,N_8958,N_8725);
nor U9128 (N_9128,N_8956,N_8967);
and U9129 (N_9129,N_8996,N_8735);
xnor U9130 (N_9130,N_8745,N_8929);
xnor U9131 (N_9131,N_8876,N_8790);
nand U9132 (N_9132,N_8738,N_8802);
nand U9133 (N_9133,N_8976,N_8785);
and U9134 (N_9134,N_8768,N_8899);
or U9135 (N_9135,N_8898,N_8801);
nand U9136 (N_9136,N_8943,N_8702);
nor U9137 (N_9137,N_8825,N_8723);
xor U9138 (N_9138,N_8910,N_8765);
or U9139 (N_9139,N_8822,N_8890);
nor U9140 (N_9140,N_8954,N_8923);
nand U9141 (N_9141,N_8754,N_8841);
or U9142 (N_9142,N_8713,N_8894);
xor U9143 (N_9143,N_8997,N_8788);
nor U9144 (N_9144,N_8776,N_8766);
nor U9145 (N_9145,N_8951,N_8916);
and U9146 (N_9146,N_8852,N_8907);
nand U9147 (N_9147,N_8853,N_8839);
xnor U9148 (N_9148,N_8865,N_8848);
or U9149 (N_9149,N_8847,N_8770);
nor U9150 (N_9150,N_8844,N_8847);
nand U9151 (N_9151,N_8961,N_8800);
xnor U9152 (N_9152,N_8817,N_8971);
nor U9153 (N_9153,N_8833,N_8999);
nand U9154 (N_9154,N_8925,N_8705);
nor U9155 (N_9155,N_8750,N_8936);
nor U9156 (N_9156,N_8901,N_8965);
and U9157 (N_9157,N_8829,N_8874);
and U9158 (N_9158,N_8734,N_8869);
nor U9159 (N_9159,N_8707,N_8881);
xor U9160 (N_9160,N_8942,N_8808);
nor U9161 (N_9161,N_8949,N_8960);
nor U9162 (N_9162,N_8859,N_8737);
xor U9163 (N_9163,N_8919,N_8770);
or U9164 (N_9164,N_8953,N_8989);
nor U9165 (N_9165,N_8772,N_8920);
xnor U9166 (N_9166,N_8993,N_8952);
xor U9167 (N_9167,N_8954,N_8879);
and U9168 (N_9168,N_8953,N_8806);
or U9169 (N_9169,N_8866,N_8790);
nand U9170 (N_9170,N_8980,N_8901);
and U9171 (N_9171,N_8998,N_8988);
nand U9172 (N_9172,N_8851,N_8973);
nand U9173 (N_9173,N_8881,N_8896);
nor U9174 (N_9174,N_8784,N_8793);
and U9175 (N_9175,N_8727,N_8966);
or U9176 (N_9176,N_8845,N_8911);
and U9177 (N_9177,N_8817,N_8946);
or U9178 (N_9178,N_8871,N_8727);
or U9179 (N_9179,N_8909,N_8850);
and U9180 (N_9180,N_8877,N_8808);
nand U9181 (N_9181,N_8962,N_8717);
xor U9182 (N_9182,N_8766,N_8785);
and U9183 (N_9183,N_8889,N_8776);
and U9184 (N_9184,N_8900,N_8831);
nand U9185 (N_9185,N_8709,N_8910);
nand U9186 (N_9186,N_8890,N_8755);
nand U9187 (N_9187,N_8740,N_8848);
xor U9188 (N_9188,N_8707,N_8765);
nand U9189 (N_9189,N_8887,N_8777);
nor U9190 (N_9190,N_8733,N_8839);
nand U9191 (N_9191,N_8847,N_8972);
nor U9192 (N_9192,N_8998,N_8727);
and U9193 (N_9193,N_8802,N_8808);
or U9194 (N_9194,N_8853,N_8794);
and U9195 (N_9195,N_8960,N_8858);
and U9196 (N_9196,N_8945,N_8787);
and U9197 (N_9197,N_8861,N_8937);
nor U9198 (N_9198,N_8998,N_8957);
and U9199 (N_9199,N_8766,N_8770);
nand U9200 (N_9200,N_8725,N_8888);
nand U9201 (N_9201,N_8818,N_8947);
xnor U9202 (N_9202,N_8927,N_8775);
nand U9203 (N_9203,N_8886,N_8723);
nand U9204 (N_9204,N_8851,N_8780);
and U9205 (N_9205,N_8937,N_8752);
xor U9206 (N_9206,N_8821,N_8872);
nor U9207 (N_9207,N_8788,N_8897);
nand U9208 (N_9208,N_8950,N_8817);
nor U9209 (N_9209,N_8866,N_8878);
xor U9210 (N_9210,N_8791,N_8835);
xor U9211 (N_9211,N_8777,N_8719);
or U9212 (N_9212,N_8947,N_8762);
and U9213 (N_9213,N_8774,N_8980);
or U9214 (N_9214,N_8997,N_8736);
xnor U9215 (N_9215,N_8872,N_8733);
or U9216 (N_9216,N_8913,N_8909);
nand U9217 (N_9217,N_8926,N_8976);
xnor U9218 (N_9218,N_8951,N_8929);
and U9219 (N_9219,N_8718,N_8715);
nor U9220 (N_9220,N_8859,N_8862);
nand U9221 (N_9221,N_8787,N_8768);
nor U9222 (N_9222,N_8928,N_8811);
nand U9223 (N_9223,N_8781,N_8767);
and U9224 (N_9224,N_8965,N_8911);
nor U9225 (N_9225,N_8902,N_8772);
xnor U9226 (N_9226,N_8749,N_8852);
nor U9227 (N_9227,N_8812,N_8714);
nand U9228 (N_9228,N_8812,N_8762);
or U9229 (N_9229,N_8824,N_8820);
or U9230 (N_9230,N_8813,N_8799);
xnor U9231 (N_9231,N_8926,N_8830);
or U9232 (N_9232,N_8778,N_8978);
or U9233 (N_9233,N_8704,N_8713);
and U9234 (N_9234,N_8755,N_8907);
or U9235 (N_9235,N_8904,N_8930);
xnor U9236 (N_9236,N_8942,N_8946);
or U9237 (N_9237,N_8843,N_8706);
and U9238 (N_9238,N_8992,N_8850);
and U9239 (N_9239,N_8980,N_8721);
xor U9240 (N_9240,N_8850,N_8895);
xnor U9241 (N_9241,N_8702,N_8767);
and U9242 (N_9242,N_8775,N_8710);
and U9243 (N_9243,N_8887,N_8757);
and U9244 (N_9244,N_8875,N_8829);
xor U9245 (N_9245,N_8931,N_8730);
nand U9246 (N_9246,N_8923,N_8971);
xnor U9247 (N_9247,N_8909,N_8883);
nand U9248 (N_9248,N_8916,N_8884);
or U9249 (N_9249,N_8924,N_8776);
and U9250 (N_9250,N_8988,N_8962);
xnor U9251 (N_9251,N_8853,N_8968);
or U9252 (N_9252,N_8943,N_8970);
or U9253 (N_9253,N_8920,N_8710);
xor U9254 (N_9254,N_8745,N_8967);
or U9255 (N_9255,N_8841,N_8808);
nor U9256 (N_9256,N_8897,N_8988);
xor U9257 (N_9257,N_8846,N_8711);
nand U9258 (N_9258,N_8968,N_8731);
or U9259 (N_9259,N_8719,N_8756);
or U9260 (N_9260,N_8757,N_8768);
nor U9261 (N_9261,N_8915,N_8968);
or U9262 (N_9262,N_8919,N_8912);
nor U9263 (N_9263,N_8900,N_8775);
or U9264 (N_9264,N_8810,N_8855);
nand U9265 (N_9265,N_8837,N_8944);
and U9266 (N_9266,N_8847,N_8719);
or U9267 (N_9267,N_8944,N_8991);
nor U9268 (N_9268,N_8962,N_8863);
nand U9269 (N_9269,N_8840,N_8935);
nor U9270 (N_9270,N_8797,N_8958);
or U9271 (N_9271,N_8978,N_8837);
or U9272 (N_9272,N_8850,N_8812);
nor U9273 (N_9273,N_8755,N_8759);
nand U9274 (N_9274,N_8870,N_8854);
and U9275 (N_9275,N_8928,N_8776);
xor U9276 (N_9276,N_8772,N_8794);
xor U9277 (N_9277,N_8715,N_8950);
and U9278 (N_9278,N_8975,N_8720);
or U9279 (N_9279,N_8927,N_8792);
nand U9280 (N_9280,N_8949,N_8785);
and U9281 (N_9281,N_8866,N_8976);
nand U9282 (N_9282,N_8713,N_8969);
xor U9283 (N_9283,N_8805,N_8795);
xor U9284 (N_9284,N_8924,N_8707);
or U9285 (N_9285,N_8789,N_8856);
nor U9286 (N_9286,N_8865,N_8845);
nor U9287 (N_9287,N_8985,N_8872);
and U9288 (N_9288,N_8871,N_8943);
nand U9289 (N_9289,N_8821,N_8981);
or U9290 (N_9290,N_8716,N_8770);
and U9291 (N_9291,N_8911,N_8897);
or U9292 (N_9292,N_8838,N_8845);
and U9293 (N_9293,N_8848,N_8976);
or U9294 (N_9294,N_8751,N_8942);
and U9295 (N_9295,N_8972,N_8798);
nor U9296 (N_9296,N_8772,N_8972);
or U9297 (N_9297,N_8763,N_8824);
xnor U9298 (N_9298,N_8711,N_8865);
or U9299 (N_9299,N_8899,N_8813);
and U9300 (N_9300,N_9158,N_9230);
and U9301 (N_9301,N_9101,N_9252);
nand U9302 (N_9302,N_9105,N_9091);
nand U9303 (N_9303,N_9040,N_9197);
xor U9304 (N_9304,N_9085,N_9056);
nor U9305 (N_9305,N_9275,N_9129);
and U9306 (N_9306,N_9073,N_9015);
and U9307 (N_9307,N_9006,N_9140);
or U9308 (N_9308,N_9164,N_9118);
or U9309 (N_9309,N_9210,N_9179);
and U9310 (N_9310,N_9237,N_9013);
or U9311 (N_9311,N_9251,N_9087);
nand U9312 (N_9312,N_9298,N_9069);
xor U9313 (N_9313,N_9026,N_9176);
or U9314 (N_9314,N_9083,N_9242);
xnor U9315 (N_9315,N_9038,N_9148);
and U9316 (N_9316,N_9020,N_9080);
or U9317 (N_9317,N_9191,N_9059);
or U9318 (N_9318,N_9260,N_9066);
and U9319 (N_9319,N_9103,N_9106);
nor U9320 (N_9320,N_9246,N_9049);
and U9321 (N_9321,N_9084,N_9008);
nor U9322 (N_9322,N_9193,N_9220);
and U9323 (N_9323,N_9181,N_9294);
nor U9324 (N_9324,N_9109,N_9266);
nand U9325 (N_9325,N_9155,N_9007);
nor U9326 (N_9326,N_9009,N_9055);
or U9327 (N_9327,N_9136,N_9258);
nand U9328 (N_9328,N_9272,N_9283);
or U9329 (N_9329,N_9281,N_9172);
nand U9330 (N_9330,N_9153,N_9028);
xnor U9331 (N_9331,N_9088,N_9152);
or U9332 (N_9332,N_9250,N_9057);
nor U9333 (N_9333,N_9295,N_9269);
and U9334 (N_9334,N_9198,N_9174);
xor U9335 (N_9335,N_9003,N_9284);
nor U9336 (N_9336,N_9233,N_9122);
nor U9337 (N_9337,N_9097,N_9139);
nor U9338 (N_9338,N_9192,N_9029);
nor U9339 (N_9339,N_9182,N_9170);
xnor U9340 (N_9340,N_9067,N_9200);
or U9341 (N_9341,N_9257,N_9245);
nor U9342 (N_9342,N_9060,N_9099);
and U9343 (N_9343,N_9188,N_9141);
xnor U9344 (N_9344,N_9162,N_9030);
and U9345 (N_9345,N_9231,N_9157);
and U9346 (N_9346,N_9204,N_9100);
nand U9347 (N_9347,N_9079,N_9282);
or U9348 (N_9348,N_9256,N_9022);
or U9349 (N_9349,N_9286,N_9163);
nand U9350 (N_9350,N_9092,N_9238);
or U9351 (N_9351,N_9019,N_9265);
xor U9352 (N_9352,N_9199,N_9160);
and U9353 (N_9353,N_9119,N_9190);
xnor U9354 (N_9354,N_9063,N_9146);
nor U9355 (N_9355,N_9127,N_9035);
nor U9356 (N_9356,N_9014,N_9223);
or U9357 (N_9357,N_9090,N_9244);
nand U9358 (N_9358,N_9142,N_9229);
or U9359 (N_9359,N_9046,N_9297);
and U9360 (N_9360,N_9065,N_9096);
and U9361 (N_9361,N_9041,N_9051);
xor U9362 (N_9362,N_9267,N_9165);
or U9363 (N_9363,N_9288,N_9262);
xnor U9364 (N_9364,N_9173,N_9205);
xnor U9365 (N_9365,N_9005,N_9023);
nor U9366 (N_9366,N_9017,N_9212);
and U9367 (N_9367,N_9064,N_9075);
nor U9368 (N_9368,N_9135,N_9137);
nand U9369 (N_9369,N_9234,N_9123);
and U9370 (N_9370,N_9226,N_9240);
and U9371 (N_9371,N_9280,N_9243);
or U9372 (N_9372,N_9044,N_9032);
and U9373 (N_9373,N_9249,N_9034);
and U9374 (N_9374,N_9027,N_9228);
or U9375 (N_9375,N_9126,N_9113);
or U9376 (N_9376,N_9048,N_9270);
or U9377 (N_9377,N_9211,N_9293);
xnor U9378 (N_9378,N_9292,N_9068);
xnor U9379 (N_9379,N_9150,N_9130);
nand U9380 (N_9380,N_9254,N_9151);
or U9381 (N_9381,N_9222,N_9112);
nand U9382 (N_9382,N_9183,N_9031);
or U9383 (N_9383,N_9154,N_9241);
nand U9384 (N_9384,N_9248,N_9093);
nor U9385 (N_9385,N_9202,N_9004);
nand U9386 (N_9386,N_9255,N_9070);
nor U9387 (N_9387,N_9052,N_9108);
nand U9388 (N_9388,N_9120,N_9208);
and U9389 (N_9389,N_9061,N_9058);
and U9390 (N_9390,N_9062,N_9121);
xnor U9391 (N_9391,N_9094,N_9116);
nand U9392 (N_9392,N_9102,N_9247);
and U9393 (N_9393,N_9177,N_9268);
and U9394 (N_9394,N_9178,N_9166);
and U9395 (N_9395,N_9232,N_9104);
xor U9396 (N_9396,N_9156,N_9071);
nand U9397 (N_9397,N_9296,N_9081);
and U9398 (N_9398,N_9253,N_9117);
and U9399 (N_9399,N_9147,N_9239);
nor U9400 (N_9400,N_9168,N_9215);
nor U9401 (N_9401,N_9018,N_9145);
or U9402 (N_9402,N_9209,N_9175);
xnor U9403 (N_9403,N_9225,N_9289);
nand U9404 (N_9404,N_9167,N_9125);
and U9405 (N_9405,N_9287,N_9203);
nand U9406 (N_9406,N_9235,N_9050);
xnor U9407 (N_9407,N_9072,N_9276);
and U9408 (N_9408,N_9076,N_9138);
xor U9409 (N_9409,N_9011,N_9277);
xnor U9410 (N_9410,N_9290,N_9033);
xnor U9411 (N_9411,N_9047,N_9264);
xnor U9412 (N_9412,N_9001,N_9201);
xnor U9413 (N_9413,N_9189,N_9124);
and U9414 (N_9414,N_9227,N_9186);
xnor U9415 (N_9415,N_9133,N_9037);
xor U9416 (N_9416,N_9187,N_9213);
xnor U9417 (N_9417,N_9180,N_9131);
xnor U9418 (N_9418,N_9278,N_9086);
nor U9419 (N_9419,N_9236,N_9036);
or U9420 (N_9420,N_9194,N_9074);
or U9421 (N_9421,N_9010,N_9077);
nand U9422 (N_9422,N_9196,N_9111);
xnor U9423 (N_9423,N_9207,N_9043);
or U9424 (N_9424,N_9218,N_9271);
xnor U9425 (N_9425,N_9024,N_9279);
xor U9426 (N_9426,N_9221,N_9114);
and U9427 (N_9427,N_9016,N_9261);
or U9428 (N_9428,N_9285,N_9143);
nor U9429 (N_9429,N_9053,N_9291);
xor U9430 (N_9430,N_9098,N_9144);
nor U9431 (N_9431,N_9002,N_9159);
xnor U9432 (N_9432,N_9128,N_9000);
and U9433 (N_9433,N_9206,N_9042);
nor U9434 (N_9434,N_9219,N_9132);
xnor U9435 (N_9435,N_9195,N_9107);
xor U9436 (N_9436,N_9171,N_9110);
and U9437 (N_9437,N_9095,N_9012);
or U9438 (N_9438,N_9054,N_9224);
nand U9439 (N_9439,N_9299,N_9045);
nor U9440 (N_9440,N_9185,N_9025);
or U9441 (N_9441,N_9078,N_9259);
nor U9442 (N_9442,N_9274,N_9089);
and U9443 (N_9443,N_9263,N_9273);
or U9444 (N_9444,N_9217,N_9134);
xor U9445 (N_9445,N_9149,N_9021);
and U9446 (N_9446,N_9214,N_9082);
nand U9447 (N_9447,N_9161,N_9115);
nor U9448 (N_9448,N_9184,N_9216);
nor U9449 (N_9449,N_9039,N_9169);
nand U9450 (N_9450,N_9261,N_9247);
nor U9451 (N_9451,N_9125,N_9291);
nor U9452 (N_9452,N_9243,N_9287);
xor U9453 (N_9453,N_9233,N_9082);
nand U9454 (N_9454,N_9148,N_9008);
nor U9455 (N_9455,N_9267,N_9090);
nand U9456 (N_9456,N_9148,N_9120);
nand U9457 (N_9457,N_9117,N_9162);
nor U9458 (N_9458,N_9154,N_9029);
xnor U9459 (N_9459,N_9278,N_9251);
xnor U9460 (N_9460,N_9017,N_9290);
nor U9461 (N_9461,N_9062,N_9173);
nor U9462 (N_9462,N_9139,N_9127);
nand U9463 (N_9463,N_9210,N_9145);
nor U9464 (N_9464,N_9267,N_9030);
nand U9465 (N_9465,N_9014,N_9018);
nand U9466 (N_9466,N_9241,N_9094);
or U9467 (N_9467,N_9275,N_9270);
xnor U9468 (N_9468,N_9270,N_9068);
and U9469 (N_9469,N_9076,N_9152);
xor U9470 (N_9470,N_9040,N_9001);
nand U9471 (N_9471,N_9180,N_9064);
and U9472 (N_9472,N_9034,N_9044);
xor U9473 (N_9473,N_9174,N_9196);
and U9474 (N_9474,N_9170,N_9166);
nor U9475 (N_9475,N_9179,N_9147);
nand U9476 (N_9476,N_9277,N_9123);
or U9477 (N_9477,N_9243,N_9091);
or U9478 (N_9478,N_9146,N_9258);
or U9479 (N_9479,N_9031,N_9200);
or U9480 (N_9480,N_9293,N_9126);
and U9481 (N_9481,N_9125,N_9098);
nand U9482 (N_9482,N_9195,N_9053);
or U9483 (N_9483,N_9251,N_9095);
or U9484 (N_9484,N_9299,N_9115);
or U9485 (N_9485,N_9248,N_9037);
xor U9486 (N_9486,N_9126,N_9060);
and U9487 (N_9487,N_9182,N_9052);
xnor U9488 (N_9488,N_9251,N_9028);
xnor U9489 (N_9489,N_9234,N_9182);
and U9490 (N_9490,N_9036,N_9275);
xnor U9491 (N_9491,N_9055,N_9234);
nand U9492 (N_9492,N_9043,N_9041);
and U9493 (N_9493,N_9177,N_9251);
nor U9494 (N_9494,N_9217,N_9242);
or U9495 (N_9495,N_9261,N_9267);
nor U9496 (N_9496,N_9051,N_9175);
nor U9497 (N_9497,N_9055,N_9012);
and U9498 (N_9498,N_9124,N_9083);
xor U9499 (N_9499,N_9171,N_9124);
nand U9500 (N_9500,N_9223,N_9118);
or U9501 (N_9501,N_9266,N_9202);
nand U9502 (N_9502,N_9269,N_9090);
xnor U9503 (N_9503,N_9099,N_9284);
nand U9504 (N_9504,N_9106,N_9214);
or U9505 (N_9505,N_9001,N_9079);
xor U9506 (N_9506,N_9033,N_9161);
nor U9507 (N_9507,N_9033,N_9296);
xnor U9508 (N_9508,N_9108,N_9107);
and U9509 (N_9509,N_9252,N_9163);
xor U9510 (N_9510,N_9284,N_9119);
xor U9511 (N_9511,N_9160,N_9213);
xor U9512 (N_9512,N_9135,N_9005);
or U9513 (N_9513,N_9204,N_9150);
or U9514 (N_9514,N_9276,N_9214);
or U9515 (N_9515,N_9077,N_9252);
nand U9516 (N_9516,N_9232,N_9025);
xnor U9517 (N_9517,N_9128,N_9056);
nor U9518 (N_9518,N_9002,N_9121);
xnor U9519 (N_9519,N_9234,N_9197);
or U9520 (N_9520,N_9116,N_9132);
or U9521 (N_9521,N_9104,N_9239);
or U9522 (N_9522,N_9111,N_9104);
xnor U9523 (N_9523,N_9102,N_9049);
or U9524 (N_9524,N_9148,N_9147);
nand U9525 (N_9525,N_9156,N_9030);
xor U9526 (N_9526,N_9171,N_9138);
nand U9527 (N_9527,N_9163,N_9142);
nor U9528 (N_9528,N_9136,N_9191);
and U9529 (N_9529,N_9257,N_9206);
nand U9530 (N_9530,N_9096,N_9243);
or U9531 (N_9531,N_9261,N_9200);
and U9532 (N_9532,N_9025,N_9168);
nor U9533 (N_9533,N_9152,N_9228);
xor U9534 (N_9534,N_9249,N_9108);
or U9535 (N_9535,N_9031,N_9161);
nand U9536 (N_9536,N_9059,N_9053);
xnor U9537 (N_9537,N_9155,N_9272);
and U9538 (N_9538,N_9131,N_9245);
and U9539 (N_9539,N_9063,N_9260);
nor U9540 (N_9540,N_9269,N_9144);
and U9541 (N_9541,N_9267,N_9059);
or U9542 (N_9542,N_9214,N_9012);
nor U9543 (N_9543,N_9232,N_9208);
nor U9544 (N_9544,N_9289,N_9093);
xnor U9545 (N_9545,N_9108,N_9240);
or U9546 (N_9546,N_9003,N_9050);
xnor U9547 (N_9547,N_9069,N_9112);
and U9548 (N_9548,N_9153,N_9255);
or U9549 (N_9549,N_9026,N_9190);
and U9550 (N_9550,N_9211,N_9009);
and U9551 (N_9551,N_9017,N_9063);
or U9552 (N_9552,N_9271,N_9156);
xnor U9553 (N_9553,N_9150,N_9112);
xor U9554 (N_9554,N_9065,N_9178);
xor U9555 (N_9555,N_9255,N_9256);
xor U9556 (N_9556,N_9129,N_9056);
nor U9557 (N_9557,N_9159,N_9097);
nor U9558 (N_9558,N_9292,N_9213);
nand U9559 (N_9559,N_9250,N_9295);
xor U9560 (N_9560,N_9067,N_9274);
or U9561 (N_9561,N_9086,N_9005);
nor U9562 (N_9562,N_9159,N_9204);
nor U9563 (N_9563,N_9059,N_9127);
nand U9564 (N_9564,N_9018,N_9150);
nor U9565 (N_9565,N_9282,N_9269);
and U9566 (N_9566,N_9038,N_9212);
or U9567 (N_9567,N_9006,N_9274);
xor U9568 (N_9568,N_9290,N_9114);
and U9569 (N_9569,N_9099,N_9035);
xor U9570 (N_9570,N_9175,N_9031);
and U9571 (N_9571,N_9052,N_9028);
xnor U9572 (N_9572,N_9159,N_9137);
and U9573 (N_9573,N_9077,N_9079);
nand U9574 (N_9574,N_9190,N_9046);
nand U9575 (N_9575,N_9125,N_9226);
or U9576 (N_9576,N_9197,N_9105);
nand U9577 (N_9577,N_9121,N_9175);
nor U9578 (N_9578,N_9204,N_9226);
nand U9579 (N_9579,N_9097,N_9075);
and U9580 (N_9580,N_9225,N_9047);
or U9581 (N_9581,N_9273,N_9247);
nand U9582 (N_9582,N_9230,N_9086);
or U9583 (N_9583,N_9003,N_9072);
nand U9584 (N_9584,N_9255,N_9148);
xor U9585 (N_9585,N_9281,N_9080);
and U9586 (N_9586,N_9234,N_9140);
and U9587 (N_9587,N_9122,N_9176);
nand U9588 (N_9588,N_9024,N_9246);
xor U9589 (N_9589,N_9038,N_9183);
xor U9590 (N_9590,N_9201,N_9085);
and U9591 (N_9591,N_9184,N_9138);
nor U9592 (N_9592,N_9261,N_9179);
nand U9593 (N_9593,N_9229,N_9203);
nand U9594 (N_9594,N_9279,N_9256);
xnor U9595 (N_9595,N_9227,N_9209);
xor U9596 (N_9596,N_9177,N_9035);
nand U9597 (N_9597,N_9134,N_9165);
xor U9598 (N_9598,N_9117,N_9144);
nand U9599 (N_9599,N_9193,N_9119);
nand U9600 (N_9600,N_9325,N_9469);
nand U9601 (N_9601,N_9538,N_9352);
nand U9602 (N_9602,N_9332,N_9315);
or U9603 (N_9603,N_9370,N_9560);
nand U9604 (N_9604,N_9443,N_9437);
or U9605 (N_9605,N_9450,N_9458);
and U9606 (N_9606,N_9438,N_9494);
nor U9607 (N_9607,N_9320,N_9564);
xor U9608 (N_9608,N_9574,N_9519);
nor U9609 (N_9609,N_9527,N_9484);
xnor U9610 (N_9610,N_9451,N_9379);
or U9611 (N_9611,N_9403,N_9361);
xor U9612 (N_9612,N_9595,N_9313);
nand U9613 (N_9613,N_9396,N_9512);
or U9614 (N_9614,N_9553,N_9517);
or U9615 (N_9615,N_9504,N_9501);
xor U9616 (N_9616,N_9580,N_9555);
xnor U9617 (N_9617,N_9552,N_9535);
xnor U9618 (N_9618,N_9427,N_9529);
or U9619 (N_9619,N_9426,N_9369);
and U9620 (N_9620,N_9497,N_9373);
or U9621 (N_9621,N_9586,N_9544);
nand U9622 (N_9622,N_9381,N_9360);
nor U9623 (N_9623,N_9337,N_9387);
nand U9624 (N_9624,N_9431,N_9404);
and U9625 (N_9625,N_9490,N_9408);
or U9626 (N_9626,N_9333,N_9572);
nand U9627 (N_9627,N_9472,N_9323);
or U9628 (N_9628,N_9415,N_9353);
and U9629 (N_9629,N_9356,N_9465);
and U9630 (N_9630,N_9423,N_9392);
xnor U9631 (N_9631,N_9375,N_9319);
nand U9632 (N_9632,N_9336,N_9406);
or U9633 (N_9633,N_9581,N_9471);
xnor U9634 (N_9634,N_9479,N_9347);
nor U9635 (N_9635,N_9433,N_9416);
or U9636 (N_9636,N_9329,N_9314);
nor U9637 (N_9637,N_9418,N_9350);
nor U9638 (N_9638,N_9513,N_9394);
nor U9639 (N_9639,N_9478,N_9410);
or U9640 (N_9640,N_9578,N_9341);
nand U9641 (N_9641,N_9358,N_9326);
and U9642 (N_9642,N_9594,N_9597);
or U9643 (N_9643,N_9533,N_9598);
or U9644 (N_9644,N_9317,N_9429);
nor U9645 (N_9645,N_9354,N_9474);
xor U9646 (N_9646,N_9335,N_9521);
nor U9647 (N_9647,N_9412,N_9436);
or U9648 (N_9648,N_9508,N_9328);
or U9649 (N_9649,N_9346,N_9321);
nor U9650 (N_9650,N_9435,N_9434);
nand U9651 (N_9651,N_9561,N_9393);
nor U9652 (N_9652,N_9491,N_9349);
nand U9653 (N_9653,N_9587,N_9308);
or U9654 (N_9654,N_9417,N_9300);
nor U9655 (N_9655,N_9307,N_9330);
and U9656 (N_9656,N_9331,N_9540);
xnor U9657 (N_9657,N_9562,N_9445);
or U9658 (N_9658,N_9407,N_9316);
and U9659 (N_9659,N_9411,N_9523);
xnor U9660 (N_9660,N_9481,N_9419);
nor U9661 (N_9661,N_9441,N_9453);
or U9662 (N_9662,N_9596,N_9505);
or U9663 (N_9663,N_9312,N_9367);
xnor U9664 (N_9664,N_9537,N_9592);
xor U9665 (N_9665,N_9386,N_9391);
or U9666 (N_9666,N_9455,N_9304);
xor U9667 (N_9667,N_9444,N_9591);
nand U9668 (N_9668,N_9382,N_9351);
and U9669 (N_9669,N_9534,N_9452);
and U9670 (N_9670,N_9301,N_9302);
xor U9671 (N_9671,N_9510,N_9524);
xor U9672 (N_9672,N_9390,N_9520);
or U9673 (N_9673,N_9547,N_9432);
xnor U9674 (N_9674,N_9364,N_9528);
or U9675 (N_9675,N_9460,N_9480);
nand U9676 (N_9676,N_9327,N_9475);
xor U9677 (N_9677,N_9464,N_9448);
nor U9678 (N_9678,N_9339,N_9402);
or U9679 (N_9679,N_9357,N_9593);
nand U9680 (N_9680,N_9377,N_9362);
nor U9681 (N_9681,N_9371,N_9470);
or U9682 (N_9682,N_9495,N_9548);
nand U9683 (N_9683,N_9509,N_9384);
nor U9684 (N_9684,N_9368,N_9563);
xnor U9685 (N_9685,N_9483,N_9305);
or U9686 (N_9686,N_9456,N_9549);
xor U9687 (N_9687,N_9522,N_9303);
or U9688 (N_9688,N_9543,N_9311);
xor U9689 (N_9689,N_9401,N_9421);
nand U9690 (N_9690,N_9345,N_9467);
xnor U9691 (N_9691,N_9439,N_9388);
nand U9692 (N_9692,N_9589,N_9590);
xnor U9693 (N_9693,N_9468,N_9568);
and U9694 (N_9694,N_9420,N_9556);
nand U9695 (N_9695,N_9366,N_9338);
nand U9696 (N_9696,N_9503,N_9385);
xnor U9697 (N_9697,N_9372,N_9461);
nand U9698 (N_9698,N_9343,N_9511);
and U9699 (N_9699,N_9506,N_9395);
xor U9700 (N_9700,N_9526,N_9342);
xnor U9701 (N_9701,N_9536,N_9447);
nand U9702 (N_9702,N_9584,N_9378);
or U9703 (N_9703,N_9422,N_9355);
nor U9704 (N_9704,N_9348,N_9565);
nand U9705 (N_9705,N_9413,N_9551);
and U9706 (N_9706,N_9324,N_9488);
xnor U9707 (N_9707,N_9399,N_9566);
or U9708 (N_9708,N_9485,N_9365);
and U9709 (N_9709,N_9486,N_9489);
nand U9710 (N_9710,N_9430,N_9516);
nor U9711 (N_9711,N_9459,N_9310);
xor U9712 (N_9712,N_9477,N_9567);
and U9713 (N_9713,N_9466,N_9463);
or U9714 (N_9714,N_9500,N_9554);
and U9715 (N_9715,N_9577,N_9583);
xnor U9716 (N_9716,N_9473,N_9454);
nor U9717 (N_9717,N_9359,N_9446);
or U9718 (N_9718,N_9409,N_9424);
and U9719 (N_9719,N_9405,N_9492);
and U9720 (N_9720,N_9531,N_9318);
nand U9721 (N_9721,N_9414,N_9340);
nand U9722 (N_9722,N_9542,N_9462);
nor U9723 (N_9723,N_9425,N_9398);
or U9724 (N_9724,N_9493,N_9571);
nand U9725 (N_9725,N_9334,N_9374);
nor U9726 (N_9726,N_9557,N_9309);
xnor U9727 (N_9727,N_9363,N_9502);
nand U9728 (N_9728,N_9440,N_9442);
nand U9729 (N_9729,N_9579,N_9532);
xnor U9730 (N_9730,N_9482,N_9476);
nand U9731 (N_9731,N_9545,N_9400);
or U9732 (N_9732,N_9573,N_9582);
nand U9733 (N_9733,N_9507,N_9499);
xor U9734 (N_9734,N_9496,N_9397);
xnor U9735 (N_9735,N_9515,N_9306);
nand U9736 (N_9736,N_9383,N_9376);
and U9737 (N_9737,N_9498,N_9569);
nand U9738 (N_9738,N_9550,N_9558);
and U9739 (N_9739,N_9570,N_9530);
nand U9740 (N_9740,N_9546,N_9487);
nand U9741 (N_9741,N_9576,N_9457);
and U9742 (N_9742,N_9380,N_9585);
nand U9743 (N_9743,N_9428,N_9449);
and U9744 (N_9744,N_9322,N_9518);
nand U9745 (N_9745,N_9575,N_9525);
xnor U9746 (N_9746,N_9539,N_9344);
or U9747 (N_9747,N_9599,N_9389);
nor U9748 (N_9748,N_9588,N_9514);
nand U9749 (N_9749,N_9559,N_9541);
and U9750 (N_9750,N_9455,N_9480);
xnor U9751 (N_9751,N_9363,N_9537);
or U9752 (N_9752,N_9310,N_9484);
nand U9753 (N_9753,N_9535,N_9540);
xnor U9754 (N_9754,N_9433,N_9513);
xor U9755 (N_9755,N_9372,N_9355);
nor U9756 (N_9756,N_9456,N_9472);
nand U9757 (N_9757,N_9471,N_9510);
nand U9758 (N_9758,N_9587,N_9352);
nor U9759 (N_9759,N_9572,N_9353);
nor U9760 (N_9760,N_9352,N_9338);
or U9761 (N_9761,N_9428,N_9562);
xor U9762 (N_9762,N_9551,N_9301);
and U9763 (N_9763,N_9499,N_9522);
xnor U9764 (N_9764,N_9332,N_9482);
nand U9765 (N_9765,N_9443,N_9430);
nand U9766 (N_9766,N_9396,N_9552);
xor U9767 (N_9767,N_9305,N_9350);
nor U9768 (N_9768,N_9521,N_9312);
xor U9769 (N_9769,N_9318,N_9360);
xor U9770 (N_9770,N_9413,N_9347);
nor U9771 (N_9771,N_9313,N_9421);
xor U9772 (N_9772,N_9532,N_9369);
and U9773 (N_9773,N_9465,N_9440);
and U9774 (N_9774,N_9596,N_9362);
and U9775 (N_9775,N_9451,N_9398);
and U9776 (N_9776,N_9300,N_9533);
nand U9777 (N_9777,N_9501,N_9471);
xor U9778 (N_9778,N_9377,N_9593);
and U9779 (N_9779,N_9586,N_9527);
xnor U9780 (N_9780,N_9320,N_9436);
xor U9781 (N_9781,N_9493,N_9575);
or U9782 (N_9782,N_9496,N_9380);
or U9783 (N_9783,N_9504,N_9583);
and U9784 (N_9784,N_9309,N_9536);
and U9785 (N_9785,N_9472,N_9311);
nor U9786 (N_9786,N_9468,N_9587);
and U9787 (N_9787,N_9536,N_9367);
nor U9788 (N_9788,N_9411,N_9359);
xor U9789 (N_9789,N_9395,N_9528);
or U9790 (N_9790,N_9328,N_9391);
nor U9791 (N_9791,N_9474,N_9571);
and U9792 (N_9792,N_9359,N_9504);
or U9793 (N_9793,N_9346,N_9594);
xnor U9794 (N_9794,N_9560,N_9493);
xnor U9795 (N_9795,N_9370,N_9467);
nand U9796 (N_9796,N_9569,N_9521);
or U9797 (N_9797,N_9494,N_9422);
and U9798 (N_9798,N_9367,N_9539);
or U9799 (N_9799,N_9401,N_9428);
nor U9800 (N_9800,N_9587,N_9397);
nand U9801 (N_9801,N_9383,N_9524);
and U9802 (N_9802,N_9539,N_9444);
xor U9803 (N_9803,N_9459,N_9499);
and U9804 (N_9804,N_9542,N_9310);
xnor U9805 (N_9805,N_9393,N_9335);
or U9806 (N_9806,N_9345,N_9375);
nor U9807 (N_9807,N_9397,N_9497);
xor U9808 (N_9808,N_9525,N_9568);
xor U9809 (N_9809,N_9548,N_9375);
nand U9810 (N_9810,N_9330,N_9358);
or U9811 (N_9811,N_9320,N_9332);
and U9812 (N_9812,N_9564,N_9400);
nor U9813 (N_9813,N_9340,N_9418);
nor U9814 (N_9814,N_9500,N_9499);
nor U9815 (N_9815,N_9502,N_9493);
nand U9816 (N_9816,N_9590,N_9555);
nor U9817 (N_9817,N_9363,N_9491);
or U9818 (N_9818,N_9395,N_9341);
or U9819 (N_9819,N_9564,N_9318);
nand U9820 (N_9820,N_9598,N_9418);
xor U9821 (N_9821,N_9323,N_9403);
nand U9822 (N_9822,N_9369,N_9586);
nand U9823 (N_9823,N_9566,N_9571);
nor U9824 (N_9824,N_9440,N_9357);
nor U9825 (N_9825,N_9488,N_9445);
or U9826 (N_9826,N_9396,N_9341);
and U9827 (N_9827,N_9306,N_9545);
and U9828 (N_9828,N_9357,N_9386);
nor U9829 (N_9829,N_9413,N_9545);
and U9830 (N_9830,N_9309,N_9541);
xnor U9831 (N_9831,N_9379,N_9385);
and U9832 (N_9832,N_9380,N_9591);
or U9833 (N_9833,N_9568,N_9413);
nand U9834 (N_9834,N_9400,N_9450);
xor U9835 (N_9835,N_9477,N_9301);
or U9836 (N_9836,N_9302,N_9307);
nor U9837 (N_9837,N_9500,N_9571);
nand U9838 (N_9838,N_9405,N_9382);
and U9839 (N_9839,N_9439,N_9370);
or U9840 (N_9840,N_9557,N_9342);
nor U9841 (N_9841,N_9460,N_9386);
nand U9842 (N_9842,N_9341,N_9477);
and U9843 (N_9843,N_9372,N_9416);
or U9844 (N_9844,N_9406,N_9537);
or U9845 (N_9845,N_9541,N_9362);
nor U9846 (N_9846,N_9500,N_9439);
xor U9847 (N_9847,N_9581,N_9469);
or U9848 (N_9848,N_9392,N_9550);
xor U9849 (N_9849,N_9466,N_9538);
xor U9850 (N_9850,N_9542,N_9514);
xor U9851 (N_9851,N_9495,N_9457);
nor U9852 (N_9852,N_9443,N_9408);
xor U9853 (N_9853,N_9308,N_9338);
nand U9854 (N_9854,N_9331,N_9407);
nor U9855 (N_9855,N_9337,N_9397);
nor U9856 (N_9856,N_9366,N_9469);
xor U9857 (N_9857,N_9531,N_9437);
and U9858 (N_9858,N_9445,N_9426);
xnor U9859 (N_9859,N_9451,N_9485);
nor U9860 (N_9860,N_9506,N_9423);
nand U9861 (N_9861,N_9469,N_9328);
xnor U9862 (N_9862,N_9532,N_9481);
xnor U9863 (N_9863,N_9522,N_9519);
xor U9864 (N_9864,N_9332,N_9457);
nor U9865 (N_9865,N_9334,N_9333);
nand U9866 (N_9866,N_9327,N_9402);
and U9867 (N_9867,N_9308,N_9390);
nor U9868 (N_9868,N_9550,N_9541);
xnor U9869 (N_9869,N_9358,N_9560);
and U9870 (N_9870,N_9499,N_9539);
and U9871 (N_9871,N_9476,N_9538);
nor U9872 (N_9872,N_9446,N_9539);
or U9873 (N_9873,N_9397,N_9560);
xor U9874 (N_9874,N_9531,N_9388);
nand U9875 (N_9875,N_9327,N_9434);
nor U9876 (N_9876,N_9574,N_9476);
nand U9877 (N_9877,N_9499,N_9544);
xor U9878 (N_9878,N_9302,N_9536);
nand U9879 (N_9879,N_9402,N_9591);
and U9880 (N_9880,N_9558,N_9594);
or U9881 (N_9881,N_9462,N_9530);
or U9882 (N_9882,N_9540,N_9597);
nand U9883 (N_9883,N_9542,N_9384);
and U9884 (N_9884,N_9499,N_9528);
and U9885 (N_9885,N_9334,N_9342);
or U9886 (N_9886,N_9334,N_9397);
and U9887 (N_9887,N_9433,N_9534);
xor U9888 (N_9888,N_9402,N_9522);
or U9889 (N_9889,N_9417,N_9516);
nor U9890 (N_9890,N_9454,N_9363);
or U9891 (N_9891,N_9486,N_9501);
and U9892 (N_9892,N_9429,N_9465);
xnor U9893 (N_9893,N_9553,N_9523);
and U9894 (N_9894,N_9504,N_9388);
nand U9895 (N_9895,N_9480,N_9443);
nand U9896 (N_9896,N_9450,N_9366);
xnor U9897 (N_9897,N_9571,N_9594);
or U9898 (N_9898,N_9480,N_9560);
xor U9899 (N_9899,N_9573,N_9391);
nor U9900 (N_9900,N_9689,N_9736);
xor U9901 (N_9901,N_9677,N_9723);
xor U9902 (N_9902,N_9665,N_9766);
nor U9903 (N_9903,N_9806,N_9738);
and U9904 (N_9904,N_9732,N_9747);
or U9905 (N_9905,N_9785,N_9618);
xor U9906 (N_9906,N_9840,N_9722);
and U9907 (N_9907,N_9740,N_9894);
or U9908 (N_9908,N_9849,N_9694);
xnor U9909 (N_9909,N_9892,N_9811);
xor U9910 (N_9910,N_9782,N_9667);
or U9911 (N_9911,N_9824,N_9690);
nand U9912 (N_9912,N_9706,N_9854);
and U9913 (N_9913,N_9749,N_9669);
and U9914 (N_9914,N_9695,N_9674);
or U9915 (N_9915,N_9767,N_9726);
nor U9916 (N_9916,N_9636,N_9693);
nand U9917 (N_9917,N_9872,N_9897);
nand U9918 (N_9918,N_9691,N_9616);
and U9919 (N_9919,N_9875,N_9713);
xnor U9920 (N_9920,N_9896,N_9720);
and U9921 (N_9921,N_9705,N_9868);
nor U9922 (N_9922,N_9680,N_9630);
or U9923 (N_9923,N_9818,N_9718);
xnor U9924 (N_9924,N_9790,N_9735);
and U9925 (N_9925,N_9654,N_9804);
xnor U9926 (N_9926,N_9893,N_9859);
nor U9927 (N_9927,N_9681,N_9675);
nor U9928 (N_9928,N_9870,N_9865);
and U9929 (N_9929,N_9710,N_9881);
nor U9930 (N_9930,N_9627,N_9628);
and U9931 (N_9931,N_9678,N_9823);
or U9932 (N_9932,N_9838,N_9728);
xnor U9933 (N_9933,N_9753,N_9679);
nand U9934 (N_9934,N_9642,N_9692);
and U9935 (N_9935,N_9602,N_9676);
and U9936 (N_9936,N_9714,N_9653);
nor U9937 (N_9937,N_9891,N_9787);
nand U9938 (N_9938,N_9709,N_9621);
nor U9939 (N_9939,N_9671,N_9883);
nor U9940 (N_9940,N_9834,N_9808);
or U9941 (N_9941,N_9762,N_9833);
nor U9942 (N_9942,N_9827,N_9741);
and U9943 (N_9943,N_9719,N_9622);
xnor U9944 (N_9944,N_9615,N_9794);
and U9945 (N_9945,N_9686,N_9770);
nand U9946 (N_9946,N_9876,N_9848);
xor U9947 (N_9947,N_9874,N_9898);
or U9948 (N_9948,N_9668,N_9845);
nand U9949 (N_9949,N_9605,N_9700);
nor U9950 (N_9950,N_9841,N_9836);
xnor U9951 (N_9951,N_9776,N_9864);
and U9952 (N_9952,N_9816,N_9708);
nor U9953 (N_9953,N_9842,N_9620);
and U9954 (N_9954,N_9717,N_9660);
or U9955 (N_9955,N_9743,N_9635);
nand U9956 (N_9956,N_9814,N_9604);
and U9957 (N_9957,N_9666,N_9822);
or U9958 (N_9958,N_9869,N_9831);
xnor U9959 (N_9959,N_9886,N_9895);
nor U9960 (N_9960,N_9798,N_9637);
xnor U9961 (N_9961,N_9853,N_9832);
nor U9962 (N_9962,N_9796,N_9783);
nand U9963 (N_9963,N_9737,N_9803);
nand U9964 (N_9964,N_9711,N_9861);
nor U9965 (N_9965,N_9880,N_9752);
or U9966 (N_9966,N_9884,N_9825);
and U9967 (N_9967,N_9820,N_9855);
xor U9968 (N_9968,N_9611,N_9657);
and U9969 (N_9969,N_9744,N_9843);
nand U9970 (N_9970,N_9704,N_9813);
nand U9971 (N_9971,N_9867,N_9658);
nor U9972 (N_9972,N_9769,N_9651);
and U9973 (N_9973,N_9670,N_9756);
nor U9974 (N_9974,N_9850,N_9606);
xor U9975 (N_9975,N_9697,N_9812);
nor U9976 (N_9976,N_9879,N_9885);
xor U9977 (N_9977,N_9858,N_9638);
and U9978 (N_9978,N_9707,N_9648);
or U9979 (N_9979,N_9779,N_9784);
and U9980 (N_9980,N_9647,N_9712);
nor U9981 (N_9981,N_9634,N_9742);
nand U9982 (N_9982,N_9751,N_9835);
nor U9983 (N_9983,N_9830,N_9807);
or U9984 (N_9984,N_9768,N_9729);
and U9985 (N_9985,N_9629,N_9765);
xor U9986 (N_9986,N_9600,N_9809);
nand U9987 (N_9987,N_9801,N_9847);
or U9988 (N_9988,N_9758,N_9890);
and U9989 (N_9989,N_9640,N_9655);
nor U9990 (N_9990,N_9778,N_9791);
nand U9991 (N_9991,N_9727,N_9601);
and U9992 (N_9992,N_9702,N_9802);
nand U9993 (N_9993,N_9703,N_9795);
and U9994 (N_9994,N_9805,N_9613);
and U9995 (N_9995,N_9641,N_9750);
nor U9996 (N_9996,N_9672,N_9773);
xor U9997 (N_9997,N_9856,N_9746);
or U9998 (N_9998,N_9715,N_9788);
or U9999 (N_9999,N_9873,N_9661);
and U10000 (N_10000,N_9772,N_9698);
nand U10001 (N_10001,N_9644,N_9817);
or U10002 (N_10002,N_9828,N_9650);
nand U10003 (N_10003,N_9757,N_9730);
or U10004 (N_10004,N_9739,N_9781);
nand U10005 (N_10005,N_9839,N_9780);
nand U10006 (N_10006,N_9610,N_9731);
or U10007 (N_10007,N_9725,N_9878);
and U10008 (N_10008,N_9862,N_9761);
or U10009 (N_10009,N_9685,N_9664);
xor U10010 (N_10010,N_9643,N_9877);
xnor U10011 (N_10011,N_9759,N_9748);
nand U10012 (N_10012,N_9624,N_9649);
nor U10013 (N_10013,N_9774,N_9734);
and U10014 (N_10014,N_9603,N_9721);
nor U10015 (N_10015,N_9701,N_9777);
or U10016 (N_10016,N_9646,N_9846);
nand U10017 (N_10017,N_9716,N_9754);
or U10018 (N_10018,N_9626,N_9612);
nand U10019 (N_10019,N_9607,N_9829);
nor U10020 (N_10020,N_9888,N_9887);
nor U10021 (N_10021,N_9863,N_9682);
xor U10022 (N_10022,N_9793,N_9889);
or U10023 (N_10023,N_9652,N_9683);
xnor U10024 (N_10024,N_9687,N_9851);
or U10025 (N_10025,N_9819,N_9662);
nand U10026 (N_10026,N_9786,N_9815);
xnor U10027 (N_10027,N_9631,N_9837);
nor U10028 (N_10028,N_9775,N_9724);
and U10029 (N_10029,N_9800,N_9755);
xnor U10030 (N_10030,N_9771,N_9645);
nor U10031 (N_10031,N_9639,N_9609);
nand U10032 (N_10032,N_9899,N_9614);
xnor U10033 (N_10033,N_9684,N_9871);
or U10034 (N_10034,N_9821,N_9633);
nor U10035 (N_10035,N_9623,N_9760);
and U10036 (N_10036,N_9764,N_9882);
xor U10037 (N_10037,N_9797,N_9826);
nand U10038 (N_10038,N_9663,N_9763);
nor U10039 (N_10039,N_9659,N_9852);
xor U10040 (N_10040,N_9844,N_9688);
or U10041 (N_10041,N_9789,N_9799);
nand U10042 (N_10042,N_9792,N_9632);
nor U10043 (N_10043,N_9733,N_9860);
nor U10044 (N_10044,N_9866,N_9617);
xor U10045 (N_10045,N_9656,N_9608);
or U10046 (N_10046,N_9625,N_9619);
xor U10047 (N_10047,N_9810,N_9857);
xnor U10048 (N_10048,N_9696,N_9699);
nand U10049 (N_10049,N_9673,N_9745);
xor U10050 (N_10050,N_9833,N_9781);
xor U10051 (N_10051,N_9752,N_9712);
nor U10052 (N_10052,N_9727,N_9635);
nor U10053 (N_10053,N_9756,N_9675);
or U10054 (N_10054,N_9726,N_9741);
xnor U10055 (N_10055,N_9679,N_9840);
or U10056 (N_10056,N_9840,N_9838);
and U10057 (N_10057,N_9714,N_9875);
nand U10058 (N_10058,N_9660,N_9624);
or U10059 (N_10059,N_9604,N_9724);
nand U10060 (N_10060,N_9729,N_9814);
nand U10061 (N_10061,N_9742,N_9728);
nor U10062 (N_10062,N_9822,N_9801);
xor U10063 (N_10063,N_9616,N_9898);
or U10064 (N_10064,N_9727,N_9661);
or U10065 (N_10065,N_9680,N_9828);
xnor U10066 (N_10066,N_9849,N_9852);
and U10067 (N_10067,N_9804,N_9768);
xnor U10068 (N_10068,N_9830,N_9785);
nor U10069 (N_10069,N_9676,N_9700);
and U10070 (N_10070,N_9831,N_9736);
nand U10071 (N_10071,N_9886,N_9877);
and U10072 (N_10072,N_9705,N_9866);
nor U10073 (N_10073,N_9642,N_9730);
nor U10074 (N_10074,N_9733,N_9785);
nand U10075 (N_10075,N_9628,N_9617);
or U10076 (N_10076,N_9711,N_9697);
or U10077 (N_10077,N_9870,N_9620);
or U10078 (N_10078,N_9634,N_9664);
xnor U10079 (N_10079,N_9827,N_9723);
or U10080 (N_10080,N_9794,N_9839);
xor U10081 (N_10081,N_9818,N_9603);
nor U10082 (N_10082,N_9653,N_9828);
nand U10083 (N_10083,N_9754,N_9626);
and U10084 (N_10084,N_9646,N_9869);
xor U10085 (N_10085,N_9827,N_9861);
nand U10086 (N_10086,N_9832,N_9645);
xor U10087 (N_10087,N_9611,N_9860);
xor U10088 (N_10088,N_9705,N_9810);
nand U10089 (N_10089,N_9730,N_9816);
nand U10090 (N_10090,N_9884,N_9751);
nor U10091 (N_10091,N_9838,N_9702);
nor U10092 (N_10092,N_9638,N_9720);
nor U10093 (N_10093,N_9716,N_9759);
and U10094 (N_10094,N_9728,N_9765);
and U10095 (N_10095,N_9757,N_9623);
nand U10096 (N_10096,N_9813,N_9622);
nand U10097 (N_10097,N_9812,N_9771);
nand U10098 (N_10098,N_9638,N_9669);
nor U10099 (N_10099,N_9842,N_9826);
xnor U10100 (N_10100,N_9792,N_9633);
and U10101 (N_10101,N_9813,N_9694);
and U10102 (N_10102,N_9670,N_9715);
nand U10103 (N_10103,N_9827,N_9784);
or U10104 (N_10104,N_9818,N_9828);
nand U10105 (N_10105,N_9869,N_9884);
and U10106 (N_10106,N_9675,N_9724);
nand U10107 (N_10107,N_9670,N_9850);
nand U10108 (N_10108,N_9715,N_9684);
nand U10109 (N_10109,N_9891,N_9779);
and U10110 (N_10110,N_9718,N_9875);
or U10111 (N_10111,N_9707,N_9602);
and U10112 (N_10112,N_9871,N_9623);
nand U10113 (N_10113,N_9885,N_9741);
nand U10114 (N_10114,N_9693,N_9898);
and U10115 (N_10115,N_9834,N_9851);
xor U10116 (N_10116,N_9741,N_9645);
nor U10117 (N_10117,N_9857,N_9849);
and U10118 (N_10118,N_9816,N_9628);
nor U10119 (N_10119,N_9752,N_9804);
nand U10120 (N_10120,N_9851,N_9603);
xnor U10121 (N_10121,N_9879,N_9610);
xnor U10122 (N_10122,N_9806,N_9699);
nor U10123 (N_10123,N_9814,N_9807);
nand U10124 (N_10124,N_9632,N_9876);
and U10125 (N_10125,N_9873,N_9687);
nor U10126 (N_10126,N_9834,N_9832);
and U10127 (N_10127,N_9660,N_9845);
and U10128 (N_10128,N_9621,N_9720);
and U10129 (N_10129,N_9643,N_9677);
and U10130 (N_10130,N_9897,N_9778);
xnor U10131 (N_10131,N_9696,N_9660);
and U10132 (N_10132,N_9627,N_9825);
and U10133 (N_10133,N_9834,N_9607);
and U10134 (N_10134,N_9896,N_9863);
nand U10135 (N_10135,N_9805,N_9701);
and U10136 (N_10136,N_9838,N_9800);
and U10137 (N_10137,N_9784,N_9602);
and U10138 (N_10138,N_9764,N_9738);
and U10139 (N_10139,N_9647,N_9859);
nor U10140 (N_10140,N_9897,N_9719);
nand U10141 (N_10141,N_9610,N_9651);
nand U10142 (N_10142,N_9770,N_9644);
nor U10143 (N_10143,N_9714,N_9845);
nor U10144 (N_10144,N_9764,N_9774);
nor U10145 (N_10145,N_9740,N_9899);
xor U10146 (N_10146,N_9713,N_9867);
xnor U10147 (N_10147,N_9605,N_9845);
and U10148 (N_10148,N_9860,N_9789);
nor U10149 (N_10149,N_9814,N_9853);
nand U10150 (N_10150,N_9717,N_9718);
nand U10151 (N_10151,N_9884,N_9712);
nand U10152 (N_10152,N_9741,N_9671);
nand U10153 (N_10153,N_9729,N_9715);
nor U10154 (N_10154,N_9806,N_9770);
or U10155 (N_10155,N_9793,N_9841);
and U10156 (N_10156,N_9646,N_9677);
and U10157 (N_10157,N_9769,N_9753);
nor U10158 (N_10158,N_9786,N_9661);
xnor U10159 (N_10159,N_9616,N_9640);
xor U10160 (N_10160,N_9797,N_9791);
and U10161 (N_10161,N_9685,N_9714);
xnor U10162 (N_10162,N_9864,N_9663);
nor U10163 (N_10163,N_9832,N_9810);
and U10164 (N_10164,N_9759,N_9619);
xnor U10165 (N_10165,N_9857,N_9866);
nor U10166 (N_10166,N_9873,N_9733);
or U10167 (N_10167,N_9803,N_9656);
nor U10168 (N_10168,N_9629,N_9894);
xor U10169 (N_10169,N_9602,N_9630);
nand U10170 (N_10170,N_9701,N_9882);
nand U10171 (N_10171,N_9850,N_9684);
or U10172 (N_10172,N_9762,N_9679);
and U10173 (N_10173,N_9810,N_9667);
xnor U10174 (N_10174,N_9755,N_9813);
nor U10175 (N_10175,N_9873,N_9858);
xor U10176 (N_10176,N_9819,N_9862);
nand U10177 (N_10177,N_9846,N_9712);
and U10178 (N_10178,N_9604,N_9614);
nor U10179 (N_10179,N_9708,N_9656);
xor U10180 (N_10180,N_9632,N_9754);
nand U10181 (N_10181,N_9747,N_9641);
or U10182 (N_10182,N_9814,N_9676);
or U10183 (N_10183,N_9694,N_9612);
and U10184 (N_10184,N_9868,N_9628);
nor U10185 (N_10185,N_9766,N_9875);
or U10186 (N_10186,N_9600,N_9738);
and U10187 (N_10187,N_9868,N_9741);
and U10188 (N_10188,N_9744,N_9633);
nor U10189 (N_10189,N_9665,N_9849);
nor U10190 (N_10190,N_9845,N_9872);
xor U10191 (N_10191,N_9689,N_9774);
nand U10192 (N_10192,N_9776,N_9649);
and U10193 (N_10193,N_9761,N_9745);
nand U10194 (N_10194,N_9866,N_9782);
nand U10195 (N_10195,N_9655,N_9813);
nand U10196 (N_10196,N_9828,N_9717);
and U10197 (N_10197,N_9854,N_9699);
nor U10198 (N_10198,N_9628,N_9805);
xnor U10199 (N_10199,N_9831,N_9862);
xnor U10200 (N_10200,N_10091,N_10184);
or U10201 (N_10201,N_9955,N_10089);
xor U10202 (N_10202,N_10194,N_10067);
and U10203 (N_10203,N_10077,N_9997);
xnor U10204 (N_10204,N_9908,N_9935);
xor U10205 (N_10205,N_10008,N_9918);
and U10206 (N_10206,N_10095,N_9901);
xnor U10207 (N_10207,N_9968,N_9970);
xnor U10208 (N_10208,N_10148,N_10144);
nand U10209 (N_10209,N_9957,N_10103);
and U10210 (N_10210,N_10139,N_10051);
nor U10211 (N_10211,N_9939,N_9911);
xnor U10212 (N_10212,N_10141,N_9927);
nor U10213 (N_10213,N_9921,N_9941);
or U10214 (N_10214,N_10004,N_9906);
nand U10215 (N_10215,N_10080,N_10136);
and U10216 (N_10216,N_10185,N_9948);
xor U10217 (N_10217,N_10199,N_10150);
nand U10218 (N_10218,N_10035,N_9987);
nor U10219 (N_10219,N_10181,N_10132);
and U10220 (N_10220,N_9949,N_10093);
and U10221 (N_10221,N_10134,N_10063);
nand U10222 (N_10222,N_10171,N_9936);
or U10223 (N_10223,N_10085,N_9933);
nand U10224 (N_10224,N_10078,N_9914);
and U10225 (N_10225,N_10118,N_10043);
and U10226 (N_10226,N_10005,N_9972);
or U10227 (N_10227,N_9903,N_10092);
and U10228 (N_10228,N_9990,N_10086);
nor U10229 (N_10229,N_9980,N_9938);
or U10230 (N_10230,N_10082,N_10117);
nor U10231 (N_10231,N_10022,N_10119);
or U10232 (N_10232,N_10129,N_10057);
and U10233 (N_10233,N_10017,N_10110);
or U10234 (N_10234,N_9964,N_9996);
nor U10235 (N_10235,N_9985,N_10153);
nor U10236 (N_10236,N_10161,N_10042);
nand U10237 (N_10237,N_10099,N_10052);
nand U10238 (N_10238,N_10100,N_9913);
or U10239 (N_10239,N_9988,N_10021);
nand U10240 (N_10240,N_9925,N_10047);
and U10241 (N_10241,N_9969,N_10124);
and U10242 (N_10242,N_10176,N_9954);
or U10243 (N_10243,N_9962,N_10106);
xor U10244 (N_10244,N_10175,N_9993);
and U10245 (N_10245,N_10088,N_10104);
or U10246 (N_10246,N_10019,N_9909);
and U10247 (N_10247,N_9930,N_10115);
and U10248 (N_10248,N_10002,N_10174);
nand U10249 (N_10249,N_10135,N_10112);
and U10250 (N_10250,N_9944,N_9934);
or U10251 (N_10251,N_9951,N_10189);
or U10252 (N_10252,N_9994,N_10036);
nor U10253 (N_10253,N_10000,N_9940);
or U10254 (N_10254,N_9977,N_10101);
nor U10255 (N_10255,N_10169,N_10123);
nand U10256 (N_10256,N_9942,N_10127);
or U10257 (N_10257,N_10108,N_9971);
or U10258 (N_10258,N_10071,N_9960);
and U10259 (N_10259,N_10128,N_10041);
and U10260 (N_10260,N_10162,N_10030);
nand U10261 (N_10261,N_9947,N_10152);
or U10262 (N_10262,N_10014,N_9963);
or U10263 (N_10263,N_10087,N_10040);
or U10264 (N_10264,N_9979,N_10061);
nor U10265 (N_10265,N_9943,N_9950);
or U10266 (N_10266,N_10191,N_10186);
xnor U10267 (N_10267,N_10049,N_10183);
or U10268 (N_10268,N_10156,N_10166);
xor U10269 (N_10269,N_10026,N_10146);
xor U10270 (N_10270,N_9961,N_10125);
nand U10271 (N_10271,N_10151,N_10034);
nand U10272 (N_10272,N_9975,N_9917);
nor U10273 (N_10273,N_10037,N_10193);
xor U10274 (N_10274,N_10032,N_10066);
and U10275 (N_10275,N_10094,N_10168);
or U10276 (N_10276,N_9976,N_10160);
or U10277 (N_10277,N_10053,N_10016);
nor U10278 (N_10278,N_9999,N_10065);
and U10279 (N_10279,N_10081,N_9989);
nor U10280 (N_10280,N_10069,N_10133);
and U10281 (N_10281,N_10131,N_9926);
or U10282 (N_10282,N_10044,N_10113);
nand U10283 (N_10283,N_9912,N_9922);
nand U10284 (N_10284,N_10097,N_10149);
nand U10285 (N_10285,N_9965,N_10074);
nor U10286 (N_10286,N_10006,N_10114);
nand U10287 (N_10287,N_10011,N_10137);
xor U10288 (N_10288,N_9945,N_10056);
and U10289 (N_10289,N_9998,N_9953);
or U10290 (N_10290,N_9983,N_10157);
nand U10291 (N_10291,N_10012,N_10158);
and U10292 (N_10292,N_10182,N_10130);
nor U10293 (N_10293,N_10084,N_10060);
nand U10294 (N_10294,N_10028,N_9946);
nor U10295 (N_10295,N_9931,N_9982);
nor U10296 (N_10296,N_10031,N_9995);
nand U10297 (N_10297,N_10007,N_10179);
xor U10298 (N_10298,N_9932,N_10073);
xnor U10299 (N_10299,N_10009,N_10059);
nand U10300 (N_10300,N_10172,N_10165);
or U10301 (N_10301,N_9937,N_10190);
nand U10302 (N_10302,N_10198,N_9986);
or U10303 (N_10303,N_10062,N_10173);
xnor U10304 (N_10304,N_10138,N_9904);
nand U10305 (N_10305,N_10102,N_9923);
or U10306 (N_10306,N_10048,N_10107);
nand U10307 (N_10307,N_10033,N_9905);
or U10308 (N_10308,N_9956,N_10195);
and U10309 (N_10309,N_9958,N_10072);
xor U10310 (N_10310,N_10058,N_9924);
or U10311 (N_10311,N_10079,N_10163);
or U10312 (N_10312,N_10120,N_9915);
or U10313 (N_10313,N_10159,N_9900);
nor U10314 (N_10314,N_9992,N_10121);
or U10315 (N_10315,N_9916,N_10178);
nand U10316 (N_10316,N_10145,N_10055);
nand U10317 (N_10317,N_10096,N_10083);
nor U10318 (N_10318,N_10003,N_10167);
and U10319 (N_10319,N_10054,N_10064);
or U10320 (N_10320,N_10177,N_9967);
nand U10321 (N_10321,N_9974,N_10126);
nor U10322 (N_10322,N_10155,N_10111);
nor U10323 (N_10323,N_10045,N_10116);
or U10324 (N_10324,N_10013,N_10001);
or U10325 (N_10325,N_10010,N_10109);
and U10326 (N_10326,N_9981,N_10039);
nand U10327 (N_10327,N_10105,N_10122);
and U10328 (N_10328,N_10098,N_10038);
nand U10329 (N_10329,N_10075,N_9973);
or U10330 (N_10330,N_10020,N_10188);
nor U10331 (N_10331,N_9919,N_10140);
xnor U10332 (N_10332,N_10027,N_10024);
and U10333 (N_10333,N_9910,N_9929);
nand U10334 (N_10334,N_10070,N_10143);
and U10335 (N_10335,N_9907,N_9959);
and U10336 (N_10336,N_10023,N_9984);
and U10337 (N_10337,N_10180,N_10076);
or U10338 (N_10338,N_10029,N_10025);
nor U10339 (N_10339,N_10196,N_10068);
nor U10340 (N_10340,N_10050,N_10018);
nand U10341 (N_10341,N_9966,N_9952);
and U10342 (N_10342,N_10164,N_10090);
and U10343 (N_10343,N_10170,N_10046);
or U10344 (N_10344,N_10147,N_10197);
nor U10345 (N_10345,N_9991,N_10192);
xor U10346 (N_10346,N_10142,N_9920);
or U10347 (N_10347,N_9928,N_10154);
xnor U10348 (N_10348,N_9978,N_10015);
nand U10349 (N_10349,N_10187,N_9902);
nand U10350 (N_10350,N_9986,N_10090);
nor U10351 (N_10351,N_10057,N_9906);
nor U10352 (N_10352,N_10012,N_9961);
and U10353 (N_10353,N_9969,N_10081);
or U10354 (N_10354,N_10147,N_9970);
and U10355 (N_10355,N_10199,N_10013);
and U10356 (N_10356,N_10125,N_10168);
nand U10357 (N_10357,N_10088,N_9949);
nor U10358 (N_10358,N_10081,N_10155);
nor U10359 (N_10359,N_10020,N_10119);
or U10360 (N_10360,N_10005,N_9990);
nand U10361 (N_10361,N_10134,N_9946);
xor U10362 (N_10362,N_10096,N_10133);
and U10363 (N_10363,N_9950,N_10059);
nor U10364 (N_10364,N_10052,N_10073);
nand U10365 (N_10365,N_10051,N_9999);
nand U10366 (N_10366,N_10173,N_10178);
nor U10367 (N_10367,N_9919,N_10127);
xnor U10368 (N_10368,N_10089,N_10039);
xnor U10369 (N_10369,N_10174,N_10079);
xor U10370 (N_10370,N_10082,N_10058);
and U10371 (N_10371,N_9993,N_10058);
and U10372 (N_10372,N_10172,N_9938);
xor U10373 (N_10373,N_9952,N_9974);
nand U10374 (N_10374,N_10065,N_9968);
nor U10375 (N_10375,N_9941,N_10091);
nor U10376 (N_10376,N_9944,N_10078);
nor U10377 (N_10377,N_9927,N_9924);
xnor U10378 (N_10378,N_10048,N_10060);
xnor U10379 (N_10379,N_10029,N_9962);
or U10380 (N_10380,N_9967,N_9949);
nor U10381 (N_10381,N_9930,N_9948);
xor U10382 (N_10382,N_10037,N_10125);
and U10383 (N_10383,N_10055,N_9968);
xor U10384 (N_10384,N_10160,N_10082);
or U10385 (N_10385,N_10100,N_9921);
or U10386 (N_10386,N_10184,N_10132);
xnor U10387 (N_10387,N_9928,N_10033);
and U10388 (N_10388,N_9904,N_9927);
and U10389 (N_10389,N_10041,N_10029);
and U10390 (N_10390,N_10061,N_10005);
xor U10391 (N_10391,N_10029,N_10050);
nor U10392 (N_10392,N_10198,N_9925);
nor U10393 (N_10393,N_10172,N_9995);
nand U10394 (N_10394,N_10162,N_9933);
xnor U10395 (N_10395,N_10114,N_9926);
xor U10396 (N_10396,N_10182,N_10096);
nand U10397 (N_10397,N_9975,N_10157);
or U10398 (N_10398,N_9940,N_10039);
nor U10399 (N_10399,N_10000,N_9999);
or U10400 (N_10400,N_10128,N_10113);
nor U10401 (N_10401,N_10146,N_10064);
nand U10402 (N_10402,N_10061,N_10181);
xnor U10403 (N_10403,N_10005,N_9995);
or U10404 (N_10404,N_9983,N_10051);
and U10405 (N_10405,N_10116,N_10118);
nor U10406 (N_10406,N_10103,N_9929);
xnor U10407 (N_10407,N_9957,N_9998);
and U10408 (N_10408,N_10065,N_9917);
and U10409 (N_10409,N_10072,N_9932);
nand U10410 (N_10410,N_9970,N_10176);
or U10411 (N_10411,N_10167,N_9963);
nand U10412 (N_10412,N_9993,N_10022);
nand U10413 (N_10413,N_9954,N_9991);
nand U10414 (N_10414,N_10044,N_10101);
or U10415 (N_10415,N_10159,N_10075);
and U10416 (N_10416,N_9946,N_10126);
or U10417 (N_10417,N_10162,N_10007);
nor U10418 (N_10418,N_9924,N_10078);
or U10419 (N_10419,N_10052,N_10017);
xor U10420 (N_10420,N_10185,N_9914);
and U10421 (N_10421,N_9991,N_9932);
or U10422 (N_10422,N_10156,N_10112);
nor U10423 (N_10423,N_10187,N_10181);
nor U10424 (N_10424,N_10036,N_10082);
xnor U10425 (N_10425,N_10195,N_10043);
nand U10426 (N_10426,N_10172,N_10054);
or U10427 (N_10427,N_9976,N_10008);
or U10428 (N_10428,N_10068,N_10052);
nand U10429 (N_10429,N_10127,N_10134);
and U10430 (N_10430,N_9948,N_10004);
and U10431 (N_10431,N_9964,N_9932);
nor U10432 (N_10432,N_10146,N_9965);
and U10433 (N_10433,N_10053,N_10085);
nand U10434 (N_10434,N_10100,N_10083);
nor U10435 (N_10435,N_9996,N_9908);
nand U10436 (N_10436,N_9977,N_9942);
xnor U10437 (N_10437,N_9931,N_9969);
xnor U10438 (N_10438,N_10133,N_10079);
xor U10439 (N_10439,N_10083,N_10054);
nand U10440 (N_10440,N_9954,N_10159);
nor U10441 (N_10441,N_10003,N_10162);
xnor U10442 (N_10442,N_10176,N_10172);
nand U10443 (N_10443,N_9914,N_10069);
xor U10444 (N_10444,N_10120,N_9918);
nand U10445 (N_10445,N_10017,N_9926);
nor U10446 (N_10446,N_10090,N_9918);
nand U10447 (N_10447,N_10176,N_10161);
or U10448 (N_10448,N_10196,N_10125);
nand U10449 (N_10449,N_9963,N_10111);
or U10450 (N_10450,N_9913,N_9964);
and U10451 (N_10451,N_10098,N_10184);
or U10452 (N_10452,N_9911,N_10095);
nor U10453 (N_10453,N_10162,N_10194);
nand U10454 (N_10454,N_10117,N_10028);
nand U10455 (N_10455,N_9931,N_10012);
nor U10456 (N_10456,N_9949,N_9992);
and U10457 (N_10457,N_10063,N_9918);
or U10458 (N_10458,N_10004,N_9934);
nor U10459 (N_10459,N_10026,N_9964);
xnor U10460 (N_10460,N_10174,N_9912);
xnor U10461 (N_10461,N_9925,N_9953);
and U10462 (N_10462,N_10117,N_10048);
nor U10463 (N_10463,N_10195,N_10017);
nor U10464 (N_10464,N_10196,N_10120);
nand U10465 (N_10465,N_10062,N_9992);
nand U10466 (N_10466,N_10034,N_9947);
and U10467 (N_10467,N_10071,N_10110);
xor U10468 (N_10468,N_10047,N_9937);
xnor U10469 (N_10469,N_10165,N_9931);
and U10470 (N_10470,N_10142,N_10060);
and U10471 (N_10471,N_10051,N_10037);
xor U10472 (N_10472,N_10103,N_10174);
nand U10473 (N_10473,N_9920,N_9961);
nand U10474 (N_10474,N_10024,N_10190);
nor U10475 (N_10475,N_10120,N_9967);
xnor U10476 (N_10476,N_9989,N_9973);
xor U10477 (N_10477,N_10055,N_9966);
xnor U10478 (N_10478,N_10008,N_9957);
nor U10479 (N_10479,N_10046,N_9967);
and U10480 (N_10480,N_10042,N_10119);
xnor U10481 (N_10481,N_10107,N_9930);
xor U10482 (N_10482,N_10088,N_10027);
nor U10483 (N_10483,N_10008,N_10040);
and U10484 (N_10484,N_10037,N_10151);
nand U10485 (N_10485,N_10191,N_10105);
or U10486 (N_10486,N_9985,N_10123);
xnor U10487 (N_10487,N_9981,N_10079);
xor U10488 (N_10488,N_9991,N_10140);
xnor U10489 (N_10489,N_9951,N_10009);
nor U10490 (N_10490,N_10178,N_10106);
nor U10491 (N_10491,N_9981,N_10104);
or U10492 (N_10492,N_9973,N_10027);
and U10493 (N_10493,N_9905,N_10132);
nand U10494 (N_10494,N_10032,N_9943);
nand U10495 (N_10495,N_10097,N_10136);
nand U10496 (N_10496,N_9997,N_10030);
and U10497 (N_10497,N_10050,N_10160);
xor U10498 (N_10498,N_9969,N_9902);
and U10499 (N_10499,N_10022,N_10041);
xnor U10500 (N_10500,N_10477,N_10384);
or U10501 (N_10501,N_10247,N_10283);
nor U10502 (N_10502,N_10498,N_10469);
nor U10503 (N_10503,N_10497,N_10290);
and U10504 (N_10504,N_10307,N_10319);
nor U10505 (N_10505,N_10474,N_10436);
xor U10506 (N_10506,N_10422,N_10246);
or U10507 (N_10507,N_10397,N_10243);
xnor U10508 (N_10508,N_10252,N_10267);
xor U10509 (N_10509,N_10266,N_10381);
nor U10510 (N_10510,N_10285,N_10295);
nand U10511 (N_10511,N_10364,N_10428);
or U10512 (N_10512,N_10265,N_10219);
and U10513 (N_10513,N_10483,N_10459);
nand U10514 (N_10514,N_10217,N_10250);
nand U10515 (N_10515,N_10216,N_10401);
xor U10516 (N_10516,N_10248,N_10276);
nor U10517 (N_10517,N_10417,N_10411);
nor U10518 (N_10518,N_10371,N_10271);
or U10519 (N_10519,N_10288,N_10305);
or U10520 (N_10520,N_10341,N_10286);
nor U10521 (N_10521,N_10398,N_10240);
and U10522 (N_10522,N_10235,N_10444);
or U10523 (N_10523,N_10351,N_10495);
and U10524 (N_10524,N_10275,N_10414);
or U10525 (N_10525,N_10209,N_10245);
nor U10526 (N_10526,N_10408,N_10470);
nor U10527 (N_10527,N_10278,N_10377);
and U10528 (N_10528,N_10499,N_10238);
or U10529 (N_10529,N_10274,N_10450);
and U10530 (N_10530,N_10204,N_10310);
xor U10531 (N_10531,N_10329,N_10405);
or U10532 (N_10532,N_10303,N_10257);
nand U10533 (N_10533,N_10325,N_10343);
and U10534 (N_10534,N_10468,N_10404);
and U10535 (N_10535,N_10440,N_10452);
xor U10536 (N_10536,N_10254,N_10447);
nand U10537 (N_10537,N_10306,N_10268);
xnor U10538 (N_10538,N_10324,N_10231);
xor U10539 (N_10539,N_10352,N_10300);
and U10540 (N_10540,N_10223,N_10369);
nand U10541 (N_10541,N_10317,N_10347);
and U10542 (N_10542,N_10476,N_10438);
and U10543 (N_10543,N_10225,N_10368);
and U10544 (N_10544,N_10349,N_10302);
nor U10545 (N_10545,N_10342,N_10393);
xor U10546 (N_10546,N_10228,N_10270);
nor U10547 (N_10547,N_10487,N_10361);
xnor U10548 (N_10548,N_10312,N_10353);
or U10549 (N_10549,N_10453,N_10413);
nor U10550 (N_10550,N_10456,N_10359);
nand U10551 (N_10551,N_10385,N_10392);
or U10552 (N_10552,N_10213,N_10493);
nor U10553 (N_10553,N_10331,N_10466);
xor U10554 (N_10554,N_10242,N_10211);
or U10555 (N_10555,N_10399,N_10451);
or U10556 (N_10556,N_10279,N_10481);
xor U10557 (N_10557,N_10313,N_10261);
nor U10558 (N_10558,N_10269,N_10472);
and U10559 (N_10559,N_10362,N_10210);
and U10560 (N_10560,N_10258,N_10222);
and U10561 (N_10561,N_10350,N_10395);
xnor U10562 (N_10562,N_10373,N_10332);
and U10563 (N_10563,N_10354,N_10215);
and U10564 (N_10564,N_10296,N_10284);
nand U10565 (N_10565,N_10454,N_10383);
or U10566 (N_10566,N_10253,N_10496);
nand U10567 (N_10567,N_10449,N_10280);
nand U10568 (N_10568,N_10461,N_10202);
nor U10569 (N_10569,N_10382,N_10433);
or U10570 (N_10570,N_10200,N_10434);
nor U10571 (N_10571,N_10425,N_10479);
nor U10572 (N_10572,N_10322,N_10244);
or U10573 (N_10573,N_10293,N_10489);
nor U10574 (N_10574,N_10338,N_10323);
nor U10575 (N_10575,N_10336,N_10214);
nand U10576 (N_10576,N_10441,N_10443);
xnor U10577 (N_10577,N_10442,N_10437);
xnor U10578 (N_10578,N_10237,N_10294);
and U10579 (N_10579,N_10301,N_10335);
xor U10580 (N_10580,N_10208,N_10423);
or U10581 (N_10581,N_10212,N_10221);
or U10582 (N_10582,N_10415,N_10389);
xor U10583 (N_10583,N_10282,N_10486);
nor U10584 (N_10584,N_10446,N_10412);
and U10585 (N_10585,N_10419,N_10345);
nand U10586 (N_10586,N_10344,N_10473);
or U10587 (N_10587,N_10363,N_10460);
and U10588 (N_10588,N_10320,N_10201);
nor U10589 (N_10589,N_10471,N_10367);
or U10590 (N_10590,N_10492,N_10339);
nand U10591 (N_10591,N_10328,N_10218);
nor U10592 (N_10592,N_10475,N_10488);
xnor U10593 (N_10593,N_10403,N_10375);
xor U10594 (N_10594,N_10220,N_10249);
xnor U10595 (N_10595,N_10448,N_10366);
xor U10596 (N_10596,N_10480,N_10239);
or U10597 (N_10597,N_10234,N_10251);
or U10598 (N_10598,N_10365,N_10467);
xor U10599 (N_10599,N_10327,N_10431);
or U10600 (N_10600,N_10314,N_10387);
xnor U10601 (N_10601,N_10462,N_10334);
nand U10602 (N_10602,N_10355,N_10407);
and U10603 (N_10603,N_10264,N_10358);
nor U10604 (N_10604,N_10277,N_10484);
and U10605 (N_10605,N_10346,N_10236);
or U10606 (N_10606,N_10402,N_10232);
and U10607 (N_10607,N_10348,N_10356);
nand U10608 (N_10608,N_10260,N_10337);
and U10609 (N_10609,N_10309,N_10439);
nand U10610 (N_10610,N_10273,N_10410);
nand U10611 (N_10611,N_10406,N_10321);
nand U10612 (N_10612,N_10435,N_10292);
nand U10613 (N_10613,N_10259,N_10330);
nor U10614 (N_10614,N_10409,N_10360);
or U10615 (N_10615,N_10207,N_10340);
or U10616 (N_10616,N_10427,N_10463);
nor U10617 (N_10617,N_10227,N_10263);
and U10618 (N_10618,N_10304,N_10465);
nand U10619 (N_10619,N_10308,N_10291);
nand U10620 (N_10620,N_10429,N_10396);
nand U10621 (N_10621,N_10316,N_10255);
or U10622 (N_10622,N_10432,N_10491);
nand U10623 (N_10623,N_10430,N_10455);
nor U10624 (N_10624,N_10230,N_10226);
and U10625 (N_10625,N_10424,N_10376);
nor U10626 (N_10626,N_10318,N_10485);
nor U10627 (N_10627,N_10394,N_10372);
or U10628 (N_10628,N_10464,N_10478);
nor U10629 (N_10629,N_10391,N_10206);
and U10630 (N_10630,N_10241,N_10357);
nor U10631 (N_10631,N_10421,N_10445);
xor U10632 (N_10632,N_10378,N_10458);
nor U10633 (N_10633,N_10379,N_10420);
and U10634 (N_10634,N_10457,N_10482);
nand U10635 (N_10635,N_10400,N_10386);
xor U10636 (N_10636,N_10203,N_10299);
nand U10637 (N_10637,N_10262,N_10494);
xor U10638 (N_10638,N_10289,N_10333);
nand U10639 (N_10639,N_10426,N_10370);
nor U10640 (N_10640,N_10380,N_10298);
nor U10641 (N_10641,N_10297,N_10256);
xnor U10642 (N_10642,N_10315,N_10311);
or U10643 (N_10643,N_10326,N_10287);
and U10644 (N_10644,N_10416,N_10281);
and U10645 (N_10645,N_10388,N_10490);
nand U10646 (N_10646,N_10272,N_10224);
xor U10647 (N_10647,N_10390,N_10418);
nor U10648 (N_10648,N_10233,N_10229);
nand U10649 (N_10649,N_10374,N_10205);
or U10650 (N_10650,N_10255,N_10306);
nand U10651 (N_10651,N_10393,N_10373);
nor U10652 (N_10652,N_10419,N_10398);
nor U10653 (N_10653,N_10414,N_10290);
nor U10654 (N_10654,N_10246,N_10200);
or U10655 (N_10655,N_10354,N_10252);
nor U10656 (N_10656,N_10335,N_10345);
nand U10657 (N_10657,N_10360,N_10435);
nand U10658 (N_10658,N_10380,N_10291);
and U10659 (N_10659,N_10280,N_10496);
nand U10660 (N_10660,N_10283,N_10285);
nand U10661 (N_10661,N_10392,N_10370);
and U10662 (N_10662,N_10303,N_10481);
nand U10663 (N_10663,N_10468,N_10497);
or U10664 (N_10664,N_10348,N_10279);
nor U10665 (N_10665,N_10267,N_10372);
xor U10666 (N_10666,N_10323,N_10215);
nor U10667 (N_10667,N_10259,N_10405);
and U10668 (N_10668,N_10407,N_10224);
nor U10669 (N_10669,N_10240,N_10360);
xnor U10670 (N_10670,N_10354,N_10206);
and U10671 (N_10671,N_10456,N_10413);
and U10672 (N_10672,N_10330,N_10280);
nand U10673 (N_10673,N_10375,N_10316);
nor U10674 (N_10674,N_10399,N_10268);
or U10675 (N_10675,N_10493,N_10498);
and U10676 (N_10676,N_10255,N_10372);
nand U10677 (N_10677,N_10306,N_10383);
or U10678 (N_10678,N_10218,N_10258);
or U10679 (N_10679,N_10265,N_10317);
nor U10680 (N_10680,N_10452,N_10380);
nand U10681 (N_10681,N_10270,N_10332);
and U10682 (N_10682,N_10416,N_10265);
nand U10683 (N_10683,N_10233,N_10223);
nor U10684 (N_10684,N_10216,N_10381);
and U10685 (N_10685,N_10296,N_10381);
xor U10686 (N_10686,N_10333,N_10215);
nor U10687 (N_10687,N_10454,N_10487);
or U10688 (N_10688,N_10362,N_10477);
or U10689 (N_10689,N_10459,N_10324);
xor U10690 (N_10690,N_10489,N_10336);
nand U10691 (N_10691,N_10421,N_10225);
xnor U10692 (N_10692,N_10254,N_10292);
nand U10693 (N_10693,N_10363,N_10421);
and U10694 (N_10694,N_10208,N_10451);
or U10695 (N_10695,N_10468,N_10484);
nand U10696 (N_10696,N_10286,N_10420);
nand U10697 (N_10697,N_10398,N_10274);
nor U10698 (N_10698,N_10371,N_10499);
nor U10699 (N_10699,N_10234,N_10231);
xnor U10700 (N_10700,N_10220,N_10400);
xor U10701 (N_10701,N_10317,N_10409);
and U10702 (N_10702,N_10480,N_10358);
nor U10703 (N_10703,N_10474,N_10486);
xor U10704 (N_10704,N_10415,N_10339);
nand U10705 (N_10705,N_10284,N_10211);
or U10706 (N_10706,N_10349,N_10213);
nand U10707 (N_10707,N_10308,N_10297);
and U10708 (N_10708,N_10438,N_10354);
xnor U10709 (N_10709,N_10481,N_10419);
xnor U10710 (N_10710,N_10474,N_10275);
nor U10711 (N_10711,N_10328,N_10478);
or U10712 (N_10712,N_10249,N_10379);
nand U10713 (N_10713,N_10445,N_10226);
and U10714 (N_10714,N_10482,N_10264);
or U10715 (N_10715,N_10399,N_10470);
and U10716 (N_10716,N_10334,N_10401);
nand U10717 (N_10717,N_10419,N_10450);
nor U10718 (N_10718,N_10397,N_10409);
nor U10719 (N_10719,N_10214,N_10395);
or U10720 (N_10720,N_10294,N_10477);
nand U10721 (N_10721,N_10229,N_10445);
nand U10722 (N_10722,N_10451,N_10411);
xor U10723 (N_10723,N_10495,N_10420);
nor U10724 (N_10724,N_10365,N_10217);
nor U10725 (N_10725,N_10416,N_10235);
xnor U10726 (N_10726,N_10287,N_10343);
nand U10727 (N_10727,N_10376,N_10406);
and U10728 (N_10728,N_10346,N_10452);
or U10729 (N_10729,N_10489,N_10311);
or U10730 (N_10730,N_10387,N_10287);
nor U10731 (N_10731,N_10389,N_10316);
or U10732 (N_10732,N_10419,N_10330);
nand U10733 (N_10733,N_10329,N_10386);
nor U10734 (N_10734,N_10332,N_10392);
nor U10735 (N_10735,N_10383,N_10251);
nand U10736 (N_10736,N_10346,N_10420);
or U10737 (N_10737,N_10464,N_10339);
and U10738 (N_10738,N_10296,N_10287);
nor U10739 (N_10739,N_10392,N_10447);
and U10740 (N_10740,N_10293,N_10288);
nor U10741 (N_10741,N_10333,N_10444);
nand U10742 (N_10742,N_10339,N_10397);
xnor U10743 (N_10743,N_10222,N_10421);
and U10744 (N_10744,N_10380,N_10478);
nand U10745 (N_10745,N_10401,N_10356);
nor U10746 (N_10746,N_10326,N_10302);
nor U10747 (N_10747,N_10449,N_10260);
nor U10748 (N_10748,N_10455,N_10249);
and U10749 (N_10749,N_10324,N_10427);
xnor U10750 (N_10750,N_10365,N_10279);
nand U10751 (N_10751,N_10408,N_10296);
nand U10752 (N_10752,N_10203,N_10297);
or U10753 (N_10753,N_10498,N_10366);
nand U10754 (N_10754,N_10460,N_10463);
and U10755 (N_10755,N_10266,N_10346);
nand U10756 (N_10756,N_10247,N_10323);
nand U10757 (N_10757,N_10339,N_10304);
nand U10758 (N_10758,N_10327,N_10281);
or U10759 (N_10759,N_10328,N_10398);
and U10760 (N_10760,N_10381,N_10314);
or U10761 (N_10761,N_10241,N_10393);
or U10762 (N_10762,N_10319,N_10256);
nor U10763 (N_10763,N_10316,N_10226);
nand U10764 (N_10764,N_10316,N_10435);
or U10765 (N_10765,N_10346,N_10239);
nand U10766 (N_10766,N_10315,N_10282);
and U10767 (N_10767,N_10258,N_10387);
nand U10768 (N_10768,N_10320,N_10427);
xor U10769 (N_10769,N_10218,N_10346);
nand U10770 (N_10770,N_10277,N_10486);
nor U10771 (N_10771,N_10492,N_10367);
nand U10772 (N_10772,N_10303,N_10271);
nand U10773 (N_10773,N_10406,N_10235);
nor U10774 (N_10774,N_10307,N_10365);
and U10775 (N_10775,N_10309,N_10243);
or U10776 (N_10776,N_10347,N_10291);
xor U10777 (N_10777,N_10364,N_10279);
or U10778 (N_10778,N_10228,N_10420);
nor U10779 (N_10779,N_10253,N_10344);
or U10780 (N_10780,N_10213,N_10323);
and U10781 (N_10781,N_10327,N_10334);
nor U10782 (N_10782,N_10209,N_10283);
or U10783 (N_10783,N_10211,N_10400);
or U10784 (N_10784,N_10424,N_10312);
nand U10785 (N_10785,N_10304,N_10308);
nor U10786 (N_10786,N_10330,N_10349);
or U10787 (N_10787,N_10322,N_10313);
xnor U10788 (N_10788,N_10460,N_10426);
xnor U10789 (N_10789,N_10249,N_10233);
xor U10790 (N_10790,N_10230,N_10436);
nand U10791 (N_10791,N_10274,N_10336);
nand U10792 (N_10792,N_10422,N_10374);
or U10793 (N_10793,N_10467,N_10378);
nor U10794 (N_10794,N_10413,N_10393);
nor U10795 (N_10795,N_10231,N_10219);
xnor U10796 (N_10796,N_10317,N_10414);
nand U10797 (N_10797,N_10396,N_10222);
and U10798 (N_10798,N_10344,N_10225);
or U10799 (N_10799,N_10257,N_10432);
xor U10800 (N_10800,N_10759,N_10767);
nor U10801 (N_10801,N_10603,N_10775);
and U10802 (N_10802,N_10743,N_10750);
nor U10803 (N_10803,N_10503,N_10586);
nand U10804 (N_10804,N_10629,N_10647);
xor U10805 (N_10805,N_10650,N_10730);
nand U10806 (N_10806,N_10600,N_10688);
and U10807 (N_10807,N_10536,N_10745);
nand U10808 (N_10808,N_10649,N_10614);
and U10809 (N_10809,N_10703,N_10786);
and U10810 (N_10810,N_10512,N_10712);
or U10811 (N_10811,N_10606,N_10686);
nand U10812 (N_10812,N_10726,N_10569);
xor U10813 (N_10813,N_10792,N_10694);
and U10814 (N_10814,N_10768,N_10798);
or U10815 (N_10815,N_10681,N_10526);
or U10816 (N_10816,N_10770,N_10504);
xor U10817 (N_10817,N_10696,N_10608);
xor U10818 (N_10818,N_10797,N_10630);
xnor U10819 (N_10819,N_10772,N_10642);
or U10820 (N_10820,N_10550,N_10563);
and U10821 (N_10821,N_10723,N_10584);
and U10822 (N_10822,N_10794,N_10746);
xnor U10823 (N_10823,N_10667,N_10501);
xor U10824 (N_10824,N_10622,N_10725);
or U10825 (N_10825,N_10539,N_10678);
nor U10826 (N_10826,N_10538,N_10543);
or U10827 (N_10827,N_10788,N_10721);
nand U10828 (N_10828,N_10533,N_10716);
nand U10829 (N_10829,N_10588,N_10714);
or U10830 (N_10830,N_10579,N_10732);
xor U10831 (N_10831,N_10661,N_10640);
and U10832 (N_10832,N_10796,N_10598);
xor U10833 (N_10833,N_10578,N_10632);
nor U10834 (N_10834,N_10790,N_10664);
nand U10835 (N_10835,N_10619,N_10548);
or U10836 (N_10836,N_10717,N_10523);
nand U10837 (N_10837,N_10633,N_10655);
and U10838 (N_10838,N_10735,N_10789);
xor U10839 (N_10839,N_10634,N_10668);
or U10840 (N_10840,N_10645,N_10528);
or U10841 (N_10841,N_10752,N_10657);
nor U10842 (N_10842,N_10542,N_10659);
and U10843 (N_10843,N_10627,N_10507);
xnor U10844 (N_10844,N_10757,N_10689);
or U10845 (N_10845,N_10782,N_10502);
nor U10846 (N_10846,N_10763,N_10621);
nor U10847 (N_10847,N_10566,N_10613);
or U10848 (N_10848,N_10535,N_10623);
nor U10849 (N_10849,N_10776,N_10665);
nor U10850 (N_10850,N_10524,N_10568);
nand U10851 (N_10851,N_10561,N_10595);
nor U10852 (N_10852,N_10615,N_10604);
nand U10853 (N_10853,N_10741,N_10643);
and U10854 (N_10854,N_10679,N_10652);
or U10855 (N_10855,N_10654,N_10761);
nor U10856 (N_10856,N_10670,N_10774);
nor U10857 (N_10857,N_10666,N_10559);
and U10858 (N_10858,N_10702,N_10541);
xor U10859 (N_10859,N_10585,N_10522);
nand U10860 (N_10860,N_10519,N_10571);
xor U10861 (N_10861,N_10517,N_10708);
nor U10862 (N_10862,N_10637,N_10748);
nor U10863 (N_10863,N_10506,N_10656);
or U10864 (N_10864,N_10651,N_10581);
nor U10865 (N_10865,N_10739,N_10699);
and U10866 (N_10866,N_10554,N_10513);
nor U10867 (N_10867,N_10760,N_10660);
nor U10868 (N_10868,N_10589,N_10631);
xnor U10869 (N_10869,N_10580,N_10527);
or U10870 (N_10870,N_10625,N_10572);
xnor U10871 (N_10871,N_10762,N_10676);
nor U10872 (N_10872,N_10769,N_10754);
xor U10873 (N_10873,N_10720,N_10744);
and U10874 (N_10874,N_10599,N_10715);
nand U10875 (N_10875,N_10567,N_10555);
nand U10876 (N_10876,N_10758,N_10574);
and U10877 (N_10877,N_10766,N_10673);
nand U10878 (N_10878,N_10648,N_10718);
nand U10879 (N_10879,N_10791,N_10658);
xnor U10880 (N_10880,N_10687,N_10587);
nand U10881 (N_10881,N_10693,N_10709);
nor U10882 (N_10882,N_10707,N_10755);
nand U10883 (N_10883,N_10764,N_10662);
xor U10884 (N_10884,N_10565,N_10609);
xor U10885 (N_10885,N_10537,N_10500);
and U10886 (N_10886,N_10530,N_10518);
and U10887 (N_10887,N_10675,N_10793);
and U10888 (N_10888,N_10635,N_10620);
nor U10889 (N_10889,N_10624,N_10698);
nand U10890 (N_10890,N_10781,N_10592);
and U10891 (N_10891,N_10795,N_10749);
nor U10892 (N_10892,N_10510,N_10515);
nor U10893 (N_10893,N_10784,N_10618);
nand U10894 (N_10894,N_10783,N_10582);
xnor U10895 (N_10895,N_10737,N_10765);
xor U10896 (N_10896,N_10540,N_10644);
nor U10897 (N_10897,N_10529,N_10593);
and U10898 (N_10898,N_10607,N_10697);
nor U10899 (N_10899,N_10516,N_10602);
xor U10900 (N_10900,N_10575,N_10583);
and U10901 (N_10901,N_10646,N_10753);
or U10902 (N_10902,N_10734,N_10638);
nor U10903 (N_10903,N_10549,N_10552);
xor U10904 (N_10904,N_10771,N_10610);
or U10905 (N_10905,N_10573,N_10672);
or U10906 (N_10906,N_10706,N_10773);
or U10907 (N_10907,N_10534,N_10545);
xnor U10908 (N_10908,N_10785,N_10596);
nand U10909 (N_10909,N_10557,N_10711);
and U10910 (N_10910,N_10591,N_10663);
nor U10911 (N_10911,N_10570,N_10511);
or U10912 (N_10912,N_10546,N_10677);
xor U10913 (N_10913,N_10605,N_10779);
xnor U10914 (N_10914,N_10558,N_10671);
xor U10915 (N_10915,N_10727,N_10616);
nor U10916 (N_10916,N_10551,N_10756);
xnor U10917 (N_10917,N_10617,N_10611);
xor U10918 (N_10918,N_10628,N_10682);
nor U10919 (N_10919,N_10553,N_10626);
nor U10920 (N_10920,N_10701,N_10564);
nand U10921 (N_10921,N_10612,N_10547);
xor U10922 (N_10922,N_10729,N_10713);
nor U10923 (N_10923,N_10742,N_10639);
xnor U10924 (N_10924,N_10731,N_10722);
nor U10925 (N_10925,N_10692,N_10705);
or U10926 (N_10926,N_10521,N_10780);
nor U10927 (N_10927,N_10724,N_10594);
and U10928 (N_10928,N_10560,N_10747);
nor U10929 (N_10929,N_10532,N_10799);
nand U10930 (N_10930,N_10691,N_10733);
nor U10931 (N_10931,N_10669,N_10751);
nand U10932 (N_10932,N_10778,N_10577);
or U10933 (N_10933,N_10787,N_10514);
xnor U10934 (N_10934,N_10680,N_10740);
nand U10935 (N_10935,N_10700,N_10576);
or U10936 (N_10936,N_10728,N_10508);
nor U10937 (N_10937,N_10636,N_10684);
or U10938 (N_10938,N_10520,N_10544);
or U10939 (N_10939,N_10525,N_10710);
and U10940 (N_10940,N_10509,N_10683);
or U10941 (N_10941,N_10674,N_10531);
nand U10942 (N_10942,N_10601,N_10562);
nand U10943 (N_10943,N_10695,N_10704);
and U10944 (N_10944,N_10653,N_10685);
nand U10945 (N_10945,N_10719,N_10690);
xnor U10946 (N_10946,N_10641,N_10738);
nor U10947 (N_10947,N_10590,N_10505);
and U10948 (N_10948,N_10736,N_10597);
xor U10949 (N_10949,N_10556,N_10777);
nor U10950 (N_10950,N_10700,N_10708);
nand U10951 (N_10951,N_10706,N_10782);
xnor U10952 (N_10952,N_10667,N_10623);
nor U10953 (N_10953,N_10564,N_10594);
or U10954 (N_10954,N_10568,N_10757);
and U10955 (N_10955,N_10579,N_10504);
or U10956 (N_10956,N_10745,N_10763);
or U10957 (N_10957,N_10648,N_10515);
nand U10958 (N_10958,N_10748,N_10562);
nor U10959 (N_10959,N_10571,N_10602);
nand U10960 (N_10960,N_10696,N_10648);
nor U10961 (N_10961,N_10716,N_10556);
and U10962 (N_10962,N_10559,N_10648);
xnor U10963 (N_10963,N_10602,N_10712);
and U10964 (N_10964,N_10595,N_10708);
nor U10965 (N_10965,N_10740,N_10570);
nor U10966 (N_10966,N_10649,N_10729);
xnor U10967 (N_10967,N_10767,N_10577);
nor U10968 (N_10968,N_10588,N_10612);
xnor U10969 (N_10969,N_10608,N_10569);
or U10970 (N_10970,N_10517,N_10715);
nor U10971 (N_10971,N_10596,N_10744);
nor U10972 (N_10972,N_10504,N_10578);
nor U10973 (N_10973,N_10554,N_10657);
nor U10974 (N_10974,N_10615,N_10684);
and U10975 (N_10975,N_10611,N_10758);
and U10976 (N_10976,N_10572,N_10793);
nand U10977 (N_10977,N_10778,N_10560);
nor U10978 (N_10978,N_10664,N_10588);
or U10979 (N_10979,N_10777,N_10669);
or U10980 (N_10980,N_10528,N_10629);
nand U10981 (N_10981,N_10677,N_10689);
or U10982 (N_10982,N_10739,N_10727);
xor U10983 (N_10983,N_10748,N_10696);
or U10984 (N_10984,N_10761,N_10642);
and U10985 (N_10985,N_10727,N_10719);
nor U10986 (N_10986,N_10796,N_10619);
nor U10987 (N_10987,N_10776,N_10630);
nand U10988 (N_10988,N_10613,N_10569);
xor U10989 (N_10989,N_10506,N_10732);
nor U10990 (N_10990,N_10576,N_10729);
or U10991 (N_10991,N_10608,N_10736);
nor U10992 (N_10992,N_10757,N_10733);
xnor U10993 (N_10993,N_10629,N_10500);
and U10994 (N_10994,N_10548,N_10683);
and U10995 (N_10995,N_10582,N_10717);
nor U10996 (N_10996,N_10728,N_10500);
and U10997 (N_10997,N_10796,N_10538);
or U10998 (N_10998,N_10502,N_10512);
nand U10999 (N_10999,N_10795,N_10791);
or U11000 (N_11000,N_10704,N_10675);
and U11001 (N_11001,N_10582,N_10780);
nor U11002 (N_11002,N_10602,N_10543);
and U11003 (N_11003,N_10644,N_10588);
or U11004 (N_11004,N_10720,N_10786);
or U11005 (N_11005,N_10533,N_10787);
xnor U11006 (N_11006,N_10593,N_10750);
nor U11007 (N_11007,N_10649,N_10529);
and U11008 (N_11008,N_10721,N_10728);
and U11009 (N_11009,N_10538,N_10731);
nand U11010 (N_11010,N_10680,N_10721);
or U11011 (N_11011,N_10675,N_10507);
or U11012 (N_11012,N_10768,N_10677);
xor U11013 (N_11013,N_10689,N_10769);
nand U11014 (N_11014,N_10723,N_10535);
nor U11015 (N_11015,N_10762,N_10542);
nor U11016 (N_11016,N_10573,N_10733);
or U11017 (N_11017,N_10635,N_10535);
nand U11018 (N_11018,N_10782,N_10507);
and U11019 (N_11019,N_10701,N_10550);
and U11020 (N_11020,N_10631,N_10663);
xnor U11021 (N_11021,N_10507,N_10637);
xnor U11022 (N_11022,N_10772,N_10572);
nor U11023 (N_11023,N_10757,N_10613);
or U11024 (N_11024,N_10755,N_10757);
and U11025 (N_11025,N_10771,N_10553);
and U11026 (N_11026,N_10558,N_10764);
nand U11027 (N_11027,N_10607,N_10781);
or U11028 (N_11028,N_10616,N_10724);
nor U11029 (N_11029,N_10641,N_10522);
or U11030 (N_11030,N_10679,N_10521);
nor U11031 (N_11031,N_10578,N_10677);
nor U11032 (N_11032,N_10508,N_10727);
nand U11033 (N_11033,N_10799,N_10671);
and U11034 (N_11034,N_10556,N_10582);
and U11035 (N_11035,N_10588,N_10772);
and U11036 (N_11036,N_10613,N_10671);
or U11037 (N_11037,N_10512,N_10750);
nand U11038 (N_11038,N_10670,N_10680);
xor U11039 (N_11039,N_10591,N_10609);
or U11040 (N_11040,N_10715,N_10704);
nand U11041 (N_11041,N_10673,N_10648);
xnor U11042 (N_11042,N_10783,N_10704);
and U11043 (N_11043,N_10748,N_10526);
xor U11044 (N_11044,N_10572,N_10771);
and U11045 (N_11045,N_10562,N_10651);
nor U11046 (N_11046,N_10676,N_10633);
nand U11047 (N_11047,N_10684,N_10664);
and U11048 (N_11048,N_10761,N_10611);
nor U11049 (N_11049,N_10552,N_10598);
nor U11050 (N_11050,N_10522,N_10764);
or U11051 (N_11051,N_10554,N_10705);
or U11052 (N_11052,N_10603,N_10651);
or U11053 (N_11053,N_10608,N_10713);
nand U11054 (N_11054,N_10599,N_10578);
or U11055 (N_11055,N_10614,N_10550);
nand U11056 (N_11056,N_10701,N_10768);
nor U11057 (N_11057,N_10704,N_10563);
xor U11058 (N_11058,N_10732,N_10689);
and U11059 (N_11059,N_10757,N_10790);
and U11060 (N_11060,N_10687,N_10628);
xor U11061 (N_11061,N_10625,N_10621);
nor U11062 (N_11062,N_10612,N_10700);
nor U11063 (N_11063,N_10549,N_10761);
and U11064 (N_11064,N_10673,N_10552);
nor U11065 (N_11065,N_10568,N_10603);
and U11066 (N_11066,N_10612,N_10537);
and U11067 (N_11067,N_10685,N_10584);
xor U11068 (N_11068,N_10535,N_10689);
and U11069 (N_11069,N_10722,N_10726);
and U11070 (N_11070,N_10624,N_10719);
or U11071 (N_11071,N_10701,N_10546);
nand U11072 (N_11072,N_10585,N_10634);
or U11073 (N_11073,N_10589,N_10645);
nand U11074 (N_11074,N_10556,N_10754);
nor U11075 (N_11075,N_10654,N_10754);
xnor U11076 (N_11076,N_10518,N_10652);
nand U11077 (N_11077,N_10612,N_10761);
nand U11078 (N_11078,N_10717,N_10651);
xnor U11079 (N_11079,N_10537,N_10519);
nor U11080 (N_11080,N_10553,N_10526);
nor U11081 (N_11081,N_10667,N_10578);
xnor U11082 (N_11082,N_10785,N_10548);
xor U11083 (N_11083,N_10790,N_10709);
or U11084 (N_11084,N_10629,N_10717);
or U11085 (N_11085,N_10538,N_10588);
nand U11086 (N_11086,N_10692,N_10757);
xor U11087 (N_11087,N_10581,N_10565);
nor U11088 (N_11088,N_10567,N_10608);
and U11089 (N_11089,N_10792,N_10697);
nor U11090 (N_11090,N_10796,N_10757);
nor U11091 (N_11091,N_10718,N_10553);
or U11092 (N_11092,N_10558,N_10667);
xor U11093 (N_11093,N_10643,N_10601);
nand U11094 (N_11094,N_10662,N_10538);
nor U11095 (N_11095,N_10563,N_10625);
and U11096 (N_11096,N_10579,N_10699);
or U11097 (N_11097,N_10585,N_10552);
and U11098 (N_11098,N_10524,N_10645);
and U11099 (N_11099,N_10747,N_10558);
nor U11100 (N_11100,N_10964,N_10840);
nand U11101 (N_11101,N_10875,N_11095);
or U11102 (N_11102,N_11096,N_11066);
nand U11103 (N_11103,N_10994,N_10930);
or U11104 (N_11104,N_11083,N_10958);
or U11105 (N_11105,N_10857,N_11032);
xnor U11106 (N_11106,N_10814,N_10916);
nor U11107 (N_11107,N_11000,N_10886);
nand U11108 (N_11108,N_10982,N_11076);
nand U11109 (N_11109,N_10981,N_10949);
nand U11110 (N_11110,N_10844,N_10929);
nor U11111 (N_11111,N_10895,N_10806);
nor U11112 (N_11112,N_10934,N_10810);
nor U11113 (N_11113,N_11084,N_10990);
nand U11114 (N_11114,N_11019,N_11021);
xnor U11115 (N_11115,N_11028,N_11049);
and U11116 (N_11116,N_11082,N_10816);
or U11117 (N_11117,N_10802,N_10885);
nor U11118 (N_11118,N_11048,N_10980);
and U11119 (N_11119,N_10880,N_11051);
nor U11120 (N_11120,N_11094,N_10950);
nor U11121 (N_11121,N_11090,N_11069);
or U11122 (N_11122,N_10925,N_10825);
or U11123 (N_11123,N_11073,N_10951);
and U11124 (N_11124,N_11039,N_10853);
and U11125 (N_11125,N_10942,N_11018);
or U11126 (N_11126,N_11006,N_10968);
and U11127 (N_11127,N_11068,N_11097);
nor U11128 (N_11128,N_10901,N_10907);
xnor U11129 (N_11129,N_11031,N_10993);
nor U11130 (N_11130,N_10939,N_10888);
xor U11131 (N_11131,N_10996,N_11022);
and U11132 (N_11132,N_10971,N_10881);
or U11133 (N_11133,N_10931,N_11026);
nor U11134 (N_11134,N_10910,N_10887);
nand U11135 (N_11135,N_10804,N_10893);
xnor U11136 (N_11136,N_10920,N_11091);
xnor U11137 (N_11137,N_10860,N_11078);
xor U11138 (N_11138,N_10803,N_10998);
and U11139 (N_11139,N_10969,N_11012);
or U11140 (N_11140,N_11043,N_10827);
or U11141 (N_11141,N_10850,N_10923);
nor U11142 (N_11142,N_10876,N_11017);
nand U11143 (N_11143,N_10936,N_11002);
or U11144 (N_11144,N_11054,N_10935);
nand U11145 (N_11145,N_10890,N_10984);
nor U11146 (N_11146,N_10823,N_10926);
nand U11147 (N_11147,N_10903,N_10955);
nand U11148 (N_11148,N_10906,N_10927);
nand U11149 (N_11149,N_10952,N_11020);
xor U11150 (N_11150,N_11070,N_10999);
nor U11151 (N_11151,N_10959,N_11099);
nor U11152 (N_11152,N_11052,N_11001);
or U11153 (N_11153,N_10828,N_11014);
xnor U11154 (N_11154,N_10983,N_10948);
nor U11155 (N_11155,N_10889,N_10855);
nor U11156 (N_11156,N_10834,N_10856);
xor U11157 (N_11157,N_10922,N_10818);
nor U11158 (N_11158,N_10902,N_11040);
nand U11159 (N_11159,N_10933,N_11065);
nand U11160 (N_11160,N_10878,N_10928);
xnor U11161 (N_11161,N_10868,N_11057);
nor U11162 (N_11162,N_10973,N_10905);
nand U11163 (N_11163,N_11058,N_10986);
or U11164 (N_11164,N_10833,N_10947);
nand U11165 (N_11165,N_11038,N_11041);
or U11166 (N_11166,N_10918,N_10943);
and U11167 (N_11167,N_10820,N_10912);
nand U11168 (N_11168,N_10869,N_10863);
or U11169 (N_11169,N_10897,N_10892);
or U11170 (N_11170,N_11081,N_11074);
nand U11171 (N_11171,N_10865,N_10894);
nand U11172 (N_11172,N_10849,N_10976);
nor U11173 (N_11173,N_10807,N_11061);
xor U11174 (N_11174,N_11004,N_10962);
or U11175 (N_11175,N_10846,N_10979);
or U11176 (N_11176,N_11029,N_10908);
and U11177 (N_11177,N_10891,N_10870);
or U11178 (N_11178,N_10956,N_11008);
and U11179 (N_11179,N_10985,N_10867);
and U11180 (N_11180,N_11015,N_10842);
nor U11181 (N_11181,N_11089,N_11071);
xnor U11182 (N_11182,N_10841,N_10917);
or U11183 (N_11183,N_10921,N_10831);
or U11184 (N_11184,N_11013,N_10970);
xnor U11185 (N_11185,N_10861,N_10899);
xor U11186 (N_11186,N_10837,N_10997);
nor U11187 (N_11187,N_11007,N_10848);
xor U11188 (N_11188,N_10961,N_11093);
nor U11189 (N_11189,N_10859,N_10932);
and U11190 (N_11190,N_11010,N_11036);
or U11191 (N_11191,N_11085,N_11053);
or U11192 (N_11192,N_10957,N_10896);
xnor U11193 (N_11193,N_10966,N_10826);
xor U11194 (N_11194,N_10954,N_11087);
nor U11195 (N_11195,N_10974,N_10824);
xnor U11196 (N_11196,N_11045,N_10967);
and U11197 (N_11197,N_10978,N_10862);
nand U11198 (N_11198,N_10829,N_11016);
nand U11199 (N_11199,N_10815,N_11034);
xnor U11200 (N_11200,N_11044,N_10904);
nand U11201 (N_11201,N_11072,N_10911);
or U11202 (N_11202,N_10822,N_10805);
or U11203 (N_11203,N_10882,N_10924);
and U11204 (N_11204,N_10900,N_10812);
nor U11205 (N_11205,N_10858,N_11050);
xor U11206 (N_11206,N_11037,N_10879);
and U11207 (N_11207,N_11062,N_10987);
or U11208 (N_11208,N_10909,N_10965);
nor U11209 (N_11209,N_10946,N_11060);
or U11210 (N_11210,N_11025,N_11088);
and U11211 (N_11211,N_10937,N_10864);
or U11212 (N_11212,N_10851,N_11011);
nor U11213 (N_11213,N_10836,N_10877);
nand U11214 (N_11214,N_10898,N_11009);
xor U11215 (N_11215,N_10972,N_10871);
xnor U11216 (N_11216,N_11024,N_10873);
xnor U11217 (N_11217,N_10832,N_11059);
nor U11218 (N_11218,N_11063,N_10817);
nand U11219 (N_11219,N_10975,N_10913);
nor U11220 (N_11220,N_10977,N_11005);
nor U11221 (N_11221,N_11098,N_11067);
nand U11222 (N_11222,N_10801,N_10830);
and U11223 (N_11223,N_10800,N_10960);
or U11224 (N_11224,N_11047,N_10847);
or U11225 (N_11225,N_10835,N_10839);
and U11226 (N_11226,N_10953,N_10838);
xor U11227 (N_11227,N_11055,N_10988);
xnor U11228 (N_11228,N_10845,N_11027);
nor U11229 (N_11229,N_10872,N_10914);
or U11230 (N_11230,N_11064,N_11023);
and U11231 (N_11231,N_10940,N_10944);
xnor U11232 (N_11232,N_11075,N_10919);
nor U11233 (N_11233,N_11042,N_10915);
xor U11234 (N_11234,N_11080,N_10963);
xor U11235 (N_11235,N_11046,N_10813);
and U11236 (N_11236,N_10992,N_11035);
xnor U11237 (N_11237,N_10938,N_10874);
and U11238 (N_11238,N_10821,N_10854);
nor U11239 (N_11239,N_10883,N_11003);
nand U11240 (N_11240,N_10843,N_10808);
nand U11241 (N_11241,N_10866,N_10945);
nor U11242 (N_11242,N_11092,N_10995);
nand U11243 (N_11243,N_11056,N_10811);
xnor U11244 (N_11244,N_10819,N_11077);
xnor U11245 (N_11245,N_10852,N_10941);
xnor U11246 (N_11246,N_11086,N_10884);
or U11247 (N_11247,N_10809,N_11033);
xor U11248 (N_11248,N_11079,N_10991);
nand U11249 (N_11249,N_10989,N_11030);
or U11250 (N_11250,N_11099,N_10910);
nor U11251 (N_11251,N_10895,N_10907);
or U11252 (N_11252,N_11071,N_10975);
nand U11253 (N_11253,N_10901,N_11062);
nand U11254 (N_11254,N_11043,N_10883);
nor U11255 (N_11255,N_10907,N_10854);
xnor U11256 (N_11256,N_10941,N_10913);
or U11257 (N_11257,N_10869,N_10995);
or U11258 (N_11258,N_10867,N_10955);
nand U11259 (N_11259,N_10856,N_10995);
xnor U11260 (N_11260,N_11067,N_11083);
or U11261 (N_11261,N_11012,N_11065);
and U11262 (N_11262,N_10950,N_10824);
xor U11263 (N_11263,N_10848,N_11042);
and U11264 (N_11264,N_11056,N_11047);
nand U11265 (N_11265,N_11014,N_10900);
nor U11266 (N_11266,N_10882,N_11009);
xnor U11267 (N_11267,N_10959,N_10826);
xnor U11268 (N_11268,N_11089,N_10998);
xor U11269 (N_11269,N_11023,N_11069);
nor U11270 (N_11270,N_10933,N_11031);
nor U11271 (N_11271,N_11035,N_10926);
xor U11272 (N_11272,N_10904,N_10831);
nand U11273 (N_11273,N_10867,N_11099);
or U11274 (N_11274,N_11078,N_11016);
nor U11275 (N_11275,N_10910,N_10855);
xnor U11276 (N_11276,N_10877,N_10892);
xnor U11277 (N_11277,N_10977,N_11019);
and U11278 (N_11278,N_11008,N_11058);
or U11279 (N_11279,N_10831,N_10987);
nor U11280 (N_11280,N_10908,N_10900);
nand U11281 (N_11281,N_10868,N_11083);
nor U11282 (N_11282,N_11018,N_11041);
nor U11283 (N_11283,N_10871,N_10939);
or U11284 (N_11284,N_10913,N_10919);
nand U11285 (N_11285,N_10968,N_10817);
nor U11286 (N_11286,N_10863,N_11057);
nor U11287 (N_11287,N_10979,N_10901);
and U11288 (N_11288,N_10973,N_10970);
nor U11289 (N_11289,N_10949,N_10888);
xnor U11290 (N_11290,N_10953,N_11058);
xor U11291 (N_11291,N_11027,N_10894);
nand U11292 (N_11292,N_11078,N_10844);
and U11293 (N_11293,N_10935,N_11079);
nand U11294 (N_11294,N_11034,N_10875);
or U11295 (N_11295,N_10980,N_11092);
and U11296 (N_11296,N_10984,N_10973);
xor U11297 (N_11297,N_10892,N_10960);
nand U11298 (N_11298,N_10818,N_10909);
nor U11299 (N_11299,N_11023,N_11006);
and U11300 (N_11300,N_11068,N_11007);
or U11301 (N_11301,N_11080,N_10911);
or U11302 (N_11302,N_10876,N_10849);
and U11303 (N_11303,N_10899,N_11001);
or U11304 (N_11304,N_10956,N_10905);
nor U11305 (N_11305,N_11085,N_10867);
or U11306 (N_11306,N_10897,N_11073);
nand U11307 (N_11307,N_10862,N_11070);
and U11308 (N_11308,N_11040,N_10866);
nor U11309 (N_11309,N_10888,N_10964);
xor U11310 (N_11310,N_10946,N_11002);
and U11311 (N_11311,N_10908,N_10904);
nor U11312 (N_11312,N_10812,N_10999);
and U11313 (N_11313,N_10832,N_11054);
or U11314 (N_11314,N_10951,N_10906);
and U11315 (N_11315,N_10886,N_10836);
nand U11316 (N_11316,N_10904,N_10982);
or U11317 (N_11317,N_10936,N_11090);
nor U11318 (N_11318,N_10880,N_11067);
or U11319 (N_11319,N_11097,N_10849);
xor U11320 (N_11320,N_10877,N_10852);
xnor U11321 (N_11321,N_10886,N_10895);
nor U11322 (N_11322,N_11075,N_11096);
or U11323 (N_11323,N_10911,N_11088);
nand U11324 (N_11324,N_10897,N_10990);
xor U11325 (N_11325,N_11087,N_11098);
and U11326 (N_11326,N_11001,N_10875);
and U11327 (N_11327,N_11094,N_10903);
and U11328 (N_11328,N_10859,N_11023);
xnor U11329 (N_11329,N_11066,N_11055);
nand U11330 (N_11330,N_10952,N_10803);
nand U11331 (N_11331,N_11031,N_11044);
xor U11332 (N_11332,N_11083,N_10959);
and U11333 (N_11333,N_10850,N_10984);
nand U11334 (N_11334,N_10916,N_11095);
xor U11335 (N_11335,N_11037,N_10998);
and U11336 (N_11336,N_11033,N_10997);
and U11337 (N_11337,N_10829,N_10968);
or U11338 (N_11338,N_10990,N_10911);
or U11339 (N_11339,N_11050,N_11067);
nand U11340 (N_11340,N_10953,N_11019);
xnor U11341 (N_11341,N_11056,N_11019);
xor U11342 (N_11342,N_11036,N_11098);
nor U11343 (N_11343,N_11061,N_10838);
nor U11344 (N_11344,N_10909,N_11027);
nand U11345 (N_11345,N_11071,N_10804);
nand U11346 (N_11346,N_11060,N_10812);
nand U11347 (N_11347,N_11090,N_10851);
xor U11348 (N_11348,N_11074,N_11041);
or U11349 (N_11349,N_10951,N_10853);
xnor U11350 (N_11350,N_11025,N_10876);
nor U11351 (N_11351,N_10828,N_10983);
xnor U11352 (N_11352,N_11019,N_10963);
and U11353 (N_11353,N_10914,N_10984);
nand U11354 (N_11354,N_10801,N_11069);
xnor U11355 (N_11355,N_10965,N_10912);
xor U11356 (N_11356,N_10801,N_11080);
nand U11357 (N_11357,N_10914,N_10885);
or U11358 (N_11358,N_10976,N_10853);
nor U11359 (N_11359,N_10825,N_11046);
and U11360 (N_11360,N_11053,N_10998);
nor U11361 (N_11361,N_10977,N_11080);
nor U11362 (N_11362,N_11010,N_11011);
nand U11363 (N_11363,N_11060,N_10976);
or U11364 (N_11364,N_10881,N_11049);
and U11365 (N_11365,N_11077,N_10956);
or U11366 (N_11366,N_10835,N_10862);
xnor U11367 (N_11367,N_10985,N_11086);
nor U11368 (N_11368,N_10966,N_11067);
or U11369 (N_11369,N_10800,N_10828);
nand U11370 (N_11370,N_10852,N_11009);
nor U11371 (N_11371,N_11044,N_11026);
xor U11372 (N_11372,N_10903,N_11001);
nor U11373 (N_11373,N_11060,N_10965);
nor U11374 (N_11374,N_10846,N_11049);
xnor U11375 (N_11375,N_11065,N_10804);
xnor U11376 (N_11376,N_10862,N_10914);
or U11377 (N_11377,N_10836,N_10942);
nand U11378 (N_11378,N_10939,N_10912);
xor U11379 (N_11379,N_10955,N_10901);
xor U11380 (N_11380,N_10940,N_11013);
nor U11381 (N_11381,N_11055,N_10965);
or U11382 (N_11382,N_11086,N_11070);
xnor U11383 (N_11383,N_11031,N_11026);
nor U11384 (N_11384,N_10824,N_10886);
or U11385 (N_11385,N_10809,N_10827);
nand U11386 (N_11386,N_10944,N_11010);
nor U11387 (N_11387,N_11001,N_10811);
xor U11388 (N_11388,N_11065,N_11070);
nand U11389 (N_11389,N_10996,N_11031);
nor U11390 (N_11390,N_10991,N_11020);
xnor U11391 (N_11391,N_10966,N_10866);
or U11392 (N_11392,N_11004,N_10939);
and U11393 (N_11393,N_10847,N_10969);
and U11394 (N_11394,N_10933,N_11091);
and U11395 (N_11395,N_11087,N_11071);
and U11396 (N_11396,N_10931,N_10871);
nor U11397 (N_11397,N_11091,N_11036);
or U11398 (N_11398,N_10981,N_10897);
xnor U11399 (N_11399,N_11079,N_11084);
xor U11400 (N_11400,N_11241,N_11251);
xnor U11401 (N_11401,N_11105,N_11178);
and U11402 (N_11402,N_11231,N_11235);
nand U11403 (N_11403,N_11173,N_11308);
nand U11404 (N_11404,N_11379,N_11287);
and U11405 (N_11405,N_11152,N_11243);
nand U11406 (N_11406,N_11238,N_11326);
and U11407 (N_11407,N_11355,N_11188);
or U11408 (N_11408,N_11371,N_11330);
or U11409 (N_11409,N_11316,N_11224);
and U11410 (N_11410,N_11199,N_11254);
or U11411 (N_11411,N_11212,N_11121);
xnor U11412 (N_11412,N_11168,N_11358);
or U11413 (N_11413,N_11365,N_11205);
or U11414 (N_11414,N_11177,N_11234);
nor U11415 (N_11415,N_11338,N_11163);
and U11416 (N_11416,N_11342,N_11386);
and U11417 (N_11417,N_11298,N_11372);
xor U11418 (N_11418,N_11219,N_11380);
or U11419 (N_11419,N_11128,N_11108);
or U11420 (N_11420,N_11391,N_11135);
or U11421 (N_11421,N_11174,N_11248);
nand U11422 (N_11422,N_11214,N_11293);
nand U11423 (N_11423,N_11154,N_11189);
nor U11424 (N_11424,N_11116,N_11215);
nand U11425 (N_11425,N_11156,N_11290);
nor U11426 (N_11426,N_11385,N_11132);
nand U11427 (N_11427,N_11155,N_11267);
nor U11428 (N_11428,N_11321,N_11252);
nand U11429 (N_11429,N_11120,N_11382);
xor U11430 (N_11430,N_11111,N_11150);
or U11431 (N_11431,N_11305,N_11276);
xor U11432 (N_11432,N_11323,N_11302);
xor U11433 (N_11433,N_11273,N_11172);
nor U11434 (N_11434,N_11149,N_11226);
or U11435 (N_11435,N_11364,N_11137);
or U11436 (N_11436,N_11280,N_11192);
nor U11437 (N_11437,N_11158,N_11312);
xnor U11438 (N_11438,N_11117,N_11347);
nand U11439 (N_11439,N_11229,N_11264);
xnor U11440 (N_11440,N_11327,N_11161);
and U11441 (N_11441,N_11249,N_11307);
nand U11442 (N_11442,N_11381,N_11239);
xnor U11443 (N_11443,N_11141,N_11360);
nand U11444 (N_11444,N_11310,N_11339);
and U11445 (N_11445,N_11233,N_11340);
nand U11446 (N_11446,N_11196,N_11201);
xor U11447 (N_11447,N_11294,N_11395);
or U11448 (N_11448,N_11329,N_11289);
xnor U11449 (N_11449,N_11257,N_11160);
nor U11450 (N_11450,N_11216,N_11170);
nand U11451 (N_11451,N_11328,N_11232);
nor U11452 (N_11452,N_11245,N_11122);
nor U11453 (N_11453,N_11143,N_11180);
xor U11454 (N_11454,N_11221,N_11222);
and U11455 (N_11455,N_11181,N_11322);
xor U11456 (N_11456,N_11203,N_11344);
and U11457 (N_11457,N_11228,N_11106);
xor U11458 (N_11458,N_11225,N_11124);
and U11459 (N_11459,N_11230,N_11333);
nor U11460 (N_11460,N_11145,N_11166);
nor U11461 (N_11461,N_11281,N_11348);
xnor U11462 (N_11462,N_11263,N_11259);
nand U11463 (N_11463,N_11275,N_11282);
and U11464 (N_11464,N_11204,N_11377);
nor U11465 (N_11465,N_11208,N_11262);
xnor U11466 (N_11466,N_11388,N_11139);
nand U11467 (N_11467,N_11361,N_11151);
and U11468 (N_11468,N_11311,N_11357);
xnor U11469 (N_11469,N_11304,N_11335);
nand U11470 (N_11470,N_11112,N_11260);
nor U11471 (N_11471,N_11183,N_11350);
nor U11472 (N_11472,N_11283,N_11284);
nand U11473 (N_11473,N_11153,N_11223);
and U11474 (N_11474,N_11114,N_11134);
nor U11475 (N_11475,N_11261,N_11167);
nand U11476 (N_11476,N_11270,N_11140);
xnor U11477 (N_11477,N_11297,N_11291);
or U11478 (N_11478,N_11113,N_11367);
and U11479 (N_11479,N_11250,N_11109);
nand U11480 (N_11480,N_11383,N_11397);
nor U11481 (N_11481,N_11246,N_11240);
nand U11482 (N_11482,N_11354,N_11123);
nand U11483 (N_11483,N_11220,N_11295);
xnor U11484 (N_11484,N_11198,N_11147);
xor U11485 (N_11485,N_11255,N_11186);
nor U11486 (N_11486,N_11370,N_11162);
nand U11487 (N_11487,N_11272,N_11176);
nand U11488 (N_11488,N_11387,N_11271);
xnor U11489 (N_11489,N_11258,N_11366);
and U11490 (N_11490,N_11115,N_11296);
and U11491 (N_11491,N_11236,N_11269);
or U11492 (N_11492,N_11210,N_11369);
nor U11493 (N_11493,N_11389,N_11318);
and U11494 (N_11494,N_11138,N_11392);
or U11495 (N_11495,N_11319,N_11375);
nor U11496 (N_11496,N_11268,N_11285);
and U11497 (N_11497,N_11373,N_11256);
nand U11498 (N_11498,N_11336,N_11213);
xnor U11499 (N_11499,N_11393,N_11303);
or U11500 (N_11500,N_11274,N_11202);
nor U11501 (N_11501,N_11126,N_11356);
or U11502 (N_11502,N_11104,N_11179);
nor U11503 (N_11503,N_11211,N_11345);
and U11504 (N_11504,N_11206,N_11110);
nand U11505 (N_11505,N_11107,N_11394);
or U11506 (N_11506,N_11184,N_11253);
xor U11507 (N_11507,N_11129,N_11159);
nor U11508 (N_11508,N_11374,N_11144);
nand U11509 (N_11509,N_11195,N_11207);
nor U11510 (N_11510,N_11351,N_11378);
and U11511 (N_11511,N_11127,N_11324);
nand U11512 (N_11512,N_11242,N_11314);
nand U11513 (N_11513,N_11299,N_11396);
nand U11514 (N_11514,N_11278,N_11193);
xor U11515 (N_11515,N_11157,N_11277);
nand U11516 (N_11516,N_11301,N_11306);
or U11517 (N_11517,N_11164,N_11325);
and U11518 (N_11518,N_11349,N_11266);
nor U11519 (N_11519,N_11398,N_11352);
or U11520 (N_11520,N_11288,N_11146);
or U11521 (N_11521,N_11300,N_11265);
and U11522 (N_11522,N_11368,N_11165);
xor U11523 (N_11523,N_11102,N_11399);
nor U11524 (N_11524,N_11244,N_11315);
nand U11525 (N_11525,N_11171,N_11175);
and U11526 (N_11526,N_11237,N_11341);
xnor U11527 (N_11527,N_11148,N_11182);
nor U11528 (N_11528,N_11119,N_11317);
xnor U11529 (N_11529,N_11362,N_11169);
nand U11530 (N_11530,N_11247,N_11194);
xnor U11531 (N_11531,N_11118,N_11130);
xor U11532 (N_11532,N_11332,N_11101);
or U11533 (N_11533,N_11343,N_11359);
and U11534 (N_11534,N_11133,N_11103);
nor U11535 (N_11535,N_11320,N_11218);
or U11536 (N_11536,N_11190,N_11334);
xnor U11537 (N_11537,N_11136,N_11191);
nor U11538 (N_11538,N_11185,N_11309);
nor U11539 (N_11539,N_11353,N_11384);
nor U11540 (N_11540,N_11363,N_11313);
or U11541 (N_11541,N_11331,N_11187);
nor U11542 (N_11542,N_11131,N_11100);
or U11543 (N_11543,N_11200,N_11390);
and U11544 (N_11544,N_11125,N_11279);
nor U11545 (N_11545,N_11217,N_11209);
and U11546 (N_11546,N_11227,N_11197);
xor U11547 (N_11547,N_11292,N_11337);
nor U11548 (N_11548,N_11346,N_11286);
or U11549 (N_11549,N_11376,N_11142);
or U11550 (N_11550,N_11368,N_11161);
and U11551 (N_11551,N_11386,N_11308);
nor U11552 (N_11552,N_11280,N_11187);
or U11553 (N_11553,N_11339,N_11345);
xnor U11554 (N_11554,N_11235,N_11164);
nand U11555 (N_11555,N_11363,N_11364);
nand U11556 (N_11556,N_11192,N_11235);
or U11557 (N_11557,N_11275,N_11134);
or U11558 (N_11558,N_11353,N_11263);
and U11559 (N_11559,N_11180,N_11290);
or U11560 (N_11560,N_11150,N_11284);
and U11561 (N_11561,N_11343,N_11116);
or U11562 (N_11562,N_11213,N_11299);
or U11563 (N_11563,N_11130,N_11214);
nand U11564 (N_11564,N_11265,N_11374);
and U11565 (N_11565,N_11180,N_11231);
and U11566 (N_11566,N_11337,N_11170);
or U11567 (N_11567,N_11134,N_11168);
or U11568 (N_11568,N_11259,N_11223);
and U11569 (N_11569,N_11316,N_11153);
xnor U11570 (N_11570,N_11219,N_11365);
nor U11571 (N_11571,N_11306,N_11140);
or U11572 (N_11572,N_11253,N_11327);
and U11573 (N_11573,N_11108,N_11216);
and U11574 (N_11574,N_11296,N_11362);
xor U11575 (N_11575,N_11281,N_11181);
nor U11576 (N_11576,N_11258,N_11240);
nor U11577 (N_11577,N_11271,N_11110);
and U11578 (N_11578,N_11258,N_11289);
xnor U11579 (N_11579,N_11221,N_11258);
xnor U11580 (N_11580,N_11208,N_11235);
xnor U11581 (N_11581,N_11161,N_11106);
and U11582 (N_11582,N_11151,N_11314);
nor U11583 (N_11583,N_11224,N_11277);
nor U11584 (N_11584,N_11141,N_11165);
nor U11585 (N_11585,N_11320,N_11284);
or U11586 (N_11586,N_11390,N_11155);
nand U11587 (N_11587,N_11314,N_11371);
nor U11588 (N_11588,N_11372,N_11147);
nor U11589 (N_11589,N_11103,N_11240);
xnor U11590 (N_11590,N_11312,N_11326);
xnor U11591 (N_11591,N_11157,N_11308);
nor U11592 (N_11592,N_11222,N_11232);
or U11593 (N_11593,N_11274,N_11201);
nor U11594 (N_11594,N_11392,N_11386);
nor U11595 (N_11595,N_11274,N_11352);
and U11596 (N_11596,N_11291,N_11312);
and U11597 (N_11597,N_11343,N_11104);
and U11598 (N_11598,N_11166,N_11277);
or U11599 (N_11599,N_11332,N_11201);
nand U11600 (N_11600,N_11286,N_11231);
or U11601 (N_11601,N_11321,N_11235);
nand U11602 (N_11602,N_11225,N_11325);
nand U11603 (N_11603,N_11256,N_11115);
nand U11604 (N_11604,N_11326,N_11105);
xor U11605 (N_11605,N_11354,N_11389);
nand U11606 (N_11606,N_11249,N_11124);
nand U11607 (N_11607,N_11116,N_11179);
or U11608 (N_11608,N_11199,N_11193);
or U11609 (N_11609,N_11306,N_11125);
xnor U11610 (N_11610,N_11316,N_11335);
nand U11611 (N_11611,N_11313,N_11338);
and U11612 (N_11612,N_11378,N_11216);
xnor U11613 (N_11613,N_11216,N_11305);
nor U11614 (N_11614,N_11335,N_11250);
xnor U11615 (N_11615,N_11153,N_11301);
xnor U11616 (N_11616,N_11282,N_11208);
and U11617 (N_11617,N_11132,N_11231);
xor U11618 (N_11618,N_11174,N_11205);
xnor U11619 (N_11619,N_11352,N_11299);
and U11620 (N_11620,N_11126,N_11289);
xor U11621 (N_11621,N_11281,N_11167);
and U11622 (N_11622,N_11340,N_11259);
nor U11623 (N_11623,N_11228,N_11150);
or U11624 (N_11624,N_11302,N_11289);
nand U11625 (N_11625,N_11283,N_11243);
nand U11626 (N_11626,N_11351,N_11386);
xnor U11627 (N_11627,N_11345,N_11338);
nand U11628 (N_11628,N_11307,N_11233);
xnor U11629 (N_11629,N_11169,N_11340);
nor U11630 (N_11630,N_11292,N_11162);
nand U11631 (N_11631,N_11149,N_11398);
xnor U11632 (N_11632,N_11267,N_11374);
nand U11633 (N_11633,N_11190,N_11284);
nand U11634 (N_11634,N_11202,N_11109);
or U11635 (N_11635,N_11116,N_11391);
nor U11636 (N_11636,N_11329,N_11390);
and U11637 (N_11637,N_11186,N_11383);
nor U11638 (N_11638,N_11169,N_11207);
nor U11639 (N_11639,N_11296,N_11210);
nor U11640 (N_11640,N_11308,N_11365);
and U11641 (N_11641,N_11263,N_11308);
nor U11642 (N_11642,N_11291,N_11296);
and U11643 (N_11643,N_11386,N_11353);
or U11644 (N_11644,N_11259,N_11172);
and U11645 (N_11645,N_11365,N_11210);
and U11646 (N_11646,N_11225,N_11214);
nand U11647 (N_11647,N_11371,N_11105);
or U11648 (N_11648,N_11277,N_11393);
xor U11649 (N_11649,N_11349,N_11317);
nand U11650 (N_11650,N_11144,N_11133);
or U11651 (N_11651,N_11223,N_11256);
and U11652 (N_11652,N_11137,N_11197);
nor U11653 (N_11653,N_11330,N_11127);
nor U11654 (N_11654,N_11334,N_11134);
or U11655 (N_11655,N_11305,N_11226);
xnor U11656 (N_11656,N_11251,N_11305);
and U11657 (N_11657,N_11112,N_11128);
xor U11658 (N_11658,N_11107,N_11178);
xor U11659 (N_11659,N_11161,N_11170);
xnor U11660 (N_11660,N_11376,N_11206);
and U11661 (N_11661,N_11255,N_11247);
xor U11662 (N_11662,N_11113,N_11286);
or U11663 (N_11663,N_11200,N_11218);
nand U11664 (N_11664,N_11143,N_11164);
xor U11665 (N_11665,N_11341,N_11333);
nor U11666 (N_11666,N_11108,N_11344);
and U11667 (N_11667,N_11185,N_11231);
and U11668 (N_11668,N_11322,N_11210);
or U11669 (N_11669,N_11388,N_11258);
and U11670 (N_11670,N_11177,N_11227);
and U11671 (N_11671,N_11333,N_11231);
nand U11672 (N_11672,N_11168,N_11278);
nand U11673 (N_11673,N_11266,N_11148);
xnor U11674 (N_11674,N_11206,N_11240);
xnor U11675 (N_11675,N_11196,N_11329);
and U11676 (N_11676,N_11136,N_11347);
nand U11677 (N_11677,N_11234,N_11111);
xor U11678 (N_11678,N_11174,N_11127);
xnor U11679 (N_11679,N_11222,N_11243);
or U11680 (N_11680,N_11393,N_11306);
xnor U11681 (N_11681,N_11341,N_11163);
and U11682 (N_11682,N_11372,N_11395);
xnor U11683 (N_11683,N_11343,N_11304);
xor U11684 (N_11684,N_11332,N_11374);
nand U11685 (N_11685,N_11382,N_11236);
xor U11686 (N_11686,N_11352,N_11343);
or U11687 (N_11687,N_11380,N_11116);
and U11688 (N_11688,N_11121,N_11389);
nand U11689 (N_11689,N_11193,N_11207);
nand U11690 (N_11690,N_11387,N_11380);
or U11691 (N_11691,N_11398,N_11375);
xor U11692 (N_11692,N_11241,N_11382);
nand U11693 (N_11693,N_11190,N_11174);
xnor U11694 (N_11694,N_11299,N_11382);
xor U11695 (N_11695,N_11132,N_11144);
xnor U11696 (N_11696,N_11385,N_11397);
xor U11697 (N_11697,N_11398,N_11167);
or U11698 (N_11698,N_11299,N_11302);
and U11699 (N_11699,N_11356,N_11138);
or U11700 (N_11700,N_11428,N_11489);
xor U11701 (N_11701,N_11622,N_11585);
nor U11702 (N_11702,N_11564,N_11560);
nor U11703 (N_11703,N_11532,N_11644);
xor U11704 (N_11704,N_11597,N_11422);
nor U11705 (N_11705,N_11522,N_11575);
and U11706 (N_11706,N_11627,N_11660);
and U11707 (N_11707,N_11623,N_11494);
or U11708 (N_11708,N_11565,N_11440);
or U11709 (N_11709,N_11536,N_11482);
or U11710 (N_11710,N_11443,N_11436);
xnor U11711 (N_11711,N_11453,N_11520);
nand U11712 (N_11712,N_11439,N_11652);
nor U11713 (N_11713,N_11444,N_11679);
and U11714 (N_11714,N_11691,N_11461);
nor U11715 (N_11715,N_11550,N_11603);
nand U11716 (N_11716,N_11562,N_11406);
xnor U11717 (N_11717,N_11629,N_11570);
nor U11718 (N_11718,N_11492,N_11561);
xor U11719 (N_11719,N_11526,N_11613);
and U11720 (N_11720,N_11531,N_11563);
nor U11721 (N_11721,N_11466,N_11689);
nand U11722 (N_11722,N_11432,N_11499);
nand U11723 (N_11723,N_11574,N_11437);
nand U11724 (N_11724,N_11468,N_11673);
xnor U11725 (N_11725,N_11586,N_11480);
nor U11726 (N_11726,N_11556,N_11577);
nand U11727 (N_11727,N_11557,N_11464);
nand U11728 (N_11728,N_11458,N_11505);
and U11729 (N_11729,N_11447,N_11533);
and U11730 (N_11730,N_11553,N_11469);
and U11731 (N_11731,N_11698,N_11488);
nor U11732 (N_11732,N_11455,N_11477);
and U11733 (N_11733,N_11683,N_11457);
xnor U11734 (N_11734,N_11471,N_11655);
or U11735 (N_11735,N_11415,N_11583);
xor U11736 (N_11736,N_11446,N_11528);
and U11737 (N_11737,N_11490,N_11659);
nand U11738 (N_11738,N_11452,N_11558);
xnor U11739 (N_11739,N_11518,N_11636);
nand U11740 (N_11740,N_11530,N_11584);
nand U11741 (N_11741,N_11405,N_11654);
and U11742 (N_11742,N_11669,N_11671);
xnor U11743 (N_11743,N_11545,N_11427);
nand U11744 (N_11744,N_11497,N_11667);
or U11745 (N_11745,N_11620,N_11632);
xor U11746 (N_11746,N_11605,N_11408);
nand U11747 (N_11747,N_11692,N_11596);
xor U11748 (N_11748,N_11510,N_11664);
nor U11749 (N_11749,N_11571,N_11687);
or U11750 (N_11750,N_11548,N_11551);
and U11751 (N_11751,N_11684,N_11607);
nor U11752 (N_11752,N_11529,N_11481);
xor U11753 (N_11753,N_11677,N_11699);
nand U11754 (N_11754,N_11573,N_11690);
or U11755 (N_11755,N_11676,N_11628);
and U11756 (N_11756,N_11695,N_11540);
nand U11757 (N_11757,N_11448,N_11552);
nand U11758 (N_11758,N_11618,N_11610);
or U11759 (N_11759,N_11537,N_11435);
xor U11760 (N_11760,N_11418,N_11549);
xor U11761 (N_11761,N_11624,N_11598);
xor U11762 (N_11762,N_11416,N_11486);
nand U11763 (N_11763,N_11547,N_11515);
xor U11764 (N_11764,N_11512,N_11697);
nand U11765 (N_11765,N_11639,N_11493);
nor U11766 (N_11766,N_11485,N_11483);
nand U11767 (N_11767,N_11402,N_11625);
or U11768 (N_11768,N_11590,N_11543);
xor U11769 (N_11769,N_11542,N_11535);
nor U11770 (N_11770,N_11412,N_11403);
or U11771 (N_11771,N_11686,N_11592);
nor U11772 (N_11772,N_11612,N_11582);
nor U11773 (N_11773,N_11631,N_11630);
nand U11774 (N_11774,N_11424,N_11595);
or U11775 (N_11775,N_11539,N_11475);
and U11776 (N_11776,N_11410,N_11640);
xor U11777 (N_11777,N_11524,N_11496);
and U11778 (N_11778,N_11682,N_11409);
or U11779 (N_11779,N_11445,N_11470);
and U11780 (N_11780,N_11509,N_11567);
nor U11781 (N_11781,N_11606,N_11619);
nor U11782 (N_11782,N_11538,N_11525);
nor U11783 (N_11783,N_11463,N_11450);
or U11784 (N_11784,N_11546,N_11454);
or U11785 (N_11785,N_11616,N_11656);
nand U11786 (N_11786,N_11576,N_11429);
or U11787 (N_11787,N_11611,N_11414);
nor U11788 (N_11788,N_11608,N_11465);
and U11789 (N_11789,N_11498,N_11693);
xor U11790 (N_11790,N_11642,N_11675);
and U11791 (N_11791,N_11491,N_11508);
nand U11792 (N_11792,N_11479,N_11637);
and U11793 (N_11793,N_11568,N_11609);
or U11794 (N_11794,N_11511,N_11665);
or U11795 (N_11795,N_11407,N_11413);
or U11796 (N_11796,N_11467,N_11600);
nand U11797 (N_11797,N_11670,N_11516);
xnor U11798 (N_11798,N_11650,N_11502);
and U11799 (N_11799,N_11476,N_11681);
and U11800 (N_11800,N_11604,N_11459);
or U11801 (N_11801,N_11419,N_11504);
or U11802 (N_11802,N_11517,N_11503);
and U11803 (N_11803,N_11534,N_11641);
xnor U11804 (N_11804,N_11513,N_11581);
and U11805 (N_11805,N_11694,N_11462);
nand U11806 (N_11806,N_11643,N_11417);
or U11807 (N_11807,N_11580,N_11472);
nor U11808 (N_11808,N_11400,N_11626);
or U11809 (N_11809,N_11514,N_11487);
or U11810 (N_11810,N_11651,N_11500);
nand U11811 (N_11811,N_11634,N_11589);
and U11812 (N_11812,N_11425,N_11599);
or U11813 (N_11813,N_11633,N_11451);
or U11814 (N_11814,N_11478,N_11555);
nand U11815 (N_11815,N_11460,N_11666);
and U11816 (N_11816,N_11663,N_11420);
nand U11817 (N_11817,N_11507,N_11411);
nor U11818 (N_11818,N_11614,N_11617);
xor U11819 (N_11819,N_11523,N_11685);
nor U11820 (N_11820,N_11646,N_11431);
or U11821 (N_11821,N_11519,N_11401);
nor U11822 (N_11822,N_11456,N_11569);
nor U11823 (N_11823,N_11449,N_11442);
nand U11824 (N_11824,N_11657,N_11602);
or U11825 (N_11825,N_11566,N_11678);
nor U11826 (N_11826,N_11423,N_11438);
or U11827 (N_11827,N_11615,N_11501);
nand U11828 (N_11828,N_11591,N_11527);
nand U11829 (N_11829,N_11648,N_11638);
nor U11830 (N_11830,N_11541,N_11621);
and U11831 (N_11831,N_11674,N_11601);
nand U11832 (N_11832,N_11430,N_11578);
nor U11833 (N_11833,N_11662,N_11649);
nor U11834 (N_11834,N_11645,N_11688);
and U11835 (N_11835,N_11572,N_11661);
and U11836 (N_11836,N_11404,N_11588);
nor U11837 (N_11837,N_11495,N_11658);
xnor U11838 (N_11838,N_11473,N_11594);
and U11839 (N_11839,N_11506,N_11559);
or U11840 (N_11840,N_11647,N_11579);
xnor U11841 (N_11841,N_11441,N_11421);
nor U11842 (N_11842,N_11544,N_11474);
nand U11843 (N_11843,N_11554,N_11426);
nand U11844 (N_11844,N_11635,N_11672);
nor U11845 (N_11845,N_11668,N_11680);
nor U11846 (N_11846,N_11434,N_11521);
nand U11847 (N_11847,N_11484,N_11653);
nor U11848 (N_11848,N_11587,N_11696);
and U11849 (N_11849,N_11433,N_11593);
nor U11850 (N_11850,N_11571,N_11463);
nand U11851 (N_11851,N_11490,N_11671);
nor U11852 (N_11852,N_11404,N_11473);
xnor U11853 (N_11853,N_11681,N_11660);
nor U11854 (N_11854,N_11578,N_11407);
xnor U11855 (N_11855,N_11546,N_11482);
nand U11856 (N_11856,N_11490,N_11608);
or U11857 (N_11857,N_11572,N_11588);
xor U11858 (N_11858,N_11410,N_11590);
nand U11859 (N_11859,N_11591,N_11693);
nand U11860 (N_11860,N_11630,N_11507);
and U11861 (N_11861,N_11440,N_11588);
nor U11862 (N_11862,N_11606,N_11494);
or U11863 (N_11863,N_11550,N_11572);
nand U11864 (N_11864,N_11492,N_11596);
and U11865 (N_11865,N_11450,N_11631);
nand U11866 (N_11866,N_11686,N_11602);
nand U11867 (N_11867,N_11502,N_11436);
xor U11868 (N_11868,N_11533,N_11438);
and U11869 (N_11869,N_11468,N_11609);
nand U11870 (N_11870,N_11677,N_11659);
and U11871 (N_11871,N_11630,N_11670);
xnor U11872 (N_11872,N_11699,N_11412);
xor U11873 (N_11873,N_11653,N_11448);
nand U11874 (N_11874,N_11570,N_11688);
xor U11875 (N_11875,N_11560,N_11517);
nand U11876 (N_11876,N_11662,N_11453);
nand U11877 (N_11877,N_11557,N_11630);
or U11878 (N_11878,N_11500,N_11504);
or U11879 (N_11879,N_11646,N_11589);
xnor U11880 (N_11880,N_11642,N_11667);
or U11881 (N_11881,N_11559,N_11609);
or U11882 (N_11882,N_11547,N_11478);
nor U11883 (N_11883,N_11680,N_11546);
nor U11884 (N_11884,N_11533,N_11479);
or U11885 (N_11885,N_11465,N_11555);
and U11886 (N_11886,N_11447,N_11500);
xnor U11887 (N_11887,N_11575,N_11685);
and U11888 (N_11888,N_11694,N_11442);
nor U11889 (N_11889,N_11657,N_11600);
nor U11890 (N_11890,N_11693,N_11683);
xnor U11891 (N_11891,N_11401,N_11598);
nand U11892 (N_11892,N_11541,N_11577);
xor U11893 (N_11893,N_11489,N_11613);
nor U11894 (N_11894,N_11448,N_11686);
or U11895 (N_11895,N_11629,N_11441);
xor U11896 (N_11896,N_11405,N_11604);
nor U11897 (N_11897,N_11444,N_11434);
and U11898 (N_11898,N_11461,N_11672);
nor U11899 (N_11899,N_11654,N_11455);
nor U11900 (N_11900,N_11685,N_11424);
nor U11901 (N_11901,N_11431,N_11635);
or U11902 (N_11902,N_11453,N_11517);
xor U11903 (N_11903,N_11533,N_11625);
nor U11904 (N_11904,N_11564,N_11614);
nand U11905 (N_11905,N_11453,N_11428);
nand U11906 (N_11906,N_11431,N_11475);
and U11907 (N_11907,N_11599,N_11546);
nor U11908 (N_11908,N_11612,N_11605);
nand U11909 (N_11909,N_11656,N_11443);
or U11910 (N_11910,N_11591,N_11494);
nand U11911 (N_11911,N_11459,N_11579);
or U11912 (N_11912,N_11586,N_11414);
xor U11913 (N_11913,N_11531,N_11605);
nor U11914 (N_11914,N_11670,N_11618);
xnor U11915 (N_11915,N_11504,N_11664);
and U11916 (N_11916,N_11696,N_11679);
xor U11917 (N_11917,N_11622,N_11663);
nor U11918 (N_11918,N_11610,N_11429);
and U11919 (N_11919,N_11523,N_11605);
and U11920 (N_11920,N_11432,N_11479);
nand U11921 (N_11921,N_11658,N_11510);
nor U11922 (N_11922,N_11501,N_11654);
nand U11923 (N_11923,N_11407,N_11405);
and U11924 (N_11924,N_11427,N_11579);
and U11925 (N_11925,N_11441,N_11581);
and U11926 (N_11926,N_11479,N_11696);
or U11927 (N_11927,N_11529,N_11616);
and U11928 (N_11928,N_11548,N_11479);
and U11929 (N_11929,N_11429,N_11402);
nor U11930 (N_11930,N_11468,N_11472);
or U11931 (N_11931,N_11657,N_11662);
or U11932 (N_11932,N_11534,N_11448);
and U11933 (N_11933,N_11580,N_11429);
and U11934 (N_11934,N_11643,N_11658);
and U11935 (N_11935,N_11695,N_11405);
nand U11936 (N_11936,N_11496,N_11690);
nor U11937 (N_11937,N_11454,N_11589);
or U11938 (N_11938,N_11433,N_11662);
nand U11939 (N_11939,N_11621,N_11641);
xor U11940 (N_11940,N_11555,N_11558);
nor U11941 (N_11941,N_11638,N_11510);
or U11942 (N_11942,N_11635,N_11461);
and U11943 (N_11943,N_11567,N_11696);
or U11944 (N_11944,N_11585,N_11443);
and U11945 (N_11945,N_11456,N_11521);
xnor U11946 (N_11946,N_11429,N_11459);
xor U11947 (N_11947,N_11644,N_11409);
and U11948 (N_11948,N_11489,N_11570);
xor U11949 (N_11949,N_11602,N_11608);
nand U11950 (N_11950,N_11618,N_11542);
or U11951 (N_11951,N_11405,N_11673);
or U11952 (N_11952,N_11638,N_11678);
and U11953 (N_11953,N_11631,N_11485);
nand U11954 (N_11954,N_11589,N_11411);
nor U11955 (N_11955,N_11472,N_11603);
and U11956 (N_11956,N_11540,N_11418);
nor U11957 (N_11957,N_11601,N_11530);
or U11958 (N_11958,N_11653,N_11642);
nand U11959 (N_11959,N_11686,N_11581);
or U11960 (N_11960,N_11625,N_11571);
xnor U11961 (N_11961,N_11685,N_11483);
nor U11962 (N_11962,N_11559,N_11546);
nand U11963 (N_11963,N_11590,N_11606);
and U11964 (N_11964,N_11643,N_11403);
or U11965 (N_11965,N_11595,N_11526);
and U11966 (N_11966,N_11401,N_11427);
nand U11967 (N_11967,N_11633,N_11499);
nand U11968 (N_11968,N_11671,N_11448);
xor U11969 (N_11969,N_11633,N_11604);
xnor U11970 (N_11970,N_11487,N_11628);
xnor U11971 (N_11971,N_11522,N_11648);
nand U11972 (N_11972,N_11698,N_11676);
nor U11973 (N_11973,N_11697,N_11413);
nand U11974 (N_11974,N_11604,N_11553);
nand U11975 (N_11975,N_11588,N_11487);
nand U11976 (N_11976,N_11625,N_11629);
nand U11977 (N_11977,N_11482,N_11648);
nor U11978 (N_11978,N_11667,N_11634);
nand U11979 (N_11979,N_11452,N_11643);
and U11980 (N_11980,N_11479,N_11547);
nor U11981 (N_11981,N_11645,N_11500);
and U11982 (N_11982,N_11585,N_11514);
or U11983 (N_11983,N_11682,N_11666);
nand U11984 (N_11984,N_11544,N_11631);
or U11985 (N_11985,N_11439,N_11511);
nor U11986 (N_11986,N_11585,N_11629);
nor U11987 (N_11987,N_11652,N_11615);
nor U11988 (N_11988,N_11602,N_11643);
or U11989 (N_11989,N_11566,N_11599);
and U11990 (N_11990,N_11456,N_11476);
xor U11991 (N_11991,N_11409,N_11449);
nor U11992 (N_11992,N_11567,N_11413);
nor U11993 (N_11993,N_11513,N_11659);
xor U11994 (N_11994,N_11670,N_11643);
nand U11995 (N_11995,N_11500,N_11502);
nor U11996 (N_11996,N_11430,N_11672);
nand U11997 (N_11997,N_11474,N_11497);
and U11998 (N_11998,N_11697,N_11497);
and U11999 (N_11999,N_11504,N_11650);
xor U12000 (N_12000,N_11725,N_11837);
and U12001 (N_12001,N_11959,N_11854);
or U12002 (N_12002,N_11967,N_11760);
or U12003 (N_12003,N_11727,N_11768);
xnor U12004 (N_12004,N_11731,N_11993);
xor U12005 (N_12005,N_11847,N_11905);
nand U12006 (N_12006,N_11702,N_11941);
or U12007 (N_12007,N_11998,N_11876);
or U12008 (N_12008,N_11881,N_11978);
or U12009 (N_12009,N_11816,N_11804);
nand U12010 (N_12010,N_11705,N_11851);
and U12011 (N_12011,N_11735,N_11802);
nand U12012 (N_12012,N_11829,N_11992);
nor U12013 (N_12013,N_11711,N_11806);
xnor U12014 (N_12014,N_11773,N_11758);
or U12015 (N_12015,N_11872,N_11703);
or U12016 (N_12016,N_11817,N_11868);
and U12017 (N_12017,N_11845,N_11891);
and U12018 (N_12018,N_11843,N_11771);
nand U12019 (N_12019,N_11996,N_11729);
and U12020 (N_12020,N_11910,N_11820);
nand U12021 (N_12021,N_11732,N_11908);
or U12022 (N_12022,N_11764,N_11999);
nor U12023 (N_12023,N_11841,N_11956);
xnor U12024 (N_12024,N_11792,N_11793);
nor U12025 (N_12025,N_11983,N_11809);
nor U12026 (N_12026,N_11823,N_11950);
and U12027 (N_12027,N_11995,N_11762);
xnor U12028 (N_12028,N_11885,N_11953);
and U12029 (N_12029,N_11917,N_11896);
nor U12030 (N_12030,N_11946,N_11733);
nand U12031 (N_12031,N_11719,N_11710);
or U12032 (N_12032,N_11890,N_11763);
or U12033 (N_12033,N_11898,N_11799);
or U12034 (N_12034,N_11869,N_11757);
xnor U12035 (N_12035,N_11954,N_11990);
nand U12036 (N_12036,N_11826,N_11895);
xnor U12037 (N_12037,N_11870,N_11775);
xor U12038 (N_12038,N_11740,N_11747);
and U12039 (N_12039,N_11730,N_11759);
nor U12040 (N_12040,N_11962,N_11884);
and U12041 (N_12041,N_11737,N_11780);
nand U12042 (N_12042,N_11973,N_11700);
xnor U12043 (N_12043,N_11778,N_11932);
xnor U12044 (N_12044,N_11736,N_11850);
and U12045 (N_12045,N_11926,N_11818);
nand U12046 (N_12046,N_11723,N_11975);
nor U12047 (N_12047,N_11787,N_11742);
and U12048 (N_12048,N_11933,N_11810);
nor U12049 (N_12049,N_11960,N_11788);
or U12050 (N_12050,N_11937,N_11925);
and U12051 (N_12051,N_11923,N_11899);
and U12052 (N_12052,N_11708,N_11852);
xor U12053 (N_12053,N_11716,N_11942);
xnor U12054 (N_12054,N_11879,N_11838);
or U12055 (N_12055,N_11864,N_11940);
or U12056 (N_12056,N_11738,N_11987);
nor U12057 (N_12057,N_11914,N_11722);
nand U12058 (N_12058,N_11991,N_11903);
xnor U12059 (N_12059,N_11726,N_11715);
or U12060 (N_12060,N_11979,N_11801);
nand U12061 (N_12061,N_11791,N_11704);
and U12062 (N_12062,N_11860,N_11958);
nor U12063 (N_12063,N_11880,N_11745);
xnor U12064 (N_12064,N_11794,N_11938);
and U12065 (N_12065,N_11821,N_11935);
nand U12066 (N_12066,N_11915,N_11964);
nor U12067 (N_12067,N_11728,N_11893);
or U12068 (N_12068,N_11706,N_11886);
and U12069 (N_12069,N_11774,N_11988);
and U12070 (N_12070,N_11786,N_11835);
and U12071 (N_12071,N_11779,N_11980);
nand U12072 (N_12072,N_11795,N_11798);
nor U12073 (N_12073,N_11877,N_11752);
nor U12074 (N_12074,N_11782,N_11948);
and U12075 (N_12075,N_11883,N_11741);
nor U12076 (N_12076,N_11772,N_11836);
or U12077 (N_12077,N_11986,N_11753);
and U12078 (N_12078,N_11750,N_11709);
xnor U12079 (N_12079,N_11907,N_11921);
nand U12080 (N_12080,N_11856,N_11811);
nand U12081 (N_12081,N_11784,N_11963);
xnor U12082 (N_12082,N_11800,N_11918);
or U12083 (N_12083,N_11858,N_11862);
xor U12084 (N_12084,N_11743,N_11913);
and U12085 (N_12085,N_11825,N_11930);
xnor U12086 (N_12086,N_11849,N_11828);
nor U12087 (N_12087,N_11961,N_11906);
nor U12088 (N_12088,N_11734,N_11989);
or U12089 (N_12089,N_11756,N_11892);
nand U12090 (N_12090,N_11968,N_11803);
xnor U12091 (N_12091,N_11985,N_11807);
xor U12092 (N_12092,N_11859,N_11931);
and U12093 (N_12093,N_11922,N_11984);
xnor U12094 (N_12094,N_11927,N_11754);
nor U12095 (N_12095,N_11839,N_11969);
and U12096 (N_12096,N_11974,N_11744);
xor U12097 (N_12097,N_11952,N_11904);
and U12098 (N_12098,N_11808,N_11977);
nand U12099 (N_12099,N_11769,N_11749);
nand U12100 (N_12100,N_11949,N_11902);
nand U12101 (N_12101,N_11761,N_11878);
and U12102 (N_12102,N_11765,N_11824);
nand U12103 (N_12103,N_11945,N_11944);
xnor U12104 (N_12104,N_11965,N_11713);
nor U12105 (N_12105,N_11842,N_11827);
and U12106 (N_12106,N_11901,N_11982);
nor U12107 (N_12107,N_11909,N_11831);
xnor U12108 (N_12108,N_11981,N_11746);
nand U12109 (N_12109,N_11939,N_11928);
nor U12110 (N_12110,N_11848,N_11776);
and U12111 (N_12111,N_11781,N_11897);
nor U12112 (N_12112,N_11861,N_11943);
nand U12113 (N_12113,N_11790,N_11853);
or U12114 (N_12114,N_11796,N_11815);
and U12115 (N_12115,N_11783,N_11819);
nor U12116 (N_12116,N_11936,N_11739);
and U12117 (N_12117,N_11971,N_11846);
and U12118 (N_12118,N_11844,N_11766);
nand U12119 (N_12119,N_11721,N_11707);
xor U12120 (N_12120,N_11830,N_11916);
and U12121 (N_12121,N_11822,N_11976);
nand U12122 (N_12122,N_11701,N_11966);
xor U12123 (N_12123,N_11972,N_11751);
or U12124 (N_12124,N_11957,N_11871);
and U12125 (N_12125,N_11748,N_11805);
xnor U12126 (N_12126,N_11785,N_11994);
nand U12127 (N_12127,N_11863,N_11840);
or U12128 (N_12128,N_11934,N_11789);
and U12129 (N_12129,N_11894,N_11718);
xor U12130 (N_12130,N_11873,N_11867);
or U12131 (N_12131,N_11833,N_11767);
nand U12132 (N_12132,N_11919,N_11712);
nand U12133 (N_12133,N_11924,N_11770);
and U12134 (N_12134,N_11911,N_11812);
or U12135 (N_12135,N_11813,N_11724);
nand U12136 (N_12136,N_11814,N_11797);
nand U12137 (N_12137,N_11951,N_11882);
or U12138 (N_12138,N_11929,N_11855);
or U12139 (N_12139,N_11834,N_11900);
xor U12140 (N_12140,N_11920,N_11832);
and U12141 (N_12141,N_11714,N_11889);
xnor U12142 (N_12142,N_11866,N_11997);
nand U12143 (N_12143,N_11720,N_11912);
xor U12144 (N_12144,N_11947,N_11955);
or U12145 (N_12145,N_11875,N_11887);
and U12146 (N_12146,N_11717,N_11777);
nor U12147 (N_12147,N_11755,N_11970);
and U12148 (N_12148,N_11874,N_11857);
xor U12149 (N_12149,N_11865,N_11888);
and U12150 (N_12150,N_11876,N_11874);
or U12151 (N_12151,N_11781,N_11839);
nor U12152 (N_12152,N_11750,N_11714);
xor U12153 (N_12153,N_11771,N_11759);
and U12154 (N_12154,N_11811,N_11866);
nand U12155 (N_12155,N_11857,N_11971);
nand U12156 (N_12156,N_11997,N_11796);
nand U12157 (N_12157,N_11781,N_11865);
nand U12158 (N_12158,N_11985,N_11853);
xor U12159 (N_12159,N_11800,N_11913);
nand U12160 (N_12160,N_11794,N_11992);
and U12161 (N_12161,N_11770,N_11961);
nand U12162 (N_12162,N_11943,N_11834);
xnor U12163 (N_12163,N_11821,N_11997);
nor U12164 (N_12164,N_11768,N_11911);
and U12165 (N_12165,N_11703,N_11738);
nand U12166 (N_12166,N_11924,N_11853);
and U12167 (N_12167,N_11804,N_11885);
nand U12168 (N_12168,N_11797,N_11768);
nor U12169 (N_12169,N_11706,N_11757);
and U12170 (N_12170,N_11964,N_11830);
xnor U12171 (N_12171,N_11756,N_11908);
xor U12172 (N_12172,N_11738,N_11734);
xnor U12173 (N_12173,N_11828,N_11928);
nand U12174 (N_12174,N_11787,N_11923);
nor U12175 (N_12175,N_11749,N_11783);
nand U12176 (N_12176,N_11890,N_11962);
and U12177 (N_12177,N_11704,N_11932);
nand U12178 (N_12178,N_11923,N_11833);
xnor U12179 (N_12179,N_11891,N_11820);
or U12180 (N_12180,N_11862,N_11716);
nor U12181 (N_12181,N_11918,N_11732);
nor U12182 (N_12182,N_11861,N_11957);
xor U12183 (N_12183,N_11947,N_11861);
or U12184 (N_12184,N_11781,N_11747);
or U12185 (N_12185,N_11730,N_11829);
nand U12186 (N_12186,N_11972,N_11885);
or U12187 (N_12187,N_11716,N_11877);
or U12188 (N_12188,N_11779,N_11836);
or U12189 (N_12189,N_11771,N_11906);
nor U12190 (N_12190,N_11710,N_11726);
nor U12191 (N_12191,N_11761,N_11809);
and U12192 (N_12192,N_11973,N_11966);
xor U12193 (N_12193,N_11722,N_11830);
xnor U12194 (N_12194,N_11740,N_11781);
xnor U12195 (N_12195,N_11715,N_11932);
xnor U12196 (N_12196,N_11819,N_11948);
nand U12197 (N_12197,N_11928,N_11762);
nor U12198 (N_12198,N_11909,N_11725);
nor U12199 (N_12199,N_11749,N_11868);
xor U12200 (N_12200,N_11984,N_11946);
nor U12201 (N_12201,N_11936,N_11828);
or U12202 (N_12202,N_11758,N_11989);
or U12203 (N_12203,N_11866,N_11867);
nand U12204 (N_12204,N_11809,N_11744);
nor U12205 (N_12205,N_11783,N_11856);
xnor U12206 (N_12206,N_11915,N_11835);
nor U12207 (N_12207,N_11901,N_11732);
nor U12208 (N_12208,N_11711,N_11946);
nor U12209 (N_12209,N_11715,N_11746);
nor U12210 (N_12210,N_11928,N_11783);
or U12211 (N_12211,N_11923,N_11723);
nand U12212 (N_12212,N_11904,N_11962);
nand U12213 (N_12213,N_11777,N_11967);
or U12214 (N_12214,N_11812,N_11843);
nor U12215 (N_12215,N_11771,N_11900);
or U12216 (N_12216,N_11716,N_11832);
and U12217 (N_12217,N_11858,N_11868);
nand U12218 (N_12218,N_11835,N_11975);
xnor U12219 (N_12219,N_11982,N_11967);
or U12220 (N_12220,N_11723,N_11875);
or U12221 (N_12221,N_11955,N_11940);
nand U12222 (N_12222,N_11802,N_11726);
or U12223 (N_12223,N_11883,N_11996);
and U12224 (N_12224,N_11910,N_11791);
xor U12225 (N_12225,N_11989,N_11784);
nand U12226 (N_12226,N_11957,N_11892);
and U12227 (N_12227,N_11888,N_11809);
nand U12228 (N_12228,N_11966,N_11901);
nand U12229 (N_12229,N_11756,N_11905);
xor U12230 (N_12230,N_11945,N_11989);
xor U12231 (N_12231,N_11830,N_11998);
nand U12232 (N_12232,N_11769,N_11739);
xor U12233 (N_12233,N_11848,N_11868);
and U12234 (N_12234,N_11781,N_11908);
and U12235 (N_12235,N_11784,N_11896);
nor U12236 (N_12236,N_11824,N_11774);
and U12237 (N_12237,N_11873,N_11959);
nor U12238 (N_12238,N_11964,N_11853);
and U12239 (N_12239,N_11910,N_11715);
xor U12240 (N_12240,N_11860,N_11702);
xnor U12241 (N_12241,N_11808,N_11755);
or U12242 (N_12242,N_11781,N_11861);
nor U12243 (N_12243,N_11706,N_11966);
nand U12244 (N_12244,N_11717,N_11895);
or U12245 (N_12245,N_11908,N_11989);
nor U12246 (N_12246,N_11800,N_11840);
xor U12247 (N_12247,N_11829,N_11781);
nor U12248 (N_12248,N_11758,N_11949);
and U12249 (N_12249,N_11900,N_11722);
nand U12250 (N_12250,N_11934,N_11893);
and U12251 (N_12251,N_11714,N_11906);
and U12252 (N_12252,N_11919,N_11792);
xor U12253 (N_12253,N_11938,N_11857);
and U12254 (N_12254,N_11796,N_11992);
nor U12255 (N_12255,N_11996,N_11911);
nand U12256 (N_12256,N_11788,N_11802);
nand U12257 (N_12257,N_11917,N_11907);
nor U12258 (N_12258,N_11922,N_11937);
and U12259 (N_12259,N_11776,N_11764);
or U12260 (N_12260,N_11946,N_11906);
or U12261 (N_12261,N_11981,N_11888);
nor U12262 (N_12262,N_11812,N_11759);
nand U12263 (N_12263,N_11748,N_11779);
and U12264 (N_12264,N_11943,N_11724);
nor U12265 (N_12265,N_11945,N_11743);
nand U12266 (N_12266,N_11903,N_11761);
or U12267 (N_12267,N_11959,N_11878);
xnor U12268 (N_12268,N_11892,N_11797);
and U12269 (N_12269,N_11882,N_11704);
or U12270 (N_12270,N_11705,N_11815);
nand U12271 (N_12271,N_11903,N_11889);
and U12272 (N_12272,N_11708,N_11728);
nor U12273 (N_12273,N_11705,N_11727);
xor U12274 (N_12274,N_11905,N_11924);
nor U12275 (N_12275,N_11992,N_11787);
nand U12276 (N_12276,N_11742,N_11958);
xor U12277 (N_12277,N_11986,N_11847);
nand U12278 (N_12278,N_11819,N_11865);
xnor U12279 (N_12279,N_11814,N_11756);
xor U12280 (N_12280,N_11878,N_11745);
nand U12281 (N_12281,N_11895,N_11938);
nor U12282 (N_12282,N_11703,N_11750);
and U12283 (N_12283,N_11837,N_11809);
or U12284 (N_12284,N_11796,N_11775);
xor U12285 (N_12285,N_11822,N_11872);
or U12286 (N_12286,N_11963,N_11733);
nor U12287 (N_12287,N_11794,N_11711);
or U12288 (N_12288,N_11799,N_11724);
xnor U12289 (N_12289,N_11866,N_11880);
or U12290 (N_12290,N_11730,N_11874);
nand U12291 (N_12291,N_11716,N_11807);
nand U12292 (N_12292,N_11995,N_11930);
or U12293 (N_12293,N_11830,N_11846);
nand U12294 (N_12294,N_11865,N_11780);
nand U12295 (N_12295,N_11706,N_11779);
or U12296 (N_12296,N_11975,N_11865);
or U12297 (N_12297,N_11750,N_11896);
and U12298 (N_12298,N_11796,N_11733);
nand U12299 (N_12299,N_11709,N_11930);
or U12300 (N_12300,N_12125,N_12216);
or U12301 (N_12301,N_12042,N_12090);
nand U12302 (N_12302,N_12073,N_12193);
or U12303 (N_12303,N_12143,N_12139);
and U12304 (N_12304,N_12018,N_12298);
and U12305 (N_12305,N_12126,N_12207);
nand U12306 (N_12306,N_12180,N_12050);
xnor U12307 (N_12307,N_12176,N_12147);
and U12308 (N_12308,N_12247,N_12135);
xnor U12309 (N_12309,N_12036,N_12181);
nand U12310 (N_12310,N_12007,N_12124);
and U12311 (N_12311,N_12159,N_12149);
xnor U12312 (N_12312,N_12145,N_12259);
xor U12313 (N_12313,N_12081,N_12170);
nor U12314 (N_12314,N_12102,N_12238);
nand U12315 (N_12315,N_12201,N_12106);
nand U12316 (N_12316,N_12215,N_12168);
xnor U12317 (N_12317,N_12178,N_12160);
nor U12318 (N_12318,N_12224,N_12142);
and U12319 (N_12319,N_12228,N_12058);
xor U12320 (N_12320,N_12000,N_12039);
or U12321 (N_12321,N_12233,N_12295);
nand U12322 (N_12322,N_12283,N_12164);
nor U12323 (N_12323,N_12221,N_12138);
and U12324 (N_12324,N_12251,N_12189);
or U12325 (N_12325,N_12163,N_12148);
xor U12326 (N_12326,N_12144,N_12172);
xor U12327 (N_12327,N_12061,N_12108);
or U12328 (N_12328,N_12047,N_12112);
nor U12329 (N_12329,N_12263,N_12162);
xnor U12330 (N_12330,N_12218,N_12060);
and U12331 (N_12331,N_12158,N_12296);
or U12332 (N_12332,N_12231,N_12115);
nand U12333 (N_12333,N_12219,N_12129);
and U12334 (N_12334,N_12062,N_12241);
nand U12335 (N_12335,N_12211,N_12134);
or U12336 (N_12336,N_12196,N_12026);
xor U12337 (N_12337,N_12019,N_12087);
or U12338 (N_12338,N_12071,N_12271);
and U12339 (N_12339,N_12099,N_12130);
nand U12340 (N_12340,N_12287,N_12120);
nor U12341 (N_12341,N_12273,N_12105);
and U12342 (N_12342,N_12014,N_12117);
nand U12343 (N_12343,N_12028,N_12136);
xnor U12344 (N_12344,N_12140,N_12002);
xnor U12345 (N_12345,N_12264,N_12269);
nor U12346 (N_12346,N_12070,N_12184);
and U12347 (N_12347,N_12153,N_12185);
or U12348 (N_12348,N_12030,N_12079);
or U12349 (N_12349,N_12024,N_12059);
and U12350 (N_12350,N_12278,N_12013);
xnor U12351 (N_12351,N_12232,N_12246);
and U12352 (N_12352,N_12100,N_12223);
nor U12353 (N_12353,N_12072,N_12092);
xor U12354 (N_12354,N_12281,N_12165);
nor U12355 (N_12355,N_12239,N_12171);
xor U12356 (N_12356,N_12006,N_12235);
or U12357 (N_12357,N_12230,N_12118);
and U12358 (N_12358,N_12107,N_12009);
and U12359 (N_12359,N_12226,N_12057);
and U12360 (N_12360,N_12209,N_12022);
nand U12361 (N_12361,N_12121,N_12186);
or U12362 (N_12362,N_12203,N_12222);
and U12363 (N_12363,N_12110,N_12292);
xor U12364 (N_12364,N_12015,N_12294);
xor U12365 (N_12365,N_12109,N_12175);
or U12366 (N_12366,N_12236,N_12086);
nand U12367 (N_12367,N_12151,N_12182);
nor U12368 (N_12368,N_12104,N_12097);
nand U12369 (N_12369,N_12284,N_12082);
nand U12370 (N_12370,N_12192,N_12198);
or U12371 (N_12371,N_12285,N_12008);
nor U12372 (N_12372,N_12217,N_12208);
xor U12373 (N_12373,N_12077,N_12225);
or U12374 (N_12374,N_12122,N_12080);
nand U12375 (N_12375,N_12020,N_12031);
or U12376 (N_12376,N_12242,N_12085);
nor U12377 (N_12377,N_12046,N_12156);
or U12378 (N_12378,N_12279,N_12034);
nor U12379 (N_12379,N_12248,N_12213);
and U12380 (N_12380,N_12132,N_12141);
or U12381 (N_12381,N_12265,N_12229);
xor U12382 (N_12382,N_12252,N_12037);
xor U12383 (N_12383,N_12040,N_12154);
xnor U12384 (N_12384,N_12256,N_12299);
or U12385 (N_12385,N_12114,N_12214);
nand U12386 (N_12386,N_12183,N_12029);
nor U12387 (N_12387,N_12297,N_12074);
nor U12388 (N_12388,N_12255,N_12267);
nor U12389 (N_12389,N_12258,N_12174);
nand U12390 (N_12390,N_12237,N_12257);
nand U12391 (N_12391,N_12068,N_12202);
nor U12392 (N_12392,N_12051,N_12101);
and U12393 (N_12393,N_12091,N_12274);
or U12394 (N_12394,N_12291,N_12069);
or U12395 (N_12395,N_12155,N_12244);
xor U12396 (N_12396,N_12035,N_12103);
and U12397 (N_12397,N_12290,N_12157);
nor U12398 (N_12398,N_12270,N_12190);
and U12399 (N_12399,N_12240,N_12001);
nor U12400 (N_12400,N_12063,N_12179);
nor U12401 (N_12401,N_12243,N_12277);
nor U12402 (N_12402,N_12245,N_12005);
xor U12403 (N_12403,N_12021,N_12056);
and U12404 (N_12404,N_12041,N_12261);
xor U12405 (N_12405,N_12187,N_12043);
xnor U12406 (N_12406,N_12131,N_12268);
nor U12407 (N_12407,N_12276,N_12250);
nand U12408 (N_12408,N_12054,N_12096);
and U12409 (N_12409,N_12094,N_12032);
xor U12410 (N_12410,N_12194,N_12065);
nor U12411 (N_12411,N_12012,N_12111);
or U12412 (N_12412,N_12127,N_12067);
nand U12413 (N_12413,N_12188,N_12146);
xnor U12414 (N_12414,N_12260,N_12084);
nand U12415 (N_12415,N_12275,N_12003);
nor U12416 (N_12416,N_12010,N_12289);
nor U12417 (N_12417,N_12293,N_12173);
nor U12418 (N_12418,N_12075,N_12137);
xnor U12419 (N_12419,N_12152,N_12078);
nor U12420 (N_12420,N_12044,N_12280);
xor U12421 (N_12421,N_12288,N_12016);
xnor U12422 (N_12422,N_12053,N_12045);
nor U12423 (N_12423,N_12089,N_12048);
or U12424 (N_12424,N_12197,N_12027);
nand U12425 (N_12425,N_12093,N_12166);
and U12426 (N_12426,N_12249,N_12205);
nand U12427 (N_12427,N_12023,N_12234);
and U12428 (N_12428,N_12286,N_12049);
nand U12429 (N_12429,N_12083,N_12095);
nor U12430 (N_12430,N_12038,N_12220);
nand U12431 (N_12431,N_12254,N_12191);
xnor U12432 (N_12432,N_12055,N_12064);
nand U12433 (N_12433,N_12195,N_12017);
or U12434 (N_12434,N_12011,N_12025);
nor U12435 (N_12435,N_12262,N_12253);
nand U12436 (N_12436,N_12098,N_12076);
nand U12437 (N_12437,N_12133,N_12123);
xnor U12438 (N_12438,N_12210,N_12128);
nor U12439 (N_12439,N_12004,N_12167);
nand U12440 (N_12440,N_12161,N_12033);
and U12441 (N_12441,N_12266,N_12227);
or U12442 (N_12442,N_12116,N_12204);
xor U12443 (N_12443,N_12200,N_12272);
xnor U12444 (N_12444,N_12066,N_12177);
xor U12445 (N_12445,N_12088,N_12212);
nor U12446 (N_12446,N_12169,N_12206);
and U12447 (N_12447,N_12119,N_12282);
xor U12448 (N_12448,N_12150,N_12052);
xnor U12449 (N_12449,N_12199,N_12113);
nor U12450 (N_12450,N_12135,N_12283);
nand U12451 (N_12451,N_12174,N_12170);
or U12452 (N_12452,N_12219,N_12022);
nand U12453 (N_12453,N_12223,N_12249);
xnor U12454 (N_12454,N_12087,N_12233);
xor U12455 (N_12455,N_12070,N_12026);
and U12456 (N_12456,N_12132,N_12126);
xnor U12457 (N_12457,N_12197,N_12132);
xor U12458 (N_12458,N_12138,N_12038);
and U12459 (N_12459,N_12076,N_12258);
xor U12460 (N_12460,N_12199,N_12032);
nor U12461 (N_12461,N_12176,N_12266);
nor U12462 (N_12462,N_12215,N_12273);
xor U12463 (N_12463,N_12102,N_12277);
xnor U12464 (N_12464,N_12161,N_12091);
nand U12465 (N_12465,N_12239,N_12208);
nor U12466 (N_12466,N_12127,N_12184);
nand U12467 (N_12467,N_12066,N_12256);
xnor U12468 (N_12468,N_12065,N_12062);
and U12469 (N_12469,N_12232,N_12253);
nor U12470 (N_12470,N_12143,N_12027);
xor U12471 (N_12471,N_12187,N_12128);
and U12472 (N_12472,N_12125,N_12088);
xor U12473 (N_12473,N_12224,N_12257);
nor U12474 (N_12474,N_12006,N_12156);
nand U12475 (N_12475,N_12272,N_12295);
nor U12476 (N_12476,N_12269,N_12118);
xnor U12477 (N_12477,N_12221,N_12163);
or U12478 (N_12478,N_12126,N_12046);
xor U12479 (N_12479,N_12035,N_12021);
nor U12480 (N_12480,N_12138,N_12270);
nand U12481 (N_12481,N_12192,N_12048);
xor U12482 (N_12482,N_12124,N_12246);
nand U12483 (N_12483,N_12189,N_12039);
and U12484 (N_12484,N_12252,N_12217);
and U12485 (N_12485,N_12111,N_12004);
nor U12486 (N_12486,N_12095,N_12136);
nand U12487 (N_12487,N_12183,N_12193);
nand U12488 (N_12488,N_12049,N_12235);
and U12489 (N_12489,N_12126,N_12108);
xor U12490 (N_12490,N_12077,N_12268);
nand U12491 (N_12491,N_12232,N_12211);
and U12492 (N_12492,N_12013,N_12018);
nand U12493 (N_12493,N_12105,N_12228);
xor U12494 (N_12494,N_12299,N_12072);
and U12495 (N_12495,N_12081,N_12242);
nand U12496 (N_12496,N_12100,N_12198);
nor U12497 (N_12497,N_12281,N_12206);
nand U12498 (N_12498,N_12187,N_12143);
nand U12499 (N_12499,N_12153,N_12228);
nand U12500 (N_12500,N_12047,N_12160);
and U12501 (N_12501,N_12075,N_12080);
nor U12502 (N_12502,N_12137,N_12179);
or U12503 (N_12503,N_12121,N_12125);
or U12504 (N_12504,N_12240,N_12174);
nor U12505 (N_12505,N_12183,N_12265);
and U12506 (N_12506,N_12036,N_12087);
xnor U12507 (N_12507,N_12022,N_12288);
and U12508 (N_12508,N_12075,N_12030);
nand U12509 (N_12509,N_12294,N_12211);
or U12510 (N_12510,N_12025,N_12209);
or U12511 (N_12511,N_12103,N_12016);
or U12512 (N_12512,N_12262,N_12196);
or U12513 (N_12513,N_12159,N_12225);
xor U12514 (N_12514,N_12106,N_12056);
or U12515 (N_12515,N_12076,N_12000);
or U12516 (N_12516,N_12252,N_12081);
or U12517 (N_12517,N_12003,N_12054);
xor U12518 (N_12518,N_12063,N_12142);
or U12519 (N_12519,N_12270,N_12263);
nand U12520 (N_12520,N_12213,N_12030);
or U12521 (N_12521,N_12179,N_12097);
xor U12522 (N_12522,N_12077,N_12095);
nand U12523 (N_12523,N_12237,N_12026);
and U12524 (N_12524,N_12152,N_12181);
or U12525 (N_12525,N_12090,N_12150);
nor U12526 (N_12526,N_12030,N_12056);
or U12527 (N_12527,N_12080,N_12165);
nand U12528 (N_12528,N_12247,N_12232);
and U12529 (N_12529,N_12009,N_12203);
or U12530 (N_12530,N_12028,N_12005);
xnor U12531 (N_12531,N_12288,N_12186);
or U12532 (N_12532,N_12179,N_12266);
nand U12533 (N_12533,N_12175,N_12185);
xnor U12534 (N_12534,N_12235,N_12229);
xor U12535 (N_12535,N_12009,N_12285);
or U12536 (N_12536,N_12002,N_12092);
xor U12537 (N_12537,N_12094,N_12086);
nand U12538 (N_12538,N_12239,N_12097);
nand U12539 (N_12539,N_12276,N_12182);
nand U12540 (N_12540,N_12299,N_12241);
and U12541 (N_12541,N_12227,N_12123);
nand U12542 (N_12542,N_12276,N_12037);
nor U12543 (N_12543,N_12287,N_12087);
or U12544 (N_12544,N_12299,N_12096);
nand U12545 (N_12545,N_12010,N_12093);
xor U12546 (N_12546,N_12155,N_12081);
and U12547 (N_12547,N_12297,N_12054);
nand U12548 (N_12548,N_12102,N_12000);
or U12549 (N_12549,N_12106,N_12179);
xnor U12550 (N_12550,N_12120,N_12168);
nor U12551 (N_12551,N_12020,N_12206);
and U12552 (N_12552,N_12202,N_12294);
nand U12553 (N_12553,N_12013,N_12002);
nand U12554 (N_12554,N_12037,N_12017);
xnor U12555 (N_12555,N_12010,N_12134);
nor U12556 (N_12556,N_12079,N_12208);
and U12557 (N_12557,N_12002,N_12132);
nor U12558 (N_12558,N_12008,N_12211);
xor U12559 (N_12559,N_12274,N_12264);
xnor U12560 (N_12560,N_12163,N_12268);
or U12561 (N_12561,N_12214,N_12169);
nor U12562 (N_12562,N_12092,N_12284);
nand U12563 (N_12563,N_12202,N_12044);
xor U12564 (N_12564,N_12211,N_12226);
xnor U12565 (N_12565,N_12141,N_12095);
or U12566 (N_12566,N_12247,N_12028);
nor U12567 (N_12567,N_12014,N_12281);
and U12568 (N_12568,N_12172,N_12207);
or U12569 (N_12569,N_12036,N_12295);
and U12570 (N_12570,N_12234,N_12283);
xor U12571 (N_12571,N_12263,N_12238);
or U12572 (N_12572,N_12289,N_12048);
or U12573 (N_12573,N_12237,N_12041);
nor U12574 (N_12574,N_12275,N_12132);
nor U12575 (N_12575,N_12128,N_12142);
nand U12576 (N_12576,N_12050,N_12049);
nand U12577 (N_12577,N_12091,N_12267);
and U12578 (N_12578,N_12055,N_12206);
nor U12579 (N_12579,N_12208,N_12229);
or U12580 (N_12580,N_12022,N_12057);
xnor U12581 (N_12581,N_12115,N_12182);
nor U12582 (N_12582,N_12076,N_12056);
nand U12583 (N_12583,N_12147,N_12270);
xnor U12584 (N_12584,N_12277,N_12209);
or U12585 (N_12585,N_12283,N_12203);
nor U12586 (N_12586,N_12213,N_12072);
nand U12587 (N_12587,N_12180,N_12035);
xnor U12588 (N_12588,N_12143,N_12264);
xor U12589 (N_12589,N_12176,N_12046);
or U12590 (N_12590,N_12281,N_12044);
or U12591 (N_12591,N_12069,N_12293);
or U12592 (N_12592,N_12025,N_12232);
or U12593 (N_12593,N_12140,N_12118);
and U12594 (N_12594,N_12101,N_12230);
xnor U12595 (N_12595,N_12234,N_12091);
or U12596 (N_12596,N_12293,N_12116);
and U12597 (N_12597,N_12227,N_12221);
xor U12598 (N_12598,N_12259,N_12072);
nand U12599 (N_12599,N_12171,N_12006);
nor U12600 (N_12600,N_12429,N_12326);
and U12601 (N_12601,N_12550,N_12598);
nand U12602 (N_12602,N_12522,N_12407);
nor U12603 (N_12603,N_12350,N_12483);
or U12604 (N_12604,N_12389,N_12312);
nand U12605 (N_12605,N_12333,N_12591);
nand U12606 (N_12606,N_12451,N_12322);
or U12607 (N_12607,N_12530,N_12464);
and U12608 (N_12608,N_12357,N_12549);
nor U12609 (N_12609,N_12475,N_12538);
nor U12610 (N_12610,N_12551,N_12335);
xor U12611 (N_12611,N_12452,N_12492);
nor U12612 (N_12612,N_12569,N_12554);
and U12613 (N_12613,N_12432,N_12526);
or U12614 (N_12614,N_12566,N_12568);
nand U12615 (N_12615,N_12321,N_12380);
nor U12616 (N_12616,N_12360,N_12574);
nor U12617 (N_12617,N_12556,N_12485);
nand U12618 (N_12618,N_12307,N_12457);
and U12619 (N_12619,N_12552,N_12359);
and U12620 (N_12620,N_12560,N_12570);
xnor U12621 (N_12621,N_12364,N_12511);
nand U12622 (N_12622,N_12513,N_12400);
nor U12623 (N_12623,N_12503,N_12417);
and U12624 (N_12624,N_12414,N_12355);
or U12625 (N_12625,N_12544,N_12583);
nand U12626 (N_12626,N_12430,N_12501);
xnor U12627 (N_12627,N_12301,N_12521);
nor U12628 (N_12628,N_12494,N_12339);
nor U12629 (N_12629,N_12433,N_12519);
or U12630 (N_12630,N_12361,N_12499);
nor U12631 (N_12631,N_12514,N_12518);
or U12632 (N_12632,N_12427,N_12394);
nor U12633 (N_12633,N_12349,N_12565);
nand U12634 (N_12634,N_12453,N_12356);
and U12635 (N_12635,N_12527,N_12428);
or U12636 (N_12636,N_12450,N_12564);
xnor U12637 (N_12637,N_12468,N_12311);
nand U12638 (N_12638,N_12454,N_12529);
and U12639 (N_12639,N_12398,N_12548);
nor U12640 (N_12640,N_12510,N_12336);
nand U12641 (N_12641,N_12406,N_12539);
xnor U12642 (N_12642,N_12575,N_12484);
nand U12643 (N_12643,N_12490,N_12379);
nand U12644 (N_12644,N_12441,N_12386);
nand U12645 (N_12645,N_12422,N_12334);
nand U12646 (N_12646,N_12448,N_12354);
nand U12647 (N_12647,N_12381,N_12313);
xor U12648 (N_12648,N_12592,N_12416);
and U12649 (N_12649,N_12491,N_12547);
nor U12650 (N_12650,N_12474,N_12347);
or U12651 (N_12651,N_12532,N_12588);
nand U12652 (N_12652,N_12505,N_12535);
and U12653 (N_12653,N_12515,N_12376);
xor U12654 (N_12654,N_12531,N_12303);
and U12655 (N_12655,N_12328,N_12319);
nand U12656 (N_12656,N_12533,N_12498);
or U12657 (N_12657,N_12467,N_12412);
or U12658 (N_12658,N_12344,N_12345);
nand U12659 (N_12659,N_12572,N_12542);
or U12660 (N_12660,N_12472,N_12446);
nand U12661 (N_12661,N_12504,N_12310);
nor U12662 (N_12662,N_12496,N_12488);
or U12663 (N_12663,N_12413,N_12597);
nor U12664 (N_12664,N_12593,N_12573);
nor U12665 (N_12665,N_12403,N_12351);
xnor U12666 (N_12666,N_12404,N_12383);
nand U12667 (N_12667,N_12579,N_12393);
nor U12668 (N_12668,N_12558,N_12302);
and U12669 (N_12669,N_12595,N_12445);
or U12670 (N_12670,N_12424,N_12371);
or U12671 (N_12671,N_12462,N_12368);
and U12672 (N_12672,N_12308,N_12395);
nor U12673 (N_12673,N_12426,N_12399);
xor U12674 (N_12674,N_12325,N_12392);
nand U12675 (N_12675,N_12497,N_12523);
nand U12676 (N_12676,N_12377,N_12409);
nor U12677 (N_12677,N_12461,N_12540);
and U12678 (N_12678,N_12423,N_12402);
and U12679 (N_12679,N_12337,N_12365);
and U12680 (N_12680,N_12374,N_12341);
or U12681 (N_12681,N_12500,N_12517);
or U12682 (N_12682,N_12459,N_12306);
nand U12683 (N_12683,N_12370,N_12508);
nand U12684 (N_12684,N_12358,N_12304);
nand U12685 (N_12685,N_12553,N_12495);
nor U12686 (N_12686,N_12463,N_12562);
nand U12687 (N_12687,N_12353,N_12329);
and U12688 (N_12688,N_12528,N_12323);
or U12689 (N_12689,N_12545,N_12343);
nor U12690 (N_12690,N_12408,N_12431);
nor U12691 (N_12691,N_12596,N_12330);
nor U12692 (N_12692,N_12561,N_12581);
or U12693 (N_12693,N_12520,N_12584);
and U12694 (N_12694,N_12480,N_12576);
and U12695 (N_12695,N_12541,N_12410);
and U12696 (N_12696,N_12314,N_12418);
and U12697 (N_12697,N_12362,N_12387);
nand U12698 (N_12698,N_12512,N_12477);
and U12699 (N_12699,N_12587,N_12435);
or U12700 (N_12700,N_12439,N_12324);
nor U12701 (N_12701,N_12401,N_12546);
nor U12702 (N_12702,N_12486,N_12420);
nor U12703 (N_12703,N_12411,N_12559);
xnor U12704 (N_12704,N_12440,N_12397);
xnor U12705 (N_12705,N_12525,N_12375);
nor U12706 (N_12706,N_12436,N_12524);
or U12707 (N_12707,N_12444,N_12388);
xor U12708 (N_12708,N_12434,N_12363);
xor U12709 (N_12709,N_12465,N_12366);
nor U12710 (N_12710,N_12537,N_12405);
xnor U12711 (N_12711,N_12590,N_12470);
nor U12712 (N_12712,N_12384,N_12578);
and U12713 (N_12713,N_12317,N_12469);
nand U12714 (N_12714,N_12309,N_12471);
xor U12715 (N_12715,N_12481,N_12346);
nand U12716 (N_12716,N_12352,N_12502);
or U12717 (N_12717,N_12385,N_12458);
and U12718 (N_12718,N_12478,N_12373);
or U12719 (N_12719,N_12449,N_12594);
and U12720 (N_12720,N_12442,N_12419);
xor U12721 (N_12721,N_12557,N_12367);
or U12722 (N_12722,N_12487,N_12320);
xor U12723 (N_12723,N_12331,N_12318);
and U12724 (N_12724,N_12421,N_12577);
and U12725 (N_12725,N_12555,N_12332);
and U12726 (N_12726,N_12567,N_12582);
and U12727 (N_12727,N_12447,N_12599);
or U12728 (N_12728,N_12585,N_12580);
and U12729 (N_12729,N_12390,N_12563);
and U12730 (N_12730,N_12438,N_12536);
nand U12731 (N_12731,N_12516,N_12460);
nor U12732 (N_12732,N_12479,N_12473);
xnor U12733 (N_12733,N_12571,N_12305);
and U12734 (N_12734,N_12455,N_12415);
xnor U12735 (N_12735,N_12534,N_12586);
and U12736 (N_12736,N_12382,N_12507);
nand U12737 (N_12737,N_12315,N_12327);
or U12738 (N_12738,N_12378,N_12443);
nand U12739 (N_12739,N_12340,N_12589);
or U12740 (N_12740,N_12342,N_12482);
nand U12741 (N_12741,N_12369,N_12543);
or U12742 (N_12742,N_12509,N_12437);
nor U12743 (N_12743,N_12493,N_12425);
nor U12744 (N_12744,N_12396,N_12348);
or U12745 (N_12745,N_12506,N_12489);
xnor U12746 (N_12746,N_12338,N_12316);
and U12747 (N_12747,N_12476,N_12391);
or U12748 (N_12748,N_12372,N_12300);
and U12749 (N_12749,N_12466,N_12456);
and U12750 (N_12750,N_12370,N_12464);
or U12751 (N_12751,N_12446,N_12404);
nand U12752 (N_12752,N_12587,N_12472);
or U12753 (N_12753,N_12467,N_12386);
nor U12754 (N_12754,N_12475,N_12544);
and U12755 (N_12755,N_12520,N_12425);
or U12756 (N_12756,N_12554,N_12441);
nor U12757 (N_12757,N_12366,N_12417);
or U12758 (N_12758,N_12385,N_12560);
nand U12759 (N_12759,N_12569,N_12377);
xor U12760 (N_12760,N_12596,N_12353);
or U12761 (N_12761,N_12513,N_12449);
xor U12762 (N_12762,N_12485,N_12476);
nor U12763 (N_12763,N_12387,N_12528);
nand U12764 (N_12764,N_12440,N_12349);
nor U12765 (N_12765,N_12376,N_12588);
nor U12766 (N_12766,N_12462,N_12451);
or U12767 (N_12767,N_12494,N_12303);
xnor U12768 (N_12768,N_12327,N_12418);
xnor U12769 (N_12769,N_12319,N_12335);
and U12770 (N_12770,N_12400,N_12385);
and U12771 (N_12771,N_12381,N_12427);
or U12772 (N_12772,N_12492,N_12382);
or U12773 (N_12773,N_12322,N_12427);
and U12774 (N_12774,N_12374,N_12459);
or U12775 (N_12775,N_12531,N_12445);
xor U12776 (N_12776,N_12355,N_12526);
nor U12777 (N_12777,N_12559,N_12339);
xnor U12778 (N_12778,N_12552,N_12587);
and U12779 (N_12779,N_12379,N_12429);
or U12780 (N_12780,N_12553,N_12341);
or U12781 (N_12781,N_12499,N_12381);
nand U12782 (N_12782,N_12473,N_12509);
xnor U12783 (N_12783,N_12524,N_12449);
nand U12784 (N_12784,N_12328,N_12492);
or U12785 (N_12785,N_12349,N_12524);
and U12786 (N_12786,N_12371,N_12304);
nor U12787 (N_12787,N_12439,N_12401);
nor U12788 (N_12788,N_12365,N_12343);
and U12789 (N_12789,N_12486,N_12307);
nor U12790 (N_12790,N_12581,N_12489);
and U12791 (N_12791,N_12454,N_12561);
nor U12792 (N_12792,N_12461,N_12410);
nor U12793 (N_12793,N_12363,N_12583);
and U12794 (N_12794,N_12494,N_12393);
and U12795 (N_12795,N_12354,N_12587);
or U12796 (N_12796,N_12316,N_12450);
nor U12797 (N_12797,N_12506,N_12333);
xor U12798 (N_12798,N_12526,N_12366);
xor U12799 (N_12799,N_12301,N_12527);
nand U12800 (N_12800,N_12572,N_12302);
nor U12801 (N_12801,N_12433,N_12312);
or U12802 (N_12802,N_12499,N_12320);
and U12803 (N_12803,N_12408,N_12380);
and U12804 (N_12804,N_12402,N_12384);
nor U12805 (N_12805,N_12309,N_12304);
xnor U12806 (N_12806,N_12323,N_12554);
xnor U12807 (N_12807,N_12379,N_12450);
and U12808 (N_12808,N_12527,N_12328);
nor U12809 (N_12809,N_12523,N_12467);
or U12810 (N_12810,N_12373,N_12420);
xnor U12811 (N_12811,N_12574,N_12418);
xnor U12812 (N_12812,N_12564,N_12395);
nand U12813 (N_12813,N_12592,N_12438);
xnor U12814 (N_12814,N_12506,N_12375);
xnor U12815 (N_12815,N_12544,N_12507);
nand U12816 (N_12816,N_12431,N_12580);
nand U12817 (N_12817,N_12504,N_12459);
xnor U12818 (N_12818,N_12566,N_12574);
xnor U12819 (N_12819,N_12400,N_12542);
or U12820 (N_12820,N_12535,N_12503);
or U12821 (N_12821,N_12368,N_12303);
nand U12822 (N_12822,N_12355,N_12471);
and U12823 (N_12823,N_12386,N_12438);
nor U12824 (N_12824,N_12456,N_12426);
and U12825 (N_12825,N_12329,N_12325);
and U12826 (N_12826,N_12504,N_12441);
nor U12827 (N_12827,N_12372,N_12441);
nand U12828 (N_12828,N_12340,N_12419);
and U12829 (N_12829,N_12474,N_12331);
nand U12830 (N_12830,N_12450,N_12526);
or U12831 (N_12831,N_12349,N_12491);
nor U12832 (N_12832,N_12496,N_12339);
or U12833 (N_12833,N_12383,N_12418);
xor U12834 (N_12834,N_12474,N_12311);
nor U12835 (N_12835,N_12322,N_12510);
or U12836 (N_12836,N_12509,N_12512);
nor U12837 (N_12837,N_12586,N_12590);
xor U12838 (N_12838,N_12381,N_12501);
nor U12839 (N_12839,N_12341,N_12433);
nor U12840 (N_12840,N_12517,N_12450);
nor U12841 (N_12841,N_12448,N_12362);
and U12842 (N_12842,N_12389,N_12381);
and U12843 (N_12843,N_12499,N_12378);
and U12844 (N_12844,N_12484,N_12362);
xor U12845 (N_12845,N_12451,N_12402);
xor U12846 (N_12846,N_12512,N_12569);
nand U12847 (N_12847,N_12474,N_12561);
and U12848 (N_12848,N_12540,N_12401);
nand U12849 (N_12849,N_12552,N_12373);
or U12850 (N_12850,N_12424,N_12367);
xnor U12851 (N_12851,N_12352,N_12558);
and U12852 (N_12852,N_12419,N_12472);
nor U12853 (N_12853,N_12320,N_12361);
nor U12854 (N_12854,N_12566,N_12353);
nor U12855 (N_12855,N_12558,N_12409);
xor U12856 (N_12856,N_12441,N_12346);
and U12857 (N_12857,N_12479,N_12315);
nand U12858 (N_12858,N_12464,N_12584);
nand U12859 (N_12859,N_12493,N_12313);
or U12860 (N_12860,N_12447,N_12531);
or U12861 (N_12861,N_12330,N_12443);
and U12862 (N_12862,N_12430,N_12373);
or U12863 (N_12863,N_12438,N_12532);
and U12864 (N_12864,N_12465,N_12487);
or U12865 (N_12865,N_12420,N_12541);
or U12866 (N_12866,N_12595,N_12470);
nand U12867 (N_12867,N_12554,N_12369);
and U12868 (N_12868,N_12397,N_12444);
and U12869 (N_12869,N_12596,N_12367);
nor U12870 (N_12870,N_12491,N_12435);
nor U12871 (N_12871,N_12456,N_12474);
and U12872 (N_12872,N_12507,N_12328);
xor U12873 (N_12873,N_12417,N_12530);
nor U12874 (N_12874,N_12354,N_12317);
nand U12875 (N_12875,N_12353,N_12365);
xor U12876 (N_12876,N_12389,N_12463);
xor U12877 (N_12877,N_12312,N_12318);
and U12878 (N_12878,N_12356,N_12565);
nand U12879 (N_12879,N_12304,N_12556);
nor U12880 (N_12880,N_12550,N_12560);
nor U12881 (N_12881,N_12568,N_12371);
xnor U12882 (N_12882,N_12485,N_12416);
and U12883 (N_12883,N_12425,N_12532);
and U12884 (N_12884,N_12427,N_12450);
and U12885 (N_12885,N_12347,N_12346);
xor U12886 (N_12886,N_12378,N_12558);
nor U12887 (N_12887,N_12331,N_12363);
nand U12888 (N_12888,N_12425,N_12463);
and U12889 (N_12889,N_12320,N_12485);
or U12890 (N_12890,N_12538,N_12585);
and U12891 (N_12891,N_12348,N_12486);
xnor U12892 (N_12892,N_12350,N_12451);
nand U12893 (N_12893,N_12332,N_12410);
nand U12894 (N_12894,N_12304,N_12344);
nand U12895 (N_12895,N_12541,N_12333);
and U12896 (N_12896,N_12519,N_12373);
or U12897 (N_12897,N_12327,N_12387);
nand U12898 (N_12898,N_12375,N_12405);
nand U12899 (N_12899,N_12362,N_12423);
or U12900 (N_12900,N_12773,N_12712);
and U12901 (N_12901,N_12653,N_12792);
or U12902 (N_12902,N_12617,N_12696);
xor U12903 (N_12903,N_12723,N_12725);
and U12904 (N_12904,N_12663,N_12673);
and U12905 (N_12905,N_12684,N_12754);
nand U12906 (N_12906,N_12707,N_12685);
nand U12907 (N_12907,N_12644,N_12742);
and U12908 (N_12908,N_12740,N_12724);
nor U12909 (N_12909,N_12711,N_12769);
nand U12910 (N_12910,N_12844,N_12841);
and U12911 (N_12911,N_12749,N_12816);
nor U12912 (N_12912,N_12858,N_12872);
and U12913 (N_12913,N_12869,N_12619);
xnor U12914 (N_12914,N_12873,N_12806);
and U12915 (N_12915,N_12656,N_12836);
and U12916 (N_12916,N_12652,N_12860);
nand U12917 (N_12917,N_12659,N_12842);
nand U12918 (N_12918,N_12857,N_12667);
or U12919 (N_12919,N_12881,N_12618);
and U12920 (N_12920,N_12756,N_12813);
xnor U12921 (N_12921,N_12654,N_12819);
nor U12922 (N_12922,N_12794,N_12761);
xnor U12923 (N_12923,N_12796,N_12829);
nand U12924 (N_12924,N_12783,N_12892);
xor U12925 (N_12925,N_12665,N_12605);
or U12926 (N_12926,N_12637,N_12787);
or U12927 (N_12927,N_12864,N_12720);
or U12928 (N_12928,N_12847,N_12870);
nor U12929 (N_12929,N_12811,N_12885);
nand U12930 (N_12930,N_12833,N_12607);
xnor U12931 (N_12931,N_12883,N_12779);
and U12932 (N_12932,N_12768,N_12703);
nand U12933 (N_12933,N_12780,N_12630);
nor U12934 (N_12934,N_12709,N_12649);
nor U12935 (N_12935,N_12736,N_12631);
nand U12936 (N_12936,N_12784,N_12716);
nand U12937 (N_12937,N_12683,N_12710);
nand U12938 (N_12938,N_12651,N_12731);
nor U12939 (N_12939,N_12638,N_12837);
nor U12940 (N_12940,N_12640,N_12775);
or U12941 (N_12941,N_12818,N_12625);
xor U12942 (N_12942,N_12626,N_12863);
xor U12943 (N_12943,N_12650,N_12601);
nand U12944 (N_12944,N_12647,N_12865);
nand U12945 (N_12945,N_12717,N_12868);
and U12946 (N_12946,N_12680,N_12692);
or U12947 (N_12947,N_12760,N_12677);
and U12948 (N_12948,N_12835,N_12800);
or U12949 (N_12949,N_12895,N_12610);
nand U12950 (N_12950,N_12614,N_12602);
nor U12951 (N_12951,N_12695,N_12777);
nor U12952 (N_12952,N_12606,N_12643);
nand U12953 (N_12953,N_12808,N_12743);
nor U12954 (N_12954,N_12834,N_12661);
and U12955 (N_12955,N_12746,N_12893);
and U12956 (N_12956,N_12752,N_12627);
or U12957 (N_12957,N_12802,N_12807);
xnor U12958 (N_12958,N_12785,N_12702);
or U12959 (N_12959,N_12660,N_12826);
nor U12960 (N_12960,N_12759,N_12822);
nor U12961 (N_12961,N_12762,N_12713);
nand U12962 (N_12962,N_12899,N_12662);
or U12963 (N_12963,N_12880,N_12706);
and U12964 (N_12964,N_12827,N_12632);
nor U12965 (N_12965,N_12633,N_12877);
nor U12966 (N_12966,N_12718,N_12634);
or U12967 (N_12967,N_12642,N_12855);
nand U12968 (N_12968,N_12790,N_12821);
and U12969 (N_12969,N_12705,N_12600);
nand U12970 (N_12970,N_12879,N_12799);
xnor U12971 (N_12971,N_12828,N_12719);
or U12972 (N_12972,N_12699,N_12727);
nand U12973 (N_12973,N_12830,N_12615);
nor U12974 (N_12974,N_12876,N_12809);
or U12975 (N_12975,N_12668,N_12646);
or U12976 (N_12976,N_12636,N_12886);
and U12977 (N_12977,N_12776,N_12875);
nand U12978 (N_12978,N_12758,N_12698);
xor U12979 (N_12979,N_12884,N_12622);
nand U12980 (N_12980,N_12823,N_12657);
nand U12981 (N_12981,N_12609,N_12658);
or U12982 (N_12982,N_12798,N_12848);
nor U12983 (N_12983,N_12890,N_12669);
nand U12984 (N_12984,N_12846,N_12812);
or U12985 (N_12985,N_12898,N_12878);
xnor U12986 (N_12986,N_12810,N_12641);
xnor U12987 (N_12987,N_12803,N_12735);
nand U12988 (N_12988,N_12889,N_12664);
xor U12989 (N_12989,N_12738,N_12888);
and U12990 (N_12990,N_12845,N_12722);
nor U12991 (N_12991,N_12786,N_12882);
nand U12992 (N_12992,N_12734,N_12897);
or U12993 (N_12993,N_12781,N_12804);
nand U12994 (N_12994,N_12853,N_12817);
nor U12995 (N_12995,N_12850,N_12831);
or U12996 (N_12996,N_12765,N_12616);
nand U12997 (N_12997,N_12732,N_12894);
or U12998 (N_12998,N_12851,N_12655);
xor U12999 (N_12999,N_12681,N_12825);
nand U13000 (N_13000,N_12679,N_12690);
and U13001 (N_13001,N_12748,N_12701);
and U13002 (N_13002,N_12603,N_12852);
nor U13003 (N_13003,N_12763,N_12820);
nor U13004 (N_13004,N_12688,N_12824);
nor U13005 (N_13005,N_12739,N_12671);
nor U13006 (N_13006,N_12635,N_12689);
or U13007 (N_13007,N_12861,N_12874);
or U13008 (N_13008,N_12726,N_12862);
and U13009 (N_13009,N_12849,N_12871);
or U13010 (N_13010,N_12751,N_12840);
xor U13011 (N_13011,N_12628,N_12621);
nor U13012 (N_13012,N_12687,N_12791);
nor U13013 (N_13013,N_12793,N_12854);
xnor U13014 (N_13014,N_12623,N_12772);
nand U13015 (N_13015,N_12757,N_12691);
nand U13016 (N_13016,N_12737,N_12859);
and U13017 (N_13017,N_12747,N_12839);
and U13018 (N_13018,N_12715,N_12838);
or U13019 (N_13019,N_12694,N_12867);
and U13020 (N_13020,N_12797,N_12753);
nor U13021 (N_13021,N_12891,N_12782);
nor U13022 (N_13022,N_12645,N_12708);
nand U13023 (N_13023,N_12604,N_12801);
nor U13024 (N_13024,N_12789,N_12704);
nand U13025 (N_13025,N_12730,N_12744);
and U13026 (N_13026,N_12714,N_12729);
xnor U13027 (N_13027,N_12771,N_12612);
or U13028 (N_13028,N_12728,N_12613);
or U13029 (N_13029,N_12805,N_12832);
and U13030 (N_13030,N_12620,N_12896);
and U13031 (N_13031,N_12755,N_12686);
nand U13032 (N_13032,N_12676,N_12750);
nor U13033 (N_13033,N_12624,N_12815);
and U13034 (N_13034,N_12697,N_12672);
nor U13035 (N_13035,N_12678,N_12682);
xnor U13036 (N_13036,N_12741,N_12670);
or U13037 (N_13037,N_12774,N_12629);
nor U13038 (N_13038,N_12611,N_12674);
nand U13039 (N_13039,N_12733,N_12766);
or U13040 (N_13040,N_12666,N_12778);
and U13041 (N_13041,N_12675,N_12795);
nand U13042 (N_13042,N_12745,N_12843);
or U13043 (N_13043,N_12767,N_12770);
nor U13044 (N_13044,N_12887,N_12856);
and U13045 (N_13045,N_12814,N_12648);
nor U13046 (N_13046,N_12788,N_12608);
or U13047 (N_13047,N_12764,N_12700);
nand U13048 (N_13048,N_12639,N_12693);
nand U13049 (N_13049,N_12866,N_12721);
xnor U13050 (N_13050,N_12852,N_12672);
and U13051 (N_13051,N_12707,N_12679);
xnor U13052 (N_13052,N_12732,N_12862);
or U13053 (N_13053,N_12687,N_12711);
and U13054 (N_13054,N_12683,N_12796);
and U13055 (N_13055,N_12738,N_12695);
xor U13056 (N_13056,N_12654,N_12710);
and U13057 (N_13057,N_12605,N_12835);
or U13058 (N_13058,N_12687,N_12807);
xor U13059 (N_13059,N_12747,N_12620);
nor U13060 (N_13060,N_12694,N_12863);
nand U13061 (N_13061,N_12747,N_12864);
xor U13062 (N_13062,N_12862,N_12835);
xnor U13063 (N_13063,N_12671,N_12663);
xor U13064 (N_13064,N_12635,N_12646);
nand U13065 (N_13065,N_12876,N_12756);
or U13066 (N_13066,N_12864,N_12712);
and U13067 (N_13067,N_12648,N_12842);
nand U13068 (N_13068,N_12615,N_12827);
nand U13069 (N_13069,N_12687,N_12835);
nand U13070 (N_13070,N_12770,N_12688);
nor U13071 (N_13071,N_12824,N_12609);
nor U13072 (N_13072,N_12721,N_12623);
nand U13073 (N_13073,N_12688,N_12706);
nand U13074 (N_13074,N_12609,N_12874);
xor U13075 (N_13075,N_12876,N_12764);
xor U13076 (N_13076,N_12875,N_12710);
and U13077 (N_13077,N_12811,N_12707);
xnor U13078 (N_13078,N_12610,N_12879);
or U13079 (N_13079,N_12886,N_12774);
nor U13080 (N_13080,N_12746,N_12801);
or U13081 (N_13081,N_12699,N_12684);
xnor U13082 (N_13082,N_12632,N_12740);
nand U13083 (N_13083,N_12776,N_12882);
or U13084 (N_13084,N_12614,N_12858);
xnor U13085 (N_13085,N_12813,N_12743);
nand U13086 (N_13086,N_12734,N_12723);
or U13087 (N_13087,N_12844,N_12698);
or U13088 (N_13088,N_12790,N_12710);
nand U13089 (N_13089,N_12868,N_12643);
nand U13090 (N_13090,N_12891,N_12762);
and U13091 (N_13091,N_12699,N_12781);
and U13092 (N_13092,N_12724,N_12881);
or U13093 (N_13093,N_12604,N_12830);
or U13094 (N_13094,N_12793,N_12808);
nand U13095 (N_13095,N_12646,N_12822);
and U13096 (N_13096,N_12667,N_12607);
nor U13097 (N_13097,N_12757,N_12649);
nand U13098 (N_13098,N_12830,N_12814);
or U13099 (N_13099,N_12636,N_12637);
or U13100 (N_13100,N_12711,N_12700);
or U13101 (N_13101,N_12712,N_12683);
nand U13102 (N_13102,N_12899,N_12793);
nand U13103 (N_13103,N_12892,N_12810);
nand U13104 (N_13104,N_12662,N_12890);
and U13105 (N_13105,N_12732,N_12688);
nand U13106 (N_13106,N_12663,N_12846);
or U13107 (N_13107,N_12780,N_12786);
nor U13108 (N_13108,N_12666,N_12868);
and U13109 (N_13109,N_12832,N_12885);
nor U13110 (N_13110,N_12667,N_12688);
nand U13111 (N_13111,N_12763,N_12672);
nand U13112 (N_13112,N_12699,N_12824);
and U13113 (N_13113,N_12616,N_12770);
nand U13114 (N_13114,N_12724,N_12673);
and U13115 (N_13115,N_12679,N_12686);
nor U13116 (N_13116,N_12726,N_12779);
nor U13117 (N_13117,N_12789,N_12624);
nor U13118 (N_13118,N_12883,N_12861);
nand U13119 (N_13119,N_12607,N_12726);
or U13120 (N_13120,N_12732,N_12714);
xnor U13121 (N_13121,N_12759,N_12652);
xnor U13122 (N_13122,N_12719,N_12696);
nand U13123 (N_13123,N_12656,N_12892);
or U13124 (N_13124,N_12625,N_12899);
and U13125 (N_13125,N_12733,N_12640);
or U13126 (N_13126,N_12624,N_12670);
and U13127 (N_13127,N_12778,N_12688);
nor U13128 (N_13128,N_12669,N_12635);
and U13129 (N_13129,N_12651,N_12807);
nor U13130 (N_13130,N_12654,N_12877);
nor U13131 (N_13131,N_12833,N_12862);
nand U13132 (N_13132,N_12721,N_12705);
and U13133 (N_13133,N_12642,N_12846);
and U13134 (N_13134,N_12890,N_12774);
nand U13135 (N_13135,N_12862,N_12675);
xnor U13136 (N_13136,N_12607,N_12658);
and U13137 (N_13137,N_12787,N_12746);
nor U13138 (N_13138,N_12631,N_12616);
nand U13139 (N_13139,N_12667,N_12657);
and U13140 (N_13140,N_12713,N_12614);
xnor U13141 (N_13141,N_12832,N_12772);
nor U13142 (N_13142,N_12766,N_12838);
nor U13143 (N_13143,N_12809,N_12625);
xor U13144 (N_13144,N_12845,N_12864);
nor U13145 (N_13145,N_12809,N_12741);
xor U13146 (N_13146,N_12664,N_12776);
nor U13147 (N_13147,N_12806,N_12693);
or U13148 (N_13148,N_12616,N_12665);
nand U13149 (N_13149,N_12888,N_12883);
nor U13150 (N_13150,N_12736,N_12615);
or U13151 (N_13151,N_12865,N_12746);
nor U13152 (N_13152,N_12889,N_12635);
nand U13153 (N_13153,N_12766,N_12854);
xor U13154 (N_13154,N_12619,N_12708);
xnor U13155 (N_13155,N_12865,N_12718);
or U13156 (N_13156,N_12788,N_12684);
and U13157 (N_13157,N_12757,N_12602);
nor U13158 (N_13158,N_12743,N_12774);
xor U13159 (N_13159,N_12656,N_12762);
xor U13160 (N_13160,N_12719,N_12667);
or U13161 (N_13161,N_12741,N_12663);
nand U13162 (N_13162,N_12891,N_12850);
xnor U13163 (N_13163,N_12886,N_12793);
or U13164 (N_13164,N_12825,N_12787);
xor U13165 (N_13165,N_12644,N_12661);
nand U13166 (N_13166,N_12652,N_12665);
nand U13167 (N_13167,N_12893,N_12614);
and U13168 (N_13168,N_12689,N_12641);
or U13169 (N_13169,N_12654,N_12632);
and U13170 (N_13170,N_12751,N_12882);
xnor U13171 (N_13171,N_12603,N_12624);
xor U13172 (N_13172,N_12739,N_12889);
nor U13173 (N_13173,N_12819,N_12757);
xnor U13174 (N_13174,N_12677,N_12846);
xor U13175 (N_13175,N_12709,N_12725);
xor U13176 (N_13176,N_12694,N_12895);
nor U13177 (N_13177,N_12791,N_12621);
nand U13178 (N_13178,N_12788,N_12805);
nor U13179 (N_13179,N_12843,N_12651);
nand U13180 (N_13180,N_12750,N_12881);
or U13181 (N_13181,N_12692,N_12800);
nand U13182 (N_13182,N_12826,N_12881);
and U13183 (N_13183,N_12822,N_12708);
nand U13184 (N_13184,N_12693,N_12648);
or U13185 (N_13185,N_12765,N_12804);
or U13186 (N_13186,N_12826,N_12864);
nand U13187 (N_13187,N_12691,N_12614);
and U13188 (N_13188,N_12737,N_12785);
and U13189 (N_13189,N_12786,N_12751);
and U13190 (N_13190,N_12601,N_12740);
or U13191 (N_13191,N_12796,N_12692);
and U13192 (N_13192,N_12736,N_12646);
xor U13193 (N_13193,N_12806,N_12704);
xnor U13194 (N_13194,N_12805,N_12721);
or U13195 (N_13195,N_12836,N_12811);
and U13196 (N_13196,N_12611,N_12711);
nand U13197 (N_13197,N_12761,N_12724);
or U13198 (N_13198,N_12788,N_12629);
or U13199 (N_13199,N_12784,N_12796);
nand U13200 (N_13200,N_13085,N_13069);
nor U13201 (N_13201,N_13164,N_13084);
nand U13202 (N_13202,N_13010,N_13186);
or U13203 (N_13203,N_12935,N_13181);
and U13204 (N_13204,N_13185,N_13045);
or U13205 (N_13205,N_13016,N_13126);
or U13206 (N_13206,N_12946,N_12918);
nand U13207 (N_13207,N_12930,N_12968);
xnor U13208 (N_13208,N_12965,N_13090);
or U13209 (N_13209,N_13188,N_12914);
or U13210 (N_13210,N_12923,N_13110);
and U13211 (N_13211,N_12979,N_13158);
nand U13212 (N_13212,N_12901,N_13091);
or U13213 (N_13213,N_12949,N_12953);
or U13214 (N_13214,N_13075,N_13159);
xnor U13215 (N_13215,N_12992,N_12943);
and U13216 (N_13216,N_13190,N_12947);
nor U13217 (N_13217,N_12950,N_12927);
and U13218 (N_13218,N_12996,N_13080);
and U13219 (N_13219,N_13049,N_13003);
or U13220 (N_13220,N_13054,N_13172);
nand U13221 (N_13221,N_13020,N_13169);
nor U13222 (N_13222,N_13098,N_13155);
and U13223 (N_13223,N_13025,N_12998);
xor U13224 (N_13224,N_13150,N_13099);
nand U13225 (N_13225,N_13145,N_12959);
nor U13226 (N_13226,N_12920,N_13013);
nand U13227 (N_13227,N_12937,N_12915);
nand U13228 (N_13228,N_13177,N_13064);
nor U13229 (N_13229,N_13160,N_13102);
and U13230 (N_13230,N_13122,N_13133);
nand U13231 (N_13231,N_13047,N_13026);
nor U13232 (N_13232,N_13115,N_12912);
nor U13233 (N_13233,N_13193,N_13142);
and U13234 (N_13234,N_13140,N_13079);
nor U13235 (N_13235,N_13139,N_13125);
nand U13236 (N_13236,N_12907,N_12986);
nor U13237 (N_13237,N_12906,N_12970);
or U13238 (N_13238,N_12972,N_13093);
xnor U13239 (N_13239,N_12989,N_13116);
or U13240 (N_13240,N_12981,N_13006);
xnor U13241 (N_13241,N_13004,N_13101);
nor U13242 (N_13242,N_12971,N_13118);
or U13243 (N_13243,N_12969,N_13008);
xnor U13244 (N_13244,N_13103,N_13019);
and U13245 (N_13245,N_13015,N_13114);
or U13246 (N_13246,N_12908,N_13053);
xnor U13247 (N_13247,N_13162,N_13048);
nor U13248 (N_13248,N_12929,N_13073);
xor U13249 (N_13249,N_12917,N_13127);
nor U13250 (N_13250,N_12911,N_13152);
and U13251 (N_13251,N_13123,N_13174);
xor U13252 (N_13252,N_12940,N_12980);
and U13253 (N_13253,N_13119,N_12990);
and U13254 (N_13254,N_12994,N_13149);
and U13255 (N_13255,N_13061,N_13068);
or U13256 (N_13256,N_13144,N_13024);
or U13257 (N_13257,N_13043,N_13196);
and U13258 (N_13258,N_12904,N_13167);
xor U13259 (N_13259,N_12941,N_13021);
nand U13260 (N_13260,N_13011,N_13175);
nor U13261 (N_13261,N_13154,N_13109);
or U13262 (N_13262,N_13082,N_12932);
nor U13263 (N_13263,N_13179,N_13106);
and U13264 (N_13264,N_13183,N_13141);
xor U13265 (N_13265,N_12956,N_12945);
nand U13266 (N_13266,N_13129,N_12955);
xor U13267 (N_13267,N_12985,N_12926);
nand U13268 (N_13268,N_12963,N_13178);
nand U13269 (N_13269,N_13131,N_12976);
xnor U13270 (N_13270,N_13198,N_13124);
xor U13271 (N_13271,N_12988,N_12997);
or U13272 (N_13272,N_12952,N_13030);
xnor U13273 (N_13273,N_12944,N_13072);
nor U13274 (N_13274,N_12948,N_13143);
xor U13275 (N_13275,N_13094,N_13096);
and U13276 (N_13276,N_12987,N_12924);
nand U13277 (N_13277,N_12903,N_13168);
or U13278 (N_13278,N_13166,N_12999);
nor U13279 (N_13279,N_13088,N_12993);
or U13280 (N_13280,N_13022,N_13074);
and U13281 (N_13281,N_12922,N_12966);
nor U13282 (N_13282,N_12919,N_12916);
or U13283 (N_13283,N_13033,N_13037);
and U13284 (N_13284,N_12982,N_12954);
xor U13285 (N_13285,N_13042,N_12960);
and U13286 (N_13286,N_13121,N_12905);
nor U13287 (N_13287,N_13182,N_13194);
and U13288 (N_13288,N_13189,N_13039);
or U13289 (N_13289,N_12995,N_13113);
xor U13290 (N_13290,N_12974,N_13146);
nand U13291 (N_13291,N_13195,N_12962);
or U13292 (N_13292,N_13184,N_13040);
xor U13293 (N_13293,N_13062,N_13029);
or U13294 (N_13294,N_12925,N_13035);
nor U13295 (N_13295,N_13086,N_13031);
or U13296 (N_13296,N_12967,N_13170);
and U13297 (N_13297,N_13161,N_13067);
xnor U13298 (N_13298,N_13057,N_12913);
nand U13299 (N_13299,N_12957,N_12991);
nor U13300 (N_13300,N_13055,N_13180);
nand U13301 (N_13301,N_12951,N_13009);
xor U13302 (N_13302,N_13136,N_12977);
nand U13303 (N_13303,N_13134,N_13089);
xor U13304 (N_13304,N_13078,N_13001);
nand U13305 (N_13305,N_13100,N_13017);
nand U13306 (N_13306,N_13128,N_13192);
and U13307 (N_13307,N_13148,N_13111);
or U13308 (N_13308,N_12938,N_12961);
or U13309 (N_13309,N_12909,N_13081);
or U13310 (N_13310,N_13032,N_13063);
nand U13311 (N_13311,N_13046,N_13151);
nand U13312 (N_13312,N_12942,N_13171);
xor U13313 (N_13313,N_13105,N_13130);
and U13314 (N_13314,N_13058,N_13157);
xor U13315 (N_13315,N_12984,N_13066);
and U13316 (N_13316,N_13012,N_13176);
or U13317 (N_13317,N_13147,N_12936);
nand U13318 (N_13318,N_13059,N_12900);
and U13319 (N_13319,N_13197,N_13137);
and U13320 (N_13320,N_13095,N_13076);
nor U13321 (N_13321,N_13056,N_12933);
xnor U13322 (N_13322,N_12939,N_13187);
xor U13323 (N_13323,N_13087,N_13117);
and U13324 (N_13324,N_13173,N_12958);
nand U13325 (N_13325,N_13191,N_12983);
or U13326 (N_13326,N_13156,N_12902);
nand U13327 (N_13327,N_13052,N_12934);
or U13328 (N_13328,N_13071,N_13000);
nand U13329 (N_13329,N_13153,N_13051);
nand U13330 (N_13330,N_12964,N_13097);
or U13331 (N_13331,N_13018,N_12973);
or U13332 (N_13332,N_13034,N_13135);
nor U13333 (N_13333,N_13038,N_13023);
nand U13334 (N_13334,N_12975,N_13104);
nand U13335 (N_13335,N_13036,N_13112);
nand U13336 (N_13336,N_13083,N_13007);
xor U13337 (N_13337,N_13060,N_13107);
nor U13338 (N_13338,N_13028,N_12978);
xnor U13339 (N_13339,N_13005,N_13044);
and U13340 (N_13340,N_13138,N_13132);
nor U13341 (N_13341,N_13065,N_13050);
or U13342 (N_13342,N_13163,N_13077);
nor U13343 (N_13343,N_12928,N_13041);
nand U13344 (N_13344,N_13120,N_12931);
nand U13345 (N_13345,N_13002,N_13014);
nand U13346 (N_13346,N_13027,N_12910);
and U13347 (N_13347,N_13092,N_13108);
or U13348 (N_13348,N_13165,N_13070);
nor U13349 (N_13349,N_12921,N_13199);
or U13350 (N_13350,N_12906,N_12983);
and U13351 (N_13351,N_13086,N_13173);
nor U13352 (N_13352,N_12975,N_13052);
nor U13353 (N_13353,N_12951,N_12945);
or U13354 (N_13354,N_13143,N_13112);
xnor U13355 (N_13355,N_13142,N_13043);
or U13356 (N_13356,N_13179,N_13093);
or U13357 (N_13357,N_12923,N_12924);
and U13358 (N_13358,N_12908,N_12945);
and U13359 (N_13359,N_12909,N_13163);
nor U13360 (N_13360,N_13132,N_13066);
or U13361 (N_13361,N_13175,N_12984);
nand U13362 (N_13362,N_12962,N_13031);
xor U13363 (N_13363,N_12907,N_13078);
and U13364 (N_13364,N_13164,N_13111);
and U13365 (N_13365,N_13045,N_13071);
nand U13366 (N_13366,N_13121,N_13159);
xor U13367 (N_13367,N_12919,N_13038);
xnor U13368 (N_13368,N_13161,N_13182);
or U13369 (N_13369,N_12954,N_13044);
nor U13370 (N_13370,N_13133,N_12948);
and U13371 (N_13371,N_13002,N_12933);
nor U13372 (N_13372,N_13070,N_13062);
or U13373 (N_13373,N_13113,N_12918);
xnor U13374 (N_13374,N_13088,N_13121);
nor U13375 (N_13375,N_13026,N_13129);
and U13376 (N_13376,N_12936,N_12916);
or U13377 (N_13377,N_13052,N_12953);
and U13378 (N_13378,N_13108,N_12959);
or U13379 (N_13379,N_13034,N_12948);
or U13380 (N_13380,N_12904,N_13124);
nand U13381 (N_13381,N_12938,N_12914);
xnor U13382 (N_13382,N_13035,N_13026);
and U13383 (N_13383,N_13175,N_13096);
and U13384 (N_13384,N_13058,N_12932);
nor U13385 (N_13385,N_13031,N_13188);
nand U13386 (N_13386,N_13055,N_12917);
and U13387 (N_13387,N_12928,N_13155);
nor U13388 (N_13388,N_12917,N_12960);
or U13389 (N_13389,N_13190,N_13127);
or U13390 (N_13390,N_12908,N_12990);
or U13391 (N_13391,N_13188,N_12994);
or U13392 (N_13392,N_12963,N_12903);
xnor U13393 (N_13393,N_13002,N_13053);
nand U13394 (N_13394,N_13063,N_13195);
xnor U13395 (N_13395,N_13177,N_13086);
or U13396 (N_13396,N_13104,N_12946);
xnor U13397 (N_13397,N_13023,N_13099);
nand U13398 (N_13398,N_13177,N_12900);
or U13399 (N_13399,N_13104,N_12933);
nand U13400 (N_13400,N_13170,N_13153);
xor U13401 (N_13401,N_13113,N_13080);
and U13402 (N_13402,N_13156,N_13165);
nor U13403 (N_13403,N_12938,N_12904);
nand U13404 (N_13404,N_13016,N_12962);
or U13405 (N_13405,N_12956,N_13181);
nand U13406 (N_13406,N_13098,N_12945);
xor U13407 (N_13407,N_13023,N_12985);
or U13408 (N_13408,N_13167,N_13042);
or U13409 (N_13409,N_12927,N_13163);
xnor U13410 (N_13410,N_13199,N_13160);
nor U13411 (N_13411,N_13161,N_12947);
and U13412 (N_13412,N_13091,N_12912);
and U13413 (N_13413,N_13076,N_13105);
and U13414 (N_13414,N_12953,N_13024);
and U13415 (N_13415,N_13181,N_12965);
nand U13416 (N_13416,N_13078,N_12944);
nand U13417 (N_13417,N_12984,N_13130);
and U13418 (N_13418,N_13096,N_13015);
nand U13419 (N_13419,N_13188,N_13085);
xor U13420 (N_13420,N_13168,N_13055);
xnor U13421 (N_13421,N_13150,N_13158);
nand U13422 (N_13422,N_13195,N_12910);
nor U13423 (N_13423,N_12951,N_13080);
and U13424 (N_13424,N_13140,N_12941);
xor U13425 (N_13425,N_13170,N_13199);
or U13426 (N_13426,N_13068,N_13026);
or U13427 (N_13427,N_12926,N_12994);
nor U13428 (N_13428,N_12971,N_13102);
nand U13429 (N_13429,N_13005,N_12985);
and U13430 (N_13430,N_13019,N_12911);
nor U13431 (N_13431,N_12965,N_13010);
nand U13432 (N_13432,N_13104,N_12953);
or U13433 (N_13433,N_13181,N_13083);
or U13434 (N_13434,N_12943,N_12903);
or U13435 (N_13435,N_13050,N_13075);
nand U13436 (N_13436,N_13120,N_13042);
nand U13437 (N_13437,N_12963,N_13008);
nor U13438 (N_13438,N_12965,N_13041);
or U13439 (N_13439,N_12908,N_12942);
and U13440 (N_13440,N_12915,N_13032);
or U13441 (N_13441,N_12908,N_13140);
nor U13442 (N_13442,N_13178,N_12966);
or U13443 (N_13443,N_12996,N_12994);
nand U13444 (N_13444,N_13039,N_13119);
or U13445 (N_13445,N_13196,N_13111);
nor U13446 (N_13446,N_13181,N_13088);
or U13447 (N_13447,N_12976,N_13185);
nand U13448 (N_13448,N_13072,N_12969);
and U13449 (N_13449,N_13146,N_12929);
nor U13450 (N_13450,N_12968,N_13064);
nand U13451 (N_13451,N_12951,N_13167);
nor U13452 (N_13452,N_13043,N_13097);
and U13453 (N_13453,N_13003,N_13183);
or U13454 (N_13454,N_13039,N_12928);
xor U13455 (N_13455,N_12907,N_13072);
nand U13456 (N_13456,N_13171,N_13180);
nor U13457 (N_13457,N_12954,N_13073);
and U13458 (N_13458,N_13038,N_12900);
and U13459 (N_13459,N_13012,N_12948);
xor U13460 (N_13460,N_13126,N_13168);
and U13461 (N_13461,N_13071,N_13148);
and U13462 (N_13462,N_13049,N_13052);
xor U13463 (N_13463,N_13176,N_12928);
nand U13464 (N_13464,N_13035,N_12956);
nand U13465 (N_13465,N_13117,N_13191);
or U13466 (N_13466,N_13120,N_12937);
xnor U13467 (N_13467,N_13102,N_13082);
nor U13468 (N_13468,N_13155,N_13080);
and U13469 (N_13469,N_13189,N_13062);
or U13470 (N_13470,N_13000,N_13173);
and U13471 (N_13471,N_13086,N_13084);
or U13472 (N_13472,N_13078,N_13138);
xnor U13473 (N_13473,N_13054,N_13176);
nor U13474 (N_13474,N_13165,N_13074);
nand U13475 (N_13475,N_13087,N_12982);
or U13476 (N_13476,N_12958,N_13154);
nor U13477 (N_13477,N_12900,N_12978);
and U13478 (N_13478,N_12959,N_13033);
nor U13479 (N_13479,N_13148,N_13176);
and U13480 (N_13480,N_12993,N_12927);
or U13481 (N_13481,N_13134,N_12900);
nor U13482 (N_13482,N_13161,N_12964);
or U13483 (N_13483,N_12936,N_12990);
nor U13484 (N_13484,N_12987,N_12995);
xnor U13485 (N_13485,N_12921,N_12960);
nor U13486 (N_13486,N_13035,N_13021);
or U13487 (N_13487,N_13105,N_13047);
nand U13488 (N_13488,N_13096,N_13198);
and U13489 (N_13489,N_13171,N_12927);
xnor U13490 (N_13490,N_13014,N_13024);
nor U13491 (N_13491,N_13006,N_12954);
nor U13492 (N_13492,N_13055,N_13054);
nor U13493 (N_13493,N_13098,N_13001);
nand U13494 (N_13494,N_12983,N_13180);
and U13495 (N_13495,N_13188,N_13009);
xor U13496 (N_13496,N_13141,N_13120);
and U13497 (N_13497,N_13104,N_12921);
or U13498 (N_13498,N_13088,N_12973);
nor U13499 (N_13499,N_12950,N_13152);
and U13500 (N_13500,N_13348,N_13469);
and U13501 (N_13501,N_13374,N_13308);
nand U13502 (N_13502,N_13331,N_13358);
or U13503 (N_13503,N_13325,N_13262);
xnor U13504 (N_13504,N_13444,N_13216);
xor U13505 (N_13505,N_13356,N_13496);
xnor U13506 (N_13506,N_13386,N_13457);
xnor U13507 (N_13507,N_13284,N_13230);
and U13508 (N_13508,N_13468,N_13416);
or U13509 (N_13509,N_13210,N_13251);
nand U13510 (N_13510,N_13245,N_13345);
nand U13511 (N_13511,N_13406,N_13476);
xnor U13512 (N_13512,N_13277,N_13229);
nand U13513 (N_13513,N_13253,N_13322);
xnor U13514 (N_13514,N_13340,N_13353);
nand U13515 (N_13515,N_13368,N_13419);
nand U13516 (N_13516,N_13391,N_13381);
nor U13517 (N_13517,N_13370,N_13414);
nor U13518 (N_13518,N_13423,N_13236);
and U13519 (N_13519,N_13385,N_13479);
and U13520 (N_13520,N_13237,N_13227);
and U13521 (N_13521,N_13217,N_13330);
and U13522 (N_13522,N_13213,N_13267);
and U13523 (N_13523,N_13394,N_13300);
or U13524 (N_13524,N_13412,N_13280);
nand U13525 (N_13525,N_13393,N_13424);
and U13526 (N_13526,N_13256,N_13328);
and U13527 (N_13527,N_13366,N_13221);
and U13528 (N_13528,N_13460,N_13373);
xnor U13529 (N_13529,N_13465,N_13302);
or U13530 (N_13530,N_13248,N_13379);
nand U13531 (N_13531,N_13288,N_13321);
nor U13532 (N_13532,N_13411,N_13413);
or U13533 (N_13533,N_13326,N_13360);
nand U13534 (N_13534,N_13285,N_13390);
or U13535 (N_13535,N_13304,N_13456);
or U13536 (N_13536,N_13455,N_13486);
and U13537 (N_13537,N_13264,N_13266);
and U13538 (N_13538,N_13343,N_13427);
and U13539 (N_13539,N_13259,N_13276);
and U13540 (N_13540,N_13305,N_13231);
xnor U13541 (N_13541,N_13323,N_13378);
nand U13542 (N_13542,N_13405,N_13293);
xnor U13543 (N_13543,N_13403,N_13281);
nand U13544 (N_13544,N_13319,N_13338);
xor U13545 (N_13545,N_13329,N_13399);
or U13546 (N_13546,N_13498,N_13470);
xnor U13547 (N_13547,N_13382,N_13337);
xor U13548 (N_13548,N_13438,N_13485);
nor U13549 (N_13549,N_13417,N_13309);
nand U13550 (N_13550,N_13472,N_13449);
and U13551 (N_13551,N_13223,N_13235);
or U13552 (N_13552,N_13362,N_13436);
or U13553 (N_13553,N_13240,N_13349);
nand U13554 (N_13554,N_13352,N_13278);
or U13555 (N_13555,N_13257,N_13234);
or U13556 (N_13556,N_13467,N_13206);
nor U13557 (N_13557,N_13282,N_13314);
or U13558 (N_13558,N_13272,N_13415);
or U13559 (N_13559,N_13222,N_13320);
nor U13560 (N_13560,N_13224,N_13484);
xor U13561 (N_13561,N_13474,N_13493);
or U13562 (N_13562,N_13312,N_13473);
or U13563 (N_13563,N_13260,N_13471);
xor U13564 (N_13564,N_13303,N_13376);
and U13565 (N_13565,N_13487,N_13244);
and U13566 (N_13566,N_13316,N_13355);
and U13567 (N_13567,N_13464,N_13211);
or U13568 (N_13568,N_13334,N_13269);
nand U13569 (N_13569,N_13202,N_13425);
nor U13570 (N_13570,N_13250,N_13418);
nor U13571 (N_13571,N_13261,N_13357);
nor U13572 (N_13572,N_13387,N_13306);
or U13573 (N_13573,N_13365,N_13480);
xnor U13574 (N_13574,N_13341,N_13311);
and U13575 (N_13575,N_13428,N_13238);
nor U13576 (N_13576,N_13246,N_13317);
xor U13577 (N_13577,N_13454,N_13453);
and U13578 (N_13578,N_13431,N_13220);
xnor U13579 (N_13579,N_13388,N_13380);
xnor U13580 (N_13580,N_13344,N_13233);
and U13581 (N_13581,N_13258,N_13483);
xnor U13582 (N_13582,N_13494,N_13429);
nand U13583 (N_13583,N_13273,N_13361);
nor U13584 (N_13584,N_13342,N_13477);
xnor U13585 (N_13585,N_13478,N_13315);
or U13586 (N_13586,N_13441,N_13292);
xor U13587 (N_13587,N_13402,N_13241);
nor U13588 (N_13588,N_13283,N_13327);
xnor U13589 (N_13589,N_13203,N_13219);
nor U13590 (N_13590,N_13201,N_13296);
or U13591 (N_13591,N_13243,N_13249);
nand U13592 (N_13592,N_13218,N_13286);
xor U13593 (N_13593,N_13497,N_13482);
or U13594 (N_13594,N_13268,N_13437);
nor U13595 (N_13595,N_13481,N_13205);
nand U13596 (N_13596,N_13270,N_13377);
or U13597 (N_13597,N_13242,N_13462);
and U13598 (N_13598,N_13452,N_13488);
and U13599 (N_13599,N_13422,N_13265);
nor U13600 (N_13600,N_13208,N_13332);
or U13601 (N_13601,N_13207,N_13212);
nor U13602 (N_13602,N_13301,N_13499);
nor U13603 (N_13603,N_13410,N_13463);
and U13604 (N_13604,N_13297,N_13307);
or U13605 (N_13605,N_13400,N_13447);
nand U13606 (N_13606,N_13346,N_13398);
or U13607 (N_13607,N_13299,N_13443);
nand U13608 (N_13608,N_13274,N_13290);
and U13609 (N_13609,N_13351,N_13430);
and U13610 (N_13610,N_13445,N_13458);
and U13611 (N_13611,N_13318,N_13433);
and U13612 (N_13612,N_13407,N_13310);
nor U13613 (N_13613,N_13263,N_13448);
xnor U13614 (N_13614,N_13408,N_13369);
nor U13615 (N_13615,N_13459,N_13492);
xor U13616 (N_13616,N_13275,N_13409);
nand U13617 (N_13617,N_13215,N_13295);
xor U13618 (N_13618,N_13232,N_13367);
or U13619 (N_13619,N_13491,N_13435);
xor U13620 (N_13620,N_13350,N_13446);
xnor U13621 (N_13621,N_13324,N_13466);
and U13622 (N_13622,N_13279,N_13461);
xor U13623 (N_13623,N_13371,N_13384);
nand U13624 (N_13624,N_13333,N_13354);
nand U13625 (N_13625,N_13298,N_13372);
xnor U13626 (N_13626,N_13420,N_13252);
nor U13627 (N_13627,N_13395,N_13247);
nand U13628 (N_13628,N_13255,N_13363);
xnor U13629 (N_13629,N_13432,N_13439);
or U13630 (N_13630,N_13375,N_13383);
nand U13631 (N_13631,N_13495,N_13440);
nand U13632 (N_13632,N_13397,N_13294);
and U13633 (N_13633,N_13489,N_13287);
and U13634 (N_13634,N_13359,N_13347);
nor U13635 (N_13635,N_13271,N_13339);
xor U13636 (N_13636,N_13313,N_13214);
nand U13637 (N_13637,N_13291,N_13204);
xor U13638 (N_13638,N_13426,N_13404);
and U13639 (N_13639,N_13451,N_13401);
nand U13640 (N_13640,N_13434,N_13209);
and U13641 (N_13641,N_13392,N_13364);
nand U13642 (N_13642,N_13254,N_13226);
xor U13643 (N_13643,N_13475,N_13421);
nor U13644 (N_13644,N_13289,N_13239);
or U13645 (N_13645,N_13442,N_13450);
xor U13646 (N_13646,N_13200,N_13228);
nand U13647 (N_13647,N_13225,N_13336);
and U13648 (N_13648,N_13389,N_13396);
nor U13649 (N_13649,N_13490,N_13335);
or U13650 (N_13650,N_13318,N_13361);
nand U13651 (N_13651,N_13433,N_13315);
and U13652 (N_13652,N_13318,N_13423);
and U13653 (N_13653,N_13238,N_13491);
nor U13654 (N_13654,N_13495,N_13431);
and U13655 (N_13655,N_13264,N_13297);
or U13656 (N_13656,N_13315,N_13262);
or U13657 (N_13657,N_13234,N_13496);
or U13658 (N_13658,N_13404,N_13441);
or U13659 (N_13659,N_13388,N_13426);
and U13660 (N_13660,N_13248,N_13260);
and U13661 (N_13661,N_13499,N_13351);
nand U13662 (N_13662,N_13247,N_13308);
and U13663 (N_13663,N_13465,N_13456);
or U13664 (N_13664,N_13215,N_13484);
xor U13665 (N_13665,N_13294,N_13461);
or U13666 (N_13666,N_13419,N_13427);
and U13667 (N_13667,N_13364,N_13214);
nor U13668 (N_13668,N_13311,N_13498);
nand U13669 (N_13669,N_13451,N_13415);
nand U13670 (N_13670,N_13309,N_13429);
and U13671 (N_13671,N_13399,N_13289);
xnor U13672 (N_13672,N_13307,N_13352);
nor U13673 (N_13673,N_13423,N_13266);
nand U13674 (N_13674,N_13289,N_13246);
and U13675 (N_13675,N_13365,N_13282);
nand U13676 (N_13676,N_13458,N_13338);
and U13677 (N_13677,N_13317,N_13316);
xor U13678 (N_13678,N_13434,N_13495);
nor U13679 (N_13679,N_13303,N_13413);
xor U13680 (N_13680,N_13427,N_13371);
and U13681 (N_13681,N_13285,N_13327);
or U13682 (N_13682,N_13358,N_13381);
nand U13683 (N_13683,N_13201,N_13491);
or U13684 (N_13684,N_13275,N_13407);
and U13685 (N_13685,N_13463,N_13270);
or U13686 (N_13686,N_13235,N_13421);
or U13687 (N_13687,N_13360,N_13240);
xnor U13688 (N_13688,N_13288,N_13475);
and U13689 (N_13689,N_13373,N_13240);
nor U13690 (N_13690,N_13280,N_13238);
nor U13691 (N_13691,N_13257,N_13497);
or U13692 (N_13692,N_13400,N_13267);
xnor U13693 (N_13693,N_13231,N_13395);
and U13694 (N_13694,N_13464,N_13345);
and U13695 (N_13695,N_13412,N_13474);
xor U13696 (N_13696,N_13452,N_13203);
nand U13697 (N_13697,N_13306,N_13470);
xnor U13698 (N_13698,N_13279,N_13411);
or U13699 (N_13699,N_13496,N_13434);
and U13700 (N_13700,N_13456,N_13275);
and U13701 (N_13701,N_13489,N_13357);
nor U13702 (N_13702,N_13419,N_13391);
xnor U13703 (N_13703,N_13217,N_13237);
and U13704 (N_13704,N_13217,N_13218);
nor U13705 (N_13705,N_13254,N_13261);
xor U13706 (N_13706,N_13344,N_13468);
and U13707 (N_13707,N_13329,N_13210);
nand U13708 (N_13708,N_13330,N_13444);
nor U13709 (N_13709,N_13391,N_13480);
and U13710 (N_13710,N_13235,N_13230);
nor U13711 (N_13711,N_13284,N_13232);
xor U13712 (N_13712,N_13465,N_13497);
or U13713 (N_13713,N_13372,N_13379);
and U13714 (N_13714,N_13440,N_13208);
nand U13715 (N_13715,N_13228,N_13324);
nand U13716 (N_13716,N_13490,N_13329);
xnor U13717 (N_13717,N_13429,N_13371);
nand U13718 (N_13718,N_13302,N_13482);
nor U13719 (N_13719,N_13313,N_13334);
nor U13720 (N_13720,N_13302,N_13471);
and U13721 (N_13721,N_13395,N_13451);
or U13722 (N_13722,N_13490,N_13203);
xor U13723 (N_13723,N_13419,N_13428);
and U13724 (N_13724,N_13205,N_13225);
or U13725 (N_13725,N_13379,N_13252);
nand U13726 (N_13726,N_13413,N_13323);
and U13727 (N_13727,N_13278,N_13399);
xnor U13728 (N_13728,N_13287,N_13349);
and U13729 (N_13729,N_13416,N_13450);
xnor U13730 (N_13730,N_13429,N_13317);
or U13731 (N_13731,N_13448,N_13336);
nor U13732 (N_13732,N_13208,N_13397);
nand U13733 (N_13733,N_13377,N_13399);
nand U13734 (N_13734,N_13442,N_13245);
nand U13735 (N_13735,N_13275,N_13376);
or U13736 (N_13736,N_13430,N_13378);
nor U13737 (N_13737,N_13299,N_13498);
nor U13738 (N_13738,N_13394,N_13319);
or U13739 (N_13739,N_13212,N_13215);
xnor U13740 (N_13740,N_13469,N_13287);
nand U13741 (N_13741,N_13438,N_13240);
nor U13742 (N_13742,N_13467,N_13248);
or U13743 (N_13743,N_13490,N_13257);
xor U13744 (N_13744,N_13485,N_13399);
or U13745 (N_13745,N_13343,N_13455);
or U13746 (N_13746,N_13296,N_13430);
or U13747 (N_13747,N_13212,N_13420);
or U13748 (N_13748,N_13488,N_13334);
or U13749 (N_13749,N_13499,N_13345);
and U13750 (N_13750,N_13362,N_13275);
nand U13751 (N_13751,N_13411,N_13325);
nor U13752 (N_13752,N_13498,N_13277);
or U13753 (N_13753,N_13429,N_13302);
and U13754 (N_13754,N_13228,N_13345);
nand U13755 (N_13755,N_13493,N_13491);
nand U13756 (N_13756,N_13257,N_13498);
nand U13757 (N_13757,N_13477,N_13236);
nor U13758 (N_13758,N_13405,N_13251);
and U13759 (N_13759,N_13418,N_13275);
nand U13760 (N_13760,N_13320,N_13417);
and U13761 (N_13761,N_13468,N_13466);
and U13762 (N_13762,N_13489,N_13484);
and U13763 (N_13763,N_13426,N_13213);
and U13764 (N_13764,N_13327,N_13313);
xor U13765 (N_13765,N_13283,N_13221);
and U13766 (N_13766,N_13314,N_13456);
or U13767 (N_13767,N_13268,N_13229);
or U13768 (N_13768,N_13419,N_13326);
and U13769 (N_13769,N_13388,N_13210);
or U13770 (N_13770,N_13439,N_13456);
nand U13771 (N_13771,N_13411,N_13457);
xnor U13772 (N_13772,N_13322,N_13409);
or U13773 (N_13773,N_13383,N_13363);
and U13774 (N_13774,N_13383,N_13285);
xnor U13775 (N_13775,N_13311,N_13444);
and U13776 (N_13776,N_13306,N_13461);
xnor U13777 (N_13777,N_13295,N_13492);
or U13778 (N_13778,N_13427,N_13330);
nor U13779 (N_13779,N_13233,N_13225);
xor U13780 (N_13780,N_13475,N_13383);
and U13781 (N_13781,N_13368,N_13249);
nor U13782 (N_13782,N_13367,N_13221);
and U13783 (N_13783,N_13276,N_13294);
nor U13784 (N_13784,N_13331,N_13405);
and U13785 (N_13785,N_13338,N_13253);
xor U13786 (N_13786,N_13331,N_13284);
and U13787 (N_13787,N_13452,N_13219);
and U13788 (N_13788,N_13218,N_13465);
and U13789 (N_13789,N_13222,N_13245);
or U13790 (N_13790,N_13208,N_13472);
xor U13791 (N_13791,N_13287,N_13451);
xnor U13792 (N_13792,N_13365,N_13405);
or U13793 (N_13793,N_13293,N_13354);
nand U13794 (N_13794,N_13307,N_13461);
or U13795 (N_13795,N_13300,N_13274);
and U13796 (N_13796,N_13209,N_13416);
nor U13797 (N_13797,N_13335,N_13421);
nor U13798 (N_13798,N_13260,N_13253);
nor U13799 (N_13799,N_13477,N_13436);
and U13800 (N_13800,N_13692,N_13736);
xnor U13801 (N_13801,N_13639,N_13771);
and U13802 (N_13802,N_13636,N_13670);
nand U13803 (N_13803,N_13594,N_13596);
nor U13804 (N_13804,N_13511,N_13703);
nor U13805 (N_13805,N_13529,N_13524);
nand U13806 (N_13806,N_13651,N_13604);
xor U13807 (N_13807,N_13548,N_13641);
xor U13808 (N_13808,N_13740,N_13502);
or U13809 (N_13809,N_13514,N_13583);
nor U13810 (N_13810,N_13522,N_13676);
nor U13811 (N_13811,N_13645,N_13743);
or U13812 (N_13812,N_13684,N_13680);
xnor U13813 (N_13813,N_13669,N_13735);
or U13814 (N_13814,N_13555,N_13565);
nand U13815 (N_13815,N_13712,N_13527);
nand U13816 (N_13816,N_13600,N_13500);
nand U13817 (N_13817,N_13616,N_13661);
and U13818 (N_13818,N_13628,N_13697);
xor U13819 (N_13819,N_13586,N_13612);
or U13820 (N_13820,N_13722,N_13662);
and U13821 (N_13821,N_13578,N_13655);
nand U13822 (N_13822,N_13775,N_13768);
or U13823 (N_13823,N_13672,N_13696);
or U13824 (N_13824,N_13531,N_13598);
and U13825 (N_13825,N_13741,N_13799);
nand U13826 (N_13826,N_13691,N_13790);
nor U13827 (N_13827,N_13738,N_13556);
and U13828 (N_13828,N_13552,N_13631);
or U13829 (N_13829,N_13613,N_13789);
nor U13830 (N_13830,N_13558,N_13732);
nor U13831 (N_13831,N_13719,N_13751);
xnor U13832 (N_13832,N_13637,N_13601);
or U13833 (N_13833,N_13623,N_13709);
or U13834 (N_13834,N_13593,N_13671);
and U13835 (N_13835,N_13777,N_13678);
nor U13836 (N_13836,N_13614,N_13758);
and U13837 (N_13837,N_13528,N_13649);
nor U13838 (N_13838,N_13507,N_13615);
nand U13839 (N_13839,N_13650,N_13508);
xnor U13840 (N_13840,N_13513,N_13699);
nor U13841 (N_13841,N_13674,N_13536);
nand U13842 (N_13842,N_13749,N_13792);
or U13843 (N_13843,N_13647,N_13668);
nor U13844 (N_13844,N_13549,N_13546);
or U13845 (N_13845,N_13626,N_13695);
nand U13846 (N_13846,N_13505,N_13515);
nand U13847 (N_13847,N_13659,N_13609);
nand U13848 (N_13848,N_13664,N_13787);
xor U13849 (N_13849,N_13657,N_13525);
nand U13850 (N_13850,N_13763,N_13690);
or U13851 (N_13851,N_13731,N_13627);
and U13852 (N_13852,N_13724,N_13520);
or U13853 (N_13853,N_13591,N_13617);
xor U13854 (N_13854,N_13764,N_13534);
xor U13855 (N_13855,N_13605,N_13791);
and U13856 (N_13856,N_13660,N_13750);
and U13857 (N_13857,N_13715,N_13711);
xnor U13858 (N_13858,N_13747,N_13761);
or U13859 (N_13859,N_13642,N_13510);
xor U13860 (N_13860,N_13793,N_13726);
nor U13861 (N_13861,N_13652,N_13550);
and U13862 (N_13862,N_13501,N_13648);
nand U13863 (N_13863,N_13778,N_13506);
nand U13864 (N_13864,N_13559,N_13653);
and U13865 (N_13865,N_13767,N_13533);
xor U13866 (N_13866,N_13752,N_13599);
nor U13867 (N_13867,N_13720,N_13638);
and U13868 (N_13868,N_13770,N_13545);
nor U13869 (N_13869,N_13710,N_13579);
nand U13870 (N_13870,N_13602,N_13694);
xnor U13871 (N_13871,N_13585,N_13728);
nor U13872 (N_13872,N_13630,N_13713);
or U13873 (N_13873,N_13781,N_13721);
nor U13874 (N_13874,N_13759,N_13798);
nor U13875 (N_13875,N_13526,N_13519);
xor U13876 (N_13876,N_13788,N_13568);
nand U13877 (N_13877,N_13704,N_13667);
and U13878 (N_13878,N_13621,N_13797);
nor U13879 (N_13879,N_13622,N_13733);
nor U13880 (N_13880,N_13608,N_13683);
nand U13881 (N_13881,N_13716,N_13517);
and U13882 (N_13882,N_13682,N_13698);
nand U13883 (N_13883,N_13581,N_13574);
and U13884 (N_13884,N_13625,N_13705);
and U13885 (N_13885,N_13737,N_13765);
nand U13886 (N_13886,N_13576,N_13782);
nor U13887 (N_13887,N_13706,N_13512);
nand U13888 (N_13888,N_13756,N_13665);
nor U13889 (N_13889,N_13532,N_13727);
or U13890 (N_13890,N_13656,N_13755);
xnor U13891 (N_13891,N_13634,N_13553);
xnor U13892 (N_13892,N_13557,N_13739);
nor U13893 (N_13893,N_13772,N_13685);
nor U13894 (N_13894,N_13701,N_13624);
or U13895 (N_13895,N_13589,N_13729);
xor U13896 (N_13896,N_13688,N_13644);
xor U13897 (N_13897,N_13780,N_13539);
or U13898 (N_13898,N_13643,N_13730);
or U13899 (N_13899,N_13551,N_13746);
xnor U13900 (N_13900,N_13795,N_13663);
or U13901 (N_13901,N_13745,N_13542);
and U13902 (N_13902,N_13566,N_13714);
nand U13903 (N_13903,N_13783,N_13689);
and U13904 (N_13904,N_13571,N_13588);
or U13905 (N_13905,N_13646,N_13618);
nand U13906 (N_13906,N_13597,N_13516);
and U13907 (N_13907,N_13734,N_13773);
and U13908 (N_13908,N_13521,N_13776);
nand U13909 (N_13909,N_13580,N_13707);
and U13910 (N_13910,N_13769,N_13504);
and U13911 (N_13911,N_13547,N_13666);
nand U13912 (N_13912,N_13717,N_13658);
and U13913 (N_13913,N_13779,N_13561);
nand U13914 (N_13914,N_13748,N_13744);
nand U13915 (N_13915,N_13774,N_13753);
and U13916 (N_13916,N_13702,N_13560);
nor U13917 (N_13917,N_13693,N_13562);
xnor U13918 (N_13918,N_13754,N_13723);
nor U13919 (N_13919,N_13619,N_13687);
or U13920 (N_13920,N_13530,N_13592);
or U13921 (N_13921,N_13794,N_13607);
or U13922 (N_13922,N_13785,N_13718);
or U13923 (N_13923,N_13544,N_13606);
or U13924 (N_13924,N_13575,N_13503);
nor U13925 (N_13925,N_13543,N_13603);
nor U13926 (N_13926,N_13677,N_13675);
or U13927 (N_13927,N_13632,N_13654);
or U13928 (N_13928,N_13595,N_13541);
and U13929 (N_13929,N_13620,N_13766);
nand U13930 (N_13930,N_13563,N_13635);
nor U13931 (N_13931,N_13610,N_13582);
and U13932 (N_13932,N_13518,N_13784);
xor U13933 (N_13933,N_13577,N_13564);
nand U13934 (N_13934,N_13786,N_13537);
and U13935 (N_13935,N_13569,N_13629);
nor U13936 (N_13936,N_13673,N_13640);
nor U13937 (N_13937,N_13572,N_13573);
nor U13938 (N_13938,N_13587,N_13757);
and U13939 (N_13939,N_13509,N_13760);
and U13940 (N_13940,N_13681,N_13742);
and U13941 (N_13941,N_13700,N_13590);
and U13942 (N_13942,N_13535,N_13554);
and U13943 (N_13943,N_13679,N_13762);
or U13944 (N_13944,N_13584,N_13633);
nor U13945 (N_13945,N_13540,N_13570);
xor U13946 (N_13946,N_13567,N_13686);
nor U13947 (N_13947,N_13708,N_13796);
and U13948 (N_13948,N_13538,N_13611);
and U13949 (N_13949,N_13725,N_13523);
and U13950 (N_13950,N_13593,N_13703);
xor U13951 (N_13951,N_13626,N_13703);
and U13952 (N_13952,N_13635,N_13706);
or U13953 (N_13953,N_13538,N_13532);
nand U13954 (N_13954,N_13714,N_13666);
nor U13955 (N_13955,N_13520,N_13690);
nor U13956 (N_13956,N_13714,N_13573);
or U13957 (N_13957,N_13675,N_13783);
xnor U13958 (N_13958,N_13700,N_13520);
nand U13959 (N_13959,N_13696,N_13622);
xnor U13960 (N_13960,N_13687,N_13639);
xnor U13961 (N_13961,N_13595,N_13733);
or U13962 (N_13962,N_13505,N_13672);
nand U13963 (N_13963,N_13700,N_13515);
and U13964 (N_13964,N_13612,N_13537);
or U13965 (N_13965,N_13775,N_13549);
or U13966 (N_13966,N_13729,N_13524);
xor U13967 (N_13967,N_13739,N_13697);
nand U13968 (N_13968,N_13779,N_13508);
or U13969 (N_13969,N_13799,N_13647);
xor U13970 (N_13970,N_13771,N_13743);
or U13971 (N_13971,N_13653,N_13580);
xor U13972 (N_13972,N_13757,N_13657);
xor U13973 (N_13973,N_13512,N_13597);
nand U13974 (N_13974,N_13797,N_13796);
and U13975 (N_13975,N_13775,N_13789);
nor U13976 (N_13976,N_13751,N_13709);
nor U13977 (N_13977,N_13577,N_13753);
nand U13978 (N_13978,N_13763,N_13781);
nand U13979 (N_13979,N_13679,N_13500);
xnor U13980 (N_13980,N_13734,N_13605);
or U13981 (N_13981,N_13654,N_13506);
xor U13982 (N_13982,N_13613,N_13544);
nand U13983 (N_13983,N_13722,N_13734);
xor U13984 (N_13984,N_13552,N_13744);
xor U13985 (N_13985,N_13702,N_13672);
or U13986 (N_13986,N_13614,N_13784);
or U13987 (N_13987,N_13754,N_13717);
xnor U13988 (N_13988,N_13553,N_13740);
or U13989 (N_13989,N_13697,N_13680);
xnor U13990 (N_13990,N_13674,N_13762);
nor U13991 (N_13991,N_13640,N_13515);
and U13992 (N_13992,N_13742,N_13791);
nand U13993 (N_13993,N_13618,N_13753);
and U13994 (N_13994,N_13597,N_13588);
nand U13995 (N_13995,N_13692,N_13748);
nand U13996 (N_13996,N_13529,N_13613);
nand U13997 (N_13997,N_13642,N_13519);
nand U13998 (N_13998,N_13564,N_13575);
nor U13999 (N_13999,N_13660,N_13531);
xnor U14000 (N_14000,N_13763,N_13641);
nand U14001 (N_14001,N_13566,N_13584);
xor U14002 (N_14002,N_13625,N_13511);
nand U14003 (N_14003,N_13572,N_13691);
and U14004 (N_14004,N_13506,N_13509);
xnor U14005 (N_14005,N_13637,N_13554);
nand U14006 (N_14006,N_13566,N_13530);
nand U14007 (N_14007,N_13659,N_13587);
nor U14008 (N_14008,N_13586,N_13516);
nand U14009 (N_14009,N_13742,N_13712);
and U14010 (N_14010,N_13580,N_13619);
and U14011 (N_14011,N_13786,N_13793);
nand U14012 (N_14012,N_13793,N_13510);
or U14013 (N_14013,N_13729,N_13713);
nand U14014 (N_14014,N_13798,N_13569);
nor U14015 (N_14015,N_13788,N_13618);
and U14016 (N_14016,N_13677,N_13561);
or U14017 (N_14017,N_13716,N_13518);
nor U14018 (N_14018,N_13650,N_13560);
nor U14019 (N_14019,N_13619,N_13793);
and U14020 (N_14020,N_13565,N_13543);
nor U14021 (N_14021,N_13526,N_13520);
nor U14022 (N_14022,N_13520,N_13628);
and U14023 (N_14023,N_13667,N_13581);
and U14024 (N_14024,N_13601,N_13530);
nor U14025 (N_14025,N_13730,N_13526);
or U14026 (N_14026,N_13577,N_13529);
and U14027 (N_14027,N_13607,N_13640);
or U14028 (N_14028,N_13677,N_13686);
or U14029 (N_14029,N_13661,N_13781);
nand U14030 (N_14030,N_13583,N_13711);
xnor U14031 (N_14031,N_13684,N_13730);
or U14032 (N_14032,N_13529,N_13770);
nor U14033 (N_14033,N_13516,N_13517);
nand U14034 (N_14034,N_13617,N_13729);
and U14035 (N_14035,N_13783,N_13716);
nor U14036 (N_14036,N_13772,N_13559);
nor U14037 (N_14037,N_13636,N_13573);
xnor U14038 (N_14038,N_13573,N_13677);
nand U14039 (N_14039,N_13553,N_13617);
and U14040 (N_14040,N_13594,N_13578);
nor U14041 (N_14041,N_13721,N_13664);
nand U14042 (N_14042,N_13657,N_13679);
nand U14043 (N_14043,N_13635,N_13551);
xnor U14044 (N_14044,N_13771,N_13530);
nor U14045 (N_14045,N_13626,N_13596);
nand U14046 (N_14046,N_13559,N_13591);
nand U14047 (N_14047,N_13698,N_13706);
nand U14048 (N_14048,N_13692,N_13540);
nor U14049 (N_14049,N_13513,N_13725);
and U14050 (N_14050,N_13539,N_13509);
or U14051 (N_14051,N_13574,N_13762);
or U14052 (N_14052,N_13703,N_13698);
and U14053 (N_14053,N_13555,N_13596);
nor U14054 (N_14054,N_13593,N_13625);
or U14055 (N_14055,N_13692,N_13772);
xor U14056 (N_14056,N_13760,N_13516);
nor U14057 (N_14057,N_13761,N_13652);
nor U14058 (N_14058,N_13521,N_13698);
or U14059 (N_14059,N_13643,N_13792);
nor U14060 (N_14060,N_13692,N_13728);
nor U14061 (N_14061,N_13707,N_13570);
or U14062 (N_14062,N_13643,N_13634);
xor U14063 (N_14063,N_13754,N_13627);
nor U14064 (N_14064,N_13567,N_13602);
nor U14065 (N_14065,N_13720,N_13767);
and U14066 (N_14066,N_13727,N_13652);
or U14067 (N_14067,N_13773,N_13650);
nor U14068 (N_14068,N_13608,N_13782);
nand U14069 (N_14069,N_13514,N_13758);
nand U14070 (N_14070,N_13740,N_13526);
or U14071 (N_14071,N_13635,N_13523);
or U14072 (N_14072,N_13507,N_13605);
or U14073 (N_14073,N_13508,N_13539);
or U14074 (N_14074,N_13625,N_13744);
and U14075 (N_14075,N_13758,N_13607);
nand U14076 (N_14076,N_13723,N_13534);
nor U14077 (N_14077,N_13616,N_13573);
and U14078 (N_14078,N_13534,N_13779);
nand U14079 (N_14079,N_13649,N_13667);
xnor U14080 (N_14080,N_13643,N_13517);
or U14081 (N_14081,N_13610,N_13502);
xor U14082 (N_14082,N_13576,N_13622);
or U14083 (N_14083,N_13776,N_13606);
nor U14084 (N_14084,N_13748,N_13746);
or U14085 (N_14085,N_13685,N_13655);
nor U14086 (N_14086,N_13639,N_13596);
xor U14087 (N_14087,N_13696,N_13754);
and U14088 (N_14088,N_13541,N_13725);
xor U14089 (N_14089,N_13522,N_13702);
xnor U14090 (N_14090,N_13637,N_13593);
xor U14091 (N_14091,N_13605,N_13515);
and U14092 (N_14092,N_13690,N_13776);
xnor U14093 (N_14093,N_13795,N_13780);
and U14094 (N_14094,N_13532,N_13621);
nor U14095 (N_14095,N_13540,N_13589);
nor U14096 (N_14096,N_13785,N_13585);
and U14097 (N_14097,N_13681,N_13617);
nor U14098 (N_14098,N_13694,N_13563);
nor U14099 (N_14099,N_13568,N_13515);
nand U14100 (N_14100,N_13948,N_14047);
nand U14101 (N_14101,N_13967,N_13894);
and U14102 (N_14102,N_13842,N_14017);
xor U14103 (N_14103,N_13964,N_13959);
nor U14104 (N_14104,N_14070,N_14037);
and U14105 (N_14105,N_14065,N_13830);
and U14106 (N_14106,N_13804,N_13923);
nand U14107 (N_14107,N_13871,N_13810);
xor U14108 (N_14108,N_13997,N_14095);
nand U14109 (N_14109,N_13926,N_13819);
nand U14110 (N_14110,N_13867,N_14078);
or U14111 (N_14111,N_13850,N_14056);
and U14112 (N_14112,N_13902,N_14052);
and U14113 (N_14113,N_14024,N_13825);
xor U14114 (N_14114,N_13972,N_13837);
xnor U14115 (N_14115,N_13855,N_13803);
or U14116 (N_14116,N_13878,N_14021);
or U14117 (N_14117,N_13900,N_13989);
nand U14118 (N_14118,N_13932,N_14075);
xor U14119 (N_14119,N_13838,N_13991);
xor U14120 (N_14120,N_13915,N_13857);
and U14121 (N_14121,N_13962,N_13927);
xor U14122 (N_14122,N_13879,N_14002);
nor U14123 (N_14123,N_13899,N_13998);
nand U14124 (N_14124,N_13916,N_13924);
nor U14125 (N_14125,N_13884,N_13917);
and U14126 (N_14126,N_13977,N_13937);
or U14127 (N_14127,N_13890,N_13930);
nand U14128 (N_14128,N_14081,N_14044);
nor U14129 (N_14129,N_14043,N_13911);
nor U14130 (N_14130,N_13844,N_13860);
and U14131 (N_14131,N_13816,N_14060);
nor U14132 (N_14132,N_13986,N_14040);
or U14133 (N_14133,N_13812,N_13841);
nor U14134 (N_14134,N_13935,N_13958);
xor U14135 (N_14135,N_13815,N_13995);
xnor U14136 (N_14136,N_14091,N_13897);
xor U14137 (N_14137,N_13843,N_13978);
nor U14138 (N_14138,N_13808,N_13827);
nand U14139 (N_14139,N_13955,N_14059);
xnor U14140 (N_14140,N_13851,N_13934);
xor U14141 (N_14141,N_13954,N_13829);
nor U14142 (N_14142,N_13875,N_13903);
and U14143 (N_14143,N_14036,N_14085);
nor U14144 (N_14144,N_14099,N_13859);
xnor U14145 (N_14145,N_13912,N_13922);
nor U14146 (N_14146,N_14010,N_13858);
nand U14147 (N_14147,N_13946,N_13814);
xor U14148 (N_14148,N_13953,N_13872);
xor U14149 (N_14149,N_14022,N_13846);
and U14150 (N_14150,N_14098,N_13870);
or U14151 (N_14151,N_14003,N_13869);
or U14152 (N_14152,N_13945,N_13887);
xnor U14153 (N_14153,N_13951,N_13913);
or U14154 (N_14154,N_13863,N_13847);
nand U14155 (N_14155,N_13982,N_14009);
and U14156 (N_14156,N_13833,N_14079);
xor U14157 (N_14157,N_14026,N_13940);
nand U14158 (N_14158,N_13892,N_13906);
xnor U14159 (N_14159,N_13936,N_14058);
and U14160 (N_14160,N_14086,N_14093);
xnor U14161 (N_14161,N_13888,N_14082);
and U14162 (N_14162,N_13952,N_13868);
nand U14163 (N_14163,N_13919,N_14004);
nor U14164 (N_14164,N_13966,N_13832);
or U14165 (N_14165,N_14030,N_13993);
or U14166 (N_14166,N_14051,N_14072);
or U14167 (N_14167,N_14066,N_13933);
or U14168 (N_14168,N_13885,N_13968);
xor U14169 (N_14169,N_14050,N_14028);
xnor U14170 (N_14170,N_13985,N_13987);
xnor U14171 (N_14171,N_14013,N_14031);
nor U14172 (N_14172,N_13811,N_14008);
nor U14173 (N_14173,N_13957,N_13961);
nand U14174 (N_14174,N_13802,N_13981);
or U14175 (N_14175,N_14006,N_13990);
or U14176 (N_14176,N_14011,N_14048);
and U14177 (N_14177,N_14007,N_14020);
or U14178 (N_14178,N_13918,N_14094);
xnor U14179 (N_14179,N_13914,N_13910);
or U14180 (N_14180,N_13891,N_13874);
nand U14181 (N_14181,N_13896,N_14063);
xor U14182 (N_14182,N_13849,N_14083);
or U14183 (N_14183,N_13820,N_13988);
or U14184 (N_14184,N_14067,N_13974);
nor U14185 (N_14185,N_13980,N_13960);
or U14186 (N_14186,N_13928,N_14023);
or U14187 (N_14187,N_14087,N_13862);
and U14188 (N_14188,N_13886,N_13999);
nor U14189 (N_14189,N_13949,N_13800);
nand U14190 (N_14190,N_14025,N_14016);
and U14191 (N_14191,N_13823,N_13876);
nand U14192 (N_14192,N_14038,N_13809);
xnor U14193 (N_14193,N_14071,N_13861);
xnor U14194 (N_14194,N_14064,N_13921);
and U14195 (N_14195,N_13947,N_13853);
xnor U14196 (N_14196,N_14062,N_14033);
or U14197 (N_14197,N_14074,N_13941);
or U14198 (N_14198,N_14045,N_13856);
and U14199 (N_14199,N_13983,N_14053);
xnor U14200 (N_14200,N_13965,N_13956);
xor U14201 (N_14201,N_14034,N_13822);
or U14202 (N_14202,N_14001,N_14029);
nand U14203 (N_14203,N_13938,N_13866);
nand U14204 (N_14204,N_13994,N_14057);
xor U14205 (N_14205,N_14019,N_13865);
xnor U14206 (N_14206,N_14097,N_14073);
or U14207 (N_14207,N_13801,N_13817);
nand U14208 (N_14208,N_14032,N_13831);
or U14209 (N_14209,N_14080,N_14068);
nand U14210 (N_14210,N_14089,N_13824);
nor U14211 (N_14211,N_13805,N_13909);
nand U14212 (N_14212,N_14014,N_13939);
or U14213 (N_14213,N_13979,N_13854);
or U14214 (N_14214,N_14046,N_14039);
and U14215 (N_14215,N_14042,N_13828);
nor U14216 (N_14216,N_13806,N_13904);
or U14217 (N_14217,N_14076,N_13845);
and U14218 (N_14218,N_13996,N_13807);
or U14219 (N_14219,N_13834,N_14088);
or U14220 (N_14220,N_13840,N_13852);
nor U14221 (N_14221,N_13839,N_14054);
xor U14222 (N_14222,N_14035,N_14012);
nand U14223 (N_14223,N_13929,N_13908);
nand U14224 (N_14224,N_13898,N_13835);
and U14225 (N_14225,N_13905,N_14092);
nor U14226 (N_14226,N_13907,N_14027);
or U14227 (N_14227,N_13942,N_13848);
and U14228 (N_14228,N_13901,N_13893);
nand U14229 (N_14229,N_13973,N_14077);
and U14230 (N_14230,N_13943,N_13826);
xnor U14231 (N_14231,N_13920,N_14084);
and U14232 (N_14232,N_13895,N_13873);
nor U14233 (N_14233,N_13883,N_14069);
nor U14234 (N_14234,N_13975,N_14005);
nor U14235 (N_14235,N_14000,N_13950);
xnor U14236 (N_14236,N_13992,N_13925);
or U14237 (N_14237,N_13984,N_13970);
nand U14238 (N_14238,N_13864,N_13944);
nor U14239 (N_14239,N_13931,N_13881);
and U14240 (N_14240,N_14041,N_14015);
xnor U14241 (N_14241,N_14090,N_14049);
nor U14242 (N_14242,N_13969,N_13889);
or U14243 (N_14243,N_13818,N_13836);
xnor U14244 (N_14244,N_14055,N_14061);
nor U14245 (N_14245,N_13963,N_13976);
xnor U14246 (N_14246,N_13821,N_13813);
xor U14247 (N_14247,N_14096,N_14018);
nor U14248 (N_14248,N_13971,N_13877);
and U14249 (N_14249,N_13880,N_13882);
nand U14250 (N_14250,N_14002,N_14021);
and U14251 (N_14251,N_14069,N_13977);
and U14252 (N_14252,N_13939,N_13841);
or U14253 (N_14253,N_14088,N_13958);
and U14254 (N_14254,N_14070,N_14064);
nand U14255 (N_14255,N_13822,N_14030);
nor U14256 (N_14256,N_13914,N_13947);
nor U14257 (N_14257,N_13850,N_14074);
xor U14258 (N_14258,N_14052,N_13998);
or U14259 (N_14259,N_14069,N_13947);
xor U14260 (N_14260,N_13873,N_14038);
nand U14261 (N_14261,N_13930,N_14029);
nor U14262 (N_14262,N_13919,N_13828);
nor U14263 (N_14263,N_14069,N_14000);
or U14264 (N_14264,N_14003,N_13831);
nor U14265 (N_14265,N_13830,N_14061);
and U14266 (N_14266,N_13839,N_14090);
and U14267 (N_14267,N_13852,N_13814);
or U14268 (N_14268,N_13887,N_13930);
or U14269 (N_14269,N_13825,N_13977);
nor U14270 (N_14270,N_13890,N_14018);
xnor U14271 (N_14271,N_13904,N_13858);
or U14272 (N_14272,N_13952,N_13813);
xor U14273 (N_14273,N_14015,N_14054);
and U14274 (N_14274,N_14067,N_13973);
nand U14275 (N_14275,N_13920,N_14058);
nand U14276 (N_14276,N_13901,N_13924);
nand U14277 (N_14277,N_13957,N_14093);
or U14278 (N_14278,N_13881,N_13917);
nor U14279 (N_14279,N_13964,N_13855);
and U14280 (N_14280,N_13899,N_14082);
nor U14281 (N_14281,N_13863,N_13843);
nand U14282 (N_14282,N_13943,N_13976);
and U14283 (N_14283,N_13967,N_14065);
nor U14284 (N_14284,N_13934,N_13842);
and U14285 (N_14285,N_13881,N_13871);
nand U14286 (N_14286,N_14062,N_13877);
or U14287 (N_14287,N_14020,N_13973);
and U14288 (N_14288,N_13847,N_13893);
xnor U14289 (N_14289,N_13961,N_14010);
nor U14290 (N_14290,N_14073,N_13946);
nor U14291 (N_14291,N_13839,N_13911);
nand U14292 (N_14292,N_13812,N_13888);
and U14293 (N_14293,N_14045,N_13957);
nand U14294 (N_14294,N_13803,N_13817);
or U14295 (N_14295,N_13980,N_13818);
nand U14296 (N_14296,N_13973,N_13863);
nand U14297 (N_14297,N_13877,N_13992);
or U14298 (N_14298,N_14089,N_13833);
nor U14299 (N_14299,N_13918,N_13922);
or U14300 (N_14300,N_13904,N_14007);
and U14301 (N_14301,N_14015,N_13894);
and U14302 (N_14302,N_13876,N_13846);
xor U14303 (N_14303,N_14087,N_14019);
nand U14304 (N_14304,N_13909,N_13871);
or U14305 (N_14305,N_13965,N_13863);
nand U14306 (N_14306,N_14051,N_13860);
and U14307 (N_14307,N_13941,N_13944);
xnor U14308 (N_14308,N_13892,N_14044);
nor U14309 (N_14309,N_13917,N_13821);
xor U14310 (N_14310,N_13947,N_13966);
or U14311 (N_14311,N_13930,N_14038);
nor U14312 (N_14312,N_14078,N_13948);
nor U14313 (N_14313,N_13825,N_13815);
nor U14314 (N_14314,N_14036,N_13974);
or U14315 (N_14315,N_14018,N_13922);
xnor U14316 (N_14316,N_14051,N_13869);
or U14317 (N_14317,N_13821,N_13865);
nand U14318 (N_14318,N_13948,N_14091);
xnor U14319 (N_14319,N_14042,N_13831);
nor U14320 (N_14320,N_13843,N_13891);
and U14321 (N_14321,N_14037,N_13900);
nor U14322 (N_14322,N_13921,N_13938);
xnor U14323 (N_14323,N_13877,N_13985);
xor U14324 (N_14324,N_13962,N_13832);
nor U14325 (N_14325,N_13838,N_13873);
nor U14326 (N_14326,N_13960,N_13925);
or U14327 (N_14327,N_13868,N_13910);
xor U14328 (N_14328,N_13933,N_14011);
or U14329 (N_14329,N_14055,N_13989);
or U14330 (N_14330,N_13913,N_14070);
or U14331 (N_14331,N_14012,N_14056);
nand U14332 (N_14332,N_13873,N_13812);
or U14333 (N_14333,N_13820,N_14064);
or U14334 (N_14334,N_13949,N_13968);
nor U14335 (N_14335,N_13845,N_14028);
nor U14336 (N_14336,N_14002,N_13949);
xor U14337 (N_14337,N_13970,N_14022);
nand U14338 (N_14338,N_14013,N_14081);
or U14339 (N_14339,N_14035,N_14027);
and U14340 (N_14340,N_13822,N_14061);
nor U14341 (N_14341,N_14092,N_13888);
and U14342 (N_14342,N_14076,N_13901);
and U14343 (N_14343,N_13913,N_13864);
xor U14344 (N_14344,N_13808,N_13982);
and U14345 (N_14345,N_13871,N_13882);
xor U14346 (N_14346,N_13974,N_13963);
nand U14347 (N_14347,N_14059,N_13868);
xnor U14348 (N_14348,N_14007,N_13841);
or U14349 (N_14349,N_13843,N_14060);
and U14350 (N_14350,N_13930,N_13994);
and U14351 (N_14351,N_13870,N_13900);
nor U14352 (N_14352,N_14024,N_13900);
nand U14353 (N_14353,N_13863,N_13813);
or U14354 (N_14354,N_14012,N_14010);
and U14355 (N_14355,N_14087,N_13951);
or U14356 (N_14356,N_14040,N_13987);
or U14357 (N_14357,N_13811,N_14038);
nor U14358 (N_14358,N_14078,N_13817);
nand U14359 (N_14359,N_13967,N_13858);
nor U14360 (N_14360,N_14085,N_14082);
nand U14361 (N_14361,N_13957,N_13863);
and U14362 (N_14362,N_14039,N_13891);
xor U14363 (N_14363,N_14079,N_13869);
and U14364 (N_14364,N_13891,N_14090);
xor U14365 (N_14365,N_13870,N_13840);
or U14366 (N_14366,N_13899,N_14044);
or U14367 (N_14367,N_14022,N_14012);
and U14368 (N_14368,N_13917,N_14080);
or U14369 (N_14369,N_13878,N_13973);
and U14370 (N_14370,N_14064,N_13985);
xor U14371 (N_14371,N_14099,N_13837);
nand U14372 (N_14372,N_13855,N_13853);
and U14373 (N_14373,N_13881,N_14076);
xor U14374 (N_14374,N_13803,N_14096);
and U14375 (N_14375,N_13908,N_13966);
nor U14376 (N_14376,N_14059,N_14035);
or U14377 (N_14377,N_13802,N_13887);
or U14378 (N_14378,N_14010,N_13977);
or U14379 (N_14379,N_14046,N_14096);
and U14380 (N_14380,N_14017,N_13921);
nor U14381 (N_14381,N_14089,N_13973);
or U14382 (N_14382,N_14009,N_13995);
nand U14383 (N_14383,N_13923,N_13999);
or U14384 (N_14384,N_14001,N_13823);
nor U14385 (N_14385,N_13804,N_14043);
nor U14386 (N_14386,N_13921,N_13908);
and U14387 (N_14387,N_13915,N_14078);
and U14388 (N_14388,N_13953,N_14096);
or U14389 (N_14389,N_13813,N_13907);
xnor U14390 (N_14390,N_14069,N_14023);
nand U14391 (N_14391,N_14061,N_13881);
nor U14392 (N_14392,N_13943,N_13811);
nor U14393 (N_14393,N_13821,N_13814);
or U14394 (N_14394,N_14034,N_14013);
nor U14395 (N_14395,N_13903,N_13850);
nor U14396 (N_14396,N_14062,N_14073);
nand U14397 (N_14397,N_13901,N_14035);
and U14398 (N_14398,N_14067,N_14066);
or U14399 (N_14399,N_13820,N_13979);
nand U14400 (N_14400,N_14374,N_14302);
or U14401 (N_14401,N_14313,N_14394);
xor U14402 (N_14402,N_14327,N_14399);
nor U14403 (N_14403,N_14289,N_14259);
nor U14404 (N_14404,N_14128,N_14255);
and U14405 (N_14405,N_14326,N_14323);
and U14406 (N_14406,N_14395,N_14160);
and U14407 (N_14407,N_14359,N_14219);
xor U14408 (N_14408,N_14251,N_14239);
and U14409 (N_14409,N_14362,N_14348);
or U14410 (N_14410,N_14354,N_14306);
xnor U14411 (N_14411,N_14349,N_14281);
nand U14412 (N_14412,N_14310,N_14233);
nor U14413 (N_14413,N_14120,N_14378);
or U14414 (N_14414,N_14163,N_14198);
nand U14415 (N_14415,N_14110,N_14262);
xnor U14416 (N_14416,N_14147,N_14333);
nor U14417 (N_14417,N_14383,N_14246);
or U14418 (N_14418,N_14142,N_14154);
nor U14419 (N_14419,N_14254,N_14318);
or U14420 (N_14420,N_14125,N_14155);
nand U14421 (N_14421,N_14191,N_14340);
nand U14422 (N_14422,N_14182,N_14269);
nor U14423 (N_14423,N_14353,N_14217);
xnor U14424 (N_14424,N_14307,N_14238);
and U14425 (N_14425,N_14250,N_14207);
xor U14426 (N_14426,N_14371,N_14339);
and U14427 (N_14427,N_14369,N_14242);
or U14428 (N_14428,N_14391,N_14235);
xnor U14429 (N_14429,N_14351,N_14230);
nand U14430 (N_14430,N_14277,N_14256);
and U14431 (N_14431,N_14122,N_14266);
and U14432 (N_14432,N_14267,N_14180);
and U14433 (N_14433,N_14222,N_14196);
or U14434 (N_14434,N_14271,N_14335);
nor U14435 (N_14435,N_14317,N_14344);
nor U14436 (N_14436,N_14216,N_14261);
or U14437 (N_14437,N_14388,N_14106);
nor U14438 (N_14438,N_14153,N_14101);
and U14439 (N_14439,N_14345,N_14161);
nor U14440 (N_14440,N_14393,N_14260);
nand U14441 (N_14441,N_14370,N_14316);
nand U14442 (N_14442,N_14165,N_14293);
nand U14443 (N_14443,N_14325,N_14263);
and U14444 (N_14444,N_14305,N_14381);
nor U14445 (N_14445,N_14140,N_14249);
nand U14446 (N_14446,N_14214,N_14205);
nand U14447 (N_14447,N_14194,N_14361);
nand U14448 (N_14448,N_14272,N_14195);
nor U14449 (N_14449,N_14220,N_14279);
or U14450 (N_14450,N_14273,N_14121);
xnor U14451 (N_14451,N_14257,N_14276);
nand U14452 (N_14452,N_14150,N_14188);
or U14453 (N_14453,N_14108,N_14126);
and U14454 (N_14454,N_14319,N_14105);
nor U14455 (N_14455,N_14355,N_14295);
nand U14456 (N_14456,N_14303,N_14322);
or U14457 (N_14457,N_14146,N_14365);
or U14458 (N_14458,N_14236,N_14177);
or U14459 (N_14459,N_14173,N_14285);
nand U14460 (N_14460,N_14258,N_14223);
nand U14461 (N_14461,N_14336,N_14200);
or U14462 (N_14462,N_14226,N_14342);
or U14463 (N_14463,N_14385,N_14224);
xor U14464 (N_14464,N_14157,N_14159);
and U14465 (N_14465,N_14175,N_14286);
or U14466 (N_14466,N_14245,N_14347);
xor U14467 (N_14467,N_14169,N_14199);
or U14468 (N_14468,N_14145,N_14375);
and U14469 (N_14469,N_14275,N_14178);
or U14470 (N_14470,N_14185,N_14320);
or U14471 (N_14471,N_14297,N_14210);
xnor U14472 (N_14472,N_14117,N_14240);
xnor U14473 (N_14473,N_14171,N_14166);
nor U14474 (N_14474,N_14270,N_14193);
or U14475 (N_14475,N_14290,N_14184);
and U14476 (N_14476,N_14209,N_14232);
and U14477 (N_14477,N_14148,N_14283);
nor U14478 (N_14478,N_14301,N_14189);
or U14479 (N_14479,N_14156,N_14168);
and U14480 (N_14480,N_14139,N_14231);
nor U14481 (N_14481,N_14366,N_14127);
xnor U14482 (N_14482,N_14389,N_14206);
xnor U14483 (N_14483,N_14253,N_14215);
nor U14484 (N_14484,N_14364,N_14397);
nor U14485 (N_14485,N_14329,N_14321);
nor U14486 (N_14486,N_14292,N_14304);
nor U14487 (N_14487,N_14186,N_14387);
and U14488 (N_14488,N_14331,N_14134);
nor U14489 (N_14489,N_14268,N_14352);
or U14490 (N_14490,N_14109,N_14358);
and U14491 (N_14491,N_14234,N_14299);
and U14492 (N_14492,N_14225,N_14390);
and U14493 (N_14493,N_14386,N_14133);
xnor U14494 (N_14494,N_14131,N_14123);
nor U14495 (N_14495,N_14149,N_14204);
or U14496 (N_14496,N_14346,N_14213);
xor U14497 (N_14497,N_14172,N_14298);
nand U14498 (N_14498,N_14202,N_14158);
xnor U14499 (N_14499,N_14167,N_14384);
and U14500 (N_14500,N_14124,N_14228);
nor U14501 (N_14501,N_14192,N_14315);
nor U14502 (N_14502,N_14143,N_14137);
nand U14503 (N_14503,N_14328,N_14356);
xor U14504 (N_14504,N_14119,N_14201);
or U14505 (N_14505,N_14118,N_14382);
and U14506 (N_14506,N_14187,N_14392);
and U14507 (N_14507,N_14308,N_14132);
nand U14508 (N_14508,N_14265,N_14291);
or U14509 (N_14509,N_14114,N_14112);
nand U14510 (N_14510,N_14294,N_14115);
or U14511 (N_14511,N_14130,N_14288);
nor U14512 (N_14512,N_14376,N_14343);
nand U14513 (N_14513,N_14183,N_14312);
xor U14514 (N_14514,N_14176,N_14377);
nor U14515 (N_14515,N_14380,N_14247);
xnor U14516 (N_14516,N_14197,N_14311);
and U14517 (N_14517,N_14138,N_14373);
xor U14518 (N_14518,N_14170,N_14181);
nor U14519 (N_14519,N_14129,N_14179);
nor U14520 (N_14520,N_14284,N_14162);
nor U14521 (N_14521,N_14135,N_14107);
xnor U14522 (N_14522,N_14221,N_14372);
nor U14523 (N_14523,N_14244,N_14337);
and U14524 (N_14524,N_14264,N_14332);
nand U14525 (N_14525,N_14296,N_14237);
or U14526 (N_14526,N_14368,N_14309);
nor U14527 (N_14527,N_14252,N_14229);
and U14528 (N_14528,N_14104,N_14360);
nor U14529 (N_14529,N_14208,N_14100);
xnor U14530 (N_14530,N_14152,N_14330);
and U14531 (N_14531,N_14341,N_14227);
nand U14532 (N_14532,N_14203,N_14111);
nor U14533 (N_14533,N_14398,N_14103);
nand U14534 (N_14534,N_14280,N_14248);
nand U14535 (N_14535,N_14113,N_14190);
or U14536 (N_14536,N_14396,N_14274);
xnor U14537 (N_14537,N_14324,N_14363);
or U14538 (N_14538,N_14357,N_14212);
nor U14539 (N_14539,N_14300,N_14164);
xor U14540 (N_14540,N_14338,N_14282);
or U14541 (N_14541,N_14367,N_14136);
xnor U14542 (N_14542,N_14287,N_14116);
nor U14543 (N_14543,N_14218,N_14314);
and U14544 (N_14544,N_14151,N_14141);
and U14545 (N_14545,N_14144,N_14102);
or U14546 (N_14546,N_14174,N_14278);
or U14547 (N_14547,N_14243,N_14334);
nor U14548 (N_14548,N_14379,N_14241);
nor U14549 (N_14549,N_14350,N_14211);
xnor U14550 (N_14550,N_14309,N_14338);
nand U14551 (N_14551,N_14106,N_14297);
xnor U14552 (N_14552,N_14279,N_14118);
or U14553 (N_14553,N_14144,N_14168);
nand U14554 (N_14554,N_14255,N_14187);
or U14555 (N_14555,N_14122,N_14310);
nand U14556 (N_14556,N_14394,N_14249);
nand U14557 (N_14557,N_14371,N_14214);
or U14558 (N_14558,N_14187,N_14210);
nor U14559 (N_14559,N_14136,N_14272);
nand U14560 (N_14560,N_14113,N_14142);
or U14561 (N_14561,N_14186,N_14301);
xor U14562 (N_14562,N_14302,N_14387);
xor U14563 (N_14563,N_14367,N_14282);
and U14564 (N_14564,N_14281,N_14311);
or U14565 (N_14565,N_14100,N_14270);
nand U14566 (N_14566,N_14115,N_14141);
nor U14567 (N_14567,N_14247,N_14241);
or U14568 (N_14568,N_14295,N_14251);
nor U14569 (N_14569,N_14179,N_14203);
or U14570 (N_14570,N_14275,N_14223);
nand U14571 (N_14571,N_14312,N_14221);
xor U14572 (N_14572,N_14198,N_14322);
and U14573 (N_14573,N_14119,N_14272);
and U14574 (N_14574,N_14109,N_14284);
or U14575 (N_14575,N_14156,N_14305);
and U14576 (N_14576,N_14349,N_14231);
or U14577 (N_14577,N_14116,N_14181);
and U14578 (N_14578,N_14333,N_14358);
or U14579 (N_14579,N_14310,N_14170);
nor U14580 (N_14580,N_14117,N_14245);
or U14581 (N_14581,N_14133,N_14294);
or U14582 (N_14582,N_14177,N_14306);
xor U14583 (N_14583,N_14316,N_14247);
xnor U14584 (N_14584,N_14286,N_14221);
and U14585 (N_14585,N_14340,N_14106);
nand U14586 (N_14586,N_14276,N_14247);
and U14587 (N_14587,N_14360,N_14298);
or U14588 (N_14588,N_14164,N_14315);
xnor U14589 (N_14589,N_14378,N_14290);
nand U14590 (N_14590,N_14344,N_14225);
xor U14591 (N_14591,N_14126,N_14295);
or U14592 (N_14592,N_14346,N_14337);
or U14593 (N_14593,N_14327,N_14163);
and U14594 (N_14594,N_14321,N_14133);
nand U14595 (N_14595,N_14142,N_14229);
or U14596 (N_14596,N_14250,N_14204);
nor U14597 (N_14597,N_14397,N_14356);
nand U14598 (N_14598,N_14296,N_14183);
or U14599 (N_14599,N_14341,N_14136);
or U14600 (N_14600,N_14349,N_14211);
xnor U14601 (N_14601,N_14191,N_14377);
and U14602 (N_14602,N_14304,N_14393);
or U14603 (N_14603,N_14137,N_14144);
and U14604 (N_14604,N_14144,N_14187);
nand U14605 (N_14605,N_14105,N_14179);
or U14606 (N_14606,N_14258,N_14322);
nand U14607 (N_14607,N_14274,N_14251);
and U14608 (N_14608,N_14153,N_14217);
xnor U14609 (N_14609,N_14132,N_14307);
nor U14610 (N_14610,N_14359,N_14243);
nor U14611 (N_14611,N_14370,N_14381);
xor U14612 (N_14612,N_14210,N_14282);
xnor U14613 (N_14613,N_14232,N_14352);
or U14614 (N_14614,N_14332,N_14275);
and U14615 (N_14615,N_14225,N_14238);
or U14616 (N_14616,N_14340,N_14163);
or U14617 (N_14617,N_14278,N_14213);
or U14618 (N_14618,N_14189,N_14317);
and U14619 (N_14619,N_14160,N_14208);
and U14620 (N_14620,N_14369,N_14122);
and U14621 (N_14621,N_14267,N_14393);
nor U14622 (N_14622,N_14290,N_14216);
and U14623 (N_14623,N_14190,N_14225);
or U14624 (N_14624,N_14113,N_14256);
nand U14625 (N_14625,N_14255,N_14101);
and U14626 (N_14626,N_14390,N_14168);
and U14627 (N_14627,N_14285,N_14162);
nand U14628 (N_14628,N_14347,N_14171);
and U14629 (N_14629,N_14377,N_14217);
and U14630 (N_14630,N_14239,N_14147);
or U14631 (N_14631,N_14324,N_14260);
or U14632 (N_14632,N_14210,N_14260);
or U14633 (N_14633,N_14161,N_14351);
or U14634 (N_14634,N_14168,N_14110);
xnor U14635 (N_14635,N_14324,N_14140);
nand U14636 (N_14636,N_14228,N_14176);
xor U14637 (N_14637,N_14208,N_14167);
or U14638 (N_14638,N_14384,N_14158);
or U14639 (N_14639,N_14134,N_14393);
xor U14640 (N_14640,N_14165,N_14243);
and U14641 (N_14641,N_14278,N_14322);
nor U14642 (N_14642,N_14382,N_14398);
xnor U14643 (N_14643,N_14248,N_14225);
xor U14644 (N_14644,N_14339,N_14121);
nand U14645 (N_14645,N_14377,N_14366);
nor U14646 (N_14646,N_14367,N_14109);
and U14647 (N_14647,N_14323,N_14114);
nand U14648 (N_14648,N_14366,N_14309);
or U14649 (N_14649,N_14356,N_14181);
nor U14650 (N_14650,N_14116,N_14237);
and U14651 (N_14651,N_14167,N_14120);
and U14652 (N_14652,N_14263,N_14346);
nand U14653 (N_14653,N_14372,N_14367);
or U14654 (N_14654,N_14194,N_14205);
xnor U14655 (N_14655,N_14299,N_14269);
or U14656 (N_14656,N_14394,N_14381);
or U14657 (N_14657,N_14276,N_14303);
and U14658 (N_14658,N_14392,N_14330);
xor U14659 (N_14659,N_14199,N_14175);
nand U14660 (N_14660,N_14152,N_14393);
nand U14661 (N_14661,N_14308,N_14323);
nand U14662 (N_14662,N_14324,N_14361);
and U14663 (N_14663,N_14237,N_14139);
xnor U14664 (N_14664,N_14184,N_14102);
xor U14665 (N_14665,N_14187,N_14361);
or U14666 (N_14666,N_14291,N_14290);
nor U14667 (N_14667,N_14307,N_14390);
nand U14668 (N_14668,N_14335,N_14382);
or U14669 (N_14669,N_14112,N_14262);
or U14670 (N_14670,N_14352,N_14144);
and U14671 (N_14671,N_14374,N_14390);
or U14672 (N_14672,N_14119,N_14231);
or U14673 (N_14673,N_14241,N_14314);
xnor U14674 (N_14674,N_14291,N_14280);
nand U14675 (N_14675,N_14232,N_14230);
nor U14676 (N_14676,N_14211,N_14163);
xor U14677 (N_14677,N_14103,N_14286);
and U14678 (N_14678,N_14311,N_14131);
nor U14679 (N_14679,N_14361,N_14146);
nor U14680 (N_14680,N_14194,N_14135);
nand U14681 (N_14681,N_14308,N_14377);
nand U14682 (N_14682,N_14321,N_14161);
nor U14683 (N_14683,N_14278,N_14292);
nand U14684 (N_14684,N_14252,N_14285);
nor U14685 (N_14685,N_14171,N_14320);
nand U14686 (N_14686,N_14192,N_14144);
or U14687 (N_14687,N_14320,N_14331);
nor U14688 (N_14688,N_14179,N_14209);
or U14689 (N_14689,N_14364,N_14385);
xnor U14690 (N_14690,N_14271,N_14210);
nor U14691 (N_14691,N_14181,N_14363);
and U14692 (N_14692,N_14229,N_14382);
nand U14693 (N_14693,N_14300,N_14185);
xor U14694 (N_14694,N_14307,N_14163);
or U14695 (N_14695,N_14278,N_14308);
nor U14696 (N_14696,N_14113,N_14246);
or U14697 (N_14697,N_14328,N_14269);
and U14698 (N_14698,N_14250,N_14373);
nor U14699 (N_14699,N_14102,N_14116);
nor U14700 (N_14700,N_14448,N_14595);
and U14701 (N_14701,N_14434,N_14651);
nand U14702 (N_14702,N_14517,N_14691);
and U14703 (N_14703,N_14426,N_14523);
nand U14704 (N_14704,N_14419,N_14462);
nand U14705 (N_14705,N_14473,N_14600);
and U14706 (N_14706,N_14458,N_14605);
xnor U14707 (N_14707,N_14487,N_14513);
nor U14708 (N_14708,N_14541,N_14597);
xnor U14709 (N_14709,N_14417,N_14413);
and U14710 (N_14710,N_14418,N_14657);
and U14711 (N_14711,N_14546,N_14670);
xnor U14712 (N_14712,N_14680,N_14437);
or U14713 (N_14713,N_14469,N_14669);
and U14714 (N_14714,N_14537,N_14624);
nor U14715 (N_14715,N_14536,N_14620);
xor U14716 (N_14716,N_14578,N_14555);
nor U14717 (N_14717,N_14671,N_14672);
and U14718 (N_14718,N_14539,N_14653);
or U14719 (N_14719,N_14443,N_14564);
nand U14720 (N_14720,N_14629,N_14580);
or U14721 (N_14721,N_14401,N_14614);
nor U14722 (N_14722,N_14404,N_14694);
xor U14723 (N_14723,N_14489,N_14545);
and U14724 (N_14724,N_14674,N_14442);
or U14725 (N_14725,N_14479,N_14526);
nor U14726 (N_14726,N_14444,N_14400);
nand U14727 (N_14727,N_14650,N_14529);
nor U14728 (N_14728,N_14409,N_14570);
and U14729 (N_14729,N_14515,N_14626);
nand U14730 (N_14730,N_14652,N_14408);
nand U14731 (N_14731,N_14505,N_14630);
xnor U14732 (N_14732,N_14598,N_14607);
or U14733 (N_14733,N_14538,N_14440);
and U14734 (N_14734,N_14682,N_14554);
nor U14735 (N_14735,N_14410,N_14456);
and U14736 (N_14736,N_14445,N_14528);
nand U14737 (N_14737,N_14599,N_14435);
and U14738 (N_14738,N_14592,N_14449);
or U14739 (N_14739,N_14665,N_14695);
xor U14740 (N_14740,N_14430,N_14659);
nand U14741 (N_14741,N_14549,N_14460);
or U14742 (N_14742,N_14533,N_14478);
and U14743 (N_14743,N_14502,N_14678);
and U14744 (N_14744,N_14496,N_14468);
and U14745 (N_14745,N_14684,N_14634);
nor U14746 (N_14746,N_14527,N_14640);
or U14747 (N_14747,N_14494,N_14575);
nor U14748 (N_14748,N_14696,N_14590);
nor U14749 (N_14749,N_14459,N_14572);
xnor U14750 (N_14750,N_14571,N_14608);
nand U14751 (N_14751,N_14690,N_14604);
xor U14752 (N_14752,N_14493,N_14509);
and U14753 (N_14753,N_14455,N_14510);
nor U14754 (N_14754,N_14542,N_14519);
xnor U14755 (N_14755,N_14481,N_14616);
xor U14756 (N_14756,N_14622,N_14514);
or U14757 (N_14757,N_14467,N_14503);
or U14758 (N_14758,N_14559,N_14658);
or U14759 (N_14759,N_14594,N_14577);
or U14760 (N_14760,N_14532,N_14433);
nand U14761 (N_14761,N_14476,N_14406);
nand U14762 (N_14762,N_14490,N_14641);
xor U14763 (N_14763,N_14475,N_14560);
nand U14764 (N_14764,N_14454,N_14615);
nor U14765 (N_14765,N_14558,N_14477);
or U14766 (N_14766,N_14450,N_14466);
and U14767 (N_14767,N_14429,N_14416);
nand U14768 (N_14768,N_14464,N_14488);
nand U14769 (N_14769,N_14483,N_14663);
nand U14770 (N_14770,N_14569,N_14550);
nand U14771 (N_14771,N_14667,N_14415);
xor U14772 (N_14772,N_14561,N_14683);
xor U14773 (N_14773,N_14579,N_14495);
or U14774 (N_14774,N_14662,N_14606);
nor U14775 (N_14775,N_14453,N_14441);
or U14776 (N_14776,N_14525,N_14422);
nor U14777 (N_14777,N_14500,N_14508);
and U14778 (N_14778,N_14628,N_14648);
nand U14779 (N_14779,N_14501,N_14438);
nor U14780 (N_14780,N_14655,N_14676);
and U14781 (N_14781,N_14436,N_14463);
or U14782 (N_14782,N_14618,N_14613);
xnor U14783 (N_14783,N_14625,N_14432);
and U14784 (N_14784,N_14645,N_14635);
xor U14785 (N_14785,N_14576,N_14551);
or U14786 (N_14786,N_14499,N_14461);
nand U14787 (N_14787,N_14506,N_14587);
xnor U14788 (N_14788,N_14405,N_14689);
nor U14789 (N_14789,N_14544,N_14636);
xnor U14790 (N_14790,N_14567,N_14507);
or U14791 (N_14791,N_14698,N_14685);
xnor U14792 (N_14792,N_14639,N_14687);
or U14793 (N_14793,N_14424,N_14638);
or U14794 (N_14794,N_14675,N_14504);
nor U14795 (N_14795,N_14589,N_14585);
and U14796 (N_14796,N_14439,N_14414);
nor U14797 (N_14797,N_14565,N_14543);
and U14798 (N_14798,N_14553,N_14516);
and U14799 (N_14799,N_14548,N_14556);
and U14800 (N_14800,N_14511,N_14593);
or U14801 (N_14801,N_14446,N_14535);
or U14802 (N_14802,N_14661,N_14692);
and U14803 (N_14803,N_14531,N_14582);
nor U14804 (N_14804,N_14451,N_14699);
nand U14805 (N_14805,N_14562,N_14520);
nand U14806 (N_14806,N_14644,N_14447);
nor U14807 (N_14807,N_14497,N_14465);
nand U14808 (N_14808,N_14573,N_14492);
nand U14809 (N_14809,N_14552,N_14407);
xnor U14810 (N_14810,N_14581,N_14411);
and U14811 (N_14811,N_14623,N_14522);
or U14812 (N_14812,N_14660,N_14491);
xor U14813 (N_14813,N_14583,N_14427);
xor U14814 (N_14814,N_14485,N_14612);
or U14815 (N_14815,N_14591,N_14617);
or U14816 (N_14816,N_14470,N_14677);
nand U14817 (N_14817,N_14633,N_14596);
nand U14818 (N_14818,N_14656,N_14512);
nand U14819 (N_14819,N_14412,N_14524);
nand U14820 (N_14820,N_14610,N_14679);
xnor U14821 (N_14821,N_14471,N_14654);
nor U14822 (N_14822,N_14588,N_14697);
nand U14823 (N_14823,N_14566,N_14563);
or U14824 (N_14824,N_14482,N_14646);
xnor U14825 (N_14825,N_14431,N_14688);
nor U14826 (N_14826,N_14457,N_14498);
or U14827 (N_14827,N_14681,N_14642);
or U14828 (N_14828,N_14621,N_14666);
nand U14829 (N_14829,N_14425,N_14586);
nand U14830 (N_14830,N_14557,N_14472);
nand U14831 (N_14831,N_14568,N_14693);
xor U14832 (N_14832,N_14480,N_14619);
or U14833 (N_14833,N_14420,N_14664);
and U14834 (N_14834,N_14609,N_14530);
xnor U14835 (N_14835,N_14611,N_14403);
xor U14836 (N_14836,N_14584,N_14428);
xnor U14837 (N_14837,N_14423,N_14574);
or U14838 (N_14838,N_14637,N_14649);
xor U14839 (N_14839,N_14421,N_14452);
or U14840 (N_14840,N_14668,N_14673);
xnor U14841 (N_14841,N_14643,N_14534);
xnor U14842 (N_14842,N_14601,N_14632);
nand U14843 (N_14843,N_14602,N_14540);
nor U14844 (N_14844,N_14518,N_14627);
nand U14845 (N_14845,N_14521,N_14486);
or U14846 (N_14846,N_14603,N_14402);
or U14847 (N_14847,N_14474,N_14547);
nor U14848 (N_14848,N_14484,N_14631);
or U14849 (N_14849,N_14647,N_14686);
and U14850 (N_14850,N_14460,N_14439);
nor U14851 (N_14851,N_14508,N_14592);
and U14852 (N_14852,N_14562,N_14429);
xor U14853 (N_14853,N_14502,N_14681);
xnor U14854 (N_14854,N_14526,N_14571);
or U14855 (N_14855,N_14475,N_14691);
or U14856 (N_14856,N_14670,N_14651);
and U14857 (N_14857,N_14618,N_14607);
nand U14858 (N_14858,N_14645,N_14584);
nand U14859 (N_14859,N_14471,N_14494);
and U14860 (N_14860,N_14507,N_14603);
xnor U14861 (N_14861,N_14557,N_14437);
or U14862 (N_14862,N_14671,N_14402);
nor U14863 (N_14863,N_14618,N_14555);
nor U14864 (N_14864,N_14520,N_14425);
and U14865 (N_14865,N_14517,N_14428);
nor U14866 (N_14866,N_14414,N_14552);
nor U14867 (N_14867,N_14534,N_14414);
nor U14868 (N_14868,N_14684,N_14560);
or U14869 (N_14869,N_14543,N_14448);
nand U14870 (N_14870,N_14545,N_14418);
nor U14871 (N_14871,N_14560,N_14601);
nor U14872 (N_14872,N_14487,N_14534);
nand U14873 (N_14873,N_14693,N_14427);
or U14874 (N_14874,N_14465,N_14484);
nand U14875 (N_14875,N_14511,N_14601);
nand U14876 (N_14876,N_14578,N_14469);
and U14877 (N_14877,N_14689,N_14538);
nor U14878 (N_14878,N_14423,N_14623);
nand U14879 (N_14879,N_14512,N_14681);
or U14880 (N_14880,N_14541,N_14692);
nand U14881 (N_14881,N_14469,N_14490);
and U14882 (N_14882,N_14664,N_14515);
nand U14883 (N_14883,N_14461,N_14506);
nor U14884 (N_14884,N_14670,N_14518);
nor U14885 (N_14885,N_14416,N_14525);
and U14886 (N_14886,N_14636,N_14417);
nor U14887 (N_14887,N_14691,N_14417);
xor U14888 (N_14888,N_14470,N_14505);
nor U14889 (N_14889,N_14498,N_14674);
nor U14890 (N_14890,N_14402,N_14665);
and U14891 (N_14891,N_14459,N_14579);
xor U14892 (N_14892,N_14692,N_14485);
nor U14893 (N_14893,N_14529,N_14618);
nand U14894 (N_14894,N_14567,N_14670);
xor U14895 (N_14895,N_14510,N_14575);
nand U14896 (N_14896,N_14645,N_14681);
and U14897 (N_14897,N_14510,N_14587);
and U14898 (N_14898,N_14611,N_14498);
nor U14899 (N_14899,N_14578,N_14529);
xnor U14900 (N_14900,N_14417,N_14615);
nand U14901 (N_14901,N_14508,N_14449);
nand U14902 (N_14902,N_14536,N_14493);
or U14903 (N_14903,N_14536,N_14517);
nor U14904 (N_14904,N_14616,N_14620);
or U14905 (N_14905,N_14409,N_14487);
xor U14906 (N_14906,N_14638,N_14410);
or U14907 (N_14907,N_14685,N_14612);
xor U14908 (N_14908,N_14417,N_14590);
xor U14909 (N_14909,N_14617,N_14534);
nand U14910 (N_14910,N_14539,N_14406);
xnor U14911 (N_14911,N_14664,N_14691);
and U14912 (N_14912,N_14699,N_14552);
nor U14913 (N_14913,N_14641,N_14628);
nor U14914 (N_14914,N_14570,N_14472);
xnor U14915 (N_14915,N_14692,N_14633);
xor U14916 (N_14916,N_14566,N_14640);
and U14917 (N_14917,N_14670,N_14603);
and U14918 (N_14918,N_14643,N_14457);
nand U14919 (N_14919,N_14669,N_14519);
xor U14920 (N_14920,N_14606,N_14473);
xnor U14921 (N_14921,N_14515,N_14425);
or U14922 (N_14922,N_14542,N_14582);
xor U14923 (N_14923,N_14689,N_14465);
xnor U14924 (N_14924,N_14605,N_14590);
nand U14925 (N_14925,N_14579,N_14626);
xor U14926 (N_14926,N_14544,N_14425);
and U14927 (N_14927,N_14648,N_14521);
and U14928 (N_14928,N_14680,N_14564);
xor U14929 (N_14929,N_14445,N_14542);
or U14930 (N_14930,N_14541,N_14664);
xor U14931 (N_14931,N_14639,N_14440);
nand U14932 (N_14932,N_14497,N_14678);
and U14933 (N_14933,N_14600,N_14542);
xor U14934 (N_14934,N_14693,N_14624);
and U14935 (N_14935,N_14470,N_14635);
and U14936 (N_14936,N_14462,N_14439);
or U14937 (N_14937,N_14491,N_14400);
or U14938 (N_14938,N_14515,N_14692);
nand U14939 (N_14939,N_14543,N_14664);
or U14940 (N_14940,N_14490,N_14669);
xnor U14941 (N_14941,N_14585,N_14551);
xor U14942 (N_14942,N_14419,N_14424);
and U14943 (N_14943,N_14586,N_14637);
xor U14944 (N_14944,N_14510,N_14452);
nor U14945 (N_14945,N_14512,N_14426);
and U14946 (N_14946,N_14427,N_14546);
xor U14947 (N_14947,N_14515,N_14404);
and U14948 (N_14948,N_14664,N_14488);
nand U14949 (N_14949,N_14552,N_14491);
and U14950 (N_14950,N_14646,N_14519);
or U14951 (N_14951,N_14425,N_14552);
nor U14952 (N_14952,N_14431,N_14619);
nand U14953 (N_14953,N_14588,N_14510);
nor U14954 (N_14954,N_14556,N_14407);
nand U14955 (N_14955,N_14514,N_14469);
nor U14956 (N_14956,N_14583,N_14441);
nor U14957 (N_14957,N_14506,N_14598);
nor U14958 (N_14958,N_14523,N_14451);
and U14959 (N_14959,N_14481,N_14543);
nor U14960 (N_14960,N_14624,N_14452);
xor U14961 (N_14961,N_14557,N_14457);
or U14962 (N_14962,N_14487,N_14592);
nor U14963 (N_14963,N_14673,N_14464);
or U14964 (N_14964,N_14532,N_14523);
and U14965 (N_14965,N_14502,N_14461);
and U14966 (N_14966,N_14401,N_14460);
xor U14967 (N_14967,N_14618,N_14547);
and U14968 (N_14968,N_14695,N_14552);
or U14969 (N_14969,N_14535,N_14439);
xor U14970 (N_14970,N_14654,N_14418);
nor U14971 (N_14971,N_14542,N_14682);
nor U14972 (N_14972,N_14435,N_14647);
and U14973 (N_14973,N_14421,N_14590);
nand U14974 (N_14974,N_14662,N_14418);
or U14975 (N_14975,N_14617,N_14661);
xor U14976 (N_14976,N_14656,N_14614);
nor U14977 (N_14977,N_14643,N_14444);
and U14978 (N_14978,N_14541,N_14405);
or U14979 (N_14979,N_14432,N_14579);
and U14980 (N_14980,N_14671,N_14400);
and U14981 (N_14981,N_14687,N_14670);
or U14982 (N_14982,N_14552,N_14484);
and U14983 (N_14983,N_14568,N_14500);
and U14984 (N_14984,N_14438,N_14619);
xnor U14985 (N_14985,N_14642,N_14540);
nor U14986 (N_14986,N_14594,N_14616);
xor U14987 (N_14987,N_14439,N_14684);
nor U14988 (N_14988,N_14445,N_14441);
or U14989 (N_14989,N_14411,N_14545);
or U14990 (N_14990,N_14420,N_14408);
xnor U14991 (N_14991,N_14520,N_14616);
nand U14992 (N_14992,N_14485,N_14585);
xor U14993 (N_14993,N_14429,N_14462);
nand U14994 (N_14994,N_14575,N_14478);
and U14995 (N_14995,N_14607,N_14436);
nand U14996 (N_14996,N_14602,N_14515);
nor U14997 (N_14997,N_14478,N_14549);
nand U14998 (N_14998,N_14656,N_14627);
and U14999 (N_14999,N_14641,N_14405);
or UO_0 (O_0,N_14744,N_14772);
and UO_1 (O_1,N_14887,N_14912);
nand UO_2 (O_2,N_14839,N_14818);
xnor UO_3 (O_3,N_14988,N_14925);
nor UO_4 (O_4,N_14823,N_14817);
and UO_5 (O_5,N_14845,N_14796);
and UO_6 (O_6,N_14940,N_14997);
or UO_7 (O_7,N_14707,N_14765);
or UO_8 (O_8,N_14907,N_14703);
and UO_9 (O_9,N_14749,N_14780);
nand UO_10 (O_10,N_14728,N_14806);
and UO_11 (O_11,N_14775,N_14730);
nor UO_12 (O_12,N_14939,N_14785);
or UO_13 (O_13,N_14978,N_14945);
nand UO_14 (O_14,N_14754,N_14769);
or UO_15 (O_15,N_14941,N_14974);
xor UO_16 (O_16,N_14899,N_14748);
and UO_17 (O_17,N_14724,N_14864);
nand UO_18 (O_18,N_14727,N_14853);
xor UO_19 (O_19,N_14846,N_14898);
xnor UO_20 (O_20,N_14992,N_14778);
nand UO_21 (O_21,N_14783,N_14847);
xnor UO_22 (O_22,N_14920,N_14874);
or UO_23 (O_23,N_14950,N_14848);
nor UO_24 (O_24,N_14731,N_14762);
and UO_25 (O_25,N_14927,N_14779);
and UO_26 (O_26,N_14811,N_14975);
or UO_27 (O_27,N_14715,N_14968);
nand UO_28 (O_28,N_14850,N_14717);
nand UO_29 (O_29,N_14756,N_14800);
and UO_30 (O_30,N_14725,N_14931);
xor UO_31 (O_31,N_14856,N_14757);
and UO_32 (O_32,N_14809,N_14700);
and UO_33 (O_33,N_14802,N_14930);
and UO_34 (O_34,N_14781,N_14739);
xnor UO_35 (O_35,N_14750,N_14770);
xor UO_36 (O_36,N_14958,N_14763);
or UO_37 (O_37,N_14753,N_14702);
xor UO_38 (O_38,N_14921,N_14840);
xnor UO_39 (O_39,N_14999,N_14886);
or UO_40 (O_40,N_14760,N_14943);
or UO_41 (O_41,N_14926,N_14877);
nand UO_42 (O_42,N_14909,N_14803);
or UO_43 (O_43,N_14878,N_14949);
xnor UO_44 (O_44,N_14734,N_14929);
nor UO_45 (O_45,N_14774,N_14977);
or UO_46 (O_46,N_14922,N_14953);
or UO_47 (O_47,N_14746,N_14913);
and UO_48 (O_48,N_14880,N_14837);
xnor UO_49 (O_49,N_14870,N_14918);
nand UO_50 (O_50,N_14808,N_14732);
and UO_51 (O_51,N_14881,N_14736);
nand UO_52 (O_52,N_14790,N_14793);
and UO_53 (O_53,N_14718,N_14733);
xor UO_54 (O_54,N_14832,N_14914);
xor UO_55 (O_55,N_14807,N_14709);
or UO_56 (O_56,N_14984,N_14743);
and UO_57 (O_57,N_14737,N_14726);
nor UO_58 (O_58,N_14972,N_14860);
nand UO_59 (O_59,N_14982,N_14901);
or UO_60 (O_60,N_14966,N_14956);
nand UO_61 (O_61,N_14824,N_14720);
xnor UO_62 (O_62,N_14712,N_14986);
and UO_63 (O_63,N_14841,N_14723);
nor UO_64 (O_64,N_14721,N_14863);
and UO_65 (O_65,N_14771,N_14890);
nand UO_66 (O_66,N_14962,N_14871);
xnor UO_67 (O_67,N_14891,N_14810);
nor UO_68 (O_68,N_14758,N_14934);
and UO_69 (O_69,N_14716,N_14825);
nor UO_70 (O_70,N_14829,N_14704);
nor UO_71 (O_71,N_14843,N_14916);
or UO_72 (O_72,N_14741,N_14838);
nor UO_73 (O_73,N_14936,N_14998);
nand UO_74 (O_74,N_14814,N_14820);
nand UO_75 (O_75,N_14745,N_14861);
xnor UO_76 (O_76,N_14791,N_14852);
nor UO_77 (O_77,N_14917,N_14714);
nor UO_78 (O_78,N_14713,N_14967);
or UO_79 (O_79,N_14964,N_14928);
xnor UO_80 (O_80,N_14855,N_14888);
or UO_81 (O_81,N_14862,N_14875);
or UO_82 (O_82,N_14834,N_14924);
xor UO_83 (O_83,N_14904,N_14902);
or UO_84 (O_84,N_14854,N_14897);
nor UO_85 (O_85,N_14900,N_14859);
and UO_86 (O_86,N_14797,N_14767);
xor UO_87 (O_87,N_14844,N_14946);
nand UO_88 (O_88,N_14873,N_14755);
nand UO_89 (O_89,N_14794,N_14867);
nand UO_90 (O_90,N_14786,N_14995);
xnor UO_91 (O_91,N_14915,N_14932);
or UO_92 (O_92,N_14935,N_14799);
nand UO_93 (O_93,N_14944,N_14951);
and UO_94 (O_94,N_14827,N_14816);
nand UO_95 (O_95,N_14990,N_14910);
xor UO_96 (O_96,N_14719,N_14801);
nand UO_97 (O_97,N_14961,N_14911);
or UO_98 (O_98,N_14759,N_14821);
or UO_99 (O_99,N_14869,N_14789);
and UO_100 (O_100,N_14895,N_14994);
nand UO_101 (O_101,N_14815,N_14738);
nor UO_102 (O_102,N_14740,N_14960);
or UO_103 (O_103,N_14706,N_14747);
or UO_104 (O_104,N_14849,N_14711);
xnor UO_105 (O_105,N_14865,N_14812);
nand UO_106 (O_106,N_14828,N_14947);
or UO_107 (O_107,N_14937,N_14908);
nand UO_108 (O_108,N_14868,N_14955);
nor UO_109 (O_109,N_14858,N_14882);
nor UO_110 (O_110,N_14776,N_14701);
or UO_111 (O_111,N_14708,N_14792);
nand UO_112 (O_112,N_14833,N_14831);
xor UO_113 (O_113,N_14954,N_14896);
nand UO_114 (O_114,N_14764,N_14948);
nor UO_115 (O_115,N_14784,N_14836);
or UO_116 (O_116,N_14872,N_14893);
nand UO_117 (O_117,N_14813,N_14766);
nor UO_118 (O_118,N_14826,N_14980);
nor UO_119 (O_119,N_14705,N_14795);
xor UO_120 (O_120,N_14959,N_14979);
or UO_121 (O_121,N_14787,N_14965);
nand UO_122 (O_122,N_14842,N_14903);
or UO_123 (O_123,N_14991,N_14782);
and UO_124 (O_124,N_14798,N_14761);
and UO_125 (O_125,N_14710,N_14957);
nand UO_126 (O_126,N_14989,N_14788);
or UO_127 (O_127,N_14851,N_14866);
nand UO_128 (O_128,N_14973,N_14805);
and UO_129 (O_129,N_14996,N_14933);
nand UO_130 (O_130,N_14889,N_14768);
or UO_131 (O_131,N_14987,N_14981);
xnor UO_132 (O_132,N_14735,N_14777);
or UO_133 (O_133,N_14751,N_14883);
nor UO_134 (O_134,N_14876,N_14976);
nand UO_135 (O_135,N_14970,N_14919);
nand UO_136 (O_136,N_14938,N_14985);
nand UO_137 (O_137,N_14905,N_14722);
and UO_138 (O_138,N_14742,N_14923);
or UO_139 (O_139,N_14804,N_14971);
nand UO_140 (O_140,N_14952,N_14773);
or UO_141 (O_141,N_14963,N_14892);
xor UO_142 (O_142,N_14894,N_14822);
or UO_143 (O_143,N_14983,N_14819);
and UO_144 (O_144,N_14969,N_14942);
or UO_145 (O_145,N_14906,N_14830);
nand UO_146 (O_146,N_14993,N_14835);
and UO_147 (O_147,N_14884,N_14729);
xor UO_148 (O_148,N_14879,N_14857);
nor UO_149 (O_149,N_14752,N_14885);
nand UO_150 (O_150,N_14893,N_14745);
xnor UO_151 (O_151,N_14719,N_14893);
nand UO_152 (O_152,N_14905,N_14711);
xor UO_153 (O_153,N_14958,N_14909);
or UO_154 (O_154,N_14967,N_14813);
or UO_155 (O_155,N_14808,N_14847);
nor UO_156 (O_156,N_14792,N_14842);
xnor UO_157 (O_157,N_14788,N_14896);
nor UO_158 (O_158,N_14878,N_14966);
nor UO_159 (O_159,N_14988,N_14768);
and UO_160 (O_160,N_14931,N_14901);
and UO_161 (O_161,N_14831,N_14834);
or UO_162 (O_162,N_14739,N_14727);
and UO_163 (O_163,N_14870,N_14773);
or UO_164 (O_164,N_14944,N_14937);
and UO_165 (O_165,N_14917,N_14867);
xnor UO_166 (O_166,N_14832,N_14713);
nor UO_167 (O_167,N_14838,N_14789);
and UO_168 (O_168,N_14959,N_14712);
xor UO_169 (O_169,N_14922,N_14712);
xnor UO_170 (O_170,N_14823,N_14992);
nand UO_171 (O_171,N_14876,N_14883);
xnor UO_172 (O_172,N_14810,N_14722);
nand UO_173 (O_173,N_14815,N_14702);
or UO_174 (O_174,N_14938,N_14740);
nor UO_175 (O_175,N_14755,N_14743);
or UO_176 (O_176,N_14706,N_14872);
xnor UO_177 (O_177,N_14818,N_14945);
and UO_178 (O_178,N_14835,N_14817);
xor UO_179 (O_179,N_14746,N_14825);
and UO_180 (O_180,N_14752,N_14837);
or UO_181 (O_181,N_14923,N_14833);
and UO_182 (O_182,N_14960,N_14895);
xnor UO_183 (O_183,N_14740,N_14996);
nand UO_184 (O_184,N_14876,N_14715);
xor UO_185 (O_185,N_14956,N_14811);
nand UO_186 (O_186,N_14813,N_14925);
and UO_187 (O_187,N_14774,N_14943);
and UO_188 (O_188,N_14746,N_14720);
or UO_189 (O_189,N_14732,N_14901);
nor UO_190 (O_190,N_14812,N_14735);
nand UO_191 (O_191,N_14700,N_14715);
nor UO_192 (O_192,N_14863,N_14892);
and UO_193 (O_193,N_14878,N_14772);
nand UO_194 (O_194,N_14742,N_14701);
or UO_195 (O_195,N_14791,N_14736);
nand UO_196 (O_196,N_14750,N_14775);
and UO_197 (O_197,N_14746,N_14776);
or UO_198 (O_198,N_14995,N_14725);
or UO_199 (O_199,N_14832,N_14850);
nand UO_200 (O_200,N_14948,N_14803);
nand UO_201 (O_201,N_14838,N_14962);
xnor UO_202 (O_202,N_14992,N_14716);
nand UO_203 (O_203,N_14792,N_14767);
nor UO_204 (O_204,N_14708,N_14942);
xor UO_205 (O_205,N_14942,N_14994);
xor UO_206 (O_206,N_14773,N_14772);
xnor UO_207 (O_207,N_14901,N_14813);
nand UO_208 (O_208,N_14961,N_14938);
nor UO_209 (O_209,N_14935,N_14940);
nor UO_210 (O_210,N_14867,N_14770);
xor UO_211 (O_211,N_14830,N_14834);
or UO_212 (O_212,N_14994,N_14729);
or UO_213 (O_213,N_14715,N_14738);
xor UO_214 (O_214,N_14728,N_14853);
nor UO_215 (O_215,N_14808,N_14878);
nand UO_216 (O_216,N_14744,N_14852);
or UO_217 (O_217,N_14935,N_14763);
nor UO_218 (O_218,N_14771,N_14880);
or UO_219 (O_219,N_14826,N_14769);
or UO_220 (O_220,N_14991,N_14833);
nand UO_221 (O_221,N_14899,N_14942);
and UO_222 (O_222,N_14940,N_14930);
and UO_223 (O_223,N_14881,N_14792);
xor UO_224 (O_224,N_14910,N_14851);
or UO_225 (O_225,N_14973,N_14825);
and UO_226 (O_226,N_14717,N_14780);
or UO_227 (O_227,N_14950,N_14745);
and UO_228 (O_228,N_14757,N_14967);
xnor UO_229 (O_229,N_14724,N_14725);
and UO_230 (O_230,N_14745,N_14946);
xnor UO_231 (O_231,N_14738,N_14833);
and UO_232 (O_232,N_14781,N_14810);
nor UO_233 (O_233,N_14807,N_14819);
and UO_234 (O_234,N_14762,N_14867);
nor UO_235 (O_235,N_14909,N_14717);
xnor UO_236 (O_236,N_14893,N_14914);
nor UO_237 (O_237,N_14891,N_14732);
and UO_238 (O_238,N_14922,N_14914);
or UO_239 (O_239,N_14881,N_14837);
xor UO_240 (O_240,N_14720,N_14956);
nor UO_241 (O_241,N_14902,N_14758);
xnor UO_242 (O_242,N_14832,N_14794);
nor UO_243 (O_243,N_14983,N_14833);
nor UO_244 (O_244,N_14725,N_14819);
or UO_245 (O_245,N_14981,N_14894);
or UO_246 (O_246,N_14784,N_14729);
and UO_247 (O_247,N_14843,N_14780);
nand UO_248 (O_248,N_14981,N_14926);
and UO_249 (O_249,N_14914,N_14713);
nand UO_250 (O_250,N_14757,N_14732);
or UO_251 (O_251,N_14981,N_14831);
or UO_252 (O_252,N_14971,N_14995);
or UO_253 (O_253,N_14787,N_14917);
or UO_254 (O_254,N_14910,N_14814);
or UO_255 (O_255,N_14978,N_14813);
or UO_256 (O_256,N_14971,N_14953);
or UO_257 (O_257,N_14937,N_14883);
nand UO_258 (O_258,N_14802,N_14755);
xor UO_259 (O_259,N_14953,N_14744);
nor UO_260 (O_260,N_14846,N_14950);
nand UO_261 (O_261,N_14974,N_14872);
or UO_262 (O_262,N_14799,N_14833);
or UO_263 (O_263,N_14842,N_14998);
and UO_264 (O_264,N_14724,N_14998);
nor UO_265 (O_265,N_14948,N_14808);
nand UO_266 (O_266,N_14961,N_14773);
nand UO_267 (O_267,N_14863,N_14994);
nand UO_268 (O_268,N_14870,N_14855);
or UO_269 (O_269,N_14916,N_14869);
nand UO_270 (O_270,N_14827,N_14859);
or UO_271 (O_271,N_14712,N_14807);
or UO_272 (O_272,N_14706,N_14770);
nand UO_273 (O_273,N_14768,N_14837);
or UO_274 (O_274,N_14880,N_14867);
nand UO_275 (O_275,N_14979,N_14962);
and UO_276 (O_276,N_14761,N_14952);
and UO_277 (O_277,N_14918,N_14923);
xnor UO_278 (O_278,N_14752,N_14955);
or UO_279 (O_279,N_14707,N_14824);
or UO_280 (O_280,N_14831,N_14867);
nand UO_281 (O_281,N_14786,N_14836);
nand UO_282 (O_282,N_14837,N_14999);
or UO_283 (O_283,N_14999,N_14896);
or UO_284 (O_284,N_14868,N_14731);
and UO_285 (O_285,N_14798,N_14805);
nor UO_286 (O_286,N_14790,N_14775);
nand UO_287 (O_287,N_14805,N_14993);
and UO_288 (O_288,N_14819,N_14705);
nor UO_289 (O_289,N_14884,N_14916);
or UO_290 (O_290,N_14711,N_14900);
nand UO_291 (O_291,N_14730,N_14983);
xor UO_292 (O_292,N_14726,N_14970);
and UO_293 (O_293,N_14795,N_14939);
nand UO_294 (O_294,N_14870,N_14958);
nor UO_295 (O_295,N_14776,N_14949);
nand UO_296 (O_296,N_14869,N_14895);
xnor UO_297 (O_297,N_14962,N_14707);
nand UO_298 (O_298,N_14972,N_14703);
nor UO_299 (O_299,N_14898,N_14988);
nor UO_300 (O_300,N_14896,N_14998);
and UO_301 (O_301,N_14803,N_14934);
nor UO_302 (O_302,N_14920,N_14944);
and UO_303 (O_303,N_14844,N_14881);
or UO_304 (O_304,N_14775,N_14909);
xnor UO_305 (O_305,N_14915,N_14751);
or UO_306 (O_306,N_14865,N_14782);
and UO_307 (O_307,N_14963,N_14948);
xor UO_308 (O_308,N_14863,N_14714);
xor UO_309 (O_309,N_14799,N_14832);
and UO_310 (O_310,N_14842,N_14754);
nor UO_311 (O_311,N_14996,N_14806);
xor UO_312 (O_312,N_14936,N_14810);
nand UO_313 (O_313,N_14971,N_14783);
nand UO_314 (O_314,N_14996,N_14787);
or UO_315 (O_315,N_14792,N_14706);
nand UO_316 (O_316,N_14862,N_14712);
nand UO_317 (O_317,N_14732,N_14906);
or UO_318 (O_318,N_14969,N_14834);
and UO_319 (O_319,N_14969,N_14724);
nor UO_320 (O_320,N_14845,N_14826);
or UO_321 (O_321,N_14789,N_14926);
xnor UO_322 (O_322,N_14985,N_14970);
xor UO_323 (O_323,N_14837,N_14706);
nand UO_324 (O_324,N_14728,N_14776);
or UO_325 (O_325,N_14852,N_14814);
and UO_326 (O_326,N_14833,N_14931);
xnor UO_327 (O_327,N_14724,N_14852);
nor UO_328 (O_328,N_14837,N_14948);
xnor UO_329 (O_329,N_14945,N_14812);
nor UO_330 (O_330,N_14942,N_14882);
nor UO_331 (O_331,N_14776,N_14967);
nand UO_332 (O_332,N_14837,N_14702);
and UO_333 (O_333,N_14890,N_14915);
and UO_334 (O_334,N_14726,N_14778);
xor UO_335 (O_335,N_14821,N_14893);
and UO_336 (O_336,N_14969,N_14702);
xnor UO_337 (O_337,N_14834,N_14780);
or UO_338 (O_338,N_14998,N_14871);
nand UO_339 (O_339,N_14730,N_14812);
nor UO_340 (O_340,N_14861,N_14986);
and UO_341 (O_341,N_14915,N_14972);
nand UO_342 (O_342,N_14722,N_14889);
nor UO_343 (O_343,N_14915,N_14863);
nor UO_344 (O_344,N_14774,N_14956);
xor UO_345 (O_345,N_14943,N_14733);
and UO_346 (O_346,N_14838,N_14777);
and UO_347 (O_347,N_14900,N_14869);
and UO_348 (O_348,N_14754,N_14733);
nand UO_349 (O_349,N_14945,N_14888);
xor UO_350 (O_350,N_14747,N_14878);
nand UO_351 (O_351,N_14994,N_14776);
or UO_352 (O_352,N_14983,N_14957);
xnor UO_353 (O_353,N_14858,N_14714);
nand UO_354 (O_354,N_14869,N_14961);
and UO_355 (O_355,N_14957,N_14892);
or UO_356 (O_356,N_14769,N_14850);
nor UO_357 (O_357,N_14958,N_14934);
and UO_358 (O_358,N_14897,N_14852);
or UO_359 (O_359,N_14974,N_14796);
nor UO_360 (O_360,N_14762,N_14803);
or UO_361 (O_361,N_14961,N_14956);
or UO_362 (O_362,N_14861,N_14871);
xor UO_363 (O_363,N_14703,N_14929);
nand UO_364 (O_364,N_14917,N_14896);
xnor UO_365 (O_365,N_14860,N_14923);
or UO_366 (O_366,N_14936,N_14834);
nand UO_367 (O_367,N_14842,N_14733);
or UO_368 (O_368,N_14925,N_14706);
and UO_369 (O_369,N_14792,N_14852);
or UO_370 (O_370,N_14812,N_14738);
and UO_371 (O_371,N_14741,N_14971);
and UO_372 (O_372,N_14948,N_14759);
or UO_373 (O_373,N_14796,N_14732);
nand UO_374 (O_374,N_14804,N_14911);
or UO_375 (O_375,N_14781,N_14755);
and UO_376 (O_376,N_14859,N_14726);
nand UO_377 (O_377,N_14881,N_14853);
and UO_378 (O_378,N_14961,N_14738);
and UO_379 (O_379,N_14712,N_14795);
and UO_380 (O_380,N_14753,N_14950);
xor UO_381 (O_381,N_14927,N_14837);
xnor UO_382 (O_382,N_14815,N_14919);
xnor UO_383 (O_383,N_14748,N_14808);
xnor UO_384 (O_384,N_14837,N_14832);
xnor UO_385 (O_385,N_14917,N_14791);
nor UO_386 (O_386,N_14842,N_14962);
xnor UO_387 (O_387,N_14891,N_14721);
or UO_388 (O_388,N_14897,N_14836);
xnor UO_389 (O_389,N_14901,N_14967);
nand UO_390 (O_390,N_14828,N_14857);
and UO_391 (O_391,N_14801,N_14973);
xor UO_392 (O_392,N_14936,N_14978);
xnor UO_393 (O_393,N_14769,N_14861);
nand UO_394 (O_394,N_14815,N_14938);
nand UO_395 (O_395,N_14779,N_14965);
nand UO_396 (O_396,N_14944,N_14909);
or UO_397 (O_397,N_14920,N_14953);
xnor UO_398 (O_398,N_14984,N_14965);
nor UO_399 (O_399,N_14941,N_14830);
nor UO_400 (O_400,N_14974,N_14750);
nand UO_401 (O_401,N_14793,N_14826);
or UO_402 (O_402,N_14728,N_14899);
nor UO_403 (O_403,N_14708,N_14924);
nor UO_404 (O_404,N_14927,N_14986);
and UO_405 (O_405,N_14960,N_14915);
nand UO_406 (O_406,N_14895,N_14773);
nand UO_407 (O_407,N_14740,N_14987);
or UO_408 (O_408,N_14774,N_14959);
or UO_409 (O_409,N_14877,N_14793);
xnor UO_410 (O_410,N_14877,N_14706);
nand UO_411 (O_411,N_14873,N_14859);
and UO_412 (O_412,N_14767,N_14836);
or UO_413 (O_413,N_14802,N_14959);
xnor UO_414 (O_414,N_14825,N_14803);
nor UO_415 (O_415,N_14804,N_14977);
nor UO_416 (O_416,N_14729,N_14957);
and UO_417 (O_417,N_14837,N_14734);
xnor UO_418 (O_418,N_14731,N_14843);
xor UO_419 (O_419,N_14950,N_14971);
or UO_420 (O_420,N_14894,N_14939);
xnor UO_421 (O_421,N_14757,N_14907);
and UO_422 (O_422,N_14759,N_14974);
xnor UO_423 (O_423,N_14928,N_14861);
xor UO_424 (O_424,N_14734,N_14913);
and UO_425 (O_425,N_14879,N_14756);
and UO_426 (O_426,N_14992,N_14709);
and UO_427 (O_427,N_14766,N_14941);
nor UO_428 (O_428,N_14859,N_14951);
or UO_429 (O_429,N_14934,N_14724);
nor UO_430 (O_430,N_14796,N_14717);
nor UO_431 (O_431,N_14722,N_14794);
and UO_432 (O_432,N_14759,N_14918);
nor UO_433 (O_433,N_14784,N_14831);
or UO_434 (O_434,N_14944,N_14835);
nand UO_435 (O_435,N_14817,N_14971);
nand UO_436 (O_436,N_14726,N_14777);
or UO_437 (O_437,N_14861,N_14960);
and UO_438 (O_438,N_14931,N_14709);
xnor UO_439 (O_439,N_14813,N_14870);
xor UO_440 (O_440,N_14998,N_14994);
and UO_441 (O_441,N_14727,N_14903);
nand UO_442 (O_442,N_14729,N_14733);
and UO_443 (O_443,N_14835,N_14735);
and UO_444 (O_444,N_14751,N_14877);
nor UO_445 (O_445,N_14853,N_14779);
nor UO_446 (O_446,N_14985,N_14818);
and UO_447 (O_447,N_14792,N_14942);
and UO_448 (O_448,N_14722,N_14977);
xnor UO_449 (O_449,N_14807,N_14925);
nor UO_450 (O_450,N_14897,N_14982);
nand UO_451 (O_451,N_14851,N_14751);
nand UO_452 (O_452,N_14726,N_14815);
and UO_453 (O_453,N_14798,N_14804);
or UO_454 (O_454,N_14942,N_14802);
nand UO_455 (O_455,N_14741,N_14743);
nor UO_456 (O_456,N_14857,N_14785);
xnor UO_457 (O_457,N_14786,N_14756);
xnor UO_458 (O_458,N_14913,N_14806);
and UO_459 (O_459,N_14944,N_14924);
nand UO_460 (O_460,N_14772,N_14719);
nor UO_461 (O_461,N_14812,N_14833);
or UO_462 (O_462,N_14996,N_14954);
and UO_463 (O_463,N_14978,N_14916);
xor UO_464 (O_464,N_14863,N_14749);
and UO_465 (O_465,N_14708,N_14990);
or UO_466 (O_466,N_14926,N_14818);
nor UO_467 (O_467,N_14839,N_14786);
and UO_468 (O_468,N_14756,N_14704);
and UO_469 (O_469,N_14981,N_14915);
or UO_470 (O_470,N_14820,N_14798);
and UO_471 (O_471,N_14897,N_14806);
and UO_472 (O_472,N_14967,N_14851);
xor UO_473 (O_473,N_14814,N_14783);
xor UO_474 (O_474,N_14965,N_14700);
or UO_475 (O_475,N_14940,N_14926);
xor UO_476 (O_476,N_14834,N_14846);
nor UO_477 (O_477,N_14711,N_14716);
xor UO_478 (O_478,N_14955,N_14978);
xnor UO_479 (O_479,N_14947,N_14819);
or UO_480 (O_480,N_14826,N_14836);
or UO_481 (O_481,N_14810,N_14964);
nor UO_482 (O_482,N_14722,N_14715);
xnor UO_483 (O_483,N_14976,N_14865);
or UO_484 (O_484,N_14845,N_14940);
nor UO_485 (O_485,N_14917,N_14743);
nand UO_486 (O_486,N_14706,N_14990);
nor UO_487 (O_487,N_14701,N_14876);
nand UO_488 (O_488,N_14966,N_14777);
and UO_489 (O_489,N_14818,N_14857);
nand UO_490 (O_490,N_14781,N_14797);
nor UO_491 (O_491,N_14903,N_14999);
and UO_492 (O_492,N_14790,N_14798);
and UO_493 (O_493,N_14923,N_14813);
nor UO_494 (O_494,N_14925,N_14798);
nor UO_495 (O_495,N_14913,N_14861);
nor UO_496 (O_496,N_14919,N_14972);
nor UO_497 (O_497,N_14713,N_14812);
or UO_498 (O_498,N_14787,N_14971);
and UO_499 (O_499,N_14743,N_14894);
xnor UO_500 (O_500,N_14765,N_14744);
or UO_501 (O_501,N_14802,N_14923);
nand UO_502 (O_502,N_14768,N_14913);
nand UO_503 (O_503,N_14851,N_14746);
nand UO_504 (O_504,N_14896,N_14955);
nor UO_505 (O_505,N_14827,N_14855);
and UO_506 (O_506,N_14836,N_14930);
xor UO_507 (O_507,N_14852,N_14745);
or UO_508 (O_508,N_14849,N_14792);
nor UO_509 (O_509,N_14926,N_14815);
nand UO_510 (O_510,N_14852,N_14949);
xor UO_511 (O_511,N_14808,N_14707);
nor UO_512 (O_512,N_14785,N_14751);
nor UO_513 (O_513,N_14923,N_14768);
or UO_514 (O_514,N_14770,N_14989);
nand UO_515 (O_515,N_14881,N_14845);
and UO_516 (O_516,N_14825,N_14960);
nand UO_517 (O_517,N_14851,N_14777);
xor UO_518 (O_518,N_14844,N_14912);
and UO_519 (O_519,N_14825,N_14879);
or UO_520 (O_520,N_14758,N_14909);
xnor UO_521 (O_521,N_14753,N_14996);
xnor UO_522 (O_522,N_14846,N_14789);
and UO_523 (O_523,N_14838,N_14793);
nor UO_524 (O_524,N_14756,N_14826);
xor UO_525 (O_525,N_14830,N_14829);
nand UO_526 (O_526,N_14915,N_14737);
or UO_527 (O_527,N_14775,N_14830);
nand UO_528 (O_528,N_14786,N_14804);
nand UO_529 (O_529,N_14703,N_14991);
xor UO_530 (O_530,N_14854,N_14923);
or UO_531 (O_531,N_14799,N_14959);
xnor UO_532 (O_532,N_14918,N_14768);
or UO_533 (O_533,N_14848,N_14856);
xor UO_534 (O_534,N_14784,N_14940);
nor UO_535 (O_535,N_14880,N_14815);
or UO_536 (O_536,N_14920,N_14933);
xor UO_537 (O_537,N_14886,N_14977);
nand UO_538 (O_538,N_14911,N_14742);
xor UO_539 (O_539,N_14850,N_14872);
and UO_540 (O_540,N_14955,N_14876);
xnor UO_541 (O_541,N_14950,N_14733);
xnor UO_542 (O_542,N_14705,N_14992);
or UO_543 (O_543,N_14948,N_14899);
and UO_544 (O_544,N_14737,N_14794);
nand UO_545 (O_545,N_14714,N_14872);
or UO_546 (O_546,N_14896,N_14720);
xnor UO_547 (O_547,N_14813,N_14799);
xnor UO_548 (O_548,N_14829,N_14918);
and UO_549 (O_549,N_14947,N_14826);
and UO_550 (O_550,N_14723,N_14872);
or UO_551 (O_551,N_14961,N_14732);
nor UO_552 (O_552,N_14857,N_14795);
nor UO_553 (O_553,N_14722,N_14984);
and UO_554 (O_554,N_14807,N_14719);
xnor UO_555 (O_555,N_14791,N_14949);
nor UO_556 (O_556,N_14791,N_14794);
nor UO_557 (O_557,N_14947,N_14910);
nand UO_558 (O_558,N_14707,N_14860);
nor UO_559 (O_559,N_14976,N_14739);
or UO_560 (O_560,N_14792,N_14858);
and UO_561 (O_561,N_14934,N_14756);
and UO_562 (O_562,N_14938,N_14882);
nand UO_563 (O_563,N_14893,N_14918);
nand UO_564 (O_564,N_14727,N_14966);
and UO_565 (O_565,N_14794,N_14746);
and UO_566 (O_566,N_14789,N_14882);
xor UO_567 (O_567,N_14709,N_14987);
xor UO_568 (O_568,N_14721,N_14816);
and UO_569 (O_569,N_14854,N_14752);
or UO_570 (O_570,N_14724,N_14857);
nand UO_571 (O_571,N_14811,N_14939);
or UO_572 (O_572,N_14974,N_14810);
or UO_573 (O_573,N_14769,N_14705);
or UO_574 (O_574,N_14794,N_14914);
nor UO_575 (O_575,N_14755,N_14787);
nand UO_576 (O_576,N_14873,N_14754);
nor UO_577 (O_577,N_14901,N_14842);
nand UO_578 (O_578,N_14776,N_14941);
nand UO_579 (O_579,N_14934,N_14740);
or UO_580 (O_580,N_14756,N_14773);
or UO_581 (O_581,N_14911,N_14960);
nand UO_582 (O_582,N_14854,N_14813);
nand UO_583 (O_583,N_14829,N_14812);
and UO_584 (O_584,N_14717,N_14797);
xor UO_585 (O_585,N_14794,N_14865);
or UO_586 (O_586,N_14759,N_14868);
xnor UO_587 (O_587,N_14736,N_14849);
or UO_588 (O_588,N_14725,N_14957);
nor UO_589 (O_589,N_14911,N_14821);
nor UO_590 (O_590,N_14799,N_14765);
xnor UO_591 (O_591,N_14930,N_14911);
nand UO_592 (O_592,N_14725,N_14996);
xor UO_593 (O_593,N_14849,N_14870);
xnor UO_594 (O_594,N_14775,N_14861);
and UO_595 (O_595,N_14758,N_14729);
nand UO_596 (O_596,N_14892,N_14979);
nor UO_597 (O_597,N_14717,N_14875);
nand UO_598 (O_598,N_14843,N_14745);
nor UO_599 (O_599,N_14988,N_14971);
nand UO_600 (O_600,N_14913,N_14932);
nor UO_601 (O_601,N_14919,N_14784);
nand UO_602 (O_602,N_14890,N_14842);
nor UO_603 (O_603,N_14991,N_14936);
or UO_604 (O_604,N_14780,N_14727);
and UO_605 (O_605,N_14946,N_14982);
nand UO_606 (O_606,N_14778,N_14826);
nand UO_607 (O_607,N_14825,N_14703);
and UO_608 (O_608,N_14970,N_14889);
nor UO_609 (O_609,N_14833,N_14971);
nand UO_610 (O_610,N_14791,N_14838);
and UO_611 (O_611,N_14918,N_14772);
nand UO_612 (O_612,N_14941,N_14808);
nand UO_613 (O_613,N_14820,N_14911);
or UO_614 (O_614,N_14958,N_14840);
and UO_615 (O_615,N_14885,N_14828);
xor UO_616 (O_616,N_14748,N_14893);
nand UO_617 (O_617,N_14970,N_14759);
xor UO_618 (O_618,N_14851,N_14729);
and UO_619 (O_619,N_14934,N_14714);
xor UO_620 (O_620,N_14740,N_14847);
nor UO_621 (O_621,N_14987,N_14888);
xor UO_622 (O_622,N_14923,N_14974);
nand UO_623 (O_623,N_14985,N_14900);
xor UO_624 (O_624,N_14936,N_14919);
and UO_625 (O_625,N_14822,N_14762);
xor UO_626 (O_626,N_14878,N_14841);
nor UO_627 (O_627,N_14995,N_14945);
nand UO_628 (O_628,N_14861,N_14839);
nand UO_629 (O_629,N_14875,N_14912);
nor UO_630 (O_630,N_14811,N_14898);
nand UO_631 (O_631,N_14831,N_14936);
or UO_632 (O_632,N_14777,N_14724);
nand UO_633 (O_633,N_14987,N_14790);
xor UO_634 (O_634,N_14953,N_14771);
nor UO_635 (O_635,N_14821,N_14917);
and UO_636 (O_636,N_14925,N_14702);
and UO_637 (O_637,N_14811,N_14989);
or UO_638 (O_638,N_14952,N_14812);
xor UO_639 (O_639,N_14863,N_14810);
nor UO_640 (O_640,N_14866,N_14923);
nor UO_641 (O_641,N_14762,N_14941);
or UO_642 (O_642,N_14731,N_14806);
or UO_643 (O_643,N_14992,N_14703);
nand UO_644 (O_644,N_14787,N_14707);
or UO_645 (O_645,N_14997,N_14946);
nor UO_646 (O_646,N_14719,N_14916);
xor UO_647 (O_647,N_14873,N_14955);
or UO_648 (O_648,N_14723,N_14818);
and UO_649 (O_649,N_14857,N_14892);
xor UO_650 (O_650,N_14955,N_14911);
nand UO_651 (O_651,N_14851,N_14757);
or UO_652 (O_652,N_14974,N_14808);
and UO_653 (O_653,N_14716,N_14970);
and UO_654 (O_654,N_14939,N_14918);
and UO_655 (O_655,N_14972,N_14786);
nand UO_656 (O_656,N_14872,N_14861);
nand UO_657 (O_657,N_14860,N_14988);
xor UO_658 (O_658,N_14840,N_14775);
xor UO_659 (O_659,N_14920,N_14923);
and UO_660 (O_660,N_14908,N_14817);
nand UO_661 (O_661,N_14752,N_14897);
nor UO_662 (O_662,N_14926,N_14705);
xnor UO_663 (O_663,N_14986,N_14925);
and UO_664 (O_664,N_14835,N_14852);
and UO_665 (O_665,N_14949,N_14824);
nand UO_666 (O_666,N_14914,N_14963);
or UO_667 (O_667,N_14820,N_14805);
nor UO_668 (O_668,N_14920,N_14771);
xnor UO_669 (O_669,N_14839,N_14925);
and UO_670 (O_670,N_14981,N_14875);
and UO_671 (O_671,N_14937,N_14860);
nor UO_672 (O_672,N_14843,N_14929);
and UO_673 (O_673,N_14804,N_14772);
nor UO_674 (O_674,N_14882,N_14821);
and UO_675 (O_675,N_14995,N_14752);
nor UO_676 (O_676,N_14835,N_14877);
or UO_677 (O_677,N_14831,N_14934);
xor UO_678 (O_678,N_14882,N_14829);
xnor UO_679 (O_679,N_14718,N_14822);
and UO_680 (O_680,N_14901,N_14983);
nand UO_681 (O_681,N_14717,N_14771);
or UO_682 (O_682,N_14794,N_14721);
nand UO_683 (O_683,N_14798,N_14894);
nand UO_684 (O_684,N_14903,N_14938);
nor UO_685 (O_685,N_14813,N_14746);
nand UO_686 (O_686,N_14943,N_14953);
and UO_687 (O_687,N_14861,N_14908);
nor UO_688 (O_688,N_14946,N_14937);
and UO_689 (O_689,N_14999,N_14843);
and UO_690 (O_690,N_14979,N_14714);
nor UO_691 (O_691,N_14725,N_14796);
and UO_692 (O_692,N_14804,N_14720);
nand UO_693 (O_693,N_14778,N_14741);
nand UO_694 (O_694,N_14770,N_14992);
xor UO_695 (O_695,N_14720,N_14903);
nand UO_696 (O_696,N_14796,N_14804);
and UO_697 (O_697,N_14926,N_14892);
nand UO_698 (O_698,N_14853,N_14816);
nand UO_699 (O_699,N_14984,N_14987);
xnor UO_700 (O_700,N_14855,N_14792);
and UO_701 (O_701,N_14776,N_14720);
nor UO_702 (O_702,N_14907,N_14794);
and UO_703 (O_703,N_14955,N_14793);
xnor UO_704 (O_704,N_14971,N_14954);
nand UO_705 (O_705,N_14716,N_14856);
and UO_706 (O_706,N_14739,N_14982);
and UO_707 (O_707,N_14773,N_14912);
nand UO_708 (O_708,N_14759,N_14776);
xor UO_709 (O_709,N_14837,N_14915);
nor UO_710 (O_710,N_14810,N_14902);
xor UO_711 (O_711,N_14911,N_14904);
nor UO_712 (O_712,N_14771,N_14935);
and UO_713 (O_713,N_14756,N_14943);
or UO_714 (O_714,N_14879,N_14719);
nand UO_715 (O_715,N_14963,N_14983);
xnor UO_716 (O_716,N_14768,N_14864);
or UO_717 (O_717,N_14993,N_14828);
or UO_718 (O_718,N_14723,N_14710);
or UO_719 (O_719,N_14702,N_14728);
and UO_720 (O_720,N_14756,N_14991);
or UO_721 (O_721,N_14990,N_14773);
nor UO_722 (O_722,N_14946,N_14957);
nand UO_723 (O_723,N_14919,N_14835);
or UO_724 (O_724,N_14724,N_14841);
nand UO_725 (O_725,N_14891,N_14776);
and UO_726 (O_726,N_14811,N_14998);
xnor UO_727 (O_727,N_14725,N_14898);
nand UO_728 (O_728,N_14880,N_14903);
or UO_729 (O_729,N_14701,N_14932);
and UO_730 (O_730,N_14783,N_14992);
xnor UO_731 (O_731,N_14733,N_14753);
nor UO_732 (O_732,N_14734,N_14991);
or UO_733 (O_733,N_14915,N_14831);
nor UO_734 (O_734,N_14796,N_14887);
nor UO_735 (O_735,N_14740,N_14825);
xnor UO_736 (O_736,N_14816,N_14701);
or UO_737 (O_737,N_14967,N_14812);
nor UO_738 (O_738,N_14816,N_14846);
xor UO_739 (O_739,N_14805,N_14818);
nor UO_740 (O_740,N_14927,N_14761);
xnor UO_741 (O_741,N_14901,N_14736);
or UO_742 (O_742,N_14968,N_14960);
nor UO_743 (O_743,N_14905,N_14883);
nor UO_744 (O_744,N_14879,N_14774);
or UO_745 (O_745,N_14821,N_14705);
xor UO_746 (O_746,N_14979,N_14812);
nand UO_747 (O_747,N_14981,N_14891);
and UO_748 (O_748,N_14762,N_14722);
and UO_749 (O_749,N_14901,N_14826);
nor UO_750 (O_750,N_14948,N_14881);
or UO_751 (O_751,N_14895,N_14917);
nand UO_752 (O_752,N_14894,N_14901);
xor UO_753 (O_753,N_14744,N_14816);
nor UO_754 (O_754,N_14932,N_14745);
and UO_755 (O_755,N_14802,N_14749);
or UO_756 (O_756,N_14994,N_14934);
and UO_757 (O_757,N_14945,N_14779);
nor UO_758 (O_758,N_14939,N_14946);
or UO_759 (O_759,N_14866,N_14939);
nand UO_760 (O_760,N_14821,N_14898);
or UO_761 (O_761,N_14725,N_14960);
xor UO_762 (O_762,N_14822,N_14710);
xor UO_763 (O_763,N_14749,N_14834);
and UO_764 (O_764,N_14976,N_14919);
nand UO_765 (O_765,N_14800,N_14964);
nor UO_766 (O_766,N_14959,N_14776);
or UO_767 (O_767,N_14995,N_14813);
xor UO_768 (O_768,N_14777,N_14904);
and UO_769 (O_769,N_14759,N_14834);
or UO_770 (O_770,N_14825,N_14940);
and UO_771 (O_771,N_14900,N_14956);
or UO_772 (O_772,N_14753,N_14771);
xnor UO_773 (O_773,N_14727,N_14927);
nor UO_774 (O_774,N_14788,N_14867);
and UO_775 (O_775,N_14942,N_14832);
nor UO_776 (O_776,N_14917,N_14842);
xnor UO_777 (O_777,N_14799,N_14984);
or UO_778 (O_778,N_14784,N_14928);
or UO_779 (O_779,N_14850,N_14861);
nand UO_780 (O_780,N_14761,N_14716);
or UO_781 (O_781,N_14887,N_14722);
nand UO_782 (O_782,N_14867,N_14884);
and UO_783 (O_783,N_14812,N_14987);
xnor UO_784 (O_784,N_14817,N_14809);
xor UO_785 (O_785,N_14739,N_14807);
and UO_786 (O_786,N_14988,N_14986);
or UO_787 (O_787,N_14861,N_14987);
xnor UO_788 (O_788,N_14889,N_14733);
xor UO_789 (O_789,N_14761,N_14914);
nor UO_790 (O_790,N_14706,N_14737);
xor UO_791 (O_791,N_14861,N_14901);
nand UO_792 (O_792,N_14714,N_14864);
xor UO_793 (O_793,N_14718,N_14979);
and UO_794 (O_794,N_14963,N_14775);
and UO_795 (O_795,N_14873,N_14879);
or UO_796 (O_796,N_14806,N_14792);
and UO_797 (O_797,N_14826,N_14903);
and UO_798 (O_798,N_14885,N_14768);
xor UO_799 (O_799,N_14957,N_14714);
or UO_800 (O_800,N_14969,N_14723);
nand UO_801 (O_801,N_14788,N_14713);
and UO_802 (O_802,N_14944,N_14954);
or UO_803 (O_803,N_14769,N_14729);
nor UO_804 (O_804,N_14851,N_14847);
nor UO_805 (O_805,N_14789,N_14749);
nor UO_806 (O_806,N_14769,N_14734);
nand UO_807 (O_807,N_14877,N_14813);
and UO_808 (O_808,N_14906,N_14931);
or UO_809 (O_809,N_14974,N_14916);
nor UO_810 (O_810,N_14949,N_14818);
and UO_811 (O_811,N_14890,N_14818);
nor UO_812 (O_812,N_14859,N_14782);
xor UO_813 (O_813,N_14909,N_14787);
and UO_814 (O_814,N_14953,N_14715);
nand UO_815 (O_815,N_14895,N_14837);
and UO_816 (O_816,N_14861,N_14891);
xnor UO_817 (O_817,N_14758,N_14763);
or UO_818 (O_818,N_14754,N_14898);
xor UO_819 (O_819,N_14983,N_14834);
nand UO_820 (O_820,N_14890,N_14894);
nor UO_821 (O_821,N_14764,N_14812);
nor UO_822 (O_822,N_14972,N_14795);
or UO_823 (O_823,N_14849,N_14845);
nor UO_824 (O_824,N_14789,N_14832);
xor UO_825 (O_825,N_14849,N_14956);
xor UO_826 (O_826,N_14961,N_14897);
xor UO_827 (O_827,N_14714,N_14719);
nor UO_828 (O_828,N_14799,N_14965);
xor UO_829 (O_829,N_14835,N_14861);
nor UO_830 (O_830,N_14719,N_14823);
and UO_831 (O_831,N_14774,N_14954);
nor UO_832 (O_832,N_14720,N_14792);
xnor UO_833 (O_833,N_14909,N_14723);
and UO_834 (O_834,N_14759,N_14908);
nand UO_835 (O_835,N_14930,N_14806);
xor UO_836 (O_836,N_14962,N_14992);
and UO_837 (O_837,N_14755,N_14886);
xor UO_838 (O_838,N_14886,N_14975);
nand UO_839 (O_839,N_14793,N_14919);
nor UO_840 (O_840,N_14771,N_14764);
and UO_841 (O_841,N_14829,N_14915);
xnor UO_842 (O_842,N_14749,N_14763);
or UO_843 (O_843,N_14900,N_14748);
and UO_844 (O_844,N_14729,N_14837);
nor UO_845 (O_845,N_14904,N_14912);
nor UO_846 (O_846,N_14703,N_14911);
nand UO_847 (O_847,N_14787,N_14869);
nand UO_848 (O_848,N_14730,N_14843);
nand UO_849 (O_849,N_14799,N_14986);
xnor UO_850 (O_850,N_14842,N_14918);
nor UO_851 (O_851,N_14926,N_14951);
and UO_852 (O_852,N_14720,N_14745);
or UO_853 (O_853,N_14989,N_14939);
or UO_854 (O_854,N_14853,N_14944);
nor UO_855 (O_855,N_14952,N_14729);
and UO_856 (O_856,N_14819,N_14750);
or UO_857 (O_857,N_14828,N_14776);
and UO_858 (O_858,N_14709,N_14896);
and UO_859 (O_859,N_14986,N_14736);
nand UO_860 (O_860,N_14821,N_14913);
xor UO_861 (O_861,N_14797,N_14745);
xor UO_862 (O_862,N_14709,N_14917);
nor UO_863 (O_863,N_14787,N_14788);
nor UO_864 (O_864,N_14952,N_14794);
and UO_865 (O_865,N_14820,N_14760);
nor UO_866 (O_866,N_14984,N_14875);
xor UO_867 (O_867,N_14704,N_14973);
and UO_868 (O_868,N_14893,N_14910);
and UO_869 (O_869,N_14735,N_14779);
nand UO_870 (O_870,N_14872,N_14916);
or UO_871 (O_871,N_14722,N_14949);
or UO_872 (O_872,N_14810,N_14950);
or UO_873 (O_873,N_14716,N_14887);
and UO_874 (O_874,N_14875,N_14781);
nor UO_875 (O_875,N_14994,N_14865);
and UO_876 (O_876,N_14706,N_14942);
nand UO_877 (O_877,N_14859,N_14872);
nand UO_878 (O_878,N_14949,N_14753);
or UO_879 (O_879,N_14974,N_14886);
xnor UO_880 (O_880,N_14823,N_14709);
or UO_881 (O_881,N_14972,N_14718);
nand UO_882 (O_882,N_14788,N_14905);
nor UO_883 (O_883,N_14935,N_14815);
nand UO_884 (O_884,N_14791,N_14819);
and UO_885 (O_885,N_14795,N_14755);
or UO_886 (O_886,N_14880,N_14762);
nor UO_887 (O_887,N_14704,N_14937);
and UO_888 (O_888,N_14838,N_14869);
or UO_889 (O_889,N_14947,N_14756);
or UO_890 (O_890,N_14813,N_14828);
xnor UO_891 (O_891,N_14992,N_14928);
nand UO_892 (O_892,N_14831,N_14753);
nand UO_893 (O_893,N_14861,N_14932);
or UO_894 (O_894,N_14710,N_14939);
xnor UO_895 (O_895,N_14954,N_14848);
nand UO_896 (O_896,N_14869,N_14984);
and UO_897 (O_897,N_14980,N_14713);
xnor UO_898 (O_898,N_14859,N_14792);
or UO_899 (O_899,N_14816,N_14742);
nand UO_900 (O_900,N_14817,N_14766);
or UO_901 (O_901,N_14773,N_14705);
nand UO_902 (O_902,N_14791,N_14718);
and UO_903 (O_903,N_14864,N_14771);
nor UO_904 (O_904,N_14932,N_14892);
xor UO_905 (O_905,N_14881,N_14958);
nor UO_906 (O_906,N_14869,N_14839);
nand UO_907 (O_907,N_14724,N_14929);
or UO_908 (O_908,N_14794,N_14789);
or UO_909 (O_909,N_14963,N_14929);
or UO_910 (O_910,N_14785,N_14820);
nor UO_911 (O_911,N_14787,N_14710);
nand UO_912 (O_912,N_14907,N_14848);
nor UO_913 (O_913,N_14776,N_14857);
or UO_914 (O_914,N_14955,N_14852);
or UO_915 (O_915,N_14806,N_14882);
or UO_916 (O_916,N_14783,N_14996);
xnor UO_917 (O_917,N_14891,N_14780);
nand UO_918 (O_918,N_14936,N_14986);
or UO_919 (O_919,N_14801,N_14932);
or UO_920 (O_920,N_14982,N_14885);
nor UO_921 (O_921,N_14730,N_14807);
xor UO_922 (O_922,N_14912,N_14873);
nand UO_923 (O_923,N_14946,N_14977);
nand UO_924 (O_924,N_14709,N_14979);
or UO_925 (O_925,N_14795,N_14781);
xnor UO_926 (O_926,N_14704,N_14979);
nand UO_927 (O_927,N_14904,N_14812);
and UO_928 (O_928,N_14945,N_14771);
or UO_929 (O_929,N_14979,N_14859);
nand UO_930 (O_930,N_14830,N_14958);
nand UO_931 (O_931,N_14775,N_14845);
nor UO_932 (O_932,N_14778,N_14872);
and UO_933 (O_933,N_14730,N_14849);
nor UO_934 (O_934,N_14938,N_14937);
xnor UO_935 (O_935,N_14890,N_14946);
and UO_936 (O_936,N_14744,N_14735);
xnor UO_937 (O_937,N_14710,N_14729);
nand UO_938 (O_938,N_14798,N_14727);
xnor UO_939 (O_939,N_14852,N_14896);
xnor UO_940 (O_940,N_14710,N_14915);
xor UO_941 (O_941,N_14716,N_14806);
nor UO_942 (O_942,N_14793,N_14958);
nand UO_943 (O_943,N_14713,N_14939);
or UO_944 (O_944,N_14766,N_14936);
xnor UO_945 (O_945,N_14946,N_14891);
nor UO_946 (O_946,N_14858,N_14730);
or UO_947 (O_947,N_14854,N_14827);
or UO_948 (O_948,N_14760,N_14881);
nor UO_949 (O_949,N_14801,N_14956);
xnor UO_950 (O_950,N_14865,N_14793);
nand UO_951 (O_951,N_14745,N_14905);
nand UO_952 (O_952,N_14752,N_14757);
or UO_953 (O_953,N_14928,N_14783);
or UO_954 (O_954,N_14797,N_14841);
and UO_955 (O_955,N_14732,N_14935);
or UO_956 (O_956,N_14949,N_14790);
nand UO_957 (O_957,N_14865,N_14808);
and UO_958 (O_958,N_14799,N_14954);
nor UO_959 (O_959,N_14901,N_14731);
xnor UO_960 (O_960,N_14837,N_14830);
xor UO_961 (O_961,N_14737,N_14742);
nor UO_962 (O_962,N_14870,N_14933);
xor UO_963 (O_963,N_14720,N_14897);
or UO_964 (O_964,N_14877,N_14710);
or UO_965 (O_965,N_14700,N_14929);
or UO_966 (O_966,N_14964,N_14857);
nor UO_967 (O_967,N_14854,N_14855);
and UO_968 (O_968,N_14809,N_14927);
or UO_969 (O_969,N_14939,N_14928);
or UO_970 (O_970,N_14724,N_14800);
or UO_971 (O_971,N_14797,N_14977);
xnor UO_972 (O_972,N_14924,N_14796);
nand UO_973 (O_973,N_14912,N_14808);
nor UO_974 (O_974,N_14709,N_14986);
xor UO_975 (O_975,N_14832,N_14835);
and UO_976 (O_976,N_14705,N_14846);
nand UO_977 (O_977,N_14760,N_14823);
nand UO_978 (O_978,N_14875,N_14849);
xor UO_979 (O_979,N_14778,N_14818);
xnor UO_980 (O_980,N_14866,N_14872);
nand UO_981 (O_981,N_14989,N_14986);
xor UO_982 (O_982,N_14735,N_14990);
xor UO_983 (O_983,N_14989,N_14909);
xnor UO_984 (O_984,N_14985,N_14998);
xor UO_985 (O_985,N_14982,N_14967);
and UO_986 (O_986,N_14729,N_14782);
or UO_987 (O_987,N_14972,N_14883);
and UO_988 (O_988,N_14993,N_14952);
or UO_989 (O_989,N_14782,N_14893);
nand UO_990 (O_990,N_14961,N_14814);
nor UO_991 (O_991,N_14704,N_14932);
or UO_992 (O_992,N_14707,N_14797);
xnor UO_993 (O_993,N_14882,N_14935);
xor UO_994 (O_994,N_14912,N_14870);
or UO_995 (O_995,N_14757,N_14923);
nor UO_996 (O_996,N_14759,N_14906);
nand UO_997 (O_997,N_14867,N_14791);
xor UO_998 (O_998,N_14984,N_14913);
nand UO_999 (O_999,N_14783,N_14819);
nor UO_1000 (O_1000,N_14884,N_14895);
or UO_1001 (O_1001,N_14981,N_14906);
and UO_1002 (O_1002,N_14871,N_14918);
xor UO_1003 (O_1003,N_14787,N_14799);
or UO_1004 (O_1004,N_14936,N_14900);
xor UO_1005 (O_1005,N_14883,N_14970);
xor UO_1006 (O_1006,N_14828,N_14921);
nand UO_1007 (O_1007,N_14854,N_14799);
nand UO_1008 (O_1008,N_14821,N_14967);
and UO_1009 (O_1009,N_14709,N_14799);
and UO_1010 (O_1010,N_14839,N_14993);
xnor UO_1011 (O_1011,N_14763,N_14995);
or UO_1012 (O_1012,N_14892,N_14964);
or UO_1013 (O_1013,N_14930,N_14887);
nor UO_1014 (O_1014,N_14877,N_14733);
xnor UO_1015 (O_1015,N_14750,N_14841);
or UO_1016 (O_1016,N_14833,N_14723);
xor UO_1017 (O_1017,N_14890,N_14830);
or UO_1018 (O_1018,N_14914,N_14804);
nand UO_1019 (O_1019,N_14988,N_14984);
nand UO_1020 (O_1020,N_14731,N_14899);
or UO_1021 (O_1021,N_14771,N_14955);
and UO_1022 (O_1022,N_14904,N_14735);
nand UO_1023 (O_1023,N_14811,N_14793);
nor UO_1024 (O_1024,N_14736,N_14735);
and UO_1025 (O_1025,N_14736,N_14932);
nor UO_1026 (O_1026,N_14814,N_14891);
or UO_1027 (O_1027,N_14808,N_14846);
or UO_1028 (O_1028,N_14860,N_14949);
or UO_1029 (O_1029,N_14778,N_14809);
or UO_1030 (O_1030,N_14914,N_14747);
xor UO_1031 (O_1031,N_14706,N_14783);
or UO_1032 (O_1032,N_14940,N_14923);
xor UO_1033 (O_1033,N_14790,N_14834);
and UO_1034 (O_1034,N_14874,N_14738);
xnor UO_1035 (O_1035,N_14914,N_14986);
nand UO_1036 (O_1036,N_14709,N_14996);
nand UO_1037 (O_1037,N_14866,N_14982);
and UO_1038 (O_1038,N_14995,N_14992);
or UO_1039 (O_1039,N_14955,N_14759);
nand UO_1040 (O_1040,N_14788,N_14844);
or UO_1041 (O_1041,N_14963,N_14996);
and UO_1042 (O_1042,N_14819,N_14910);
nor UO_1043 (O_1043,N_14718,N_14878);
xor UO_1044 (O_1044,N_14714,N_14828);
xor UO_1045 (O_1045,N_14843,N_14738);
nor UO_1046 (O_1046,N_14964,N_14879);
or UO_1047 (O_1047,N_14901,N_14750);
nand UO_1048 (O_1048,N_14961,N_14755);
xnor UO_1049 (O_1049,N_14839,N_14866);
and UO_1050 (O_1050,N_14984,N_14704);
xor UO_1051 (O_1051,N_14769,N_14959);
and UO_1052 (O_1052,N_14836,N_14900);
nor UO_1053 (O_1053,N_14900,N_14950);
or UO_1054 (O_1054,N_14829,N_14710);
nand UO_1055 (O_1055,N_14953,N_14891);
xnor UO_1056 (O_1056,N_14716,N_14840);
xnor UO_1057 (O_1057,N_14805,N_14861);
or UO_1058 (O_1058,N_14916,N_14752);
xor UO_1059 (O_1059,N_14946,N_14920);
nor UO_1060 (O_1060,N_14783,N_14748);
nor UO_1061 (O_1061,N_14954,N_14877);
nand UO_1062 (O_1062,N_14967,N_14920);
xor UO_1063 (O_1063,N_14975,N_14780);
and UO_1064 (O_1064,N_14742,N_14919);
nor UO_1065 (O_1065,N_14889,N_14735);
nor UO_1066 (O_1066,N_14988,N_14755);
or UO_1067 (O_1067,N_14941,N_14862);
and UO_1068 (O_1068,N_14852,N_14760);
nor UO_1069 (O_1069,N_14840,N_14842);
or UO_1070 (O_1070,N_14977,N_14778);
nand UO_1071 (O_1071,N_14721,N_14937);
and UO_1072 (O_1072,N_14801,N_14727);
nand UO_1073 (O_1073,N_14894,N_14914);
and UO_1074 (O_1074,N_14854,N_14871);
xor UO_1075 (O_1075,N_14758,N_14811);
xnor UO_1076 (O_1076,N_14706,N_14888);
nor UO_1077 (O_1077,N_14754,N_14914);
nor UO_1078 (O_1078,N_14930,N_14788);
or UO_1079 (O_1079,N_14801,N_14861);
nor UO_1080 (O_1080,N_14840,N_14993);
or UO_1081 (O_1081,N_14828,N_14818);
or UO_1082 (O_1082,N_14709,N_14946);
nand UO_1083 (O_1083,N_14966,N_14818);
nand UO_1084 (O_1084,N_14965,N_14933);
or UO_1085 (O_1085,N_14901,N_14979);
or UO_1086 (O_1086,N_14931,N_14928);
and UO_1087 (O_1087,N_14706,N_14810);
nand UO_1088 (O_1088,N_14857,N_14933);
or UO_1089 (O_1089,N_14723,N_14876);
nor UO_1090 (O_1090,N_14810,N_14806);
or UO_1091 (O_1091,N_14922,N_14826);
and UO_1092 (O_1092,N_14949,N_14825);
nor UO_1093 (O_1093,N_14997,N_14979);
or UO_1094 (O_1094,N_14860,N_14749);
and UO_1095 (O_1095,N_14880,N_14980);
nor UO_1096 (O_1096,N_14941,N_14939);
xnor UO_1097 (O_1097,N_14894,N_14875);
and UO_1098 (O_1098,N_14909,N_14886);
xor UO_1099 (O_1099,N_14955,N_14937);
xor UO_1100 (O_1100,N_14833,N_14955);
nor UO_1101 (O_1101,N_14792,N_14893);
nand UO_1102 (O_1102,N_14880,N_14736);
xor UO_1103 (O_1103,N_14911,N_14753);
nand UO_1104 (O_1104,N_14910,N_14838);
or UO_1105 (O_1105,N_14932,N_14769);
xnor UO_1106 (O_1106,N_14782,N_14708);
xor UO_1107 (O_1107,N_14897,N_14729);
and UO_1108 (O_1108,N_14994,N_14792);
and UO_1109 (O_1109,N_14805,N_14764);
or UO_1110 (O_1110,N_14968,N_14941);
nor UO_1111 (O_1111,N_14804,N_14781);
and UO_1112 (O_1112,N_14951,N_14868);
and UO_1113 (O_1113,N_14933,N_14765);
nor UO_1114 (O_1114,N_14831,N_14748);
nand UO_1115 (O_1115,N_14852,N_14923);
and UO_1116 (O_1116,N_14874,N_14823);
and UO_1117 (O_1117,N_14900,N_14928);
nor UO_1118 (O_1118,N_14700,N_14953);
nand UO_1119 (O_1119,N_14868,N_14942);
xor UO_1120 (O_1120,N_14941,N_14997);
or UO_1121 (O_1121,N_14721,N_14805);
and UO_1122 (O_1122,N_14708,N_14756);
xor UO_1123 (O_1123,N_14785,N_14838);
and UO_1124 (O_1124,N_14935,N_14876);
nand UO_1125 (O_1125,N_14910,N_14829);
or UO_1126 (O_1126,N_14969,N_14995);
xnor UO_1127 (O_1127,N_14999,N_14831);
nand UO_1128 (O_1128,N_14776,N_14847);
xor UO_1129 (O_1129,N_14805,N_14704);
and UO_1130 (O_1130,N_14982,N_14765);
nor UO_1131 (O_1131,N_14907,N_14727);
nand UO_1132 (O_1132,N_14879,N_14826);
xnor UO_1133 (O_1133,N_14994,N_14749);
nor UO_1134 (O_1134,N_14970,N_14769);
and UO_1135 (O_1135,N_14857,N_14878);
xor UO_1136 (O_1136,N_14910,N_14877);
xor UO_1137 (O_1137,N_14779,N_14823);
and UO_1138 (O_1138,N_14848,N_14720);
nand UO_1139 (O_1139,N_14964,N_14815);
or UO_1140 (O_1140,N_14759,N_14844);
xor UO_1141 (O_1141,N_14743,N_14750);
xnor UO_1142 (O_1142,N_14757,N_14897);
and UO_1143 (O_1143,N_14713,N_14919);
xnor UO_1144 (O_1144,N_14761,N_14794);
nor UO_1145 (O_1145,N_14935,N_14863);
xor UO_1146 (O_1146,N_14720,N_14968);
nand UO_1147 (O_1147,N_14838,N_14806);
or UO_1148 (O_1148,N_14804,N_14965);
nand UO_1149 (O_1149,N_14809,N_14715);
xor UO_1150 (O_1150,N_14813,N_14888);
nand UO_1151 (O_1151,N_14789,N_14973);
nand UO_1152 (O_1152,N_14803,N_14985);
or UO_1153 (O_1153,N_14981,N_14728);
xor UO_1154 (O_1154,N_14896,N_14850);
xor UO_1155 (O_1155,N_14911,N_14831);
xnor UO_1156 (O_1156,N_14948,N_14819);
nor UO_1157 (O_1157,N_14833,N_14917);
nand UO_1158 (O_1158,N_14922,N_14768);
nor UO_1159 (O_1159,N_14966,N_14888);
or UO_1160 (O_1160,N_14869,N_14973);
nand UO_1161 (O_1161,N_14925,N_14977);
and UO_1162 (O_1162,N_14908,N_14992);
and UO_1163 (O_1163,N_14770,N_14976);
or UO_1164 (O_1164,N_14941,N_14837);
nand UO_1165 (O_1165,N_14769,N_14773);
xnor UO_1166 (O_1166,N_14891,N_14769);
and UO_1167 (O_1167,N_14969,N_14990);
nand UO_1168 (O_1168,N_14829,N_14888);
xor UO_1169 (O_1169,N_14703,N_14888);
or UO_1170 (O_1170,N_14857,N_14904);
xnor UO_1171 (O_1171,N_14909,N_14862);
and UO_1172 (O_1172,N_14796,N_14733);
nor UO_1173 (O_1173,N_14733,N_14898);
xnor UO_1174 (O_1174,N_14935,N_14930);
or UO_1175 (O_1175,N_14707,N_14774);
xnor UO_1176 (O_1176,N_14820,N_14779);
and UO_1177 (O_1177,N_14880,N_14877);
xnor UO_1178 (O_1178,N_14840,N_14949);
and UO_1179 (O_1179,N_14852,N_14818);
and UO_1180 (O_1180,N_14833,N_14819);
or UO_1181 (O_1181,N_14996,N_14901);
xnor UO_1182 (O_1182,N_14996,N_14924);
or UO_1183 (O_1183,N_14739,N_14937);
nand UO_1184 (O_1184,N_14796,N_14867);
or UO_1185 (O_1185,N_14742,N_14850);
or UO_1186 (O_1186,N_14723,N_14997);
or UO_1187 (O_1187,N_14868,N_14710);
xnor UO_1188 (O_1188,N_14859,N_14812);
or UO_1189 (O_1189,N_14880,N_14775);
and UO_1190 (O_1190,N_14882,N_14737);
nor UO_1191 (O_1191,N_14773,N_14994);
nand UO_1192 (O_1192,N_14820,N_14788);
nand UO_1193 (O_1193,N_14985,N_14715);
nand UO_1194 (O_1194,N_14985,N_14989);
xnor UO_1195 (O_1195,N_14931,N_14868);
nand UO_1196 (O_1196,N_14736,N_14935);
xnor UO_1197 (O_1197,N_14789,N_14919);
and UO_1198 (O_1198,N_14733,N_14901);
and UO_1199 (O_1199,N_14797,N_14916);
xnor UO_1200 (O_1200,N_14991,N_14841);
xor UO_1201 (O_1201,N_14789,N_14904);
nor UO_1202 (O_1202,N_14980,N_14883);
nor UO_1203 (O_1203,N_14963,N_14734);
or UO_1204 (O_1204,N_14746,N_14757);
or UO_1205 (O_1205,N_14739,N_14942);
and UO_1206 (O_1206,N_14855,N_14852);
xor UO_1207 (O_1207,N_14738,N_14806);
and UO_1208 (O_1208,N_14801,N_14775);
and UO_1209 (O_1209,N_14792,N_14910);
and UO_1210 (O_1210,N_14884,N_14892);
nand UO_1211 (O_1211,N_14926,N_14780);
nor UO_1212 (O_1212,N_14729,N_14964);
nand UO_1213 (O_1213,N_14890,N_14889);
xnor UO_1214 (O_1214,N_14791,N_14704);
xor UO_1215 (O_1215,N_14870,N_14840);
and UO_1216 (O_1216,N_14764,N_14782);
or UO_1217 (O_1217,N_14851,N_14753);
or UO_1218 (O_1218,N_14769,N_14853);
and UO_1219 (O_1219,N_14887,N_14815);
nor UO_1220 (O_1220,N_14706,N_14913);
xor UO_1221 (O_1221,N_14887,N_14973);
or UO_1222 (O_1222,N_14811,N_14897);
nor UO_1223 (O_1223,N_14786,N_14943);
nor UO_1224 (O_1224,N_14847,N_14988);
or UO_1225 (O_1225,N_14709,N_14900);
xnor UO_1226 (O_1226,N_14766,N_14920);
and UO_1227 (O_1227,N_14754,N_14763);
and UO_1228 (O_1228,N_14947,N_14894);
nor UO_1229 (O_1229,N_14874,N_14810);
or UO_1230 (O_1230,N_14762,N_14750);
xnor UO_1231 (O_1231,N_14813,N_14814);
or UO_1232 (O_1232,N_14891,N_14898);
xor UO_1233 (O_1233,N_14809,N_14782);
nand UO_1234 (O_1234,N_14727,N_14874);
nand UO_1235 (O_1235,N_14874,N_14994);
or UO_1236 (O_1236,N_14942,N_14966);
or UO_1237 (O_1237,N_14801,N_14766);
xor UO_1238 (O_1238,N_14820,N_14834);
nor UO_1239 (O_1239,N_14809,N_14714);
xnor UO_1240 (O_1240,N_14803,N_14865);
xnor UO_1241 (O_1241,N_14909,N_14902);
or UO_1242 (O_1242,N_14856,N_14902);
xor UO_1243 (O_1243,N_14711,N_14735);
xnor UO_1244 (O_1244,N_14793,N_14810);
nor UO_1245 (O_1245,N_14891,N_14979);
nand UO_1246 (O_1246,N_14910,N_14807);
xnor UO_1247 (O_1247,N_14712,N_14744);
xnor UO_1248 (O_1248,N_14935,N_14826);
nor UO_1249 (O_1249,N_14912,N_14977);
nor UO_1250 (O_1250,N_14870,N_14996);
and UO_1251 (O_1251,N_14956,N_14996);
nand UO_1252 (O_1252,N_14738,N_14814);
nand UO_1253 (O_1253,N_14816,N_14996);
xor UO_1254 (O_1254,N_14705,N_14804);
nand UO_1255 (O_1255,N_14904,N_14991);
nor UO_1256 (O_1256,N_14756,N_14867);
and UO_1257 (O_1257,N_14794,N_14730);
or UO_1258 (O_1258,N_14996,N_14926);
or UO_1259 (O_1259,N_14857,N_14951);
and UO_1260 (O_1260,N_14892,N_14912);
nor UO_1261 (O_1261,N_14797,N_14831);
nand UO_1262 (O_1262,N_14781,N_14980);
nand UO_1263 (O_1263,N_14844,N_14839);
nand UO_1264 (O_1264,N_14951,N_14874);
or UO_1265 (O_1265,N_14760,N_14887);
and UO_1266 (O_1266,N_14755,N_14722);
nand UO_1267 (O_1267,N_14877,N_14937);
nor UO_1268 (O_1268,N_14787,N_14823);
nor UO_1269 (O_1269,N_14747,N_14944);
nand UO_1270 (O_1270,N_14819,N_14765);
nand UO_1271 (O_1271,N_14893,N_14798);
nor UO_1272 (O_1272,N_14986,N_14779);
and UO_1273 (O_1273,N_14973,N_14969);
nand UO_1274 (O_1274,N_14864,N_14755);
nand UO_1275 (O_1275,N_14912,N_14954);
and UO_1276 (O_1276,N_14891,N_14937);
nand UO_1277 (O_1277,N_14785,N_14987);
nand UO_1278 (O_1278,N_14850,N_14817);
or UO_1279 (O_1279,N_14862,N_14940);
nand UO_1280 (O_1280,N_14777,N_14786);
or UO_1281 (O_1281,N_14872,N_14790);
or UO_1282 (O_1282,N_14805,N_14951);
nor UO_1283 (O_1283,N_14746,N_14812);
nand UO_1284 (O_1284,N_14961,N_14715);
and UO_1285 (O_1285,N_14787,N_14930);
nor UO_1286 (O_1286,N_14899,N_14874);
or UO_1287 (O_1287,N_14846,N_14776);
xor UO_1288 (O_1288,N_14970,N_14989);
nand UO_1289 (O_1289,N_14852,N_14794);
xnor UO_1290 (O_1290,N_14785,N_14832);
xor UO_1291 (O_1291,N_14745,N_14869);
and UO_1292 (O_1292,N_14849,N_14799);
xor UO_1293 (O_1293,N_14707,N_14783);
nor UO_1294 (O_1294,N_14851,N_14968);
and UO_1295 (O_1295,N_14745,N_14703);
xnor UO_1296 (O_1296,N_14726,N_14771);
or UO_1297 (O_1297,N_14740,N_14822);
xor UO_1298 (O_1298,N_14941,N_14912);
and UO_1299 (O_1299,N_14786,N_14845);
or UO_1300 (O_1300,N_14710,N_14795);
nand UO_1301 (O_1301,N_14959,N_14889);
nand UO_1302 (O_1302,N_14828,N_14943);
or UO_1303 (O_1303,N_14826,N_14857);
xnor UO_1304 (O_1304,N_14941,N_14789);
xnor UO_1305 (O_1305,N_14891,N_14850);
or UO_1306 (O_1306,N_14965,N_14975);
xor UO_1307 (O_1307,N_14824,N_14983);
nand UO_1308 (O_1308,N_14918,N_14966);
nor UO_1309 (O_1309,N_14807,N_14963);
and UO_1310 (O_1310,N_14800,N_14796);
xnor UO_1311 (O_1311,N_14965,N_14783);
or UO_1312 (O_1312,N_14976,N_14803);
and UO_1313 (O_1313,N_14966,N_14789);
or UO_1314 (O_1314,N_14782,N_14986);
nor UO_1315 (O_1315,N_14827,N_14819);
nor UO_1316 (O_1316,N_14868,N_14997);
nor UO_1317 (O_1317,N_14967,N_14956);
or UO_1318 (O_1318,N_14738,N_14803);
or UO_1319 (O_1319,N_14966,N_14708);
xor UO_1320 (O_1320,N_14724,N_14931);
xnor UO_1321 (O_1321,N_14717,N_14814);
nor UO_1322 (O_1322,N_14703,N_14922);
nand UO_1323 (O_1323,N_14705,N_14780);
and UO_1324 (O_1324,N_14947,N_14716);
nor UO_1325 (O_1325,N_14862,N_14938);
xor UO_1326 (O_1326,N_14762,N_14729);
and UO_1327 (O_1327,N_14724,N_14778);
xnor UO_1328 (O_1328,N_14917,N_14996);
and UO_1329 (O_1329,N_14904,N_14958);
nor UO_1330 (O_1330,N_14795,N_14737);
nand UO_1331 (O_1331,N_14834,N_14730);
or UO_1332 (O_1332,N_14875,N_14930);
nand UO_1333 (O_1333,N_14736,N_14729);
or UO_1334 (O_1334,N_14837,N_14755);
xnor UO_1335 (O_1335,N_14765,N_14873);
and UO_1336 (O_1336,N_14721,N_14904);
or UO_1337 (O_1337,N_14948,N_14835);
nand UO_1338 (O_1338,N_14852,N_14806);
and UO_1339 (O_1339,N_14742,N_14998);
nor UO_1340 (O_1340,N_14882,N_14766);
xnor UO_1341 (O_1341,N_14752,N_14801);
and UO_1342 (O_1342,N_14986,N_14974);
nor UO_1343 (O_1343,N_14873,N_14981);
or UO_1344 (O_1344,N_14766,N_14945);
xnor UO_1345 (O_1345,N_14749,N_14787);
nor UO_1346 (O_1346,N_14966,N_14996);
nor UO_1347 (O_1347,N_14973,N_14765);
xor UO_1348 (O_1348,N_14867,N_14975);
nor UO_1349 (O_1349,N_14862,N_14960);
xnor UO_1350 (O_1350,N_14827,N_14768);
xor UO_1351 (O_1351,N_14829,N_14796);
or UO_1352 (O_1352,N_14914,N_14980);
nor UO_1353 (O_1353,N_14956,N_14763);
nor UO_1354 (O_1354,N_14750,N_14842);
xor UO_1355 (O_1355,N_14751,N_14934);
and UO_1356 (O_1356,N_14981,N_14970);
nand UO_1357 (O_1357,N_14996,N_14875);
and UO_1358 (O_1358,N_14723,N_14714);
or UO_1359 (O_1359,N_14705,N_14934);
xnor UO_1360 (O_1360,N_14838,N_14963);
nor UO_1361 (O_1361,N_14892,N_14814);
nand UO_1362 (O_1362,N_14837,N_14726);
nor UO_1363 (O_1363,N_14985,N_14797);
nor UO_1364 (O_1364,N_14749,N_14980);
xor UO_1365 (O_1365,N_14757,N_14726);
and UO_1366 (O_1366,N_14871,N_14922);
nand UO_1367 (O_1367,N_14733,N_14730);
nand UO_1368 (O_1368,N_14720,N_14733);
nand UO_1369 (O_1369,N_14858,N_14701);
and UO_1370 (O_1370,N_14980,N_14978);
nor UO_1371 (O_1371,N_14965,N_14709);
or UO_1372 (O_1372,N_14804,N_14783);
or UO_1373 (O_1373,N_14929,N_14835);
or UO_1374 (O_1374,N_14980,N_14761);
or UO_1375 (O_1375,N_14950,N_14813);
or UO_1376 (O_1376,N_14830,N_14925);
nand UO_1377 (O_1377,N_14978,N_14811);
and UO_1378 (O_1378,N_14986,N_14795);
nand UO_1379 (O_1379,N_14992,N_14768);
and UO_1380 (O_1380,N_14975,N_14703);
xnor UO_1381 (O_1381,N_14813,N_14826);
nor UO_1382 (O_1382,N_14821,N_14816);
or UO_1383 (O_1383,N_14763,N_14797);
or UO_1384 (O_1384,N_14737,N_14802);
and UO_1385 (O_1385,N_14877,N_14757);
xnor UO_1386 (O_1386,N_14936,N_14926);
or UO_1387 (O_1387,N_14833,N_14781);
xnor UO_1388 (O_1388,N_14748,N_14947);
or UO_1389 (O_1389,N_14786,N_14976);
nand UO_1390 (O_1390,N_14704,N_14701);
and UO_1391 (O_1391,N_14903,N_14908);
and UO_1392 (O_1392,N_14953,N_14751);
nand UO_1393 (O_1393,N_14768,N_14890);
nor UO_1394 (O_1394,N_14781,N_14919);
and UO_1395 (O_1395,N_14706,N_14953);
or UO_1396 (O_1396,N_14909,N_14969);
nor UO_1397 (O_1397,N_14967,N_14997);
and UO_1398 (O_1398,N_14705,N_14771);
or UO_1399 (O_1399,N_14753,N_14916);
nor UO_1400 (O_1400,N_14849,N_14877);
xor UO_1401 (O_1401,N_14844,N_14972);
and UO_1402 (O_1402,N_14879,N_14885);
xor UO_1403 (O_1403,N_14795,N_14808);
nand UO_1404 (O_1404,N_14801,N_14877);
or UO_1405 (O_1405,N_14767,N_14818);
xor UO_1406 (O_1406,N_14831,N_14779);
xor UO_1407 (O_1407,N_14909,N_14795);
nand UO_1408 (O_1408,N_14778,N_14717);
nor UO_1409 (O_1409,N_14786,N_14955);
or UO_1410 (O_1410,N_14829,N_14972);
nor UO_1411 (O_1411,N_14751,N_14795);
or UO_1412 (O_1412,N_14743,N_14704);
nand UO_1413 (O_1413,N_14879,N_14781);
nand UO_1414 (O_1414,N_14963,N_14945);
or UO_1415 (O_1415,N_14962,N_14787);
xnor UO_1416 (O_1416,N_14730,N_14931);
xnor UO_1417 (O_1417,N_14711,N_14890);
xnor UO_1418 (O_1418,N_14994,N_14956);
or UO_1419 (O_1419,N_14749,N_14970);
xor UO_1420 (O_1420,N_14919,N_14788);
and UO_1421 (O_1421,N_14978,N_14873);
or UO_1422 (O_1422,N_14928,N_14851);
or UO_1423 (O_1423,N_14847,N_14957);
and UO_1424 (O_1424,N_14831,N_14771);
or UO_1425 (O_1425,N_14925,N_14814);
or UO_1426 (O_1426,N_14851,N_14830);
or UO_1427 (O_1427,N_14712,N_14840);
nor UO_1428 (O_1428,N_14816,N_14961);
and UO_1429 (O_1429,N_14833,N_14887);
xor UO_1430 (O_1430,N_14866,N_14980);
or UO_1431 (O_1431,N_14873,N_14896);
or UO_1432 (O_1432,N_14894,N_14904);
nor UO_1433 (O_1433,N_14987,N_14875);
or UO_1434 (O_1434,N_14934,N_14961);
nand UO_1435 (O_1435,N_14727,N_14714);
and UO_1436 (O_1436,N_14937,N_14788);
xnor UO_1437 (O_1437,N_14724,N_14716);
xor UO_1438 (O_1438,N_14714,N_14852);
xor UO_1439 (O_1439,N_14757,N_14711);
xor UO_1440 (O_1440,N_14706,N_14859);
xnor UO_1441 (O_1441,N_14737,N_14919);
xnor UO_1442 (O_1442,N_14819,N_14939);
nor UO_1443 (O_1443,N_14752,N_14959);
nand UO_1444 (O_1444,N_14786,N_14873);
xnor UO_1445 (O_1445,N_14835,N_14816);
or UO_1446 (O_1446,N_14833,N_14829);
nand UO_1447 (O_1447,N_14884,N_14918);
nor UO_1448 (O_1448,N_14801,N_14867);
and UO_1449 (O_1449,N_14985,N_14759);
and UO_1450 (O_1450,N_14778,N_14960);
and UO_1451 (O_1451,N_14756,N_14738);
or UO_1452 (O_1452,N_14740,N_14929);
and UO_1453 (O_1453,N_14808,N_14869);
and UO_1454 (O_1454,N_14962,N_14765);
nor UO_1455 (O_1455,N_14968,N_14759);
xnor UO_1456 (O_1456,N_14745,N_14996);
xnor UO_1457 (O_1457,N_14765,N_14835);
nor UO_1458 (O_1458,N_14930,N_14997);
nor UO_1459 (O_1459,N_14816,N_14916);
or UO_1460 (O_1460,N_14770,N_14780);
xor UO_1461 (O_1461,N_14950,N_14888);
xnor UO_1462 (O_1462,N_14982,N_14839);
nor UO_1463 (O_1463,N_14982,N_14773);
or UO_1464 (O_1464,N_14744,N_14844);
nor UO_1465 (O_1465,N_14721,N_14903);
and UO_1466 (O_1466,N_14987,N_14793);
nand UO_1467 (O_1467,N_14845,N_14811);
xor UO_1468 (O_1468,N_14745,N_14757);
or UO_1469 (O_1469,N_14807,N_14708);
nand UO_1470 (O_1470,N_14791,N_14725);
nor UO_1471 (O_1471,N_14826,N_14989);
xnor UO_1472 (O_1472,N_14869,N_14812);
nor UO_1473 (O_1473,N_14900,N_14708);
and UO_1474 (O_1474,N_14810,N_14882);
or UO_1475 (O_1475,N_14870,N_14987);
xnor UO_1476 (O_1476,N_14804,N_14888);
xnor UO_1477 (O_1477,N_14758,N_14719);
xor UO_1478 (O_1478,N_14996,N_14777);
nand UO_1479 (O_1479,N_14811,N_14883);
and UO_1480 (O_1480,N_14909,N_14861);
xnor UO_1481 (O_1481,N_14738,N_14932);
nor UO_1482 (O_1482,N_14874,N_14950);
or UO_1483 (O_1483,N_14751,N_14711);
and UO_1484 (O_1484,N_14729,N_14997);
nand UO_1485 (O_1485,N_14785,N_14978);
nor UO_1486 (O_1486,N_14746,N_14821);
xnor UO_1487 (O_1487,N_14833,N_14756);
nand UO_1488 (O_1488,N_14958,N_14806);
or UO_1489 (O_1489,N_14788,N_14750);
or UO_1490 (O_1490,N_14992,N_14986);
nor UO_1491 (O_1491,N_14785,N_14796);
nand UO_1492 (O_1492,N_14834,N_14770);
nand UO_1493 (O_1493,N_14806,N_14935);
or UO_1494 (O_1494,N_14936,N_14839);
and UO_1495 (O_1495,N_14858,N_14953);
or UO_1496 (O_1496,N_14838,N_14911);
nor UO_1497 (O_1497,N_14976,N_14764);
nand UO_1498 (O_1498,N_14895,N_14725);
nor UO_1499 (O_1499,N_14901,N_14963);
or UO_1500 (O_1500,N_14849,N_14916);
xnor UO_1501 (O_1501,N_14771,N_14773);
and UO_1502 (O_1502,N_14858,N_14777);
nand UO_1503 (O_1503,N_14718,N_14931);
nand UO_1504 (O_1504,N_14986,N_14828);
xor UO_1505 (O_1505,N_14940,N_14876);
or UO_1506 (O_1506,N_14835,N_14746);
and UO_1507 (O_1507,N_14945,N_14795);
xor UO_1508 (O_1508,N_14908,N_14912);
and UO_1509 (O_1509,N_14825,N_14795);
nor UO_1510 (O_1510,N_14962,N_14840);
nand UO_1511 (O_1511,N_14931,N_14741);
nor UO_1512 (O_1512,N_14737,N_14790);
or UO_1513 (O_1513,N_14842,N_14746);
or UO_1514 (O_1514,N_14907,N_14935);
nand UO_1515 (O_1515,N_14972,N_14833);
nor UO_1516 (O_1516,N_14716,N_14986);
nand UO_1517 (O_1517,N_14701,N_14755);
nand UO_1518 (O_1518,N_14821,N_14743);
nand UO_1519 (O_1519,N_14792,N_14812);
or UO_1520 (O_1520,N_14736,N_14987);
or UO_1521 (O_1521,N_14841,N_14845);
xnor UO_1522 (O_1522,N_14950,N_14898);
or UO_1523 (O_1523,N_14839,N_14872);
or UO_1524 (O_1524,N_14906,N_14925);
nand UO_1525 (O_1525,N_14717,N_14866);
xnor UO_1526 (O_1526,N_14937,N_14706);
xor UO_1527 (O_1527,N_14849,N_14864);
or UO_1528 (O_1528,N_14887,N_14746);
and UO_1529 (O_1529,N_14725,N_14864);
xor UO_1530 (O_1530,N_14814,N_14747);
or UO_1531 (O_1531,N_14787,N_14953);
or UO_1532 (O_1532,N_14928,N_14901);
nor UO_1533 (O_1533,N_14887,N_14908);
and UO_1534 (O_1534,N_14831,N_14718);
xor UO_1535 (O_1535,N_14825,N_14796);
nand UO_1536 (O_1536,N_14879,N_14834);
nand UO_1537 (O_1537,N_14983,N_14743);
and UO_1538 (O_1538,N_14918,N_14720);
and UO_1539 (O_1539,N_14908,N_14913);
nor UO_1540 (O_1540,N_14972,N_14856);
nor UO_1541 (O_1541,N_14805,N_14726);
or UO_1542 (O_1542,N_14717,N_14910);
nand UO_1543 (O_1543,N_14991,N_14778);
and UO_1544 (O_1544,N_14810,N_14876);
nand UO_1545 (O_1545,N_14750,N_14740);
nand UO_1546 (O_1546,N_14894,N_14882);
nor UO_1547 (O_1547,N_14833,N_14784);
and UO_1548 (O_1548,N_14792,N_14993);
nand UO_1549 (O_1549,N_14991,N_14950);
or UO_1550 (O_1550,N_14724,N_14946);
nor UO_1551 (O_1551,N_14937,N_14784);
nand UO_1552 (O_1552,N_14758,N_14971);
or UO_1553 (O_1553,N_14914,N_14950);
xnor UO_1554 (O_1554,N_14742,N_14826);
or UO_1555 (O_1555,N_14862,N_14817);
xor UO_1556 (O_1556,N_14951,N_14880);
or UO_1557 (O_1557,N_14799,N_14755);
or UO_1558 (O_1558,N_14784,N_14778);
or UO_1559 (O_1559,N_14842,N_14818);
and UO_1560 (O_1560,N_14832,N_14993);
nor UO_1561 (O_1561,N_14945,N_14866);
nor UO_1562 (O_1562,N_14816,N_14923);
xnor UO_1563 (O_1563,N_14738,N_14811);
xor UO_1564 (O_1564,N_14897,N_14915);
and UO_1565 (O_1565,N_14891,N_14790);
and UO_1566 (O_1566,N_14920,N_14961);
nand UO_1567 (O_1567,N_14935,N_14773);
nor UO_1568 (O_1568,N_14823,N_14918);
or UO_1569 (O_1569,N_14847,N_14917);
nand UO_1570 (O_1570,N_14725,N_14959);
nor UO_1571 (O_1571,N_14890,N_14777);
nor UO_1572 (O_1572,N_14997,N_14857);
or UO_1573 (O_1573,N_14709,N_14852);
nor UO_1574 (O_1574,N_14767,N_14745);
nor UO_1575 (O_1575,N_14801,N_14817);
xor UO_1576 (O_1576,N_14823,N_14761);
or UO_1577 (O_1577,N_14752,N_14975);
and UO_1578 (O_1578,N_14862,N_14822);
or UO_1579 (O_1579,N_14809,N_14811);
nor UO_1580 (O_1580,N_14973,N_14945);
nand UO_1581 (O_1581,N_14900,N_14761);
or UO_1582 (O_1582,N_14886,N_14826);
nand UO_1583 (O_1583,N_14912,N_14784);
xor UO_1584 (O_1584,N_14748,N_14952);
nor UO_1585 (O_1585,N_14804,N_14753);
and UO_1586 (O_1586,N_14903,N_14865);
nand UO_1587 (O_1587,N_14920,N_14862);
and UO_1588 (O_1588,N_14864,N_14917);
nor UO_1589 (O_1589,N_14930,N_14877);
xor UO_1590 (O_1590,N_14760,N_14855);
nor UO_1591 (O_1591,N_14989,N_14784);
nand UO_1592 (O_1592,N_14934,N_14735);
and UO_1593 (O_1593,N_14957,N_14901);
xnor UO_1594 (O_1594,N_14717,N_14831);
nor UO_1595 (O_1595,N_14834,N_14962);
or UO_1596 (O_1596,N_14943,N_14941);
nand UO_1597 (O_1597,N_14838,N_14964);
or UO_1598 (O_1598,N_14839,N_14729);
nand UO_1599 (O_1599,N_14864,N_14993);
or UO_1600 (O_1600,N_14875,N_14803);
nand UO_1601 (O_1601,N_14914,N_14938);
nand UO_1602 (O_1602,N_14970,N_14876);
nor UO_1603 (O_1603,N_14839,N_14928);
nand UO_1604 (O_1604,N_14853,N_14782);
and UO_1605 (O_1605,N_14964,N_14876);
or UO_1606 (O_1606,N_14815,N_14812);
or UO_1607 (O_1607,N_14775,N_14748);
or UO_1608 (O_1608,N_14721,N_14850);
nor UO_1609 (O_1609,N_14825,N_14761);
nor UO_1610 (O_1610,N_14785,N_14813);
nand UO_1611 (O_1611,N_14879,N_14822);
nor UO_1612 (O_1612,N_14956,N_14960);
or UO_1613 (O_1613,N_14821,N_14916);
and UO_1614 (O_1614,N_14983,N_14953);
nor UO_1615 (O_1615,N_14966,N_14962);
and UO_1616 (O_1616,N_14874,N_14885);
and UO_1617 (O_1617,N_14840,N_14944);
or UO_1618 (O_1618,N_14745,N_14707);
nand UO_1619 (O_1619,N_14956,N_14708);
xnor UO_1620 (O_1620,N_14743,N_14991);
xnor UO_1621 (O_1621,N_14819,N_14773);
or UO_1622 (O_1622,N_14743,N_14966);
nor UO_1623 (O_1623,N_14765,N_14752);
nor UO_1624 (O_1624,N_14969,N_14951);
nor UO_1625 (O_1625,N_14980,N_14915);
or UO_1626 (O_1626,N_14774,N_14916);
xor UO_1627 (O_1627,N_14899,N_14820);
nor UO_1628 (O_1628,N_14944,N_14763);
xor UO_1629 (O_1629,N_14820,N_14985);
and UO_1630 (O_1630,N_14827,N_14920);
xor UO_1631 (O_1631,N_14982,N_14924);
xnor UO_1632 (O_1632,N_14921,N_14934);
nor UO_1633 (O_1633,N_14996,N_14781);
or UO_1634 (O_1634,N_14838,N_14933);
or UO_1635 (O_1635,N_14925,N_14990);
nor UO_1636 (O_1636,N_14787,N_14820);
nand UO_1637 (O_1637,N_14730,N_14999);
xor UO_1638 (O_1638,N_14763,N_14880);
xnor UO_1639 (O_1639,N_14846,N_14760);
nand UO_1640 (O_1640,N_14819,N_14992);
or UO_1641 (O_1641,N_14891,N_14798);
and UO_1642 (O_1642,N_14750,N_14792);
nand UO_1643 (O_1643,N_14901,N_14742);
nor UO_1644 (O_1644,N_14725,N_14912);
xor UO_1645 (O_1645,N_14865,N_14801);
and UO_1646 (O_1646,N_14861,N_14719);
xor UO_1647 (O_1647,N_14839,N_14740);
nand UO_1648 (O_1648,N_14875,N_14885);
and UO_1649 (O_1649,N_14999,N_14739);
xnor UO_1650 (O_1650,N_14872,N_14803);
or UO_1651 (O_1651,N_14815,N_14970);
or UO_1652 (O_1652,N_14887,N_14949);
xor UO_1653 (O_1653,N_14831,N_14760);
or UO_1654 (O_1654,N_14988,N_14934);
xor UO_1655 (O_1655,N_14747,N_14764);
or UO_1656 (O_1656,N_14988,N_14974);
nand UO_1657 (O_1657,N_14820,N_14837);
nor UO_1658 (O_1658,N_14881,N_14815);
and UO_1659 (O_1659,N_14752,N_14887);
or UO_1660 (O_1660,N_14864,N_14973);
nor UO_1661 (O_1661,N_14701,N_14889);
nor UO_1662 (O_1662,N_14970,N_14804);
nand UO_1663 (O_1663,N_14909,N_14918);
and UO_1664 (O_1664,N_14792,N_14979);
and UO_1665 (O_1665,N_14789,N_14720);
or UO_1666 (O_1666,N_14976,N_14980);
nor UO_1667 (O_1667,N_14876,N_14830);
or UO_1668 (O_1668,N_14767,N_14830);
nor UO_1669 (O_1669,N_14975,N_14774);
xnor UO_1670 (O_1670,N_14774,N_14785);
or UO_1671 (O_1671,N_14968,N_14959);
nor UO_1672 (O_1672,N_14705,N_14941);
nor UO_1673 (O_1673,N_14769,N_14723);
and UO_1674 (O_1674,N_14802,N_14887);
or UO_1675 (O_1675,N_14730,N_14795);
nand UO_1676 (O_1676,N_14980,N_14986);
nor UO_1677 (O_1677,N_14989,N_14767);
and UO_1678 (O_1678,N_14725,N_14773);
xnor UO_1679 (O_1679,N_14821,N_14753);
nor UO_1680 (O_1680,N_14790,N_14868);
xor UO_1681 (O_1681,N_14982,N_14828);
nor UO_1682 (O_1682,N_14758,N_14836);
xor UO_1683 (O_1683,N_14859,N_14865);
or UO_1684 (O_1684,N_14863,N_14725);
or UO_1685 (O_1685,N_14889,N_14977);
or UO_1686 (O_1686,N_14931,N_14772);
nand UO_1687 (O_1687,N_14930,N_14814);
or UO_1688 (O_1688,N_14871,N_14739);
and UO_1689 (O_1689,N_14735,N_14972);
nor UO_1690 (O_1690,N_14890,N_14942);
nor UO_1691 (O_1691,N_14782,N_14785);
or UO_1692 (O_1692,N_14886,N_14931);
nand UO_1693 (O_1693,N_14884,N_14881);
and UO_1694 (O_1694,N_14951,N_14973);
nand UO_1695 (O_1695,N_14876,N_14938);
or UO_1696 (O_1696,N_14769,N_14881);
nor UO_1697 (O_1697,N_14727,N_14995);
nor UO_1698 (O_1698,N_14764,N_14762);
and UO_1699 (O_1699,N_14728,N_14767);
or UO_1700 (O_1700,N_14819,N_14945);
nor UO_1701 (O_1701,N_14810,N_14757);
nor UO_1702 (O_1702,N_14936,N_14700);
nor UO_1703 (O_1703,N_14849,N_14823);
and UO_1704 (O_1704,N_14875,N_14817);
nor UO_1705 (O_1705,N_14918,N_14748);
or UO_1706 (O_1706,N_14983,N_14905);
nand UO_1707 (O_1707,N_14976,N_14819);
and UO_1708 (O_1708,N_14731,N_14720);
xnor UO_1709 (O_1709,N_14763,N_14832);
nand UO_1710 (O_1710,N_14780,N_14844);
xor UO_1711 (O_1711,N_14929,N_14996);
or UO_1712 (O_1712,N_14859,N_14909);
nor UO_1713 (O_1713,N_14915,N_14752);
nand UO_1714 (O_1714,N_14749,N_14721);
nand UO_1715 (O_1715,N_14810,N_14928);
nand UO_1716 (O_1716,N_14722,N_14840);
and UO_1717 (O_1717,N_14806,N_14780);
nand UO_1718 (O_1718,N_14754,N_14885);
nor UO_1719 (O_1719,N_14991,N_14929);
or UO_1720 (O_1720,N_14796,N_14827);
and UO_1721 (O_1721,N_14878,N_14785);
xor UO_1722 (O_1722,N_14954,N_14731);
nor UO_1723 (O_1723,N_14874,N_14700);
xnor UO_1724 (O_1724,N_14838,N_14991);
nor UO_1725 (O_1725,N_14715,N_14720);
nor UO_1726 (O_1726,N_14757,N_14848);
nand UO_1727 (O_1727,N_14727,N_14916);
nand UO_1728 (O_1728,N_14731,N_14820);
nand UO_1729 (O_1729,N_14973,N_14986);
nor UO_1730 (O_1730,N_14923,N_14914);
xnor UO_1731 (O_1731,N_14818,N_14719);
nand UO_1732 (O_1732,N_14759,N_14890);
nor UO_1733 (O_1733,N_14801,N_14997);
or UO_1734 (O_1734,N_14879,N_14932);
or UO_1735 (O_1735,N_14709,N_14744);
xnor UO_1736 (O_1736,N_14743,N_14758);
xor UO_1737 (O_1737,N_14703,N_14921);
nand UO_1738 (O_1738,N_14918,N_14781);
or UO_1739 (O_1739,N_14781,N_14937);
or UO_1740 (O_1740,N_14943,N_14933);
nand UO_1741 (O_1741,N_14926,N_14727);
xnor UO_1742 (O_1742,N_14797,N_14710);
or UO_1743 (O_1743,N_14822,N_14998);
xnor UO_1744 (O_1744,N_14867,N_14969);
nand UO_1745 (O_1745,N_14932,N_14875);
nor UO_1746 (O_1746,N_14954,N_14773);
and UO_1747 (O_1747,N_14933,N_14994);
or UO_1748 (O_1748,N_14779,N_14989);
nor UO_1749 (O_1749,N_14987,N_14980);
or UO_1750 (O_1750,N_14742,N_14753);
xnor UO_1751 (O_1751,N_14874,N_14926);
nand UO_1752 (O_1752,N_14805,N_14732);
xnor UO_1753 (O_1753,N_14739,N_14924);
and UO_1754 (O_1754,N_14779,N_14734);
nor UO_1755 (O_1755,N_14782,N_14740);
nand UO_1756 (O_1756,N_14992,N_14952);
xnor UO_1757 (O_1757,N_14868,N_14974);
or UO_1758 (O_1758,N_14928,N_14885);
or UO_1759 (O_1759,N_14712,N_14994);
xnor UO_1760 (O_1760,N_14847,N_14807);
and UO_1761 (O_1761,N_14700,N_14763);
xnor UO_1762 (O_1762,N_14728,N_14892);
xnor UO_1763 (O_1763,N_14777,N_14816);
nor UO_1764 (O_1764,N_14992,N_14939);
or UO_1765 (O_1765,N_14901,N_14701);
and UO_1766 (O_1766,N_14983,N_14789);
xnor UO_1767 (O_1767,N_14773,N_14998);
nand UO_1768 (O_1768,N_14970,N_14734);
xor UO_1769 (O_1769,N_14998,N_14973);
nor UO_1770 (O_1770,N_14876,N_14866);
or UO_1771 (O_1771,N_14852,N_14968);
nand UO_1772 (O_1772,N_14945,N_14727);
nand UO_1773 (O_1773,N_14708,N_14828);
xnor UO_1774 (O_1774,N_14728,N_14978);
nor UO_1775 (O_1775,N_14895,N_14745);
and UO_1776 (O_1776,N_14796,N_14793);
or UO_1777 (O_1777,N_14814,N_14746);
nand UO_1778 (O_1778,N_14951,N_14717);
nor UO_1779 (O_1779,N_14866,N_14924);
and UO_1780 (O_1780,N_14737,N_14966);
nor UO_1781 (O_1781,N_14807,N_14991);
xor UO_1782 (O_1782,N_14753,N_14829);
or UO_1783 (O_1783,N_14866,N_14837);
or UO_1784 (O_1784,N_14707,N_14966);
nand UO_1785 (O_1785,N_14821,N_14833);
and UO_1786 (O_1786,N_14968,N_14988);
or UO_1787 (O_1787,N_14740,N_14763);
or UO_1788 (O_1788,N_14708,N_14912);
nor UO_1789 (O_1789,N_14883,N_14728);
or UO_1790 (O_1790,N_14786,N_14754);
and UO_1791 (O_1791,N_14925,N_14734);
nand UO_1792 (O_1792,N_14832,N_14872);
xnor UO_1793 (O_1793,N_14938,N_14777);
nor UO_1794 (O_1794,N_14750,N_14747);
nand UO_1795 (O_1795,N_14787,N_14941);
nand UO_1796 (O_1796,N_14966,N_14880);
and UO_1797 (O_1797,N_14797,N_14761);
and UO_1798 (O_1798,N_14936,N_14959);
nor UO_1799 (O_1799,N_14866,N_14907);
and UO_1800 (O_1800,N_14824,N_14870);
nor UO_1801 (O_1801,N_14937,N_14947);
or UO_1802 (O_1802,N_14964,N_14852);
and UO_1803 (O_1803,N_14845,N_14879);
nand UO_1804 (O_1804,N_14958,N_14780);
nand UO_1805 (O_1805,N_14810,N_14888);
or UO_1806 (O_1806,N_14735,N_14825);
nor UO_1807 (O_1807,N_14973,N_14928);
and UO_1808 (O_1808,N_14848,N_14953);
xor UO_1809 (O_1809,N_14779,N_14780);
and UO_1810 (O_1810,N_14851,N_14904);
nand UO_1811 (O_1811,N_14802,N_14979);
or UO_1812 (O_1812,N_14985,N_14892);
xor UO_1813 (O_1813,N_14751,N_14819);
nor UO_1814 (O_1814,N_14850,N_14885);
nor UO_1815 (O_1815,N_14937,N_14736);
nand UO_1816 (O_1816,N_14758,N_14714);
nand UO_1817 (O_1817,N_14756,N_14861);
or UO_1818 (O_1818,N_14810,N_14944);
or UO_1819 (O_1819,N_14803,N_14868);
and UO_1820 (O_1820,N_14805,N_14935);
and UO_1821 (O_1821,N_14877,N_14857);
or UO_1822 (O_1822,N_14924,N_14756);
or UO_1823 (O_1823,N_14824,N_14895);
nor UO_1824 (O_1824,N_14899,N_14857);
and UO_1825 (O_1825,N_14852,N_14775);
nand UO_1826 (O_1826,N_14868,N_14893);
nor UO_1827 (O_1827,N_14788,N_14956);
and UO_1828 (O_1828,N_14777,N_14769);
or UO_1829 (O_1829,N_14798,N_14921);
xor UO_1830 (O_1830,N_14791,N_14826);
nand UO_1831 (O_1831,N_14967,N_14866);
and UO_1832 (O_1832,N_14729,N_14928);
and UO_1833 (O_1833,N_14806,N_14921);
or UO_1834 (O_1834,N_14703,N_14778);
nand UO_1835 (O_1835,N_14935,N_14714);
and UO_1836 (O_1836,N_14752,N_14922);
nor UO_1837 (O_1837,N_14873,N_14926);
nand UO_1838 (O_1838,N_14846,N_14895);
nand UO_1839 (O_1839,N_14784,N_14770);
and UO_1840 (O_1840,N_14940,N_14913);
and UO_1841 (O_1841,N_14931,N_14821);
nand UO_1842 (O_1842,N_14808,N_14861);
or UO_1843 (O_1843,N_14915,N_14849);
or UO_1844 (O_1844,N_14748,N_14797);
and UO_1845 (O_1845,N_14859,N_14893);
and UO_1846 (O_1846,N_14938,N_14833);
xor UO_1847 (O_1847,N_14994,N_14756);
and UO_1848 (O_1848,N_14712,N_14912);
xnor UO_1849 (O_1849,N_14891,N_14731);
nand UO_1850 (O_1850,N_14986,N_14812);
xor UO_1851 (O_1851,N_14772,N_14945);
nor UO_1852 (O_1852,N_14844,N_14883);
nand UO_1853 (O_1853,N_14861,N_14924);
xor UO_1854 (O_1854,N_14993,N_14895);
or UO_1855 (O_1855,N_14960,N_14822);
nor UO_1856 (O_1856,N_14959,N_14990);
xor UO_1857 (O_1857,N_14987,N_14970);
nand UO_1858 (O_1858,N_14983,N_14864);
and UO_1859 (O_1859,N_14763,N_14857);
nor UO_1860 (O_1860,N_14703,N_14767);
xnor UO_1861 (O_1861,N_14703,N_14977);
xnor UO_1862 (O_1862,N_14875,N_14918);
nand UO_1863 (O_1863,N_14923,N_14841);
nor UO_1864 (O_1864,N_14931,N_14844);
nor UO_1865 (O_1865,N_14932,N_14721);
and UO_1866 (O_1866,N_14875,N_14721);
or UO_1867 (O_1867,N_14701,N_14744);
xor UO_1868 (O_1868,N_14866,N_14750);
xor UO_1869 (O_1869,N_14855,N_14902);
or UO_1870 (O_1870,N_14871,N_14773);
or UO_1871 (O_1871,N_14719,N_14740);
xnor UO_1872 (O_1872,N_14989,N_14742);
xor UO_1873 (O_1873,N_14954,N_14919);
or UO_1874 (O_1874,N_14976,N_14757);
xnor UO_1875 (O_1875,N_14856,N_14750);
xnor UO_1876 (O_1876,N_14919,N_14714);
and UO_1877 (O_1877,N_14985,N_14934);
nand UO_1878 (O_1878,N_14719,N_14992);
nand UO_1879 (O_1879,N_14773,N_14890);
xnor UO_1880 (O_1880,N_14799,N_14786);
nand UO_1881 (O_1881,N_14886,N_14932);
nand UO_1882 (O_1882,N_14879,N_14783);
or UO_1883 (O_1883,N_14702,N_14878);
or UO_1884 (O_1884,N_14900,N_14832);
or UO_1885 (O_1885,N_14900,N_14847);
xor UO_1886 (O_1886,N_14746,N_14933);
and UO_1887 (O_1887,N_14780,N_14730);
or UO_1888 (O_1888,N_14954,N_14890);
or UO_1889 (O_1889,N_14980,N_14926);
nor UO_1890 (O_1890,N_14757,N_14751);
and UO_1891 (O_1891,N_14724,N_14804);
xnor UO_1892 (O_1892,N_14786,N_14854);
nand UO_1893 (O_1893,N_14833,N_14839);
or UO_1894 (O_1894,N_14909,N_14981);
or UO_1895 (O_1895,N_14907,N_14982);
xnor UO_1896 (O_1896,N_14770,N_14925);
xnor UO_1897 (O_1897,N_14954,N_14736);
xor UO_1898 (O_1898,N_14711,N_14936);
and UO_1899 (O_1899,N_14731,N_14858);
nor UO_1900 (O_1900,N_14705,N_14710);
and UO_1901 (O_1901,N_14728,N_14784);
or UO_1902 (O_1902,N_14982,N_14819);
xnor UO_1903 (O_1903,N_14921,N_14843);
and UO_1904 (O_1904,N_14755,N_14853);
nor UO_1905 (O_1905,N_14799,N_14837);
xnor UO_1906 (O_1906,N_14812,N_14943);
xor UO_1907 (O_1907,N_14744,N_14787);
and UO_1908 (O_1908,N_14927,N_14822);
and UO_1909 (O_1909,N_14893,N_14981);
xnor UO_1910 (O_1910,N_14986,N_14911);
nand UO_1911 (O_1911,N_14817,N_14716);
or UO_1912 (O_1912,N_14774,N_14976);
or UO_1913 (O_1913,N_14958,N_14955);
and UO_1914 (O_1914,N_14905,N_14963);
nand UO_1915 (O_1915,N_14854,N_14956);
xor UO_1916 (O_1916,N_14931,N_14753);
and UO_1917 (O_1917,N_14822,N_14926);
xor UO_1918 (O_1918,N_14709,N_14727);
nand UO_1919 (O_1919,N_14805,N_14791);
or UO_1920 (O_1920,N_14919,N_14756);
or UO_1921 (O_1921,N_14960,N_14849);
or UO_1922 (O_1922,N_14964,N_14841);
xnor UO_1923 (O_1923,N_14760,N_14900);
xnor UO_1924 (O_1924,N_14754,N_14855);
xnor UO_1925 (O_1925,N_14779,N_14876);
or UO_1926 (O_1926,N_14961,N_14721);
xor UO_1927 (O_1927,N_14944,N_14890);
and UO_1928 (O_1928,N_14711,N_14874);
nor UO_1929 (O_1929,N_14950,N_14736);
and UO_1930 (O_1930,N_14880,N_14752);
xor UO_1931 (O_1931,N_14961,N_14868);
and UO_1932 (O_1932,N_14792,N_14841);
nor UO_1933 (O_1933,N_14961,N_14900);
and UO_1934 (O_1934,N_14722,N_14868);
and UO_1935 (O_1935,N_14916,N_14875);
and UO_1936 (O_1936,N_14818,N_14739);
nor UO_1937 (O_1937,N_14716,N_14930);
nor UO_1938 (O_1938,N_14892,N_14973);
nand UO_1939 (O_1939,N_14973,N_14960);
xor UO_1940 (O_1940,N_14761,N_14983);
nor UO_1941 (O_1941,N_14975,N_14720);
or UO_1942 (O_1942,N_14932,N_14854);
or UO_1943 (O_1943,N_14888,N_14845);
nor UO_1944 (O_1944,N_14728,N_14711);
nand UO_1945 (O_1945,N_14825,N_14829);
nand UO_1946 (O_1946,N_14918,N_14754);
or UO_1947 (O_1947,N_14873,N_14904);
and UO_1948 (O_1948,N_14821,N_14869);
or UO_1949 (O_1949,N_14776,N_14991);
nor UO_1950 (O_1950,N_14759,N_14787);
nor UO_1951 (O_1951,N_14805,N_14987);
nand UO_1952 (O_1952,N_14757,N_14730);
nand UO_1953 (O_1953,N_14865,N_14844);
and UO_1954 (O_1954,N_14714,N_14980);
nor UO_1955 (O_1955,N_14933,N_14946);
and UO_1956 (O_1956,N_14758,N_14850);
xnor UO_1957 (O_1957,N_14817,N_14854);
nor UO_1958 (O_1958,N_14796,N_14868);
or UO_1959 (O_1959,N_14998,N_14832);
and UO_1960 (O_1960,N_14743,N_14745);
nand UO_1961 (O_1961,N_14763,N_14747);
or UO_1962 (O_1962,N_14867,N_14927);
xnor UO_1963 (O_1963,N_14985,N_14883);
nand UO_1964 (O_1964,N_14850,N_14709);
nor UO_1965 (O_1965,N_14822,N_14982);
and UO_1966 (O_1966,N_14950,N_14724);
nand UO_1967 (O_1967,N_14926,N_14837);
xor UO_1968 (O_1968,N_14876,N_14745);
and UO_1969 (O_1969,N_14783,N_14838);
xor UO_1970 (O_1970,N_14886,N_14718);
xor UO_1971 (O_1971,N_14767,N_14875);
and UO_1972 (O_1972,N_14779,N_14760);
nand UO_1973 (O_1973,N_14732,N_14818);
nor UO_1974 (O_1974,N_14834,N_14958);
xor UO_1975 (O_1975,N_14746,N_14700);
xnor UO_1976 (O_1976,N_14709,N_14999);
xor UO_1977 (O_1977,N_14954,N_14842);
nand UO_1978 (O_1978,N_14963,N_14811);
or UO_1979 (O_1979,N_14721,N_14825);
nor UO_1980 (O_1980,N_14824,N_14928);
or UO_1981 (O_1981,N_14942,N_14812);
nand UO_1982 (O_1982,N_14707,N_14872);
nor UO_1983 (O_1983,N_14975,N_14938);
or UO_1984 (O_1984,N_14994,N_14923);
or UO_1985 (O_1985,N_14731,N_14970);
nand UO_1986 (O_1986,N_14783,N_14743);
xnor UO_1987 (O_1987,N_14767,N_14972);
nor UO_1988 (O_1988,N_14783,N_14900);
and UO_1989 (O_1989,N_14786,N_14914);
nor UO_1990 (O_1990,N_14989,N_14979);
nor UO_1991 (O_1991,N_14768,N_14894);
and UO_1992 (O_1992,N_14778,N_14857);
or UO_1993 (O_1993,N_14796,N_14894);
and UO_1994 (O_1994,N_14865,N_14761);
nand UO_1995 (O_1995,N_14945,N_14861);
nand UO_1996 (O_1996,N_14883,N_14890);
nor UO_1997 (O_1997,N_14876,N_14804);
or UO_1998 (O_1998,N_14850,N_14972);
nor UO_1999 (O_1999,N_14919,N_14770);
endmodule