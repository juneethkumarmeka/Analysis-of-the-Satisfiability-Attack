module basic_500_3000_500_40_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_135,In_16);
nor U1 (N_1,In_394,In_379);
and U2 (N_2,In_90,In_62);
or U3 (N_3,In_300,In_23);
or U4 (N_4,In_491,In_433);
or U5 (N_5,In_281,In_488);
nand U6 (N_6,In_121,In_44);
nand U7 (N_7,In_359,In_184);
nand U8 (N_8,In_126,In_391);
nor U9 (N_9,In_89,In_479);
and U10 (N_10,In_361,In_198);
and U11 (N_11,In_154,In_145);
or U12 (N_12,In_342,In_67);
nand U13 (N_13,In_494,In_306);
nor U14 (N_14,In_478,In_167);
nand U15 (N_15,In_321,In_490);
or U16 (N_16,In_98,In_445);
nand U17 (N_17,In_327,In_70);
nand U18 (N_18,In_156,In_497);
nor U19 (N_19,In_415,In_383);
nor U20 (N_20,In_111,In_343);
and U21 (N_21,In_205,In_81);
nand U22 (N_22,In_475,In_13);
or U23 (N_23,In_458,In_416);
and U24 (N_24,In_131,In_243);
nand U25 (N_25,In_171,In_88);
and U26 (N_26,In_214,In_168);
nand U27 (N_27,In_328,In_489);
nand U28 (N_28,In_254,In_95);
and U29 (N_29,In_474,In_387);
nor U30 (N_30,In_389,In_222);
and U31 (N_31,In_79,In_194);
or U32 (N_32,In_272,In_332);
or U33 (N_33,In_467,In_166);
nand U34 (N_34,In_106,In_443);
nor U35 (N_35,In_178,In_437);
or U36 (N_36,In_333,In_316);
and U37 (N_37,In_211,In_498);
nor U38 (N_38,In_65,In_68);
nand U39 (N_39,In_124,In_364);
nand U40 (N_40,In_63,In_227);
and U41 (N_41,In_173,In_302);
xor U42 (N_42,In_353,In_418);
nor U43 (N_43,In_232,In_288);
nand U44 (N_44,In_197,In_9);
or U45 (N_45,In_151,In_230);
and U46 (N_46,In_223,In_268);
nand U47 (N_47,In_24,In_294);
or U48 (N_48,In_405,In_440);
or U49 (N_49,In_355,In_477);
nand U50 (N_50,In_141,In_301);
xor U51 (N_51,In_344,In_19);
or U52 (N_52,In_201,In_204);
nand U53 (N_53,In_77,In_114);
nand U54 (N_54,In_191,In_400);
and U55 (N_55,In_380,In_435);
nand U56 (N_56,In_384,In_107);
nor U57 (N_57,In_469,In_410);
and U58 (N_58,In_259,In_284);
nor U59 (N_59,In_202,In_92);
or U60 (N_60,In_461,In_320);
nand U61 (N_61,In_110,In_282);
nor U62 (N_62,In_319,In_221);
nor U63 (N_63,In_404,In_464);
nand U64 (N_64,In_185,In_118);
nand U65 (N_65,In_8,In_12);
and U66 (N_66,In_426,In_434);
nor U67 (N_67,In_439,In_448);
nor U68 (N_68,In_109,In_401);
nand U69 (N_69,In_462,In_451);
nand U70 (N_70,In_103,In_357);
and U71 (N_71,In_483,In_245);
and U72 (N_72,In_388,In_422);
or U73 (N_73,In_240,In_396);
xnor U74 (N_74,In_269,In_378);
nand U75 (N_75,In_363,In_480);
and U76 (N_76,N_12,In_455);
nand U77 (N_77,In_188,In_367);
and U78 (N_78,In_438,In_208);
or U79 (N_79,In_80,In_172);
nor U80 (N_80,In_279,In_399);
and U81 (N_81,In_417,N_52);
nand U82 (N_82,In_5,In_148);
nand U83 (N_83,In_72,In_161);
and U84 (N_84,In_52,N_34);
and U85 (N_85,In_429,In_116);
or U86 (N_86,In_213,In_74);
or U87 (N_87,In_348,N_43);
and U88 (N_88,In_481,N_53);
or U89 (N_89,In_49,N_46);
or U90 (N_90,N_50,In_210);
or U91 (N_91,In_220,In_340);
and U92 (N_92,In_122,In_177);
xor U93 (N_93,N_13,In_39);
and U94 (N_94,N_3,N_36);
and U95 (N_95,In_246,In_133);
or U96 (N_96,In_225,In_331);
nor U97 (N_97,In_250,In_60);
and U98 (N_98,In_249,In_432);
and U99 (N_99,In_130,In_436);
nor U100 (N_100,N_21,In_486);
or U101 (N_101,In_216,N_29);
and U102 (N_102,In_162,In_160);
and U103 (N_103,In_492,In_186);
nor U104 (N_104,In_397,In_356);
nand U105 (N_105,In_179,In_447);
nand U106 (N_106,In_1,N_14);
nor U107 (N_107,In_326,In_192);
nor U108 (N_108,In_175,In_449);
nand U109 (N_109,N_17,In_460);
and U110 (N_110,In_260,In_354);
nand U111 (N_111,In_2,In_76);
and U112 (N_112,In_466,N_74);
or U113 (N_113,In_311,In_149);
and U114 (N_114,In_127,In_142);
or U115 (N_115,N_56,In_83);
and U116 (N_116,In_85,In_253);
or U117 (N_117,N_8,N_20);
nand U118 (N_118,In_117,In_330);
nor U119 (N_119,In_105,In_123);
xnor U120 (N_120,N_42,N_59);
xor U121 (N_121,In_263,In_362);
xor U122 (N_122,In_199,In_265);
nor U123 (N_123,In_159,N_45);
or U124 (N_124,In_27,N_26);
nor U125 (N_125,In_91,In_43);
nand U126 (N_126,In_29,N_24);
nand U127 (N_127,In_459,In_390);
and U128 (N_128,In_21,In_4);
or U129 (N_129,In_351,In_406);
or U130 (N_130,In_203,In_17);
nand U131 (N_131,In_86,In_412);
and U132 (N_132,In_84,In_365);
or U133 (N_133,In_305,In_385);
xnor U134 (N_134,In_457,In_42);
nor U135 (N_135,In_495,In_102);
xor U136 (N_136,N_63,In_446);
nand U137 (N_137,In_233,N_61);
or U138 (N_138,In_180,In_442);
and U139 (N_139,In_182,In_163);
or U140 (N_140,In_82,In_235);
nor U141 (N_141,In_36,In_381);
and U142 (N_142,In_31,In_248);
nor U143 (N_143,In_61,N_10);
or U144 (N_144,In_78,In_196);
nor U145 (N_145,In_3,N_30);
nor U146 (N_146,In_408,In_270);
or U147 (N_147,In_153,In_34);
nor U148 (N_148,In_138,In_373);
and U149 (N_149,In_368,In_349);
nor U150 (N_150,In_323,In_174);
or U151 (N_151,N_7,N_25);
nor U152 (N_152,In_393,N_143);
and U153 (N_153,N_117,N_81);
nand U154 (N_154,In_339,N_23);
nor U155 (N_155,In_144,In_137);
nor U156 (N_156,In_108,N_70);
nor U157 (N_157,N_106,In_38);
and U158 (N_158,In_285,In_244);
nand U159 (N_159,In_283,N_78);
and U160 (N_160,In_150,In_193);
nand U161 (N_161,N_147,In_33);
or U162 (N_162,In_298,In_266);
nor U163 (N_163,In_18,N_65);
and U164 (N_164,N_140,N_47);
nand U165 (N_165,In_371,N_124);
nor U166 (N_166,In_10,N_98);
or U167 (N_167,In_414,In_452);
xor U168 (N_168,In_238,In_382);
nand U169 (N_169,In_45,In_25);
xnor U170 (N_170,N_108,In_471);
and U171 (N_171,In_256,N_100);
nor U172 (N_172,In_58,In_485);
or U173 (N_173,In_112,N_136);
and U174 (N_174,N_57,In_407);
nor U175 (N_175,In_409,In_375);
or U176 (N_176,In_309,N_31);
and U177 (N_177,In_465,In_87);
nand U178 (N_178,In_341,In_258);
nand U179 (N_179,N_66,In_212);
nand U180 (N_180,In_242,N_62);
nor U181 (N_181,In_48,In_73);
or U182 (N_182,In_207,In_496);
nand U183 (N_183,In_146,N_54);
nor U184 (N_184,In_54,In_20);
nand U185 (N_185,N_133,In_170);
nand U186 (N_186,In_75,In_15);
or U187 (N_187,N_67,In_484);
and U188 (N_188,In_325,N_126);
and U189 (N_189,In_470,In_181);
xor U190 (N_190,In_97,In_428);
nor U191 (N_191,In_189,N_103);
and U192 (N_192,In_66,In_420);
nand U193 (N_193,N_68,N_107);
or U194 (N_194,In_6,In_421);
nand U195 (N_195,In_28,In_337);
nand U196 (N_196,N_16,In_308);
nand U197 (N_197,In_165,N_148);
or U198 (N_198,N_123,N_122);
nand U199 (N_199,In_158,In_291);
or U200 (N_200,N_130,In_94);
nor U201 (N_201,In_136,N_39);
nand U202 (N_202,N_33,N_115);
nor U203 (N_203,In_99,In_450);
or U204 (N_204,In_219,N_60);
and U205 (N_205,N_69,In_104);
or U206 (N_206,N_146,In_274);
nand U207 (N_207,In_290,N_2);
nor U208 (N_208,In_187,In_277);
nand U209 (N_209,In_157,In_129);
nand U210 (N_210,N_138,N_22);
nand U211 (N_211,In_376,In_315);
nand U212 (N_212,In_264,In_128);
or U213 (N_213,In_476,N_125);
nand U214 (N_214,In_46,In_55);
and U215 (N_215,N_19,In_338);
nand U216 (N_216,In_231,In_329);
or U217 (N_217,N_92,In_229);
or U218 (N_218,In_424,N_51);
nand U219 (N_219,N_111,In_32);
and U220 (N_220,In_50,N_4);
nor U221 (N_221,In_345,N_149);
nand U222 (N_222,In_403,N_37);
nand U223 (N_223,In_51,In_247);
or U224 (N_224,N_80,N_28);
nor U225 (N_225,N_120,In_431);
and U226 (N_226,N_184,In_304);
and U227 (N_227,In_295,N_176);
and U228 (N_228,N_212,In_468);
nand U229 (N_229,N_104,N_102);
nand U230 (N_230,In_101,N_110);
nor U231 (N_231,N_183,In_493);
nor U232 (N_232,N_89,N_202);
nand U233 (N_233,N_142,N_160);
nor U234 (N_234,In_206,In_143);
and U235 (N_235,In_395,N_11);
nand U236 (N_236,In_47,In_287);
nor U237 (N_237,In_56,In_134);
and U238 (N_238,In_350,N_82);
or U239 (N_239,In_261,N_152);
nand U240 (N_240,N_131,N_180);
xor U241 (N_241,N_174,N_18);
nor U242 (N_242,In_226,In_377);
nand U243 (N_243,In_236,N_206);
xnor U244 (N_244,N_189,N_216);
or U245 (N_245,N_141,N_159);
and U246 (N_246,In_241,In_35);
nor U247 (N_247,In_59,In_57);
and U248 (N_248,N_150,In_237);
nand U249 (N_249,N_95,N_83);
and U250 (N_250,In_200,N_161);
nand U251 (N_251,N_190,In_402);
and U252 (N_252,N_38,In_96);
or U253 (N_253,N_204,In_366);
nor U254 (N_254,N_6,N_0);
and U255 (N_255,N_129,N_58);
or U256 (N_256,In_411,N_166);
nand U257 (N_257,In_276,N_220);
or U258 (N_258,In_322,In_358);
or U259 (N_259,In_372,N_114);
nand U260 (N_260,In_228,In_100);
nor U261 (N_261,In_352,In_299);
xnor U262 (N_262,N_93,N_145);
nor U263 (N_263,N_177,N_151);
and U264 (N_264,N_209,In_115);
nand U265 (N_265,N_5,N_96);
or U266 (N_266,N_44,In_40);
nor U267 (N_267,N_88,N_101);
or U268 (N_268,N_179,In_69);
and U269 (N_269,In_347,In_482);
or U270 (N_270,In_139,N_35);
nand U271 (N_271,N_200,N_75);
nor U272 (N_272,In_293,N_9);
or U273 (N_273,In_37,N_99);
or U274 (N_274,In_312,In_423);
nand U275 (N_275,In_317,In_297);
xor U276 (N_276,In_252,N_76);
xor U277 (N_277,N_197,N_86);
and U278 (N_278,N_210,N_48);
nand U279 (N_279,In_307,N_94);
nor U280 (N_280,N_153,In_370);
nor U281 (N_281,N_85,N_182);
or U282 (N_282,N_155,N_156);
nor U283 (N_283,N_215,N_77);
nand U284 (N_284,N_222,N_217);
or U285 (N_285,N_121,In_441);
xnor U286 (N_286,N_84,In_463);
and U287 (N_287,In_0,In_456);
nand U288 (N_288,N_139,In_454);
nand U289 (N_289,N_175,In_419);
xnor U290 (N_290,In_53,N_119);
xnor U291 (N_291,N_211,In_335);
nand U292 (N_292,In_398,N_87);
nor U293 (N_293,In_169,N_97);
nand U294 (N_294,In_22,N_214);
and U295 (N_295,N_49,N_41);
nor U296 (N_296,In_289,N_105);
and U297 (N_297,N_132,N_40);
nand U298 (N_298,In_155,N_207);
nand U299 (N_299,N_173,N_168);
or U300 (N_300,In_215,N_272);
and U301 (N_301,N_273,N_282);
or U302 (N_302,In_224,N_292);
nor U303 (N_303,In_310,N_191);
or U304 (N_304,In_71,N_154);
xor U305 (N_305,N_266,In_125);
xnor U306 (N_306,N_275,In_164);
and U307 (N_307,N_293,In_487);
nor U308 (N_308,N_240,N_196);
or U309 (N_309,N_255,In_251);
nand U310 (N_310,In_120,N_285);
nor U311 (N_311,N_251,N_268);
nand U312 (N_312,N_278,N_223);
and U313 (N_313,N_192,In_93);
and U314 (N_314,N_172,N_257);
nor U315 (N_315,N_187,N_205);
xnor U316 (N_316,In_11,In_499);
nor U317 (N_317,In_113,N_232);
or U318 (N_318,N_269,In_292);
and U319 (N_319,In_41,In_64);
nand U320 (N_320,N_64,N_198);
or U321 (N_321,In_346,N_298);
nand U322 (N_322,N_165,N_260);
or U323 (N_323,N_291,N_241);
and U324 (N_324,N_118,N_283);
nor U325 (N_325,N_163,In_132);
xnor U326 (N_326,N_242,N_201);
nor U327 (N_327,In_430,N_297);
nand U328 (N_328,N_73,In_234);
xnor U329 (N_329,N_279,N_229);
nand U330 (N_330,N_277,In_255);
and U331 (N_331,In_183,In_303);
nor U332 (N_332,N_258,N_246);
xnor U333 (N_333,In_195,N_109);
nand U334 (N_334,N_195,N_224);
nand U335 (N_335,In_296,N_226);
or U336 (N_336,N_264,N_267);
nor U337 (N_337,In_14,N_274);
nor U338 (N_338,In_7,N_134);
and U339 (N_339,In_119,N_238);
xor U340 (N_340,N_27,N_91);
and U341 (N_341,N_55,N_213);
nand U342 (N_342,N_243,In_209);
or U343 (N_343,N_271,N_233);
nor U344 (N_344,N_171,N_254);
or U345 (N_345,N_208,In_473);
and U346 (N_346,N_181,N_249);
nand U347 (N_347,In_190,In_392);
nand U348 (N_348,N_221,In_217);
nand U349 (N_349,In_273,In_453);
nor U350 (N_350,N_71,N_250);
nand U351 (N_351,N_234,In_313);
or U352 (N_352,In_444,N_244);
and U353 (N_353,N_236,N_199);
nand U354 (N_354,N_186,N_79);
nor U355 (N_355,N_90,In_369);
or U356 (N_356,In_314,N_157);
nor U357 (N_357,In_280,In_336);
and U358 (N_358,In_386,N_15);
nor U359 (N_359,In_286,N_265);
xor U360 (N_360,In_262,N_287);
or U361 (N_361,In_30,N_281);
and U362 (N_362,N_135,In_278);
nor U363 (N_363,N_170,In_324);
nor U364 (N_364,In_472,N_270);
xnor U365 (N_365,In_267,N_230);
and U366 (N_366,N_167,N_158);
nand U367 (N_367,N_294,N_263);
or U368 (N_368,N_288,N_296);
nand U369 (N_369,N_137,N_164);
nor U370 (N_370,In_26,N_185);
nand U371 (N_371,N_280,N_1);
nand U372 (N_372,In_374,N_290);
or U373 (N_373,In_140,N_162);
nor U374 (N_374,N_261,N_32);
nor U375 (N_375,N_231,N_72);
nor U376 (N_376,N_353,N_188);
nand U377 (N_377,N_300,N_235);
nand U378 (N_378,N_365,N_326);
or U379 (N_379,N_304,N_262);
and U380 (N_380,N_350,N_370);
or U381 (N_381,N_256,N_314);
nand U382 (N_382,N_349,N_308);
and U383 (N_383,In_360,N_144);
nor U384 (N_384,N_363,N_253);
nand U385 (N_385,N_301,N_219);
nor U386 (N_386,In_334,N_307);
or U387 (N_387,N_323,N_343);
or U388 (N_388,In_318,N_374);
or U389 (N_389,N_329,N_237);
or U390 (N_390,N_335,N_295);
and U391 (N_391,N_276,N_284);
and U392 (N_392,N_360,N_316);
xnor U393 (N_393,N_194,N_356);
and U394 (N_394,N_310,N_245);
xor U395 (N_395,N_342,N_324);
nor U396 (N_396,N_302,N_228);
nand U397 (N_397,N_127,N_112);
and U398 (N_398,N_252,N_259);
nor U399 (N_399,In_147,In_275);
or U400 (N_400,N_346,N_289);
or U401 (N_401,N_367,N_321);
and U402 (N_402,N_334,N_325);
and U403 (N_403,N_337,N_322);
and U404 (N_404,N_341,N_303);
or U405 (N_405,N_313,N_354);
or U406 (N_406,N_225,N_352);
nand U407 (N_407,N_169,N_369);
and U408 (N_408,N_318,N_128);
nor U409 (N_409,N_371,N_351);
nor U410 (N_410,N_339,N_327);
or U411 (N_411,N_203,N_372);
nor U412 (N_412,N_286,N_193);
nand U413 (N_413,N_306,In_239);
nand U414 (N_414,In_271,N_340);
and U415 (N_415,N_348,N_239);
and U416 (N_416,N_248,N_317);
and U417 (N_417,In_425,N_366);
and U418 (N_418,N_358,In_257);
or U419 (N_419,N_336,N_328);
nand U420 (N_420,In_176,N_311);
and U421 (N_421,N_320,N_315);
nand U422 (N_422,N_368,N_309);
and U423 (N_423,In_152,N_338);
and U424 (N_424,N_178,In_413);
and U425 (N_425,N_361,N_359);
and U426 (N_426,N_312,N_362);
nor U427 (N_427,N_227,N_333);
nand U428 (N_428,N_344,N_116);
or U429 (N_429,N_305,N_319);
or U430 (N_430,N_331,N_332);
or U431 (N_431,N_355,In_427);
and U432 (N_432,N_373,N_345);
xor U433 (N_433,In_218,N_347);
and U434 (N_434,N_364,N_113);
nand U435 (N_435,N_299,N_247);
or U436 (N_436,N_218,N_330);
xnor U437 (N_437,N_357,N_371);
xnor U438 (N_438,N_322,N_371);
and U439 (N_439,N_334,N_193);
nor U440 (N_440,N_364,N_354);
or U441 (N_441,N_253,N_218);
or U442 (N_442,N_313,N_347);
nor U443 (N_443,N_307,N_237);
nand U444 (N_444,N_239,In_257);
nor U445 (N_445,In_318,N_373);
and U446 (N_446,N_333,N_356);
and U447 (N_447,N_349,N_307);
nor U448 (N_448,N_335,N_338);
nor U449 (N_449,N_364,N_331);
nand U450 (N_450,N_433,N_397);
nand U451 (N_451,N_447,N_432);
and U452 (N_452,N_386,N_427);
xnor U453 (N_453,N_377,N_403);
nor U454 (N_454,N_434,N_394);
nand U455 (N_455,N_418,N_429);
nand U456 (N_456,N_446,N_428);
and U457 (N_457,N_420,N_399);
xnor U458 (N_458,N_392,N_405);
xnor U459 (N_459,N_407,N_415);
nor U460 (N_460,N_390,N_402);
or U461 (N_461,N_422,N_381);
nor U462 (N_462,N_417,N_401);
and U463 (N_463,N_435,N_404);
and U464 (N_464,N_388,N_442);
nand U465 (N_465,N_389,N_449);
nor U466 (N_466,N_400,N_436);
nor U467 (N_467,N_426,N_382);
nor U468 (N_468,N_385,N_412);
or U469 (N_469,N_414,N_443);
xor U470 (N_470,N_395,N_376);
nor U471 (N_471,N_387,N_416);
and U472 (N_472,N_413,N_380);
nor U473 (N_473,N_406,N_378);
and U474 (N_474,N_411,N_384);
or U475 (N_475,N_409,N_408);
nand U476 (N_476,N_424,N_430);
or U477 (N_477,N_410,N_419);
nand U478 (N_478,N_448,N_421);
and U479 (N_479,N_379,N_391);
or U480 (N_480,N_439,N_431);
nand U481 (N_481,N_444,N_423);
nand U482 (N_482,N_437,N_383);
xnor U483 (N_483,N_438,N_393);
nand U484 (N_484,N_425,N_441);
xor U485 (N_485,N_375,N_398);
or U486 (N_486,N_396,N_445);
and U487 (N_487,N_440,N_446);
xnor U488 (N_488,N_444,N_410);
and U489 (N_489,N_388,N_413);
or U490 (N_490,N_441,N_380);
or U491 (N_491,N_426,N_431);
xnor U492 (N_492,N_421,N_383);
or U493 (N_493,N_413,N_428);
nor U494 (N_494,N_446,N_432);
xnor U495 (N_495,N_432,N_449);
nor U496 (N_496,N_419,N_420);
nand U497 (N_497,N_399,N_400);
or U498 (N_498,N_412,N_378);
and U499 (N_499,N_432,N_434);
nand U500 (N_500,N_445,N_404);
or U501 (N_501,N_400,N_402);
or U502 (N_502,N_420,N_439);
xnor U503 (N_503,N_409,N_418);
nor U504 (N_504,N_430,N_386);
and U505 (N_505,N_414,N_429);
or U506 (N_506,N_390,N_388);
nand U507 (N_507,N_417,N_447);
nor U508 (N_508,N_446,N_397);
nand U509 (N_509,N_428,N_384);
nand U510 (N_510,N_442,N_407);
nor U511 (N_511,N_405,N_377);
nor U512 (N_512,N_423,N_438);
nand U513 (N_513,N_425,N_378);
and U514 (N_514,N_434,N_435);
xor U515 (N_515,N_409,N_379);
and U516 (N_516,N_432,N_386);
nor U517 (N_517,N_441,N_402);
nor U518 (N_518,N_430,N_406);
or U519 (N_519,N_439,N_416);
and U520 (N_520,N_400,N_412);
or U521 (N_521,N_419,N_416);
nand U522 (N_522,N_425,N_389);
or U523 (N_523,N_389,N_432);
and U524 (N_524,N_388,N_408);
or U525 (N_525,N_504,N_523);
or U526 (N_526,N_519,N_455);
or U527 (N_527,N_482,N_492);
and U528 (N_528,N_489,N_452);
nor U529 (N_529,N_491,N_463);
or U530 (N_530,N_465,N_467);
and U531 (N_531,N_469,N_458);
and U532 (N_532,N_511,N_515);
nand U533 (N_533,N_484,N_490);
nor U534 (N_534,N_468,N_456);
and U535 (N_535,N_501,N_507);
and U536 (N_536,N_518,N_477);
nor U537 (N_537,N_481,N_450);
xor U538 (N_538,N_462,N_510);
and U539 (N_539,N_460,N_497);
nor U540 (N_540,N_459,N_483);
or U541 (N_541,N_505,N_521);
or U542 (N_542,N_499,N_478);
and U543 (N_543,N_457,N_498);
nand U544 (N_544,N_486,N_516);
and U545 (N_545,N_520,N_470);
and U546 (N_546,N_496,N_495);
and U547 (N_547,N_464,N_451);
and U548 (N_548,N_475,N_517);
nor U549 (N_549,N_487,N_509);
nand U550 (N_550,N_500,N_474);
nand U551 (N_551,N_479,N_471);
nand U552 (N_552,N_508,N_514);
xnor U553 (N_553,N_512,N_488);
nor U554 (N_554,N_494,N_454);
nand U555 (N_555,N_522,N_472);
nor U556 (N_556,N_524,N_476);
or U557 (N_557,N_502,N_493);
nand U558 (N_558,N_506,N_473);
nor U559 (N_559,N_513,N_485);
and U560 (N_560,N_453,N_480);
and U561 (N_561,N_466,N_503);
nor U562 (N_562,N_461,N_494);
nor U563 (N_563,N_501,N_450);
nand U564 (N_564,N_497,N_487);
nand U565 (N_565,N_484,N_503);
or U566 (N_566,N_496,N_501);
and U567 (N_567,N_519,N_486);
nand U568 (N_568,N_493,N_483);
nand U569 (N_569,N_486,N_460);
or U570 (N_570,N_455,N_493);
or U571 (N_571,N_510,N_491);
nand U572 (N_572,N_523,N_453);
xnor U573 (N_573,N_481,N_520);
or U574 (N_574,N_489,N_493);
or U575 (N_575,N_510,N_477);
nor U576 (N_576,N_462,N_458);
and U577 (N_577,N_522,N_453);
and U578 (N_578,N_499,N_522);
or U579 (N_579,N_466,N_493);
nand U580 (N_580,N_474,N_480);
nor U581 (N_581,N_521,N_453);
and U582 (N_582,N_468,N_458);
and U583 (N_583,N_476,N_495);
nand U584 (N_584,N_481,N_519);
nor U585 (N_585,N_512,N_501);
xnor U586 (N_586,N_501,N_509);
nor U587 (N_587,N_473,N_515);
nor U588 (N_588,N_463,N_486);
nor U589 (N_589,N_519,N_482);
and U590 (N_590,N_477,N_457);
nand U591 (N_591,N_479,N_496);
xnor U592 (N_592,N_508,N_451);
and U593 (N_593,N_511,N_523);
xnor U594 (N_594,N_476,N_515);
nand U595 (N_595,N_523,N_498);
nor U596 (N_596,N_494,N_476);
xnor U597 (N_597,N_462,N_474);
and U598 (N_598,N_506,N_496);
and U599 (N_599,N_463,N_494);
nor U600 (N_600,N_528,N_584);
or U601 (N_601,N_539,N_552);
or U602 (N_602,N_551,N_564);
or U603 (N_603,N_550,N_529);
or U604 (N_604,N_566,N_570);
nand U605 (N_605,N_571,N_587);
and U606 (N_606,N_560,N_596);
and U607 (N_607,N_592,N_533);
nor U608 (N_608,N_562,N_535);
or U609 (N_609,N_599,N_561);
or U610 (N_610,N_559,N_579);
and U611 (N_611,N_526,N_578);
xor U612 (N_612,N_567,N_591);
or U613 (N_613,N_582,N_577);
or U614 (N_614,N_553,N_540);
or U615 (N_615,N_542,N_537);
or U616 (N_616,N_536,N_574);
or U617 (N_617,N_597,N_545);
nand U618 (N_618,N_530,N_594);
and U619 (N_619,N_590,N_556);
nor U620 (N_620,N_549,N_557);
nor U621 (N_621,N_583,N_569);
or U622 (N_622,N_598,N_593);
or U623 (N_623,N_527,N_558);
nor U624 (N_624,N_580,N_547);
nor U625 (N_625,N_572,N_588);
xnor U626 (N_626,N_581,N_543);
nand U627 (N_627,N_585,N_565);
and U628 (N_628,N_576,N_532);
or U629 (N_629,N_531,N_586);
and U630 (N_630,N_548,N_563);
nor U631 (N_631,N_554,N_589);
nand U632 (N_632,N_575,N_544);
or U633 (N_633,N_555,N_568);
nor U634 (N_634,N_541,N_573);
xor U635 (N_635,N_534,N_525);
or U636 (N_636,N_546,N_595);
nor U637 (N_637,N_538,N_531);
nor U638 (N_638,N_585,N_534);
or U639 (N_639,N_597,N_525);
or U640 (N_640,N_589,N_560);
or U641 (N_641,N_598,N_555);
or U642 (N_642,N_596,N_559);
nor U643 (N_643,N_538,N_540);
or U644 (N_644,N_556,N_535);
or U645 (N_645,N_558,N_567);
and U646 (N_646,N_583,N_551);
nor U647 (N_647,N_577,N_588);
nand U648 (N_648,N_567,N_543);
or U649 (N_649,N_588,N_534);
and U650 (N_650,N_549,N_590);
nor U651 (N_651,N_542,N_556);
or U652 (N_652,N_589,N_563);
nand U653 (N_653,N_567,N_535);
and U654 (N_654,N_532,N_548);
nand U655 (N_655,N_551,N_528);
or U656 (N_656,N_586,N_596);
xor U657 (N_657,N_592,N_565);
nand U658 (N_658,N_557,N_526);
and U659 (N_659,N_597,N_559);
and U660 (N_660,N_538,N_535);
or U661 (N_661,N_566,N_572);
nor U662 (N_662,N_588,N_533);
nor U663 (N_663,N_526,N_558);
nor U664 (N_664,N_570,N_552);
nor U665 (N_665,N_554,N_525);
nand U666 (N_666,N_530,N_590);
or U667 (N_667,N_564,N_552);
nand U668 (N_668,N_553,N_539);
nor U669 (N_669,N_557,N_565);
and U670 (N_670,N_547,N_559);
nand U671 (N_671,N_581,N_530);
nor U672 (N_672,N_588,N_583);
xor U673 (N_673,N_560,N_584);
and U674 (N_674,N_576,N_538);
xor U675 (N_675,N_647,N_639);
nand U676 (N_676,N_608,N_600);
nand U677 (N_677,N_613,N_619);
or U678 (N_678,N_657,N_655);
or U679 (N_679,N_610,N_666);
nor U680 (N_680,N_660,N_603);
nand U681 (N_681,N_605,N_645);
nand U682 (N_682,N_636,N_635);
and U683 (N_683,N_656,N_625);
nand U684 (N_684,N_658,N_626);
xor U685 (N_685,N_620,N_629);
nand U686 (N_686,N_640,N_601);
nor U687 (N_687,N_644,N_643);
nand U688 (N_688,N_641,N_634);
nor U689 (N_689,N_607,N_671);
nand U690 (N_690,N_617,N_632);
nand U691 (N_691,N_668,N_672);
nor U692 (N_692,N_628,N_663);
and U693 (N_693,N_623,N_618);
or U694 (N_694,N_651,N_638);
nor U695 (N_695,N_611,N_630);
nand U696 (N_696,N_653,N_669);
nand U697 (N_697,N_648,N_664);
xnor U698 (N_698,N_612,N_631);
nor U699 (N_699,N_650,N_609);
and U700 (N_700,N_674,N_614);
and U701 (N_701,N_602,N_665);
nor U702 (N_702,N_670,N_662);
nand U703 (N_703,N_621,N_673);
or U704 (N_704,N_661,N_659);
and U705 (N_705,N_646,N_616);
nand U706 (N_706,N_624,N_633);
nor U707 (N_707,N_667,N_652);
or U708 (N_708,N_642,N_615);
xnor U709 (N_709,N_649,N_654);
nand U710 (N_710,N_637,N_627);
and U711 (N_711,N_606,N_622);
and U712 (N_712,N_604,N_612);
nor U713 (N_713,N_665,N_627);
or U714 (N_714,N_601,N_600);
or U715 (N_715,N_657,N_670);
and U716 (N_716,N_635,N_634);
nand U717 (N_717,N_672,N_644);
or U718 (N_718,N_622,N_666);
nor U719 (N_719,N_673,N_641);
nor U720 (N_720,N_656,N_616);
and U721 (N_721,N_674,N_649);
and U722 (N_722,N_667,N_602);
nor U723 (N_723,N_620,N_662);
nand U724 (N_724,N_643,N_656);
nor U725 (N_725,N_621,N_648);
or U726 (N_726,N_621,N_670);
nand U727 (N_727,N_654,N_631);
nand U728 (N_728,N_600,N_647);
nand U729 (N_729,N_614,N_646);
or U730 (N_730,N_644,N_653);
or U731 (N_731,N_604,N_667);
or U732 (N_732,N_642,N_667);
nand U733 (N_733,N_624,N_664);
nand U734 (N_734,N_612,N_649);
nor U735 (N_735,N_639,N_619);
or U736 (N_736,N_607,N_604);
nand U737 (N_737,N_632,N_601);
nor U738 (N_738,N_660,N_649);
and U739 (N_739,N_618,N_605);
nand U740 (N_740,N_648,N_671);
xor U741 (N_741,N_648,N_622);
nand U742 (N_742,N_608,N_609);
and U743 (N_743,N_606,N_611);
and U744 (N_744,N_622,N_639);
and U745 (N_745,N_635,N_660);
nand U746 (N_746,N_642,N_660);
or U747 (N_747,N_652,N_603);
nand U748 (N_748,N_664,N_626);
nor U749 (N_749,N_604,N_625);
and U750 (N_750,N_723,N_675);
nor U751 (N_751,N_710,N_731);
or U752 (N_752,N_748,N_680);
or U753 (N_753,N_724,N_698);
nor U754 (N_754,N_699,N_735);
nand U755 (N_755,N_712,N_742);
and U756 (N_756,N_738,N_719);
nand U757 (N_757,N_708,N_693);
and U758 (N_758,N_703,N_711);
and U759 (N_759,N_716,N_689);
and U760 (N_760,N_688,N_704);
nor U761 (N_761,N_739,N_714);
and U762 (N_762,N_700,N_733);
and U763 (N_763,N_691,N_747);
and U764 (N_764,N_745,N_736);
nor U765 (N_765,N_705,N_702);
nand U766 (N_766,N_717,N_707);
xor U767 (N_767,N_740,N_722);
or U768 (N_768,N_695,N_730);
nand U769 (N_769,N_681,N_718);
nor U770 (N_770,N_679,N_741);
and U771 (N_771,N_732,N_706);
and U772 (N_772,N_697,N_720);
and U773 (N_773,N_726,N_729);
nor U774 (N_774,N_682,N_677);
and U775 (N_775,N_685,N_694);
nand U776 (N_776,N_728,N_713);
nand U777 (N_777,N_725,N_686);
or U778 (N_778,N_678,N_696);
or U779 (N_779,N_683,N_690);
or U780 (N_780,N_715,N_744);
xor U781 (N_781,N_727,N_709);
and U782 (N_782,N_734,N_749);
and U783 (N_783,N_701,N_721);
and U784 (N_784,N_684,N_676);
xnor U785 (N_785,N_743,N_687);
and U786 (N_786,N_737,N_692);
nor U787 (N_787,N_746,N_697);
nor U788 (N_788,N_723,N_721);
xor U789 (N_789,N_700,N_703);
and U790 (N_790,N_733,N_720);
nor U791 (N_791,N_701,N_697);
or U792 (N_792,N_744,N_718);
and U793 (N_793,N_737,N_738);
nand U794 (N_794,N_732,N_747);
or U795 (N_795,N_739,N_702);
xnor U796 (N_796,N_731,N_743);
nor U797 (N_797,N_734,N_714);
nand U798 (N_798,N_706,N_681);
and U799 (N_799,N_733,N_707);
or U800 (N_800,N_695,N_697);
nand U801 (N_801,N_748,N_700);
xnor U802 (N_802,N_680,N_706);
nand U803 (N_803,N_693,N_707);
nand U804 (N_804,N_726,N_689);
nor U805 (N_805,N_718,N_722);
nor U806 (N_806,N_675,N_714);
nand U807 (N_807,N_700,N_711);
and U808 (N_808,N_688,N_721);
or U809 (N_809,N_721,N_745);
nor U810 (N_810,N_704,N_702);
and U811 (N_811,N_738,N_740);
or U812 (N_812,N_683,N_679);
and U813 (N_813,N_746,N_686);
nor U814 (N_814,N_685,N_717);
nor U815 (N_815,N_708,N_744);
nor U816 (N_816,N_682,N_730);
xnor U817 (N_817,N_739,N_744);
and U818 (N_818,N_745,N_718);
nand U819 (N_819,N_717,N_691);
nor U820 (N_820,N_749,N_690);
nand U821 (N_821,N_719,N_679);
or U822 (N_822,N_682,N_694);
and U823 (N_823,N_693,N_697);
or U824 (N_824,N_746,N_703);
nand U825 (N_825,N_799,N_804);
nand U826 (N_826,N_754,N_751);
nor U827 (N_827,N_755,N_802);
or U828 (N_828,N_774,N_797);
or U829 (N_829,N_811,N_764);
xnor U830 (N_830,N_814,N_810);
nand U831 (N_831,N_781,N_801);
nor U832 (N_832,N_790,N_786);
xor U833 (N_833,N_794,N_778);
nor U834 (N_834,N_808,N_758);
or U835 (N_835,N_792,N_793);
and U836 (N_836,N_787,N_779);
and U837 (N_837,N_757,N_818);
or U838 (N_838,N_783,N_767);
or U839 (N_839,N_760,N_776);
and U840 (N_840,N_782,N_772);
nor U841 (N_841,N_800,N_759);
xnor U842 (N_842,N_821,N_807);
or U843 (N_843,N_785,N_775);
nand U844 (N_844,N_773,N_763);
and U845 (N_845,N_756,N_769);
nor U846 (N_846,N_780,N_777);
nand U847 (N_847,N_798,N_753);
and U848 (N_848,N_796,N_750);
and U849 (N_849,N_812,N_813);
and U850 (N_850,N_809,N_823);
or U851 (N_851,N_765,N_771);
xor U852 (N_852,N_768,N_824);
xor U853 (N_853,N_761,N_784);
or U854 (N_854,N_819,N_789);
or U855 (N_855,N_766,N_791);
nor U856 (N_856,N_817,N_770);
and U857 (N_857,N_762,N_806);
or U858 (N_858,N_752,N_820);
nor U859 (N_859,N_795,N_822);
or U860 (N_860,N_816,N_805);
nor U861 (N_861,N_788,N_815);
or U862 (N_862,N_803,N_801);
xnor U863 (N_863,N_750,N_799);
nor U864 (N_864,N_795,N_807);
nor U865 (N_865,N_751,N_762);
and U866 (N_866,N_796,N_807);
nor U867 (N_867,N_819,N_785);
nor U868 (N_868,N_808,N_815);
or U869 (N_869,N_786,N_803);
nor U870 (N_870,N_767,N_751);
nand U871 (N_871,N_800,N_822);
or U872 (N_872,N_755,N_818);
and U873 (N_873,N_752,N_775);
nand U874 (N_874,N_819,N_815);
xor U875 (N_875,N_791,N_755);
nor U876 (N_876,N_789,N_821);
nand U877 (N_877,N_790,N_804);
and U878 (N_878,N_775,N_795);
nand U879 (N_879,N_788,N_761);
xor U880 (N_880,N_769,N_798);
nor U881 (N_881,N_814,N_818);
nand U882 (N_882,N_819,N_804);
nor U883 (N_883,N_758,N_786);
or U884 (N_884,N_807,N_770);
or U885 (N_885,N_752,N_762);
nor U886 (N_886,N_771,N_752);
or U887 (N_887,N_767,N_762);
nor U888 (N_888,N_814,N_756);
nor U889 (N_889,N_794,N_752);
nor U890 (N_890,N_770,N_811);
nor U891 (N_891,N_758,N_789);
nor U892 (N_892,N_750,N_758);
xor U893 (N_893,N_783,N_757);
nor U894 (N_894,N_819,N_756);
nor U895 (N_895,N_795,N_809);
or U896 (N_896,N_799,N_805);
nand U897 (N_897,N_759,N_755);
or U898 (N_898,N_809,N_801);
or U899 (N_899,N_755,N_773);
or U900 (N_900,N_834,N_833);
nand U901 (N_901,N_890,N_830);
or U902 (N_902,N_827,N_845);
or U903 (N_903,N_862,N_851);
or U904 (N_904,N_891,N_835);
nor U905 (N_905,N_870,N_888);
or U906 (N_906,N_874,N_855);
or U907 (N_907,N_825,N_884);
or U908 (N_908,N_886,N_866);
or U909 (N_909,N_899,N_889);
and U910 (N_910,N_864,N_857);
nor U911 (N_911,N_844,N_826);
nor U912 (N_912,N_887,N_876);
nor U913 (N_913,N_877,N_892);
nand U914 (N_914,N_831,N_841);
and U915 (N_915,N_850,N_846);
and U916 (N_916,N_883,N_828);
and U917 (N_917,N_868,N_839);
or U918 (N_918,N_895,N_852);
or U919 (N_919,N_865,N_867);
nor U920 (N_920,N_836,N_842);
nor U921 (N_921,N_881,N_898);
nor U922 (N_922,N_878,N_856);
or U923 (N_923,N_853,N_882);
and U924 (N_924,N_837,N_863);
or U925 (N_925,N_893,N_858);
and U926 (N_926,N_840,N_832);
nor U927 (N_927,N_843,N_869);
nor U928 (N_928,N_838,N_829);
and U929 (N_929,N_879,N_854);
or U930 (N_930,N_897,N_885);
nor U931 (N_931,N_861,N_873);
and U932 (N_932,N_880,N_849);
or U933 (N_933,N_848,N_875);
and U934 (N_934,N_872,N_894);
nand U935 (N_935,N_847,N_896);
and U936 (N_936,N_859,N_860);
and U937 (N_937,N_871,N_855);
nor U938 (N_938,N_882,N_836);
nor U939 (N_939,N_865,N_877);
xor U940 (N_940,N_853,N_893);
nor U941 (N_941,N_894,N_867);
nor U942 (N_942,N_858,N_866);
or U943 (N_943,N_843,N_863);
or U944 (N_944,N_832,N_856);
and U945 (N_945,N_899,N_878);
nor U946 (N_946,N_854,N_826);
and U947 (N_947,N_833,N_847);
nor U948 (N_948,N_841,N_890);
nand U949 (N_949,N_898,N_888);
and U950 (N_950,N_893,N_841);
nand U951 (N_951,N_854,N_893);
nand U952 (N_952,N_861,N_899);
or U953 (N_953,N_866,N_837);
xnor U954 (N_954,N_863,N_891);
and U955 (N_955,N_859,N_844);
nand U956 (N_956,N_867,N_848);
or U957 (N_957,N_835,N_863);
nor U958 (N_958,N_882,N_840);
or U959 (N_959,N_846,N_834);
nand U960 (N_960,N_879,N_839);
nand U961 (N_961,N_844,N_850);
and U962 (N_962,N_887,N_870);
nand U963 (N_963,N_862,N_876);
or U964 (N_964,N_875,N_888);
nor U965 (N_965,N_858,N_837);
xor U966 (N_966,N_874,N_890);
or U967 (N_967,N_878,N_896);
or U968 (N_968,N_868,N_858);
xor U969 (N_969,N_888,N_828);
and U970 (N_970,N_849,N_889);
nor U971 (N_971,N_879,N_844);
or U972 (N_972,N_825,N_891);
nor U973 (N_973,N_848,N_880);
nand U974 (N_974,N_876,N_881);
nand U975 (N_975,N_924,N_950);
nand U976 (N_976,N_928,N_964);
nor U977 (N_977,N_919,N_945);
and U978 (N_978,N_901,N_915);
nor U979 (N_979,N_908,N_937);
xnor U980 (N_980,N_943,N_947);
and U981 (N_981,N_960,N_955);
nand U982 (N_982,N_935,N_916);
or U983 (N_983,N_949,N_904);
or U984 (N_984,N_923,N_951);
nor U985 (N_985,N_953,N_927);
or U986 (N_986,N_938,N_962);
nand U987 (N_987,N_914,N_940);
nand U988 (N_988,N_965,N_948);
xnor U989 (N_989,N_925,N_946);
and U990 (N_990,N_903,N_918);
or U991 (N_991,N_972,N_929);
nand U992 (N_992,N_966,N_963);
or U993 (N_993,N_930,N_917);
nand U994 (N_994,N_968,N_933);
nand U995 (N_995,N_974,N_952);
nand U996 (N_996,N_922,N_939);
nand U997 (N_997,N_909,N_971);
and U998 (N_998,N_958,N_913);
or U999 (N_999,N_973,N_931);
nor U1000 (N_1000,N_912,N_905);
xor U1001 (N_1001,N_970,N_920);
xor U1002 (N_1002,N_959,N_954);
or U1003 (N_1003,N_934,N_936);
or U1004 (N_1004,N_902,N_900);
nor U1005 (N_1005,N_907,N_957);
and U1006 (N_1006,N_932,N_967);
nand U1007 (N_1007,N_969,N_944);
nor U1008 (N_1008,N_941,N_921);
nand U1009 (N_1009,N_910,N_926);
nand U1010 (N_1010,N_911,N_906);
nand U1011 (N_1011,N_956,N_961);
nand U1012 (N_1012,N_942,N_918);
and U1013 (N_1013,N_952,N_931);
nand U1014 (N_1014,N_911,N_916);
or U1015 (N_1015,N_929,N_957);
and U1016 (N_1016,N_946,N_974);
or U1017 (N_1017,N_959,N_932);
and U1018 (N_1018,N_971,N_906);
and U1019 (N_1019,N_947,N_919);
nor U1020 (N_1020,N_909,N_933);
nand U1021 (N_1021,N_919,N_933);
nand U1022 (N_1022,N_937,N_920);
or U1023 (N_1023,N_944,N_953);
nand U1024 (N_1024,N_912,N_910);
nor U1025 (N_1025,N_916,N_921);
and U1026 (N_1026,N_972,N_953);
nand U1027 (N_1027,N_971,N_962);
or U1028 (N_1028,N_926,N_961);
and U1029 (N_1029,N_969,N_929);
xor U1030 (N_1030,N_968,N_950);
nand U1031 (N_1031,N_972,N_932);
xnor U1032 (N_1032,N_908,N_902);
or U1033 (N_1033,N_900,N_903);
or U1034 (N_1034,N_948,N_906);
and U1035 (N_1035,N_943,N_909);
nand U1036 (N_1036,N_906,N_956);
nor U1037 (N_1037,N_966,N_933);
nand U1038 (N_1038,N_935,N_964);
or U1039 (N_1039,N_949,N_947);
nand U1040 (N_1040,N_928,N_952);
xor U1041 (N_1041,N_913,N_965);
or U1042 (N_1042,N_972,N_962);
and U1043 (N_1043,N_931,N_911);
nand U1044 (N_1044,N_936,N_928);
nor U1045 (N_1045,N_939,N_957);
and U1046 (N_1046,N_901,N_947);
nand U1047 (N_1047,N_908,N_950);
nand U1048 (N_1048,N_937,N_925);
nand U1049 (N_1049,N_920,N_962);
and U1050 (N_1050,N_1012,N_1024);
and U1051 (N_1051,N_1042,N_988);
or U1052 (N_1052,N_980,N_1038);
or U1053 (N_1053,N_993,N_1044);
or U1054 (N_1054,N_1014,N_982);
nand U1055 (N_1055,N_984,N_999);
nor U1056 (N_1056,N_1015,N_1039);
or U1057 (N_1057,N_1046,N_1035);
nand U1058 (N_1058,N_1031,N_991);
or U1059 (N_1059,N_1000,N_1040);
nand U1060 (N_1060,N_1020,N_1048);
or U1061 (N_1061,N_1017,N_1008);
or U1062 (N_1062,N_983,N_1034);
nand U1063 (N_1063,N_986,N_1018);
or U1064 (N_1064,N_1003,N_976);
nand U1065 (N_1065,N_985,N_1036);
nand U1066 (N_1066,N_995,N_1033);
nor U1067 (N_1067,N_1006,N_996);
nor U1068 (N_1068,N_1045,N_1025);
nand U1069 (N_1069,N_981,N_1026);
nand U1070 (N_1070,N_998,N_1016);
nor U1071 (N_1071,N_1010,N_1011);
xor U1072 (N_1072,N_990,N_1047);
nand U1073 (N_1073,N_1049,N_1032);
or U1074 (N_1074,N_1009,N_1002);
nor U1075 (N_1075,N_1007,N_1028);
nand U1076 (N_1076,N_987,N_1030);
and U1077 (N_1077,N_1013,N_1022);
nand U1078 (N_1078,N_1041,N_1019);
or U1079 (N_1079,N_1004,N_1021);
nor U1080 (N_1080,N_975,N_989);
or U1081 (N_1081,N_1001,N_1027);
and U1082 (N_1082,N_979,N_978);
xnor U1083 (N_1083,N_1029,N_1037);
nand U1084 (N_1084,N_994,N_997);
nand U1085 (N_1085,N_992,N_977);
or U1086 (N_1086,N_1005,N_1023);
and U1087 (N_1087,N_1043,N_1004);
and U1088 (N_1088,N_1033,N_1005);
xnor U1089 (N_1089,N_990,N_1001);
nor U1090 (N_1090,N_975,N_1035);
and U1091 (N_1091,N_993,N_1015);
nor U1092 (N_1092,N_1014,N_983);
xnor U1093 (N_1093,N_1020,N_1018);
or U1094 (N_1094,N_1039,N_1035);
xor U1095 (N_1095,N_1037,N_981);
and U1096 (N_1096,N_1020,N_1038);
and U1097 (N_1097,N_982,N_976);
or U1098 (N_1098,N_1033,N_988);
and U1099 (N_1099,N_976,N_975);
and U1100 (N_1100,N_1030,N_993);
nand U1101 (N_1101,N_1018,N_1000);
xor U1102 (N_1102,N_1049,N_1003);
xor U1103 (N_1103,N_1013,N_1028);
nand U1104 (N_1104,N_1009,N_1026);
or U1105 (N_1105,N_976,N_993);
nand U1106 (N_1106,N_983,N_997);
nand U1107 (N_1107,N_1049,N_1037);
nor U1108 (N_1108,N_1033,N_1013);
or U1109 (N_1109,N_1014,N_975);
nand U1110 (N_1110,N_993,N_1040);
nor U1111 (N_1111,N_988,N_1001);
and U1112 (N_1112,N_989,N_1012);
xnor U1113 (N_1113,N_990,N_992);
nand U1114 (N_1114,N_1046,N_996);
or U1115 (N_1115,N_1007,N_1032);
nor U1116 (N_1116,N_991,N_1049);
nor U1117 (N_1117,N_980,N_1028);
nor U1118 (N_1118,N_1019,N_1009);
and U1119 (N_1119,N_991,N_1032);
xor U1120 (N_1120,N_1042,N_993);
and U1121 (N_1121,N_1018,N_1026);
xor U1122 (N_1122,N_1039,N_1021);
or U1123 (N_1123,N_1036,N_1012);
or U1124 (N_1124,N_1010,N_997);
and U1125 (N_1125,N_1091,N_1114);
nand U1126 (N_1126,N_1121,N_1090);
or U1127 (N_1127,N_1122,N_1088);
and U1128 (N_1128,N_1120,N_1105);
or U1129 (N_1129,N_1124,N_1115);
nand U1130 (N_1130,N_1110,N_1083);
nor U1131 (N_1131,N_1109,N_1078);
and U1132 (N_1132,N_1064,N_1094);
and U1133 (N_1133,N_1074,N_1084);
nor U1134 (N_1134,N_1066,N_1111);
nand U1135 (N_1135,N_1076,N_1060);
and U1136 (N_1136,N_1059,N_1063);
nand U1137 (N_1137,N_1068,N_1051);
nor U1138 (N_1138,N_1101,N_1099);
nor U1139 (N_1139,N_1055,N_1065);
nand U1140 (N_1140,N_1070,N_1100);
and U1141 (N_1141,N_1097,N_1058);
xnor U1142 (N_1142,N_1102,N_1103);
and U1143 (N_1143,N_1081,N_1050);
and U1144 (N_1144,N_1113,N_1112);
xor U1145 (N_1145,N_1107,N_1093);
nand U1146 (N_1146,N_1073,N_1096);
nor U1147 (N_1147,N_1098,N_1057);
nand U1148 (N_1148,N_1069,N_1123);
and U1149 (N_1149,N_1061,N_1054);
nand U1150 (N_1150,N_1082,N_1095);
xnor U1151 (N_1151,N_1072,N_1075);
or U1152 (N_1152,N_1079,N_1056);
nand U1153 (N_1153,N_1106,N_1116);
and U1154 (N_1154,N_1117,N_1085);
nand U1155 (N_1155,N_1118,N_1104);
or U1156 (N_1156,N_1080,N_1108);
nor U1157 (N_1157,N_1071,N_1086);
and U1158 (N_1158,N_1089,N_1067);
and U1159 (N_1159,N_1062,N_1052);
nor U1160 (N_1160,N_1087,N_1053);
nor U1161 (N_1161,N_1119,N_1077);
and U1162 (N_1162,N_1092,N_1052);
or U1163 (N_1163,N_1056,N_1084);
nor U1164 (N_1164,N_1112,N_1117);
and U1165 (N_1165,N_1122,N_1107);
xor U1166 (N_1166,N_1111,N_1112);
and U1167 (N_1167,N_1063,N_1070);
nand U1168 (N_1168,N_1092,N_1075);
xor U1169 (N_1169,N_1113,N_1073);
nor U1170 (N_1170,N_1120,N_1050);
nor U1171 (N_1171,N_1101,N_1056);
and U1172 (N_1172,N_1059,N_1080);
nor U1173 (N_1173,N_1076,N_1071);
nand U1174 (N_1174,N_1084,N_1124);
nand U1175 (N_1175,N_1084,N_1063);
and U1176 (N_1176,N_1096,N_1122);
xor U1177 (N_1177,N_1073,N_1057);
or U1178 (N_1178,N_1110,N_1106);
or U1179 (N_1179,N_1110,N_1107);
or U1180 (N_1180,N_1078,N_1107);
nand U1181 (N_1181,N_1059,N_1094);
nor U1182 (N_1182,N_1085,N_1099);
nor U1183 (N_1183,N_1085,N_1083);
or U1184 (N_1184,N_1104,N_1100);
nor U1185 (N_1185,N_1105,N_1090);
and U1186 (N_1186,N_1085,N_1062);
or U1187 (N_1187,N_1117,N_1101);
or U1188 (N_1188,N_1107,N_1080);
nand U1189 (N_1189,N_1101,N_1058);
and U1190 (N_1190,N_1119,N_1078);
nand U1191 (N_1191,N_1075,N_1056);
and U1192 (N_1192,N_1088,N_1072);
and U1193 (N_1193,N_1093,N_1072);
nor U1194 (N_1194,N_1088,N_1059);
nand U1195 (N_1195,N_1094,N_1122);
or U1196 (N_1196,N_1104,N_1098);
or U1197 (N_1197,N_1055,N_1066);
nor U1198 (N_1198,N_1112,N_1085);
xor U1199 (N_1199,N_1050,N_1085);
and U1200 (N_1200,N_1129,N_1142);
or U1201 (N_1201,N_1180,N_1127);
and U1202 (N_1202,N_1195,N_1161);
and U1203 (N_1203,N_1130,N_1143);
nand U1204 (N_1204,N_1136,N_1137);
xor U1205 (N_1205,N_1169,N_1198);
or U1206 (N_1206,N_1128,N_1135);
or U1207 (N_1207,N_1189,N_1164);
nor U1208 (N_1208,N_1176,N_1186);
or U1209 (N_1209,N_1182,N_1192);
and U1210 (N_1210,N_1144,N_1184);
xnor U1211 (N_1211,N_1185,N_1152);
xnor U1212 (N_1212,N_1149,N_1181);
nand U1213 (N_1213,N_1125,N_1183);
or U1214 (N_1214,N_1179,N_1158);
nand U1215 (N_1215,N_1190,N_1154);
xnor U1216 (N_1216,N_1132,N_1162);
and U1217 (N_1217,N_1168,N_1146);
or U1218 (N_1218,N_1150,N_1171);
and U1219 (N_1219,N_1191,N_1174);
nand U1220 (N_1220,N_1145,N_1147);
nand U1221 (N_1221,N_1133,N_1170);
nor U1222 (N_1222,N_1138,N_1166);
or U1223 (N_1223,N_1153,N_1193);
or U1224 (N_1224,N_1134,N_1178);
and U1225 (N_1225,N_1167,N_1177);
nand U1226 (N_1226,N_1160,N_1126);
and U1227 (N_1227,N_1156,N_1199);
nand U1228 (N_1228,N_1163,N_1148);
and U1229 (N_1229,N_1188,N_1131);
nand U1230 (N_1230,N_1172,N_1196);
nor U1231 (N_1231,N_1155,N_1197);
nand U1232 (N_1232,N_1194,N_1187);
nor U1233 (N_1233,N_1140,N_1159);
xor U1234 (N_1234,N_1151,N_1173);
and U1235 (N_1235,N_1141,N_1157);
nand U1236 (N_1236,N_1139,N_1175);
nor U1237 (N_1237,N_1165,N_1156);
or U1238 (N_1238,N_1132,N_1181);
or U1239 (N_1239,N_1183,N_1146);
or U1240 (N_1240,N_1129,N_1150);
nand U1241 (N_1241,N_1157,N_1128);
nand U1242 (N_1242,N_1183,N_1156);
or U1243 (N_1243,N_1126,N_1171);
nor U1244 (N_1244,N_1196,N_1138);
and U1245 (N_1245,N_1186,N_1178);
nor U1246 (N_1246,N_1132,N_1184);
or U1247 (N_1247,N_1140,N_1157);
nor U1248 (N_1248,N_1145,N_1191);
nor U1249 (N_1249,N_1195,N_1157);
and U1250 (N_1250,N_1170,N_1165);
nand U1251 (N_1251,N_1129,N_1192);
nor U1252 (N_1252,N_1151,N_1155);
xor U1253 (N_1253,N_1133,N_1156);
and U1254 (N_1254,N_1162,N_1126);
and U1255 (N_1255,N_1151,N_1142);
xnor U1256 (N_1256,N_1199,N_1133);
nor U1257 (N_1257,N_1179,N_1152);
xor U1258 (N_1258,N_1133,N_1128);
and U1259 (N_1259,N_1182,N_1145);
xnor U1260 (N_1260,N_1134,N_1153);
or U1261 (N_1261,N_1161,N_1150);
nand U1262 (N_1262,N_1135,N_1125);
nor U1263 (N_1263,N_1167,N_1138);
nand U1264 (N_1264,N_1126,N_1174);
and U1265 (N_1265,N_1141,N_1127);
and U1266 (N_1266,N_1126,N_1168);
nor U1267 (N_1267,N_1158,N_1166);
or U1268 (N_1268,N_1138,N_1154);
or U1269 (N_1269,N_1172,N_1156);
nor U1270 (N_1270,N_1179,N_1159);
nand U1271 (N_1271,N_1165,N_1150);
or U1272 (N_1272,N_1150,N_1145);
nand U1273 (N_1273,N_1126,N_1133);
and U1274 (N_1274,N_1146,N_1162);
and U1275 (N_1275,N_1250,N_1225);
or U1276 (N_1276,N_1215,N_1272);
or U1277 (N_1277,N_1253,N_1263);
nor U1278 (N_1278,N_1268,N_1213);
and U1279 (N_1279,N_1223,N_1258);
nand U1280 (N_1280,N_1243,N_1202);
xor U1281 (N_1281,N_1214,N_1230);
nor U1282 (N_1282,N_1209,N_1246);
nor U1283 (N_1283,N_1255,N_1231);
and U1284 (N_1284,N_1249,N_1247);
nor U1285 (N_1285,N_1204,N_1203);
nor U1286 (N_1286,N_1236,N_1242);
nor U1287 (N_1287,N_1219,N_1221);
nand U1288 (N_1288,N_1251,N_1265);
nand U1289 (N_1289,N_1208,N_1254);
and U1290 (N_1290,N_1257,N_1228);
nor U1291 (N_1291,N_1205,N_1274);
or U1292 (N_1292,N_1267,N_1248);
and U1293 (N_1293,N_1232,N_1207);
xnor U1294 (N_1294,N_1212,N_1262);
and U1295 (N_1295,N_1238,N_1234);
and U1296 (N_1296,N_1220,N_1222);
and U1297 (N_1297,N_1271,N_1269);
xor U1298 (N_1298,N_1260,N_1211);
or U1299 (N_1299,N_1245,N_1229);
xor U1300 (N_1300,N_1235,N_1226);
and U1301 (N_1301,N_1256,N_1244);
nor U1302 (N_1302,N_1216,N_1270);
and U1303 (N_1303,N_1206,N_1233);
nor U1304 (N_1304,N_1210,N_1264);
and U1305 (N_1305,N_1224,N_1252);
or U1306 (N_1306,N_1266,N_1239);
and U1307 (N_1307,N_1241,N_1200);
and U1308 (N_1308,N_1261,N_1259);
and U1309 (N_1309,N_1237,N_1227);
nor U1310 (N_1310,N_1217,N_1240);
and U1311 (N_1311,N_1273,N_1201);
nand U1312 (N_1312,N_1218,N_1272);
or U1313 (N_1313,N_1228,N_1238);
nor U1314 (N_1314,N_1250,N_1265);
or U1315 (N_1315,N_1266,N_1267);
nand U1316 (N_1316,N_1259,N_1203);
xnor U1317 (N_1317,N_1221,N_1238);
nor U1318 (N_1318,N_1255,N_1238);
nand U1319 (N_1319,N_1234,N_1218);
xnor U1320 (N_1320,N_1260,N_1249);
and U1321 (N_1321,N_1255,N_1212);
or U1322 (N_1322,N_1238,N_1254);
or U1323 (N_1323,N_1205,N_1265);
and U1324 (N_1324,N_1230,N_1207);
nor U1325 (N_1325,N_1248,N_1240);
and U1326 (N_1326,N_1257,N_1203);
and U1327 (N_1327,N_1227,N_1217);
or U1328 (N_1328,N_1258,N_1239);
nand U1329 (N_1329,N_1274,N_1213);
xnor U1330 (N_1330,N_1253,N_1227);
xnor U1331 (N_1331,N_1245,N_1231);
and U1332 (N_1332,N_1224,N_1259);
and U1333 (N_1333,N_1260,N_1254);
nand U1334 (N_1334,N_1206,N_1213);
and U1335 (N_1335,N_1244,N_1246);
nand U1336 (N_1336,N_1236,N_1227);
nand U1337 (N_1337,N_1214,N_1200);
and U1338 (N_1338,N_1224,N_1216);
and U1339 (N_1339,N_1263,N_1238);
and U1340 (N_1340,N_1227,N_1231);
nand U1341 (N_1341,N_1270,N_1240);
or U1342 (N_1342,N_1214,N_1247);
and U1343 (N_1343,N_1223,N_1243);
nor U1344 (N_1344,N_1245,N_1214);
or U1345 (N_1345,N_1254,N_1200);
or U1346 (N_1346,N_1209,N_1263);
and U1347 (N_1347,N_1260,N_1248);
and U1348 (N_1348,N_1244,N_1265);
nor U1349 (N_1349,N_1265,N_1270);
nand U1350 (N_1350,N_1277,N_1348);
or U1351 (N_1351,N_1284,N_1275);
nand U1352 (N_1352,N_1282,N_1292);
nand U1353 (N_1353,N_1318,N_1299);
nor U1354 (N_1354,N_1293,N_1312);
nor U1355 (N_1355,N_1339,N_1304);
xnor U1356 (N_1356,N_1332,N_1290);
nor U1357 (N_1357,N_1280,N_1346);
or U1358 (N_1358,N_1337,N_1333);
nor U1359 (N_1359,N_1307,N_1345);
nand U1360 (N_1360,N_1326,N_1287);
and U1361 (N_1361,N_1310,N_1283);
or U1362 (N_1362,N_1328,N_1316);
xor U1363 (N_1363,N_1330,N_1279);
or U1364 (N_1364,N_1303,N_1334);
nand U1365 (N_1365,N_1296,N_1329);
and U1366 (N_1366,N_1321,N_1327);
and U1367 (N_1367,N_1347,N_1340);
or U1368 (N_1368,N_1317,N_1331);
nor U1369 (N_1369,N_1324,N_1349);
and U1370 (N_1370,N_1295,N_1276);
nand U1371 (N_1371,N_1342,N_1281);
nor U1372 (N_1372,N_1308,N_1291);
nor U1373 (N_1373,N_1344,N_1322);
nor U1374 (N_1374,N_1314,N_1320);
or U1375 (N_1375,N_1323,N_1300);
and U1376 (N_1376,N_1302,N_1278);
or U1377 (N_1377,N_1305,N_1298);
nand U1378 (N_1378,N_1338,N_1341);
and U1379 (N_1379,N_1311,N_1289);
xnor U1380 (N_1380,N_1319,N_1285);
and U1381 (N_1381,N_1301,N_1343);
or U1382 (N_1382,N_1297,N_1286);
xor U1383 (N_1383,N_1325,N_1294);
or U1384 (N_1384,N_1335,N_1336);
and U1385 (N_1385,N_1309,N_1288);
nor U1386 (N_1386,N_1306,N_1315);
nand U1387 (N_1387,N_1313,N_1282);
nand U1388 (N_1388,N_1280,N_1331);
xnor U1389 (N_1389,N_1317,N_1285);
or U1390 (N_1390,N_1308,N_1336);
nor U1391 (N_1391,N_1334,N_1338);
and U1392 (N_1392,N_1327,N_1329);
and U1393 (N_1393,N_1293,N_1289);
nor U1394 (N_1394,N_1276,N_1275);
and U1395 (N_1395,N_1299,N_1275);
and U1396 (N_1396,N_1288,N_1287);
nand U1397 (N_1397,N_1294,N_1285);
nand U1398 (N_1398,N_1330,N_1280);
nand U1399 (N_1399,N_1348,N_1281);
or U1400 (N_1400,N_1307,N_1337);
nor U1401 (N_1401,N_1296,N_1338);
or U1402 (N_1402,N_1285,N_1315);
or U1403 (N_1403,N_1279,N_1308);
or U1404 (N_1404,N_1325,N_1315);
xnor U1405 (N_1405,N_1347,N_1342);
nand U1406 (N_1406,N_1280,N_1309);
nor U1407 (N_1407,N_1336,N_1299);
nor U1408 (N_1408,N_1322,N_1328);
nand U1409 (N_1409,N_1283,N_1290);
nand U1410 (N_1410,N_1289,N_1332);
nor U1411 (N_1411,N_1293,N_1275);
or U1412 (N_1412,N_1311,N_1298);
or U1413 (N_1413,N_1343,N_1313);
nor U1414 (N_1414,N_1331,N_1282);
nand U1415 (N_1415,N_1348,N_1334);
nor U1416 (N_1416,N_1281,N_1286);
and U1417 (N_1417,N_1343,N_1310);
and U1418 (N_1418,N_1281,N_1339);
or U1419 (N_1419,N_1325,N_1278);
nor U1420 (N_1420,N_1283,N_1287);
nand U1421 (N_1421,N_1327,N_1296);
or U1422 (N_1422,N_1315,N_1276);
nand U1423 (N_1423,N_1302,N_1323);
nand U1424 (N_1424,N_1302,N_1291);
nor U1425 (N_1425,N_1358,N_1403);
nand U1426 (N_1426,N_1357,N_1359);
nor U1427 (N_1427,N_1394,N_1384);
and U1428 (N_1428,N_1354,N_1410);
or U1429 (N_1429,N_1414,N_1383);
nor U1430 (N_1430,N_1366,N_1371);
and U1431 (N_1431,N_1395,N_1405);
nand U1432 (N_1432,N_1377,N_1421);
or U1433 (N_1433,N_1364,N_1417);
or U1434 (N_1434,N_1422,N_1350);
nand U1435 (N_1435,N_1373,N_1396);
nor U1436 (N_1436,N_1352,N_1398);
nor U1437 (N_1437,N_1355,N_1390);
and U1438 (N_1438,N_1391,N_1416);
nor U1439 (N_1439,N_1356,N_1420);
nand U1440 (N_1440,N_1389,N_1388);
and U1441 (N_1441,N_1353,N_1368);
or U1442 (N_1442,N_1419,N_1406);
or U1443 (N_1443,N_1412,N_1404);
nand U1444 (N_1444,N_1411,N_1408);
nand U1445 (N_1445,N_1363,N_1379);
and U1446 (N_1446,N_1351,N_1374);
or U1447 (N_1447,N_1392,N_1380);
or U1448 (N_1448,N_1369,N_1381);
nor U1449 (N_1449,N_1401,N_1407);
and U1450 (N_1450,N_1386,N_1365);
nand U1451 (N_1451,N_1370,N_1378);
and U1452 (N_1452,N_1360,N_1376);
nor U1453 (N_1453,N_1385,N_1415);
nand U1454 (N_1454,N_1400,N_1382);
nand U1455 (N_1455,N_1387,N_1361);
or U1456 (N_1456,N_1372,N_1424);
or U1457 (N_1457,N_1397,N_1402);
and U1458 (N_1458,N_1393,N_1423);
and U1459 (N_1459,N_1409,N_1413);
or U1460 (N_1460,N_1399,N_1362);
nor U1461 (N_1461,N_1418,N_1375);
or U1462 (N_1462,N_1367,N_1399);
and U1463 (N_1463,N_1388,N_1422);
nand U1464 (N_1464,N_1371,N_1397);
and U1465 (N_1465,N_1415,N_1414);
nand U1466 (N_1466,N_1409,N_1382);
nand U1467 (N_1467,N_1407,N_1354);
and U1468 (N_1468,N_1421,N_1419);
and U1469 (N_1469,N_1416,N_1350);
and U1470 (N_1470,N_1407,N_1373);
and U1471 (N_1471,N_1366,N_1395);
or U1472 (N_1472,N_1376,N_1387);
and U1473 (N_1473,N_1351,N_1407);
nand U1474 (N_1474,N_1357,N_1387);
nor U1475 (N_1475,N_1385,N_1409);
nand U1476 (N_1476,N_1378,N_1364);
and U1477 (N_1477,N_1402,N_1379);
or U1478 (N_1478,N_1387,N_1399);
nor U1479 (N_1479,N_1365,N_1380);
nand U1480 (N_1480,N_1405,N_1394);
and U1481 (N_1481,N_1422,N_1402);
and U1482 (N_1482,N_1390,N_1421);
nand U1483 (N_1483,N_1423,N_1365);
and U1484 (N_1484,N_1405,N_1421);
or U1485 (N_1485,N_1356,N_1364);
and U1486 (N_1486,N_1366,N_1417);
and U1487 (N_1487,N_1350,N_1398);
nor U1488 (N_1488,N_1384,N_1422);
nor U1489 (N_1489,N_1358,N_1417);
nor U1490 (N_1490,N_1386,N_1411);
nor U1491 (N_1491,N_1384,N_1420);
nor U1492 (N_1492,N_1358,N_1410);
or U1493 (N_1493,N_1359,N_1413);
or U1494 (N_1494,N_1357,N_1406);
xnor U1495 (N_1495,N_1410,N_1378);
nor U1496 (N_1496,N_1360,N_1390);
nor U1497 (N_1497,N_1399,N_1413);
nor U1498 (N_1498,N_1357,N_1378);
and U1499 (N_1499,N_1386,N_1417);
and U1500 (N_1500,N_1446,N_1451);
or U1501 (N_1501,N_1480,N_1489);
nor U1502 (N_1502,N_1431,N_1455);
xnor U1503 (N_1503,N_1433,N_1436);
nor U1504 (N_1504,N_1485,N_1430);
and U1505 (N_1505,N_1432,N_1435);
nand U1506 (N_1506,N_1457,N_1466);
or U1507 (N_1507,N_1439,N_1498);
nand U1508 (N_1508,N_1488,N_1444);
nor U1509 (N_1509,N_1456,N_1499);
or U1510 (N_1510,N_1450,N_1458);
and U1511 (N_1511,N_1441,N_1461);
xnor U1512 (N_1512,N_1464,N_1484);
nand U1513 (N_1513,N_1495,N_1448);
and U1514 (N_1514,N_1438,N_1453);
nor U1515 (N_1515,N_1469,N_1496);
nand U1516 (N_1516,N_1473,N_1465);
and U1517 (N_1517,N_1478,N_1427);
or U1518 (N_1518,N_1463,N_1447);
xnor U1519 (N_1519,N_1491,N_1476);
xnor U1520 (N_1520,N_1493,N_1490);
nor U1521 (N_1521,N_1486,N_1477);
nand U1522 (N_1522,N_1487,N_1471);
or U1523 (N_1523,N_1497,N_1470);
or U1524 (N_1524,N_1462,N_1483);
nor U1525 (N_1525,N_1475,N_1426);
nand U1526 (N_1526,N_1429,N_1474);
or U1527 (N_1527,N_1482,N_1460);
or U1528 (N_1528,N_1449,N_1481);
nor U1529 (N_1529,N_1437,N_1472);
nand U1530 (N_1530,N_1442,N_1459);
nand U1531 (N_1531,N_1468,N_1425);
and U1532 (N_1532,N_1434,N_1494);
and U1533 (N_1533,N_1479,N_1440);
and U1534 (N_1534,N_1467,N_1445);
or U1535 (N_1535,N_1454,N_1452);
or U1536 (N_1536,N_1428,N_1443);
nor U1537 (N_1537,N_1492,N_1435);
or U1538 (N_1538,N_1428,N_1495);
nand U1539 (N_1539,N_1434,N_1425);
or U1540 (N_1540,N_1452,N_1447);
and U1541 (N_1541,N_1432,N_1448);
and U1542 (N_1542,N_1428,N_1451);
and U1543 (N_1543,N_1473,N_1441);
xor U1544 (N_1544,N_1438,N_1471);
nand U1545 (N_1545,N_1450,N_1479);
xnor U1546 (N_1546,N_1480,N_1442);
nand U1547 (N_1547,N_1488,N_1485);
nor U1548 (N_1548,N_1487,N_1431);
or U1549 (N_1549,N_1465,N_1479);
and U1550 (N_1550,N_1471,N_1492);
nor U1551 (N_1551,N_1461,N_1471);
nand U1552 (N_1552,N_1481,N_1498);
nand U1553 (N_1553,N_1463,N_1476);
nor U1554 (N_1554,N_1493,N_1462);
or U1555 (N_1555,N_1461,N_1478);
and U1556 (N_1556,N_1479,N_1438);
nor U1557 (N_1557,N_1451,N_1472);
xnor U1558 (N_1558,N_1470,N_1437);
xor U1559 (N_1559,N_1497,N_1466);
xor U1560 (N_1560,N_1483,N_1484);
nand U1561 (N_1561,N_1469,N_1475);
or U1562 (N_1562,N_1461,N_1446);
nand U1563 (N_1563,N_1471,N_1430);
nand U1564 (N_1564,N_1461,N_1458);
nor U1565 (N_1565,N_1458,N_1495);
or U1566 (N_1566,N_1491,N_1470);
nand U1567 (N_1567,N_1477,N_1442);
or U1568 (N_1568,N_1453,N_1436);
nor U1569 (N_1569,N_1467,N_1448);
xnor U1570 (N_1570,N_1487,N_1430);
nand U1571 (N_1571,N_1436,N_1482);
or U1572 (N_1572,N_1484,N_1482);
and U1573 (N_1573,N_1485,N_1429);
nand U1574 (N_1574,N_1439,N_1441);
xor U1575 (N_1575,N_1511,N_1554);
nand U1576 (N_1576,N_1528,N_1501);
or U1577 (N_1577,N_1564,N_1571);
nor U1578 (N_1578,N_1562,N_1525);
nand U1579 (N_1579,N_1503,N_1539);
or U1580 (N_1580,N_1573,N_1533);
and U1581 (N_1581,N_1536,N_1561);
and U1582 (N_1582,N_1506,N_1552);
and U1583 (N_1583,N_1568,N_1548);
nand U1584 (N_1584,N_1553,N_1518);
or U1585 (N_1585,N_1569,N_1523);
and U1586 (N_1586,N_1534,N_1517);
and U1587 (N_1587,N_1566,N_1530);
and U1588 (N_1588,N_1547,N_1500);
and U1589 (N_1589,N_1551,N_1549);
xnor U1590 (N_1590,N_1559,N_1529);
or U1591 (N_1591,N_1509,N_1520);
and U1592 (N_1592,N_1557,N_1516);
or U1593 (N_1593,N_1572,N_1574);
and U1594 (N_1594,N_1512,N_1550);
or U1595 (N_1595,N_1543,N_1541);
or U1596 (N_1596,N_1527,N_1519);
xnor U1597 (N_1597,N_1555,N_1514);
and U1598 (N_1598,N_1510,N_1535);
nand U1599 (N_1599,N_1565,N_1542);
or U1600 (N_1600,N_1502,N_1545);
nor U1601 (N_1601,N_1532,N_1556);
and U1602 (N_1602,N_1563,N_1546);
nor U1603 (N_1603,N_1540,N_1513);
or U1604 (N_1604,N_1526,N_1567);
and U1605 (N_1605,N_1570,N_1538);
or U1606 (N_1606,N_1521,N_1524);
or U1607 (N_1607,N_1515,N_1531);
and U1608 (N_1608,N_1544,N_1505);
xor U1609 (N_1609,N_1504,N_1507);
and U1610 (N_1610,N_1537,N_1558);
and U1611 (N_1611,N_1508,N_1560);
and U1612 (N_1612,N_1522,N_1551);
nand U1613 (N_1613,N_1529,N_1525);
nand U1614 (N_1614,N_1525,N_1519);
nand U1615 (N_1615,N_1573,N_1568);
nand U1616 (N_1616,N_1500,N_1544);
nand U1617 (N_1617,N_1539,N_1545);
nand U1618 (N_1618,N_1501,N_1559);
and U1619 (N_1619,N_1536,N_1560);
nand U1620 (N_1620,N_1557,N_1572);
and U1621 (N_1621,N_1529,N_1528);
nor U1622 (N_1622,N_1535,N_1564);
nand U1623 (N_1623,N_1507,N_1519);
and U1624 (N_1624,N_1545,N_1522);
or U1625 (N_1625,N_1527,N_1541);
nor U1626 (N_1626,N_1501,N_1541);
or U1627 (N_1627,N_1560,N_1512);
nor U1628 (N_1628,N_1558,N_1501);
nor U1629 (N_1629,N_1512,N_1518);
or U1630 (N_1630,N_1515,N_1560);
and U1631 (N_1631,N_1535,N_1500);
and U1632 (N_1632,N_1509,N_1567);
xor U1633 (N_1633,N_1530,N_1541);
nor U1634 (N_1634,N_1512,N_1563);
or U1635 (N_1635,N_1562,N_1519);
nand U1636 (N_1636,N_1518,N_1571);
or U1637 (N_1637,N_1538,N_1553);
and U1638 (N_1638,N_1568,N_1508);
or U1639 (N_1639,N_1546,N_1515);
or U1640 (N_1640,N_1536,N_1566);
nand U1641 (N_1641,N_1508,N_1524);
nand U1642 (N_1642,N_1514,N_1572);
nand U1643 (N_1643,N_1524,N_1569);
xor U1644 (N_1644,N_1523,N_1535);
nand U1645 (N_1645,N_1515,N_1547);
and U1646 (N_1646,N_1538,N_1529);
nor U1647 (N_1647,N_1568,N_1566);
and U1648 (N_1648,N_1571,N_1546);
or U1649 (N_1649,N_1510,N_1539);
nand U1650 (N_1650,N_1602,N_1639);
or U1651 (N_1651,N_1630,N_1588);
and U1652 (N_1652,N_1585,N_1577);
and U1653 (N_1653,N_1619,N_1648);
xor U1654 (N_1654,N_1611,N_1628);
xor U1655 (N_1655,N_1641,N_1626);
or U1656 (N_1656,N_1597,N_1589);
nor U1657 (N_1657,N_1627,N_1649);
xor U1658 (N_1658,N_1580,N_1631);
and U1659 (N_1659,N_1593,N_1613);
nor U1660 (N_1660,N_1578,N_1612);
nor U1661 (N_1661,N_1618,N_1615);
or U1662 (N_1662,N_1645,N_1587);
nor U1663 (N_1663,N_1616,N_1586);
nand U1664 (N_1664,N_1591,N_1596);
nor U1665 (N_1665,N_1579,N_1600);
or U1666 (N_1666,N_1621,N_1643);
nand U1667 (N_1667,N_1620,N_1617);
xnor U1668 (N_1668,N_1601,N_1583);
and U1669 (N_1669,N_1635,N_1637);
or U1670 (N_1670,N_1575,N_1609);
xor U1671 (N_1671,N_1576,N_1605);
or U1672 (N_1672,N_1642,N_1623);
nor U1673 (N_1673,N_1634,N_1644);
nand U1674 (N_1674,N_1598,N_1622);
xnor U1675 (N_1675,N_1603,N_1582);
nand U1676 (N_1676,N_1607,N_1638);
nor U1677 (N_1677,N_1633,N_1590);
xnor U1678 (N_1678,N_1624,N_1610);
or U1679 (N_1679,N_1646,N_1604);
nand U1680 (N_1680,N_1636,N_1632);
or U1681 (N_1681,N_1614,N_1594);
xor U1682 (N_1682,N_1647,N_1595);
nand U1683 (N_1683,N_1592,N_1608);
nand U1684 (N_1684,N_1629,N_1584);
nor U1685 (N_1685,N_1640,N_1599);
or U1686 (N_1686,N_1606,N_1581);
nand U1687 (N_1687,N_1625,N_1606);
nor U1688 (N_1688,N_1587,N_1638);
nor U1689 (N_1689,N_1647,N_1589);
nor U1690 (N_1690,N_1636,N_1584);
or U1691 (N_1691,N_1641,N_1645);
nand U1692 (N_1692,N_1641,N_1630);
nor U1693 (N_1693,N_1636,N_1638);
and U1694 (N_1694,N_1619,N_1603);
nand U1695 (N_1695,N_1626,N_1631);
and U1696 (N_1696,N_1600,N_1640);
or U1697 (N_1697,N_1591,N_1635);
and U1698 (N_1698,N_1607,N_1582);
nor U1699 (N_1699,N_1641,N_1600);
or U1700 (N_1700,N_1642,N_1612);
and U1701 (N_1701,N_1649,N_1589);
nor U1702 (N_1702,N_1635,N_1584);
nand U1703 (N_1703,N_1606,N_1644);
xor U1704 (N_1704,N_1639,N_1587);
nand U1705 (N_1705,N_1608,N_1622);
nor U1706 (N_1706,N_1639,N_1624);
or U1707 (N_1707,N_1615,N_1644);
xnor U1708 (N_1708,N_1597,N_1630);
or U1709 (N_1709,N_1606,N_1594);
or U1710 (N_1710,N_1643,N_1629);
xor U1711 (N_1711,N_1641,N_1578);
xor U1712 (N_1712,N_1638,N_1576);
and U1713 (N_1713,N_1595,N_1592);
nor U1714 (N_1714,N_1576,N_1626);
nand U1715 (N_1715,N_1607,N_1631);
or U1716 (N_1716,N_1630,N_1635);
nor U1717 (N_1717,N_1591,N_1643);
or U1718 (N_1718,N_1589,N_1634);
or U1719 (N_1719,N_1578,N_1624);
nand U1720 (N_1720,N_1643,N_1619);
nor U1721 (N_1721,N_1601,N_1604);
nor U1722 (N_1722,N_1591,N_1587);
nand U1723 (N_1723,N_1596,N_1612);
nand U1724 (N_1724,N_1585,N_1619);
nand U1725 (N_1725,N_1658,N_1704);
nand U1726 (N_1726,N_1667,N_1701);
nor U1727 (N_1727,N_1664,N_1711);
nor U1728 (N_1728,N_1714,N_1713);
and U1729 (N_1729,N_1687,N_1696);
nor U1730 (N_1730,N_1655,N_1668);
or U1731 (N_1731,N_1659,N_1680);
or U1732 (N_1732,N_1705,N_1690);
nor U1733 (N_1733,N_1700,N_1672);
xor U1734 (N_1734,N_1721,N_1712);
nor U1735 (N_1735,N_1676,N_1698);
nand U1736 (N_1736,N_1710,N_1716);
or U1737 (N_1737,N_1675,N_1684);
nand U1738 (N_1738,N_1651,N_1720);
or U1739 (N_1739,N_1656,N_1715);
and U1740 (N_1740,N_1708,N_1654);
and U1741 (N_1741,N_1691,N_1685);
nand U1742 (N_1742,N_1723,N_1673);
nand U1743 (N_1743,N_1652,N_1666);
xnor U1744 (N_1744,N_1661,N_1693);
nand U1745 (N_1745,N_1699,N_1695);
or U1746 (N_1746,N_1707,N_1670);
and U1747 (N_1747,N_1702,N_1683);
or U1748 (N_1748,N_1657,N_1706);
or U1749 (N_1749,N_1686,N_1679);
and U1750 (N_1750,N_1719,N_1703);
nor U1751 (N_1751,N_1671,N_1660);
nand U1752 (N_1752,N_1718,N_1709);
nor U1753 (N_1753,N_1669,N_1688);
nand U1754 (N_1754,N_1674,N_1697);
and U1755 (N_1755,N_1678,N_1682);
or U1756 (N_1756,N_1677,N_1724);
and U1757 (N_1757,N_1681,N_1663);
and U1758 (N_1758,N_1653,N_1665);
nand U1759 (N_1759,N_1662,N_1692);
nor U1760 (N_1760,N_1722,N_1650);
xor U1761 (N_1761,N_1694,N_1717);
or U1762 (N_1762,N_1689,N_1673);
xor U1763 (N_1763,N_1690,N_1719);
or U1764 (N_1764,N_1711,N_1656);
nor U1765 (N_1765,N_1703,N_1674);
or U1766 (N_1766,N_1715,N_1665);
and U1767 (N_1767,N_1669,N_1662);
and U1768 (N_1768,N_1682,N_1694);
or U1769 (N_1769,N_1656,N_1654);
and U1770 (N_1770,N_1657,N_1653);
and U1771 (N_1771,N_1719,N_1701);
or U1772 (N_1772,N_1722,N_1716);
or U1773 (N_1773,N_1661,N_1695);
nand U1774 (N_1774,N_1714,N_1691);
or U1775 (N_1775,N_1720,N_1717);
xor U1776 (N_1776,N_1711,N_1678);
nor U1777 (N_1777,N_1694,N_1654);
nor U1778 (N_1778,N_1670,N_1700);
or U1779 (N_1779,N_1650,N_1721);
nand U1780 (N_1780,N_1714,N_1696);
and U1781 (N_1781,N_1695,N_1658);
or U1782 (N_1782,N_1685,N_1703);
xor U1783 (N_1783,N_1704,N_1698);
or U1784 (N_1784,N_1698,N_1653);
nor U1785 (N_1785,N_1658,N_1670);
and U1786 (N_1786,N_1698,N_1718);
xnor U1787 (N_1787,N_1685,N_1669);
xnor U1788 (N_1788,N_1682,N_1674);
and U1789 (N_1789,N_1673,N_1663);
nand U1790 (N_1790,N_1658,N_1676);
nor U1791 (N_1791,N_1709,N_1695);
nand U1792 (N_1792,N_1675,N_1674);
nor U1793 (N_1793,N_1721,N_1696);
nand U1794 (N_1794,N_1691,N_1724);
nor U1795 (N_1795,N_1717,N_1659);
nand U1796 (N_1796,N_1695,N_1712);
and U1797 (N_1797,N_1670,N_1715);
xor U1798 (N_1798,N_1681,N_1654);
nor U1799 (N_1799,N_1692,N_1721);
nor U1800 (N_1800,N_1782,N_1728);
nand U1801 (N_1801,N_1738,N_1764);
xor U1802 (N_1802,N_1795,N_1791);
and U1803 (N_1803,N_1757,N_1758);
nand U1804 (N_1804,N_1792,N_1775);
nor U1805 (N_1805,N_1781,N_1742);
and U1806 (N_1806,N_1763,N_1780);
nand U1807 (N_1807,N_1765,N_1730);
nand U1808 (N_1808,N_1743,N_1770);
or U1809 (N_1809,N_1799,N_1762);
and U1810 (N_1810,N_1741,N_1760);
xor U1811 (N_1811,N_1725,N_1747);
nand U1812 (N_1812,N_1727,N_1783);
nor U1813 (N_1813,N_1787,N_1731);
and U1814 (N_1814,N_1754,N_1766);
xnor U1815 (N_1815,N_1755,N_1746);
nor U1816 (N_1816,N_1773,N_1793);
nand U1817 (N_1817,N_1786,N_1744);
or U1818 (N_1818,N_1756,N_1789);
nor U1819 (N_1819,N_1798,N_1751);
or U1820 (N_1820,N_1733,N_1736);
nand U1821 (N_1821,N_1752,N_1790);
nor U1822 (N_1822,N_1767,N_1772);
and U1823 (N_1823,N_1726,N_1774);
nand U1824 (N_1824,N_1768,N_1784);
nand U1825 (N_1825,N_1776,N_1748);
and U1826 (N_1826,N_1732,N_1749);
nand U1827 (N_1827,N_1769,N_1737);
nor U1828 (N_1828,N_1761,N_1777);
and U1829 (N_1829,N_1759,N_1735);
nor U1830 (N_1830,N_1779,N_1750);
and U1831 (N_1831,N_1788,N_1778);
and U1832 (N_1832,N_1729,N_1796);
and U1833 (N_1833,N_1734,N_1771);
nor U1834 (N_1834,N_1740,N_1739);
and U1835 (N_1835,N_1753,N_1785);
or U1836 (N_1836,N_1794,N_1797);
xnor U1837 (N_1837,N_1745,N_1764);
or U1838 (N_1838,N_1774,N_1788);
nand U1839 (N_1839,N_1777,N_1732);
nor U1840 (N_1840,N_1752,N_1798);
and U1841 (N_1841,N_1750,N_1737);
and U1842 (N_1842,N_1744,N_1729);
xor U1843 (N_1843,N_1767,N_1787);
nor U1844 (N_1844,N_1799,N_1790);
or U1845 (N_1845,N_1798,N_1777);
nand U1846 (N_1846,N_1764,N_1749);
and U1847 (N_1847,N_1754,N_1780);
nor U1848 (N_1848,N_1781,N_1728);
or U1849 (N_1849,N_1784,N_1747);
or U1850 (N_1850,N_1766,N_1760);
nand U1851 (N_1851,N_1768,N_1792);
nand U1852 (N_1852,N_1757,N_1766);
or U1853 (N_1853,N_1757,N_1782);
and U1854 (N_1854,N_1739,N_1795);
and U1855 (N_1855,N_1796,N_1756);
nand U1856 (N_1856,N_1757,N_1753);
nor U1857 (N_1857,N_1745,N_1767);
nor U1858 (N_1858,N_1775,N_1737);
or U1859 (N_1859,N_1798,N_1731);
or U1860 (N_1860,N_1749,N_1793);
nand U1861 (N_1861,N_1759,N_1789);
and U1862 (N_1862,N_1769,N_1733);
nor U1863 (N_1863,N_1773,N_1731);
nand U1864 (N_1864,N_1753,N_1739);
or U1865 (N_1865,N_1758,N_1767);
and U1866 (N_1866,N_1785,N_1740);
xor U1867 (N_1867,N_1740,N_1779);
nand U1868 (N_1868,N_1791,N_1726);
xor U1869 (N_1869,N_1774,N_1736);
nor U1870 (N_1870,N_1761,N_1731);
or U1871 (N_1871,N_1741,N_1790);
nor U1872 (N_1872,N_1737,N_1735);
nor U1873 (N_1873,N_1760,N_1739);
nand U1874 (N_1874,N_1755,N_1794);
or U1875 (N_1875,N_1874,N_1855);
nor U1876 (N_1876,N_1802,N_1838);
nand U1877 (N_1877,N_1810,N_1800);
nand U1878 (N_1878,N_1832,N_1865);
nand U1879 (N_1879,N_1830,N_1822);
nand U1880 (N_1880,N_1866,N_1853);
nor U1881 (N_1881,N_1867,N_1816);
xnor U1882 (N_1882,N_1854,N_1837);
or U1883 (N_1883,N_1847,N_1873);
nand U1884 (N_1884,N_1851,N_1823);
nor U1885 (N_1885,N_1860,N_1859);
nand U1886 (N_1886,N_1808,N_1850);
and U1887 (N_1887,N_1818,N_1840);
nor U1888 (N_1888,N_1813,N_1829);
xnor U1889 (N_1889,N_1841,N_1868);
nor U1890 (N_1890,N_1805,N_1870);
or U1891 (N_1891,N_1819,N_1836);
nor U1892 (N_1892,N_1825,N_1869);
xor U1893 (N_1893,N_1844,N_1839);
or U1894 (N_1894,N_1801,N_1871);
nor U1895 (N_1895,N_1803,N_1809);
and U1896 (N_1896,N_1852,N_1804);
nand U1897 (N_1897,N_1814,N_1846);
xor U1898 (N_1898,N_1831,N_1833);
xor U1899 (N_1899,N_1812,N_1817);
nand U1900 (N_1900,N_1862,N_1828);
nand U1901 (N_1901,N_1856,N_1827);
and U1902 (N_1902,N_1834,N_1857);
and U1903 (N_1903,N_1826,N_1842);
nand U1904 (N_1904,N_1849,N_1820);
nor U1905 (N_1905,N_1843,N_1872);
nor U1906 (N_1906,N_1845,N_1824);
nor U1907 (N_1907,N_1835,N_1821);
and U1908 (N_1908,N_1811,N_1807);
nor U1909 (N_1909,N_1848,N_1864);
and U1910 (N_1910,N_1858,N_1863);
nor U1911 (N_1911,N_1806,N_1815);
xor U1912 (N_1912,N_1861,N_1817);
and U1913 (N_1913,N_1844,N_1815);
xor U1914 (N_1914,N_1863,N_1803);
or U1915 (N_1915,N_1847,N_1854);
nor U1916 (N_1916,N_1858,N_1871);
xor U1917 (N_1917,N_1812,N_1824);
and U1918 (N_1918,N_1850,N_1873);
nand U1919 (N_1919,N_1838,N_1814);
or U1920 (N_1920,N_1827,N_1857);
or U1921 (N_1921,N_1823,N_1807);
and U1922 (N_1922,N_1860,N_1841);
nor U1923 (N_1923,N_1843,N_1828);
or U1924 (N_1924,N_1839,N_1825);
nand U1925 (N_1925,N_1830,N_1858);
or U1926 (N_1926,N_1858,N_1821);
and U1927 (N_1927,N_1836,N_1809);
or U1928 (N_1928,N_1856,N_1846);
and U1929 (N_1929,N_1807,N_1861);
or U1930 (N_1930,N_1808,N_1815);
or U1931 (N_1931,N_1843,N_1864);
nor U1932 (N_1932,N_1835,N_1833);
and U1933 (N_1933,N_1834,N_1845);
nand U1934 (N_1934,N_1845,N_1833);
nor U1935 (N_1935,N_1838,N_1861);
and U1936 (N_1936,N_1838,N_1856);
nor U1937 (N_1937,N_1805,N_1836);
nand U1938 (N_1938,N_1829,N_1846);
nand U1939 (N_1939,N_1804,N_1813);
nand U1940 (N_1940,N_1872,N_1856);
or U1941 (N_1941,N_1842,N_1851);
nand U1942 (N_1942,N_1823,N_1811);
or U1943 (N_1943,N_1801,N_1851);
nand U1944 (N_1944,N_1809,N_1858);
nand U1945 (N_1945,N_1840,N_1810);
nor U1946 (N_1946,N_1873,N_1803);
or U1947 (N_1947,N_1871,N_1837);
nand U1948 (N_1948,N_1829,N_1800);
xnor U1949 (N_1949,N_1851,N_1810);
or U1950 (N_1950,N_1930,N_1891);
nor U1951 (N_1951,N_1921,N_1943);
or U1952 (N_1952,N_1926,N_1878);
or U1953 (N_1953,N_1882,N_1918);
or U1954 (N_1954,N_1933,N_1929);
or U1955 (N_1955,N_1913,N_1911);
or U1956 (N_1956,N_1935,N_1886);
or U1957 (N_1957,N_1914,N_1949);
or U1958 (N_1958,N_1934,N_1875);
nand U1959 (N_1959,N_1944,N_1895);
nor U1960 (N_1960,N_1924,N_1917);
or U1961 (N_1961,N_1912,N_1940);
xor U1962 (N_1962,N_1900,N_1880);
nand U1963 (N_1963,N_1919,N_1899);
nand U1964 (N_1964,N_1881,N_1931);
xor U1965 (N_1965,N_1910,N_1908);
nand U1966 (N_1966,N_1920,N_1906);
or U1967 (N_1967,N_1927,N_1887);
nor U1968 (N_1968,N_1937,N_1894);
nand U1969 (N_1969,N_1907,N_1945);
or U1970 (N_1970,N_1902,N_1936);
or U1971 (N_1971,N_1890,N_1883);
nand U1972 (N_1972,N_1905,N_1901);
and U1973 (N_1973,N_1939,N_1904);
nand U1974 (N_1974,N_1879,N_1885);
nor U1975 (N_1975,N_1892,N_1946);
nand U1976 (N_1976,N_1889,N_1893);
and U1977 (N_1977,N_1888,N_1876);
or U1978 (N_1978,N_1942,N_1916);
nand U1979 (N_1979,N_1877,N_1923);
and U1980 (N_1980,N_1941,N_1897);
and U1981 (N_1981,N_1898,N_1948);
nor U1982 (N_1982,N_1903,N_1915);
or U1983 (N_1983,N_1928,N_1925);
and U1984 (N_1984,N_1884,N_1938);
nor U1985 (N_1985,N_1932,N_1909);
nor U1986 (N_1986,N_1922,N_1896);
xor U1987 (N_1987,N_1947,N_1906);
and U1988 (N_1988,N_1901,N_1892);
nor U1989 (N_1989,N_1919,N_1947);
nand U1990 (N_1990,N_1913,N_1914);
nand U1991 (N_1991,N_1903,N_1875);
or U1992 (N_1992,N_1884,N_1913);
nand U1993 (N_1993,N_1900,N_1899);
nand U1994 (N_1994,N_1932,N_1940);
nand U1995 (N_1995,N_1889,N_1899);
or U1996 (N_1996,N_1893,N_1898);
nor U1997 (N_1997,N_1934,N_1930);
nor U1998 (N_1998,N_1910,N_1930);
or U1999 (N_1999,N_1926,N_1912);
nor U2000 (N_2000,N_1935,N_1921);
nand U2001 (N_2001,N_1914,N_1878);
and U2002 (N_2002,N_1898,N_1946);
or U2003 (N_2003,N_1892,N_1879);
or U2004 (N_2004,N_1910,N_1920);
nor U2005 (N_2005,N_1939,N_1940);
nor U2006 (N_2006,N_1882,N_1885);
and U2007 (N_2007,N_1917,N_1949);
and U2008 (N_2008,N_1900,N_1929);
and U2009 (N_2009,N_1877,N_1895);
and U2010 (N_2010,N_1939,N_1945);
or U2011 (N_2011,N_1921,N_1923);
nor U2012 (N_2012,N_1904,N_1941);
nand U2013 (N_2013,N_1936,N_1898);
nand U2014 (N_2014,N_1889,N_1940);
nand U2015 (N_2015,N_1941,N_1896);
nand U2016 (N_2016,N_1875,N_1910);
and U2017 (N_2017,N_1925,N_1892);
nand U2018 (N_2018,N_1947,N_1914);
and U2019 (N_2019,N_1941,N_1932);
nand U2020 (N_2020,N_1942,N_1930);
or U2021 (N_2021,N_1943,N_1935);
nor U2022 (N_2022,N_1890,N_1911);
and U2023 (N_2023,N_1929,N_1943);
and U2024 (N_2024,N_1889,N_1904);
or U2025 (N_2025,N_1960,N_1968);
and U2026 (N_2026,N_1994,N_2024);
nor U2027 (N_2027,N_2010,N_1979);
or U2028 (N_2028,N_1971,N_1954);
nand U2029 (N_2029,N_1967,N_1980);
nor U2030 (N_2030,N_1953,N_2019);
nor U2031 (N_2031,N_1981,N_1950);
nand U2032 (N_2032,N_1990,N_1999);
or U2033 (N_2033,N_1996,N_1987);
nor U2034 (N_2034,N_2016,N_1985);
and U2035 (N_2035,N_2023,N_2020);
nor U2036 (N_2036,N_1992,N_1951);
and U2037 (N_2037,N_1997,N_1958);
nand U2038 (N_2038,N_1991,N_2012);
or U2039 (N_2039,N_1955,N_1964);
nor U2040 (N_2040,N_1982,N_1976);
and U2041 (N_2041,N_1977,N_2018);
xnor U2042 (N_2042,N_1973,N_1956);
or U2043 (N_2043,N_2000,N_1963);
or U2044 (N_2044,N_1965,N_1998);
or U2045 (N_2045,N_2017,N_1975);
nand U2046 (N_2046,N_1993,N_2005);
nand U2047 (N_2047,N_2011,N_1970);
or U2048 (N_2048,N_2021,N_1961);
nor U2049 (N_2049,N_1952,N_2008);
or U2050 (N_2050,N_1962,N_2001);
nor U2051 (N_2051,N_1966,N_2014);
nand U2052 (N_2052,N_1957,N_2022);
and U2053 (N_2053,N_1974,N_1986);
and U2054 (N_2054,N_1959,N_2013);
or U2055 (N_2055,N_2009,N_2003);
or U2056 (N_2056,N_1978,N_1969);
nand U2057 (N_2057,N_2006,N_2015);
and U2058 (N_2058,N_1989,N_2004);
or U2059 (N_2059,N_1995,N_2002);
and U2060 (N_2060,N_1983,N_1972);
and U2061 (N_2061,N_2007,N_1988);
xor U2062 (N_2062,N_1984,N_1976);
nand U2063 (N_2063,N_2010,N_2002);
and U2064 (N_2064,N_1989,N_1983);
xor U2065 (N_2065,N_2023,N_1984);
nor U2066 (N_2066,N_2019,N_1993);
or U2067 (N_2067,N_2003,N_1988);
and U2068 (N_2068,N_2009,N_2024);
nand U2069 (N_2069,N_1962,N_1982);
or U2070 (N_2070,N_1965,N_2021);
nor U2071 (N_2071,N_1963,N_2006);
xnor U2072 (N_2072,N_2016,N_2015);
and U2073 (N_2073,N_1975,N_1978);
nor U2074 (N_2074,N_2004,N_1972);
and U2075 (N_2075,N_2018,N_1965);
and U2076 (N_2076,N_2018,N_1979);
nand U2077 (N_2077,N_2003,N_2004);
and U2078 (N_2078,N_2012,N_1963);
or U2079 (N_2079,N_1966,N_1970);
nor U2080 (N_2080,N_1951,N_2011);
and U2081 (N_2081,N_1971,N_1979);
or U2082 (N_2082,N_2017,N_1966);
nor U2083 (N_2083,N_1976,N_2013);
nor U2084 (N_2084,N_2016,N_1997);
nor U2085 (N_2085,N_1972,N_1985);
and U2086 (N_2086,N_2003,N_1978);
or U2087 (N_2087,N_2017,N_1973);
nor U2088 (N_2088,N_1997,N_1999);
nor U2089 (N_2089,N_2017,N_1984);
xnor U2090 (N_2090,N_2016,N_1955);
nand U2091 (N_2091,N_1963,N_1977);
or U2092 (N_2092,N_1999,N_2007);
nor U2093 (N_2093,N_1954,N_2018);
and U2094 (N_2094,N_1978,N_2019);
and U2095 (N_2095,N_2022,N_1996);
nor U2096 (N_2096,N_1958,N_1969);
nand U2097 (N_2097,N_1953,N_2013);
and U2098 (N_2098,N_1951,N_1980);
nor U2099 (N_2099,N_1998,N_2021);
or U2100 (N_2100,N_2037,N_2090);
nand U2101 (N_2101,N_2043,N_2066);
nand U2102 (N_2102,N_2064,N_2088);
or U2103 (N_2103,N_2029,N_2082);
nor U2104 (N_2104,N_2034,N_2027);
xor U2105 (N_2105,N_2050,N_2093);
xnor U2106 (N_2106,N_2047,N_2026);
or U2107 (N_2107,N_2058,N_2033);
xor U2108 (N_2108,N_2056,N_2076);
and U2109 (N_2109,N_2089,N_2036);
and U2110 (N_2110,N_2052,N_2067);
or U2111 (N_2111,N_2060,N_2038);
nor U2112 (N_2112,N_2040,N_2091);
nand U2113 (N_2113,N_2053,N_2079);
nand U2114 (N_2114,N_2055,N_2080);
nor U2115 (N_2115,N_2045,N_2030);
and U2116 (N_2116,N_2084,N_2046);
and U2117 (N_2117,N_2097,N_2041);
nor U2118 (N_2118,N_2072,N_2096);
or U2119 (N_2119,N_2081,N_2070);
nand U2120 (N_2120,N_2094,N_2085);
nand U2121 (N_2121,N_2075,N_2025);
or U2122 (N_2122,N_2042,N_2032);
and U2123 (N_2123,N_2065,N_2054);
and U2124 (N_2124,N_2031,N_2069);
nand U2125 (N_2125,N_2083,N_2057);
and U2126 (N_2126,N_2044,N_2078);
and U2127 (N_2127,N_2098,N_2077);
or U2128 (N_2128,N_2087,N_2059);
nor U2129 (N_2129,N_2074,N_2073);
nor U2130 (N_2130,N_2063,N_2068);
nor U2131 (N_2131,N_2061,N_2095);
xor U2132 (N_2132,N_2039,N_2062);
nand U2133 (N_2133,N_2049,N_2086);
nand U2134 (N_2134,N_2051,N_2035);
and U2135 (N_2135,N_2048,N_2099);
or U2136 (N_2136,N_2071,N_2028);
nor U2137 (N_2137,N_2092,N_2055);
and U2138 (N_2138,N_2033,N_2088);
nor U2139 (N_2139,N_2054,N_2074);
and U2140 (N_2140,N_2027,N_2081);
and U2141 (N_2141,N_2092,N_2029);
nand U2142 (N_2142,N_2037,N_2066);
nor U2143 (N_2143,N_2083,N_2072);
and U2144 (N_2144,N_2071,N_2035);
or U2145 (N_2145,N_2049,N_2062);
or U2146 (N_2146,N_2055,N_2096);
nand U2147 (N_2147,N_2077,N_2027);
or U2148 (N_2148,N_2096,N_2086);
nor U2149 (N_2149,N_2039,N_2049);
and U2150 (N_2150,N_2066,N_2048);
nor U2151 (N_2151,N_2034,N_2099);
nor U2152 (N_2152,N_2025,N_2052);
and U2153 (N_2153,N_2063,N_2053);
xor U2154 (N_2154,N_2067,N_2090);
nand U2155 (N_2155,N_2046,N_2073);
nor U2156 (N_2156,N_2051,N_2048);
nor U2157 (N_2157,N_2030,N_2034);
xor U2158 (N_2158,N_2027,N_2060);
or U2159 (N_2159,N_2030,N_2031);
xor U2160 (N_2160,N_2061,N_2052);
and U2161 (N_2161,N_2051,N_2053);
nor U2162 (N_2162,N_2058,N_2051);
nand U2163 (N_2163,N_2042,N_2068);
nor U2164 (N_2164,N_2042,N_2093);
nor U2165 (N_2165,N_2067,N_2098);
xnor U2166 (N_2166,N_2094,N_2099);
or U2167 (N_2167,N_2060,N_2094);
xor U2168 (N_2168,N_2035,N_2076);
or U2169 (N_2169,N_2047,N_2069);
nand U2170 (N_2170,N_2075,N_2093);
nor U2171 (N_2171,N_2062,N_2052);
nor U2172 (N_2172,N_2068,N_2080);
xnor U2173 (N_2173,N_2071,N_2065);
and U2174 (N_2174,N_2082,N_2026);
and U2175 (N_2175,N_2108,N_2156);
or U2176 (N_2176,N_2155,N_2101);
nor U2177 (N_2177,N_2147,N_2121);
or U2178 (N_2178,N_2161,N_2170);
xor U2179 (N_2179,N_2174,N_2141);
and U2180 (N_2180,N_2102,N_2111);
or U2181 (N_2181,N_2106,N_2136);
and U2182 (N_2182,N_2139,N_2138);
xnor U2183 (N_2183,N_2112,N_2152);
nor U2184 (N_2184,N_2127,N_2162);
nor U2185 (N_2185,N_2126,N_2103);
nor U2186 (N_2186,N_2142,N_2144);
or U2187 (N_2187,N_2135,N_2157);
and U2188 (N_2188,N_2129,N_2173);
nand U2189 (N_2189,N_2110,N_2105);
xor U2190 (N_2190,N_2154,N_2107);
xor U2191 (N_2191,N_2163,N_2150);
and U2192 (N_2192,N_2125,N_2172);
nand U2193 (N_2193,N_2109,N_2122);
nor U2194 (N_2194,N_2143,N_2160);
nor U2195 (N_2195,N_2146,N_2158);
nand U2196 (N_2196,N_2114,N_2140);
nor U2197 (N_2197,N_2131,N_2171);
xor U2198 (N_2198,N_2132,N_2149);
or U2199 (N_2199,N_2159,N_2119);
nand U2200 (N_2200,N_2134,N_2133);
or U2201 (N_2201,N_2165,N_2120);
nor U2202 (N_2202,N_2153,N_2166);
nor U2203 (N_2203,N_2130,N_2123);
nand U2204 (N_2204,N_2118,N_2117);
or U2205 (N_2205,N_2100,N_2169);
nand U2206 (N_2206,N_2116,N_2137);
xnor U2207 (N_2207,N_2115,N_2151);
nand U2208 (N_2208,N_2128,N_2104);
or U2209 (N_2209,N_2148,N_2168);
or U2210 (N_2210,N_2145,N_2164);
nand U2211 (N_2211,N_2113,N_2167);
and U2212 (N_2212,N_2124,N_2132);
nor U2213 (N_2213,N_2108,N_2122);
nand U2214 (N_2214,N_2129,N_2126);
xor U2215 (N_2215,N_2142,N_2147);
and U2216 (N_2216,N_2103,N_2136);
and U2217 (N_2217,N_2145,N_2133);
and U2218 (N_2218,N_2106,N_2107);
or U2219 (N_2219,N_2149,N_2173);
or U2220 (N_2220,N_2172,N_2104);
and U2221 (N_2221,N_2106,N_2101);
nand U2222 (N_2222,N_2142,N_2103);
nand U2223 (N_2223,N_2115,N_2156);
nand U2224 (N_2224,N_2117,N_2151);
or U2225 (N_2225,N_2152,N_2163);
nand U2226 (N_2226,N_2134,N_2116);
and U2227 (N_2227,N_2135,N_2158);
nand U2228 (N_2228,N_2120,N_2140);
and U2229 (N_2229,N_2161,N_2134);
or U2230 (N_2230,N_2165,N_2132);
nand U2231 (N_2231,N_2127,N_2156);
nor U2232 (N_2232,N_2118,N_2150);
nor U2233 (N_2233,N_2163,N_2139);
xnor U2234 (N_2234,N_2135,N_2105);
nor U2235 (N_2235,N_2137,N_2105);
nor U2236 (N_2236,N_2154,N_2135);
or U2237 (N_2237,N_2143,N_2112);
nor U2238 (N_2238,N_2125,N_2121);
nand U2239 (N_2239,N_2149,N_2161);
or U2240 (N_2240,N_2156,N_2104);
nor U2241 (N_2241,N_2156,N_2129);
and U2242 (N_2242,N_2162,N_2123);
or U2243 (N_2243,N_2164,N_2154);
nor U2244 (N_2244,N_2103,N_2132);
nor U2245 (N_2245,N_2150,N_2141);
and U2246 (N_2246,N_2140,N_2103);
nor U2247 (N_2247,N_2158,N_2104);
and U2248 (N_2248,N_2147,N_2119);
nand U2249 (N_2249,N_2149,N_2118);
xnor U2250 (N_2250,N_2183,N_2190);
or U2251 (N_2251,N_2245,N_2186);
or U2252 (N_2252,N_2225,N_2232);
nor U2253 (N_2253,N_2210,N_2185);
nor U2254 (N_2254,N_2182,N_2218);
nand U2255 (N_2255,N_2196,N_2179);
nand U2256 (N_2256,N_2181,N_2220);
nor U2257 (N_2257,N_2200,N_2243);
or U2258 (N_2258,N_2201,N_2208);
nor U2259 (N_2259,N_2189,N_2211);
nor U2260 (N_2260,N_2244,N_2228);
or U2261 (N_2261,N_2176,N_2202);
or U2262 (N_2262,N_2205,N_2177);
or U2263 (N_2263,N_2235,N_2199);
nand U2264 (N_2264,N_2242,N_2236);
or U2265 (N_2265,N_2229,N_2194);
or U2266 (N_2266,N_2207,N_2233);
nor U2267 (N_2267,N_2240,N_2215);
or U2268 (N_2268,N_2191,N_2184);
nor U2269 (N_2269,N_2192,N_2213);
nand U2270 (N_2270,N_2221,N_2188);
nand U2271 (N_2271,N_2231,N_2249);
nand U2272 (N_2272,N_2195,N_2238);
or U2273 (N_2273,N_2178,N_2217);
or U2274 (N_2274,N_2247,N_2237);
and U2275 (N_2275,N_2204,N_2175);
and U2276 (N_2276,N_2234,N_2219);
and U2277 (N_2277,N_2241,N_2187);
or U2278 (N_2278,N_2223,N_2206);
or U2279 (N_2279,N_2180,N_2227);
nand U2280 (N_2280,N_2198,N_2197);
and U2281 (N_2281,N_2209,N_2224);
or U2282 (N_2282,N_2246,N_2248);
or U2283 (N_2283,N_2193,N_2222);
and U2284 (N_2284,N_2212,N_2230);
nand U2285 (N_2285,N_2214,N_2203);
nor U2286 (N_2286,N_2239,N_2226);
or U2287 (N_2287,N_2216,N_2236);
nor U2288 (N_2288,N_2224,N_2240);
nand U2289 (N_2289,N_2211,N_2177);
nor U2290 (N_2290,N_2197,N_2227);
xnor U2291 (N_2291,N_2186,N_2226);
nor U2292 (N_2292,N_2225,N_2200);
xnor U2293 (N_2293,N_2233,N_2177);
xor U2294 (N_2294,N_2206,N_2212);
and U2295 (N_2295,N_2241,N_2216);
or U2296 (N_2296,N_2235,N_2232);
and U2297 (N_2297,N_2235,N_2238);
nor U2298 (N_2298,N_2241,N_2218);
nor U2299 (N_2299,N_2212,N_2198);
or U2300 (N_2300,N_2219,N_2205);
or U2301 (N_2301,N_2209,N_2242);
nand U2302 (N_2302,N_2189,N_2213);
xor U2303 (N_2303,N_2247,N_2205);
and U2304 (N_2304,N_2184,N_2220);
or U2305 (N_2305,N_2216,N_2248);
and U2306 (N_2306,N_2249,N_2215);
nor U2307 (N_2307,N_2189,N_2203);
or U2308 (N_2308,N_2185,N_2198);
and U2309 (N_2309,N_2193,N_2178);
or U2310 (N_2310,N_2197,N_2230);
nor U2311 (N_2311,N_2198,N_2242);
and U2312 (N_2312,N_2194,N_2186);
nor U2313 (N_2313,N_2227,N_2218);
or U2314 (N_2314,N_2205,N_2195);
nor U2315 (N_2315,N_2186,N_2234);
or U2316 (N_2316,N_2209,N_2190);
and U2317 (N_2317,N_2192,N_2210);
nor U2318 (N_2318,N_2199,N_2219);
and U2319 (N_2319,N_2204,N_2218);
or U2320 (N_2320,N_2220,N_2208);
or U2321 (N_2321,N_2184,N_2188);
and U2322 (N_2322,N_2195,N_2211);
nor U2323 (N_2323,N_2209,N_2192);
and U2324 (N_2324,N_2249,N_2223);
and U2325 (N_2325,N_2287,N_2262);
nand U2326 (N_2326,N_2264,N_2304);
nor U2327 (N_2327,N_2282,N_2316);
xnor U2328 (N_2328,N_2277,N_2305);
and U2329 (N_2329,N_2271,N_2279);
nor U2330 (N_2330,N_2286,N_2270);
and U2331 (N_2331,N_2315,N_2299);
nand U2332 (N_2332,N_2256,N_2312);
nor U2333 (N_2333,N_2284,N_2250);
nor U2334 (N_2334,N_2319,N_2311);
nor U2335 (N_2335,N_2281,N_2322);
xor U2336 (N_2336,N_2320,N_2296);
or U2337 (N_2337,N_2295,N_2290);
and U2338 (N_2338,N_2273,N_2318);
or U2339 (N_2339,N_2269,N_2275);
nand U2340 (N_2340,N_2258,N_2260);
nand U2341 (N_2341,N_2255,N_2272);
nor U2342 (N_2342,N_2268,N_2298);
nor U2343 (N_2343,N_2288,N_2261);
nand U2344 (N_2344,N_2292,N_2297);
nor U2345 (N_2345,N_2291,N_2263);
and U2346 (N_2346,N_2254,N_2265);
or U2347 (N_2347,N_2302,N_2293);
nand U2348 (N_2348,N_2259,N_2323);
nor U2349 (N_2349,N_2257,N_2267);
xor U2350 (N_2350,N_2294,N_2314);
and U2351 (N_2351,N_2274,N_2283);
or U2352 (N_2352,N_2313,N_2276);
nand U2353 (N_2353,N_2285,N_2251);
nand U2354 (N_2354,N_2321,N_2306);
nand U2355 (N_2355,N_2317,N_2253);
and U2356 (N_2356,N_2301,N_2300);
or U2357 (N_2357,N_2309,N_2303);
or U2358 (N_2358,N_2289,N_2266);
nor U2359 (N_2359,N_2310,N_2280);
nand U2360 (N_2360,N_2308,N_2278);
and U2361 (N_2361,N_2252,N_2324);
or U2362 (N_2362,N_2307,N_2298);
and U2363 (N_2363,N_2275,N_2314);
xnor U2364 (N_2364,N_2291,N_2312);
or U2365 (N_2365,N_2276,N_2272);
nand U2366 (N_2366,N_2301,N_2322);
and U2367 (N_2367,N_2321,N_2278);
or U2368 (N_2368,N_2279,N_2286);
xor U2369 (N_2369,N_2321,N_2277);
nor U2370 (N_2370,N_2279,N_2319);
and U2371 (N_2371,N_2274,N_2298);
and U2372 (N_2372,N_2260,N_2324);
or U2373 (N_2373,N_2291,N_2273);
and U2374 (N_2374,N_2324,N_2322);
or U2375 (N_2375,N_2264,N_2287);
and U2376 (N_2376,N_2252,N_2286);
or U2377 (N_2377,N_2318,N_2258);
nor U2378 (N_2378,N_2324,N_2265);
nand U2379 (N_2379,N_2307,N_2286);
nor U2380 (N_2380,N_2319,N_2317);
nor U2381 (N_2381,N_2269,N_2291);
and U2382 (N_2382,N_2284,N_2306);
xnor U2383 (N_2383,N_2254,N_2298);
or U2384 (N_2384,N_2265,N_2309);
and U2385 (N_2385,N_2311,N_2253);
nand U2386 (N_2386,N_2317,N_2318);
nand U2387 (N_2387,N_2313,N_2318);
nand U2388 (N_2388,N_2307,N_2322);
nand U2389 (N_2389,N_2320,N_2252);
nor U2390 (N_2390,N_2275,N_2285);
nand U2391 (N_2391,N_2251,N_2253);
xor U2392 (N_2392,N_2284,N_2304);
xor U2393 (N_2393,N_2294,N_2272);
nor U2394 (N_2394,N_2278,N_2298);
or U2395 (N_2395,N_2303,N_2279);
and U2396 (N_2396,N_2302,N_2263);
nand U2397 (N_2397,N_2253,N_2292);
and U2398 (N_2398,N_2315,N_2311);
xor U2399 (N_2399,N_2269,N_2255);
xnor U2400 (N_2400,N_2341,N_2343);
nor U2401 (N_2401,N_2354,N_2383);
xor U2402 (N_2402,N_2349,N_2330);
nand U2403 (N_2403,N_2393,N_2334);
and U2404 (N_2404,N_2398,N_2328);
nor U2405 (N_2405,N_2346,N_2386);
nor U2406 (N_2406,N_2353,N_2381);
nand U2407 (N_2407,N_2384,N_2352);
nand U2408 (N_2408,N_2376,N_2377);
and U2409 (N_2409,N_2361,N_2332);
nor U2410 (N_2410,N_2366,N_2365);
or U2411 (N_2411,N_2333,N_2358);
nor U2412 (N_2412,N_2347,N_2378);
nor U2413 (N_2413,N_2337,N_2395);
nor U2414 (N_2414,N_2369,N_2382);
or U2415 (N_2415,N_2335,N_2355);
nand U2416 (N_2416,N_2331,N_2360);
nand U2417 (N_2417,N_2345,N_2371);
nor U2418 (N_2418,N_2364,N_2342);
and U2419 (N_2419,N_2326,N_2372);
and U2420 (N_2420,N_2368,N_2388);
xor U2421 (N_2421,N_2390,N_2374);
xor U2422 (N_2422,N_2380,N_2344);
and U2423 (N_2423,N_2336,N_2339);
nor U2424 (N_2424,N_2394,N_2325);
xnor U2425 (N_2425,N_2399,N_2389);
nand U2426 (N_2426,N_2385,N_2387);
or U2427 (N_2427,N_2391,N_2356);
xor U2428 (N_2428,N_2363,N_2367);
nor U2429 (N_2429,N_2340,N_2397);
or U2430 (N_2430,N_2329,N_2338);
and U2431 (N_2431,N_2348,N_2357);
or U2432 (N_2432,N_2351,N_2327);
nor U2433 (N_2433,N_2350,N_2359);
and U2434 (N_2434,N_2396,N_2373);
nand U2435 (N_2435,N_2379,N_2362);
xnor U2436 (N_2436,N_2370,N_2392);
or U2437 (N_2437,N_2375,N_2373);
nand U2438 (N_2438,N_2354,N_2331);
nor U2439 (N_2439,N_2393,N_2375);
nor U2440 (N_2440,N_2337,N_2364);
xor U2441 (N_2441,N_2365,N_2385);
or U2442 (N_2442,N_2353,N_2366);
nand U2443 (N_2443,N_2371,N_2368);
nand U2444 (N_2444,N_2373,N_2370);
nand U2445 (N_2445,N_2325,N_2395);
nand U2446 (N_2446,N_2332,N_2378);
nor U2447 (N_2447,N_2328,N_2365);
nor U2448 (N_2448,N_2384,N_2360);
or U2449 (N_2449,N_2396,N_2371);
and U2450 (N_2450,N_2382,N_2354);
or U2451 (N_2451,N_2361,N_2374);
nor U2452 (N_2452,N_2338,N_2363);
or U2453 (N_2453,N_2333,N_2361);
or U2454 (N_2454,N_2380,N_2326);
nor U2455 (N_2455,N_2384,N_2391);
nor U2456 (N_2456,N_2376,N_2367);
and U2457 (N_2457,N_2389,N_2374);
or U2458 (N_2458,N_2331,N_2329);
or U2459 (N_2459,N_2341,N_2340);
or U2460 (N_2460,N_2340,N_2339);
nor U2461 (N_2461,N_2339,N_2369);
or U2462 (N_2462,N_2382,N_2330);
nor U2463 (N_2463,N_2371,N_2387);
and U2464 (N_2464,N_2360,N_2332);
nor U2465 (N_2465,N_2348,N_2349);
xor U2466 (N_2466,N_2353,N_2359);
or U2467 (N_2467,N_2350,N_2395);
nor U2468 (N_2468,N_2346,N_2385);
or U2469 (N_2469,N_2391,N_2326);
nand U2470 (N_2470,N_2357,N_2386);
or U2471 (N_2471,N_2399,N_2338);
nor U2472 (N_2472,N_2397,N_2343);
and U2473 (N_2473,N_2378,N_2385);
nor U2474 (N_2474,N_2392,N_2396);
nand U2475 (N_2475,N_2400,N_2424);
or U2476 (N_2476,N_2418,N_2441);
and U2477 (N_2477,N_2430,N_2453);
and U2478 (N_2478,N_2433,N_2474);
nor U2479 (N_2479,N_2419,N_2442);
nand U2480 (N_2480,N_2455,N_2408);
nor U2481 (N_2481,N_2405,N_2473);
nor U2482 (N_2482,N_2440,N_2411);
nor U2483 (N_2483,N_2445,N_2409);
nand U2484 (N_2484,N_2471,N_2466);
or U2485 (N_2485,N_2464,N_2446);
xnor U2486 (N_2486,N_2416,N_2417);
nand U2487 (N_2487,N_2401,N_2429);
nand U2488 (N_2488,N_2447,N_2470);
nor U2489 (N_2489,N_2406,N_2467);
nand U2490 (N_2490,N_2459,N_2438);
and U2491 (N_2491,N_2461,N_2436);
xor U2492 (N_2492,N_2427,N_2437);
nand U2493 (N_2493,N_2444,N_2454);
nor U2494 (N_2494,N_2462,N_2413);
or U2495 (N_2495,N_2422,N_2402);
or U2496 (N_2496,N_2463,N_2449);
or U2497 (N_2497,N_2421,N_2410);
nand U2498 (N_2498,N_2423,N_2443);
and U2499 (N_2499,N_2472,N_2468);
nor U2500 (N_2500,N_2439,N_2426);
nor U2501 (N_2501,N_2414,N_2457);
and U2502 (N_2502,N_2460,N_2448);
or U2503 (N_2503,N_2403,N_2415);
nor U2504 (N_2504,N_2432,N_2465);
or U2505 (N_2505,N_2452,N_2451);
nand U2506 (N_2506,N_2431,N_2450);
and U2507 (N_2507,N_2458,N_2407);
nor U2508 (N_2508,N_2456,N_2420);
and U2509 (N_2509,N_2428,N_2469);
nor U2510 (N_2510,N_2425,N_2435);
nand U2511 (N_2511,N_2412,N_2404);
and U2512 (N_2512,N_2434,N_2456);
or U2513 (N_2513,N_2473,N_2468);
nand U2514 (N_2514,N_2440,N_2435);
nor U2515 (N_2515,N_2421,N_2402);
or U2516 (N_2516,N_2423,N_2472);
nand U2517 (N_2517,N_2437,N_2419);
nor U2518 (N_2518,N_2448,N_2447);
and U2519 (N_2519,N_2440,N_2437);
and U2520 (N_2520,N_2437,N_2418);
nor U2521 (N_2521,N_2402,N_2466);
nor U2522 (N_2522,N_2403,N_2461);
and U2523 (N_2523,N_2440,N_2453);
xnor U2524 (N_2524,N_2457,N_2462);
xor U2525 (N_2525,N_2422,N_2468);
nor U2526 (N_2526,N_2433,N_2405);
nor U2527 (N_2527,N_2413,N_2405);
or U2528 (N_2528,N_2427,N_2436);
and U2529 (N_2529,N_2459,N_2458);
nor U2530 (N_2530,N_2402,N_2433);
nor U2531 (N_2531,N_2467,N_2418);
or U2532 (N_2532,N_2442,N_2405);
or U2533 (N_2533,N_2426,N_2435);
and U2534 (N_2534,N_2466,N_2413);
xor U2535 (N_2535,N_2445,N_2430);
nand U2536 (N_2536,N_2441,N_2462);
and U2537 (N_2537,N_2435,N_2433);
nand U2538 (N_2538,N_2453,N_2437);
or U2539 (N_2539,N_2418,N_2438);
nand U2540 (N_2540,N_2462,N_2437);
nand U2541 (N_2541,N_2474,N_2449);
or U2542 (N_2542,N_2421,N_2435);
or U2543 (N_2543,N_2427,N_2466);
and U2544 (N_2544,N_2443,N_2456);
nand U2545 (N_2545,N_2405,N_2412);
nand U2546 (N_2546,N_2466,N_2417);
nand U2547 (N_2547,N_2426,N_2445);
nand U2548 (N_2548,N_2425,N_2440);
nor U2549 (N_2549,N_2458,N_2420);
nor U2550 (N_2550,N_2509,N_2508);
xor U2551 (N_2551,N_2502,N_2503);
and U2552 (N_2552,N_2530,N_2486);
or U2553 (N_2553,N_2515,N_2525);
xnor U2554 (N_2554,N_2548,N_2538);
or U2555 (N_2555,N_2487,N_2543);
nand U2556 (N_2556,N_2517,N_2483);
nand U2557 (N_2557,N_2540,N_2500);
or U2558 (N_2558,N_2534,N_2488);
or U2559 (N_2559,N_2533,N_2510);
or U2560 (N_2560,N_2507,N_2535);
nor U2561 (N_2561,N_2477,N_2523);
and U2562 (N_2562,N_2512,N_2498);
xnor U2563 (N_2563,N_2531,N_2489);
nand U2564 (N_2564,N_2490,N_2478);
nor U2565 (N_2565,N_2482,N_2484);
nor U2566 (N_2566,N_2505,N_2521);
and U2567 (N_2567,N_2549,N_2491);
and U2568 (N_2568,N_2496,N_2511);
nor U2569 (N_2569,N_2514,N_2493);
and U2570 (N_2570,N_2546,N_2528);
xnor U2571 (N_2571,N_2516,N_2495);
nor U2572 (N_2572,N_2524,N_2481);
nand U2573 (N_2573,N_2479,N_2544);
and U2574 (N_2574,N_2539,N_2541);
nand U2575 (N_2575,N_2526,N_2529);
and U2576 (N_2576,N_2504,N_2513);
nor U2577 (N_2577,N_2542,N_2501);
and U2578 (N_2578,N_2499,N_2497);
nor U2579 (N_2579,N_2520,N_2545);
nor U2580 (N_2580,N_2475,N_2480);
or U2581 (N_2581,N_2492,N_2494);
or U2582 (N_2582,N_2532,N_2522);
xnor U2583 (N_2583,N_2537,N_2518);
or U2584 (N_2584,N_2485,N_2547);
or U2585 (N_2585,N_2519,N_2527);
nor U2586 (N_2586,N_2476,N_2536);
and U2587 (N_2587,N_2506,N_2488);
or U2588 (N_2588,N_2515,N_2534);
or U2589 (N_2589,N_2496,N_2488);
xnor U2590 (N_2590,N_2531,N_2526);
nand U2591 (N_2591,N_2534,N_2545);
nor U2592 (N_2592,N_2523,N_2544);
or U2593 (N_2593,N_2505,N_2546);
and U2594 (N_2594,N_2505,N_2477);
nor U2595 (N_2595,N_2506,N_2492);
or U2596 (N_2596,N_2477,N_2489);
nor U2597 (N_2597,N_2486,N_2517);
xor U2598 (N_2598,N_2491,N_2539);
nand U2599 (N_2599,N_2549,N_2539);
or U2600 (N_2600,N_2527,N_2479);
nor U2601 (N_2601,N_2536,N_2518);
nor U2602 (N_2602,N_2492,N_2524);
nand U2603 (N_2603,N_2516,N_2480);
or U2604 (N_2604,N_2499,N_2529);
xor U2605 (N_2605,N_2525,N_2483);
and U2606 (N_2606,N_2515,N_2477);
or U2607 (N_2607,N_2478,N_2477);
and U2608 (N_2608,N_2506,N_2530);
nand U2609 (N_2609,N_2487,N_2511);
and U2610 (N_2610,N_2548,N_2544);
nand U2611 (N_2611,N_2475,N_2517);
and U2612 (N_2612,N_2519,N_2501);
and U2613 (N_2613,N_2529,N_2532);
nor U2614 (N_2614,N_2546,N_2518);
nor U2615 (N_2615,N_2522,N_2511);
nand U2616 (N_2616,N_2529,N_2490);
nor U2617 (N_2617,N_2488,N_2546);
and U2618 (N_2618,N_2543,N_2479);
and U2619 (N_2619,N_2526,N_2506);
or U2620 (N_2620,N_2537,N_2475);
xnor U2621 (N_2621,N_2502,N_2499);
xnor U2622 (N_2622,N_2543,N_2488);
nor U2623 (N_2623,N_2488,N_2518);
nand U2624 (N_2624,N_2482,N_2499);
nand U2625 (N_2625,N_2593,N_2598);
and U2626 (N_2626,N_2585,N_2570);
or U2627 (N_2627,N_2557,N_2581);
nor U2628 (N_2628,N_2555,N_2573);
nand U2629 (N_2629,N_2571,N_2580);
nand U2630 (N_2630,N_2591,N_2586);
xnor U2631 (N_2631,N_2582,N_2603);
nor U2632 (N_2632,N_2552,N_2597);
or U2633 (N_2633,N_2588,N_2604);
and U2634 (N_2634,N_2620,N_2596);
nor U2635 (N_2635,N_2601,N_2583);
or U2636 (N_2636,N_2575,N_2567);
and U2637 (N_2637,N_2613,N_2616);
or U2638 (N_2638,N_2599,N_2594);
or U2639 (N_2639,N_2622,N_2558);
nor U2640 (N_2640,N_2587,N_2589);
or U2641 (N_2641,N_2605,N_2595);
nand U2642 (N_2642,N_2553,N_2615);
nor U2643 (N_2643,N_2561,N_2564);
xnor U2644 (N_2644,N_2617,N_2554);
nor U2645 (N_2645,N_2584,N_2614);
nand U2646 (N_2646,N_2563,N_2611);
nor U2647 (N_2647,N_2574,N_2556);
or U2648 (N_2648,N_2569,N_2577);
or U2649 (N_2649,N_2576,N_2607);
nor U2650 (N_2650,N_2562,N_2623);
nor U2651 (N_2651,N_2568,N_2560);
nor U2652 (N_2652,N_2559,N_2624);
or U2653 (N_2653,N_2612,N_2610);
nand U2654 (N_2654,N_2565,N_2608);
or U2655 (N_2655,N_2551,N_2619);
nand U2656 (N_2656,N_2618,N_2566);
or U2657 (N_2657,N_2578,N_2602);
or U2658 (N_2658,N_2600,N_2590);
nor U2659 (N_2659,N_2572,N_2579);
nor U2660 (N_2660,N_2592,N_2606);
or U2661 (N_2661,N_2550,N_2621);
xor U2662 (N_2662,N_2609,N_2588);
nor U2663 (N_2663,N_2566,N_2600);
nand U2664 (N_2664,N_2592,N_2614);
or U2665 (N_2665,N_2606,N_2620);
and U2666 (N_2666,N_2621,N_2603);
or U2667 (N_2667,N_2613,N_2586);
and U2668 (N_2668,N_2552,N_2594);
and U2669 (N_2669,N_2583,N_2568);
and U2670 (N_2670,N_2550,N_2584);
nand U2671 (N_2671,N_2619,N_2550);
nor U2672 (N_2672,N_2553,N_2578);
or U2673 (N_2673,N_2567,N_2616);
nor U2674 (N_2674,N_2580,N_2621);
nor U2675 (N_2675,N_2575,N_2576);
nand U2676 (N_2676,N_2606,N_2611);
nor U2677 (N_2677,N_2589,N_2583);
xor U2678 (N_2678,N_2610,N_2558);
xor U2679 (N_2679,N_2557,N_2592);
xor U2680 (N_2680,N_2557,N_2559);
or U2681 (N_2681,N_2623,N_2580);
and U2682 (N_2682,N_2600,N_2574);
nor U2683 (N_2683,N_2596,N_2581);
nand U2684 (N_2684,N_2617,N_2605);
nor U2685 (N_2685,N_2612,N_2578);
or U2686 (N_2686,N_2566,N_2615);
nand U2687 (N_2687,N_2587,N_2597);
or U2688 (N_2688,N_2586,N_2553);
or U2689 (N_2689,N_2618,N_2613);
nand U2690 (N_2690,N_2598,N_2614);
nor U2691 (N_2691,N_2618,N_2575);
xor U2692 (N_2692,N_2552,N_2601);
or U2693 (N_2693,N_2582,N_2558);
or U2694 (N_2694,N_2586,N_2624);
or U2695 (N_2695,N_2575,N_2569);
nor U2696 (N_2696,N_2552,N_2578);
or U2697 (N_2697,N_2559,N_2598);
nor U2698 (N_2698,N_2623,N_2554);
and U2699 (N_2699,N_2572,N_2557);
nand U2700 (N_2700,N_2675,N_2689);
nor U2701 (N_2701,N_2658,N_2630);
and U2702 (N_2702,N_2633,N_2664);
xnor U2703 (N_2703,N_2699,N_2693);
nand U2704 (N_2704,N_2634,N_2668);
or U2705 (N_2705,N_2666,N_2690);
nand U2706 (N_2706,N_2661,N_2655);
nand U2707 (N_2707,N_2679,N_2644);
or U2708 (N_2708,N_2687,N_2695);
nor U2709 (N_2709,N_2694,N_2692);
and U2710 (N_2710,N_2626,N_2645);
and U2711 (N_2711,N_2691,N_2659);
or U2712 (N_2712,N_2641,N_2651);
and U2713 (N_2713,N_2680,N_2677);
or U2714 (N_2714,N_2642,N_2698);
nor U2715 (N_2715,N_2647,N_2681);
or U2716 (N_2716,N_2696,N_2672);
or U2717 (N_2717,N_2636,N_2652);
and U2718 (N_2718,N_2654,N_2629);
nor U2719 (N_2719,N_2678,N_2631);
xnor U2720 (N_2720,N_2684,N_2628);
nand U2721 (N_2721,N_2640,N_2697);
nor U2722 (N_2722,N_2635,N_2673);
or U2723 (N_2723,N_2669,N_2627);
and U2724 (N_2724,N_2667,N_2648);
nand U2725 (N_2725,N_2656,N_2649);
or U2726 (N_2726,N_2663,N_2632);
nand U2727 (N_2727,N_2657,N_2639);
xor U2728 (N_2728,N_2625,N_2637);
nand U2729 (N_2729,N_2674,N_2670);
or U2730 (N_2730,N_2643,N_2665);
or U2731 (N_2731,N_2688,N_2650);
xor U2732 (N_2732,N_2660,N_2676);
or U2733 (N_2733,N_2638,N_2646);
xor U2734 (N_2734,N_2685,N_2653);
nand U2735 (N_2735,N_2686,N_2682);
or U2736 (N_2736,N_2671,N_2662);
or U2737 (N_2737,N_2683,N_2655);
nand U2738 (N_2738,N_2644,N_2630);
nand U2739 (N_2739,N_2693,N_2667);
nand U2740 (N_2740,N_2644,N_2699);
or U2741 (N_2741,N_2681,N_2653);
or U2742 (N_2742,N_2693,N_2631);
and U2743 (N_2743,N_2664,N_2671);
and U2744 (N_2744,N_2669,N_2691);
nand U2745 (N_2745,N_2641,N_2659);
nor U2746 (N_2746,N_2646,N_2692);
or U2747 (N_2747,N_2696,N_2666);
and U2748 (N_2748,N_2655,N_2641);
nand U2749 (N_2749,N_2643,N_2651);
nor U2750 (N_2750,N_2697,N_2632);
nor U2751 (N_2751,N_2660,N_2625);
or U2752 (N_2752,N_2682,N_2688);
and U2753 (N_2753,N_2634,N_2695);
and U2754 (N_2754,N_2673,N_2694);
nor U2755 (N_2755,N_2695,N_2657);
or U2756 (N_2756,N_2694,N_2677);
nand U2757 (N_2757,N_2655,N_2637);
and U2758 (N_2758,N_2642,N_2635);
xnor U2759 (N_2759,N_2674,N_2640);
or U2760 (N_2760,N_2672,N_2656);
or U2761 (N_2761,N_2668,N_2633);
nand U2762 (N_2762,N_2628,N_2642);
and U2763 (N_2763,N_2678,N_2681);
or U2764 (N_2764,N_2656,N_2697);
or U2765 (N_2765,N_2664,N_2662);
nor U2766 (N_2766,N_2653,N_2670);
and U2767 (N_2767,N_2647,N_2672);
and U2768 (N_2768,N_2634,N_2694);
nor U2769 (N_2769,N_2673,N_2689);
nand U2770 (N_2770,N_2691,N_2645);
and U2771 (N_2771,N_2670,N_2696);
and U2772 (N_2772,N_2673,N_2684);
or U2773 (N_2773,N_2656,N_2653);
or U2774 (N_2774,N_2685,N_2676);
nand U2775 (N_2775,N_2705,N_2758);
nand U2776 (N_2776,N_2750,N_2716);
or U2777 (N_2777,N_2757,N_2751);
and U2778 (N_2778,N_2710,N_2768);
nor U2779 (N_2779,N_2717,N_2735);
and U2780 (N_2780,N_2743,N_2737);
nor U2781 (N_2781,N_2729,N_2766);
xor U2782 (N_2782,N_2709,N_2772);
or U2783 (N_2783,N_2714,N_2731);
and U2784 (N_2784,N_2707,N_2715);
or U2785 (N_2785,N_2747,N_2769);
and U2786 (N_2786,N_2721,N_2754);
xor U2787 (N_2787,N_2755,N_2718);
nor U2788 (N_2788,N_2703,N_2700);
and U2789 (N_2789,N_2704,N_2761);
nor U2790 (N_2790,N_2736,N_2738);
and U2791 (N_2791,N_2765,N_2763);
nand U2792 (N_2792,N_2701,N_2726);
and U2793 (N_2793,N_2774,N_2764);
nand U2794 (N_2794,N_2746,N_2712);
nor U2795 (N_2795,N_2760,N_2748);
or U2796 (N_2796,N_2730,N_2752);
and U2797 (N_2797,N_2732,N_2702);
or U2798 (N_2798,N_2741,N_2739);
nor U2799 (N_2799,N_2745,N_2767);
and U2800 (N_2800,N_2706,N_2756);
nand U2801 (N_2801,N_2734,N_2762);
and U2802 (N_2802,N_2740,N_2722);
nand U2803 (N_2803,N_2727,N_2742);
nand U2804 (N_2804,N_2725,N_2759);
nor U2805 (N_2805,N_2713,N_2711);
or U2806 (N_2806,N_2720,N_2770);
and U2807 (N_2807,N_2728,N_2753);
nand U2808 (N_2808,N_2723,N_2744);
and U2809 (N_2809,N_2724,N_2773);
or U2810 (N_2810,N_2771,N_2719);
and U2811 (N_2811,N_2733,N_2708);
nor U2812 (N_2812,N_2749,N_2751);
nand U2813 (N_2813,N_2770,N_2750);
nand U2814 (N_2814,N_2767,N_2737);
and U2815 (N_2815,N_2713,N_2744);
nor U2816 (N_2816,N_2744,N_2738);
nand U2817 (N_2817,N_2705,N_2771);
and U2818 (N_2818,N_2726,N_2734);
xnor U2819 (N_2819,N_2765,N_2743);
nor U2820 (N_2820,N_2714,N_2748);
xor U2821 (N_2821,N_2730,N_2734);
nand U2822 (N_2822,N_2725,N_2727);
nand U2823 (N_2823,N_2757,N_2761);
and U2824 (N_2824,N_2762,N_2703);
or U2825 (N_2825,N_2736,N_2744);
and U2826 (N_2826,N_2741,N_2736);
nor U2827 (N_2827,N_2721,N_2709);
nor U2828 (N_2828,N_2774,N_2738);
nor U2829 (N_2829,N_2710,N_2724);
or U2830 (N_2830,N_2723,N_2740);
and U2831 (N_2831,N_2722,N_2756);
and U2832 (N_2832,N_2704,N_2772);
or U2833 (N_2833,N_2761,N_2700);
xnor U2834 (N_2834,N_2743,N_2706);
xnor U2835 (N_2835,N_2773,N_2762);
nor U2836 (N_2836,N_2711,N_2753);
nor U2837 (N_2837,N_2723,N_2743);
nor U2838 (N_2838,N_2769,N_2705);
and U2839 (N_2839,N_2701,N_2732);
xor U2840 (N_2840,N_2731,N_2702);
or U2841 (N_2841,N_2704,N_2751);
nor U2842 (N_2842,N_2748,N_2724);
or U2843 (N_2843,N_2747,N_2716);
and U2844 (N_2844,N_2752,N_2741);
or U2845 (N_2845,N_2716,N_2719);
nand U2846 (N_2846,N_2716,N_2752);
nand U2847 (N_2847,N_2728,N_2751);
or U2848 (N_2848,N_2740,N_2766);
xor U2849 (N_2849,N_2754,N_2735);
or U2850 (N_2850,N_2833,N_2783);
nand U2851 (N_2851,N_2803,N_2793);
nand U2852 (N_2852,N_2825,N_2820);
nand U2853 (N_2853,N_2776,N_2812);
nor U2854 (N_2854,N_2824,N_2777);
or U2855 (N_2855,N_2837,N_2804);
or U2856 (N_2856,N_2838,N_2828);
and U2857 (N_2857,N_2781,N_2818);
nand U2858 (N_2858,N_2835,N_2841);
nor U2859 (N_2859,N_2827,N_2836);
nor U2860 (N_2860,N_2821,N_2849);
nor U2861 (N_2861,N_2780,N_2813);
nand U2862 (N_2862,N_2834,N_2801);
and U2863 (N_2863,N_2811,N_2847);
and U2864 (N_2864,N_2778,N_2815);
and U2865 (N_2865,N_2846,N_2782);
and U2866 (N_2866,N_2805,N_2848);
nor U2867 (N_2867,N_2843,N_2819);
nor U2868 (N_2868,N_2845,N_2794);
nand U2869 (N_2869,N_2814,N_2786);
nand U2870 (N_2870,N_2788,N_2817);
nor U2871 (N_2871,N_2799,N_2829);
xnor U2872 (N_2872,N_2816,N_2798);
nand U2873 (N_2873,N_2807,N_2787);
nor U2874 (N_2874,N_2826,N_2810);
nand U2875 (N_2875,N_2789,N_2802);
or U2876 (N_2876,N_2839,N_2823);
nand U2877 (N_2877,N_2800,N_2795);
and U2878 (N_2878,N_2775,N_2779);
xnor U2879 (N_2879,N_2822,N_2796);
nor U2880 (N_2880,N_2808,N_2840);
nand U2881 (N_2881,N_2790,N_2809);
or U2882 (N_2882,N_2831,N_2791);
and U2883 (N_2883,N_2844,N_2832);
nor U2884 (N_2884,N_2785,N_2797);
nor U2885 (N_2885,N_2784,N_2842);
and U2886 (N_2886,N_2830,N_2792);
nor U2887 (N_2887,N_2806,N_2811);
nand U2888 (N_2888,N_2815,N_2837);
nor U2889 (N_2889,N_2803,N_2823);
and U2890 (N_2890,N_2792,N_2802);
nand U2891 (N_2891,N_2819,N_2814);
xor U2892 (N_2892,N_2794,N_2832);
and U2893 (N_2893,N_2812,N_2790);
or U2894 (N_2894,N_2787,N_2836);
nor U2895 (N_2895,N_2792,N_2839);
or U2896 (N_2896,N_2777,N_2847);
nor U2897 (N_2897,N_2787,N_2822);
and U2898 (N_2898,N_2840,N_2823);
nor U2899 (N_2899,N_2777,N_2815);
nor U2900 (N_2900,N_2844,N_2801);
xor U2901 (N_2901,N_2796,N_2801);
or U2902 (N_2902,N_2809,N_2778);
nand U2903 (N_2903,N_2821,N_2795);
nor U2904 (N_2904,N_2821,N_2820);
nor U2905 (N_2905,N_2778,N_2834);
nand U2906 (N_2906,N_2798,N_2792);
nand U2907 (N_2907,N_2826,N_2817);
nand U2908 (N_2908,N_2846,N_2843);
and U2909 (N_2909,N_2846,N_2839);
xnor U2910 (N_2910,N_2825,N_2783);
xor U2911 (N_2911,N_2835,N_2848);
nor U2912 (N_2912,N_2810,N_2823);
or U2913 (N_2913,N_2830,N_2833);
nor U2914 (N_2914,N_2840,N_2839);
nor U2915 (N_2915,N_2842,N_2827);
nand U2916 (N_2916,N_2785,N_2794);
nor U2917 (N_2917,N_2825,N_2776);
nand U2918 (N_2918,N_2826,N_2791);
or U2919 (N_2919,N_2801,N_2802);
xnor U2920 (N_2920,N_2784,N_2809);
nand U2921 (N_2921,N_2786,N_2846);
nor U2922 (N_2922,N_2823,N_2789);
nor U2923 (N_2923,N_2784,N_2793);
and U2924 (N_2924,N_2809,N_2816);
and U2925 (N_2925,N_2860,N_2855);
nor U2926 (N_2926,N_2873,N_2906);
nand U2927 (N_2927,N_2851,N_2911);
or U2928 (N_2928,N_2915,N_2905);
and U2929 (N_2929,N_2882,N_2852);
nand U2930 (N_2930,N_2912,N_2922);
nor U2931 (N_2931,N_2854,N_2864);
or U2932 (N_2932,N_2874,N_2878);
nand U2933 (N_2933,N_2885,N_2892);
and U2934 (N_2934,N_2895,N_2861);
nor U2935 (N_2935,N_2857,N_2897);
nand U2936 (N_2936,N_2877,N_2862);
or U2937 (N_2937,N_2871,N_2868);
nor U2938 (N_2938,N_2881,N_2883);
xor U2939 (N_2939,N_2924,N_2914);
nand U2940 (N_2940,N_2894,N_2888);
nor U2941 (N_2941,N_2853,N_2904);
and U2942 (N_2942,N_2867,N_2907);
and U2943 (N_2943,N_2916,N_2887);
nor U2944 (N_2944,N_2923,N_2858);
nand U2945 (N_2945,N_2875,N_2890);
and U2946 (N_2946,N_2921,N_2901);
nor U2947 (N_2947,N_2896,N_2876);
nor U2948 (N_2948,N_2886,N_2908);
nand U2949 (N_2949,N_2893,N_2910);
or U2950 (N_2950,N_2900,N_2870);
nor U2951 (N_2951,N_2899,N_2913);
and U2952 (N_2952,N_2889,N_2863);
nand U2953 (N_2953,N_2869,N_2859);
nand U2954 (N_2954,N_2879,N_2919);
nor U2955 (N_2955,N_2918,N_2866);
and U2956 (N_2956,N_2850,N_2903);
and U2957 (N_2957,N_2902,N_2872);
and U2958 (N_2958,N_2856,N_2909);
or U2959 (N_2959,N_2865,N_2920);
and U2960 (N_2960,N_2898,N_2884);
and U2961 (N_2961,N_2880,N_2917);
or U2962 (N_2962,N_2891,N_2864);
or U2963 (N_2963,N_2893,N_2868);
or U2964 (N_2964,N_2868,N_2907);
nand U2965 (N_2965,N_2923,N_2908);
and U2966 (N_2966,N_2883,N_2915);
nor U2967 (N_2967,N_2886,N_2865);
or U2968 (N_2968,N_2874,N_2886);
and U2969 (N_2969,N_2874,N_2860);
xnor U2970 (N_2970,N_2883,N_2895);
or U2971 (N_2971,N_2907,N_2880);
or U2972 (N_2972,N_2915,N_2917);
nor U2973 (N_2973,N_2899,N_2872);
or U2974 (N_2974,N_2913,N_2896);
and U2975 (N_2975,N_2865,N_2863);
or U2976 (N_2976,N_2904,N_2880);
nor U2977 (N_2977,N_2910,N_2851);
and U2978 (N_2978,N_2916,N_2854);
nand U2979 (N_2979,N_2903,N_2901);
nor U2980 (N_2980,N_2924,N_2915);
nor U2981 (N_2981,N_2919,N_2882);
or U2982 (N_2982,N_2900,N_2914);
nand U2983 (N_2983,N_2857,N_2858);
or U2984 (N_2984,N_2852,N_2924);
nand U2985 (N_2985,N_2852,N_2865);
or U2986 (N_2986,N_2880,N_2872);
nand U2987 (N_2987,N_2896,N_2894);
and U2988 (N_2988,N_2886,N_2924);
or U2989 (N_2989,N_2865,N_2850);
and U2990 (N_2990,N_2861,N_2894);
nor U2991 (N_2991,N_2921,N_2858);
xor U2992 (N_2992,N_2878,N_2857);
nor U2993 (N_2993,N_2869,N_2887);
xnor U2994 (N_2994,N_2895,N_2914);
and U2995 (N_2995,N_2920,N_2889);
or U2996 (N_2996,N_2912,N_2870);
nand U2997 (N_2997,N_2882,N_2912);
or U2998 (N_2998,N_2896,N_2889);
or U2999 (N_2999,N_2873,N_2887);
and UO_0 (O_0,N_2941,N_2952);
nor UO_1 (O_1,N_2983,N_2929);
nand UO_2 (O_2,N_2979,N_2982);
and UO_3 (O_3,N_2964,N_2945);
and UO_4 (O_4,N_2933,N_2932);
xor UO_5 (O_5,N_2928,N_2944);
and UO_6 (O_6,N_2930,N_2963);
nor UO_7 (O_7,N_2981,N_2965);
xor UO_8 (O_8,N_2975,N_2988);
and UO_9 (O_9,N_2967,N_2958);
or UO_10 (O_10,N_2971,N_2956);
and UO_11 (O_11,N_2977,N_2940);
nand UO_12 (O_12,N_2994,N_2931);
nand UO_13 (O_13,N_2974,N_2991);
or UO_14 (O_14,N_2987,N_2978);
nor UO_15 (O_15,N_2939,N_2984);
nand UO_16 (O_16,N_2989,N_2969);
xor UO_17 (O_17,N_2960,N_2976);
xnor UO_18 (O_18,N_2934,N_2951);
nand UO_19 (O_19,N_2942,N_2937);
nand UO_20 (O_20,N_2986,N_2938);
nor UO_21 (O_21,N_2997,N_2955);
nor UO_22 (O_22,N_2980,N_2949);
nor UO_23 (O_23,N_2927,N_2966);
nor UO_24 (O_24,N_2935,N_2990);
and UO_25 (O_25,N_2999,N_2985);
nor UO_26 (O_26,N_2993,N_2948);
and UO_27 (O_27,N_2953,N_2995);
xor UO_28 (O_28,N_2954,N_2992);
nand UO_29 (O_29,N_2998,N_2970);
nand UO_30 (O_30,N_2957,N_2968);
or UO_31 (O_31,N_2936,N_2996);
and UO_32 (O_32,N_2961,N_2959);
nor UO_33 (O_33,N_2947,N_2926);
and UO_34 (O_34,N_2973,N_2946);
or UO_35 (O_35,N_2962,N_2950);
nand UO_36 (O_36,N_2972,N_2943);
or UO_37 (O_37,N_2925,N_2975);
xor UO_38 (O_38,N_2963,N_2984);
nand UO_39 (O_39,N_2942,N_2991);
nor UO_40 (O_40,N_2949,N_2972);
and UO_41 (O_41,N_2973,N_2936);
and UO_42 (O_42,N_2964,N_2958);
and UO_43 (O_43,N_2960,N_2945);
nor UO_44 (O_44,N_2966,N_2983);
nand UO_45 (O_45,N_2942,N_2947);
nor UO_46 (O_46,N_2957,N_2938);
or UO_47 (O_47,N_2940,N_2961);
and UO_48 (O_48,N_2974,N_2965);
nor UO_49 (O_49,N_2932,N_2958);
and UO_50 (O_50,N_2925,N_2983);
and UO_51 (O_51,N_2992,N_2980);
nor UO_52 (O_52,N_2943,N_2951);
or UO_53 (O_53,N_2970,N_2983);
or UO_54 (O_54,N_2938,N_2937);
nand UO_55 (O_55,N_2968,N_2991);
and UO_56 (O_56,N_2960,N_2991);
or UO_57 (O_57,N_2965,N_2953);
and UO_58 (O_58,N_2981,N_2925);
nor UO_59 (O_59,N_2927,N_2939);
nand UO_60 (O_60,N_2985,N_2981);
nand UO_61 (O_61,N_2969,N_2998);
or UO_62 (O_62,N_2956,N_2976);
xor UO_63 (O_63,N_2965,N_2958);
nand UO_64 (O_64,N_2974,N_2971);
or UO_65 (O_65,N_2956,N_2979);
xnor UO_66 (O_66,N_2951,N_2947);
nor UO_67 (O_67,N_2961,N_2930);
and UO_68 (O_68,N_2984,N_2928);
and UO_69 (O_69,N_2955,N_2936);
nor UO_70 (O_70,N_2987,N_2955);
and UO_71 (O_71,N_2952,N_2959);
and UO_72 (O_72,N_2959,N_2996);
nand UO_73 (O_73,N_2987,N_2931);
nand UO_74 (O_74,N_2941,N_2933);
nor UO_75 (O_75,N_2931,N_2937);
or UO_76 (O_76,N_2960,N_2930);
and UO_77 (O_77,N_2981,N_2982);
and UO_78 (O_78,N_2944,N_2971);
or UO_79 (O_79,N_2948,N_2942);
nor UO_80 (O_80,N_2971,N_2999);
nor UO_81 (O_81,N_2950,N_2985);
and UO_82 (O_82,N_2928,N_2942);
or UO_83 (O_83,N_2979,N_2965);
nand UO_84 (O_84,N_2936,N_2952);
nand UO_85 (O_85,N_2933,N_2967);
and UO_86 (O_86,N_2972,N_2966);
and UO_87 (O_87,N_2943,N_2963);
and UO_88 (O_88,N_2952,N_2935);
and UO_89 (O_89,N_2963,N_2942);
or UO_90 (O_90,N_2977,N_2935);
nor UO_91 (O_91,N_2980,N_2967);
nor UO_92 (O_92,N_2968,N_2998);
and UO_93 (O_93,N_2942,N_2951);
or UO_94 (O_94,N_2970,N_2944);
nand UO_95 (O_95,N_2993,N_2959);
xnor UO_96 (O_96,N_2989,N_2984);
nor UO_97 (O_97,N_2996,N_2931);
and UO_98 (O_98,N_2939,N_2960);
nand UO_99 (O_99,N_2940,N_2981);
xor UO_100 (O_100,N_2945,N_2925);
nor UO_101 (O_101,N_2943,N_2961);
or UO_102 (O_102,N_2990,N_2936);
or UO_103 (O_103,N_2981,N_2939);
and UO_104 (O_104,N_2971,N_2928);
and UO_105 (O_105,N_2928,N_2939);
nor UO_106 (O_106,N_2955,N_2928);
nor UO_107 (O_107,N_2948,N_2960);
nor UO_108 (O_108,N_2962,N_2965);
nor UO_109 (O_109,N_2962,N_2988);
or UO_110 (O_110,N_2960,N_2996);
or UO_111 (O_111,N_2982,N_2955);
and UO_112 (O_112,N_2942,N_2975);
and UO_113 (O_113,N_2997,N_2944);
nor UO_114 (O_114,N_2980,N_2993);
nor UO_115 (O_115,N_2995,N_2941);
or UO_116 (O_116,N_2999,N_2943);
and UO_117 (O_117,N_2999,N_2941);
and UO_118 (O_118,N_2980,N_2954);
or UO_119 (O_119,N_2974,N_2941);
nand UO_120 (O_120,N_2953,N_2960);
or UO_121 (O_121,N_2962,N_2954);
nor UO_122 (O_122,N_2949,N_2948);
or UO_123 (O_123,N_2941,N_2989);
nor UO_124 (O_124,N_2942,N_2940);
or UO_125 (O_125,N_2928,N_2974);
nor UO_126 (O_126,N_2953,N_2979);
nand UO_127 (O_127,N_2973,N_2996);
nor UO_128 (O_128,N_2981,N_2943);
or UO_129 (O_129,N_2934,N_2995);
and UO_130 (O_130,N_2935,N_2967);
nand UO_131 (O_131,N_2948,N_2989);
nor UO_132 (O_132,N_2980,N_2948);
nor UO_133 (O_133,N_2929,N_2981);
and UO_134 (O_134,N_2939,N_2995);
nand UO_135 (O_135,N_2986,N_2990);
or UO_136 (O_136,N_2947,N_2981);
nand UO_137 (O_137,N_2973,N_2939);
and UO_138 (O_138,N_2987,N_2946);
nand UO_139 (O_139,N_2974,N_2976);
or UO_140 (O_140,N_2937,N_2953);
or UO_141 (O_141,N_2975,N_2974);
or UO_142 (O_142,N_2961,N_2979);
nor UO_143 (O_143,N_2989,N_2991);
nor UO_144 (O_144,N_2935,N_2968);
and UO_145 (O_145,N_2971,N_2930);
nor UO_146 (O_146,N_2973,N_2961);
xor UO_147 (O_147,N_2949,N_2927);
or UO_148 (O_148,N_2981,N_2944);
nand UO_149 (O_149,N_2998,N_2932);
nand UO_150 (O_150,N_2932,N_2968);
nor UO_151 (O_151,N_2959,N_2980);
nor UO_152 (O_152,N_2929,N_2926);
xnor UO_153 (O_153,N_2986,N_2948);
and UO_154 (O_154,N_2940,N_2954);
nor UO_155 (O_155,N_2970,N_2927);
xnor UO_156 (O_156,N_2990,N_2959);
and UO_157 (O_157,N_2925,N_2987);
or UO_158 (O_158,N_2960,N_2966);
or UO_159 (O_159,N_2993,N_2935);
or UO_160 (O_160,N_2960,N_2997);
nand UO_161 (O_161,N_2988,N_2969);
or UO_162 (O_162,N_2996,N_2925);
nand UO_163 (O_163,N_2949,N_2963);
xor UO_164 (O_164,N_2944,N_2946);
nor UO_165 (O_165,N_2941,N_2947);
nor UO_166 (O_166,N_2993,N_2952);
nor UO_167 (O_167,N_2934,N_2944);
xor UO_168 (O_168,N_2964,N_2988);
or UO_169 (O_169,N_2949,N_2975);
and UO_170 (O_170,N_2991,N_2998);
and UO_171 (O_171,N_2954,N_2986);
nor UO_172 (O_172,N_2987,N_2959);
nor UO_173 (O_173,N_2982,N_2975);
nor UO_174 (O_174,N_2930,N_2998);
nand UO_175 (O_175,N_2955,N_2971);
nand UO_176 (O_176,N_2980,N_2964);
or UO_177 (O_177,N_2939,N_2999);
and UO_178 (O_178,N_2954,N_2959);
and UO_179 (O_179,N_2937,N_2966);
xnor UO_180 (O_180,N_2999,N_2970);
and UO_181 (O_181,N_2925,N_2938);
and UO_182 (O_182,N_2941,N_2968);
or UO_183 (O_183,N_2989,N_2942);
or UO_184 (O_184,N_2943,N_2993);
or UO_185 (O_185,N_2952,N_2960);
nand UO_186 (O_186,N_2969,N_2964);
nand UO_187 (O_187,N_2970,N_2980);
nor UO_188 (O_188,N_2995,N_2952);
or UO_189 (O_189,N_2977,N_2996);
nor UO_190 (O_190,N_2952,N_2974);
nand UO_191 (O_191,N_2957,N_2986);
nor UO_192 (O_192,N_2980,N_2999);
nand UO_193 (O_193,N_2944,N_2974);
or UO_194 (O_194,N_2961,N_2985);
nor UO_195 (O_195,N_2927,N_2998);
or UO_196 (O_196,N_2981,N_2997);
or UO_197 (O_197,N_2932,N_2999);
or UO_198 (O_198,N_2950,N_2977);
and UO_199 (O_199,N_2968,N_2992);
or UO_200 (O_200,N_2980,N_2930);
xor UO_201 (O_201,N_2998,N_2959);
nor UO_202 (O_202,N_2964,N_2944);
and UO_203 (O_203,N_2925,N_2933);
or UO_204 (O_204,N_2929,N_2978);
or UO_205 (O_205,N_2982,N_2957);
and UO_206 (O_206,N_2995,N_2943);
nor UO_207 (O_207,N_2972,N_2938);
and UO_208 (O_208,N_2992,N_2965);
nand UO_209 (O_209,N_2963,N_2944);
and UO_210 (O_210,N_2952,N_2981);
or UO_211 (O_211,N_2937,N_2993);
nand UO_212 (O_212,N_2966,N_2935);
nand UO_213 (O_213,N_2930,N_2991);
nand UO_214 (O_214,N_2999,N_2979);
or UO_215 (O_215,N_2935,N_2936);
xnor UO_216 (O_216,N_2948,N_2992);
and UO_217 (O_217,N_2930,N_2964);
nand UO_218 (O_218,N_2945,N_2984);
nor UO_219 (O_219,N_2973,N_2972);
or UO_220 (O_220,N_2967,N_2939);
and UO_221 (O_221,N_2946,N_2937);
and UO_222 (O_222,N_2994,N_2933);
nor UO_223 (O_223,N_2993,N_2964);
nand UO_224 (O_224,N_2959,N_2929);
nor UO_225 (O_225,N_2972,N_2976);
nand UO_226 (O_226,N_2992,N_2986);
nor UO_227 (O_227,N_2984,N_2950);
xor UO_228 (O_228,N_2961,N_2926);
xnor UO_229 (O_229,N_2943,N_2982);
and UO_230 (O_230,N_2989,N_2986);
or UO_231 (O_231,N_2968,N_2962);
nand UO_232 (O_232,N_2930,N_2937);
or UO_233 (O_233,N_2963,N_2934);
nor UO_234 (O_234,N_2964,N_2960);
nor UO_235 (O_235,N_2993,N_2949);
nor UO_236 (O_236,N_2931,N_2930);
or UO_237 (O_237,N_2994,N_2986);
or UO_238 (O_238,N_2967,N_2959);
nor UO_239 (O_239,N_2993,N_2995);
or UO_240 (O_240,N_2970,N_2968);
and UO_241 (O_241,N_2958,N_2945);
and UO_242 (O_242,N_2997,N_2950);
nand UO_243 (O_243,N_2974,N_2978);
nand UO_244 (O_244,N_2983,N_2959);
nand UO_245 (O_245,N_2963,N_2957);
nand UO_246 (O_246,N_2926,N_2927);
or UO_247 (O_247,N_2930,N_2926);
nand UO_248 (O_248,N_2970,N_2991);
and UO_249 (O_249,N_2950,N_2925);
and UO_250 (O_250,N_2965,N_2935);
or UO_251 (O_251,N_2988,N_2940);
and UO_252 (O_252,N_2939,N_2968);
or UO_253 (O_253,N_2958,N_2980);
and UO_254 (O_254,N_2987,N_2928);
nand UO_255 (O_255,N_2927,N_2962);
or UO_256 (O_256,N_2944,N_2977);
nor UO_257 (O_257,N_2973,N_2938);
or UO_258 (O_258,N_2985,N_2969);
and UO_259 (O_259,N_2998,N_2975);
nor UO_260 (O_260,N_2930,N_2936);
nand UO_261 (O_261,N_2947,N_2953);
nor UO_262 (O_262,N_2969,N_2966);
nor UO_263 (O_263,N_2960,N_2975);
or UO_264 (O_264,N_2985,N_2972);
or UO_265 (O_265,N_2955,N_2937);
nor UO_266 (O_266,N_2966,N_2938);
and UO_267 (O_267,N_2941,N_2950);
nor UO_268 (O_268,N_2968,N_2966);
xor UO_269 (O_269,N_2994,N_2962);
or UO_270 (O_270,N_2943,N_2964);
nand UO_271 (O_271,N_2989,N_2993);
and UO_272 (O_272,N_2989,N_2950);
nand UO_273 (O_273,N_2962,N_2972);
xnor UO_274 (O_274,N_2954,N_2995);
or UO_275 (O_275,N_2996,N_2956);
or UO_276 (O_276,N_2955,N_2990);
or UO_277 (O_277,N_2978,N_2928);
and UO_278 (O_278,N_2984,N_2982);
xnor UO_279 (O_279,N_2989,N_2982);
and UO_280 (O_280,N_2981,N_2999);
and UO_281 (O_281,N_2956,N_2947);
nor UO_282 (O_282,N_2971,N_2986);
nor UO_283 (O_283,N_2954,N_2982);
or UO_284 (O_284,N_2998,N_2939);
xnor UO_285 (O_285,N_2949,N_2999);
or UO_286 (O_286,N_2988,N_2968);
and UO_287 (O_287,N_2943,N_2930);
and UO_288 (O_288,N_2991,N_2962);
nand UO_289 (O_289,N_2959,N_2946);
and UO_290 (O_290,N_2965,N_2943);
and UO_291 (O_291,N_2948,N_2964);
and UO_292 (O_292,N_2928,N_2956);
nand UO_293 (O_293,N_2990,N_2950);
or UO_294 (O_294,N_2932,N_2970);
or UO_295 (O_295,N_2951,N_2928);
and UO_296 (O_296,N_2932,N_2926);
nand UO_297 (O_297,N_2987,N_2984);
and UO_298 (O_298,N_2943,N_2957);
nand UO_299 (O_299,N_2927,N_2980);
nor UO_300 (O_300,N_2937,N_2980);
nand UO_301 (O_301,N_2931,N_2938);
nand UO_302 (O_302,N_2983,N_2965);
nand UO_303 (O_303,N_2988,N_2997);
nor UO_304 (O_304,N_2954,N_2957);
nand UO_305 (O_305,N_2933,N_2993);
or UO_306 (O_306,N_2939,N_2936);
or UO_307 (O_307,N_2973,N_2993);
or UO_308 (O_308,N_2953,N_2959);
xor UO_309 (O_309,N_2925,N_2973);
or UO_310 (O_310,N_2984,N_2966);
nand UO_311 (O_311,N_2982,N_2932);
and UO_312 (O_312,N_2970,N_2948);
and UO_313 (O_313,N_2979,N_2958);
nor UO_314 (O_314,N_2978,N_2932);
nand UO_315 (O_315,N_2974,N_2999);
or UO_316 (O_316,N_2947,N_2965);
and UO_317 (O_317,N_2994,N_2978);
nand UO_318 (O_318,N_2949,N_2957);
or UO_319 (O_319,N_2988,N_2945);
xnor UO_320 (O_320,N_2935,N_2962);
nand UO_321 (O_321,N_2998,N_2940);
nand UO_322 (O_322,N_2974,N_2980);
or UO_323 (O_323,N_2945,N_2948);
nand UO_324 (O_324,N_2960,N_2993);
nand UO_325 (O_325,N_2987,N_2998);
nor UO_326 (O_326,N_2948,N_2943);
nand UO_327 (O_327,N_2974,N_2925);
xor UO_328 (O_328,N_2985,N_2980);
nand UO_329 (O_329,N_2932,N_2997);
xnor UO_330 (O_330,N_2929,N_2995);
or UO_331 (O_331,N_2935,N_2955);
and UO_332 (O_332,N_2967,N_2961);
and UO_333 (O_333,N_2993,N_2946);
and UO_334 (O_334,N_2999,N_2964);
nor UO_335 (O_335,N_2983,N_2962);
nor UO_336 (O_336,N_2955,N_2966);
nand UO_337 (O_337,N_2937,N_2968);
or UO_338 (O_338,N_2971,N_2962);
xor UO_339 (O_339,N_2927,N_2968);
nand UO_340 (O_340,N_2951,N_2941);
and UO_341 (O_341,N_2983,N_2930);
nor UO_342 (O_342,N_2941,N_2926);
xor UO_343 (O_343,N_2971,N_2990);
or UO_344 (O_344,N_2929,N_2988);
nor UO_345 (O_345,N_2987,N_2983);
and UO_346 (O_346,N_2954,N_2929);
and UO_347 (O_347,N_2982,N_2929);
or UO_348 (O_348,N_2968,N_2973);
or UO_349 (O_349,N_2988,N_2955);
or UO_350 (O_350,N_2933,N_2950);
nor UO_351 (O_351,N_2929,N_2969);
xor UO_352 (O_352,N_2942,N_2990);
nor UO_353 (O_353,N_2930,N_2985);
nand UO_354 (O_354,N_2934,N_2997);
nand UO_355 (O_355,N_2964,N_2961);
and UO_356 (O_356,N_2972,N_2988);
and UO_357 (O_357,N_2941,N_2937);
xnor UO_358 (O_358,N_2951,N_2971);
nor UO_359 (O_359,N_2987,N_2992);
nor UO_360 (O_360,N_2952,N_2971);
or UO_361 (O_361,N_2974,N_2988);
xnor UO_362 (O_362,N_2986,N_2974);
and UO_363 (O_363,N_2943,N_2938);
nor UO_364 (O_364,N_2953,N_2935);
nor UO_365 (O_365,N_2959,N_2972);
or UO_366 (O_366,N_2951,N_2968);
or UO_367 (O_367,N_2943,N_2927);
nor UO_368 (O_368,N_2954,N_2964);
nand UO_369 (O_369,N_2971,N_2972);
and UO_370 (O_370,N_2936,N_2940);
nand UO_371 (O_371,N_2953,N_2983);
or UO_372 (O_372,N_2949,N_2990);
nand UO_373 (O_373,N_2976,N_2979);
nor UO_374 (O_374,N_2973,N_2955);
and UO_375 (O_375,N_2987,N_2994);
and UO_376 (O_376,N_2941,N_2994);
nand UO_377 (O_377,N_2947,N_2961);
and UO_378 (O_378,N_2981,N_2963);
or UO_379 (O_379,N_2953,N_2987);
xor UO_380 (O_380,N_2967,N_2938);
nor UO_381 (O_381,N_2986,N_2970);
xor UO_382 (O_382,N_2932,N_2947);
or UO_383 (O_383,N_2965,N_2969);
or UO_384 (O_384,N_2937,N_2999);
nand UO_385 (O_385,N_2989,N_2959);
or UO_386 (O_386,N_2960,N_2982);
nand UO_387 (O_387,N_2999,N_2986);
nand UO_388 (O_388,N_2937,N_2977);
xor UO_389 (O_389,N_2983,N_2963);
nand UO_390 (O_390,N_2965,N_2941);
nand UO_391 (O_391,N_2945,N_2940);
or UO_392 (O_392,N_2987,N_2932);
nor UO_393 (O_393,N_2964,N_2995);
nand UO_394 (O_394,N_2927,N_2954);
xor UO_395 (O_395,N_2978,N_2963);
nor UO_396 (O_396,N_2936,N_2951);
and UO_397 (O_397,N_2944,N_2978);
nor UO_398 (O_398,N_2985,N_2990);
nand UO_399 (O_399,N_2942,N_2952);
and UO_400 (O_400,N_2971,N_2959);
nand UO_401 (O_401,N_2937,N_2962);
nand UO_402 (O_402,N_2998,N_2993);
nand UO_403 (O_403,N_2994,N_2995);
and UO_404 (O_404,N_2972,N_2970);
nand UO_405 (O_405,N_2978,N_2956);
or UO_406 (O_406,N_2935,N_2987);
nor UO_407 (O_407,N_2931,N_2939);
xor UO_408 (O_408,N_2947,N_2969);
nand UO_409 (O_409,N_2954,N_2991);
or UO_410 (O_410,N_2960,N_2926);
and UO_411 (O_411,N_2963,N_2964);
or UO_412 (O_412,N_2972,N_2975);
or UO_413 (O_413,N_2960,N_2929);
nor UO_414 (O_414,N_2945,N_2989);
nor UO_415 (O_415,N_2951,N_2996);
or UO_416 (O_416,N_2942,N_2934);
and UO_417 (O_417,N_2973,N_2964);
and UO_418 (O_418,N_2988,N_2947);
nand UO_419 (O_419,N_2983,N_2968);
and UO_420 (O_420,N_2964,N_2966);
or UO_421 (O_421,N_2986,N_2926);
nor UO_422 (O_422,N_2942,N_2945);
nand UO_423 (O_423,N_2954,N_2978);
nor UO_424 (O_424,N_2963,N_2974);
and UO_425 (O_425,N_2998,N_2981);
nand UO_426 (O_426,N_2964,N_2984);
nand UO_427 (O_427,N_2969,N_2956);
nor UO_428 (O_428,N_2971,N_2969);
nand UO_429 (O_429,N_2942,N_2968);
xnor UO_430 (O_430,N_2989,N_2936);
nor UO_431 (O_431,N_2985,N_2943);
nand UO_432 (O_432,N_2949,N_2976);
and UO_433 (O_433,N_2999,N_2947);
and UO_434 (O_434,N_2984,N_2953);
nor UO_435 (O_435,N_2933,N_2999);
xnor UO_436 (O_436,N_2975,N_2932);
nand UO_437 (O_437,N_2925,N_2978);
and UO_438 (O_438,N_2959,N_2973);
and UO_439 (O_439,N_2953,N_2939);
xor UO_440 (O_440,N_2928,N_2960);
nor UO_441 (O_441,N_2945,N_2934);
or UO_442 (O_442,N_2986,N_2952);
nand UO_443 (O_443,N_2941,N_2963);
nor UO_444 (O_444,N_2937,N_2948);
nor UO_445 (O_445,N_2968,N_2977);
nor UO_446 (O_446,N_2926,N_2984);
nor UO_447 (O_447,N_2977,N_2974);
nand UO_448 (O_448,N_2975,N_2928);
or UO_449 (O_449,N_2980,N_2973);
nand UO_450 (O_450,N_2931,N_2998);
nor UO_451 (O_451,N_2989,N_2981);
xnor UO_452 (O_452,N_2974,N_2943);
and UO_453 (O_453,N_2951,N_2988);
or UO_454 (O_454,N_2957,N_2956);
or UO_455 (O_455,N_2986,N_2949);
nand UO_456 (O_456,N_2960,N_2968);
or UO_457 (O_457,N_2996,N_2927);
nand UO_458 (O_458,N_2973,N_2927);
or UO_459 (O_459,N_2954,N_2930);
and UO_460 (O_460,N_2971,N_2983);
xnor UO_461 (O_461,N_2985,N_2938);
and UO_462 (O_462,N_2976,N_2933);
xor UO_463 (O_463,N_2948,N_2953);
nand UO_464 (O_464,N_2936,N_2956);
nand UO_465 (O_465,N_2957,N_2975);
or UO_466 (O_466,N_2937,N_2982);
nand UO_467 (O_467,N_2942,N_2976);
or UO_468 (O_468,N_2963,N_2979);
xnor UO_469 (O_469,N_2991,N_2949);
or UO_470 (O_470,N_2940,N_2999);
nand UO_471 (O_471,N_2938,N_2933);
nand UO_472 (O_472,N_2990,N_2972);
nor UO_473 (O_473,N_2970,N_2955);
and UO_474 (O_474,N_2976,N_2939);
and UO_475 (O_475,N_2974,N_2949);
xor UO_476 (O_476,N_2930,N_2932);
nor UO_477 (O_477,N_2993,N_2940);
xor UO_478 (O_478,N_2980,N_2947);
nor UO_479 (O_479,N_2976,N_2951);
and UO_480 (O_480,N_2975,N_2973);
or UO_481 (O_481,N_2931,N_2977);
nor UO_482 (O_482,N_2995,N_2979);
and UO_483 (O_483,N_2997,N_2980);
nand UO_484 (O_484,N_2934,N_2952);
and UO_485 (O_485,N_2974,N_2989);
or UO_486 (O_486,N_2986,N_2965);
nand UO_487 (O_487,N_2983,N_2990);
nor UO_488 (O_488,N_2992,N_2945);
and UO_489 (O_489,N_2978,N_2976);
and UO_490 (O_490,N_2991,N_2955);
nand UO_491 (O_491,N_2962,N_2985);
nand UO_492 (O_492,N_2984,N_2959);
xnor UO_493 (O_493,N_2949,N_2964);
and UO_494 (O_494,N_2932,N_2934);
nor UO_495 (O_495,N_2985,N_2944);
or UO_496 (O_496,N_2972,N_2984);
or UO_497 (O_497,N_2994,N_2973);
nor UO_498 (O_498,N_2998,N_2949);
nor UO_499 (O_499,N_2988,N_2939);
endmodule