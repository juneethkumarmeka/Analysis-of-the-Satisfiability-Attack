module basic_500_3000_500_5_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
and U0 (N_0,In_172,In_332);
nand U1 (N_1,In_387,In_276);
nor U2 (N_2,In_17,In_2);
xnor U3 (N_3,In_296,In_429);
nand U4 (N_4,In_383,In_430);
and U5 (N_5,In_490,In_201);
and U6 (N_6,In_465,In_63);
nor U7 (N_7,In_377,In_27);
and U8 (N_8,In_420,In_141);
and U9 (N_9,In_102,In_93);
nand U10 (N_10,In_174,In_125);
nand U11 (N_11,In_135,In_266);
nand U12 (N_12,In_223,In_319);
nand U13 (N_13,In_12,In_385);
nor U14 (N_14,In_391,In_483);
nand U15 (N_15,In_106,In_225);
and U16 (N_16,In_448,In_340);
nand U17 (N_17,In_426,In_15);
nand U18 (N_18,In_386,In_226);
nor U19 (N_19,In_488,In_124);
and U20 (N_20,In_357,In_424);
or U21 (N_21,In_220,In_161);
and U22 (N_22,In_209,In_51);
nor U23 (N_23,In_344,In_140);
or U24 (N_24,In_303,In_212);
nor U25 (N_25,In_41,In_360);
nand U26 (N_26,In_192,In_193);
nor U27 (N_27,In_302,In_300);
nand U28 (N_28,In_86,In_283);
nand U29 (N_29,In_455,In_261);
or U30 (N_30,In_312,In_180);
and U31 (N_31,In_458,In_177);
nand U32 (N_32,In_454,In_11);
or U33 (N_33,In_217,In_197);
or U34 (N_34,In_148,In_482);
nor U35 (N_35,In_3,In_229);
nand U36 (N_36,In_37,In_423);
nand U37 (N_37,In_290,In_356);
or U38 (N_38,In_309,In_122);
nor U39 (N_39,In_292,In_390);
and U40 (N_40,In_61,In_85);
or U41 (N_41,In_145,In_6);
or U42 (N_42,In_405,In_313);
xnor U43 (N_43,In_108,In_453);
nor U44 (N_44,In_185,In_471);
nand U45 (N_45,In_165,In_13);
nor U46 (N_46,In_128,In_379);
nor U47 (N_47,In_236,In_411);
and U48 (N_48,In_282,In_477);
nand U49 (N_49,In_474,In_353);
and U50 (N_50,In_263,In_243);
or U51 (N_51,In_358,In_33);
or U52 (N_52,In_475,In_421);
nor U53 (N_53,In_468,In_191);
nor U54 (N_54,In_327,In_381);
nor U55 (N_55,In_246,In_50);
and U56 (N_56,In_1,In_259);
or U57 (N_57,In_160,In_244);
and U58 (N_58,In_162,In_378);
nor U59 (N_59,In_368,In_324);
nand U60 (N_60,In_175,In_239);
and U61 (N_61,In_214,In_142);
or U62 (N_62,In_401,In_485);
nor U63 (N_63,In_186,In_402);
and U64 (N_64,In_345,In_395);
or U65 (N_65,In_484,In_205);
nor U66 (N_66,In_204,In_4);
nor U67 (N_67,In_10,In_370);
nor U68 (N_68,In_473,In_157);
nor U69 (N_69,In_417,In_317);
nand U70 (N_70,In_167,In_275);
nand U71 (N_71,In_406,In_288);
or U72 (N_72,In_121,In_469);
or U73 (N_73,In_437,In_211);
nor U74 (N_74,In_447,In_190);
nor U75 (N_75,In_457,In_235);
nor U76 (N_76,In_334,In_278);
and U77 (N_77,In_419,In_99);
nor U78 (N_78,In_376,In_154);
nand U79 (N_79,In_168,In_48);
and U80 (N_80,In_431,In_388);
nor U81 (N_81,In_155,In_80);
and U82 (N_82,In_22,In_316);
or U83 (N_83,In_314,In_260);
nand U84 (N_84,In_100,In_361);
nor U85 (N_85,In_77,In_371);
and U86 (N_86,In_144,In_151);
and U87 (N_87,In_202,In_75);
nand U88 (N_88,In_240,In_364);
nor U89 (N_89,In_291,In_68);
nor U90 (N_90,In_28,In_335);
or U91 (N_91,In_216,In_105);
nor U92 (N_92,In_92,In_5);
and U93 (N_93,In_481,In_224);
or U94 (N_94,In_67,In_72);
nor U95 (N_95,In_306,In_115);
nor U96 (N_96,In_228,In_264);
and U97 (N_97,In_479,In_416);
nor U98 (N_98,In_436,In_251);
and U99 (N_99,In_445,In_427);
and U100 (N_100,In_103,In_491);
and U101 (N_101,In_472,In_396);
nand U102 (N_102,In_196,In_298);
or U103 (N_103,In_34,In_389);
or U104 (N_104,In_284,In_373);
and U105 (N_105,In_267,In_362);
or U106 (N_106,In_495,In_494);
nand U107 (N_107,In_158,In_16);
nor U108 (N_108,In_59,In_42);
or U109 (N_109,In_60,In_98);
and U110 (N_110,In_54,In_435);
or U111 (N_111,In_375,In_127);
nor U112 (N_112,In_394,In_255);
nor U113 (N_113,In_78,In_207);
or U114 (N_114,In_354,In_408);
nand U115 (N_115,In_338,In_150);
xor U116 (N_116,In_110,In_176);
or U117 (N_117,In_130,In_412);
or U118 (N_118,In_82,In_287);
or U119 (N_119,In_463,In_136);
nor U120 (N_120,In_210,In_308);
or U121 (N_121,In_182,In_164);
nor U122 (N_122,In_297,In_462);
nand U123 (N_123,In_315,In_109);
and U124 (N_124,In_333,In_199);
or U125 (N_125,In_45,In_97);
or U126 (N_126,In_258,In_111);
or U127 (N_127,In_64,In_400);
nor U128 (N_128,In_194,In_83);
and U129 (N_129,In_200,In_21);
and U130 (N_130,In_112,In_183);
or U131 (N_131,In_245,In_178);
and U132 (N_132,In_152,In_66);
and U133 (N_133,In_466,In_318);
nor U134 (N_134,In_407,In_137);
or U135 (N_135,In_262,In_337);
nand U136 (N_136,In_404,In_277);
and U137 (N_137,In_90,In_399);
nor U138 (N_138,In_114,In_269);
nor U139 (N_139,In_286,In_215);
or U140 (N_140,In_329,In_163);
and U141 (N_141,In_230,In_374);
nor U142 (N_142,In_38,In_169);
nand U143 (N_143,In_131,In_166);
or U144 (N_144,In_272,In_227);
nor U145 (N_145,In_91,In_76);
or U146 (N_146,In_233,In_134);
and U147 (N_147,In_498,In_460);
and U148 (N_148,In_330,In_149);
nor U149 (N_149,In_281,In_119);
nor U150 (N_150,In_222,In_380);
or U151 (N_151,In_118,In_311);
and U152 (N_152,In_273,In_349);
nor U153 (N_153,In_486,In_359);
nor U154 (N_154,In_237,In_31);
nor U155 (N_155,In_451,In_257);
nand U156 (N_156,In_30,In_449);
nand U157 (N_157,In_0,In_304);
or U158 (N_158,In_123,In_295);
or U159 (N_159,In_250,In_139);
nand U160 (N_160,In_331,In_265);
and U161 (N_161,In_171,In_52);
or U162 (N_162,In_428,In_397);
nor U163 (N_163,In_84,In_274);
nand U164 (N_164,In_293,In_73);
nand U165 (N_165,In_241,In_415);
and U166 (N_166,In_188,In_206);
and U167 (N_167,In_443,In_328);
or U168 (N_168,In_96,In_232);
nor U169 (N_169,In_46,In_289);
nor U170 (N_170,In_476,In_366);
and U171 (N_171,In_307,In_94);
nor U172 (N_172,In_231,In_170);
nor U173 (N_173,In_414,In_325);
nor U174 (N_174,In_104,In_489);
nand U175 (N_175,In_467,In_184);
nor U176 (N_176,In_497,In_35);
or U177 (N_177,In_20,In_252);
or U178 (N_178,In_310,In_441);
nand U179 (N_179,In_18,In_446);
nor U180 (N_180,In_280,In_496);
or U181 (N_181,In_153,In_74);
nand U182 (N_182,In_363,In_321);
nand U183 (N_183,In_81,In_242);
nand U184 (N_184,In_187,In_234);
nand U185 (N_185,In_351,In_343);
nor U186 (N_186,In_179,In_254);
or U187 (N_187,In_117,In_159);
nor U188 (N_188,In_355,In_470);
or U189 (N_189,In_203,In_24);
nand U190 (N_190,In_299,In_53);
nand U191 (N_191,In_219,In_101);
and U192 (N_192,In_221,In_478);
or U193 (N_193,In_14,In_39);
and U194 (N_194,In_464,In_392);
nor U195 (N_195,In_36,In_26);
or U196 (N_196,In_301,In_372);
and U197 (N_197,In_294,In_433);
or U198 (N_198,In_320,In_238);
or U199 (N_199,In_322,In_339);
nor U200 (N_200,In_365,In_456);
nand U201 (N_201,In_253,In_249);
or U202 (N_202,In_285,In_393);
or U203 (N_203,In_323,In_347);
nand U204 (N_204,In_70,In_132);
and U205 (N_205,In_146,In_352);
nand U206 (N_206,In_7,In_55);
nand U207 (N_207,In_450,In_218);
and U208 (N_208,In_247,In_422);
nor U209 (N_209,In_369,In_29);
nand U210 (N_210,In_346,In_65);
and U211 (N_211,In_189,In_107);
or U212 (N_212,In_348,In_87);
or U213 (N_213,In_147,In_116);
and U214 (N_214,In_425,In_181);
and U215 (N_215,In_47,In_129);
and U216 (N_216,In_58,In_213);
or U217 (N_217,In_133,In_440);
nand U218 (N_218,In_25,In_268);
nor U219 (N_219,In_499,In_195);
or U220 (N_220,In_382,In_62);
nor U221 (N_221,In_88,In_432);
nand U222 (N_222,In_126,In_57);
nor U223 (N_223,In_270,In_89);
nor U224 (N_224,In_492,In_438);
or U225 (N_225,In_49,In_208);
and U226 (N_226,In_198,In_350);
and U227 (N_227,In_156,In_409);
and U228 (N_228,In_9,In_23);
and U229 (N_229,In_44,In_410);
nor U230 (N_230,In_32,In_40);
nor U231 (N_231,In_69,In_487);
nor U232 (N_232,In_113,In_143);
and U233 (N_233,In_138,In_367);
or U234 (N_234,In_19,In_120);
or U235 (N_235,In_442,In_384);
nor U236 (N_236,In_403,In_279);
or U237 (N_237,In_341,In_342);
nor U238 (N_238,In_413,In_493);
and U239 (N_239,In_43,In_173);
and U240 (N_240,In_326,In_444);
nor U241 (N_241,In_459,In_56);
nor U242 (N_242,In_398,In_461);
and U243 (N_243,In_256,In_452);
or U244 (N_244,In_271,In_434);
and U245 (N_245,In_439,In_480);
or U246 (N_246,In_95,In_305);
or U247 (N_247,In_8,In_248);
nor U248 (N_248,In_71,In_336);
nand U249 (N_249,In_418,In_79);
nand U250 (N_250,In_195,In_62);
or U251 (N_251,In_78,In_191);
and U252 (N_252,In_281,In_458);
nand U253 (N_253,In_297,In_94);
and U254 (N_254,In_58,In_379);
and U255 (N_255,In_496,In_430);
nor U256 (N_256,In_360,In_497);
and U257 (N_257,In_121,In_133);
and U258 (N_258,In_377,In_90);
nand U259 (N_259,In_234,In_27);
and U260 (N_260,In_320,In_431);
nor U261 (N_261,In_335,In_155);
or U262 (N_262,In_440,In_420);
or U263 (N_263,In_497,In_14);
nor U264 (N_264,In_101,In_183);
and U265 (N_265,In_360,In_332);
and U266 (N_266,In_328,In_157);
nand U267 (N_267,In_148,In_49);
or U268 (N_268,In_16,In_253);
nand U269 (N_269,In_403,In_204);
and U270 (N_270,In_277,In_190);
nand U271 (N_271,In_0,In_128);
and U272 (N_272,In_215,In_320);
and U273 (N_273,In_483,In_112);
and U274 (N_274,In_86,In_104);
and U275 (N_275,In_37,In_465);
nand U276 (N_276,In_124,In_164);
nor U277 (N_277,In_459,In_336);
or U278 (N_278,In_375,In_100);
and U279 (N_279,In_304,In_136);
nand U280 (N_280,In_278,In_146);
or U281 (N_281,In_17,In_88);
and U282 (N_282,In_332,In_141);
nor U283 (N_283,In_38,In_14);
and U284 (N_284,In_291,In_485);
nor U285 (N_285,In_457,In_482);
and U286 (N_286,In_380,In_429);
or U287 (N_287,In_11,In_85);
nand U288 (N_288,In_370,In_108);
and U289 (N_289,In_85,In_291);
and U290 (N_290,In_99,In_177);
nor U291 (N_291,In_9,In_279);
xnor U292 (N_292,In_411,In_197);
nor U293 (N_293,In_15,In_333);
or U294 (N_294,In_351,In_205);
and U295 (N_295,In_443,In_154);
or U296 (N_296,In_148,In_186);
nand U297 (N_297,In_90,In_388);
nor U298 (N_298,In_205,In_267);
or U299 (N_299,In_333,In_387);
xnor U300 (N_300,In_209,In_181);
nand U301 (N_301,In_235,In_86);
or U302 (N_302,In_265,In_397);
or U303 (N_303,In_96,In_267);
and U304 (N_304,In_21,In_204);
nand U305 (N_305,In_41,In_354);
or U306 (N_306,In_306,In_200);
nor U307 (N_307,In_164,In_192);
nand U308 (N_308,In_400,In_302);
nand U309 (N_309,In_480,In_282);
nor U310 (N_310,In_246,In_410);
or U311 (N_311,In_257,In_70);
nor U312 (N_312,In_483,In_58);
or U313 (N_313,In_332,In_54);
and U314 (N_314,In_303,In_291);
nand U315 (N_315,In_220,In_434);
nand U316 (N_316,In_166,In_440);
nor U317 (N_317,In_370,In_143);
xor U318 (N_318,In_158,In_143);
nand U319 (N_319,In_20,In_476);
nand U320 (N_320,In_207,In_428);
and U321 (N_321,In_308,In_322);
nor U322 (N_322,In_109,In_345);
or U323 (N_323,In_218,In_126);
or U324 (N_324,In_245,In_223);
nand U325 (N_325,In_150,In_100);
nand U326 (N_326,In_406,In_265);
or U327 (N_327,In_372,In_204);
and U328 (N_328,In_262,In_499);
nand U329 (N_329,In_308,In_468);
nand U330 (N_330,In_265,In_427);
nand U331 (N_331,In_81,In_434);
or U332 (N_332,In_189,In_301);
nand U333 (N_333,In_237,In_266);
and U334 (N_334,In_105,In_487);
nor U335 (N_335,In_226,In_230);
and U336 (N_336,In_412,In_115);
and U337 (N_337,In_98,In_4);
or U338 (N_338,In_259,In_258);
nor U339 (N_339,In_275,In_270);
nand U340 (N_340,In_426,In_393);
and U341 (N_341,In_381,In_314);
and U342 (N_342,In_376,In_364);
nor U343 (N_343,In_398,In_308);
nor U344 (N_344,In_341,In_209);
nor U345 (N_345,In_90,In_115);
or U346 (N_346,In_249,In_156);
or U347 (N_347,In_484,In_163);
nor U348 (N_348,In_279,In_280);
nand U349 (N_349,In_278,In_153);
nor U350 (N_350,In_360,In_378);
or U351 (N_351,In_158,In_345);
and U352 (N_352,In_462,In_53);
nor U353 (N_353,In_17,In_438);
nor U354 (N_354,In_414,In_458);
nand U355 (N_355,In_479,In_471);
nand U356 (N_356,In_12,In_365);
and U357 (N_357,In_370,In_105);
and U358 (N_358,In_417,In_341);
or U359 (N_359,In_55,In_412);
and U360 (N_360,In_203,In_389);
and U361 (N_361,In_129,In_94);
nor U362 (N_362,In_302,In_196);
or U363 (N_363,In_234,In_219);
nor U364 (N_364,In_441,In_474);
nand U365 (N_365,In_146,In_400);
or U366 (N_366,In_474,In_153);
nor U367 (N_367,In_202,In_229);
or U368 (N_368,In_411,In_117);
and U369 (N_369,In_496,In_174);
or U370 (N_370,In_48,In_170);
nand U371 (N_371,In_58,In_104);
and U372 (N_372,In_316,In_66);
or U373 (N_373,In_422,In_109);
nor U374 (N_374,In_334,In_284);
nand U375 (N_375,In_1,In_422);
nor U376 (N_376,In_420,In_5);
and U377 (N_377,In_48,In_355);
or U378 (N_378,In_439,In_200);
and U379 (N_379,In_150,In_125);
nand U380 (N_380,In_182,In_446);
nand U381 (N_381,In_436,In_425);
nor U382 (N_382,In_134,In_380);
nor U383 (N_383,In_207,In_166);
or U384 (N_384,In_440,In_450);
or U385 (N_385,In_188,In_353);
or U386 (N_386,In_158,In_303);
and U387 (N_387,In_16,In_458);
and U388 (N_388,In_232,In_111);
nor U389 (N_389,In_102,In_331);
nand U390 (N_390,In_132,In_359);
nor U391 (N_391,In_12,In_443);
nor U392 (N_392,In_140,In_192);
xor U393 (N_393,In_140,In_186);
nor U394 (N_394,In_203,In_354);
or U395 (N_395,In_228,In_458);
nand U396 (N_396,In_423,In_103);
nand U397 (N_397,In_51,In_359);
or U398 (N_398,In_178,In_484);
nor U399 (N_399,In_207,In_94);
and U400 (N_400,In_288,In_458);
or U401 (N_401,In_396,In_404);
nand U402 (N_402,In_28,In_89);
or U403 (N_403,In_41,In_129);
or U404 (N_404,In_19,In_259);
and U405 (N_405,In_227,In_417);
or U406 (N_406,In_70,In_457);
nand U407 (N_407,In_197,In_344);
or U408 (N_408,In_94,In_84);
or U409 (N_409,In_222,In_466);
nor U410 (N_410,In_389,In_29);
nor U411 (N_411,In_392,In_307);
nand U412 (N_412,In_347,In_419);
nor U413 (N_413,In_136,In_258);
nand U414 (N_414,In_219,In_12);
or U415 (N_415,In_69,In_359);
and U416 (N_416,In_480,In_431);
nand U417 (N_417,In_369,In_327);
nor U418 (N_418,In_24,In_165);
nor U419 (N_419,In_214,In_340);
or U420 (N_420,In_62,In_191);
nor U421 (N_421,In_285,In_413);
or U422 (N_422,In_375,In_456);
or U423 (N_423,In_338,In_120);
nor U424 (N_424,In_25,In_405);
and U425 (N_425,In_139,In_401);
nand U426 (N_426,In_294,In_426);
and U427 (N_427,In_110,In_101);
nand U428 (N_428,In_415,In_302);
nor U429 (N_429,In_258,In_141);
nand U430 (N_430,In_143,In_37);
or U431 (N_431,In_423,In_368);
and U432 (N_432,In_117,In_406);
nor U433 (N_433,In_458,In_196);
and U434 (N_434,In_199,In_411);
nor U435 (N_435,In_128,In_350);
nand U436 (N_436,In_86,In_414);
nor U437 (N_437,In_266,In_65);
or U438 (N_438,In_397,In_70);
xor U439 (N_439,In_215,In_8);
nand U440 (N_440,In_102,In_375);
and U441 (N_441,In_295,In_442);
and U442 (N_442,In_53,In_148);
nand U443 (N_443,In_17,In_325);
or U444 (N_444,In_332,In_42);
or U445 (N_445,In_243,In_439);
or U446 (N_446,In_122,In_151);
or U447 (N_447,In_146,In_299);
or U448 (N_448,In_139,In_386);
nor U449 (N_449,In_157,In_250);
nand U450 (N_450,In_429,In_302);
and U451 (N_451,In_99,In_294);
nor U452 (N_452,In_433,In_449);
or U453 (N_453,In_38,In_123);
and U454 (N_454,In_13,In_470);
and U455 (N_455,In_469,In_87);
or U456 (N_456,In_227,In_180);
nor U457 (N_457,In_328,In_212);
nand U458 (N_458,In_413,In_180);
nor U459 (N_459,In_158,In_434);
nor U460 (N_460,In_269,In_321);
and U461 (N_461,In_492,In_101);
nor U462 (N_462,In_362,In_49);
and U463 (N_463,In_341,In_459);
and U464 (N_464,In_326,In_104);
nor U465 (N_465,In_182,In_19);
nand U466 (N_466,In_417,In_313);
nor U467 (N_467,In_293,In_434);
nand U468 (N_468,In_450,In_102);
and U469 (N_469,In_73,In_453);
nor U470 (N_470,In_169,In_437);
or U471 (N_471,In_321,In_276);
nor U472 (N_472,In_172,In_155);
and U473 (N_473,In_29,In_158);
and U474 (N_474,In_147,In_318);
or U475 (N_475,In_39,In_226);
and U476 (N_476,In_224,In_275);
or U477 (N_477,In_336,In_224);
nor U478 (N_478,In_178,In_331);
nor U479 (N_479,In_409,In_275);
nand U480 (N_480,In_129,In_283);
nor U481 (N_481,In_26,In_370);
or U482 (N_482,In_376,In_73);
or U483 (N_483,In_355,In_203);
nand U484 (N_484,In_431,In_274);
nor U485 (N_485,In_389,In_303);
or U486 (N_486,In_50,In_395);
or U487 (N_487,In_131,In_463);
or U488 (N_488,In_426,In_356);
or U489 (N_489,In_66,In_74);
or U490 (N_490,In_212,In_406);
or U491 (N_491,In_90,In_423);
nor U492 (N_492,In_372,In_46);
nor U493 (N_493,In_258,In_167);
or U494 (N_494,In_428,In_359);
and U495 (N_495,In_1,In_95);
or U496 (N_496,In_472,In_2);
nor U497 (N_497,In_205,In_383);
nor U498 (N_498,In_31,In_418);
or U499 (N_499,In_311,In_352);
nor U500 (N_500,In_367,In_264);
and U501 (N_501,In_29,In_328);
nor U502 (N_502,In_478,In_146);
nor U503 (N_503,In_231,In_486);
and U504 (N_504,In_222,In_443);
or U505 (N_505,In_471,In_181);
or U506 (N_506,In_296,In_222);
nand U507 (N_507,In_171,In_486);
or U508 (N_508,In_182,In_437);
or U509 (N_509,In_294,In_122);
nor U510 (N_510,In_354,In_76);
and U511 (N_511,In_482,In_202);
nand U512 (N_512,In_426,In_28);
nor U513 (N_513,In_374,In_394);
nor U514 (N_514,In_8,In_369);
nand U515 (N_515,In_73,In_190);
or U516 (N_516,In_67,In_394);
and U517 (N_517,In_154,In_313);
or U518 (N_518,In_139,In_357);
and U519 (N_519,In_324,In_67);
and U520 (N_520,In_475,In_434);
or U521 (N_521,In_399,In_166);
nand U522 (N_522,In_143,In_291);
nand U523 (N_523,In_385,In_9);
nand U524 (N_524,In_335,In_461);
and U525 (N_525,In_153,In_211);
nand U526 (N_526,In_91,In_112);
or U527 (N_527,In_226,In_163);
and U528 (N_528,In_188,In_303);
and U529 (N_529,In_307,In_115);
and U530 (N_530,In_198,In_459);
nand U531 (N_531,In_142,In_154);
and U532 (N_532,In_442,In_11);
nor U533 (N_533,In_287,In_265);
nor U534 (N_534,In_148,In_0);
or U535 (N_535,In_450,In_160);
nor U536 (N_536,In_31,In_25);
or U537 (N_537,In_292,In_226);
nor U538 (N_538,In_463,In_376);
xnor U539 (N_539,In_366,In_255);
nand U540 (N_540,In_134,In_276);
nor U541 (N_541,In_282,In_331);
and U542 (N_542,In_460,In_477);
and U543 (N_543,In_258,In_255);
nand U544 (N_544,In_430,In_229);
or U545 (N_545,In_281,In_23);
nor U546 (N_546,In_325,In_232);
or U547 (N_547,In_177,In_65);
or U548 (N_548,In_344,In_318);
xnor U549 (N_549,In_487,In_493);
nor U550 (N_550,In_350,In_266);
or U551 (N_551,In_453,In_443);
and U552 (N_552,In_463,In_226);
or U553 (N_553,In_354,In_48);
and U554 (N_554,In_202,In_468);
nor U555 (N_555,In_433,In_448);
xnor U556 (N_556,In_29,In_120);
or U557 (N_557,In_95,In_169);
or U558 (N_558,In_347,In_369);
or U559 (N_559,In_108,In_157);
nand U560 (N_560,In_144,In_142);
or U561 (N_561,In_374,In_217);
nand U562 (N_562,In_437,In_270);
or U563 (N_563,In_161,In_156);
or U564 (N_564,In_491,In_288);
nand U565 (N_565,In_90,In_475);
nor U566 (N_566,In_371,In_45);
nand U567 (N_567,In_44,In_99);
nor U568 (N_568,In_136,In_321);
xor U569 (N_569,In_0,In_18);
or U570 (N_570,In_396,In_252);
and U571 (N_571,In_97,In_11);
xor U572 (N_572,In_86,In_29);
nor U573 (N_573,In_53,In_46);
nor U574 (N_574,In_378,In_170);
nor U575 (N_575,In_103,In_33);
nor U576 (N_576,In_166,In_176);
or U577 (N_577,In_172,In_370);
nand U578 (N_578,In_35,In_301);
nand U579 (N_579,In_246,In_347);
or U580 (N_580,In_33,In_381);
or U581 (N_581,In_460,In_147);
and U582 (N_582,In_357,In_446);
and U583 (N_583,In_410,In_230);
or U584 (N_584,In_210,In_304);
and U585 (N_585,In_128,In_479);
nand U586 (N_586,In_134,In_319);
nor U587 (N_587,In_62,In_312);
nor U588 (N_588,In_497,In_429);
nor U589 (N_589,In_327,In_11);
or U590 (N_590,In_438,In_230);
nand U591 (N_591,In_99,In_312);
nor U592 (N_592,In_179,In_332);
nand U593 (N_593,In_183,In_137);
nor U594 (N_594,In_250,In_4);
and U595 (N_595,In_244,In_206);
and U596 (N_596,In_281,In_285);
and U597 (N_597,In_341,In_151);
or U598 (N_598,In_69,In_431);
nand U599 (N_599,In_105,In_162);
nor U600 (N_600,N_40,N_407);
nand U601 (N_601,N_520,N_304);
nor U602 (N_602,N_411,N_140);
and U603 (N_603,N_591,N_508);
nor U604 (N_604,N_170,N_298);
nor U605 (N_605,N_388,N_317);
nand U606 (N_606,N_153,N_449);
and U607 (N_607,N_325,N_47);
and U608 (N_608,N_496,N_480);
nor U609 (N_609,N_578,N_124);
and U610 (N_610,N_121,N_297);
and U611 (N_611,N_143,N_289);
nand U612 (N_612,N_374,N_115);
nand U613 (N_613,N_426,N_492);
nor U614 (N_614,N_176,N_44);
nor U615 (N_615,N_77,N_250);
and U616 (N_616,N_423,N_180);
nand U617 (N_617,N_228,N_386);
and U618 (N_618,N_100,N_389);
and U619 (N_619,N_406,N_402);
nand U620 (N_620,N_31,N_96);
nand U621 (N_621,N_60,N_438);
and U622 (N_622,N_158,N_547);
nand U623 (N_623,N_391,N_584);
nand U624 (N_624,N_307,N_192);
nor U625 (N_625,N_35,N_225);
nand U626 (N_626,N_369,N_542);
nor U627 (N_627,N_71,N_95);
nand U628 (N_628,N_574,N_446);
and U629 (N_629,N_183,N_18);
or U630 (N_630,N_221,N_427);
or U631 (N_631,N_586,N_175);
and U632 (N_632,N_497,N_309);
nand U633 (N_633,N_530,N_541);
and U634 (N_634,N_569,N_570);
and U635 (N_635,N_0,N_415);
nor U636 (N_636,N_475,N_375);
or U637 (N_637,N_172,N_502);
nor U638 (N_638,N_412,N_74);
nand U639 (N_639,N_258,N_420);
nor U640 (N_640,N_107,N_169);
nand U641 (N_641,N_193,N_568);
or U642 (N_642,N_312,N_105);
nand U643 (N_643,N_13,N_99);
nor U644 (N_644,N_247,N_495);
nand U645 (N_645,N_525,N_413);
nand U646 (N_646,N_396,N_58);
nand U647 (N_647,N_352,N_589);
and U648 (N_648,N_507,N_465);
and U649 (N_649,N_248,N_83);
and U650 (N_650,N_120,N_146);
nor U651 (N_651,N_361,N_364);
nor U652 (N_652,N_365,N_379);
nor U653 (N_653,N_128,N_468);
or U654 (N_654,N_395,N_112);
nor U655 (N_655,N_363,N_417);
nand U656 (N_656,N_503,N_152);
nand U657 (N_657,N_384,N_347);
and U658 (N_658,N_259,N_433);
nand U659 (N_659,N_334,N_182);
nor U660 (N_660,N_538,N_167);
nand U661 (N_661,N_523,N_217);
nor U662 (N_662,N_15,N_42);
nand U663 (N_663,N_482,N_291);
nor U664 (N_664,N_454,N_267);
nand U665 (N_665,N_457,N_571);
or U666 (N_666,N_588,N_283);
nand U667 (N_667,N_87,N_137);
and U668 (N_668,N_491,N_102);
nor U669 (N_669,N_197,N_215);
or U670 (N_670,N_484,N_28);
or U671 (N_671,N_29,N_21);
or U672 (N_672,N_227,N_345);
nand U673 (N_673,N_200,N_108);
or U674 (N_674,N_331,N_275);
or U675 (N_675,N_561,N_80);
nand U676 (N_676,N_382,N_236);
nor U677 (N_677,N_380,N_150);
nor U678 (N_678,N_301,N_26);
or U679 (N_679,N_416,N_220);
and U680 (N_680,N_126,N_276);
nand U681 (N_681,N_323,N_230);
nor U682 (N_682,N_377,N_185);
or U683 (N_683,N_202,N_174);
and U684 (N_684,N_451,N_338);
and U685 (N_685,N_149,N_206);
nor U686 (N_686,N_414,N_277);
nor U687 (N_687,N_593,N_251);
or U688 (N_688,N_543,N_513);
and U689 (N_689,N_293,N_392);
nand U690 (N_690,N_254,N_370);
and U691 (N_691,N_478,N_544);
nor U692 (N_692,N_12,N_390);
nor U693 (N_693,N_66,N_212);
nand U694 (N_694,N_448,N_464);
and U695 (N_695,N_122,N_255);
nor U696 (N_696,N_272,N_303);
and U697 (N_697,N_4,N_597);
nand U698 (N_698,N_581,N_490);
and U699 (N_699,N_592,N_257);
or U700 (N_700,N_311,N_555);
nand U701 (N_701,N_342,N_243);
and U702 (N_702,N_210,N_245);
or U703 (N_703,N_563,N_231);
nor U704 (N_704,N_337,N_287);
or U705 (N_705,N_110,N_373);
nor U706 (N_706,N_204,N_136);
nand U707 (N_707,N_285,N_599);
nand U708 (N_708,N_385,N_1);
xnor U709 (N_709,N_548,N_50);
and U710 (N_710,N_5,N_512);
and U711 (N_711,N_177,N_346);
and U712 (N_712,N_41,N_526);
or U713 (N_713,N_239,N_145);
or U714 (N_714,N_57,N_418);
nor U715 (N_715,N_442,N_226);
nor U716 (N_716,N_559,N_32);
or U717 (N_717,N_376,N_598);
nor U718 (N_718,N_203,N_518);
and U719 (N_719,N_531,N_279);
nand U720 (N_720,N_196,N_522);
or U721 (N_721,N_359,N_408);
or U722 (N_722,N_129,N_16);
and U723 (N_723,N_280,N_378);
nand U724 (N_724,N_444,N_90);
or U725 (N_725,N_357,N_54);
xor U726 (N_726,N_216,N_349);
or U727 (N_727,N_560,N_97);
nor U728 (N_728,N_135,N_425);
nand U729 (N_729,N_333,N_314);
and U730 (N_730,N_383,N_264);
or U731 (N_731,N_493,N_51);
nor U732 (N_732,N_340,N_580);
nand U733 (N_733,N_450,N_458);
and U734 (N_734,N_144,N_274);
nor U735 (N_735,N_156,N_306);
and U736 (N_736,N_266,N_324);
nand U737 (N_737,N_8,N_515);
nor U738 (N_738,N_188,N_562);
or U739 (N_739,N_223,N_371);
nand U740 (N_740,N_56,N_461);
and U741 (N_741,N_286,N_318);
nand U742 (N_742,N_2,N_64);
or U743 (N_743,N_147,N_539);
nor U744 (N_744,N_157,N_30);
nor U745 (N_745,N_558,N_320);
nor U746 (N_746,N_62,N_394);
nand U747 (N_747,N_387,N_595);
and U748 (N_748,N_545,N_190);
nor U749 (N_749,N_269,N_114);
and U750 (N_750,N_583,N_3);
nand U751 (N_751,N_330,N_82);
or U752 (N_752,N_294,N_455);
nand U753 (N_753,N_585,N_39);
nor U754 (N_754,N_53,N_9);
nor U755 (N_755,N_315,N_399);
or U756 (N_756,N_271,N_73);
or U757 (N_757,N_473,N_381);
or U758 (N_758,N_161,N_358);
nor U759 (N_759,N_510,N_19);
nand U760 (N_760,N_155,N_205);
or U761 (N_761,N_529,N_403);
or U762 (N_762,N_339,N_404);
and U763 (N_763,N_499,N_201);
and U764 (N_764,N_445,N_93);
or U765 (N_765,N_509,N_63);
and U766 (N_766,N_38,N_437);
or U767 (N_767,N_292,N_505);
nor U768 (N_768,N_186,N_139);
or U769 (N_769,N_488,N_75);
xnor U770 (N_770,N_441,N_372);
nand U771 (N_771,N_332,N_104);
and U772 (N_772,N_244,N_327);
or U773 (N_773,N_151,N_207);
nand U774 (N_774,N_498,N_500);
or U775 (N_775,N_308,N_10);
nor U776 (N_776,N_78,N_299);
nor U777 (N_777,N_282,N_519);
nor U778 (N_778,N_23,N_256);
nand U779 (N_779,N_37,N_262);
nor U780 (N_780,N_431,N_536);
or U781 (N_781,N_296,N_288);
nor U782 (N_782,N_187,N_131);
or U783 (N_783,N_443,N_34);
nor U784 (N_784,N_224,N_46);
nand U785 (N_785,N_511,N_535);
nor U786 (N_786,N_326,N_424);
nor U787 (N_787,N_166,N_409);
nand U788 (N_788,N_240,N_472);
and U789 (N_789,N_477,N_329);
or U790 (N_790,N_86,N_527);
or U791 (N_791,N_350,N_551);
and U792 (N_792,N_469,N_577);
nor U793 (N_793,N_165,N_232);
nor U794 (N_794,N_194,N_343);
nand U795 (N_795,N_141,N_434);
nand U796 (N_796,N_134,N_321);
or U797 (N_797,N_103,N_265);
and U798 (N_798,N_397,N_302);
or U799 (N_799,N_55,N_460);
nand U800 (N_800,N_322,N_459);
and U801 (N_801,N_237,N_366);
and U802 (N_802,N_582,N_476);
nor U803 (N_803,N_516,N_351);
or U804 (N_804,N_113,N_43);
nor U805 (N_805,N_159,N_52);
nand U806 (N_806,N_341,N_70);
or U807 (N_807,N_123,N_20);
or U808 (N_808,N_181,N_25);
and U809 (N_809,N_487,N_494);
nor U810 (N_810,N_191,N_534);
nand U811 (N_811,N_504,N_118);
or U812 (N_812,N_179,N_148);
nor U813 (N_813,N_36,N_195);
or U814 (N_814,N_481,N_471);
nand U815 (N_815,N_260,N_295);
nand U816 (N_816,N_24,N_85);
nand U817 (N_817,N_436,N_211);
nor U818 (N_818,N_214,N_410);
xnor U819 (N_819,N_125,N_419);
nor U820 (N_820,N_67,N_229);
nand U821 (N_821,N_540,N_109);
nor U822 (N_822,N_142,N_7);
or U823 (N_823,N_439,N_132);
nor U824 (N_824,N_421,N_573);
nor U825 (N_825,N_72,N_6);
nand U826 (N_826,N_572,N_567);
or U827 (N_827,N_335,N_79);
and U828 (N_828,N_428,N_94);
and U829 (N_829,N_456,N_49);
and U830 (N_830,N_521,N_235);
and U831 (N_831,N_462,N_171);
or U832 (N_832,N_130,N_564);
nor U833 (N_833,N_119,N_489);
nor U834 (N_834,N_290,N_552);
nand U835 (N_835,N_241,N_501);
and U836 (N_836,N_576,N_447);
nand U837 (N_837,N_344,N_81);
and U838 (N_838,N_222,N_319);
nand U839 (N_839,N_162,N_367);
and U840 (N_840,N_353,N_14);
or U841 (N_841,N_284,N_116);
nor U842 (N_842,N_219,N_154);
and U843 (N_843,N_281,N_273);
nand U844 (N_844,N_528,N_65);
or U845 (N_845,N_430,N_98);
nor U846 (N_846,N_11,N_238);
and U847 (N_847,N_163,N_27);
nor U848 (N_848,N_336,N_33);
and U849 (N_849,N_479,N_360);
or U850 (N_850,N_483,N_278);
or U851 (N_851,N_313,N_305);
nand U852 (N_852,N_198,N_566);
or U853 (N_853,N_550,N_59);
nand U854 (N_854,N_111,N_422);
and U855 (N_855,N_253,N_533);
nand U856 (N_856,N_596,N_246);
or U857 (N_857,N_463,N_252);
and U858 (N_858,N_453,N_234);
and U859 (N_859,N_199,N_213);
or U860 (N_860,N_466,N_233);
nand U861 (N_861,N_398,N_173);
or U862 (N_862,N_486,N_160);
and U863 (N_863,N_355,N_557);
and U864 (N_864,N_164,N_117);
and U865 (N_865,N_401,N_22);
nor U866 (N_866,N_218,N_467);
or U867 (N_867,N_209,N_400);
or U868 (N_868,N_565,N_432);
or U869 (N_869,N_268,N_549);
nand U870 (N_870,N_553,N_45);
and U871 (N_871,N_506,N_133);
and U872 (N_872,N_138,N_84);
or U873 (N_873,N_554,N_590);
nand U874 (N_874,N_178,N_68);
nand U875 (N_875,N_127,N_189);
nor U876 (N_876,N_300,N_261);
nand U877 (N_877,N_356,N_91);
nand U878 (N_878,N_532,N_92);
and U879 (N_879,N_168,N_579);
xor U880 (N_880,N_89,N_310);
nor U881 (N_881,N_485,N_76);
nor U882 (N_882,N_514,N_316);
and U883 (N_883,N_575,N_88);
nor U884 (N_884,N_354,N_405);
and U885 (N_885,N_61,N_48);
and U886 (N_886,N_452,N_242);
or U887 (N_887,N_537,N_470);
nor U888 (N_888,N_524,N_270);
and U889 (N_889,N_587,N_69);
and U890 (N_890,N_556,N_368);
nand U891 (N_891,N_328,N_429);
or U892 (N_892,N_184,N_249);
nor U893 (N_893,N_17,N_474);
and U894 (N_894,N_546,N_362);
or U895 (N_895,N_517,N_106);
and U896 (N_896,N_101,N_393);
or U897 (N_897,N_208,N_435);
or U898 (N_898,N_348,N_440);
nand U899 (N_899,N_263,N_594);
or U900 (N_900,N_159,N_229);
and U901 (N_901,N_318,N_473);
or U902 (N_902,N_488,N_417);
nand U903 (N_903,N_511,N_150);
nor U904 (N_904,N_202,N_466);
nand U905 (N_905,N_63,N_495);
or U906 (N_906,N_193,N_427);
or U907 (N_907,N_312,N_187);
nand U908 (N_908,N_279,N_192);
nor U909 (N_909,N_381,N_70);
nor U910 (N_910,N_154,N_245);
nand U911 (N_911,N_484,N_269);
nor U912 (N_912,N_568,N_586);
nor U913 (N_913,N_319,N_499);
and U914 (N_914,N_424,N_73);
and U915 (N_915,N_24,N_556);
and U916 (N_916,N_29,N_393);
nor U917 (N_917,N_25,N_236);
nor U918 (N_918,N_599,N_363);
or U919 (N_919,N_167,N_556);
or U920 (N_920,N_15,N_576);
or U921 (N_921,N_220,N_361);
and U922 (N_922,N_50,N_31);
and U923 (N_923,N_492,N_388);
and U924 (N_924,N_183,N_140);
nand U925 (N_925,N_141,N_519);
or U926 (N_926,N_512,N_441);
nand U927 (N_927,N_352,N_11);
nor U928 (N_928,N_583,N_517);
or U929 (N_929,N_521,N_213);
nand U930 (N_930,N_487,N_87);
nor U931 (N_931,N_224,N_311);
nor U932 (N_932,N_106,N_416);
and U933 (N_933,N_53,N_73);
or U934 (N_934,N_50,N_569);
nand U935 (N_935,N_83,N_459);
nor U936 (N_936,N_599,N_47);
nor U937 (N_937,N_412,N_229);
or U938 (N_938,N_360,N_136);
nor U939 (N_939,N_473,N_538);
or U940 (N_940,N_520,N_456);
and U941 (N_941,N_323,N_254);
nand U942 (N_942,N_385,N_362);
or U943 (N_943,N_155,N_381);
nor U944 (N_944,N_467,N_128);
and U945 (N_945,N_314,N_303);
and U946 (N_946,N_540,N_260);
nand U947 (N_947,N_31,N_582);
and U948 (N_948,N_478,N_403);
nand U949 (N_949,N_132,N_174);
or U950 (N_950,N_438,N_301);
or U951 (N_951,N_31,N_12);
nor U952 (N_952,N_109,N_310);
or U953 (N_953,N_149,N_98);
nand U954 (N_954,N_405,N_182);
and U955 (N_955,N_17,N_385);
nand U956 (N_956,N_523,N_594);
or U957 (N_957,N_271,N_218);
nand U958 (N_958,N_209,N_499);
nand U959 (N_959,N_534,N_431);
nor U960 (N_960,N_215,N_64);
nand U961 (N_961,N_465,N_598);
nand U962 (N_962,N_496,N_454);
nor U963 (N_963,N_355,N_61);
nand U964 (N_964,N_253,N_135);
nor U965 (N_965,N_135,N_398);
or U966 (N_966,N_42,N_100);
nand U967 (N_967,N_290,N_129);
or U968 (N_968,N_241,N_296);
and U969 (N_969,N_466,N_593);
nor U970 (N_970,N_68,N_547);
nand U971 (N_971,N_433,N_133);
xor U972 (N_972,N_152,N_559);
nand U973 (N_973,N_387,N_355);
and U974 (N_974,N_472,N_6);
nand U975 (N_975,N_243,N_80);
nand U976 (N_976,N_16,N_275);
nand U977 (N_977,N_71,N_52);
nor U978 (N_978,N_500,N_281);
nand U979 (N_979,N_390,N_250);
nor U980 (N_980,N_207,N_123);
nand U981 (N_981,N_228,N_472);
nand U982 (N_982,N_149,N_59);
and U983 (N_983,N_180,N_494);
or U984 (N_984,N_112,N_364);
nand U985 (N_985,N_428,N_282);
or U986 (N_986,N_528,N_135);
nor U987 (N_987,N_62,N_120);
and U988 (N_988,N_574,N_21);
nand U989 (N_989,N_167,N_395);
nor U990 (N_990,N_422,N_454);
nand U991 (N_991,N_472,N_68);
and U992 (N_992,N_268,N_570);
nor U993 (N_993,N_595,N_25);
nor U994 (N_994,N_133,N_362);
nor U995 (N_995,N_220,N_91);
nor U996 (N_996,N_543,N_264);
nand U997 (N_997,N_213,N_413);
nand U998 (N_998,N_47,N_20);
nor U999 (N_999,N_417,N_497);
and U1000 (N_1000,N_369,N_256);
and U1001 (N_1001,N_333,N_492);
nand U1002 (N_1002,N_539,N_332);
nand U1003 (N_1003,N_103,N_318);
or U1004 (N_1004,N_344,N_291);
nor U1005 (N_1005,N_294,N_358);
nor U1006 (N_1006,N_180,N_433);
nand U1007 (N_1007,N_132,N_356);
nor U1008 (N_1008,N_179,N_525);
and U1009 (N_1009,N_586,N_267);
nor U1010 (N_1010,N_40,N_159);
nand U1011 (N_1011,N_275,N_487);
or U1012 (N_1012,N_430,N_55);
nand U1013 (N_1013,N_220,N_419);
or U1014 (N_1014,N_253,N_158);
nand U1015 (N_1015,N_63,N_590);
nor U1016 (N_1016,N_60,N_492);
or U1017 (N_1017,N_63,N_88);
nand U1018 (N_1018,N_294,N_482);
nand U1019 (N_1019,N_447,N_343);
and U1020 (N_1020,N_137,N_212);
or U1021 (N_1021,N_272,N_253);
nor U1022 (N_1022,N_512,N_308);
nor U1023 (N_1023,N_555,N_32);
and U1024 (N_1024,N_394,N_78);
and U1025 (N_1025,N_193,N_278);
nand U1026 (N_1026,N_90,N_402);
nor U1027 (N_1027,N_528,N_491);
and U1028 (N_1028,N_58,N_63);
nand U1029 (N_1029,N_459,N_12);
or U1030 (N_1030,N_46,N_38);
nor U1031 (N_1031,N_175,N_180);
or U1032 (N_1032,N_265,N_34);
and U1033 (N_1033,N_382,N_517);
nor U1034 (N_1034,N_303,N_123);
or U1035 (N_1035,N_447,N_325);
or U1036 (N_1036,N_136,N_561);
nand U1037 (N_1037,N_202,N_331);
nor U1038 (N_1038,N_452,N_431);
and U1039 (N_1039,N_407,N_536);
nand U1040 (N_1040,N_146,N_560);
and U1041 (N_1041,N_278,N_57);
and U1042 (N_1042,N_377,N_160);
nand U1043 (N_1043,N_277,N_337);
nand U1044 (N_1044,N_447,N_544);
nand U1045 (N_1045,N_448,N_391);
nand U1046 (N_1046,N_108,N_457);
nor U1047 (N_1047,N_2,N_479);
or U1048 (N_1048,N_57,N_529);
or U1049 (N_1049,N_200,N_332);
nand U1050 (N_1050,N_65,N_576);
or U1051 (N_1051,N_238,N_203);
or U1052 (N_1052,N_150,N_43);
nor U1053 (N_1053,N_467,N_280);
nand U1054 (N_1054,N_227,N_265);
and U1055 (N_1055,N_399,N_6);
nand U1056 (N_1056,N_313,N_423);
or U1057 (N_1057,N_21,N_529);
nand U1058 (N_1058,N_454,N_433);
nand U1059 (N_1059,N_553,N_33);
and U1060 (N_1060,N_350,N_587);
or U1061 (N_1061,N_522,N_153);
nor U1062 (N_1062,N_341,N_420);
xor U1063 (N_1063,N_5,N_108);
or U1064 (N_1064,N_407,N_544);
nand U1065 (N_1065,N_534,N_497);
or U1066 (N_1066,N_449,N_423);
nand U1067 (N_1067,N_561,N_506);
nand U1068 (N_1068,N_507,N_27);
nand U1069 (N_1069,N_549,N_148);
or U1070 (N_1070,N_47,N_5);
and U1071 (N_1071,N_92,N_328);
nand U1072 (N_1072,N_416,N_585);
or U1073 (N_1073,N_464,N_6);
or U1074 (N_1074,N_246,N_305);
nand U1075 (N_1075,N_317,N_441);
nor U1076 (N_1076,N_477,N_78);
and U1077 (N_1077,N_252,N_574);
nand U1078 (N_1078,N_515,N_115);
or U1079 (N_1079,N_368,N_399);
nor U1080 (N_1080,N_313,N_37);
nand U1081 (N_1081,N_188,N_50);
and U1082 (N_1082,N_32,N_218);
nand U1083 (N_1083,N_120,N_379);
xnor U1084 (N_1084,N_276,N_578);
and U1085 (N_1085,N_394,N_178);
nand U1086 (N_1086,N_516,N_412);
and U1087 (N_1087,N_292,N_90);
xor U1088 (N_1088,N_235,N_582);
nor U1089 (N_1089,N_525,N_171);
nor U1090 (N_1090,N_441,N_274);
nand U1091 (N_1091,N_357,N_106);
or U1092 (N_1092,N_519,N_153);
nand U1093 (N_1093,N_318,N_388);
and U1094 (N_1094,N_1,N_167);
nand U1095 (N_1095,N_110,N_509);
nor U1096 (N_1096,N_218,N_373);
nand U1097 (N_1097,N_428,N_589);
nor U1098 (N_1098,N_367,N_60);
or U1099 (N_1099,N_450,N_147);
and U1100 (N_1100,N_94,N_141);
or U1101 (N_1101,N_189,N_526);
and U1102 (N_1102,N_442,N_151);
or U1103 (N_1103,N_33,N_288);
nand U1104 (N_1104,N_429,N_282);
or U1105 (N_1105,N_353,N_336);
or U1106 (N_1106,N_72,N_181);
nand U1107 (N_1107,N_379,N_449);
nor U1108 (N_1108,N_231,N_35);
nor U1109 (N_1109,N_588,N_257);
nand U1110 (N_1110,N_505,N_441);
nand U1111 (N_1111,N_442,N_389);
and U1112 (N_1112,N_131,N_454);
and U1113 (N_1113,N_246,N_156);
nor U1114 (N_1114,N_386,N_265);
or U1115 (N_1115,N_536,N_209);
nand U1116 (N_1116,N_51,N_446);
and U1117 (N_1117,N_329,N_407);
or U1118 (N_1118,N_506,N_20);
and U1119 (N_1119,N_504,N_448);
nand U1120 (N_1120,N_324,N_452);
and U1121 (N_1121,N_462,N_197);
and U1122 (N_1122,N_61,N_14);
nand U1123 (N_1123,N_374,N_489);
nor U1124 (N_1124,N_56,N_595);
or U1125 (N_1125,N_373,N_158);
nand U1126 (N_1126,N_507,N_324);
nand U1127 (N_1127,N_495,N_5);
nor U1128 (N_1128,N_231,N_448);
nor U1129 (N_1129,N_59,N_576);
nor U1130 (N_1130,N_27,N_212);
nand U1131 (N_1131,N_440,N_512);
nand U1132 (N_1132,N_483,N_290);
nand U1133 (N_1133,N_204,N_284);
nand U1134 (N_1134,N_184,N_591);
nand U1135 (N_1135,N_190,N_176);
nor U1136 (N_1136,N_47,N_364);
and U1137 (N_1137,N_164,N_570);
nor U1138 (N_1138,N_295,N_551);
nand U1139 (N_1139,N_138,N_178);
or U1140 (N_1140,N_313,N_55);
and U1141 (N_1141,N_350,N_122);
nor U1142 (N_1142,N_214,N_330);
nand U1143 (N_1143,N_69,N_374);
nand U1144 (N_1144,N_531,N_517);
or U1145 (N_1145,N_171,N_146);
and U1146 (N_1146,N_89,N_172);
nand U1147 (N_1147,N_575,N_250);
nand U1148 (N_1148,N_243,N_23);
nor U1149 (N_1149,N_547,N_390);
nor U1150 (N_1150,N_443,N_285);
nor U1151 (N_1151,N_407,N_98);
nor U1152 (N_1152,N_431,N_539);
nand U1153 (N_1153,N_486,N_380);
and U1154 (N_1154,N_555,N_558);
or U1155 (N_1155,N_24,N_400);
nand U1156 (N_1156,N_520,N_455);
nand U1157 (N_1157,N_226,N_175);
nor U1158 (N_1158,N_273,N_171);
nand U1159 (N_1159,N_313,N_511);
nor U1160 (N_1160,N_532,N_16);
nor U1161 (N_1161,N_60,N_496);
and U1162 (N_1162,N_271,N_176);
nand U1163 (N_1163,N_9,N_556);
and U1164 (N_1164,N_503,N_585);
nand U1165 (N_1165,N_210,N_525);
or U1166 (N_1166,N_479,N_588);
nand U1167 (N_1167,N_137,N_88);
nand U1168 (N_1168,N_9,N_306);
or U1169 (N_1169,N_279,N_280);
nand U1170 (N_1170,N_52,N_410);
and U1171 (N_1171,N_299,N_240);
or U1172 (N_1172,N_188,N_455);
nor U1173 (N_1173,N_496,N_353);
nor U1174 (N_1174,N_427,N_575);
and U1175 (N_1175,N_237,N_29);
xor U1176 (N_1176,N_213,N_550);
nand U1177 (N_1177,N_199,N_179);
nor U1178 (N_1178,N_359,N_446);
nand U1179 (N_1179,N_274,N_348);
or U1180 (N_1180,N_115,N_471);
nor U1181 (N_1181,N_210,N_215);
or U1182 (N_1182,N_465,N_34);
nand U1183 (N_1183,N_17,N_75);
nand U1184 (N_1184,N_173,N_472);
or U1185 (N_1185,N_235,N_380);
nand U1186 (N_1186,N_310,N_201);
nor U1187 (N_1187,N_514,N_203);
nor U1188 (N_1188,N_159,N_282);
or U1189 (N_1189,N_345,N_521);
nor U1190 (N_1190,N_539,N_368);
and U1191 (N_1191,N_231,N_590);
and U1192 (N_1192,N_443,N_305);
nand U1193 (N_1193,N_345,N_384);
and U1194 (N_1194,N_279,N_564);
or U1195 (N_1195,N_524,N_520);
nand U1196 (N_1196,N_580,N_443);
nand U1197 (N_1197,N_122,N_93);
and U1198 (N_1198,N_213,N_207);
or U1199 (N_1199,N_409,N_355);
nor U1200 (N_1200,N_790,N_1138);
or U1201 (N_1201,N_931,N_1086);
nor U1202 (N_1202,N_1172,N_627);
or U1203 (N_1203,N_610,N_1165);
and U1204 (N_1204,N_1179,N_1170);
or U1205 (N_1205,N_1129,N_794);
nor U1206 (N_1206,N_1033,N_1014);
nand U1207 (N_1207,N_1122,N_999);
nand U1208 (N_1208,N_1015,N_967);
and U1209 (N_1209,N_924,N_890);
nor U1210 (N_1210,N_1012,N_944);
nor U1211 (N_1211,N_1114,N_653);
xor U1212 (N_1212,N_1069,N_756);
nand U1213 (N_1213,N_1175,N_664);
and U1214 (N_1214,N_938,N_806);
nand U1215 (N_1215,N_1188,N_702);
or U1216 (N_1216,N_1112,N_761);
and U1217 (N_1217,N_1037,N_830);
and U1218 (N_1218,N_780,N_824);
nor U1219 (N_1219,N_1124,N_1159);
nand U1220 (N_1220,N_691,N_1091);
and U1221 (N_1221,N_991,N_1022);
and U1222 (N_1222,N_990,N_1008);
or U1223 (N_1223,N_766,N_833);
nand U1224 (N_1224,N_636,N_720);
and U1225 (N_1225,N_838,N_963);
nor U1226 (N_1226,N_689,N_869);
and U1227 (N_1227,N_718,N_1043);
nor U1228 (N_1228,N_867,N_704);
nor U1229 (N_1229,N_905,N_776);
nor U1230 (N_1230,N_850,N_839);
nand U1231 (N_1231,N_980,N_754);
nand U1232 (N_1232,N_827,N_863);
nand U1233 (N_1233,N_645,N_868);
and U1234 (N_1234,N_670,N_799);
nand U1235 (N_1235,N_1173,N_1117);
nand U1236 (N_1236,N_940,N_741);
or U1237 (N_1237,N_1155,N_1064);
nor U1238 (N_1238,N_742,N_947);
and U1239 (N_1239,N_625,N_860);
nor U1240 (N_1240,N_744,N_1081);
nand U1241 (N_1241,N_1152,N_675);
or U1242 (N_1242,N_1062,N_1157);
xnor U1243 (N_1243,N_1177,N_774);
or U1244 (N_1244,N_1142,N_994);
and U1245 (N_1245,N_810,N_1098);
and U1246 (N_1246,N_783,N_808);
nand U1247 (N_1247,N_1192,N_713);
nand U1248 (N_1248,N_1058,N_881);
and U1249 (N_1249,N_976,N_677);
nand U1250 (N_1250,N_886,N_1007);
and U1251 (N_1251,N_604,N_851);
and U1252 (N_1252,N_845,N_921);
and U1253 (N_1253,N_1006,N_601);
nor U1254 (N_1254,N_753,N_727);
and U1255 (N_1255,N_646,N_656);
and U1256 (N_1256,N_789,N_688);
nand U1257 (N_1257,N_1001,N_832);
nor U1258 (N_1258,N_730,N_858);
nand U1259 (N_1259,N_966,N_1083);
and U1260 (N_1260,N_866,N_920);
and U1261 (N_1261,N_820,N_695);
nor U1262 (N_1262,N_1195,N_989);
nor U1263 (N_1263,N_975,N_913);
nor U1264 (N_1264,N_731,N_849);
or U1265 (N_1265,N_823,N_1130);
or U1266 (N_1266,N_979,N_1139);
and U1267 (N_1267,N_805,N_1029);
or U1268 (N_1268,N_1049,N_891);
or U1269 (N_1269,N_888,N_935);
and U1270 (N_1270,N_884,N_1054);
or U1271 (N_1271,N_958,N_919);
nand U1272 (N_1272,N_1087,N_959);
or U1273 (N_1273,N_781,N_791);
and U1274 (N_1274,N_986,N_1032);
or U1275 (N_1275,N_611,N_708);
or U1276 (N_1276,N_729,N_1031);
or U1277 (N_1277,N_750,N_747);
nor U1278 (N_1278,N_767,N_1044);
nand U1279 (N_1279,N_1010,N_1090);
or U1280 (N_1280,N_942,N_1060);
and U1281 (N_1281,N_1168,N_894);
nand U1282 (N_1282,N_1002,N_1028);
or U1283 (N_1283,N_900,N_957);
nor U1284 (N_1284,N_927,N_1063);
and U1285 (N_1285,N_714,N_904);
and U1286 (N_1286,N_972,N_1180);
and U1287 (N_1287,N_711,N_658);
or U1288 (N_1288,N_875,N_1061);
and U1289 (N_1289,N_661,N_1103);
nand U1290 (N_1290,N_1095,N_1106);
nand U1291 (N_1291,N_1017,N_985);
nor U1292 (N_1292,N_686,N_666);
nand U1293 (N_1293,N_786,N_699);
nand U1294 (N_1294,N_1126,N_950);
and U1295 (N_1295,N_871,N_968);
nor U1296 (N_1296,N_671,N_1038);
nor U1297 (N_1297,N_949,N_692);
or U1298 (N_1298,N_971,N_922);
and U1299 (N_1299,N_1111,N_630);
and U1300 (N_1300,N_628,N_952);
nand U1301 (N_1301,N_1162,N_1199);
or U1302 (N_1302,N_848,N_1068);
nor U1303 (N_1303,N_1020,N_910);
nor U1304 (N_1304,N_615,N_911);
nor U1305 (N_1305,N_1026,N_917);
and U1306 (N_1306,N_1134,N_703);
or U1307 (N_1307,N_934,N_733);
nor U1308 (N_1308,N_898,N_746);
nor U1309 (N_1309,N_1097,N_901);
xor U1310 (N_1310,N_983,N_1019);
nor U1311 (N_1311,N_758,N_614);
nor U1312 (N_1312,N_1151,N_698);
and U1313 (N_1313,N_785,N_1074);
nand U1314 (N_1314,N_822,N_690);
or U1315 (N_1315,N_914,N_1133);
and U1316 (N_1316,N_728,N_801);
and U1317 (N_1317,N_1071,N_640);
or U1318 (N_1318,N_1181,N_889);
or U1319 (N_1319,N_651,N_973);
nand U1320 (N_1320,N_1041,N_620);
nor U1321 (N_1321,N_907,N_932);
nor U1322 (N_1322,N_1148,N_676);
nor U1323 (N_1323,N_1137,N_723);
nand U1324 (N_1324,N_1153,N_1070);
and U1325 (N_1325,N_1120,N_683);
nor U1326 (N_1326,N_685,N_826);
nor U1327 (N_1327,N_795,N_996);
nand U1328 (N_1328,N_897,N_831);
and U1329 (N_1329,N_769,N_792);
or U1330 (N_1330,N_841,N_607);
nand U1331 (N_1331,N_709,N_879);
nor U1332 (N_1332,N_1140,N_796);
nor U1333 (N_1333,N_751,N_648);
nand U1334 (N_1334,N_853,N_818);
and U1335 (N_1335,N_925,N_998);
and U1336 (N_1336,N_768,N_665);
and U1337 (N_1337,N_837,N_700);
or U1338 (N_1338,N_735,N_1166);
or U1339 (N_1339,N_825,N_748);
nand U1340 (N_1340,N_842,N_1055);
or U1341 (N_1341,N_1123,N_779);
and U1342 (N_1342,N_715,N_777);
or U1343 (N_1343,N_762,N_1089);
nor U1344 (N_1344,N_908,N_1040);
or U1345 (N_1345,N_814,N_1021);
and U1346 (N_1346,N_1005,N_946);
nand U1347 (N_1347,N_1036,N_701);
nand U1348 (N_1348,N_706,N_1144);
nor U1349 (N_1349,N_765,N_621);
or U1350 (N_1350,N_637,N_643);
nand U1351 (N_1351,N_679,N_608);
nand U1352 (N_1352,N_918,N_693);
nor U1353 (N_1353,N_668,N_684);
nor U1354 (N_1354,N_1161,N_811);
nand U1355 (N_1355,N_835,N_784);
nor U1356 (N_1356,N_836,N_902);
or U1357 (N_1357,N_803,N_923);
and U1358 (N_1358,N_895,N_961);
nor U1359 (N_1359,N_719,N_1059);
or U1360 (N_1360,N_778,N_1102);
nand U1361 (N_1361,N_770,N_997);
or U1362 (N_1362,N_821,N_864);
nand U1363 (N_1363,N_609,N_1025);
and U1364 (N_1364,N_1051,N_605);
nor U1365 (N_1365,N_834,N_816);
nor U1366 (N_1366,N_1131,N_667);
nor U1367 (N_1367,N_1065,N_1024);
and U1368 (N_1368,N_846,N_1187);
or U1369 (N_1369,N_672,N_882);
nor U1370 (N_1370,N_612,N_1141);
nor U1371 (N_1371,N_793,N_752);
nor U1372 (N_1372,N_945,N_1035);
or U1373 (N_1373,N_981,N_697);
nand U1374 (N_1374,N_788,N_885);
and U1375 (N_1375,N_1034,N_616);
and U1376 (N_1376,N_617,N_1185);
nand U1377 (N_1377,N_862,N_937);
nand U1378 (N_1378,N_639,N_856);
and U1379 (N_1379,N_1013,N_844);
nand U1380 (N_1380,N_716,N_797);
and U1381 (N_1381,N_737,N_1009);
and U1382 (N_1382,N_1108,N_1000);
nor U1383 (N_1383,N_1042,N_798);
nand U1384 (N_1384,N_1105,N_988);
nor U1385 (N_1385,N_887,N_1132);
or U1386 (N_1386,N_977,N_1136);
or U1387 (N_1387,N_962,N_1183);
nor U1388 (N_1388,N_1078,N_1077);
nand U1389 (N_1389,N_644,N_600);
xor U1390 (N_1390,N_1154,N_1030);
and U1391 (N_1391,N_1115,N_915);
or U1392 (N_1392,N_843,N_1109);
or U1393 (N_1393,N_722,N_1169);
nor U1394 (N_1394,N_712,N_1128);
or U1395 (N_1395,N_650,N_987);
or U1396 (N_1396,N_876,N_682);
nand U1397 (N_1397,N_802,N_909);
or U1398 (N_1398,N_936,N_773);
nand U1399 (N_1399,N_1027,N_807);
or U1400 (N_1400,N_1079,N_1048);
nand U1401 (N_1401,N_1150,N_1149);
nor U1402 (N_1402,N_655,N_1056);
and U1403 (N_1403,N_1096,N_1039);
and U1404 (N_1404,N_948,N_1127);
or U1405 (N_1405,N_970,N_1164);
or U1406 (N_1406,N_622,N_1085);
nor U1407 (N_1407,N_943,N_854);
and U1408 (N_1408,N_649,N_1178);
and U1409 (N_1409,N_1046,N_726);
nand U1410 (N_1410,N_982,N_662);
nor U1411 (N_1411,N_926,N_775);
nor U1412 (N_1412,N_960,N_1092);
or U1413 (N_1413,N_642,N_740);
nor U1414 (N_1414,N_1125,N_1072);
and U1415 (N_1415,N_883,N_1163);
and U1416 (N_1416,N_893,N_828);
nor U1417 (N_1417,N_707,N_694);
nand U1418 (N_1418,N_725,N_1082);
or U1419 (N_1419,N_732,N_857);
or U1420 (N_1420,N_1107,N_659);
nor U1421 (N_1421,N_603,N_1099);
nand U1422 (N_1422,N_1057,N_1093);
nor U1423 (N_1423,N_995,N_1076);
nor U1424 (N_1424,N_1182,N_652);
or U1425 (N_1425,N_657,N_638);
nand U1426 (N_1426,N_631,N_852);
or U1427 (N_1427,N_634,N_1003);
or U1428 (N_1428,N_772,N_829);
or U1429 (N_1429,N_1135,N_955);
nor U1430 (N_1430,N_1101,N_847);
nor U1431 (N_1431,N_1053,N_984);
and U1432 (N_1432,N_606,N_929);
and U1433 (N_1433,N_1146,N_618);
nand U1434 (N_1434,N_1160,N_1047);
nand U1435 (N_1435,N_759,N_1104);
nand U1436 (N_1436,N_1156,N_1176);
or U1437 (N_1437,N_757,N_1186);
nor U1438 (N_1438,N_1066,N_755);
nand U1439 (N_1439,N_749,N_1045);
and U1440 (N_1440,N_1158,N_877);
or U1441 (N_1441,N_1080,N_654);
and U1442 (N_1442,N_930,N_705);
and U1443 (N_1443,N_632,N_928);
and U1444 (N_1444,N_1073,N_771);
or U1445 (N_1445,N_1191,N_993);
or U1446 (N_1446,N_964,N_965);
or U1447 (N_1447,N_1004,N_1094);
nand U1448 (N_1448,N_1075,N_602);
nor U1449 (N_1449,N_855,N_724);
and U1450 (N_1450,N_1147,N_669);
and U1451 (N_1451,N_870,N_912);
or U1452 (N_1452,N_1088,N_1100);
xnor U1453 (N_1453,N_969,N_819);
nor U1454 (N_1454,N_673,N_1143);
and U1455 (N_1455,N_680,N_872);
or U1456 (N_1456,N_933,N_978);
nor U1457 (N_1457,N_717,N_681);
and U1458 (N_1458,N_1190,N_626);
nand U1459 (N_1459,N_1011,N_782);
and U1460 (N_1460,N_1145,N_629);
nand U1461 (N_1461,N_1196,N_941);
and U1462 (N_1462,N_635,N_764);
nand U1463 (N_1463,N_1110,N_1016);
nand U1464 (N_1464,N_939,N_906);
nor U1465 (N_1465,N_840,N_809);
and U1466 (N_1466,N_951,N_1174);
and U1467 (N_1467,N_800,N_1121);
nor U1468 (N_1468,N_787,N_1113);
nor U1469 (N_1469,N_745,N_1116);
and U1470 (N_1470,N_1189,N_641);
and U1471 (N_1471,N_1067,N_956);
and U1472 (N_1472,N_1023,N_1018);
and U1473 (N_1473,N_743,N_663);
nand U1474 (N_1474,N_624,N_1084);
nand U1475 (N_1475,N_734,N_903);
nand U1476 (N_1476,N_804,N_815);
nor U1477 (N_1477,N_739,N_623);
and U1478 (N_1478,N_1119,N_1184);
and U1479 (N_1479,N_1050,N_1167);
nor U1480 (N_1480,N_721,N_710);
and U1481 (N_1481,N_916,N_880);
nand U1482 (N_1482,N_992,N_760);
nand U1483 (N_1483,N_660,N_861);
nand U1484 (N_1484,N_687,N_678);
or U1485 (N_1485,N_736,N_896);
nor U1486 (N_1486,N_1171,N_1118);
and U1487 (N_1487,N_674,N_874);
and U1488 (N_1488,N_812,N_899);
nand U1489 (N_1489,N_859,N_1197);
or U1490 (N_1490,N_865,N_974);
or U1491 (N_1491,N_953,N_1052);
or U1492 (N_1492,N_1193,N_878);
nand U1493 (N_1493,N_892,N_613);
or U1494 (N_1494,N_696,N_954);
or U1495 (N_1495,N_763,N_1198);
or U1496 (N_1496,N_738,N_1194);
and U1497 (N_1497,N_817,N_633);
and U1498 (N_1498,N_619,N_813);
and U1499 (N_1499,N_647,N_873);
nand U1500 (N_1500,N_1120,N_983);
nand U1501 (N_1501,N_753,N_1158);
and U1502 (N_1502,N_802,N_1087);
nand U1503 (N_1503,N_605,N_677);
nand U1504 (N_1504,N_763,N_767);
or U1505 (N_1505,N_747,N_786);
nand U1506 (N_1506,N_1107,N_861);
nor U1507 (N_1507,N_1192,N_1144);
and U1508 (N_1508,N_1136,N_1151);
or U1509 (N_1509,N_1125,N_1183);
and U1510 (N_1510,N_633,N_1042);
or U1511 (N_1511,N_814,N_1076);
and U1512 (N_1512,N_824,N_751);
nor U1513 (N_1513,N_1080,N_1166);
or U1514 (N_1514,N_962,N_832);
or U1515 (N_1515,N_888,N_1123);
nor U1516 (N_1516,N_816,N_860);
nor U1517 (N_1517,N_1004,N_995);
nor U1518 (N_1518,N_616,N_872);
nor U1519 (N_1519,N_982,N_884);
nor U1520 (N_1520,N_1024,N_1029);
and U1521 (N_1521,N_632,N_1121);
and U1522 (N_1522,N_1066,N_972);
nand U1523 (N_1523,N_1157,N_1091);
or U1524 (N_1524,N_885,N_980);
or U1525 (N_1525,N_1015,N_877);
nor U1526 (N_1526,N_792,N_607);
and U1527 (N_1527,N_796,N_1015);
nor U1528 (N_1528,N_1117,N_1090);
nor U1529 (N_1529,N_663,N_1130);
nor U1530 (N_1530,N_1162,N_905);
nand U1531 (N_1531,N_1066,N_1170);
and U1532 (N_1532,N_780,N_929);
nand U1533 (N_1533,N_1149,N_1018);
and U1534 (N_1534,N_1036,N_883);
and U1535 (N_1535,N_865,N_656);
nor U1536 (N_1536,N_735,N_805);
nor U1537 (N_1537,N_1056,N_904);
nand U1538 (N_1538,N_1053,N_1047);
and U1539 (N_1539,N_1028,N_1058);
and U1540 (N_1540,N_703,N_810);
or U1541 (N_1541,N_721,N_1040);
and U1542 (N_1542,N_1006,N_916);
nor U1543 (N_1543,N_777,N_830);
and U1544 (N_1544,N_1159,N_953);
nand U1545 (N_1545,N_902,N_768);
nor U1546 (N_1546,N_837,N_1001);
or U1547 (N_1547,N_603,N_668);
and U1548 (N_1548,N_1167,N_728);
nand U1549 (N_1549,N_681,N_602);
and U1550 (N_1550,N_1109,N_1066);
and U1551 (N_1551,N_683,N_1068);
nand U1552 (N_1552,N_973,N_914);
or U1553 (N_1553,N_1173,N_1084);
nor U1554 (N_1554,N_626,N_878);
nand U1555 (N_1555,N_830,N_989);
nor U1556 (N_1556,N_656,N_929);
nand U1557 (N_1557,N_1096,N_660);
nor U1558 (N_1558,N_1020,N_842);
nand U1559 (N_1559,N_1034,N_666);
nand U1560 (N_1560,N_719,N_811);
or U1561 (N_1561,N_910,N_798);
and U1562 (N_1562,N_971,N_1121);
nand U1563 (N_1563,N_946,N_970);
nand U1564 (N_1564,N_871,N_1099);
nand U1565 (N_1565,N_1144,N_796);
or U1566 (N_1566,N_812,N_963);
and U1567 (N_1567,N_691,N_1032);
and U1568 (N_1568,N_607,N_954);
and U1569 (N_1569,N_662,N_1170);
and U1570 (N_1570,N_795,N_1050);
or U1571 (N_1571,N_852,N_681);
nand U1572 (N_1572,N_933,N_690);
nor U1573 (N_1573,N_612,N_875);
nor U1574 (N_1574,N_1028,N_1186);
and U1575 (N_1575,N_656,N_1000);
and U1576 (N_1576,N_801,N_883);
and U1577 (N_1577,N_615,N_764);
nand U1578 (N_1578,N_904,N_647);
or U1579 (N_1579,N_1004,N_1070);
nand U1580 (N_1580,N_738,N_763);
nand U1581 (N_1581,N_823,N_1153);
or U1582 (N_1582,N_1026,N_865);
nor U1583 (N_1583,N_705,N_791);
nand U1584 (N_1584,N_626,N_918);
and U1585 (N_1585,N_835,N_644);
and U1586 (N_1586,N_979,N_850);
nor U1587 (N_1587,N_780,N_620);
or U1588 (N_1588,N_951,N_709);
nor U1589 (N_1589,N_856,N_806);
and U1590 (N_1590,N_1191,N_714);
nand U1591 (N_1591,N_941,N_617);
or U1592 (N_1592,N_1157,N_869);
nand U1593 (N_1593,N_676,N_666);
nor U1594 (N_1594,N_1055,N_609);
and U1595 (N_1595,N_914,N_613);
nor U1596 (N_1596,N_877,N_1188);
nand U1597 (N_1597,N_683,N_609);
or U1598 (N_1598,N_772,N_817);
nor U1599 (N_1599,N_1094,N_985);
and U1600 (N_1600,N_885,N_1032);
nand U1601 (N_1601,N_1073,N_652);
nand U1602 (N_1602,N_979,N_744);
nor U1603 (N_1603,N_843,N_883);
or U1604 (N_1604,N_1169,N_1006);
and U1605 (N_1605,N_615,N_612);
nand U1606 (N_1606,N_1075,N_634);
nand U1607 (N_1607,N_612,N_882);
nand U1608 (N_1608,N_933,N_1130);
nand U1609 (N_1609,N_969,N_772);
nand U1610 (N_1610,N_989,N_1170);
nand U1611 (N_1611,N_886,N_1006);
or U1612 (N_1612,N_859,N_643);
or U1613 (N_1613,N_1045,N_621);
nand U1614 (N_1614,N_1116,N_824);
or U1615 (N_1615,N_854,N_1158);
nor U1616 (N_1616,N_691,N_645);
xor U1617 (N_1617,N_1017,N_660);
and U1618 (N_1618,N_786,N_1195);
nand U1619 (N_1619,N_1055,N_601);
nor U1620 (N_1620,N_680,N_813);
nor U1621 (N_1621,N_1006,N_955);
and U1622 (N_1622,N_793,N_686);
nand U1623 (N_1623,N_851,N_1033);
nand U1624 (N_1624,N_828,N_1138);
xor U1625 (N_1625,N_689,N_931);
and U1626 (N_1626,N_956,N_1084);
nor U1627 (N_1627,N_1175,N_727);
nor U1628 (N_1628,N_1128,N_1161);
nand U1629 (N_1629,N_872,N_621);
and U1630 (N_1630,N_800,N_1019);
nor U1631 (N_1631,N_758,N_1159);
nor U1632 (N_1632,N_949,N_871);
nand U1633 (N_1633,N_1182,N_980);
or U1634 (N_1634,N_998,N_991);
and U1635 (N_1635,N_961,N_1185);
and U1636 (N_1636,N_751,N_833);
or U1637 (N_1637,N_952,N_834);
or U1638 (N_1638,N_642,N_1171);
nand U1639 (N_1639,N_726,N_1164);
and U1640 (N_1640,N_1092,N_1126);
and U1641 (N_1641,N_1081,N_862);
nand U1642 (N_1642,N_703,N_731);
and U1643 (N_1643,N_1085,N_881);
and U1644 (N_1644,N_814,N_601);
and U1645 (N_1645,N_776,N_685);
or U1646 (N_1646,N_1169,N_985);
and U1647 (N_1647,N_947,N_1000);
or U1648 (N_1648,N_1126,N_653);
nand U1649 (N_1649,N_886,N_746);
nor U1650 (N_1650,N_843,N_1182);
nand U1651 (N_1651,N_1124,N_1183);
nor U1652 (N_1652,N_627,N_755);
or U1653 (N_1653,N_998,N_658);
nand U1654 (N_1654,N_1057,N_1096);
or U1655 (N_1655,N_689,N_751);
nor U1656 (N_1656,N_1187,N_769);
and U1657 (N_1657,N_1177,N_1014);
nor U1658 (N_1658,N_1003,N_735);
nor U1659 (N_1659,N_784,N_746);
or U1660 (N_1660,N_830,N_945);
nor U1661 (N_1661,N_1057,N_774);
nand U1662 (N_1662,N_702,N_1128);
and U1663 (N_1663,N_1010,N_883);
and U1664 (N_1664,N_929,N_626);
nand U1665 (N_1665,N_637,N_777);
nor U1666 (N_1666,N_1195,N_1067);
or U1667 (N_1667,N_636,N_925);
nor U1668 (N_1668,N_630,N_894);
nor U1669 (N_1669,N_1153,N_1036);
nand U1670 (N_1670,N_886,N_1092);
and U1671 (N_1671,N_1054,N_1019);
nor U1672 (N_1672,N_1155,N_1020);
nand U1673 (N_1673,N_858,N_1039);
and U1674 (N_1674,N_1185,N_1051);
and U1675 (N_1675,N_909,N_1056);
and U1676 (N_1676,N_720,N_1105);
and U1677 (N_1677,N_864,N_774);
or U1678 (N_1678,N_782,N_868);
nor U1679 (N_1679,N_863,N_687);
or U1680 (N_1680,N_1064,N_861);
or U1681 (N_1681,N_1066,N_603);
nand U1682 (N_1682,N_913,N_760);
or U1683 (N_1683,N_1175,N_875);
or U1684 (N_1684,N_901,N_804);
nor U1685 (N_1685,N_638,N_631);
and U1686 (N_1686,N_743,N_635);
or U1687 (N_1687,N_1150,N_880);
nor U1688 (N_1688,N_778,N_623);
nor U1689 (N_1689,N_723,N_1096);
nor U1690 (N_1690,N_614,N_980);
and U1691 (N_1691,N_672,N_630);
nand U1692 (N_1692,N_684,N_718);
and U1693 (N_1693,N_1084,N_605);
and U1694 (N_1694,N_913,N_1197);
or U1695 (N_1695,N_883,N_1064);
or U1696 (N_1696,N_782,N_947);
and U1697 (N_1697,N_608,N_736);
or U1698 (N_1698,N_722,N_841);
or U1699 (N_1699,N_1141,N_913);
nand U1700 (N_1700,N_1189,N_1107);
or U1701 (N_1701,N_1104,N_1145);
nand U1702 (N_1702,N_1122,N_736);
nand U1703 (N_1703,N_760,N_966);
or U1704 (N_1704,N_1076,N_917);
nor U1705 (N_1705,N_1057,N_793);
nand U1706 (N_1706,N_711,N_731);
nor U1707 (N_1707,N_1083,N_1024);
or U1708 (N_1708,N_681,N_776);
nand U1709 (N_1709,N_758,N_785);
nand U1710 (N_1710,N_631,N_1099);
nand U1711 (N_1711,N_646,N_753);
and U1712 (N_1712,N_683,N_996);
nor U1713 (N_1713,N_700,N_611);
nand U1714 (N_1714,N_680,N_1123);
or U1715 (N_1715,N_1150,N_771);
and U1716 (N_1716,N_726,N_900);
nand U1717 (N_1717,N_1186,N_1075);
or U1718 (N_1718,N_939,N_1011);
and U1719 (N_1719,N_943,N_1167);
nand U1720 (N_1720,N_782,N_718);
nand U1721 (N_1721,N_1085,N_1127);
or U1722 (N_1722,N_712,N_1073);
nor U1723 (N_1723,N_694,N_926);
nor U1724 (N_1724,N_1109,N_939);
nand U1725 (N_1725,N_1118,N_776);
or U1726 (N_1726,N_680,N_1079);
nand U1727 (N_1727,N_841,N_1085);
nand U1728 (N_1728,N_922,N_1018);
and U1729 (N_1729,N_1122,N_973);
nand U1730 (N_1730,N_642,N_1146);
nand U1731 (N_1731,N_1042,N_810);
and U1732 (N_1732,N_856,N_1040);
or U1733 (N_1733,N_736,N_789);
and U1734 (N_1734,N_735,N_1194);
nand U1735 (N_1735,N_951,N_1137);
nor U1736 (N_1736,N_1084,N_803);
nor U1737 (N_1737,N_1197,N_819);
or U1738 (N_1738,N_782,N_1147);
and U1739 (N_1739,N_840,N_1002);
nand U1740 (N_1740,N_680,N_906);
nor U1741 (N_1741,N_937,N_1156);
and U1742 (N_1742,N_607,N_832);
and U1743 (N_1743,N_899,N_982);
and U1744 (N_1744,N_763,N_871);
nand U1745 (N_1745,N_787,N_1064);
or U1746 (N_1746,N_648,N_1106);
and U1747 (N_1747,N_714,N_1086);
or U1748 (N_1748,N_873,N_755);
nand U1749 (N_1749,N_1063,N_1016);
or U1750 (N_1750,N_716,N_659);
nand U1751 (N_1751,N_892,N_740);
or U1752 (N_1752,N_874,N_1096);
nand U1753 (N_1753,N_897,N_1083);
nor U1754 (N_1754,N_1129,N_644);
or U1755 (N_1755,N_1021,N_903);
nor U1756 (N_1756,N_890,N_904);
nand U1757 (N_1757,N_992,N_860);
or U1758 (N_1758,N_1025,N_698);
or U1759 (N_1759,N_1142,N_734);
and U1760 (N_1760,N_1147,N_885);
nor U1761 (N_1761,N_1131,N_704);
and U1762 (N_1762,N_792,N_934);
nor U1763 (N_1763,N_867,N_1177);
nand U1764 (N_1764,N_674,N_1162);
nand U1765 (N_1765,N_673,N_1168);
nor U1766 (N_1766,N_727,N_655);
nand U1767 (N_1767,N_870,N_614);
and U1768 (N_1768,N_875,N_1162);
nor U1769 (N_1769,N_1164,N_750);
or U1770 (N_1770,N_1059,N_881);
nor U1771 (N_1771,N_636,N_921);
nand U1772 (N_1772,N_887,N_812);
nand U1773 (N_1773,N_1132,N_869);
and U1774 (N_1774,N_1067,N_787);
and U1775 (N_1775,N_970,N_1130);
and U1776 (N_1776,N_966,N_847);
nor U1777 (N_1777,N_766,N_688);
and U1778 (N_1778,N_789,N_901);
or U1779 (N_1779,N_698,N_774);
or U1780 (N_1780,N_1188,N_673);
and U1781 (N_1781,N_811,N_818);
nor U1782 (N_1782,N_670,N_824);
and U1783 (N_1783,N_682,N_805);
nand U1784 (N_1784,N_891,N_1185);
and U1785 (N_1785,N_622,N_1149);
or U1786 (N_1786,N_1110,N_1122);
or U1787 (N_1787,N_809,N_1174);
nand U1788 (N_1788,N_1164,N_716);
or U1789 (N_1789,N_1047,N_1031);
and U1790 (N_1790,N_788,N_638);
or U1791 (N_1791,N_748,N_805);
nand U1792 (N_1792,N_1053,N_633);
nand U1793 (N_1793,N_813,N_935);
nand U1794 (N_1794,N_763,N_692);
or U1795 (N_1795,N_998,N_848);
nor U1796 (N_1796,N_979,N_659);
nor U1797 (N_1797,N_794,N_755);
or U1798 (N_1798,N_1199,N_908);
nand U1799 (N_1799,N_631,N_792);
and U1800 (N_1800,N_1380,N_1222);
nor U1801 (N_1801,N_1565,N_1396);
or U1802 (N_1802,N_1437,N_1470);
nor U1803 (N_1803,N_1683,N_1338);
nand U1804 (N_1804,N_1295,N_1286);
nand U1805 (N_1805,N_1799,N_1612);
nor U1806 (N_1806,N_1402,N_1452);
or U1807 (N_1807,N_1635,N_1644);
or U1808 (N_1808,N_1447,N_1462);
nor U1809 (N_1809,N_1468,N_1758);
and U1810 (N_1810,N_1495,N_1742);
and U1811 (N_1811,N_1527,N_1574);
nand U1812 (N_1812,N_1647,N_1692);
or U1813 (N_1813,N_1508,N_1326);
nor U1814 (N_1814,N_1765,N_1419);
nor U1815 (N_1815,N_1327,N_1601);
nor U1816 (N_1816,N_1250,N_1710);
and U1817 (N_1817,N_1637,N_1448);
or U1818 (N_1818,N_1507,N_1285);
and U1819 (N_1819,N_1657,N_1283);
and U1820 (N_1820,N_1522,N_1340);
or U1821 (N_1821,N_1735,N_1541);
and U1822 (N_1822,N_1444,N_1537);
or U1823 (N_1823,N_1602,N_1525);
and U1824 (N_1824,N_1685,N_1705);
and U1825 (N_1825,N_1782,N_1369);
and U1826 (N_1826,N_1757,N_1678);
xor U1827 (N_1827,N_1439,N_1709);
and U1828 (N_1828,N_1335,N_1371);
nor U1829 (N_1829,N_1309,N_1490);
nand U1830 (N_1830,N_1526,N_1467);
nand U1831 (N_1831,N_1622,N_1339);
and U1832 (N_1832,N_1551,N_1767);
and U1833 (N_1833,N_1681,N_1384);
or U1834 (N_1834,N_1484,N_1481);
nand U1835 (N_1835,N_1455,N_1229);
nor U1836 (N_1836,N_1276,N_1759);
nor U1837 (N_1837,N_1214,N_1624);
and U1838 (N_1838,N_1302,N_1723);
and U1839 (N_1839,N_1475,N_1756);
and U1840 (N_1840,N_1204,N_1400);
nand U1841 (N_1841,N_1218,N_1798);
and U1842 (N_1842,N_1228,N_1347);
xor U1843 (N_1843,N_1581,N_1307);
nor U1844 (N_1844,N_1586,N_1571);
or U1845 (N_1845,N_1255,N_1364);
and U1846 (N_1846,N_1442,N_1515);
and U1847 (N_1847,N_1252,N_1290);
or U1848 (N_1848,N_1403,N_1784);
and U1849 (N_1849,N_1698,N_1535);
nand U1850 (N_1850,N_1781,N_1769);
nand U1851 (N_1851,N_1477,N_1377);
nor U1852 (N_1852,N_1443,N_1329);
or U1853 (N_1853,N_1320,N_1634);
nor U1854 (N_1854,N_1249,N_1245);
nand U1855 (N_1855,N_1337,N_1240);
nor U1856 (N_1856,N_1568,N_1479);
nor U1857 (N_1857,N_1744,N_1207);
nand U1858 (N_1858,N_1332,N_1270);
nand U1859 (N_1859,N_1405,N_1243);
nand U1860 (N_1860,N_1621,N_1786);
nor U1861 (N_1861,N_1755,N_1203);
and U1862 (N_1862,N_1510,N_1740);
or U1863 (N_1863,N_1458,N_1609);
nor U1864 (N_1864,N_1673,N_1366);
nor U1865 (N_1865,N_1220,N_1473);
and U1866 (N_1866,N_1362,N_1517);
and U1867 (N_1867,N_1736,N_1793);
or U1868 (N_1868,N_1411,N_1753);
or U1869 (N_1869,N_1363,N_1355);
and U1870 (N_1870,N_1747,N_1259);
nand U1871 (N_1871,N_1783,N_1464);
or U1872 (N_1872,N_1393,N_1370);
nor U1873 (N_1873,N_1684,N_1227);
or U1874 (N_1874,N_1383,N_1655);
or U1875 (N_1875,N_1585,N_1548);
nor U1876 (N_1876,N_1210,N_1646);
and U1877 (N_1877,N_1534,N_1594);
nand U1878 (N_1878,N_1722,N_1668);
or U1879 (N_1879,N_1417,N_1365);
and U1880 (N_1880,N_1324,N_1712);
and U1881 (N_1881,N_1652,N_1288);
or U1882 (N_1882,N_1623,N_1351);
or U1883 (N_1883,N_1694,N_1772);
or U1884 (N_1884,N_1578,N_1472);
nor U1885 (N_1885,N_1558,N_1277);
or U1886 (N_1886,N_1592,N_1319);
nor U1887 (N_1887,N_1572,N_1717);
and U1888 (N_1888,N_1404,N_1353);
nor U1889 (N_1889,N_1361,N_1261);
nand U1890 (N_1890,N_1567,N_1432);
nor U1891 (N_1891,N_1780,N_1457);
nor U1892 (N_1892,N_1244,N_1532);
or U1893 (N_1893,N_1292,N_1459);
nand U1894 (N_1894,N_1768,N_1588);
and U1895 (N_1895,N_1566,N_1318);
nand U1896 (N_1896,N_1697,N_1346);
nor U1897 (N_1897,N_1303,N_1797);
nand U1898 (N_1898,N_1582,N_1715);
or U1899 (N_1899,N_1426,N_1381);
nand U1900 (N_1900,N_1289,N_1509);
nor U1901 (N_1901,N_1265,N_1299);
and U1902 (N_1902,N_1234,N_1570);
and U1903 (N_1903,N_1627,N_1354);
and U1904 (N_1904,N_1331,N_1616);
nor U1905 (N_1905,N_1410,N_1641);
nand U1906 (N_1906,N_1603,N_1737);
xnor U1907 (N_1907,N_1628,N_1496);
nand U1908 (N_1908,N_1390,N_1795);
nand U1909 (N_1909,N_1281,N_1375);
nand U1910 (N_1910,N_1385,N_1435);
and U1911 (N_1911,N_1438,N_1376);
nand U1912 (N_1912,N_1519,N_1626);
or U1913 (N_1913,N_1547,N_1304);
nor U1914 (N_1914,N_1675,N_1269);
nor U1915 (N_1915,N_1530,N_1284);
nor U1916 (N_1916,N_1614,N_1421);
nand U1917 (N_1917,N_1745,N_1267);
and U1918 (N_1918,N_1664,N_1341);
and U1919 (N_1919,N_1213,N_1764);
and U1920 (N_1920,N_1545,N_1241);
or U1921 (N_1921,N_1689,N_1751);
or U1922 (N_1922,N_1536,N_1590);
nand U1923 (N_1923,N_1414,N_1230);
and U1924 (N_1924,N_1445,N_1321);
nand U1925 (N_1925,N_1345,N_1311);
or U1926 (N_1926,N_1453,N_1407);
nor U1927 (N_1927,N_1555,N_1511);
and U1928 (N_1928,N_1636,N_1706);
nand U1929 (N_1929,N_1446,N_1659);
and U1930 (N_1930,N_1258,N_1776);
nand U1931 (N_1931,N_1687,N_1306);
nand U1932 (N_1932,N_1654,N_1454);
nand U1933 (N_1933,N_1556,N_1730);
and U1934 (N_1934,N_1314,N_1658);
nand U1935 (N_1935,N_1643,N_1785);
nor U1936 (N_1936,N_1696,N_1356);
nand U1937 (N_1937,N_1553,N_1499);
and U1938 (N_1938,N_1789,N_1591);
nand U1939 (N_1939,N_1246,N_1387);
nor U1940 (N_1940,N_1232,N_1278);
nand U1941 (N_1941,N_1498,N_1424);
and U1942 (N_1942,N_1373,N_1633);
nor U1943 (N_1943,N_1449,N_1703);
and U1944 (N_1944,N_1398,N_1544);
nand U1945 (N_1945,N_1262,N_1695);
nand U1946 (N_1946,N_1731,N_1313);
nand U1947 (N_1947,N_1274,N_1343);
or U1948 (N_1948,N_1580,N_1202);
or U1949 (N_1949,N_1762,N_1516);
nor U1950 (N_1950,N_1394,N_1268);
and U1951 (N_1951,N_1649,N_1300);
or U1952 (N_1952,N_1584,N_1433);
nor U1953 (N_1953,N_1266,N_1205);
or U1954 (N_1954,N_1531,N_1350);
nor U1955 (N_1955,N_1778,N_1520);
or U1956 (N_1956,N_1748,N_1349);
and U1957 (N_1957,N_1523,N_1429);
nor U1958 (N_1958,N_1334,N_1391);
nand U1959 (N_1959,N_1293,N_1330);
nor U1960 (N_1960,N_1598,N_1599);
nor U1961 (N_1961,N_1734,N_1677);
nor U1962 (N_1962,N_1233,N_1401);
nor U1963 (N_1963,N_1638,N_1587);
or U1964 (N_1964,N_1688,N_1716);
or U1965 (N_1965,N_1542,N_1450);
nor U1966 (N_1966,N_1593,N_1397);
nand U1967 (N_1967,N_1699,N_1409);
xnor U1968 (N_1968,N_1546,N_1619);
or U1969 (N_1969,N_1539,N_1482);
nand U1970 (N_1970,N_1251,N_1282);
nor U1971 (N_1971,N_1436,N_1392);
nand U1972 (N_1972,N_1679,N_1492);
nor U1973 (N_1973,N_1500,N_1691);
nand U1974 (N_1974,N_1749,N_1665);
xor U1975 (N_1975,N_1650,N_1201);
nor U1976 (N_1976,N_1298,N_1247);
nand U1977 (N_1977,N_1779,N_1763);
nor U1978 (N_1978,N_1615,N_1606);
or U1979 (N_1979,N_1231,N_1538);
or U1980 (N_1980,N_1617,N_1216);
nor U1981 (N_1981,N_1794,N_1322);
or U1982 (N_1982,N_1550,N_1474);
nand U1983 (N_1983,N_1427,N_1773);
nand U1984 (N_1984,N_1287,N_1708);
and U1985 (N_1985,N_1328,N_1771);
or U1986 (N_1986,N_1729,N_1440);
or U1987 (N_1987,N_1291,N_1388);
or U1988 (N_1988,N_1256,N_1512);
or U1989 (N_1989,N_1273,N_1235);
and U1990 (N_1990,N_1540,N_1596);
nor U1991 (N_1991,N_1333,N_1219);
and U1992 (N_1992,N_1352,N_1423);
nand U1993 (N_1993,N_1315,N_1653);
or U1994 (N_1994,N_1215,N_1465);
and U1995 (N_1995,N_1576,N_1663);
nand U1996 (N_1996,N_1260,N_1408);
nor U1997 (N_1997,N_1666,N_1728);
nand U1998 (N_1998,N_1718,N_1503);
nor U1999 (N_1999,N_1676,N_1750);
nand U2000 (N_2000,N_1790,N_1724);
nand U2001 (N_2001,N_1305,N_1554);
nand U2002 (N_2002,N_1669,N_1325);
or U2003 (N_2003,N_1721,N_1480);
or U2004 (N_2004,N_1224,N_1775);
nor U2005 (N_2005,N_1727,N_1504);
and U2006 (N_2006,N_1422,N_1359);
nor U2007 (N_2007,N_1386,N_1569);
nand U2008 (N_2008,N_1648,N_1533);
nand U2009 (N_2009,N_1752,N_1711);
nand U2010 (N_2010,N_1559,N_1577);
and U2011 (N_2011,N_1693,N_1389);
and U2012 (N_2012,N_1211,N_1713);
or U2013 (N_2013,N_1702,N_1726);
and U2014 (N_2014,N_1639,N_1733);
and U2015 (N_2015,N_1743,N_1223);
and U2016 (N_2016,N_1308,N_1682);
or U2017 (N_2017,N_1561,N_1497);
nand U2018 (N_2018,N_1301,N_1738);
and U2019 (N_2019,N_1670,N_1493);
nor U2020 (N_2020,N_1296,N_1557);
nand U2021 (N_2021,N_1760,N_1483);
or U2022 (N_2022,N_1469,N_1528);
xnor U2023 (N_2023,N_1342,N_1549);
nor U2024 (N_2024,N_1796,N_1336);
nand U2025 (N_2025,N_1506,N_1766);
nand U2026 (N_2026,N_1608,N_1264);
or U2027 (N_2027,N_1372,N_1631);
nand U2028 (N_2028,N_1310,N_1358);
and U2029 (N_2029,N_1297,N_1690);
or U2030 (N_2030,N_1257,N_1714);
nand U2031 (N_2031,N_1242,N_1275);
nand U2032 (N_2032,N_1543,N_1651);
nor U2033 (N_2033,N_1645,N_1209);
nand U2034 (N_2034,N_1254,N_1674);
xnor U2035 (N_2035,N_1378,N_1754);
nor U2036 (N_2036,N_1208,N_1348);
or U2037 (N_2037,N_1206,N_1357);
or U2038 (N_2038,N_1485,N_1595);
or U2039 (N_2039,N_1629,N_1524);
nor U2040 (N_2040,N_1788,N_1312);
nand U2041 (N_2041,N_1466,N_1662);
nand U2042 (N_2042,N_1672,N_1513);
nand U2043 (N_2043,N_1416,N_1605);
nor U2044 (N_2044,N_1271,N_1774);
nand U2045 (N_2045,N_1607,N_1611);
nor U2046 (N_2046,N_1279,N_1237);
and U2047 (N_2047,N_1478,N_1707);
and U2048 (N_2048,N_1502,N_1456);
and U2049 (N_2049,N_1604,N_1642);
and U2050 (N_2050,N_1471,N_1661);
or U2051 (N_2051,N_1518,N_1597);
nand U2052 (N_2052,N_1667,N_1430);
or U2053 (N_2053,N_1521,N_1476);
xnor U2054 (N_2054,N_1732,N_1217);
and U2055 (N_2055,N_1418,N_1494);
nor U2056 (N_2056,N_1640,N_1463);
and U2057 (N_2057,N_1441,N_1618);
and U2058 (N_2058,N_1560,N_1630);
and U2059 (N_2059,N_1399,N_1719);
nand U2060 (N_2060,N_1746,N_1344);
nor U2061 (N_2061,N_1514,N_1379);
nor U2062 (N_2062,N_1680,N_1787);
or U2063 (N_2063,N_1741,N_1704);
or U2064 (N_2064,N_1431,N_1610);
or U2065 (N_2065,N_1434,N_1671);
nand U2066 (N_2066,N_1374,N_1489);
nand U2067 (N_2067,N_1239,N_1316);
nor U2068 (N_2068,N_1294,N_1487);
or U2069 (N_2069,N_1739,N_1777);
nand U2070 (N_2070,N_1613,N_1412);
nand U2071 (N_2071,N_1563,N_1575);
or U2072 (N_2072,N_1420,N_1573);
nand U2073 (N_2073,N_1238,N_1323);
nor U2074 (N_2074,N_1200,N_1280);
nand U2075 (N_2075,N_1212,N_1367);
nand U2076 (N_2076,N_1620,N_1461);
and U2077 (N_2077,N_1488,N_1368);
or U2078 (N_2078,N_1263,N_1413);
or U2079 (N_2079,N_1460,N_1360);
nand U2080 (N_2080,N_1700,N_1701);
and U2081 (N_2081,N_1686,N_1225);
and U2082 (N_2082,N_1221,N_1725);
or U2083 (N_2083,N_1406,N_1317);
or U2084 (N_2084,N_1600,N_1564);
nand U2085 (N_2085,N_1486,N_1236);
or U2086 (N_2086,N_1562,N_1382);
and U2087 (N_2087,N_1589,N_1625);
nor U2088 (N_2088,N_1501,N_1791);
or U2089 (N_2089,N_1415,N_1552);
and U2090 (N_2090,N_1579,N_1720);
or U2091 (N_2091,N_1583,N_1226);
and U2092 (N_2092,N_1656,N_1491);
nand U2093 (N_2093,N_1792,N_1632);
nor U2094 (N_2094,N_1451,N_1428);
or U2095 (N_2095,N_1770,N_1425);
nor U2096 (N_2096,N_1529,N_1761);
nand U2097 (N_2097,N_1253,N_1248);
or U2098 (N_2098,N_1505,N_1395);
and U2099 (N_2099,N_1272,N_1660);
nor U2100 (N_2100,N_1334,N_1455);
nand U2101 (N_2101,N_1784,N_1696);
nor U2102 (N_2102,N_1690,N_1714);
and U2103 (N_2103,N_1405,N_1383);
and U2104 (N_2104,N_1504,N_1612);
and U2105 (N_2105,N_1649,N_1212);
or U2106 (N_2106,N_1294,N_1493);
nor U2107 (N_2107,N_1587,N_1769);
nor U2108 (N_2108,N_1722,N_1696);
nor U2109 (N_2109,N_1617,N_1583);
nand U2110 (N_2110,N_1624,N_1646);
and U2111 (N_2111,N_1612,N_1660);
or U2112 (N_2112,N_1347,N_1304);
nand U2113 (N_2113,N_1235,N_1479);
or U2114 (N_2114,N_1636,N_1292);
nand U2115 (N_2115,N_1435,N_1620);
nand U2116 (N_2116,N_1253,N_1478);
and U2117 (N_2117,N_1762,N_1774);
nand U2118 (N_2118,N_1502,N_1634);
and U2119 (N_2119,N_1643,N_1238);
or U2120 (N_2120,N_1284,N_1291);
and U2121 (N_2121,N_1407,N_1561);
or U2122 (N_2122,N_1774,N_1541);
nand U2123 (N_2123,N_1330,N_1269);
or U2124 (N_2124,N_1354,N_1583);
nor U2125 (N_2125,N_1710,N_1527);
and U2126 (N_2126,N_1742,N_1358);
nor U2127 (N_2127,N_1431,N_1580);
nor U2128 (N_2128,N_1560,N_1248);
and U2129 (N_2129,N_1781,N_1363);
nor U2130 (N_2130,N_1207,N_1653);
or U2131 (N_2131,N_1581,N_1467);
and U2132 (N_2132,N_1706,N_1507);
nor U2133 (N_2133,N_1694,N_1213);
and U2134 (N_2134,N_1203,N_1300);
nor U2135 (N_2135,N_1663,N_1294);
and U2136 (N_2136,N_1466,N_1319);
nand U2137 (N_2137,N_1682,N_1708);
nand U2138 (N_2138,N_1383,N_1460);
and U2139 (N_2139,N_1410,N_1362);
or U2140 (N_2140,N_1522,N_1531);
nor U2141 (N_2141,N_1562,N_1793);
and U2142 (N_2142,N_1321,N_1275);
nand U2143 (N_2143,N_1225,N_1231);
and U2144 (N_2144,N_1746,N_1354);
and U2145 (N_2145,N_1390,N_1280);
nor U2146 (N_2146,N_1214,N_1715);
and U2147 (N_2147,N_1747,N_1222);
or U2148 (N_2148,N_1613,N_1542);
nor U2149 (N_2149,N_1620,N_1488);
or U2150 (N_2150,N_1473,N_1203);
or U2151 (N_2151,N_1787,N_1201);
nor U2152 (N_2152,N_1573,N_1219);
or U2153 (N_2153,N_1225,N_1254);
nand U2154 (N_2154,N_1255,N_1343);
nor U2155 (N_2155,N_1241,N_1318);
nor U2156 (N_2156,N_1761,N_1647);
or U2157 (N_2157,N_1547,N_1395);
nor U2158 (N_2158,N_1730,N_1300);
xnor U2159 (N_2159,N_1365,N_1241);
nand U2160 (N_2160,N_1547,N_1785);
nor U2161 (N_2161,N_1771,N_1659);
and U2162 (N_2162,N_1687,N_1285);
and U2163 (N_2163,N_1672,N_1470);
nand U2164 (N_2164,N_1766,N_1624);
and U2165 (N_2165,N_1249,N_1373);
or U2166 (N_2166,N_1766,N_1794);
nor U2167 (N_2167,N_1429,N_1544);
xor U2168 (N_2168,N_1345,N_1232);
and U2169 (N_2169,N_1422,N_1557);
nor U2170 (N_2170,N_1328,N_1492);
or U2171 (N_2171,N_1276,N_1622);
nor U2172 (N_2172,N_1458,N_1577);
or U2173 (N_2173,N_1389,N_1380);
or U2174 (N_2174,N_1452,N_1495);
nand U2175 (N_2175,N_1374,N_1573);
nand U2176 (N_2176,N_1536,N_1357);
or U2177 (N_2177,N_1523,N_1273);
or U2178 (N_2178,N_1288,N_1363);
and U2179 (N_2179,N_1576,N_1348);
or U2180 (N_2180,N_1334,N_1497);
nor U2181 (N_2181,N_1399,N_1584);
nand U2182 (N_2182,N_1395,N_1556);
nor U2183 (N_2183,N_1495,N_1665);
nand U2184 (N_2184,N_1426,N_1798);
or U2185 (N_2185,N_1715,N_1419);
and U2186 (N_2186,N_1767,N_1547);
nor U2187 (N_2187,N_1442,N_1530);
and U2188 (N_2188,N_1584,N_1533);
nand U2189 (N_2189,N_1705,N_1621);
and U2190 (N_2190,N_1320,N_1696);
nand U2191 (N_2191,N_1431,N_1313);
nand U2192 (N_2192,N_1758,N_1611);
or U2193 (N_2193,N_1606,N_1388);
nor U2194 (N_2194,N_1765,N_1787);
and U2195 (N_2195,N_1664,N_1254);
nand U2196 (N_2196,N_1732,N_1682);
and U2197 (N_2197,N_1322,N_1479);
nand U2198 (N_2198,N_1336,N_1666);
or U2199 (N_2199,N_1274,N_1734);
or U2200 (N_2200,N_1641,N_1518);
or U2201 (N_2201,N_1276,N_1515);
and U2202 (N_2202,N_1792,N_1375);
nor U2203 (N_2203,N_1323,N_1688);
nor U2204 (N_2204,N_1272,N_1241);
and U2205 (N_2205,N_1394,N_1734);
nor U2206 (N_2206,N_1559,N_1598);
or U2207 (N_2207,N_1215,N_1408);
and U2208 (N_2208,N_1494,N_1724);
nand U2209 (N_2209,N_1322,N_1689);
nand U2210 (N_2210,N_1746,N_1378);
and U2211 (N_2211,N_1728,N_1491);
nor U2212 (N_2212,N_1408,N_1309);
nand U2213 (N_2213,N_1541,N_1577);
nor U2214 (N_2214,N_1466,N_1549);
nor U2215 (N_2215,N_1579,N_1426);
nor U2216 (N_2216,N_1736,N_1299);
or U2217 (N_2217,N_1317,N_1699);
or U2218 (N_2218,N_1786,N_1294);
nand U2219 (N_2219,N_1650,N_1412);
nand U2220 (N_2220,N_1758,N_1497);
nand U2221 (N_2221,N_1467,N_1627);
and U2222 (N_2222,N_1383,N_1582);
or U2223 (N_2223,N_1693,N_1350);
or U2224 (N_2224,N_1302,N_1278);
nand U2225 (N_2225,N_1445,N_1617);
nand U2226 (N_2226,N_1204,N_1403);
nor U2227 (N_2227,N_1702,N_1557);
and U2228 (N_2228,N_1412,N_1428);
and U2229 (N_2229,N_1793,N_1681);
and U2230 (N_2230,N_1522,N_1458);
or U2231 (N_2231,N_1797,N_1270);
nand U2232 (N_2232,N_1218,N_1466);
nor U2233 (N_2233,N_1522,N_1692);
nand U2234 (N_2234,N_1551,N_1742);
and U2235 (N_2235,N_1292,N_1302);
or U2236 (N_2236,N_1786,N_1582);
and U2237 (N_2237,N_1345,N_1512);
nand U2238 (N_2238,N_1624,N_1251);
and U2239 (N_2239,N_1413,N_1451);
or U2240 (N_2240,N_1755,N_1754);
and U2241 (N_2241,N_1642,N_1477);
nand U2242 (N_2242,N_1751,N_1282);
nor U2243 (N_2243,N_1259,N_1547);
nand U2244 (N_2244,N_1734,N_1532);
and U2245 (N_2245,N_1763,N_1677);
and U2246 (N_2246,N_1394,N_1528);
or U2247 (N_2247,N_1220,N_1794);
nand U2248 (N_2248,N_1321,N_1231);
and U2249 (N_2249,N_1611,N_1267);
nand U2250 (N_2250,N_1215,N_1537);
nor U2251 (N_2251,N_1455,N_1566);
and U2252 (N_2252,N_1207,N_1584);
or U2253 (N_2253,N_1708,N_1595);
or U2254 (N_2254,N_1429,N_1245);
and U2255 (N_2255,N_1392,N_1238);
and U2256 (N_2256,N_1410,N_1665);
nor U2257 (N_2257,N_1592,N_1656);
or U2258 (N_2258,N_1596,N_1346);
nor U2259 (N_2259,N_1420,N_1229);
or U2260 (N_2260,N_1303,N_1642);
or U2261 (N_2261,N_1498,N_1794);
and U2262 (N_2262,N_1727,N_1609);
and U2263 (N_2263,N_1700,N_1735);
nand U2264 (N_2264,N_1783,N_1795);
nor U2265 (N_2265,N_1726,N_1421);
nor U2266 (N_2266,N_1750,N_1376);
or U2267 (N_2267,N_1356,N_1294);
and U2268 (N_2268,N_1457,N_1645);
nand U2269 (N_2269,N_1621,N_1683);
and U2270 (N_2270,N_1567,N_1666);
nor U2271 (N_2271,N_1527,N_1399);
nor U2272 (N_2272,N_1412,N_1508);
or U2273 (N_2273,N_1228,N_1674);
nor U2274 (N_2274,N_1243,N_1651);
or U2275 (N_2275,N_1464,N_1237);
or U2276 (N_2276,N_1358,N_1327);
nor U2277 (N_2277,N_1540,N_1438);
nor U2278 (N_2278,N_1721,N_1484);
nand U2279 (N_2279,N_1302,N_1521);
nand U2280 (N_2280,N_1455,N_1500);
or U2281 (N_2281,N_1523,N_1432);
and U2282 (N_2282,N_1539,N_1485);
nor U2283 (N_2283,N_1502,N_1566);
nor U2284 (N_2284,N_1617,N_1651);
nor U2285 (N_2285,N_1531,N_1355);
nand U2286 (N_2286,N_1725,N_1782);
or U2287 (N_2287,N_1762,N_1509);
nand U2288 (N_2288,N_1208,N_1237);
and U2289 (N_2289,N_1554,N_1546);
nor U2290 (N_2290,N_1543,N_1368);
and U2291 (N_2291,N_1471,N_1656);
or U2292 (N_2292,N_1616,N_1337);
or U2293 (N_2293,N_1317,N_1614);
nor U2294 (N_2294,N_1346,N_1451);
or U2295 (N_2295,N_1750,N_1490);
nand U2296 (N_2296,N_1206,N_1762);
and U2297 (N_2297,N_1228,N_1624);
or U2298 (N_2298,N_1234,N_1223);
or U2299 (N_2299,N_1427,N_1736);
nand U2300 (N_2300,N_1431,N_1248);
and U2301 (N_2301,N_1759,N_1647);
nand U2302 (N_2302,N_1309,N_1232);
and U2303 (N_2303,N_1603,N_1720);
and U2304 (N_2304,N_1373,N_1431);
nand U2305 (N_2305,N_1521,N_1673);
or U2306 (N_2306,N_1736,N_1717);
nor U2307 (N_2307,N_1442,N_1295);
and U2308 (N_2308,N_1495,N_1209);
and U2309 (N_2309,N_1225,N_1545);
nand U2310 (N_2310,N_1574,N_1525);
nor U2311 (N_2311,N_1432,N_1653);
xnor U2312 (N_2312,N_1734,N_1355);
nand U2313 (N_2313,N_1543,N_1669);
and U2314 (N_2314,N_1650,N_1459);
nor U2315 (N_2315,N_1674,N_1576);
and U2316 (N_2316,N_1548,N_1482);
nand U2317 (N_2317,N_1601,N_1694);
nand U2318 (N_2318,N_1280,N_1407);
nand U2319 (N_2319,N_1699,N_1682);
nand U2320 (N_2320,N_1517,N_1365);
nor U2321 (N_2321,N_1672,N_1529);
nor U2322 (N_2322,N_1711,N_1796);
and U2323 (N_2323,N_1790,N_1791);
or U2324 (N_2324,N_1314,N_1426);
nor U2325 (N_2325,N_1370,N_1413);
nand U2326 (N_2326,N_1439,N_1365);
or U2327 (N_2327,N_1609,N_1206);
nand U2328 (N_2328,N_1416,N_1787);
nand U2329 (N_2329,N_1544,N_1679);
nor U2330 (N_2330,N_1506,N_1317);
nor U2331 (N_2331,N_1399,N_1793);
nor U2332 (N_2332,N_1677,N_1428);
and U2333 (N_2333,N_1575,N_1488);
nand U2334 (N_2334,N_1540,N_1319);
nor U2335 (N_2335,N_1696,N_1343);
and U2336 (N_2336,N_1722,N_1745);
nor U2337 (N_2337,N_1626,N_1749);
or U2338 (N_2338,N_1645,N_1554);
or U2339 (N_2339,N_1590,N_1343);
nor U2340 (N_2340,N_1213,N_1637);
and U2341 (N_2341,N_1348,N_1698);
nand U2342 (N_2342,N_1671,N_1695);
nand U2343 (N_2343,N_1565,N_1420);
nor U2344 (N_2344,N_1225,N_1442);
or U2345 (N_2345,N_1368,N_1304);
or U2346 (N_2346,N_1394,N_1202);
nor U2347 (N_2347,N_1524,N_1374);
and U2348 (N_2348,N_1726,N_1508);
and U2349 (N_2349,N_1315,N_1557);
or U2350 (N_2350,N_1691,N_1213);
and U2351 (N_2351,N_1334,N_1583);
nor U2352 (N_2352,N_1790,N_1627);
and U2353 (N_2353,N_1509,N_1453);
or U2354 (N_2354,N_1518,N_1434);
and U2355 (N_2355,N_1305,N_1378);
nand U2356 (N_2356,N_1629,N_1397);
and U2357 (N_2357,N_1577,N_1671);
nor U2358 (N_2358,N_1220,N_1402);
or U2359 (N_2359,N_1507,N_1312);
nor U2360 (N_2360,N_1212,N_1279);
and U2361 (N_2361,N_1405,N_1208);
and U2362 (N_2362,N_1772,N_1366);
and U2363 (N_2363,N_1658,N_1279);
nor U2364 (N_2364,N_1329,N_1601);
nand U2365 (N_2365,N_1205,N_1309);
and U2366 (N_2366,N_1267,N_1793);
nor U2367 (N_2367,N_1417,N_1404);
and U2368 (N_2368,N_1384,N_1381);
nor U2369 (N_2369,N_1718,N_1562);
or U2370 (N_2370,N_1469,N_1592);
nor U2371 (N_2371,N_1430,N_1721);
or U2372 (N_2372,N_1452,N_1674);
nor U2373 (N_2373,N_1646,N_1452);
and U2374 (N_2374,N_1326,N_1660);
or U2375 (N_2375,N_1664,N_1327);
and U2376 (N_2376,N_1793,N_1682);
and U2377 (N_2377,N_1597,N_1523);
and U2378 (N_2378,N_1322,N_1260);
nor U2379 (N_2379,N_1678,N_1338);
nor U2380 (N_2380,N_1705,N_1758);
nor U2381 (N_2381,N_1752,N_1361);
or U2382 (N_2382,N_1442,N_1726);
nor U2383 (N_2383,N_1552,N_1687);
and U2384 (N_2384,N_1483,N_1642);
or U2385 (N_2385,N_1500,N_1308);
nand U2386 (N_2386,N_1590,N_1491);
nand U2387 (N_2387,N_1380,N_1334);
and U2388 (N_2388,N_1355,N_1375);
nand U2389 (N_2389,N_1571,N_1269);
and U2390 (N_2390,N_1544,N_1455);
or U2391 (N_2391,N_1200,N_1481);
nor U2392 (N_2392,N_1483,N_1237);
nand U2393 (N_2393,N_1247,N_1321);
xor U2394 (N_2394,N_1442,N_1219);
or U2395 (N_2395,N_1580,N_1434);
nand U2396 (N_2396,N_1779,N_1388);
or U2397 (N_2397,N_1569,N_1468);
or U2398 (N_2398,N_1729,N_1609);
nand U2399 (N_2399,N_1641,N_1735);
and U2400 (N_2400,N_1834,N_1843);
and U2401 (N_2401,N_1817,N_1963);
nand U2402 (N_2402,N_1996,N_2120);
xnor U2403 (N_2403,N_2084,N_2178);
nand U2404 (N_2404,N_2358,N_1972);
or U2405 (N_2405,N_2143,N_2075);
and U2406 (N_2406,N_1997,N_1859);
and U2407 (N_2407,N_2257,N_1899);
nor U2408 (N_2408,N_2185,N_2334);
nand U2409 (N_2409,N_2187,N_1992);
and U2410 (N_2410,N_1895,N_1999);
or U2411 (N_2411,N_2138,N_2147);
nand U2412 (N_2412,N_2333,N_1954);
nand U2413 (N_2413,N_1833,N_1876);
nor U2414 (N_2414,N_1837,N_2304);
or U2415 (N_2415,N_2205,N_2037);
and U2416 (N_2416,N_2064,N_2281);
and U2417 (N_2417,N_2276,N_1922);
and U2418 (N_2418,N_1910,N_2026);
nand U2419 (N_2419,N_2305,N_1950);
and U2420 (N_2420,N_1804,N_2137);
or U2421 (N_2421,N_1840,N_1943);
and U2422 (N_2422,N_1951,N_2396);
nand U2423 (N_2423,N_2105,N_2139);
or U2424 (N_2424,N_2390,N_2322);
and U2425 (N_2425,N_2110,N_2186);
nand U2426 (N_2426,N_1983,N_2010);
nand U2427 (N_2427,N_1842,N_1932);
and U2428 (N_2428,N_2014,N_2125);
nand U2429 (N_2429,N_2274,N_2005);
nand U2430 (N_2430,N_1930,N_2371);
and U2431 (N_2431,N_2340,N_1879);
or U2432 (N_2432,N_2286,N_2073);
or U2433 (N_2433,N_1894,N_2086);
and U2434 (N_2434,N_2391,N_2270);
nand U2435 (N_2435,N_2157,N_2079);
nand U2436 (N_2436,N_1914,N_2247);
nor U2437 (N_2437,N_2040,N_1911);
and U2438 (N_2438,N_1956,N_2301);
nor U2439 (N_2439,N_2130,N_2074);
nand U2440 (N_2440,N_1891,N_2122);
or U2441 (N_2441,N_2108,N_2284);
nand U2442 (N_2442,N_2168,N_1828);
and U2443 (N_2443,N_2214,N_2345);
nor U2444 (N_2444,N_2030,N_2017);
and U2445 (N_2445,N_2045,N_1819);
nand U2446 (N_2446,N_2366,N_2271);
or U2447 (N_2447,N_2029,N_2365);
and U2448 (N_2448,N_2294,N_1856);
nor U2449 (N_2449,N_1973,N_2269);
or U2450 (N_2450,N_2090,N_1959);
nand U2451 (N_2451,N_2212,N_2023);
nor U2452 (N_2452,N_2244,N_2135);
and U2453 (N_2453,N_1903,N_2024);
nor U2454 (N_2454,N_1867,N_2250);
nand U2455 (N_2455,N_2343,N_2346);
or U2456 (N_2456,N_1800,N_2353);
and U2457 (N_2457,N_2208,N_1863);
and U2458 (N_2458,N_2044,N_2132);
nor U2459 (N_2459,N_2375,N_2394);
and U2460 (N_2460,N_2190,N_2312);
nand U2461 (N_2461,N_2240,N_2159);
or U2462 (N_2462,N_1912,N_1832);
or U2463 (N_2463,N_2133,N_1925);
nor U2464 (N_2464,N_2330,N_1822);
nor U2465 (N_2465,N_2350,N_1946);
nand U2466 (N_2466,N_2302,N_2089);
nand U2467 (N_2467,N_2359,N_2230);
nand U2468 (N_2468,N_1919,N_2326);
or U2469 (N_2469,N_2141,N_1916);
or U2470 (N_2470,N_2188,N_2162);
or U2471 (N_2471,N_2006,N_2238);
nand U2472 (N_2472,N_2287,N_2316);
and U2473 (N_2473,N_1998,N_2058);
nor U2474 (N_2474,N_2021,N_2289);
xnor U2475 (N_2475,N_2228,N_1872);
or U2476 (N_2476,N_2374,N_1862);
and U2477 (N_2477,N_2131,N_1830);
or U2478 (N_2478,N_1978,N_2171);
nor U2479 (N_2479,N_1814,N_1927);
nor U2480 (N_2480,N_2278,N_2226);
nor U2481 (N_2481,N_1926,N_1921);
nand U2482 (N_2482,N_2095,N_2013);
and U2483 (N_2483,N_1945,N_2174);
and U2484 (N_2484,N_2169,N_1934);
nor U2485 (N_2485,N_2252,N_2164);
nand U2486 (N_2486,N_1857,N_1969);
nor U2487 (N_2487,N_2210,N_2241);
nor U2488 (N_2488,N_1940,N_1929);
or U2489 (N_2489,N_2329,N_2196);
or U2490 (N_2490,N_2016,N_1836);
or U2491 (N_2491,N_2076,N_2148);
and U2492 (N_2492,N_2007,N_2096);
nor U2493 (N_2493,N_1896,N_2062);
nand U2494 (N_2494,N_2246,N_1960);
nand U2495 (N_2495,N_2236,N_1964);
nand U2496 (N_2496,N_2153,N_1952);
and U2497 (N_2497,N_2039,N_2380);
nand U2498 (N_2498,N_2221,N_2314);
and U2499 (N_2499,N_1987,N_1850);
and U2500 (N_2500,N_2383,N_1980);
and U2501 (N_2501,N_2012,N_2046);
or U2502 (N_2502,N_2170,N_1838);
nand U2503 (N_2503,N_2382,N_2160);
nand U2504 (N_2504,N_1884,N_1801);
nor U2505 (N_2505,N_2117,N_2248);
and U2506 (N_2506,N_2290,N_1824);
and U2507 (N_2507,N_1897,N_2167);
nor U2508 (N_2508,N_2140,N_1971);
or U2509 (N_2509,N_2384,N_1913);
or U2510 (N_2510,N_2348,N_2328);
and U2511 (N_2511,N_2273,N_2386);
and U2512 (N_2512,N_2027,N_2354);
nor U2513 (N_2513,N_2056,N_2088);
nor U2514 (N_2514,N_2071,N_2115);
nand U2515 (N_2515,N_2112,N_2189);
and U2516 (N_2516,N_1846,N_1851);
and U2517 (N_2517,N_2155,N_2243);
and U2518 (N_2518,N_2233,N_1957);
and U2519 (N_2519,N_2197,N_1935);
and U2520 (N_2520,N_2379,N_2003);
and U2521 (N_2521,N_1982,N_2082);
nand U2522 (N_2522,N_2259,N_2283);
and U2523 (N_2523,N_2191,N_2085);
or U2524 (N_2524,N_2194,N_2065);
nor U2525 (N_2525,N_2372,N_1803);
or U2526 (N_2526,N_2083,N_2367);
nand U2527 (N_2527,N_2063,N_2253);
or U2528 (N_2528,N_2018,N_2198);
nand U2529 (N_2529,N_1942,N_1829);
or U2530 (N_2530,N_2300,N_2267);
nor U2531 (N_2531,N_2048,N_2193);
and U2532 (N_2532,N_2227,N_2277);
nor U2533 (N_2533,N_2310,N_1809);
nand U2534 (N_2534,N_1878,N_2142);
nand U2535 (N_2535,N_2184,N_1966);
nand U2536 (N_2536,N_2091,N_1841);
or U2537 (N_2537,N_1868,N_2320);
nor U2538 (N_2538,N_1881,N_2126);
and U2539 (N_2539,N_2303,N_1818);
nand U2540 (N_2540,N_1944,N_1904);
or U2541 (N_2541,N_1870,N_2323);
nor U2542 (N_2542,N_1962,N_1941);
nor U2543 (N_2543,N_1989,N_2098);
nor U2544 (N_2544,N_2092,N_2363);
or U2545 (N_2545,N_2388,N_1816);
or U2546 (N_2546,N_1953,N_2008);
or U2547 (N_2547,N_2308,N_2035);
nor U2548 (N_2548,N_2114,N_2034);
or U2549 (N_2549,N_2009,N_2373);
and U2550 (N_2550,N_2124,N_2203);
and U2551 (N_2551,N_2195,N_2204);
or U2552 (N_2552,N_1855,N_2339);
nand U2553 (N_2553,N_2225,N_2093);
nor U2554 (N_2554,N_2172,N_2235);
nor U2555 (N_2555,N_2206,N_1958);
nor U2556 (N_2556,N_2097,N_2192);
nor U2557 (N_2557,N_2389,N_2261);
nand U2558 (N_2558,N_1835,N_1813);
nand U2559 (N_2559,N_2004,N_2150);
or U2560 (N_2560,N_2217,N_2176);
nand U2561 (N_2561,N_1948,N_1908);
nand U2562 (N_2562,N_1882,N_2166);
or U2563 (N_2563,N_2070,N_1885);
or U2564 (N_2564,N_1805,N_2033);
and U2565 (N_2565,N_2337,N_1984);
or U2566 (N_2566,N_1864,N_1890);
nor U2567 (N_2567,N_2047,N_2293);
or U2568 (N_2568,N_2213,N_2199);
nand U2569 (N_2569,N_2051,N_1923);
and U2570 (N_2570,N_1839,N_1947);
nand U2571 (N_2571,N_1924,N_2220);
and U2572 (N_2572,N_2069,N_1865);
or U2573 (N_2573,N_2218,N_2260);
nand U2574 (N_2574,N_2280,N_2202);
and U2575 (N_2575,N_2331,N_2224);
nand U2576 (N_2576,N_2352,N_2151);
nand U2577 (N_2577,N_2313,N_1853);
and U2578 (N_2578,N_2081,N_1976);
or U2579 (N_2579,N_1961,N_1931);
nand U2580 (N_2580,N_2078,N_2355);
or U2581 (N_2581,N_2041,N_2099);
nand U2582 (N_2582,N_2387,N_1938);
nor U2583 (N_2583,N_2393,N_2177);
or U2584 (N_2584,N_1986,N_2128);
and U2585 (N_2585,N_2161,N_2042);
nor U2586 (N_2586,N_2344,N_2136);
and U2587 (N_2587,N_1871,N_2275);
or U2588 (N_2588,N_2043,N_1906);
and U2589 (N_2589,N_2001,N_2307);
and U2590 (N_2590,N_2038,N_1887);
and U2591 (N_2591,N_2272,N_2002);
nor U2592 (N_2592,N_2362,N_2364);
nor U2593 (N_2593,N_2036,N_2360);
nand U2594 (N_2594,N_1848,N_2101);
nor U2595 (N_2595,N_2180,N_1854);
and U2596 (N_2596,N_2255,N_2123);
or U2597 (N_2597,N_1820,N_2298);
nand U2598 (N_2598,N_2378,N_1979);
nor U2599 (N_2599,N_2223,N_2342);
or U2600 (N_2600,N_1915,N_2067);
nor U2601 (N_2601,N_2256,N_2116);
or U2602 (N_2602,N_1985,N_2368);
and U2603 (N_2603,N_2154,N_1901);
nand U2604 (N_2604,N_2052,N_1849);
nor U2605 (N_2605,N_2315,N_1905);
or U2606 (N_2606,N_2049,N_1821);
nand U2607 (N_2607,N_1812,N_2061);
nor U2608 (N_2608,N_1852,N_2055);
nor U2609 (N_2609,N_2309,N_1810);
or U2610 (N_2610,N_2295,N_2060);
and U2611 (N_2611,N_2000,N_1808);
or U2612 (N_2612,N_2216,N_2222);
nor U2613 (N_2613,N_2183,N_2175);
and U2614 (N_2614,N_2237,N_2207);
and U2615 (N_2615,N_2392,N_1845);
nor U2616 (N_2616,N_2242,N_1807);
nand U2617 (N_2617,N_2025,N_1811);
nor U2618 (N_2618,N_1883,N_2251);
nand U2619 (N_2619,N_2182,N_1975);
nand U2620 (N_2620,N_2299,N_1893);
and U2621 (N_2621,N_2134,N_1827);
and U2622 (N_2622,N_1970,N_2209);
and U2623 (N_2623,N_2111,N_1858);
nand U2624 (N_2624,N_2361,N_2318);
nor U2625 (N_2625,N_2031,N_2011);
nor U2626 (N_2626,N_2231,N_2292);
nand U2627 (N_2627,N_2152,N_2156);
nor U2628 (N_2628,N_1918,N_2254);
and U2629 (N_2629,N_2144,N_2266);
nand U2630 (N_2630,N_1967,N_1877);
and U2631 (N_2631,N_2127,N_2102);
and U2632 (N_2632,N_2336,N_2028);
xnor U2633 (N_2633,N_2381,N_1917);
or U2634 (N_2634,N_2077,N_2129);
nor U2635 (N_2635,N_2104,N_1866);
nand U2636 (N_2636,N_1869,N_2109);
and U2637 (N_2637,N_2291,N_2219);
nor U2638 (N_2638,N_1860,N_2249);
and U2639 (N_2639,N_2398,N_2121);
nor U2640 (N_2640,N_2106,N_2215);
nand U2641 (N_2641,N_2311,N_2385);
nand U2642 (N_2642,N_2068,N_1937);
or U2643 (N_2643,N_2179,N_2211);
nor U2644 (N_2644,N_2181,N_1825);
nand U2645 (N_2645,N_1990,N_1965);
or U2646 (N_2646,N_1844,N_2370);
and U2647 (N_2647,N_2173,N_2053);
or U2648 (N_2648,N_2072,N_2019);
and U2649 (N_2649,N_2317,N_1875);
and U2650 (N_2650,N_1892,N_1907);
or U2651 (N_2651,N_2145,N_2264);
or U2652 (N_2652,N_1936,N_2015);
and U2653 (N_2653,N_2262,N_1933);
nor U2654 (N_2654,N_1928,N_2245);
or U2655 (N_2655,N_2080,N_1909);
nor U2656 (N_2656,N_1806,N_1991);
nor U2657 (N_2657,N_2032,N_1888);
or U2658 (N_2658,N_2324,N_2397);
nor U2659 (N_2659,N_2338,N_2146);
nand U2660 (N_2660,N_2113,N_2229);
nand U2661 (N_2661,N_2265,N_2327);
and U2662 (N_2662,N_1880,N_2296);
and U2663 (N_2663,N_2268,N_2376);
nand U2664 (N_2664,N_1955,N_1898);
or U2665 (N_2665,N_2232,N_2057);
nor U2666 (N_2666,N_1826,N_2347);
nand U2667 (N_2667,N_1874,N_1993);
and U2668 (N_2668,N_2297,N_2258);
nand U2669 (N_2669,N_2054,N_2059);
and U2670 (N_2670,N_2094,N_2349);
and U2671 (N_2671,N_2325,N_2022);
and U2672 (N_2672,N_1889,N_1861);
and U2673 (N_2673,N_1823,N_1988);
and U2674 (N_2674,N_2066,N_2239);
or U2675 (N_2675,N_2149,N_2288);
nand U2676 (N_2676,N_2100,N_1994);
and U2677 (N_2677,N_2351,N_2357);
and U2678 (N_2678,N_2158,N_1968);
nand U2679 (N_2679,N_2263,N_2369);
nor U2680 (N_2680,N_2395,N_1902);
and U2681 (N_2681,N_1815,N_2321);
or U2682 (N_2682,N_1949,N_1831);
nand U2683 (N_2683,N_2377,N_2103);
nor U2684 (N_2684,N_2118,N_1974);
or U2685 (N_2685,N_1886,N_1920);
nand U2686 (N_2686,N_2119,N_2306);
nor U2687 (N_2687,N_1802,N_2200);
and U2688 (N_2688,N_2201,N_2282);
nor U2689 (N_2689,N_2050,N_2279);
nand U2690 (N_2690,N_2165,N_1847);
nor U2691 (N_2691,N_2335,N_2356);
nand U2692 (N_2692,N_2332,N_2341);
nor U2693 (N_2693,N_1977,N_2163);
nor U2694 (N_2694,N_2319,N_1873);
nor U2695 (N_2695,N_1981,N_1939);
or U2696 (N_2696,N_2020,N_1900);
nand U2697 (N_2697,N_2285,N_2399);
and U2698 (N_2698,N_2087,N_2107);
and U2699 (N_2699,N_2234,N_1995);
xor U2700 (N_2700,N_2296,N_1813);
nor U2701 (N_2701,N_2199,N_2381);
or U2702 (N_2702,N_2375,N_1905);
and U2703 (N_2703,N_2233,N_1954);
and U2704 (N_2704,N_1865,N_2358);
or U2705 (N_2705,N_2284,N_1831);
or U2706 (N_2706,N_1856,N_1818);
or U2707 (N_2707,N_1947,N_2389);
nor U2708 (N_2708,N_2287,N_2115);
or U2709 (N_2709,N_1992,N_1873);
or U2710 (N_2710,N_2097,N_2379);
and U2711 (N_2711,N_1848,N_2006);
nand U2712 (N_2712,N_2166,N_2027);
nand U2713 (N_2713,N_2251,N_2180);
or U2714 (N_2714,N_2051,N_1893);
nor U2715 (N_2715,N_1966,N_1823);
or U2716 (N_2716,N_2255,N_2293);
and U2717 (N_2717,N_1812,N_2375);
or U2718 (N_2718,N_2334,N_1819);
nor U2719 (N_2719,N_1905,N_2304);
nand U2720 (N_2720,N_2139,N_2305);
and U2721 (N_2721,N_2142,N_2056);
nor U2722 (N_2722,N_2077,N_2356);
nor U2723 (N_2723,N_1805,N_1825);
or U2724 (N_2724,N_2260,N_2178);
or U2725 (N_2725,N_2229,N_2336);
and U2726 (N_2726,N_2085,N_1824);
or U2727 (N_2727,N_2377,N_2124);
nor U2728 (N_2728,N_2131,N_1995);
and U2729 (N_2729,N_2313,N_2207);
nand U2730 (N_2730,N_1856,N_1974);
and U2731 (N_2731,N_2218,N_2180);
nor U2732 (N_2732,N_1834,N_2273);
nand U2733 (N_2733,N_2350,N_1974);
nor U2734 (N_2734,N_2280,N_1826);
or U2735 (N_2735,N_2092,N_2123);
and U2736 (N_2736,N_2367,N_2332);
nor U2737 (N_2737,N_2193,N_2170);
nor U2738 (N_2738,N_2315,N_2112);
nand U2739 (N_2739,N_2089,N_2137);
or U2740 (N_2740,N_2277,N_2068);
and U2741 (N_2741,N_1850,N_1829);
and U2742 (N_2742,N_1997,N_2169);
and U2743 (N_2743,N_2197,N_1802);
nand U2744 (N_2744,N_2332,N_2297);
or U2745 (N_2745,N_2048,N_2057);
and U2746 (N_2746,N_2070,N_1854);
or U2747 (N_2747,N_1998,N_2089);
or U2748 (N_2748,N_1809,N_2329);
nor U2749 (N_2749,N_1943,N_2309);
or U2750 (N_2750,N_2229,N_1997);
nor U2751 (N_2751,N_2050,N_2247);
nand U2752 (N_2752,N_2285,N_1910);
and U2753 (N_2753,N_2263,N_1896);
and U2754 (N_2754,N_2079,N_2356);
or U2755 (N_2755,N_2236,N_2308);
nand U2756 (N_2756,N_1963,N_2358);
nor U2757 (N_2757,N_1940,N_2383);
nor U2758 (N_2758,N_2190,N_2135);
nand U2759 (N_2759,N_1875,N_2089);
and U2760 (N_2760,N_2227,N_2079);
nor U2761 (N_2761,N_2348,N_2207);
nor U2762 (N_2762,N_1946,N_2146);
nor U2763 (N_2763,N_2113,N_2158);
and U2764 (N_2764,N_2385,N_2095);
or U2765 (N_2765,N_1931,N_1960);
or U2766 (N_2766,N_2199,N_2035);
nor U2767 (N_2767,N_2107,N_2002);
nor U2768 (N_2768,N_1994,N_1913);
or U2769 (N_2769,N_2152,N_2255);
or U2770 (N_2770,N_1974,N_2164);
nand U2771 (N_2771,N_2058,N_1960);
or U2772 (N_2772,N_1951,N_2246);
and U2773 (N_2773,N_1878,N_2147);
nand U2774 (N_2774,N_1819,N_2199);
nor U2775 (N_2775,N_2276,N_1886);
or U2776 (N_2776,N_2341,N_2073);
nand U2777 (N_2777,N_2005,N_1925);
nand U2778 (N_2778,N_2192,N_2023);
nand U2779 (N_2779,N_2315,N_1894);
and U2780 (N_2780,N_1929,N_1804);
nand U2781 (N_2781,N_2306,N_1889);
nor U2782 (N_2782,N_1809,N_2191);
nand U2783 (N_2783,N_2355,N_2392);
or U2784 (N_2784,N_1826,N_2231);
and U2785 (N_2785,N_2372,N_2143);
and U2786 (N_2786,N_2102,N_2377);
and U2787 (N_2787,N_1934,N_1915);
and U2788 (N_2788,N_2025,N_2289);
and U2789 (N_2789,N_1837,N_2049);
nor U2790 (N_2790,N_1902,N_2103);
or U2791 (N_2791,N_2365,N_2042);
nor U2792 (N_2792,N_2359,N_2206);
nor U2793 (N_2793,N_1847,N_2041);
nand U2794 (N_2794,N_1988,N_2303);
and U2795 (N_2795,N_2361,N_1936);
and U2796 (N_2796,N_2082,N_1839);
nand U2797 (N_2797,N_2212,N_2155);
or U2798 (N_2798,N_1866,N_2213);
nor U2799 (N_2799,N_2115,N_1842);
and U2800 (N_2800,N_2122,N_2229);
or U2801 (N_2801,N_2235,N_2017);
nand U2802 (N_2802,N_2007,N_2310);
nand U2803 (N_2803,N_2345,N_2185);
nand U2804 (N_2804,N_2214,N_2193);
nand U2805 (N_2805,N_2278,N_1870);
nor U2806 (N_2806,N_1879,N_2287);
or U2807 (N_2807,N_2345,N_2038);
nand U2808 (N_2808,N_2309,N_2090);
nor U2809 (N_2809,N_2201,N_2126);
or U2810 (N_2810,N_2004,N_2165);
and U2811 (N_2811,N_2377,N_1967);
and U2812 (N_2812,N_2204,N_2288);
and U2813 (N_2813,N_2079,N_2144);
nand U2814 (N_2814,N_1986,N_2057);
nor U2815 (N_2815,N_2309,N_2112);
and U2816 (N_2816,N_2124,N_2339);
nor U2817 (N_2817,N_2340,N_2372);
nand U2818 (N_2818,N_2380,N_2358);
nand U2819 (N_2819,N_2141,N_1900);
or U2820 (N_2820,N_2098,N_1868);
and U2821 (N_2821,N_2225,N_2081);
nor U2822 (N_2822,N_2140,N_2377);
and U2823 (N_2823,N_1971,N_1819);
nand U2824 (N_2824,N_2101,N_1825);
or U2825 (N_2825,N_2110,N_2133);
nor U2826 (N_2826,N_2031,N_1821);
and U2827 (N_2827,N_2090,N_2231);
nor U2828 (N_2828,N_1826,N_2381);
nor U2829 (N_2829,N_1912,N_2036);
or U2830 (N_2830,N_1884,N_1866);
nand U2831 (N_2831,N_2173,N_2344);
nor U2832 (N_2832,N_2097,N_2124);
and U2833 (N_2833,N_2154,N_2223);
nor U2834 (N_2834,N_2317,N_2356);
nor U2835 (N_2835,N_2112,N_1807);
nand U2836 (N_2836,N_2227,N_2312);
nand U2837 (N_2837,N_2150,N_1981);
and U2838 (N_2838,N_1890,N_2184);
nor U2839 (N_2839,N_2027,N_1936);
and U2840 (N_2840,N_2087,N_2118);
nor U2841 (N_2841,N_2125,N_2288);
and U2842 (N_2842,N_2375,N_2045);
nor U2843 (N_2843,N_1922,N_2098);
and U2844 (N_2844,N_1822,N_1972);
nor U2845 (N_2845,N_2054,N_2271);
nand U2846 (N_2846,N_2110,N_2196);
nor U2847 (N_2847,N_2240,N_2165);
nor U2848 (N_2848,N_2303,N_1938);
or U2849 (N_2849,N_2070,N_2004);
nand U2850 (N_2850,N_2346,N_2017);
nor U2851 (N_2851,N_2102,N_1842);
and U2852 (N_2852,N_2034,N_2272);
nand U2853 (N_2853,N_2244,N_2139);
nor U2854 (N_2854,N_2310,N_2376);
and U2855 (N_2855,N_2203,N_1957);
and U2856 (N_2856,N_2335,N_2322);
nor U2857 (N_2857,N_2011,N_1866);
nor U2858 (N_2858,N_2257,N_2167);
and U2859 (N_2859,N_1903,N_1890);
and U2860 (N_2860,N_1844,N_2072);
and U2861 (N_2861,N_1846,N_1909);
nor U2862 (N_2862,N_2162,N_2339);
nand U2863 (N_2863,N_2023,N_2306);
and U2864 (N_2864,N_1842,N_1881);
nor U2865 (N_2865,N_2341,N_2061);
and U2866 (N_2866,N_1814,N_1921);
and U2867 (N_2867,N_2337,N_2144);
and U2868 (N_2868,N_2084,N_2228);
nor U2869 (N_2869,N_1846,N_2075);
nand U2870 (N_2870,N_2154,N_2245);
nor U2871 (N_2871,N_1923,N_2287);
and U2872 (N_2872,N_1867,N_2375);
or U2873 (N_2873,N_2098,N_2101);
nand U2874 (N_2874,N_2288,N_1860);
or U2875 (N_2875,N_2076,N_1819);
or U2876 (N_2876,N_1934,N_2293);
and U2877 (N_2877,N_2139,N_1881);
nor U2878 (N_2878,N_2294,N_2323);
or U2879 (N_2879,N_2371,N_2383);
nand U2880 (N_2880,N_2191,N_2091);
nand U2881 (N_2881,N_2165,N_2017);
or U2882 (N_2882,N_2241,N_1938);
nand U2883 (N_2883,N_1886,N_2280);
or U2884 (N_2884,N_2020,N_2177);
nor U2885 (N_2885,N_1822,N_1956);
and U2886 (N_2886,N_2064,N_1918);
or U2887 (N_2887,N_2144,N_2148);
or U2888 (N_2888,N_2010,N_2337);
or U2889 (N_2889,N_1879,N_2282);
or U2890 (N_2890,N_1951,N_2084);
and U2891 (N_2891,N_1996,N_2299);
nor U2892 (N_2892,N_2048,N_1802);
nor U2893 (N_2893,N_2375,N_2271);
and U2894 (N_2894,N_1855,N_2359);
nor U2895 (N_2895,N_2320,N_2258);
or U2896 (N_2896,N_1958,N_2098);
nor U2897 (N_2897,N_2310,N_2397);
nor U2898 (N_2898,N_1836,N_1881);
or U2899 (N_2899,N_1928,N_2395);
nand U2900 (N_2900,N_1963,N_2097);
nand U2901 (N_2901,N_1989,N_2363);
or U2902 (N_2902,N_2151,N_1884);
or U2903 (N_2903,N_1965,N_1800);
nor U2904 (N_2904,N_2165,N_2117);
nand U2905 (N_2905,N_1841,N_2391);
nand U2906 (N_2906,N_2363,N_1881);
nor U2907 (N_2907,N_2293,N_2137);
or U2908 (N_2908,N_2241,N_2080);
and U2909 (N_2909,N_1960,N_2136);
and U2910 (N_2910,N_2167,N_2209);
and U2911 (N_2911,N_2083,N_2076);
nor U2912 (N_2912,N_2211,N_2014);
and U2913 (N_2913,N_2288,N_1921);
nor U2914 (N_2914,N_2320,N_2127);
nor U2915 (N_2915,N_1889,N_1921);
nor U2916 (N_2916,N_2157,N_2248);
and U2917 (N_2917,N_2034,N_2302);
or U2918 (N_2918,N_1976,N_1901);
or U2919 (N_2919,N_2058,N_2391);
nand U2920 (N_2920,N_2133,N_2323);
nor U2921 (N_2921,N_2301,N_2289);
nand U2922 (N_2922,N_2120,N_2282);
or U2923 (N_2923,N_2027,N_1875);
or U2924 (N_2924,N_2364,N_2310);
nor U2925 (N_2925,N_1926,N_1915);
or U2926 (N_2926,N_2084,N_2168);
and U2927 (N_2927,N_2267,N_2152);
and U2928 (N_2928,N_1972,N_2368);
or U2929 (N_2929,N_1932,N_2375);
and U2930 (N_2930,N_2023,N_2304);
nor U2931 (N_2931,N_1860,N_2108);
nor U2932 (N_2932,N_2164,N_2246);
xor U2933 (N_2933,N_2141,N_1973);
nand U2934 (N_2934,N_1995,N_2235);
or U2935 (N_2935,N_2104,N_2386);
and U2936 (N_2936,N_2075,N_2331);
and U2937 (N_2937,N_2338,N_2373);
and U2938 (N_2938,N_2348,N_2212);
nor U2939 (N_2939,N_2367,N_2149);
nand U2940 (N_2940,N_2353,N_2119);
and U2941 (N_2941,N_1971,N_1916);
or U2942 (N_2942,N_1823,N_2240);
nor U2943 (N_2943,N_2107,N_2273);
nand U2944 (N_2944,N_1817,N_2236);
nor U2945 (N_2945,N_2197,N_1967);
and U2946 (N_2946,N_2356,N_1831);
and U2947 (N_2947,N_1882,N_2316);
nand U2948 (N_2948,N_1894,N_1933);
or U2949 (N_2949,N_1917,N_2161);
nand U2950 (N_2950,N_2078,N_2213);
nor U2951 (N_2951,N_2156,N_2004);
nor U2952 (N_2952,N_2388,N_2367);
nor U2953 (N_2953,N_1949,N_2356);
nor U2954 (N_2954,N_1858,N_2309);
or U2955 (N_2955,N_1855,N_1818);
and U2956 (N_2956,N_2127,N_1896);
or U2957 (N_2957,N_1891,N_2357);
nand U2958 (N_2958,N_2207,N_2040);
nand U2959 (N_2959,N_2198,N_1974);
and U2960 (N_2960,N_2313,N_2283);
and U2961 (N_2961,N_2140,N_2270);
nor U2962 (N_2962,N_1938,N_2126);
and U2963 (N_2963,N_1893,N_2360);
or U2964 (N_2964,N_1967,N_2221);
or U2965 (N_2965,N_2066,N_2074);
or U2966 (N_2966,N_1915,N_2095);
or U2967 (N_2967,N_2192,N_1935);
or U2968 (N_2968,N_1976,N_2294);
or U2969 (N_2969,N_2091,N_2231);
nand U2970 (N_2970,N_1932,N_2111);
nand U2971 (N_2971,N_2076,N_1912);
nand U2972 (N_2972,N_2246,N_1897);
xor U2973 (N_2973,N_2155,N_1985);
nand U2974 (N_2974,N_2002,N_2388);
nor U2975 (N_2975,N_1847,N_2070);
and U2976 (N_2976,N_1978,N_2103);
and U2977 (N_2977,N_2267,N_2342);
or U2978 (N_2978,N_2330,N_1848);
and U2979 (N_2979,N_1900,N_2109);
nand U2980 (N_2980,N_1854,N_2119);
nand U2981 (N_2981,N_2031,N_2021);
nor U2982 (N_2982,N_2296,N_2272);
or U2983 (N_2983,N_1875,N_2334);
or U2984 (N_2984,N_2040,N_2250);
nand U2985 (N_2985,N_2168,N_1919);
nand U2986 (N_2986,N_2380,N_2063);
or U2987 (N_2987,N_1993,N_1860);
nor U2988 (N_2988,N_2233,N_1989);
or U2989 (N_2989,N_2237,N_1966);
and U2990 (N_2990,N_1964,N_2008);
nor U2991 (N_2991,N_2369,N_2031);
nand U2992 (N_2992,N_2380,N_2121);
nor U2993 (N_2993,N_1992,N_1802);
or U2994 (N_2994,N_1840,N_1837);
and U2995 (N_2995,N_1898,N_2330);
and U2996 (N_2996,N_2049,N_2242);
or U2997 (N_2997,N_2171,N_2096);
or U2998 (N_2998,N_1895,N_2325);
nand U2999 (N_2999,N_2132,N_2138);
nand UO_0 (O_0,N_2729,N_2786);
nor UO_1 (O_1,N_2495,N_2583);
or UO_2 (O_2,N_2715,N_2687);
nand UO_3 (O_3,N_2817,N_2820);
nand UO_4 (O_4,N_2695,N_2730);
and UO_5 (O_5,N_2949,N_2487);
nand UO_6 (O_6,N_2684,N_2449);
nand UO_7 (O_7,N_2823,N_2785);
nor UO_8 (O_8,N_2677,N_2604);
nand UO_9 (O_9,N_2904,N_2746);
and UO_10 (O_10,N_2435,N_2411);
and UO_11 (O_11,N_2948,N_2995);
and UO_12 (O_12,N_2711,N_2963);
nor UO_13 (O_13,N_2889,N_2906);
nand UO_14 (O_14,N_2469,N_2734);
and UO_15 (O_15,N_2626,N_2918);
nor UO_16 (O_16,N_2722,N_2550);
nand UO_17 (O_17,N_2477,N_2890);
nand UO_18 (O_18,N_2821,N_2508);
or UO_19 (O_19,N_2713,N_2969);
and UO_20 (O_20,N_2933,N_2965);
or UO_21 (O_21,N_2700,N_2919);
or UO_22 (O_22,N_2607,N_2901);
and UO_23 (O_23,N_2825,N_2659);
nor UO_24 (O_24,N_2418,N_2610);
nor UO_25 (O_25,N_2750,N_2405);
or UO_26 (O_26,N_2404,N_2406);
and UO_27 (O_27,N_2788,N_2598);
and UO_28 (O_28,N_2689,N_2675);
nor UO_29 (O_29,N_2651,N_2408);
or UO_30 (O_30,N_2455,N_2961);
nand UO_31 (O_31,N_2784,N_2649);
nor UO_32 (O_32,N_2420,N_2619);
nand UO_33 (O_33,N_2543,N_2736);
nand UO_34 (O_34,N_2478,N_2662);
or UO_35 (O_35,N_2917,N_2803);
nor UO_36 (O_36,N_2433,N_2895);
and UO_37 (O_37,N_2735,N_2453);
nand UO_38 (O_38,N_2849,N_2454);
nand UO_39 (O_39,N_2505,N_2674);
nor UO_40 (O_40,N_2991,N_2912);
and UO_41 (O_41,N_2526,N_2605);
and UO_42 (O_42,N_2412,N_2828);
nand UO_43 (O_43,N_2745,N_2533);
nor UO_44 (O_44,N_2499,N_2813);
or UO_45 (O_45,N_2769,N_2504);
nand UO_46 (O_46,N_2593,N_2458);
or UO_47 (O_47,N_2709,N_2488);
nand UO_48 (O_48,N_2515,N_2576);
nand UO_49 (O_49,N_2613,N_2642);
nor UO_50 (O_50,N_2587,N_2512);
nand UO_51 (O_51,N_2548,N_2987);
nand UO_52 (O_52,N_2692,N_2871);
nor UO_53 (O_53,N_2671,N_2721);
nand UO_54 (O_54,N_2500,N_2908);
or UO_55 (O_55,N_2596,N_2847);
nor UO_56 (O_56,N_2400,N_2774);
or UO_57 (O_57,N_2936,N_2880);
or UO_58 (O_58,N_2441,N_2926);
and UO_59 (O_59,N_2415,N_2579);
nand UO_60 (O_60,N_2968,N_2795);
or UO_61 (O_61,N_2629,N_2916);
nand UO_62 (O_62,N_2616,N_2957);
and UO_63 (O_63,N_2754,N_2898);
and UO_64 (O_64,N_2866,N_2799);
and UO_65 (O_65,N_2717,N_2907);
nand UO_66 (O_66,N_2472,N_2693);
nand UO_67 (O_67,N_2718,N_2812);
nand UO_68 (O_68,N_2814,N_2585);
and UO_69 (O_69,N_2768,N_2492);
nand UO_70 (O_70,N_2705,N_2489);
nand UO_71 (O_71,N_2570,N_2402);
nand UO_72 (O_72,N_2545,N_2482);
or UO_73 (O_73,N_2714,N_2666);
nand UO_74 (O_74,N_2846,N_2839);
nand UO_75 (O_75,N_2572,N_2737);
nand UO_76 (O_76,N_2416,N_2470);
or UO_77 (O_77,N_2690,N_2959);
and UO_78 (O_78,N_2831,N_2698);
or UO_79 (O_79,N_2796,N_2565);
nor UO_80 (O_80,N_2474,N_2502);
and UO_81 (O_81,N_2511,N_2858);
and UO_82 (O_82,N_2595,N_2801);
nand UO_83 (O_83,N_2955,N_2970);
or UO_84 (O_84,N_2909,N_2465);
nand UO_85 (O_85,N_2497,N_2951);
nor UO_86 (O_86,N_2944,N_2932);
nor UO_87 (O_87,N_2707,N_2620);
nand UO_88 (O_88,N_2724,N_2732);
nand UO_89 (O_89,N_2553,N_2637);
and UO_90 (O_90,N_2998,N_2892);
nand UO_91 (O_91,N_2410,N_2804);
nor UO_92 (O_92,N_2872,N_2423);
or UO_93 (O_93,N_2845,N_2432);
and UO_94 (O_94,N_2964,N_2694);
and UO_95 (O_95,N_2986,N_2602);
or UO_96 (O_96,N_2556,N_2836);
or UO_97 (O_97,N_2739,N_2439);
nor UO_98 (O_98,N_2878,N_2855);
and UO_99 (O_99,N_2528,N_2688);
or UO_100 (O_100,N_2771,N_2573);
nand UO_101 (O_101,N_2843,N_2481);
or UO_102 (O_102,N_2925,N_2857);
nand UO_103 (O_103,N_2468,N_2905);
and UO_104 (O_104,N_2635,N_2877);
or UO_105 (O_105,N_2952,N_2655);
nand UO_106 (O_106,N_2600,N_2685);
and UO_107 (O_107,N_2757,N_2874);
and UO_108 (O_108,N_2856,N_2865);
nor UO_109 (O_109,N_2879,N_2514);
nor UO_110 (O_110,N_2743,N_2679);
and UO_111 (O_111,N_2947,N_2853);
or UO_112 (O_112,N_2984,N_2575);
and UO_113 (O_113,N_2456,N_2440);
and UO_114 (O_114,N_2424,N_2638);
nor UO_115 (O_115,N_2676,N_2726);
or UO_116 (O_116,N_2485,N_2922);
nand UO_117 (O_117,N_2574,N_2623);
xnor UO_118 (O_118,N_2667,N_2555);
nand UO_119 (O_119,N_2954,N_2973);
nor UO_120 (O_120,N_2431,N_2444);
or UO_121 (O_121,N_2884,N_2633);
or UO_122 (O_122,N_2793,N_2434);
xor UO_123 (O_123,N_2840,N_2988);
nand UO_124 (O_124,N_2997,N_2826);
or UO_125 (O_125,N_2731,N_2939);
and UO_126 (O_126,N_2742,N_2805);
nand UO_127 (O_127,N_2603,N_2807);
nor UO_128 (O_128,N_2464,N_2930);
nand UO_129 (O_129,N_2467,N_2775);
or UO_130 (O_130,N_2490,N_2868);
or UO_131 (O_131,N_2582,N_2566);
nand UO_132 (O_132,N_2647,N_2752);
and UO_133 (O_133,N_2535,N_2463);
or UO_134 (O_134,N_2850,N_2680);
nor UO_135 (O_135,N_2762,N_2891);
nor UO_136 (O_136,N_2888,N_2744);
or UO_137 (O_137,N_2668,N_2830);
or UO_138 (O_138,N_2966,N_2903);
or UO_139 (O_139,N_2521,N_2989);
and UO_140 (O_140,N_2990,N_2696);
and UO_141 (O_141,N_2981,N_2563);
nor UO_142 (O_142,N_2741,N_2802);
nand UO_143 (O_143,N_2864,N_2445);
nor UO_144 (O_144,N_2429,N_2837);
nand UO_145 (O_145,N_2417,N_2660);
nor UO_146 (O_146,N_2584,N_2827);
nor UO_147 (O_147,N_2834,N_2720);
nor UO_148 (O_148,N_2921,N_2529);
or UO_149 (O_149,N_2627,N_2710);
nand UO_150 (O_150,N_2524,N_2756);
or UO_151 (O_151,N_2539,N_2806);
and UO_152 (O_152,N_2648,N_2728);
and UO_153 (O_153,N_2611,N_2641);
and UO_154 (O_154,N_2992,N_2471);
nand UO_155 (O_155,N_2451,N_2622);
nor UO_156 (O_156,N_2751,N_2764);
or UO_157 (O_157,N_2829,N_2683);
nor UO_158 (O_158,N_2686,N_2789);
nand UO_159 (O_159,N_2776,N_2540);
nor UO_160 (O_160,N_2670,N_2673);
and UO_161 (O_161,N_2938,N_2935);
and UO_162 (O_162,N_2763,N_2994);
or UO_163 (O_163,N_2578,N_2971);
and UO_164 (O_164,N_2755,N_2811);
and UO_165 (O_165,N_2422,N_2483);
and UO_166 (O_166,N_2665,N_2496);
nor UO_167 (O_167,N_2716,N_2897);
or UO_168 (O_168,N_2953,N_2977);
nand UO_169 (O_169,N_2401,N_2428);
nor UO_170 (O_170,N_2522,N_2893);
nand UO_171 (O_171,N_2541,N_2982);
nand UO_172 (O_172,N_2597,N_2887);
or UO_173 (O_173,N_2546,N_2929);
nor UO_174 (O_174,N_2854,N_2958);
nor UO_175 (O_175,N_2475,N_2656);
or UO_176 (O_176,N_2749,N_2559);
nor UO_177 (O_177,N_2975,N_2479);
nor UO_178 (O_178,N_2661,N_2915);
and UO_179 (O_179,N_2523,N_2513);
nand UO_180 (O_180,N_2436,N_2851);
nor UO_181 (O_181,N_2678,N_2885);
or UO_182 (O_182,N_2614,N_2819);
and UO_183 (O_183,N_2520,N_2810);
or UO_184 (O_184,N_2733,N_2427);
and UO_185 (O_185,N_2704,N_2748);
or UO_186 (O_186,N_2443,N_2608);
and UO_187 (O_187,N_2738,N_2446);
nand UO_188 (O_188,N_2924,N_2530);
nand UO_189 (O_189,N_2900,N_2760);
or UO_190 (O_190,N_2910,N_2480);
and UO_191 (O_191,N_2913,N_2657);
nor UO_192 (O_192,N_2873,N_2999);
or UO_193 (O_193,N_2654,N_2632);
and UO_194 (O_194,N_2727,N_2624);
and UO_195 (O_195,N_2599,N_2549);
nor UO_196 (O_196,N_2646,N_2979);
nand UO_197 (O_197,N_2934,N_2527);
nand UO_198 (O_198,N_2794,N_2822);
and UO_199 (O_199,N_2740,N_2972);
and UO_200 (O_200,N_2409,N_2896);
or UO_201 (O_201,N_2486,N_2706);
nand UO_202 (O_202,N_2532,N_2590);
and UO_203 (O_203,N_2773,N_2708);
nand UO_204 (O_204,N_2510,N_2815);
nand UO_205 (O_205,N_2702,N_2476);
and UO_206 (O_206,N_2554,N_2861);
and UO_207 (O_207,N_2838,N_2691);
and UO_208 (O_208,N_2452,N_2517);
or UO_209 (O_209,N_2937,N_2859);
nor UO_210 (O_210,N_2832,N_2960);
nor UO_211 (O_211,N_2460,N_2493);
nor UO_212 (O_212,N_2983,N_2403);
nor UO_213 (O_213,N_2644,N_2701);
nand UO_214 (O_214,N_2664,N_2766);
nand UO_215 (O_215,N_2594,N_2609);
or UO_216 (O_216,N_2869,N_2437);
nor UO_217 (O_217,N_2781,N_2945);
and UO_218 (O_218,N_2920,N_2703);
nor UO_219 (O_219,N_2636,N_2419);
or UO_220 (O_220,N_2580,N_2426);
and UO_221 (O_221,N_2931,N_2894);
or UO_222 (O_222,N_2669,N_2881);
and UO_223 (O_223,N_2902,N_2797);
nand UO_224 (O_224,N_2777,N_2615);
nand UO_225 (O_225,N_2501,N_2645);
or UO_226 (O_226,N_2509,N_2658);
nand UO_227 (O_227,N_2985,N_2765);
and UO_228 (O_228,N_2719,N_2899);
or UO_229 (O_229,N_2833,N_2816);
nor UO_230 (O_230,N_2564,N_2980);
or UO_231 (O_231,N_2519,N_2413);
nand UO_232 (O_232,N_2558,N_2653);
nand UO_233 (O_233,N_2942,N_2557);
nor UO_234 (O_234,N_2844,N_2652);
and UO_235 (O_235,N_2650,N_2459);
nand UO_236 (O_236,N_2425,N_2551);
nor UO_237 (O_237,N_2568,N_2798);
nand UO_238 (O_238,N_2473,N_2448);
and UO_239 (O_239,N_2941,N_2770);
or UO_240 (O_240,N_2438,N_2630);
and UO_241 (O_241,N_2699,N_2824);
nand UO_242 (O_242,N_2631,N_2450);
nand UO_243 (O_243,N_2561,N_2612);
nand UO_244 (O_244,N_2852,N_2466);
or UO_245 (O_245,N_2787,N_2606);
nor UO_246 (O_246,N_2976,N_2886);
nor UO_247 (O_247,N_2634,N_2946);
nor UO_248 (O_248,N_2639,N_2753);
nor UO_249 (O_249,N_2967,N_2870);
nor UO_250 (O_250,N_2457,N_2531);
nor UO_251 (O_251,N_2491,N_2876);
nand UO_252 (O_252,N_2462,N_2536);
nand UO_253 (O_253,N_2552,N_2996);
or UO_254 (O_254,N_2911,N_2712);
or UO_255 (O_255,N_2544,N_2862);
nand UO_256 (O_256,N_2682,N_2442);
and UO_257 (O_257,N_2841,N_2978);
nor UO_258 (O_258,N_2414,N_2498);
or UO_259 (O_259,N_2778,N_2974);
nand UO_260 (O_260,N_2503,N_2618);
nor UO_261 (O_261,N_2581,N_2484);
nand UO_262 (O_262,N_2791,N_2525);
nand UO_263 (O_263,N_2421,N_2621);
nor UO_264 (O_264,N_2625,N_2617);
or UO_265 (O_265,N_2928,N_2681);
nand UO_266 (O_266,N_2993,N_2534);
or UO_267 (O_267,N_2914,N_2672);
and UO_268 (O_268,N_2790,N_2560);
nand UO_269 (O_269,N_2940,N_2780);
or UO_270 (O_270,N_2537,N_2842);
and UO_271 (O_271,N_2407,N_2950);
nand UO_272 (O_272,N_2507,N_2882);
or UO_273 (O_273,N_2818,N_2808);
and UO_274 (O_274,N_2835,N_2863);
nand UO_275 (O_275,N_2779,N_2860);
nor UO_276 (O_276,N_2589,N_2923);
nand UO_277 (O_277,N_2758,N_2591);
nand UO_278 (O_278,N_2640,N_2759);
nand UO_279 (O_279,N_2516,N_2725);
nand UO_280 (O_280,N_2783,N_2956);
or UO_281 (O_281,N_2697,N_2506);
or UO_282 (O_282,N_2761,N_2577);
nand UO_283 (O_283,N_2943,N_2800);
and UO_284 (O_284,N_2547,N_2430);
nand UO_285 (O_285,N_2848,N_2447);
or UO_286 (O_286,N_2588,N_2518);
nor UO_287 (O_287,N_2571,N_2628);
or UO_288 (O_288,N_2586,N_2782);
and UO_289 (O_289,N_2962,N_2592);
nand UO_290 (O_290,N_2867,N_2747);
nand UO_291 (O_291,N_2461,N_2883);
or UO_292 (O_292,N_2875,N_2792);
nand UO_293 (O_293,N_2927,N_2643);
and UO_294 (O_294,N_2542,N_2772);
nand UO_295 (O_295,N_2567,N_2569);
and UO_296 (O_296,N_2809,N_2494);
nand UO_297 (O_297,N_2663,N_2562);
and UO_298 (O_298,N_2601,N_2767);
or UO_299 (O_299,N_2538,N_2723);
nor UO_300 (O_300,N_2954,N_2505);
or UO_301 (O_301,N_2563,N_2707);
or UO_302 (O_302,N_2970,N_2632);
nand UO_303 (O_303,N_2424,N_2581);
nor UO_304 (O_304,N_2427,N_2831);
nand UO_305 (O_305,N_2611,N_2422);
nor UO_306 (O_306,N_2517,N_2964);
nand UO_307 (O_307,N_2845,N_2997);
nor UO_308 (O_308,N_2672,N_2524);
xnor UO_309 (O_309,N_2710,N_2495);
or UO_310 (O_310,N_2547,N_2721);
nand UO_311 (O_311,N_2414,N_2578);
and UO_312 (O_312,N_2644,N_2583);
nor UO_313 (O_313,N_2807,N_2642);
and UO_314 (O_314,N_2431,N_2741);
nor UO_315 (O_315,N_2996,N_2853);
nand UO_316 (O_316,N_2722,N_2980);
nand UO_317 (O_317,N_2866,N_2785);
nor UO_318 (O_318,N_2818,N_2709);
and UO_319 (O_319,N_2516,N_2747);
nand UO_320 (O_320,N_2646,N_2756);
or UO_321 (O_321,N_2933,N_2560);
nor UO_322 (O_322,N_2644,N_2627);
nor UO_323 (O_323,N_2853,N_2456);
nand UO_324 (O_324,N_2713,N_2670);
nand UO_325 (O_325,N_2841,N_2890);
nor UO_326 (O_326,N_2662,N_2911);
or UO_327 (O_327,N_2644,N_2408);
nor UO_328 (O_328,N_2851,N_2452);
or UO_329 (O_329,N_2861,N_2806);
nand UO_330 (O_330,N_2664,N_2486);
or UO_331 (O_331,N_2709,N_2727);
and UO_332 (O_332,N_2886,N_2493);
nor UO_333 (O_333,N_2701,N_2793);
nor UO_334 (O_334,N_2790,N_2458);
and UO_335 (O_335,N_2587,N_2758);
nor UO_336 (O_336,N_2450,N_2632);
nand UO_337 (O_337,N_2798,N_2795);
or UO_338 (O_338,N_2497,N_2918);
nor UO_339 (O_339,N_2652,N_2803);
and UO_340 (O_340,N_2822,N_2636);
or UO_341 (O_341,N_2431,N_2410);
and UO_342 (O_342,N_2919,N_2773);
or UO_343 (O_343,N_2682,N_2654);
or UO_344 (O_344,N_2457,N_2405);
nand UO_345 (O_345,N_2941,N_2680);
nand UO_346 (O_346,N_2969,N_2702);
nor UO_347 (O_347,N_2534,N_2838);
and UO_348 (O_348,N_2714,N_2554);
nand UO_349 (O_349,N_2755,N_2729);
and UO_350 (O_350,N_2747,N_2498);
nor UO_351 (O_351,N_2691,N_2546);
nand UO_352 (O_352,N_2760,N_2543);
nand UO_353 (O_353,N_2590,N_2534);
or UO_354 (O_354,N_2470,N_2778);
or UO_355 (O_355,N_2414,N_2477);
or UO_356 (O_356,N_2635,N_2955);
or UO_357 (O_357,N_2796,N_2756);
nor UO_358 (O_358,N_2427,N_2852);
and UO_359 (O_359,N_2874,N_2413);
nand UO_360 (O_360,N_2487,N_2929);
or UO_361 (O_361,N_2430,N_2768);
nand UO_362 (O_362,N_2660,N_2976);
and UO_363 (O_363,N_2463,N_2466);
xor UO_364 (O_364,N_2606,N_2572);
nor UO_365 (O_365,N_2719,N_2736);
nor UO_366 (O_366,N_2590,N_2610);
or UO_367 (O_367,N_2400,N_2449);
nor UO_368 (O_368,N_2945,N_2618);
and UO_369 (O_369,N_2528,N_2917);
nand UO_370 (O_370,N_2571,N_2753);
or UO_371 (O_371,N_2431,N_2873);
nand UO_372 (O_372,N_2841,N_2815);
and UO_373 (O_373,N_2890,N_2753);
nor UO_374 (O_374,N_2406,N_2697);
or UO_375 (O_375,N_2778,N_2615);
nor UO_376 (O_376,N_2758,N_2563);
nor UO_377 (O_377,N_2710,N_2536);
nand UO_378 (O_378,N_2673,N_2518);
and UO_379 (O_379,N_2835,N_2630);
nor UO_380 (O_380,N_2834,N_2864);
nor UO_381 (O_381,N_2546,N_2945);
or UO_382 (O_382,N_2650,N_2861);
nor UO_383 (O_383,N_2934,N_2925);
and UO_384 (O_384,N_2427,N_2874);
nand UO_385 (O_385,N_2917,N_2881);
nand UO_386 (O_386,N_2973,N_2509);
nor UO_387 (O_387,N_2406,N_2482);
nand UO_388 (O_388,N_2810,N_2780);
nor UO_389 (O_389,N_2961,N_2539);
or UO_390 (O_390,N_2793,N_2517);
or UO_391 (O_391,N_2579,N_2864);
xnor UO_392 (O_392,N_2739,N_2670);
nand UO_393 (O_393,N_2493,N_2807);
nor UO_394 (O_394,N_2487,N_2768);
and UO_395 (O_395,N_2894,N_2786);
nor UO_396 (O_396,N_2706,N_2729);
nor UO_397 (O_397,N_2821,N_2704);
nor UO_398 (O_398,N_2469,N_2400);
or UO_399 (O_399,N_2985,N_2869);
or UO_400 (O_400,N_2873,N_2488);
or UO_401 (O_401,N_2482,N_2461);
and UO_402 (O_402,N_2638,N_2944);
nand UO_403 (O_403,N_2498,N_2830);
and UO_404 (O_404,N_2560,N_2500);
or UO_405 (O_405,N_2595,N_2696);
or UO_406 (O_406,N_2556,N_2424);
nand UO_407 (O_407,N_2712,N_2599);
and UO_408 (O_408,N_2505,N_2970);
nand UO_409 (O_409,N_2413,N_2992);
nand UO_410 (O_410,N_2868,N_2791);
and UO_411 (O_411,N_2608,N_2796);
or UO_412 (O_412,N_2615,N_2752);
nand UO_413 (O_413,N_2625,N_2682);
xnor UO_414 (O_414,N_2848,N_2661);
and UO_415 (O_415,N_2673,N_2540);
nand UO_416 (O_416,N_2890,N_2750);
or UO_417 (O_417,N_2526,N_2554);
nor UO_418 (O_418,N_2868,N_2480);
nand UO_419 (O_419,N_2523,N_2738);
or UO_420 (O_420,N_2679,N_2767);
and UO_421 (O_421,N_2538,N_2925);
or UO_422 (O_422,N_2621,N_2914);
and UO_423 (O_423,N_2836,N_2589);
and UO_424 (O_424,N_2675,N_2651);
nand UO_425 (O_425,N_2652,N_2805);
nor UO_426 (O_426,N_2499,N_2629);
and UO_427 (O_427,N_2730,N_2493);
nor UO_428 (O_428,N_2898,N_2456);
nor UO_429 (O_429,N_2864,N_2724);
or UO_430 (O_430,N_2687,N_2714);
nand UO_431 (O_431,N_2482,N_2502);
nor UO_432 (O_432,N_2461,N_2622);
nor UO_433 (O_433,N_2500,N_2574);
nand UO_434 (O_434,N_2959,N_2696);
nand UO_435 (O_435,N_2525,N_2627);
nor UO_436 (O_436,N_2824,N_2558);
or UO_437 (O_437,N_2459,N_2686);
nor UO_438 (O_438,N_2508,N_2953);
nor UO_439 (O_439,N_2504,N_2519);
or UO_440 (O_440,N_2505,N_2873);
nor UO_441 (O_441,N_2815,N_2432);
or UO_442 (O_442,N_2795,N_2581);
and UO_443 (O_443,N_2937,N_2680);
nor UO_444 (O_444,N_2911,N_2892);
nand UO_445 (O_445,N_2503,N_2409);
nor UO_446 (O_446,N_2421,N_2634);
and UO_447 (O_447,N_2957,N_2736);
nand UO_448 (O_448,N_2622,N_2636);
or UO_449 (O_449,N_2437,N_2452);
and UO_450 (O_450,N_2705,N_2902);
nand UO_451 (O_451,N_2557,N_2675);
nor UO_452 (O_452,N_2802,N_2682);
or UO_453 (O_453,N_2403,N_2424);
nor UO_454 (O_454,N_2525,N_2646);
or UO_455 (O_455,N_2907,N_2960);
xor UO_456 (O_456,N_2794,N_2742);
nand UO_457 (O_457,N_2410,N_2553);
nor UO_458 (O_458,N_2678,N_2947);
nand UO_459 (O_459,N_2559,N_2866);
or UO_460 (O_460,N_2464,N_2814);
or UO_461 (O_461,N_2662,N_2872);
nand UO_462 (O_462,N_2477,N_2693);
nand UO_463 (O_463,N_2805,N_2967);
nor UO_464 (O_464,N_2548,N_2704);
or UO_465 (O_465,N_2415,N_2938);
and UO_466 (O_466,N_2995,N_2568);
and UO_467 (O_467,N_2983,N_2468);
nand UO_468 (O_468,N_2557,N_2673);
nor UO_469 (O_469,N_2913,N_2771);
and UO_470 (O_470,N_2547,N_2820);
nand UO_471 (O_471,N_2985,N_2796);
or UO_472 (O_472,N_2408,N_2631);
nand UO_473 (O_473,N_2479,N_2832);
or UO_474 (O_474,N_2617,N_2453);
or UO_475 (O_475,N_2662,N_2611);
and UO_476 (O_476,N_2975,N_2770);
nor UO_477 (O_477,N_2478,N_2853);
or UO_478 (O_478,N_2727,N_2682);
or UO_479 (O_479,N_2672,N_2570);
nor UO_480 (O_480,N_2893,N_2490);
and UO_481 (O_481,N_2666,N_2718);
nand UO_482 (O_482,N_2736,N_2927);
and UO_483 (O_483,N_2677,N_2826);
nor UO_484 (O_484,N_2949,N_2638);
or UO_485 (O_485,N_2709,N_2514);
and UO_486 (O_486,N_2599,N_2967);
nand UO_487 (O_487,N_2856,N_2439);
nand UO_488 (O_488,N_2410,N_2500);
and UO_489 (O_489,N_2417,N_2420);
and UO_490 (O_490,N_2837,N_2545);
nand UO_491 (O_491,N_2531,N_2429);
nor UO_492 (O_492,N_2516,N_2565);
or UO_493 (O_493,N_2454,N_2561);
or UO_494 (O_494,N_2631,N_2569);
and UO_495 (O_495,N_2927,N_2954);
nor UO_496 (O_496,N_2925,N_2747);
nor UO_497 (O_497,N_2781,N_2670);
nor UO_498 (O_498,N_2694,N_2575);
nor UO_499 (O_499,N_2918,N_2657);
endmodule